module top( n18 , n25 , n30 , n67 , n68 , n101 , n103 , n126 , n146 , 
n152 , n180 , n204 , n240 , n250 , n269 , n297 , n306 , n327 , n345 , 
n362 , n369 , n420 , n426 , n432 , n465 , n467 , n485 , n495 , n500 , 
n505 , n529 , n548 , n584 , n587 , n589 , n594 , n607 , n618 , n628 , 
n657 , n663 , n687 , n692 , n696 , n698 , n705 , n747 , n755 , n760 , 
n777 , n792 , n796 , n803 , n824 , n837 , n861 , n864 , n873 , n882 , 
n943 , n1016 , n1017 , n1024 , n1048 , n1052 , n1086 , n1091 , n1151 , n1168 , 
n1201 , n1208 , n1216 , n1218 , n1219 , n1220 , n1255 , n1317 , n1341 , n1381 , 
n1404 , n1413 , n1421 , n1432 , n1435 , n1443 , n1471 , n1486 , n1501 , n1512 , 
n1621 , n1654 , n1660 , n1690 , n1714 , n1760 , n1774 , n1779 , n1794 , n1803 , 
n1808 , n1813 , n1820 , n1839 , n1857 , n1860 , n1861 , n1888 , n1903 , n1905 , 
n1942 , n1958 , n1971 , n1972 , n1999 , n2004 , n2022 , n2023 , n2027 , n2093 , 
n2132 , n2142 , n2146 , n2171 , n2247 , n2262 , n2289 , n2301 , n2302 , n2318 , 
n2336 , n2419 , n2436 , n2439 , n2440 , n2511 , n2534 , n2551 , n2554 , n2563 , 
n2577 , n2598 , n2631 , n2638 , n2641 , n2714 , n2716 , n2744 , n2774 , n2804 , 
n2821 , n2836 , n2840 , n2841 , n2856 , n2884 , n2988 , n2993 , n3001 , n3030 , 
n3037 , n3053 , n3061 , n3070 , n3077 , n3084 , n3089 , n3090 , n3140 , n3164 , 
n3174 , n3245 , n3282 , n3283 , n3349 , n3360 , n3385 , n3412 , n3421 , n3430 , 
n3451 , n3455 , n3470 , n3489 , n3496 , n3519 , n3542 , n3573 , n3577 , n3587 , 
n3609 , n3626 , n3644 , n3656 , n3657 , n3681 , n3687 , n3690 , n3711 , n3717 , 
n3723 , n3728 , n3757 , n3761 , n3829 , n3892 , n3911 , n3923 , n3949 , n3955 , 
n3969 , n3982 , n3993 , n4028 , n4043 , n4049 , n4050 , n4058 , n4079 , n4098 , 
n4100 , n4114 , n4119 , n4142 , n4164 , n4168 , n4192 , n4223 , n4231 , n4237 , 
n4274 , n4303 , n4319 , n4331 , n4332 , n4336 , n4338 , n4339 , n4346 , n4347 , 
n4349 , n4353 , n4365 , n4370 , n4403 , n4410 , n4425 , n4432 , n4448 , n4451 , 
n4454 , n4467 , n4495 , n4544 , n4562 , n4575 , n4584 , n4599 , n4604 , n4615 , 
n4690 , n4702 , n4706 , n4720 , n4723 , n4735 , n4743 , n4762 , n4771 , n4777 , 
n4783 , n4799 , n4800 , n4805 , n4823 , n4826 , n4833 , n4860 , n4866 , n4875 , 
n4884 , n4888 , n4895 , n4904 , n4922 , n4925 , n4937 , n4940 , n4972 , n4991 , 
n4996 , n5007 , n5031 , n5038 , n5098 , n5102 , n5106 , n5127 , n5177 , n5190 , 
n5205 , n5233 , n5248 , n5251 , n5252 , n5258 , n5277 , n5314 , n5326 , n5333 , 
n5334 , n5363 , n5394 , n5401 , n5402 , n5426 , n5447 , n5450 , n5456 , n5490 , 
n5506 , n5509 , n5511 , n5519 , n5520 , n5521 , n5535 , n5547 , n5557 , n5567 , 
n5602 , n5624 , n5638 , n5639 , n5647 , n5654 , n5662 , n5664 , n5670 , n5717 , 
n5743 , n5774 , n5792 , n5804 , n5829 , n5848 , n5852 , n5857 , n5871 , n5883 , 
n5901 , n5902 , n5906 , n5907 , n5934 , n5954 , n5992 , n5995 , n6017 , n6025 , 
n6034 , n6038 , n6052 , n6053 , n6076 , n6128 , n6134 , n6154 , n6175 , n6187 , 
n6241 , n6282 , n6287 , n6291 );
    input n18 , n25 , n30 , n101 , n103 , n126 , n146 , n152 , n180 , 
n240 , n297 , n327 , n345 , n369 , n426 , n432 , n495 , n500 , n505 , 
n529 , n548 , n587 , n594 , n618 , n628 , n657 , n687 , n692 , n696 , 
n747 , n755 , n760 , n777 , n792 , n796 , n824 , n837 , n861 , n864 , 
n873 , n882 , n943 , n1016 , n1048 , n1052 , n1091 , n1151 , n1201 , n1216 , 
n1218 , n1220 , n1255 , n1381 , n1413 , n1432 , n1443 , n1471 , n1501 , n1512 , 
n1621 , n1654 , n1690 , n1714 , n1760 , n1774 , n1808 , n1813 , n1820 , n1861 , 
n1888 , n1903 , n1905 , n1942 , n1958 , n1971 , n1972 , n1999 , n2004 , n2022 , 
n2027 , n2093 , n2132 , n2142 , n2146 , n2247 , n2262 , n2289 , n2301 , n2318 , 
n2336 , n2419 , n2436 , n2440 , n2534 , n2551 , n2554 , n2563 , n2577 , n2638 , 
n2714 , n2744 , n2804 , n2836 , n2840 , n2841 , n2884 , n2988 , n2993 , n3001 , 
n3030 , n3037 , n3053 , n3061 , n3077 , n3084 , n3089 , n3140 , n3164 , n3174 , 
n3349 , n3360 , n3421 , n3451 , n3489 , n3519 , n3542 , n3573 , n3577 , n3644 , 
n3681 , n3687 , n3690 , n3717 , n3723 , n3728 , n3761 , n3829 , n3911 , n3955 , 
n3969 , n3993 , n4028 , n4043 , n4049 , n4050 , n4058 , n4098 , n4100 , n4119 , 
n4142 , n4164 , n4168 , n4231 , n4303 , n4319 , n4331 , n4332 , n4336 , n4338 , 
n4339 , n4346 , n4347 , n4353 , n4365 , n4370 , n4403 , n4425 , n4432 , n4448 , 
n4451 , n4454 , n4467 , n4495 , n4562 , n4575 , n4584 , n4599 , n4604 , n4615 , 
n4720 , n4723 , n4735 , n4743 , n4771 , n4777 , n4805 , n4823 , n4833 , n4866 , 
n4888 , n4922 , n4925 , n4937 , n4940 , n5031 , n5102 , n5106 , n5127 , n5177 , 
n5190 , n5205 , n5233 , n5248 , n5252 , n5258 , n5277 , n5314 , n5333 , n5363 , 
n5426 , n5450 , n5490 , n5506 , n5519 , n5521 , n5557 , n5602 , n5624 , n5638 , 
n5654 , n5662 , n5670 , n5717 , n5792 , n5829 , n5848 , n5852 , n5857 , n5883 , 
n5901 , n5906 , n5907 , n5992 , n5995 , n6017 , n6034 , n6038 , n6052 , n6053 , 
n6128 , n6154 , n6175 , n6241 , n6282 ;
    output n67 , n68 , n204 , n250 , n269 , n306 , n362 , n420 , n465 , 
n467 , n485 , n584 , n589 , n607 , n663 , n698 , n705 , n803 , n1017 , 
n1024 , n1086 , n1168 , n1208 , n1219 , n1317 , n1341 , n1404 , n1421 , n1435 , 
n1486 , n1660 , n1779 , n1794 , n1803 , n1839 , n1857 , n1860 , n2023 , n2171 , 
n2302 , n2439 , n2511 , n2598 , n2631 , n2641 , n2716 , n2774 , n2821 , n2856 , 
n3070 , n3090 , n3245 , n3282 , n3283 , n3385 , n3412 , n3430 , n3455 , n3470 , 
n3496 , n3587 , n3609 , n3626 , n3656 , n3657 , n3711 , n3757 , n3892 , n3923 , 
n3949 , n3982 , n4079 , n4114 , n4192 , n4223 , n4237 , n4274 , n4349 , n4410 , 
n4544 , n4690 , n4702 , n4706 , n4762 , n4783 , n4799 , n4800 , n4826 , n4860 , 
n4875 , n4884 , n4895 , n4904 , n4972 , n4991 , n4996 , n5007 , n5038 , n5098 , 
n5251 , n5326 , n5334 , n5394 , n5401 , n5402 , n5447 , n5456 , n5509 , n5511 , 
n5520 , n5535 , n5547 , n5567 , n5639 , n5647 , n5664 , n5743 , n5774 , n5804 , 
n5871 , n5902 , n5934 , n5954 , n6025 , n6076 , n6134 , n6187 , n6287 , n6291 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , 
n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n19 , 
n20 , n21 , n22 , n23 , n24 , n26 , n27 , n28 , n29 , n31 , 
n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , 
n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , 
n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , 
n62 , n63 , n64 , n65 , n66 , n69 , n70 , n71 , n72 , n73 , 
n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , 
n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , 
n94 , n95 , n96 , n97 , n98 , n99 , n100 , n102 , n104 , n105 , 
n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , 
n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , 
n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , 
n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n147 , 
n148 , n149 , n150 , n151 , n153 , n154 , n155 , n156 , n157 , n158 , 
n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , 
n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , 
n179 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
n200 , n201 , n202 , n203 , n205 , n206 , n207 , n208 , n209 , n210 , 
n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n241 , 
n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n251 , n252 , 
n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , 
n263 , n264 , n265 , n266 , n267 , n268 , n270 , n271 , n272 , n273 , 
n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , 
n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , 
n294 , n295 , n296 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , 
n305 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , 
n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , 
n326 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n346 , n347 , 
n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , 
n358 , n359 , n360 , n361 , n363 , n364 , n365 , n366 , n367 , n368 , 
n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
n421 , n422 , n423 , n424 , n425 , n427 , n428 , n429 , n430 , n431 , 
n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , 
n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , 
n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , 
n463 , n464 , n466 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , 
n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , 
n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n496 , 
n497 , n498 , n499 , n501 , n502 , n503 , n504 , n506 , n507 , n508 , 
n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , 
n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , 
n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n549 , n550 , 
n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , 
n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , 
n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , 
n581 , n582 , n583 , n585 , n586 , n588 , n590 , n591 , n592 , n593 , 
n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , 
n605 , n606 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , 
n616 , n617 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , 
n627 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , 
n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , 
n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n658 , 
n659 , n660 , n661 , n662 , n664 , n665 , n666 , n667 , n668 , n669 , 
n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
n680 , n681 , n682 , n683 , n684 , n685 , n686 , n688 , n689 , n690 , 
n691 , n693 , n694 , n695 , n697 , n699 , n700 , n701 , n702 , n703 , 
n704 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , 
n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , 
n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , 
n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , 
n745 , n746 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n756 , 
n757 , n758 , n759 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , 
n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n778 , 
n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , 
n789 , n790 , n791 , n793 , n794 , n795 , n797 , n798 , n799 , n800 , 
n801 , n802 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , 
n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , 
n822 , n823 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , 
n833 , n834 , n835 , n836 , n838 , n839 , n840 , n841 , n842 , n843 , 
n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , 
n854 , n855 , n856 , n857 , n858 , n859 , n860 , n862 , n863 , n865 , 
n866 , n867 , n868 , n869 , n870 , n871 , n872 , n874 , n875 , n876 , 
n877 , n878 , n879 , n880 , n881 , n883 , n884 , n885 , n886 , n887 , 
n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , 
n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , 
n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , 
n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , 
n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , 
n938 , n939 , n940 , n941 , n942 , n944 , n945 , n946 , n947 , n948 , 
n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , 
n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , 
n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , 
n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , 
n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , 
n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , 
n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1018 , n1019 , n1020 , 
n1021 , n1022 , n1023 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , 
n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , 
n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1049 , n1050 , n1051 , n1053 , 
n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , 
n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , 
n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , 
n1084 , n1085 , n1087 , n1088 , n1089 , n1090 , n1092 , n1093 , n1094 , n1095 , 
n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , 
n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , 
n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , 
n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , 
n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , 
n1146 , n1147 , n1148 , n1149 , n1150 , n1152 , n1153 , n1154 , n1155 , n1156 , 
n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , 
n1167 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , 
n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , 
n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , 
n1198 , n1199 , n1200 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1209 , 
n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1217 , n1221 , n1222 , n1223 , 
n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , 
n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , 
n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , 
n1254 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , 
n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , 
n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , 
n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , 
n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , 
n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , 
n1315 , n1316 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , 
n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , 
n1336 , n1337 , n1338 , n1339 , n1340 , n1342 , n1343 , n1344 , n1345 , n1346 , 
n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , 
n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , 
n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , 
n1377 , n1378 , n1379 , n1380 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , 
n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , 
n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1405 , n1406 , n1407 , n1408 , 
n1409 , n1410 , n1411 , n1412 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
n1420 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , 
n1431 , n1433 , n1434 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , 
n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , 
n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , 
n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1472 , n1473 , n1474 , 
n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , 
n1485 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , 
n1496 , n1497 , n1498 , n1499 , n1500 , n1502 , n1503 , n1504 , n1505 , n1506 , 
n1507 , n1508 , n1509 , n1510 , n1511 , n1513 , n1514 , n1515 , n1516 , n1517 , 
n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , 
n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , 
n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , 
n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , 
n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , 
n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , 
n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , 
n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , 
n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , 
n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , 
n1618 , n1619 , n1620 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , 
n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , 
n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , 
n1649 , n1650 , n1651 , n1652 , n1653 , n1655 , n1656 , n1657 , n1658 , n1659 , 
n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , 
n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , 
n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1691 , 
n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , 
n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , 
n1712 , n1713 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , 
n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , 
n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , 
n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , 
n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1761 , n1762 , n1763 , 
n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , 
n1775 , n1776 , n1777 , n1778 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , 
n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1795 , n1796 , 
n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1804 , n1805 , n1806 , n1807 , 
n1809 , n1810 , n1811 , n1812 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , 
n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1840 , n1841 , 
n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , 
n1852 , n1853 , n1854 , n1855 , n1856 , n1858 , n1859 , n1862 , n1863 , n1864 , 
n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , 
n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , 
n1885 , n1886 , n1887 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , 
n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1904 , n1906 , n1907 , 
n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , 
n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , 
n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , 
n1938 , n1939 , n1940 , n1941 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , 
n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1959 , 
n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
n1970 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , 
n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , 
n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n2000 , n2001 , n2002 , 
n2003 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , 
n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2024 , n2025 , 
n2026 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , 
n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , 
n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , 
n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , 
n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , 
n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , 
n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2094 , n2095 , n2096 , n2097 , 
n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , 
n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , 
n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , 
n2128 , n2129 , n2130 , n2131 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , 
n2139 , n2140 , n2141 , n2143 , n2144 , n2145 , n2147 , n2148 , n2149 , n2150 , 
n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , 
n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , 
n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , 
n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , 
n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , 
n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , 
n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , 
n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , 
n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , 
n2242 , n2243 , n2244 , n2245 , n2246 , n2248 , n2249 , n2250 , n2251 , n2252 , 
n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2263 , 
n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , 
n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , 
n2284 , n2285 , n2286 , n2287 , n2288 , n2290 , n2291 , n2292 , n2293 , n2294 , 
n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2303 , n2304 , n2305 , n2306 , 
n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , 
n2317 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , 
n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2337 , n2338 , 
n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , 
n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , 
n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , 
n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , 
n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , 
n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , 
n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , 
n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , 
n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2437 , n2438 , n2441 , n2442 , 
n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , 
n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , 
n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , 
n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , 
n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , 
n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , 
n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2512 , n2513 , 
n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , 
n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , 
n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , 
n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2552 , n2553 , n2555 , n2556 , 
n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2564 , n2565 , n2566 , n2567 , 
n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2578 , 
n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , 
n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2599 , 
n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
n2630 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2639 , n2640 , n2642 , 
n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , 
n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , 
n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , 
n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , 
n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , 
n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , 
n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , 
n2713 , n2715 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , 
n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , 
n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2745 , 
n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , 
n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , 
n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2775 , n2776 , 
n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , 
n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , 
n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2805 , n2806 , n2807 , 
n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , 
n2818 , n2819 , n2820 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , 
n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2837 , n2838 , n2839 , 
n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , 
n2852 , n2853 , n2854 , n2855 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , 
n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , 
n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , 
n2883 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , 
n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , 
n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , 
n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , 
n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , 
n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , 
n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , 
n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , 
n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , 
n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , 
n2984 , n2985 , n2986 , n2987 , n2989 , n2990 , n2991 , n2992 , n2994 , n2995 , 
n2996 , n2997 , n2998 , n2999 , n3000 , n3002 , n3003 , n3004 , n3005 , n3006 , 
n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , 
n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , 
n3027 , n3028 , n3029 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3038 , 
n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , 
n3049 , n3050 , n3051 , n3052 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
n3060 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3071 , 
n3072 , n3073 , n3074 , n3075 , n3076 , n3078 , n3079 , n3080 , n3081 , n3082 , 
n3083 , n3085 , n3086 , n3087 , n3088 , n3091 , n3092 , n3093 , n3094 , n3095 , 
n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , 
n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , 
n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , 
n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , 
n3136 , n3137 , n3138 , n3139 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , 
n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , 
n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3165 , n3166 , n3167 , 
n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3175 , n3176 , n3177 , n3178 , 
n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , 
n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , 
n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , 
n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , 
n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , 
n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , 
n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3246 , n3247 , n3248 , n3249 , 
n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
n3280 , n3281 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , 
n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , 
n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , 
n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , 
n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , 
n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , 
n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3350 , n3351 , n3352 , 
n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3361 , n3362 , n3363 , 
n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , 
n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , 
n3384 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , 
n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , 
n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3413 , n3414 , n3415 , 
n3416 , n3417 , n3418 , n3419 , n3420 , n3422 , n3423 , n3424 , n3425 , n3426 , 
n3427 , n3428 , n3429 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , 
n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , 
n3448 , n3449 , n3450 , n3452 , n3453 , n3454 , n3456 , n3457 , n3458 , n3459 , 
n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , 
n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3490 , n3491 , 
n3492 , n3493 , n3494 , n3495 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , 
n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , 
n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3520 , n3521 , n3522 , n3523 , 
n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , 
n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3543 , n3544 , 
n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , 
n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , 
n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3574 , n3575 , 
n3576 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , 
n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , 
n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , 
n3608 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , 
n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3627 , n3628 , n3629 , 
n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , 
n3640 , n3641 , n3642 , n3643 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , 
n3651 , n3652 , n3653 , n3654 , n3655 , n3658 , n3659 , n3660 , n3661 , n3662 , 
n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , 
n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3682 , n3683 , 
n3684 , n3685 , n3686 , n3688 , n3689 , n3691 , n3692 , n3693 , n3694 , n3695 , 
n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , 
n3706 , n3707 , n3708 , n3709 , n3710 , n3712 , n3713 , n3714 , n3715 , n3716 , 
n3718 , n3719 , n3720 , n3721 , n3722 , n3724 , n3725 , n3726 , n3727 , n3729 , 
n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , 
n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3758 , n3759 , n3760 , 
n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , 
n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , 
n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , 
n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , 
n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , 
n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , 
n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3830 , n3831 , n3832 , 
n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , 
n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , 
n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , 
n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , 
n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , 
n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3893 , 
n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , 
n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3912 , n3913 , n3914 , 
n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3924 , n3925 , 
n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , 
n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , 
n3946 , n3947 , n3948 , n3950 , n3951 , n3952 , n3953 , n3954 , n3956 , n3957 , 
n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , 
n3968 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , 
n3979 , n3980 , n3981 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , 
n3990 , n3991 , n3992 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , 
n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , 
n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , 
n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4029 , n4030 , n4031 , 
n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , 
n4042 , n4044 , n4045 , n4046 , n4047 , n4048 , n4051 , n4052 , n4053 , n4054 , 
n4055 , n4056 , n4057 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , 
n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , 
n4076 , n4077 , n4078 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , 
n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , 
n4097 , n4099 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , 
n4109 , n4110 , n4111 , n4112 , n4113 , n4115 , n4116 , n4117 , n4118 , n4120 , 
n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , 
n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , 
n4141 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , 
n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , 
n4162 , n4163 , n4165 , n4166 , n4167 , n4169 , n4170 , n4171 , n4172 , n4173 , 
n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , 
n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4193 , n4194 , 
n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , 
n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , 
n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4224 , n4225 , 
n4226 , n4227 , n4228 , n4229 , n4230 , n4232 , n4233 , n4234 , n4235 , n4236 , 
n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , 
n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , 
n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , 
n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4275 , n4276 , n4277 , n4278 , 
n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , 
n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , 
n4299 , n4300 , n4301 , n4302 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , 
n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4320 , 
n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
n4333 , n4334 , n4335 , n4337 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , 
n4348 , n4350 , n4351 , n4352 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , 
n4360 , n4361 , n4362 , n4363 , n4364 , n4366 , n4367 , n4368 , n4369 , n4371 , 
n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , 
n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , 
n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , 
n4402 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4411 , n4412 , n4413 , 
n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , 
n4424 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4433 , n4434 , n4435 , 
n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , 
n4446 , n4447 , n4449 , n4450 , n4452 , n4453 , n4455 , n4456 , n4457 , n4458 , 
n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4468 , n4469 , 
n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , 
n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , 
n4490 , n4491 , n4492 , n4493 , n4494 , n4496 , n4497 , n4498 , n4499 , n4500 , 
n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
n4541 , n4542 , n4543 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , 
n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , 
n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , 
n4573 , n4574 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , 
n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , 
n4595 , n4596 , n4597 , n4598 , n4600 , n4601 , n4602 , n4603 , n4605 , n4606 , 
n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4616 , n4617 , 
n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , 
n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , 
n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , 
n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , 
n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , 
n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , 
n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , 
n4688 , n4689 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , 
n4699 , n4700 , n4701 , n4703 , n4704 , n4705 , n4707 , n4708 , n4709 , n4710 , 
n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4721 , 
n4722 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , 
n4733 , n4734 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4744 , 
n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , 
n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4763 , n4764 , n4765 , 
n4766 , n4767 , n4768 , n4769 , n4770 , n4772 , n4773 , n4774 , n4775 , n4776 , 
n4778 , n4779 , n4780 , n4781 , n4782 , n4784 , n4785 , n4786 , n4787 , n4788 , 
n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , 
n4801 , n4802 , n4803 , n4804 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , 
n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , 
n4822 , n4824 , n4825 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4834 , 
n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , 
n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , 
n4855 , n4856 , n4857 , n4858 , n4859 , n4861 , n4862 , n4863 , n4864 , n4865 , 
n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4876 , n4877 , 
n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4885 , n4886 , n4887 , n4889 , 
n4890 , n4891 , n4892 , n4893 , n4894 , n4896 , n4897 , n4898 , n4899 , n4900 , 
n4901 , n4902 , n4903 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , 
n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , 
n4923 , n4924 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , 
n4934 , n4935 , n4936 , n4938 , n4939 , n4941 , n4942 , n4943 , n4944 , n4945 , 
n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , 
n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , 
n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4973 , n4974 , n4975 , n4976 , 
n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , 
n4987 , n4988 , n4989 , n4990 , n4992 , n4993 , n4994 , n4995 , n4997 , n4998 , 
n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5008 , n5009 , 
n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , 
n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , 
n5030 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5039 , n5040 , n5041 , 
n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , 
n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , 
n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , 
n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , 
n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , 
n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5099 , n5100 , n5101 , n5103 , 
n5104 , n5105 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , 
n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , 
n5125 , n5126 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , 
n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , 
n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , 
n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , 
n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , 
n5176 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , 
n5187 , n5188 , n5189 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , 
n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5206 , n5207 , n5208 , 
n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , 
n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , 
n5229 , n5230 , n5231 , n5232 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , 
n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5249 , n5250 , 
n5253 , n5254 , n5255 , n5256 , n5257 , n5259 , n5260 , n5261 , n5262 , n5263 , 
n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , 
n5274 , n5275 , n5276 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , 
n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , 
n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , 
n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5315 , 
n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , 
n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5335 , n5336 , n5337 , n5338 , 
n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , 
n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , 
n5359 , n5360 , n5361 , n5362 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , 
n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , 
n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , 
n5390 , n5391 , n5392 , n5393 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , 
n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , 
n5423 , n5424 , n5425 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , 
n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , 
n5444 , n5445 , n5446 , n5448 , n5449 , n5451 , n5452 , n5453 , n5454 , n5455 , 
n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , 
n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , 
n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , 
n5487 , n5488 , n5489 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , 
n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5507 , n5508 , 
n5510 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5522 , n5523 , 
n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , 
n5534 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , 
n5545 , n5546 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , 
n5556 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , 
n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , 
n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , 
n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , 
n5598 , n5599 , n5600 , n5601 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , 
n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , 
n5619 , n5620 , n5621 , n5622 , n5623 , n5625 , n5626 , n5627 , n5628 , n5629 , 
n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5640 , n5641 , 
n5642 , n5643 , n5644 , n5645 , n5646 , n5648 , n5649 , n5650 , n5651 , n5652 , 
n5653 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5663 , n5665 , 
n5666 , n5667 , n5668 , n5669 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , 
n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , 
n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , 
n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , 
n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , 
n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , 
n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , 
n5738 , n5739 , n5740 , n5741 , n5742 , n5744 , n5745 , n5746 , n5747 , n5748 , 
n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , 
n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , 
n5769 , n5770 , n5771 , n5772 , n5773 , n5775 , n5776 , n5777 , n5778 , n5779 , 
n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , 
n5790 , n5791 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , 
n5801 , n5802 , n5803 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , 
n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , 
n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5830 , n5831 , n5832 , 
n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , 
n5843 , n5844 , n5845 , n5846 , n5847 , n5849 , n5850 , n5851 , n5853 , n5854 , 
n5855 , n5856 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , 
n5866 , n5867 , n5868 , n5869 , n5870 , n5872 , n5873 , n5874 , n5875 , n5876 , 
n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5884 , n5885 , n5886 , n5887 , 
n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , 
n5898 , n5899 , n5900 , n5903 , n5904 , n5905 , n5908 , n5909 , n5910 , n5911 , 
n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , 
n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , 
n5932 , n5933 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , 
n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , 
n5953 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , 
n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , 
n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , 
n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5993 , n5994 , 
n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , 
n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , 
n6016 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6026 , n6027 , 
n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6035 , n6036 , n6037 , n6039 , 
n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , 
n6050 , n6051 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , 
n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , 
n6072 , n6073 , n6074 , n6075 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , 
n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , 
n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , 
n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , 
n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , 
n6123 , n6124 , n6125 , n6126 , n6127 , n6129 , n6130 , n6131 , n6132 , n6133 , 
n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , 
n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6155 , 
n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , 
n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6176 , 
n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , 
n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , 
n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , 
n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , 
n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , 
n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , 
n6238 , n6239 , n6240 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , 
n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , 
n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , 
n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , 
n6279 , n6280 , n6281 , n6283 , n6284 , n6285 , n6286 , n6288 , n6289 , n6290 , 
n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , 
n6302 , n6303 ;
    and g0 ( n2374 , n2396 , n4879 );
    or g1 ( n5255 , n6097 , n79 );
    not g2 ( n6046 , n795 );
    not g3 ( n4905 , n4925 );
    or g4 ( n4649 , n5490 , n2690 );
    not g5 ( n1538 , n1273 );
    or g6 ( n6028 , n2326 , n1323 );
    and g7 ( n1096 , n3740 , n4649 );
    not g8 ( n5777 , n858 );
    not g9 ( n867 , n5749 );
    or g10 ( n1796 , n5994 , n4457 );
    not g11 ( n3259 , n2635 );
    or g12 ( n1249 , n643 , n3526 );
    and g13 ( n5661 , n1225 , n5274 );
    and g14 ( n3668 , n3086 , n436 );
    or g15 ( n2637 , n567 , n1629 );
    and g16 ( n2776 , n1830 , n1522 );
    not g17 ( n1703 , n5258 );
    nor g18 ( n2324 , n6019 , n5869 );
    or g19 ( n2163 , n5949 , n648 );
    not g20 ( n4373 , n1767 );
    or g21 ( n2717 , n3387 , n54 );
    nor g22 ( n2252 , n4081 , n5739 );
    nor g23 ( n4296 , n4173 , n4681 );
    not g24 ( n773 , n4668 );
    nor g25 ( n2960 , n4509 , n3738 );
    and g26 ( n843 , n2274 , n4923 );
    nor g27 ( n2330 , n874 , n5669 );
    not g28 ( n5666 , n4876 );
    or g29 ( n946 , n558 , n4345 );
    nor g30 ( n3697 , n2925 , n4629 );
    not g31 ( n4929 , n1655 );
    or g32 ( n4521 , n28 , n3909 );
    or g33 ( n2869 , n1784 , n3312 );
    not g34 ( n3692 , n5662 );
    or g35 ( n4660 , n460 , n4617 );
    not g36 ( n945 , n861 );
    nor g37 ( n1134 , n3060 , n2861 );
    nor g38 ( n3946 , n4516 , n3748 );
    and g39 ( n2986 , n1912 , n1215 );
    not g40 ( n4027 , n2241 );
    not g41 ( n1799 , n1665 );
    not g42 ( n4224 , n4794 );
    and g43 ( n4421 , n1369 , n206 );
    or g44 ( n2173 , n3370 , n2677 );
    and g45 ( n700 , n5896 , n1915 );
    not g46 ( n778 , n438 );
    and g47 ( n4305 , n930 , n1849 );
    not g48 ( n4744 , n3752 );
    or g49 ( n382 , n1693 , n2433 );
    and g50 ( n730 , n3867 , n1561 );
    nor g51 ( n3317 , n1488 , n686 );
    nor g52 ( n4014 , n4923 , n5781 );
    nor g53 ( n6084 , n500 , n3391 );
    or g54 ( n3093 , n2300 , n5008 );
    not g55 ( n2618 , n4028 );
    and g56 ( n469 , n2573 , n4470 );
    or g57 ( n5094 , n1704 , n598 );
    nor g58 ( n5472 , n1337 , n1685 );
    and g59 ( n626 , n920 , n3662 );
    not g60 ( n1783 , n994 );
    nor g61 ( n4359 , n1201 , n1327 );
    and g62 ( n4144 , n5791 , n1357 );
    nor g63 ( n3422 , n594 , n4940 );
    nor g64 ( n3538 , n4467 , n2487 );
    nor g65 ( n5875 , n3553 , n5427 );
    or g66 ( n1199 , n372 , n3874 );
    and g67 ( n373 , n5121 , n5482 );
    or g68 ( n5917 , n2932 , n262 );
    nor g69 ( n6146 , n2537 , n134 );
    or g70 ( n418 , n3148 , n1003 );
    nor g71 ( n477 , n2626 , n1348 );
    or g72 ( n1427 , n5827 , n4328 );
    and g73 ( n1548 , n17 , n6249 );
    or g74 ( n3662 , n5784 , n6284 );
    nor g75 ( n4935 , n145 , n5573 );
    or g76 ( n3283 , n2938 , n1955 );
    nor g77 ( n2105 , n5662 , n3873 );
    and g78 ( n125 , n2052 , n3655 );
    and g79 ( n1792 , n4362 , n338 );
    and g80 ( n5581 , n5868 , n80 );
    or g81 ( n3930 , n5697 , n271 );
    not g82 ( n1822 , n2761 );
    not g83 ( n1840 , n4896 );
    not g84 ( n3960 , n2146 );
    not g85 ( n2915 , n3511 );
    not g86 ( n4619 , n3410 );
    and g87 ( n5496 , n2241 , n6021 );
    not g88 ( n1223 , n2393 );
    or g89 ( n5212 , n2164 , n5024 );
    or g90 ( n2083 , n2804 , n2715 );
    and g91 ( n5867 , n4408 , n3203 );
    and g92 ( n535 , n2669 , n3984 );
    or g93 ( n6196 , n439 , n3805 );
    or g94 ( n2028 , n3680 , n3505 );
    not g95 ( n5028 , n5578 );
    or g96 ( n2606 , n213 , n515 );
    not g97 ( n4251 , n4458 );
    not g98 ( n4494 , n1151 );
    not g99 ( n2029 , n5973 );
    not g100 ( n4517 , n1820 );
    and g101 ( n424 , n3932 , n3489 );
    or g102 ( n4636 , n1198 , n4902 );
    not g103 ( n6174 , n2813 );
    or g104 ( n2131 , n24 , n6173 );
    or g105 ( n1670 , n4805 , n1512 );
    and g106 ( n5818 , n3305 , n3061 );
    or g107 ( n4052 , n3297 , n1072 );
    not g108 ( n1356 , n4561 );
    and g109 ( n5614 , n1758 , n4239 );
    or g110 ( n4815 , n3746 , n1646 );
    or g111 ( n2113 , n1942 , n1655 );
    or g112 ( n1063 , n5484 , n4076 );
    or g113 ( n2184 , n1735 , n4861 );
    nor g114 ( n3746 , n2306 , n4896 );
    or g115 ( n4487 , n313 , n371 );
    or g116 ( n2944 , n2909 , n3820 );
    not g117 ( n5311 , n2777 );
    and g118 ( n2602 , n3882 , n602 );
    not g119 ( n3350 , n4812 );
    nor g120 ( n5279 , n5586 , n1022 );
    nor g121 ( n3007 , n51 , n860 );
    or g122 ( n2092 , n4222 , n1527 );
    not g123 ( n836 , n3092 );
    not g124 ( n3301 , n1802 );
    and g125 ( n1252 , n5913 , n1649 );
    nor g126 ( n771 , n5271 , n1806 );
    nor g127 ( n1889 , n1685 , n3115 );
    not g128 ( n4879 , n2097 );
    or g129 ( n3192 , n2575 , n4566 );
    not g130 ( n5888 , n5099 );
    or g131 ( n5689 , n5863 , n3605 );
    nor g132 ( n3059 , n4451 , n2993 );
    or g133 ( n1574 , n896 , n6202 );
    or g134 ( n5089 , n2165 , n93 );
    and g135 ( n3563 , n424 , n689 );
    not g136 ( n3924 , n4316 );
    not g137 ( n1061 , n4049 );
    and g138 ( n3002 , n2202 , n4005 );
    nor g139 ( n4990 , n4545 , n2446 );
    not g140 ( n3461 , n3984 );
    or g141 ( n4407 , n3147 , n949 );
    nor g142 ( n166 , n2337 , n2945 );
    or g143 ( n3726 , n6051 , n3033 );
    not g144 ( n442 , n1471 );
    not g145 ( n844 , n4937 );
    and g146 ( n3379 , n585 , n3378 );
    and g147 ( n1136 , n2067 , n4761 );
    nor g148 ( n468 , n322 , n5137 );
    and g149 ( n4405 , n5301 , n5444 );
    nor g150 ( n524 , n1448 , n4521 );
    and g151 ( n5036 , n4712 , n5672 );
    or g152 ( n2319 , n3287 , n3550 );
    not g153 ( n2615 , n3687 );
    not g154 ( n2647 , n6221 );
    not g155 ( n6147 , n469 );
    nor g156 ( n3732 , n2566 , n4513 );
    not g157 ( n5032 , n2333 );
    or g158 ( n4826 , n3219 , n3054 );
    or g159 ( n3289 , n793 , n3201 );
    and g160 ( n337 , n5140 , n998 );
    not g161 ( n1324 , n4156 );
    nor g162 ( n4387 , n1142 , n3631 );
    not g163 ( n2049 , n2918 );
    nor g164 ( n1009 , n1869 , n349 );
    or g165 ( n1297 , n5426 , n1163 );
    nor g166 ( n2876 , n261 , n1078 );
    not g167 ( n5121 , n2042 );
    not g168 ( n1263 , n2412 );
    or g169 ( n566 , n2454 , n4299 );
    nor g170 ( n3113 , n1146 , n3759 );
    or g171 ( n324 , n5296 , n1284 );
    not g172 ( n3884 , n5078 );
    or g173 ( n3901 , n2731 , n2711 );
    not g174 ( n1705 , n4888 );
    nor g175 ( n4085 , n3838 , n4917 );
    not g176 ( n2996 , n1432 );
    not g177 ( n6298 , n70 );
    not g178 ( n1763 , n1917 );
    or g179 ( n2946 , n834 , n6124 );
    or g180 ( n679 , n5901 , n3967 );
    and g181 ( n645 , n133 , n5638 );
    nor g182 ( n6097 , n3360 , n1304 );
    not g183 ( n2366 , n1458 );
    not g184 ( n106 , n1656 );
    nor g185 ( n1418 , n1324 , n3529 );
    not g186 ( n1886 , n6189 );
    not g187 ( n1854 , n4885 );
    and g188 ( n1179 , n3214 , n4136 );
    and g189 ( n3366 , n3994 , n1472 );
    nor g190 ( n2904 , n1874 , n2238 );
    nor g191 ( n2670 , n4288 , n802 );
    not g192 ( n5101 , n4483 );
    not g193 ( n3227 , n152 );
    and g194 ( n2721 , n2355 , n531 );
    not g195 ( n5712 , n1416 );
    nor g196 ( n4054 , n2114 , n5442 );
    not g197 ( n4120 , n1777 );
    not g198 ( n6051 , n5640 );
    and g199 ( n5438 , n5893 , n1984 );
    not g200 ( n4268 , n5452 );
    not g201 ( n3048 , n114 );
    and g202 ( n249 , n1362 , n3531 );
    or g203 ( n2101 , n3440 , n2122 );
    and g204 ( n1106 , n1875 , n6001 );
    and g205 ( n1337 , n2763 , n5977 );
    not g206 ( n1917 , n2109 );
    not g207 ( n4705 , n5950 );
    nor g208 ( n2214 , n4141 , n4688 );
    not g209 ( n3488 , n1734 );
    not g210 ( n3832 , n5420 );
    not g211 ( n5422 , n317 );
    nor g212 ( n2548 , n5433 , n3113 );
    not g213 ( n5562 , n1084 );
    nor g214 ( n2249 , n1503 , n2269 );
    not g215 ( n3601 , n1721 );
    nor g216 ( n1850 , n4922 , n1472 );
    or g217 ( n2627 , n766 , n2384 );
    and g218 ( n1765 , n526 , n3330 );
    or g219 ( n5708 , n5254 , n5204 );
    nor g220 ( n336 , n5416 , n2951 );
    or g221 ( n1960 , n495 , n1843 );
    nor g222 ( n3602 , n6175 , n5491 );
    and g223 ( n6086 , n5132 , n4510 );
    or g224 ( n1265 , n42 , n1198 );
    not g225 ( n554 , n5519 );
    or g226 ( n5816 , n1598 , n5579 );
    not g227 ( n1310 , n1628 );
    not g228 ( n5753 , n488 );
    and g229 ( n3082 , n1612 , n3665 );
    not g230 ( n3186 , n476 );
    nor g231 ( n6049 , n2256 , n2277 );
    or g232 ( n3695 , n1223 , n3139 );
    or g233 ( n1412 , n2226 , n3194 );
    nor g234 ( n5979 , n2915 , n757 );
    and g235 ( n668 , n5202 , n2923 );
    or g236 ( n933 , n3239 , n3005 );
    nor g237 ( n4837 , n2810 , n2662 );
    or g238 ( n3773 , n886 , n2952 );
    not g239 ( n2295 , n5927 );
    or g240 ( n1470 , n4862 , n5705 );
    nor g241 ( n6031 , n1217 , n5606 );
    or g242 ( n3830 , n2006 , n3954 );
    or g243 ( n598 , n15 , n4883 );
    or g244 ( n5758 , n1008 , n4229 );
    not g245 ( n5096 , n376 );
    and g246 ( n4228 , n1653 , n4847 );
    nor g247 ( n2718 , n1841 , n4096 );
    or g248 ( n4812 , n4487 , n4140 );
    nor g249 ( n2707 , n4425 , n1493 );
    or g250 ( n3622 , n5539 , n1840 );
    and g251 ( n5029 , n5052 , n2207 );
    or g252 ( n6279 , n351 , n4384 );
    not g253 ( n51 , n527 );
    and g254 ( n6009 , n5138 , n4172 );
    nor g255 ( n263 , n4858 , n46 );
    not g256 ( n2413 , n2534 );
    nor g257 ( n187 , n2499 , n194 );
    not g258 ( n5947 , n3378 );
    not g259 ( n4881 , n4332 );
    or g260 ( n5211 , n6128 , n403 );
    nor g261 ( n641 , n4056 , n816 );
    nor g262 ( n4715 , n6017 , n2994 );
    and g263 ( n322 , n3069 , n4067 );
    not g264 ( n5227 , n2806 );
    and g265 ( n2768 , n5613 , n4466 );
    nor g266 ( n4813 , n2383 , n553 );
    or g267 ( n4394 , n1463 , n5787 );
    or g268 ( n2595 , n6165 , n5300 );
    and g269 ( n766 , n5262 , n4658 );
    or g270 ( n4895 , n65 , n1406 );
    nor g271 ( n296 , n174 , n2855 );
    not g272 ( n3418 , n4239 );
    or g273 ( n6022 , n748 , n196 );
    nor g274 ( n5383 , n6267 , n2231 );
    or g275 ( n3020 , n2068 , n5373 );
    nor g276 ( n1053 , n3315 , n2597 );
    and g277 ( n4663 , n2049 , n308 );
    not g278 ( n931 , n5449 );
    or g279 ( n4609 , n3199 , n2298 );
    nor g280 ( n486 , n426 , n3567 );
    and g281 ( n3019 , n1417 , n3058 );
    and g282 ( n6269 , n6239 , n6289 );
    not g283 ( n963 , n1620 );
    and g284 ( n6299 , n2806 , n421 );
    nor g285 ( n2754 , n4989 , n3824 );
    or g286 ( n2662 , n2258 , n1863 );
    nor g287 ( n3327 , n6175 , n3300 );
    not g288 ( n4838 , n1399 );
    nor g289 ( n1149 , n1881 , n3769 );
    and g290 ( n4087 , n2593 , n4191 );
    or g291 ( n5710 , n6209 , n5472 );
    and g292 ( n4383 , n4759 , n1810 );
    not g293 ( n4275 , n5627 );
    or g294 ( n1229 , n437 , n3942 );
    or g295 ( n4181 , n1845 , n1736 );
    and g296 ( n5191 , n296 , n1241 );
    or g297 ( n2671 , n691 , n939 );
    nor g298 ( n6037 , n4568 , n551 );
    not g299 ( n2741 , n5730 );
    nor g300 ( n2612 , n5131 , n5197 );
    and g301 ( n5583 , n4874 , n4444 );
    or g302 ( n6119 , n2318 , n446 );
    or g303 ( n6100 , n4322 , n2522 );
    or g304 ( n4717 , n1722 , n4261 );
    nor g305 ( n1618 , n5260 , n1987 );
    or g306 ( n1573 , n5918 , n422 );
    or g307 ( n5352 , n3203 , n3857 );
    and g308 ( n3751 , n6298 , n2820 );
    not g309 ( n5461 , n657 );
    not g310 ( n4130 , n3444 );
    or g311 ( n6164 , n2726 , n1859 );
    not g312 ( n3354 , n2419 );
    nor g313 ( n2427 , n2854 , n4784 );
    not g314 ( n4046 , n462 );
    not g315 ( n1433 , n5049 );
    and g316 ( n939 , n5644 , n3629 );
    and g317 ( n1576 , n4739 , n3588 );
    or g318 ( n1490 , n4962 , n3724 );
    not g319 ( n1167 , n3488 );
    and g320 ( n5184 , n5179 , n5041 );
    or g321 ( n2338 , n6095 , n5658 );
    not g322 ( n2449 , n86 );
    or g323 ( n2235 , n4986 , n2478 );
    not g324 ( n1116 , n4556 );
    and g325 ( n3141 , n5404 , n1984 );
    or g326 ( n4254 , n5450 , n2093 );
    or g327 ( n4628 , n4292 , n1452 );
    or g328 ( n1932 , n4286 , n3708 );
    nor g329 ( n4151 , n2312 , n3176 );
    or g330 ( n3297 , n5327 , n2248 );
    and g331 ( n4156 , n136 , n4392 );
    or g332 ( n571 , n4711 , n38 );
    and g333 ( n1144 , n6026 , n2217 );
    or g334 ( n3159 , n3500 , n422 );
    or g335 ( n1711 , n4735 , n3960 );
    or g336 ( n5273 , n4218 , n3995 );
    and g337 ( n4687 , n3032 , n4922 );
    nor g338 ( n856 , n6254 , n1093 );
    not g339 ( n1997 , n859 );
    or g340 ( n2430 , n2350 , n896 );
    or g341 ( n1819 , n6255 , n4956 );
    or g342 ( n957 , n2176 , n4148 );
    not g343 ( n5596 , n4509 );
    and g344 ( n4153 , n6294 , n2957 );
    nor g345 ( n6023 , n1688 , n5085 );
    not g346 ( n5757 , n5084 );
    not g347 ( n5324 , n3534 );
    not g348 ( n3224 , n1039 );
    and g349 ( n3047 , n2609 , n1416 );
    not g350 ( n6041 , n1157 );
    not g351 ( n4683 , n4743 );
    not g352 ( n1309 , n2010 );
    not g353 ( n4997 , n3830 );
    or g354 ( n1927 , n390 , n520 );
    nor g355 ( n3787 , n4149 , n1393 );
    nor g356 ( n5093 , n2051 , n2762 );
    nor g357 ( n4883 , n581 , n979 );
    or g358 ( n3406 , n3540 , n4714 );
    and g359 ( n1977 , n4927 , n1604 );
    not g360 ( n6205 , n4102 );
    and g361 ( n3682 , n878 , n3582 );
    or g362 ( n3144 , n3723 , n4970 );
    not g363 ( n1172 , n322 );
    nor g364 ( n1600 , n631 , n276 );
    nor g365 ( n6115 , n2027 , n5622 );
    not g366 ( n1002 , n2719 );
    or g367 ( n6162 , n4236 , n1481 );
    and g368 ( n6029 , n5866 , n4390 );
    not g369 ( n464 , n6028 );
    or g370 ( n3493 , n6256 , n4711 );
    not g371 ( n6108 , n2897 );
    and g372 ( n2310 , n3594 , n5678 );
    not g373 ( n2182 , n4323 );
    and g374 ( n3279 , n1364 , n1105 );
    not g375 ( n1306 , n3443 );
    or g376 ( n1790 , n2737 , n4738 );
    not g377 ( n3256 , n645 );
    not g378 ( n967 , n4254 );
    or g379 ( n4369 , n5605 , n6193 );
    nor g380 ( n516 , n696 , n6292 );
    or g381 ( n6006 , n4179 , n4912 );
    not g382 ( n3894 , n5162 );
    not g383 ( n4887 , n791 );
    nor g384 ( n5146 , n1358 , n1532 );
    not g385 ( n37 , n4505 );
    or g386 ( n1439 , n2247 , n4049 );
    and g387 ( n5972 , n4506 , n1910 );
    nor g388 ( n619 , n861 , n1070 );
    and g389 ( n1663 , n1197 , n261 );
    or g390 ( n443 , n3068 , n2136 );
    not g391 ( n1507 , n1621 );
    not g392 ( n3932 , n6282 );
    or g393 ( n5731 , n3544 , n5674 );
    not g394 ( n5464 , n4164 );
    or g395 ( n6089 , n4940 , n796 );
    nor g396 ( n1897 , n4347 , n65 );
    or g397 ( n2408 , n6128 , n4855 );
    and g398 ( n2942 , n2842 , n3062 );
    or g399 ( n1860 , n5027 , n267 );
    nor g400 ( n2309 , n2524 , n319 );
    and g401 ( n5017 , n4183 , n6013 );
    nor g402 ( n5004 , n2266 , n603 );
    nor g403 ( n3753 , n298 , n3743 );
    nor g404 ( n4736 , n5795 , n336 );
    nor g405 ( n4415 , n4833 , n1016 );
    not g406 ( n3769 , n2860 );
    not g407 ( n4526 , n981 );
    not g408 ( n4607 , n583 );
    nor g409 ( n4343 , n523 , n186 );
    and g410 ( n1491 , n2538 , n3354 );
    or g411 ( n791 , n3374 , n3316 );
    nor g412 ( n1613 , n4168 , n2828 );
    or g413 ( n2808 , n2127 , n5718 );
    nor g414 ( n746 , n4580 , n5517 );
    not g415 ( n3532 , n2730 );
    nor g416 ( n1557 , n1064 , n2613 );
    or g417 ( n4679 , n1535 , n4893 );
    not g418 ( n5 , n3212 );
    nor g419 ( n6232 , n5260 , n4596 );
    or g420 ( n552 , n4113 , n3887 );
    or g421 ( n3126 , n2246 , n1387 );
    not g422 ( n3931 , n1297 );
    not g423 ( n5178 , n1990 );
    or g424 ( n362 , n3485 , n5236 );
    nor g425 ( n1922 , n4390 , n1199 );
    nor g426 ( n4416 , n4495 , n5940 );
    and g427 ( n1243 , n557 , n3968 );
    and g428 ( n4158 , n649 , n639 );
    nor g429 ( n1326 , n751 , n5655 );
    or g430 ( n3075 , n3197 , n6016 );
    or g431 ( n4701 , n5849 , n320 );
    nor g432 ( n1661 , n965 , n4132 );
    and g433 ( n5601 , n3081 , n4087 );
    or g434 ( n4115 , n5518 , n5719 );
    and g435 ( n1595 , n4565 , n145 );
    nor g436 ( n4064 , n5059 , n4151 );
    nor g437 ( n4230 , n369 , n3797 );
    or g438 ( n3564 , n3030 , n4317 );
    or g439 ( n2784 , n4227 , n4085 );
    or g440 ( n3459 , n463 , n1033 );
    or g441 ( n4904 , n2618 , n3868 );
    not g442 ( n3381 , n943 );
    not g443 ( n953 , n4452 );
    not g444 ( n5929 , n1269 );
    and g445 ( n1417 , n3950 , n1423 );
    not g446 ( n403 , n3360 );
    or g447 ( n4711 , n2728 , n5649 );
    and g448 ( n1081 , n4187 , n6149 );
    nor g449 ( n3879 , n4758 , n840 );
    or g450 ( n3359 , n2184 , n1174 );
    or g451 ( n2902 , n2360 , n5874 );
    or g452 ( n2349 , n5131 , n5687 );
    or g453 ( n2604 , n529 , n2366 );
    not g454 ( n2331 , n1152 );
    not g455 ( n1620 , n2347 );
    nor g456 ( n713 , n483 , n3194 );
    nor g457 ( n5429 , n3141 , n3423 );
    nor g458 ( n2134 , n3977 , n4643 );
    not g459 ( n4994 , n1097 );
    nor g460 ( n5168 , n5516 , n3152 );
    nor g461 ( n5766 , n2213 , n5225 );
    and g462 ( n2044 , n4206 , n5946 );
    and g463 ( n17 , n1041 , n4796 );
    nor g464 ( n75 , n1213 , n273 );
    nor g465 ( n809 , n1753 , n3495 );
    nor g466 ( n5018 , n734 , n1862 );
    not g467 ( n1754 , n3222 );
    or g468 ( n4664 , n855 , n1977 );
    nor g469 ( n563 , n3969 , n5062 );
    and g470 ( n2696 , n209 , n4362 );
    not g471 ( n5099 , n5929 );
    not g472 ( n3474 , n3130 );
    nor g473 ( n1325 , n3232 , n2110 );
    not g474 ( n3290 , n5728 );
    not g475 ( n3950 , n3585 );
    nor g476 ( n2822 , n1237 , n3029 );
    nor g477 ( n2193 , n251 , n651 );
    or g478 ( n739 , n3885 , n1948 );
    and g479 ( n6184 , n392 , n5852 );
    or g480 ( n4357 , n577 , n5359 );
    and g481 ( n3893 , n2929 , n5728 );
    and g482 ( n3898 , n2581 , n1388 );
    not g483 ( n3182 , n5396 );
    not g484 ( n5376 , n951 );
    and g485 ( n5773 , n5183 , n3308 );
    not g486 ( n19 , n1346 );
    nor g487 ( n5267 , n2360 , n5419 );
    and g488 ( n1668 , n564 , n347 );
    nor g489 ( n5574 , n2494 , n721 );
    buf g490 ( n1168 , n1857 );
    nor g491 ( n1194 , n4319 , n4424 );
    nor g492 ( n5812 , n3318 , n1286 );
    or g493 ( n1572 , n4311 , n3933 );
    nor g494 ( n3288 , n230 , n1056 );
    not g495 ( n2825 , n1346 );
    not g496 ( n225 , n4058 );
    not g497 ( n683 , n1974 );
    and g498 ( n2490 , n5720 , n3479 );
    or g499 ( n4634 , n4028 , n6296 );
    or g500 ( n4125 , n5935 , n2664 );
    or g501 ( n4213 , n658 , n2402 );
    not g502 ( n3767 , n1434 );
    not g503 ( n1483 , n224 );
    not g504 ( n5140 , n5059 );
    not g505 ( n1834 , n3382 );
    not g506 ( n346 , n538 );
    and g507 ( n5420 , n4444 , n3103 );
    nor g508 ( n2469 , n30 , n330 );
    nor g509 ( n5395 , n505 , n5155 );
    and g510 ( n142 , n2050 , n3831 );
    and g511 ( n5620 , n4220 , n2848 );
    not g512 ( n4906 , n1516 );
    nor g513 ( n6186 , n6038 , n1824 );
    nor g514 ( n5108 , n28 , n3056 );
    not g515 ( n5742 , n2027 );
    not g516 ( n3316 , n2767 );
    not g517 ( n3396 , n612 );
    or g518 ( n2271 , n1029 , n3049 );
    nor g519 ( n1113 , n2393 , n4127 );
    or g520 ( n4597 , n4014 , n5474 );
    and g521 ( n4256 , n3406 , n5962 );
    or g522 ( n3527 , n358 , n367 );
    or g523 ( n4063 , n3296 , n3638 );
    or g524 ( n6140 , n5485 , n1644 );
    and g525 ( n3639 , n1380 , n138 );
    and g526 ( n2002 , n5211 , n1530 );
    not g527 ( n1040 , n113 );
    and g528 ( n2437 , n5945 , n4215 );
    and g529 ( n3531 , n2863 , n2054 );
    not g530 ( n2610 , n2135 );
    or g531 ( n2937 , n142 , n3793 );
    nor g532 ( n2867 , n4344 , n939 );
    nor g533 ( n3097 , n1151 , n2391 );
    not g534 ( n4364 , n2020 );
    or g535 ( n625 , n6095 , n1145 );
    nor g536 ( n3419 , n5792 , n5996 );
    or g537 ( n6129 , n1193 , n3124 );
    or g538 ( n2227 , n808 , n408 );
    or g539 ( n6152 , n3123 , n1243 );
    not g540 ( n1099 , n5261 );
    not g541 ( n5492 , n1029 );
    nor g542 ( n5478 , n1080 , n3709 );
    and g543 ( n6112 , n2850 , n4998 );
    and g544 ( n2471 , n144 , n2487 );
    not g545 ( n2764 , n1603 );
    or g546 ( n1332 , n3845 , n1343 );
    not g547 ( n5104 , n480 );
    or g548 ( n1460 , n782 , n1589 );
    nor g549 ( n3516 , n2926 , n5689 );
    or g550 ( n4139 , n3507 , n756 );
    or g551 ( n2909 , n3104 , n2098 );
    and g552 ( n5728 , n2294 , n185 );
    and g553 ( n4053 , n1975 , n2343 );
    and g554 ( n2787 , n654 , n5027 );
    or g555 ( n1560 , n1297 , n4427 );
    not g556 ( n4892 , n6052 );
    and g557 ( n4391 , n1088 , n55 );
    nor g558 ( n4976 , n229 , n2078 );
    not g559 ( n5721 , n5293 );
    not g560 ( n2273 , n5691 );
    or g561 ( n3725 , n3869 , n3790 );
    or g562 ( n375 , n563 , n1101 );
    not g563 ( n5281 , n2797 );
    or g564 ( n4886 , n6282 , n1888 );
    nor g565 ( n2209 , n2850 , n4819 );
    and g566 ( n2180 , n767 , n5581 );
    and g567 ( n3817 , n1543 , n6018 );
    and g568 ( n5759 , n2995 , n1855 );
    or g569 ( n116 , n1169 , n3505 );
    or g570 ( n4884 , n554 , n1333 );
    or g571 ( n1644 , n555 , n4806 );
    or g572 ( n2524 , n6091 , n4149 );
    and g573 ( n832 , n492 , n2943 );
    and g574 ( n3544 , n98 , n5367 );
    not g575 ( n3734 , n2099 );
    and g576 ( n3743 , n5690 , n2800 );
    not g577 ( n3368 , n3466 );
    and g578 ( n6294 , n675 , n1686 );
    and g579 ( n321 , n5903 , n5699 );
    or g580 ( n4265 , n4386 , n6157 );
    not g581 ( n2033 , n1207 );
    and g582 ( n5173 , n5707 , n3928 );
    or g583 ( n705 , n4337 , n2079 );
    not g584 ( n5821 , n3426 );
    or g585 ( n3293 , n2497 , n973 );
    not g586 ( n3395 , n5011 );
    not g587 ( n863 , n5502 );
    not g588 ( n4281 , n3731 );
    nor g589 ( n1034 , n1048 , n2476 );
    or g590 ( n1069 , n947 , n2284 );
    not g591 ( n93 , n5686 );
    nor g592 ( n847 , n2658 , n3586 );
    nor g593 ( n4958 , n4135 , n2861 );
    nor g594 ( n5956 , n3089 , n513 );
    or g595 ( n2939 , n2395 , n5712 );
    not g596 ( n1874 , n929 );
    or g597 ( n3344 , n3203 , n542 );
    not g598 ( n1788 , n3523 );
    not g599 ( n2710 , n2666 );
    or g600 ( n5993 , n1231 , n2485 );
    not g601 ( n5865 , n2018 );
    or g602 ( n3315 , n3878 , n1539 );
    or g603 ( n196 , n372 , n15 );
    not g604 ( n956 , n4365 );
    or g605 ( n445 , n4888 , n3154 );
    not g606 ( n2032 , n4442 );
    nor g607 ( n6166 , n1820 , n5960 );
    or g608 ( n5866 , n2600 , n448 );
    not g609 ( n273 , n5099 );
    or g610 ( n4666 , n2419 , n4003 );
    or g611 ( n4786 , n198 , n1870 );
    or g612 ( n880 , n1413 , n1697 );
    not g613 ( n2266 , n1464 );
    or g614 ( n1975 , n2577 , n1768 );
    and g615 ( n4751 , n5230 , n4312 );
    not g616 ( n5026 , n1667 );
    or g617 ( n1776 , n5955 , n4526 );
    or g618 ( n5132 , n1400 , n652 );
    or g619 ( n5415 , n2659 , n6236 );
    not g620 ( n5771 , n3684 );
    or g621 ( n2125 , n4005 , n700 );
    not g622 ( n3579 , n2988 );
    not g623 ( n1125 , n2417 );
    not g624 ( n4398 , n4626 );
    or g625 ( n3962 , n268 , n3493 );
    not g626 ( n3795 , n3187 );
    nor g627 ( n5760 , n6176 , n4950 );
    and g628 ( n1419 , n2102 , n4648 );
    and g629 ( n2767 , n1065 , n2618 );
    not g630 ( n151 , n2767 );
    or g631 ( n4464 , n4111 , n2773 );
    and g632 ( n3885 , n2019 , n3895 );
    nor g633 ( n3099 , n4732 , n1600 );
    nor g634 ( n320 , n5378 , n5382 );
    and g635 ( n2153 , n3571 , n3401 );
    or g636 ( n3736 , n3554 , n2094 );
    or g637 ( n4877 , n1266 , n1610 );
    or g638 ( n5705 , n4662 , n2286 );
    or g639 ( n4778 , n4612 , n1079 );
    or g640 ( n1369 , n2153 , n947 );
    not g641 ( n60 , n1498 );
    and g642 ( n5555 , n2443 , n5464 );
    and g643 ( n285 , n3760 , n31 );
    and g644 ( n399 , n337 , n4510 );
    nor g645 ( n820 , n4633 , n3961 );
    not g646 ( n1627 , n1630 );
    not g647 ( n5091 , n6225 );
    not g648 ( n4846 , n4825 );
    or g649 ( n5301 , n5676 , n3695 );
    or g650 ( n2745 , n1251 , n884 );
    or g651 ( n3772 , n3955 , n4346 );
    and g652 ( n3606 , n3808 , n5323 );
    or g653 ( n4260 , n1572 , n4127 );
    or g654 ( n4173 , n3297 , n3678 );
    and g655 ( n4186 , n5356 , n2028 );
    not g656 ( n570 , n334 );
    or g657 ( n1148 , n5947 , n4077 );
    and g658 ( n5430 , n4106 , n594 );
    nor g659 ( n6064 , n3400 , n2556 );
    not g660 ( n268 , n3503 );
    not g661 ( n1986 , n4208 );
    not g662 ( n1909 , n2832 );
    and g663 ( n1582 , n5831 , n775 );
    or g664 ( n676 , n5753 , n6164 );
    not g665 ( n3437 , n3193 );
    or g666 ( n1542 , n5692 , n3804 );
    or g667 ( n3572 , n5848 , n3904 );
    not g668 ( n4327 , n4346 );
    and g669 ( n2759 , n3219 , n760 );
    or g670 ( n4798 , n5974 , n3351 );
    and g671 ( n5345 , n4001 , n39 );
    not g672 ( n1937 , n4283 );
    or g673 ( n2729 , n214 , n2514 );
    nor g674 ( n3649 , n572 , n6117 );
    or g675 ( n5471 , n4249 , n2629 );
    and g676 ( n4217 , n806 , n3504 );
    and g677 ( n1545 , n2981 , n3966 );
    not g678 ( n2753 , n3869 );
    and g679 ( n523 , n1960 , n6005 );
    nor g680 ( n1373 , n1140 , n3463 );
    and g681 ( n4753 , n745 , n1762 );
    or g682 ( n4668 , n3891 , n5880 );
    and g683 ( n852 , n1468 , n3957 );
    or g684 ( n6080 , n4930 , n455 );
    or g685 ( n3026 , n4953 , n5371 );
    or g686 ( n6259 , n1896 , n4122 );
    not g687 ( n1409 , n773 );
    nor g688 ( n712 , n1281 , n4840 );
    or g689 ( n1486 , n3273 , n4116 );
    nor g690 ( n2541 , n3352 , n163 );
    nor g691 ( n6062 , n5829 , n3103 );
    not g692 ( n3669 , n4605 );
    not g693 ( n3147 , n3298 );
    nor g694 ( n2892 , n374 , n4908 );
    not g695 ( n936 , n192 );
    and g696 ( n1458 , n2628 , n2705 );
    not g697 ( n1248 , n4353 );
    nor g698 ( n6102 , n4123 , n2089 );
    not g699 ( n5377 , n373 );
    and g700 ( n2425 , n2048 , n688 );
    not g701 ( n4570 , n1959 );
    nor g702 ( n4182 , n681 , n2089 );
    not g703 ( n3166 , n3664 );
    or g704 ( n4245 , n5995 , n3900 );
    or g705 ( n6180 , n2436 , n447 );
    not g706 ( n785 , n1834 );
    not g707 ( n2751 , n1527 );
    nor g708 ( n6063 , n1828 , n5133 );
    or g709 ( n4038 , n6144 , n3228 );
    nor g710 ( n2046 , n2967 , n3562 );
    not g711 ( n3509 , n4554 );
    and g712 ( n521 , n729 , n3308 );
    or g713 ( n4012 , n5362 , n1440 );
    and g714 ( n6221 , n5340 , n5665 );
    nor g715 ( n2991 , n3040 , n1134 );
    not g716 ( n892 , n260 );
    or g717 ( n2288 , n5781 , n5504 );
    not g718 ( n2129 , n1603 );
    nor g719 ( n4143 , n6051 , n4628 );
    and g720 ( n6198 , n5159 , n4713 );
    and g721 ( n6169 , n4565 , n5584 );
    or g722 ( n3095 , n2875 , n3946 );
    not g723 ( n3860 , n2732 );
    nor g724 ( n59 , n5297 , n2042 );
    and g725 ( n1906 , n3024 , n464 );
    or g726 ( n624 , n1774 , n1292 );
    not g727 ( n1918 , n1663 );
    and g728 ( n3851 , n2699 , n1954 );
    or g729 ( n1740 , n5797 , n5889 );
    and g730 ( n1866 , n6119 , n5496 );
    not g731 ( n2651 , n4651 );
    and g732 ( n1566 , n1574 , n5203 );
    not g733 ( n2570 , n825 );
    not g734 ( n1092 , n5150 );
    not g735 ( n3890 , n3235 );
    not g736 ( n2762 , n4842 );
    and g737 ( n5556 , n5674 , n5700 );
    not g738 ( n340 , n3723 );
    or g739 ( n2642 , n4992 , n3747 );
    not g740 ( n5268 , n1111 );
    nor g741 ( n2509 , n730 , n3661 );
    nor g742 ( n2038 , n2099 , n4949 );
    nor g743 ( n3306 , n1330 , n1249 );
    or g744 ( n2886 , n4379 , n2553 );
    or g745 ( n4410 , n738 , n2159 );
    and g746 ( n2190 , n4007 , n951 );
    or g747 ( n991 , n2847 , n3494 );
    and g748 ( n4215 , n6130 , n5566 );
    or g749 ( n5535 , n3111 , n375 );
    nor g750 ( n3800 , n1933 , n740 );
    or g751 ( n5374 , n4754 , n90 );
    nor g752 ( n818 , n3408 , n3850 );
    nor g753 ( n2545 , n2387 , n848 );
    or g754 ( n5166 , n4420 , n226 );
    and g755 ( n5444 , n1994 , n4824 );
    nor g756 ( n1659 , n494 , n5865 );
    or g757 ( n3420 , n3003 , n2526 );
    nor g758 ( n64 , n561 , n1280 );
    nor g759 ( n1366 , n2607 , n3465 );
    and g760 ( n5202 , n57 , n1842 );
    not g761 ( n3921 , n4278 );
    and g762 ( n1487 , n3890 , n98 );
    nor g763 ( n1733 , n4619 , n984 );
    not g764 ( n4252 , n2521 );
    not g765 ( n4781 , n3907 );
    and g766 ( n317 , n2416 , n5829 );
    not g767 ( n858 , n2499 );
    or g768 ( n2159 , n4284 , n2998 );
    or g769 ( n1691 , n5739 , n886 );
    or g770 ( n1375 , n3339 , n4004 );
    not g771 ( n4665 , n5129 );
    and g772 ( n3963 , n3338 , n2301 );
    not g773 ( n4595 , n1529 );
    and g774 ( n935 , n2983 , n5704 );
    not g775 ( n3156 , n5605 );
    not g776 ( n5322 , n1899 );
    nor g777 ( n433 , n1607 , n4204 );
    and g778 ( n2285 , n1990 , n3482 );
    or g779 ( n1732 , n1518 , n5633 );
    nor g780 ( n4103 , n45 , n1363 );
    not g781 ( n1367 , n4604 );
    and g782 ( n3613 , n3740 , n5823 );
    nor g783 ( n3264 , n2565 , n935 );
    not g784 ( n471 , n1255 );
    not g785 ( n4244 , n3006 );
    not g786 ( n3526 , n3074 );
    and g787 ( n3462 , n258 , n540 );
    not g788 ( n2911 , n32 );
    not g789 ( n984 , n2579 );
    not g790 ( n4709 , n6155 );
    or g791 ( n5143 , n905 , n2441 );
    nor g792 ( n6285 , n3360 , n3745 );
    not g793 ( n4002 , n3911 );
    and g794 ( n5305 , n4383 , n5503 );
    or g795 ( n3352 , n1054 , n1573 );
    or g796 ( n4074 , n5035 , n5123 );
    and g797 ( n2832 , n6166 , n2704 );
    nor g798 ( n709 , n5462 , n2251 );
    or g799 ( n1414 , n1657 , n579 );
    not g800 ( n2386 , n2883 );
    or g801 ( n4977 , n4419 , n4375 );
    not g802 ( n3250 , n4231 );
    nor g803 ( n156 , n3995 , n2221 );
    nor g804 ( n5060 , n3494 , n2364 );
    not g805 ( n5309 , n1563 );
    or g806 ( n623 , n2605 , n1567 );
    or g807 ( n5783 , n245 , n4022 );
    and g808 ( n1568 , n4311 , n5358 );
    not g809 ( n3667 , n5583 );
    not g810 ( n4737 , n4749 );
    not g811 ( n1952 , n5277 );
    or g812 ( n4955 , n2999 , n2591 );
    not g813 ( n228 , n5959 );
    or g814 ( n1742 , n4724 , n2683 );
    not g815 ( n673 , n2310 );
    not g816 ( n3580 , n711 );
    not g817 ( n490 , n5578 );
    and g818 ( n2958 , n6226 , n4835 );
    not g819 ( n5342 , n1717 );
    not g820 ( n5295 , n5252 );
    nor g821 ( n2384 , n5515 , n3467 );
    or g822 ( n3204 , n3894 , n3348 );
    or g823 ( n891 , n992 , n3399 );
    not g824 ( n5079 , n999 );
    not g825 ( n3188 , n1538 );
    and g826 ( n1292 , n3914 , n505 );
    not g827 ( n36 , n3063 );
    not g828 ( n4502 , n2579 );
    and g829 ( n147 , n2753 , n5505 );
    nor g830 ( n510 , n1447 , n5379 );
    not g831 ( n422 , n6195 );
    or g832 ( n5100 , n5135 , n4942 );
    and g833 ( n4638 , n4292 , n2120 );
    and g834 ( n3873 , n259 , n3519 );
    nor g835 ( n4897 , n370 , n5476 );
    and g836 ( n110 , n574 , n5172 );
    and g837 ( n5605 , n5167 , n6003 );
    nor g838 ( n4617 , n3240 , n1320 );
    and g839 ( n1103 , n6130 , n4265 );
    or g840 ( n2300 , n4324 , n831 );
    and g841 ( n3841 , n5673 , n5533 );
    not g842 ( n5973 , n4551 );
    or g843 ( n4622 , n5228 , n3789 );
    or g844 ( n3916 , n4154 , n960 );
    nor g845 ( n4682 , n2701 , n4791 );
    not g846 ( n4163 , n3394 );
    nor g847 ( n4621 , n1927 , n4107 );
    not g848 ( n3213 , n1166 );
    not g849 ( n3338 , n5102 );
    and g850 ( n2341 , n4418 , n3559 );
    or g851 ( n1445 , n151 , n2512 );
    or g852 ( n5260 , n3275 , n5587 );
    or g853 ( n5647 , n4247 , n5471 );
    or g854 ( n6005 , n4049 , n4536 );
    nor g855 ( n5786 , n2462 , n1118 );
    and g856 ( n3922 , n2903 , n2034 );
    not g857 ( n5058 , n3107 );
    nor g858 ( n674 , n5932 , n8 );
    or g859 ( n237 , n2621 , n6141 );
    not g860 ( n5739 , n3778 );
    nor g861 ( n2110 , n2215 , n2062 );
    nor g862 ( n1847 , n4581 , n916 );
    not g863 ( n3123 , n3798 );
    not g864 ( n1755 , n552 );
    not g865 ( n2115 , n1817 );
    or g866 ( n2005 , n4771 , n1967 );
    or g867 ( n5256 , n3178 , n3248 );
    not g868 ( n2954 , n2262 );
    or g869 ( n5735 , n2788 , n6023 );
    or g870 ( n4740 , n5430 , n5765 );
    and g871 ( n1111 , n2661 , n178 );
    and g872 ( n5498 , n341 , n2798 );
    not g873 ( n5293 , n6171 );
    or g874 ( n195 , n4436 , n385 );
    not g875 ( n1591 , n3918 );
    not g876 ( n2803 , n124 );
    or g877 ( n1341 , n895 , n3163 );
    or g878 ( n3416 , n6156 , n4530 );
    or g879 ( n2213 , n1638 , n5231 );
    or g880 ( n5683 , n2924 , n3310 );
    not g881 ( n3335 , n1771 );
    and g882 ( n2654 , n2218 , n3362 );
    or g883 ( n5817 , n1308 , n2898 );
    or g884 ( n4766 , n756 , n1932 );
    or g885 ( n4901 , n4098 , n3261 );
    not g886 ( n3759 , n2802 );
    and g887 ( n489 , n4980 , n3195 );
    not g888 ( n6091 , n2491 );
    nor g889 ( n3041 , n1238 , n1170 );
    nor g890 ( n1285 , n1864 , n40 );
    and g891 ( n779 , n1186 , n1201 );
    not g892 ( n1549 , n1554 );
    not g893 ( n2468 , n1162 );
    not g894 ( n2900 , n3858 );
    not g895 ( n3840 , n4242 );
    nor g896 ( n4960 , n4454 , n3219 );
    or g897 ( n3151 , n743 , n317 );
    or g898 ( n1074 , n1289 , n5732 );
    nor g899 ( n4774 , n2791 , n1795 );
    or g900 ( n1245 , n2744 , n547 );
    not g901 ( n1678 , n5975 );
    and g902 ( n4299 , n1775 , n1988 );
    nor g903 ( n3875 , n2415 , n433 );
    nor g904 ( n6240 , n5943 , n588 );
    and g905 ( n480 , n5942 , n3491 );
    or g906 ( n4817 , n5246 , n2888 );
    nor g907 ( n5845 , n249 , n3456 );
    or g908 ( n6256 , n2331 , n2780 );
    not g909 ( n182 , n2796 );
    not g910 ( n4947 , n5949 );
    not g911 ( n2069 , n1808 );
    not g912 ( n3111 , n5852 );
    not g913 ( n1388 , n4551 );
    or g914 ( n4348 , n4914 , n417 );
    nor g915 ( n5982 , n900 , n5117 );
    or g916 ( n509 , n2611 , n1638 );
    nor g917 ( n2639 , n2819 , n171 );
    or g918 ( n830 , n5614 , n3910 );
    and g919 ( n5921 , n1449 , n1899 );
    or g920 ( n2168 , n3621 , n3249 );
    not g921 ( n2369 , n4234 );
    and g922 ( n5355 , n1495 , n1929 );
    not g923 ( n4551 , n4710 );
    not g924 ( n3520 , n2423 );
    nor g925 ( n1752 , n1712 , n5840 );
    or g926 ( n3802 , n5907 , n5709 );
    and g927 ( n3821 , n3403 , n2579 );
    not g928 ( n6283 , n2752 );
    or g929 ( n243 , n5440 , n4326 );
    and g930 ( n5347 , n2912 , n4314 );
    and g931 ( n4250 , n5691 , n1741 );
    nor g932 ( n2348 , n5564 , n1883 );
    or g933 ( n2641 , n2882 , n1716 );
    nor g934 ( n74 , n2651 , n1709 );
    and g935 ( n2798 , n3749 , n3565 );
    not g936 ( n512 , n2112 );
    or g937 ( n4582 , n6293 , n5267 );
    not g938 ( n800 , n3349 );
    and g939 ( n2130 , n4938 , n2008 );
    and g940 ( n1132 , n3539 , n3774 );
    nor g941 ( n3598 , n4482 , n4630 );
    nor g942 ( n353 , n4207 , n6089 );
    or g943 ( n4023 , n3573 , n2289 );
    not g944 ( n572 , n5437 );
    not g945 ( n4436 , n1912 );
    and g946 ( n2026 , n6196 , n3480 );
    or g947 ( n560 , n2406 , n1691 );
    or g948 ( n112 , n2574 , n1392 );
    not g949 ( n2820 , n3681 );
    or g950 ( n2685 , n1993 , n2121 );
    or g951 ( n1588 , n4236 , n3619 );
    not g952 ( n3719 , n1995 );
    not g953 ( n4009 , n3667 );
    and g954 ( n551 , n1931 , n1115 );
    or g955 ( n3109 , n3237 , n694 );
    nor g956 ( n1826 , n2603 , n4048 );
    or g957 ( n3450 , n5184 , n2380 );
    and g958 ( n452 , n5603 , n3705 );
    and g959 ( n22 , n2544 , n197 );
    nor g960 ( n4257 , n1685 , n1110 );
    or g961 ( n441 , n1480 , n33 );
    not g962 ( n4136 , n5792 );
    not g963 ( n2766 , n30 );
    or g964 ( n5511 , n4695 , n1542 );
    or g965 ( n959 , n3618 , n4034 );
    or g966 ( n4490 , n4140 , n4124 );
    and g967 ( n6066 , n100 , n2381 );
    not g968 ( n6231 , n4854 );
    or g969 ( n3180 , n669 , n601 );
    and g970 ( n3813 , n5294 , n4327 );
    and g971 ( n1904 , n2442 , n5694 );
    nor g972 ( n6011 , n2030 , n3956 );
    or g973 ( n3693 , n1792 , n223 );
    and g974 ( n1323 , n365 , n3224 );
    and g975 ( n6197 , n5782 , n3206 );
    or g976 ( n2393 , n1623 , n1816 );
    and g977 ( n3740 , n3722 , n3927 );
    nor g978 ( n475 , n1514 , n993 );
    not g979 ( n3401 , n4367 );
    not g980 ( n4796 , n4100 );
    and g981 ( n49 , n5772 , n2339 );
    not g982 ( n2161 , n5689 );
    nor g983 ( n2172 , n1861 , n1005 );
    buf g984 ( n4352 , n3817 );
    or g985 ( n4934 , n685 , n3649 );
    nor g986 ( n4518 , n5950 , n1636 );
    nor g987 ( n1513 , n992 , n2100 );
    nor g988 ( n431 , n2638 , n3611 );
    not g989 ( n5909 , n5426 );
    not g990 ( n3479 , n5709 );
    or g991 ( n4878 , n5322 , n83 );
    and g992 ( n2997 , n3876 , n5698 );
    nor g993 ( n387 , n863 , n1424 );
    not g994 ( n4358 , n5558 );
    not g995 ( n904 , n2855 );
    not g996 ( n3551 , n5333 );
    or g997 ( n5284 , n2072 , n3383 );
    not g998 ( n1202 , n662 );
    not g999 ( n1805 , n3441 );
    or g1000 ( n2856 , n2996 , n5751 );
    not g1001 ( n4247 , n2247 );
    not g1002 ( n2381 , n6256 );
    nor g1003 ( n2596 , n6034 , n4796 );
    not g1004 ( n3215 , n2013 );
    nor g1005 ( n3121 , n1761 , n6132 );
    or g1006 ( n306 , n491 , n2429 );
    nor g1007 ( n4719 , n732 , n4610 );
    and g1008 ( n1478 , n1800 , n1051 );
    not g1009 ( n2267 , n2734 );
    nor g1010 ( n4080 , n5522 , n1506 );
    not g1011 ( n4266 , n991 );
    or g1012 ( n5692 , n5317 , n325 );
    or g1013 ( n4278 , n3580 , n4745 );
    nor g1014 ( n5778 , n5916 , n5374 );
    nor g1015 ( n1235 , n2878 , n3508 );
    or g1016 ( n4175 , n1876 , n6126 );
    or g1017 ( n2556 , n3872 , n530 );
    not g1018 ( n3750 , n5512 );
    not g1019 ( n5298 , n451 );
    and g1020 ( n4233 , n1754 , n2103 );
    or g1021 ( n4726 , n2440 , n5742 );
    not g1022 ( n6253 , n4402 );
    and g1023 ( n5798 , n5805 , n1245 );
    or g1024 ( n2529 , n89 , n5648 );
    not g1025 ( n1966 , n1821 );
    not g1026 ( n65 , n618 );
    nor g1027 ( n3003 , n6000 , n2002 );
    nor g1028 ( n4601 , n926 , n5473 );
    or g1029 ( n3722 , n892 , n1441 );
    or g1030 ( n5440 , n1218 , n3955 );
    and g1031 ( n2783 , n4778 , n1894 );
    not g1032 ( n5781 , n4910 );
    nor g1033 ( n6156 , n1670 , n2827 );
    or g1034 ( n3183 , n3091 , n2059 );
    or g1035 ( n46 , n2614 , n497 );
    nor g1036 ( n3083 , n2146 , n289 );
    not g1037 ( n4092 , n5555 );
    or g1038 ( n2435 , n4816 , n4756 );
    not g1039 ( n3887 , n2291 );
    or g1040 ( n2280 , n2976 , n2887 );
    or g1041 ( n5718 , n1764 , n5033 );
    not g1042 ( n5081 , n5819 );
    or g1043 ( n6033 , n2961 , n6044 );
    or g1044 ( n5312 , n5424 , n4496 );
    not g1045 ( n5516 , n3660 );
    nor g1046 ( n4121 , n1415 , n3647 );
    and g1047 ( n1166 , n3598 , n394 );
    or g1048 ( n1989 , n4823 , n5299 );
    and g1049 ( n1407 , n5285 , n3028 );
    or g1050 ( n5375 , n1805 , n4232 );
    or g1051 ( n4363 , n2215 , n5355 );
    not g1052 ( n1623 , n5813 );
    nor g1053 ( n1117 , n2085 , n845 );
    and g1054 ( n2367 , n5811 , n4306 );
    or g1055 ( n3757 , n5465 , n5783 );
    nor g1056 ( n3709 , n4503 , n2904 );
    nor g1057 ( n5916 , n2401 , n144 );
    nor g1058 ( n1221 , n180 , n4984 );
    and g1059 ( n2872 , n3333 , n4698 );
    or g1060 ( n4210 , n3643 , n4944 );
    or g1061 ( n3656 , n5877 , n5392 );
    nor g1062 ( n3371 , n1690 , n1971 );
    or g1063 ( n3556 , n3409 , n1552 );
    not g1064 ( n1751 , n1749 );
    or g1065 ( n386 , n2267 , n1920 );
    nor g1066 ( n2137 , n2109 , n6177 );
    nor g1067 ( n6007 , n4866 , n2907 );
    nor g1068 ( n354 , n3659 , n2012 );
    or g1069 ( n639 , n2836 , n5530 );
    and g1070 ( n6165 , n957 , n333 );
    nor g1071 ( n988 , n5885 , n6114 );
    or g1072 ( n1625 , n1494 , n6135 );
    or g1073 ( n1651 , n5795 , n6259 );
    and g1074 ( n4309 , n4109 , n3298 );
    or g1075 ( n1039 , n4538 , n3339 );
    or g1076 ( n5392 , n314 , n4907 );
    or g1077 ( n44 , n977 , n5259 );
    or g1078 ( n4468 , n1276 , n3352 );
    or g1079 ( n1368 , n3337 , n2280 );
    or g1080 ( n4159 , n4225 , n3208 );
    not g1081 ( n1530 , n873 );
    and g1082 ( n4754 , n3729 , n3437 );
    nor g1083 ( n794 , n1905 , n5572 );
    or g1084 ( n2402 , n6301 , n2871 );
    not g1085 ( n5584 , n4075 );
    or g1086 ( n1210 , n5956 , n2960 );
    or g1087 ( n3432 , n4196 , n5888 );
    nor g1088 ( n3762 , n4509 , n1444 );
    or g1089 ( n5240 , n1927 , n188 );
    nor g1090 ( n2838 , n5518 , n4105 );
    nor g1091 ( n2238 , n283 , n2597 );
    not g1092 ( n3679 , n413 );
    and g1093 ( n2239 , n2161 , n2185 );
    not g1094 ( n2931 , n5413 );
    not g1095 ( n4587 , n2047 );
    nor g1096 ( n5960 , n796 , n5307 );
    not g1097 ( n2632 , n6138 );
    nor g1098 ( n677 , n5 , n5839 );
    or g1099 ( n1794 , n3512 , n3126 );
    or g1100 ( n3973 , n670 , n5175 );
    nor g1101 ( n1390 , n1021 , n1970 );
    not g1102 ( n209 , n558 );
    not g1103 ( n656 , n4913 );
    and g1104 ( n5961 , n6115 , n1581 );
    and g1105 ( n3444 , n4174 , n4829 );
    not g1106 ( n3239 , n4911 );
    nor g1107 ( n134 , n5133 , n3707 );
    not g1108 ( n4234 , n3666 );
    not g1109 ( n1083 , n1836 );
    nor g1110 ( n561 , n987 , n5075 );
    or g1111 ( n4523 , n763 , n3008 );
    or g1112 ( n6300 , n101 , n4777 );
    or g1113 ( n6228 , n1937 , n862 );
    or g1114 ( n5046 , n6149 , n3795 );
    nor g1115 ( n2648 , n1420 , n2742 );
    or g1116 ( n2429 , n1766 , n3264 );
    nor g1117 ( n5428 , n4925 , n3819 );
    and g1118 ( n4129 , n85 , n850 );
    nor g1119 ( n2748 , n6053 , n875 );
    or g1120 ( n2337 , n2425 , n5921 );
    not g1121 ( n1741 , n1423 );
    not g1122 ( n1638 , n3260 );
    nor g1123 ( n2482 , n5484 , n5577 );
    and g1124 ( n2031 , n4913 , n297 );
    or g1125 ( n5590 , n2626 , n3811 );
    or g1126 ( n770 , n4969 , n1626 );
    not g1127 ( n4445 , n6128 );
    not g1128 ( n1553 , n5549 );
    and g1129 ( n1954 , n5766 , n5346 );
    and g1130 ( n394 , n5052 , n1998 );
    or g1131 ( n740 , n2782 , n203 );
    not g1132 ( n4104 , n3542 );
    not g1133 ( n3501 , n6300 );
    nor g1134 ( n6257 , n4380 , n412 );
    and g1135 ( n6123 , n3704 , n5877 );
    or g1136 ( n3076 , n1454 , n2368 );
    not g1137 ( n4828 , n2130 );
    or g1138 ( n3403 , n3785 , n4272 );
    nor g1139 ( n6043 , n3232 , n405 );
    or g1140 ( n631 , n4217 , n5093 );
    or g1141 ( n5989 , n715 , n866 );
    or g1142 ( n4273 , n826 , n3786 );
    not g1143 ( n769 , n6299 );
    not g1144 ( n937 , n6213 );
    nor g1145 ( n1729 , n3371 , n1504 );
    or g1146 ( n2746 , n346 , n1078 );
    not g1147 ( n4856 , n5792 );
    or g1148 ( n4193 , n1627 , n398 );
    not g1149 ( n3553 , n5604 );
    not g1150 ( n2765 , n4852 );
    or g1151 ( n290 , n3723 , n1052 );
    not g1152 ( n3225 , n4575 );
    not g1153 ( n3664 , n5733 );
    nor g1154 ( n358 , n5907 , n3421 );
    or g1155 ( n5219 , n3127 , n6133 );
    not g1156 ( n905 , n2559 );
    or g1157 ( n5725 , n4359 , n4293 );
    not g1158 ( n6054 , n1972 );
    not g1159 ( n2352 , n5172 );
    not g1160 ( n4229 , n2296 );
    nor g1161 ( n724 , n3415 , n5610 );
    or g1162 ( n3760 , n3170 , n4932 );
    not g1163 ( n4214 , n2091 );
    not g1164 ( n5062 , n1999 );
    or g1165 ( n2738 , n3020 , n1606 );
    not g1166 ( n1818 , n5659 );
    or g1167 ( n1467 , n4404 , n5847 );
    nor g1168 ( n3864 , n665 , n5070 );
    or g1169 ( n2255 , n687 , n1158 );
    nor g1170 ( n5589 , n6089 , n4572 );
    nor g1171 ( n2622 , n1902 , n6178 );
    not g1172 ( n985 , n2333 );
    not g1173 ( n169 , n3105 );
    not g1174 ( n2343 , n5031 );
    or g1175 ( n3070 , n4919 , n2155 );
    not g1176 ( n94 , n1052 );
    and g1177 ( n5634 , n5410 , n1890 );
    and g1178 ( n6177 , n3973 , n2781 );
    or g1179 ( n4860 , n1336 , n4540 );
    nor g1180 ( n4132 , n3204 , n2683 );
    nor g1181 ( n2284 , n373 , n6099 );
    nor g1182 ( n1597 , n2547 , n3954 );
    and g1183 ( n6143 , n2986 , n4619 );
    and g1184 ( n3919 , n5175 , n4571 );
    nor g1185 ( n3277 , n2365 , n295 );
    not g1186 ( n5237 , n3057 );
    not g1187 ( n4713 , n2301 );
    or g1188 ( n3822 , n1401 , n406 );
    and g1189 ( n542 , n5317 , n1612 );
    or g1190 ( n5672 , n3742 , n6171 );
    and g1191 ( n3895 , n1798 , n340 );
    not g1192 ( n5365 , n174 );
    or g1193 ( n1630 , n2369 , n4653 );
    or g1194 ( n4497 , n1004 , n1185 );
    and g1195 ( n4272 , n532 , n6303 );
    not g1196 ( n2496 , n5044 );
    or g1197 ( n2501 , n1099 , n4591 );
    not g1198 ( n4981 , n3717 );
    or g1199 ( n2693 , n560 , n1009 );
    not g1200 ( n1084 , n2114 );
    and g1201 ( n6265 , n1844 , n5466 );
    nor g1202 ( n2502 , n650 , n942 );
    and g1203 ( n754 , n2276 , n6208 );
    or g1204 ( n2407 , n1285 , n1274 );
    and g1205 ( n5755 , n3405 , n806 );
    or g1206 ( n3655 , n5901 , n2451 );
    and g1207 ( n886 , n4788 , n3691 );
    nor g1208 ( n1872 , n1144 , n4060 );
    nor g1209 ( n884 , n5645 , n3974 );
    not g1210 ( n2377 , n1883 );
    not g1211 ( n2519 , n481 );
    and g1212 ( n4566 , n3703 , n5681 );
    not g1213 ( n1156 , n4385 );
    nor g1214 ( n5756 , n3001 , n3579 );
    nor g1215 ( n2116 , n5448 , n5080 );
    not g1216 ( n2127 , n5370 );
    or g1217 ( n835 , n6237 , n3497 );
    not g1218 ( n3438 , n4391 );
    not g1219 ( n3546 , n3052 );
    nor g1220 ( n3877 , n665 , n3397 );
    and g1221 ( n1853 , n2014 , n3305 );
    not g1222 ( n5037 , n608 );
    nor g1223 ( n4471 , n1490 , n474 );
    not g1224 ( n1280 , n5563 );
    nor g1225 ( n5021 , n1942 , n3369 );
    nor g1226 ( n2663 , n5771 , n3252 );
    nor g1227 ( n3518 , n1081 , n2252 );
    nor g1228 ( n5200 , n1292 , n3357 );
    not g1229 ( n3105 , n4342 );
    and g1230 ( n216 , n2457 , n4713 );
    not g1231 ( n157 , n1809 );
    or g1232 ( n4195 , n3156 , n2717 );
    and g1233 ( n3476 , n5564 , n1374 );
    or g1234 ( n1420 , n2988 , n508 );
    or g1235 ( n1018 , n3409 , n3547 );
    not g1236 ( n1386 , n4077 );
    nor g1237 ( n1725 , n2017 , n425 );
    and g1238 ( n4333 , n3970 , n5283 );
    not g1239 ( n3680 , n169 );
    or g1240 ( n139 , n6082 , n1500 );
    not g1241 ( n508 , n253 );
    and g1242 ( n5843 , n3392 , n1460 );
    and g1243 ( n716 , n1188 , n3482 );
    nor g1244 ( n153 , n3200 , n1237 );
    and g1245 ( n3362 , n4201 , n4637 );
    and g1246 ( n3903 , n2568 , n1431 );
    and g1247 ( n4381 , n3934 , n5269 );
    or g1248 ( n995 , n5537 , n2376 );
    not g1249 ( n4045 , n5851 );
    or g1250 ( n5897 , n2939 , n5983 );
    and g1251 ( n323 , n6286 , n1446 );
    not g1252 ( n4773 , n1871 );
    not g1253 ( n4538 , n3380 );
    not g1254 ( n3914 , n1443 );
    not g1255 ( n3952 , n4233 );
    and g1256 ( n6103 , n4936 , n3369 );
    not g1257 ( n4598 , n4473 );
    nor g1258 ( n6110 , n2468 , n2411 );
    or g1259 ( n2702 , n360 , n5204 );
    or g1260 ( n3426 , n917 , n2077 );
    or g1261 ( n349 , n5476 , n4209 );
    or g1262 ( n1163 , n426 , n4230 );
    nor g1263 ( n3177 , n3073 , n1789 );
    and g1264 ( n4876 , n5161 , n5299 );
    not g1265 ( n1142 , n972 );
    and g1266 ( n3958 , n436 , n2915 );
    not g1267 ( n801 , n2177 );
    or g1268 ( n5619 , n3554 , n2053 );
    or g1269 ( n1722 , n4498 , n6162 );
    nor g1270 ( n1724 , n1076 , n3205 );
    not g1271 ( n2591 , n5211 );
    not g1272 ( n3281 , n5583 );
    nor g1273 ( n3867 , n3969 , n1026 );
    or g1274 ( n540 , n3202 , n518 );
    or g1275 ( n1338 , n5939 , n1569 );
    and g1276 ( n2664 , n4620 , n5522 );
    not g1277 ( n530 , n4266 );
    or g1278 ( n2613 , n3446 , n4864 );
    and g1279 ( n2725 , n3136 , n4761 );
    not g1280 ( n5702 , n887 );
    nor g1281 ( n4577 , n505 , n2385 );
    nor g1282 ( n915 , n587 , n1593 );
    nor g1283 ( n1933 , n5797 , n2179 );
    not g1284 ( n1189 , n3557 );
    nor g1285 ( n5823 , n1477 , n4779 );
    or g1286 ( n5196 , n826 , n1615 );
    and g1287 ( n2420 , n4408 , n5065 );
    not g1288 ( n342 , n1818 );
    not g1289 ( n4482 , n1246 );
    or g1290 ( n5229 , n3368 , n5710 );
    nor g1291 ( n1321 , n1734 , n2507 );
    not g1292 ( n355 , n1652 );
    and g1293 ( n97 , n569 , n1566 );
    or g1294 ( n68 , n72 , n4476 );
    not g1295 ( n1522 , n5883 );
    not g1296 ( n1797 , n4587 );
    not g1297 ( n3391 , n3174 );
    and g1298 ( n549 , n2837 , n3025 );
    or g1299 ( n1758 , n4605 , n5923 );
    or g1300 ( n4914 , n2095 , n3462 );
    not g1301 ( n239 , n2770 );
    not g1302 ( n5665 , n5992 );
    not g1303 ( n1329 , n6130 );
    or g1304 ( n3023 , n2807 , n455 );
    not g1305 ( n2145 , n4866 );
    and g1306 ( n2674 , n6056 , n284 );
    and g1307 ( n4568 , n5295 , n3728 );
    nor g1308 ( n1672 , n3748 , n2225 );
    or g1309 ( n1437 , n5531 , n3627 );
    nor g1310 ( n2594 , n2857 , n1 );
    not g1311 ( n392 , n5717 );
    or g1312 ( n1006 , n3286 , n3528 );
    not g1313 ( n2728 , n2633 );
    or g1314 ( n271 , n6068 , n3934 );
    nor g1315 ( n1133 , n1657 , n181 );
    not g1316 ( n5513 , n1314 );
    nor g1317 ( n3017 , n6203 , n3314 );
    or g1318 ( n3600 , n746 , n2011 );
    not g1319 ( n897 , n1407 );
    and g1320 ( n1355 , n5101 , n3034 );
    nor g1321 ( n3673 , n1997 , n1882 );
    and g1322 ( n1442 , n5526 , n2724 );
    and g1323 ( n2347 , n525 , n52 );
    and g1324 ( n1062 , n4308 , n1980 );
    nor g1325 ( n6060 , n1117 , n4537 );
    or g1326 ( n4712 , n3258 , n3147 );
    not g1327 ( n1781 , n3549 );
    or g1328 ( n3626 , n1525 , n622 );
    not g1329 ( n5005 , n768 );
    nor g1330 ( n2945 , n5971 , n5727 );
    not g1331 ( n2578 , n5036 );
    nor g1332 ( n3473 , n2004 , n2201 );
    or g1333 ( n1339 , n1105 , n1170 );
    not g1334 ( n3448 , n4060 );
    not g1335 ( n5090 , n3779 );
    not g1336 ( n2588 , n293 );
    and g1337 ( n3008 , n393 , n1624 );
    nor g1338 ( n4360 , n2080 , n2902 );
    and g1339 ( n314 , n4136 , n4833 );
    not g1340 ( n3770 , n538 );
    not g1341 ( n5685 , n1526 );
    not g1342 ( n5573 , n3968 );
    not g1343 ( n2893 , n2372 );
    and g1344 ( n3347 , n4061 , n1191 );
    and g1345 ( n2760 , n2069 , n1501 );
    and g1346 ( n4956 , n5144 , n364 );
    nor g1347 ( n4423 , n1877 , n3855 );
    or g1348 ( n5631 , n4166 , n326 );
    and g1349 ( n2470 , n3602 , n2124 );
    nor g1350 ( n275 , n475 , n1334 );
    and g1351 ( n4167 , n4878 , n5641 );
    nor g1352 ( n5879 , n5346 , n5932 );
    not g1353 ( n2508 , n3453 );
    or g1354 ( n569 , n434 , n5729 );
    not g1355 ( n5904 , n4276 );
    and g1356 ( n2433 , n1153 , n4954 );
    or g1357 ( n6045 , n454 , n1763 );
    nor g1358 ( n5019 , n5072 , n4077 );
    not g1359 ( n3393 , n4316 );
    nor g1360 ( n1146 , n5272 , n1263 );
    not g1361 ( n3441 , n5985 );
    and g1362 ( n4081 , n4795 , n5351 );
    not g1363 ( n2542 , n3452 );
    or g1364 ( n545 , n1852 , n4296 );
    or g1365 ( n165 , n5519 , n1218 );
    and g1366 ( n4852 , n1353 , n2270 );
    or g1367 ( n5290 , n3545 , n4988 );
    and g1368 ( n2351 , n1402 , n532 );
    nor g1369 ( n5388 , n512 , n5275 );
    or g1370 ( n341 , n2640 , n1303 );
    and g1371 ( n5396 , n2895 , n956 );
    not g1372 ( n3838 , n3951 );
    not g1373 ( n3793 , n5191 );
    or g1374 ( n1276 , n1666 , n1592 );
    not g1375 ( n2644 , n5342 );
    not g1376 ( n2873 , n2123 );
    nor g1377 ( n5454 , n618 , n6167 );
    not g1378 ( n5381 , n1671 );
    not g1379 ( n2434 , n2700 );
    nor g1380 ( n5158 , n3031 , n3828 );
    and g1381 ( n3984 , n2768 , n1507 );
    not g1382 ( n5505 , n616 );
    nor g1383 ( n3529 , n4640 , n2809 );
    nor g1384 ( n227 , n3799 , n6260 );
    not g1385 ( n4816 , n662 );
    or g1386 ( n808 , n5715 , n811 );
    and g1387 ( n5235 , n1331 , n2471 );
    or g1388 ( n940 , n4343 , n1916 );
    nor g1389 ( n2870 , n4041 , n1740 );
    nor g1390 ( n4031 , n438 , n6289 );
    or g1391 ( n194 , n2435 , n4549 );
    not g1392 ( n200 , n760 );
    not g1393 ( n1632 , n1417 );
    nor g1394 ( n1398 , n2337 , n3094 );
    or g1395 ( n5012 , n3106 , n3257 );
    or g1396 ( n419 , n5040 , n5452 );
    nor g1397 ( n722 , n744 , n4693 );
    and g1398 ( n3805 , n5910 , n707 );
    and g1399 ( n5880 , n4687 , n3225 );
    or g1400 ( n4306 , n1227 , n435 );
    not g1401 ( n1789 , n5014 );
    or g1402 ( n5954 , n5680 , n517 );
    not g1403 ( n3614 , n4593 );
    not g1404 ( n316 , n2508 );
    or g1405 ( n550 , n1640 , n1732 );
    or g1406 ( n4592 , n6295 , n4807 );
    and g1407 ( n1008 , n2776 , n4494 );
    and g1408 ( n1593 , n3273 , n4338 );
    nor g1409 ( n4654 , n2840 , n2996 );
    or g1410 ( n3319 , n2900 , n2242 );
    nor g1411 ( n6075 , n2532 , n4462 );
    not g1412 ( n1951 , n6108 );
    not g1413 ( n4899 , n3719 );
    nor g1414 ( n1948 , n6198 , n308 );
    not g1415 ( n5787 , n3593 );
    or g1416 ( n4669 , n4976 , n4846 );
    or g1417 ( n879 , n1133 , n5047 );
    not g1418 ( n55 , n755 );
    or g1419 ( n6099 , n596 , n108 );
    not g1420 ( n2406 , n3441 );
    or g1421 ( n2452 , n4616 , n2518 );
    nor g1422 ( n5407 , n4888 , n3573 );
    or g1423 ( n3718 , n4101 , n5715 );
    not g1424 ( n92 , n4886 );
    and g1425 ( n1634 , n5912 , n4872 );
    nor g1426 ( n4437 , n2146 , n1456 );
    or g1427 ( n351 , n2022 , n18 );
    or g1428 ( n802 , n2324 , n5609 );
    nor g1429 ( n5439 , n287 , n1694 );
    and g1430 ( n3630 , n457 , n4275 );
    not g1431 ( n5530 , n3751 );
    not g1432 ( n289 , n2551 );
    not g1433 ( n3199 , n5332 );
    nor g1434 ( n3738 , n1056 , n3938 );
    not g1435 ( n634 , n254 );
    not g1436 ( n4759 , n2746 );
    not g1437 ( n207 , n4631 );
    nor g1438 ( n2866 , n2758 , n6252 );
    not g1439 ( n1175 , n3275 );
    or g1440 ( n2064 , n3006 , n4733 );
    not g1441 ( n3575 , n591 );
    not g1442 ( n2287 , n3009 );
    or g1443 ( n875 , n1597 , n3023 );
    or g1444 ( n246 , n1944 , n5247 );
    not g1445 ( n4555 , n5930 );
    or g1446 ( n3925 , n1407 , n3384 );
    not g1447 ( n954 , n495 );
    not g1448 ( n1411 , n596 );
    nor g1449 ( n256 , n733 , n5493 );
    and g1450 ( n1721 , n4057 , n5641 );
    not g1451 ( n5617 , n3534 );
    not g1452 ( n5299 , n3690 );
    or g1453 ( n4527 , n2748 , n4377 );
    not g1454 ( n4131 , n1903 );
    or g1455 ( n629 , n1619 , n456 );
    or g1456 ( n2572 , n4303 , n869 );
    not g1457 ( n2782 , n2232 );
    not g1458 ( n2317 , n3279 );
    not g1459 ( n211 , n4454 );
    nor g1460 ( n640 , n236 , n2946 );
    not g1461 ( n5257 , n6255 );
    and g1462 ( n1089 , n3822 , n1464 );
    nor g1463 ( n3153 , n4335 , n4684 );
    not g1464 ( n4593 , n1623 );
    not g1465 ( n4414 , n1998 );
    or g1466 ( n765 , n2424 , n664 );
    and g1467 ( n2688 , n1277 , n2633 );
    and g1468 ( n4101 , n2513 , n2224 );
    not g1469 ( n691 , n4492 );
    and g1470 ( n3858 , n1810 , n3366 );
    or g1471 ( n1391 , n2743 , n4120 );
    nor g1472 ( n208 , n5448 , n244 );
    not g1473 ( n1198 , n5873 );
    not g1474 ( n127 , n5179 );
    nor g1475 ( n1647 , n2300 , n5335 );
    or g1476 ( n5891 , n3801 , n1252 );
    not g1477 ( n5978 , n5752 );
    nor g1478 ( n1943 , n2707 , n5585 );
    not g1479 ( n4612 , n1706 );
    or g1480 ( n3201 , n3266 , n5094 );
    nor g1481 ( n4216 , n4356 , n2862 );
    not g1482 ( n3666 , n3389 );
    and g1483 ( n4793 , n4040 , n4396 );
    and g1484 ( n272 , n907 , n4134 );
    nor g1485 ( n104 , n472 , n3091 );
    or g1486 ( n5967 , n3438 , n307 );
    not g1487 ( n4554 , n756 );
    and g1488 ( n5512 , n1298 , n479 );
    or g1489 ( n4635 , n3388 , n4011 );
    nor g1490 ( n3200 , n6283 , n4748 );
    not g1491 ( n2950 , n345 );
    nor g1492 ( n1875 , n837 , n2341 );
    and g1493 ( n2051 , n238 , n2505 );
    not g1494 ( n3487 , n617 );
    and g1495 ( n5842 , n3588 , n6091 );
    or g1496 ( n1067 , n4629 , n2086 );
    and g1497 ( n2042 , n645 , n491 );
    or g1498 ( n6289 , n892 , n3791 );
    not g1499 ( n3272 , n2095 );
    nor g1500 ( n77 , n5268 , n847 );
    nor g1501 ( n1354 , n752 , n2096 );
    not g1502 ( n1570 , n175 );
    and g1503 ( n2370 , n5498 , n4161 );
    not g1504 ( n5931 , n4823 );
    not g1505 ( n2432 , n424 );
    nor g1506 ( n6246 , n500 , n1773 );
    and g1507 ( n2231 , n105 , n3415 );
    and g1508 ( n4185 , n4764 , n3181 );
    and g1509 ( n1279 , n1511 , n850 );
    not g1510 ( n3154 , n2004 );
    not g1511 ( n5836 , n4369 );
    and g1512 ( n1603 , n470 , n4466 );
    or g1513 ( n1047 , n4745 , n1735 );
    nor g1514 ( n4891 , n1432 , n2483 );
    or g1515 ( n3263 , n1453 , n629 );
    not g1516 ( n113 , n2092 );
    not g1517 ( n3523 , n1915 );
    nor g1518 ( n3782 , n5731 , n4054 );
    and g1519 ( n1890 , n2158 , n919 );
    or g1520 ( n3091 , n1302 , n3739 );
    nor g1521 ( n1693 , n3728 , n554 );
    nor g1522 ( n3313 , n4754 , n1745 );
    not g1523 ( n544 , n3882 );
    or g1524 ( n3611 , n4687 , n4051 );
    not g1525 ( n1021 , n4458 );
    or g1526 ( n4841 , n3768 , n4210 );
    nor g1527 ( n88 , n1224 , n3350 );
    not g1528 ( n5928 , n193 );
    nor g1529 ( n95 , n2833 , n2548 );
    or g1530 ( n6236 , n319 , n396 );
    nor g1531 ( n4015 , n3059 , n5122 );
    or g1532 ( n1126 , n1717 , n772 );
    not g1533 ( n4820 , n6123 );
    not g1534 ( n4057 , n3578 );
    not g1535 ( n593 , n2797 );
    or g1536 ( n357 , n2600 , n3272 );
    or g1537 ( n4806 , n3697 , n2290 );
    nor g1538 ( n5384 , n5801 , n2388 );
    not g1539 ( n1768 , n6038 );
    nor g1540 ( n2389 , n1428 , n2978 );
    not g1541 ( n5064 , n5654 );
    and g1542 ( n845 , n3941 , n3807 );
    or g1543 ( n363 , n4472 , n713 );
    not g1544 ( n160 , n1965 );
    and g1545 ( n5549 , n912 , n3539 );
    not g1546 ( n2943 , n307 );
    and g1547 ( n3578 , n815 , n1878 );
    and g1548 ( n5837 , n3698 , n1947 );
    nor g1549 ( n1100 , n4240 , n809 );
    or g1550 ( n5116 , n2240 , n3513 );
    or g1551 ( n2 , n331 , n2249 );
    nor g1552 ( n528 , n1257 , n2140 );
    and g1553 ( n4571 , n2329 , n2174 );
    and g1554 ( n1283 , n5312 , n183 );
    and g1555 ( n4707 , n4068 , n5354 );
    and g1556 ( n470 , n5957 , n442 );
    not g1557 ( n4926 , n5241 );
    and g1558 ( n188 , n5814 , n5623 );
    not g1559 ( n6210 , n4215 );
    or g1560 ( n2322 , n2420 , n2303 );
    nor g1561 ( n2325 , n5892 , n1325 );
    nor g1562 ( n3558 , n2840 , n3543 );
    not g1563 ( n5437 , n1007 );
    nor g1564 ( n3788 , n148 , n950 );
    or g1565 ( n997 , n2135 , n3143 );
    nor g1566 ( n4949 , n1877 , n674 );
    not g1567 ( n2332 , n4486 );
    not g1568 ( n4238 , n2681 );
    or g1569 ( n2378 , n4858 , n2793 );
    nor g1570 ( n4640 , n3346 , n4394 );
    and g1571 ( n1728 , n4659 , n4683 );
    and g1572 ( n4277 , n3830 , n3629 );
    or g1573 ( n547 , n1432 , n2554 );
    not g1574 ( n3394 , n394 );
    or g1575 ( n3285 , n3912 , n4084 );
    nor g1576 ( n4105 , n4088 , n5462 );
    nor g1577 ( n2895 , n943 , n2177 );
    not g1578 ( n4169 , n807 );
    nor g1579 ( n2858 , n5813 , n1781 );
    and g1580 ( n3646 , n2842 , n4609 );
    or g1581 ( n3844 , n3825 , n680 );
    and g1582 ( n3862 , n175 , n158 );
    not g1583 ( n1965 , n1737 );
    and g1584 ( n2087 , n4342 , n2732 );
    or g1585 ( n3169 , n3622 , n4118 );
    not g1586 ( n1857 , n2970 );
    not g1587 ( n2329 , n2300 );
    not g1588 ( n4616 , n4277 );
    and g1589 ( n5711 , n5054 , n3730 );
    nor g1590 ( n3318 , n4145 , n2949 );
    or g1591 ( n3783 , n5126 , n1042 );
    not g1592 ( n2584 , n5772 );
    and g1593 ( n5330 , n1028 , n2178 );
    nor g1594 ( n3278 , n4785 , n2338 );
    not g1595 ( n3332 , n5174 );
    not g1596 ( n871 , n2311 );
    or g1597 ( n1012 , n5163 , n2512 );
    and g1598 ( n660 , n1311 , n3904 );
    or g1599 ( n4308 , n2651 , n2953 );
    and g1600 ( n3248 , n5209 , n6281 );
    not g1601 ( n2704 , n3164 );
    nor g1602 ( n5677 , n1953 , n5470 );
    or g1603 ( n1239 , n2686 , n141 );
    and g1604 ( n334 , n5461 , n1220 );
    not g1605 ( n2697 , n6059 );
    and g1606 ( n541 , n571 , n2404 );
    and g1607 ( n3586 , n3047 , n1469 );
    or g1608 ( n1384 , n673 , n242 );
    or g1609 ( n2665 , n5232 , n1487 );
    not g1610 ( n5319 , n3035 );
    nor g1611 ( n5499 , n6154 , n2336 );
    nor g1612 ( n1232 , n5387 , n4711 );
    and g1613 ( n3910 , n4839 , n937 );
    nor g1614 ( n3094 , n2989 , n4736 );
    or g1615 ( n4864 , n5933 , n1887 );
    and g1616 ( n2951 , n6294 , n940 );
    or g1617 ( n3390 , n3759 , n2373 );
    or g1618 ( n3127 , n43 , n1178 );
    not g1619 ( n5878 , n1289 );
    and g1620 ( n6201 , n4263 , n2000 );
    not g1621 ( n1371 , n2000 );
    nor g1622 ( n5832 , n3481 , n2646 );
    nor g1623 ( n952 , n4575 , n5670 );
    not g1624 ( n2979 , n2628 );
    or g1625 ( n5176 , n3607 , n170 );
    and g1626 ( n782 , n4388 , n4856 );
    and g1627 ( n3161 , n3935 , n2795 );
    or g1628 ( n581 , n5617 , n205 );
    and g1629 ( n2733 , n895 , n2563 );
    or g1630 ( n3748 , n2654 , n1190 );
    or g1631 ( n5157 , n644 , n1682 );
    nor g1632 ( n1259 , n2415 , n2920 );
    nor g1633 ( n2773 , n2894 , n4951 );
    not g1634 ( n3202 , n2340 );
    or g1635 ( n5503 , n4100 , n3546 );
    or g1636 ( n698 , n1061 , n4871 );
    not g1637 ( n76 , n4391 );
    not g1638 ( n3266 , n4435 );
    or g1639 ( n2066 , n2510 , n3211 );
    not g1640 ( n3150 , n4833 );
    or g1641 ( n4180 , n2491 , n3770 );
    not g1642 ( n5174 , n4275 );
    or g1643 ( n1345 , n4692 , n3386 );
    or g1644 ( n6170 , n4310 , n3557 );
    not g1645 ( n3685 , n2318 );
    and g1646 ( n1988 , n5432 , n5938 );
    nor g1647 ( n24 , n1968 , n4670 );
    or g1648 ( n3845 , n3720 , n215 );
    not g1649 ( n2047 , n3640 );
    nor g1650 ( n6179 , n2463 , n4859 );
    not g1651 ( n2530 , n3001 );
    not g1652 ( n3133 , n1438 );
    not g1653 ( n1171 , n3503 );
    not g1654 ( n2796 , n4618 );
    and g1655 ( n6295 , n993 , n1561 );
    and g1656 ( n2527 , n2297 , n2811 );
    nor g1657 ( n2445 , n2141 , n3788 );
    and g1658 ( n3684 , n5870 , n2766 );
    not g1659 ( n122 , n3859 );
    or g1660 ( n590 , n4262 , n1749 );
    or g1661 ( n4610 , n4993 , n942 );
    and g1662 ( n4561 , n1014 , n4131 );
    and g1663 ( n5014 , n300 , n35 );
    not g1664 ( n5761 , n3948 );
    not g1665 ( n2769 , n647 );
    not g1666 ( n2099 , n730 );
    nor g1667 ( n2672 , n241 , n5032 );
    nor g1668 ( n3198 , n6281 , n1010 );
    and g1669 ( n4399 , n1686 , n1345 );
    nor g1670 ( n5085 , n6144 , n1359 );
    not g1671 ( n5182 , n1157 );
    not g1672 ( n2626 , n3660 );
    and g1673 ( n977 , n1534 , n5230 );
    or g1674 ( n4034 , n5716 , n4558 );
    and g1675 ( n5285 , n3049 , n1637 );
    nor g1676 ( n3399 , n3157 , n3266 );
    and g1677 ( n2925 , n1328 , n999 );
    nor g1678 ( n4531 , n4289 , n4808 );
    and g1679 ( n3588 , n4977 , n3992 );
    not g1680 ( n1217 , n3195 );
    not g1681 ( n5925 , n1135 );
    nor g1682 ( n2727 , n6269 , n3816 );
    not g1683 ( n4225 , n3615 );
    nor g1684 ( n6132 , n3128 , n5222 );
    or g1685 ( n2523 , n5818 , n247 );
    or g1686 ( n1183 , n5955 , n5189 );
    or g1687 ( n3452 , n965 , n3244 );
    or g1688 ( n265 , n3639 , n2024 );
    or g1689 ( n308 , n3301 , n419 );
    nor g1690 ( n2726 , n2421 , n5872 );
    not g1691 ( n5997 , n2981 );
    and g1692 ( n5119 , n1246 , n4252 );
    and g1693 ( n737 , n1150 , n700 );
    nor g1694 ( n5183 , n25 , n5756 );
    not g1695 ( n4328 , n3448 );
    nor g1696 ( n3945 , n1760 , n4919 );
    nor g1697 ( n5593 , n2966 , n5013 );
    nor g1698 ( n4978 , n4838 , n3763 );
    or g1699 ( n726 , n1690 , n4162 );
    not g1700 ( n3951 , n4372 );
    not g1701 ( n3308 , n5638 );
    not g1702 ( n5263 , n2377 );
    not g1703 ( n1645 , n2315 );
    nor g1704 ( n1676 , n3681 , n1692 );
    or g1705 ( n5185 , n377 , n5435 );
    nor g1706 ( n6293 , n5467 , n1814 );
    and g1707 ( n924 , n4606 , n2262 );
    and g1708 ( n4334 , n2084 , n392 );
    not g1709 ( n4534 , n5252 );
    not g1710 ( n3369 , n2093 );
    or g1711 ( n2015 , n5112 , n4482 );
    nor g1712 ( n4157 , n4567 , n4522 );
    not g1713 ( n4355 , n4128 );
    and g1714 ( n3152 , n132 , n1348 );
    and g1715 ( n3271 , n2558 , n5816 );
    or g1716 ( n1335 , n2891 , n3930 );
    and g1717 ( n5481 , n22 , n2785 );
    not g1718 ( n3874 , n4452 );
    and g1719 ( n4896 , n637 , n4851 );
    or g1720 ( n4511 , n3469 , n2771 );
    or g1721 ( n3168 , n3870 , n2211 );
    nor g1722 ( n4576 , n608 , n3833 );
    or g1723 ( n2809 , n5914 , n202 );
    nor g1724 ( n2603 , n2265 , n5433 );
    or g1725 ( n2375 , n3138 , n4753 );
    not g1726 ( n2294 , n5818 );
    and g1727 ( n5459 , n4012 , n4071 );
    not g1728 ( n5390 , n1087 );
    not g1729 ( n3621 , n5160 );
    not g1730 ( n4918 , n5029 );
    or g1731 ( n1996 , n5464 , n5733 );
    or g1732 ( n4011 , n2709 , n5372 );
    nor g1733 ( n9 , n447 , n3214 );
    not g1734 ( n1224 , n3560 );
    nor g1735 ( n3710 , n3913 , n128 );
    and g1736 ( n1656 , n958 , n5850 );
    not g1737 ( n4767 , n1548 );
    nor g1738 ( n534 , n3422 , n931 );
    nor g1739 ( n3069 , n943 , n3525 );
    not g1740 ( n2599 , n693 );
    or g1741 ( n2059 , n4267 , n4594 );
    not g1742 ( n5162 , n4145 );
    not g1743 ( n5914 , n2681 );
    and g1744 ( n3905 , n2170 , n5604 );
    not g1745 ( n688 , n1484 );
    not g1746 ( n3367 , n1865 );
    not g1747 ( n576 , n5115 );
    and g1748 ( n161 , n3664 , n4881 );
    or g1749 ( n4122 , n311 , n5040 );
    nor g1750 ( n3284 , n5428 , n2261 );
    or g1751 ( n1985 , n2360 , n2829 );
    not g1752 ( n5646 , n1050 );
    not g1753 ( n5985 , n997 );
    or g1754 ( n1298 , n3048 , n70 );
    or g1755 ( n376 , n3519 , n624 );
    not g1756 ( n5291 , n1975 );
    nor g1757 ( n1968 , n18 , n1700 );
    not g1758 ( n1193 , n2498 );
    or g1759 ( n3587 , n3032 , n2917 );
    not g1760 ( n1896 , n4089 );
    nor g1761 ( n888 , n85 , n6261 );
    not g1762 ( n4378 , n2891 );
    nor g1763 ( n3175 , n760 , n6219 );
    not g1764 ( n989 , n2510 );
    nor g1765 ( n2964 , n3296 , n2756 );
    not g1766 ( n444 , n1971 );
    and g1767 ( n473 , n4623 , n5100 );
    or g1768 ( n5828 , n1496 , n1147 );
    or g1769 ( n947 , n2908 , n6205 );
    or g1770 ( n5172 , n69 , n1214 );
    and g1771 ( n2123 , n4337 , n792 );
    or g1772 ( n2723 , n5635 , n2028 );
    not g1773 ( n3505 , n1300 );
    not g1774 ( n3415 , n1898 );
    nor g1775 ( n4205 , n2634 , n1067 );
    nor g1776 ( n2356 , n2260 , n3634 );
    not g1777 ( n233 , n5537 );
    or g1778 ( n2948 , n4720 , n1138 );
    and g1779 ( n6057 , n4070 , n1287 );
    or g1780 ( n3274 , n4376 , n679 );
    not g1781 ( n866 , n4776 );
    not g1782 ( n128 , n2264 );
    not g1783 ( n3170 , n142 );
    or g1784 ( n3214 , n2436 , n5468 );
    or g1785 ( n3691 , n2369 , n4807 );
    or g1786 ( n173 , n4008 , n359 );
    not g1787 ( n3823 , n1079 );
    nor g1788 ( n2999 , n6128 , n6241 );
    or g1789 ( n430 , n4010 , n6176 );
    and g1790 ( n1869 , n5894 , n4623 );
    and g1791 ( n5500 , n1037 , n3669 );
    not g1792 ( n29 , n548 );
    or g1793 ( n1422 , n6241 , n1958 );
    nor g1794 ( n3997 , n2835 , n4465 );
    nor g1795 ( n604 , n369 , n1769 );
    or g1796 ( n5372 , n293 , n3850 );
    and g1797 ( n1669 , n1676 , n4829 );
    or g1798 ( n2868 , n26 , n5527 );
    not g1799 ( n2208 , n1391 );
    nor g1800 ( n4704 , n2997 , n3044 );
    and g1801 ( n865 , n2893 , n3022 );
    not g1802 ( n3824 , n4759 );
    not g1803 ( n2894 , n2403 );
    or g1804 ( n5455 , n1381 , n5454 );
    not g1805 ( n1589 , n6145 );
    not g1806 ( n1238 , n4524 );
    and g1807 ( n4316 , n659 , n1959 );
    not g1808 ( n1723 , n6143 );
    not g1809 ( n2968 , n4845 );
    nor g1810 ( n4861 , n281 , n3392 );
    not g1811 ( n5213 , n1578 );
    nor g1812 ( n3268 , n4046 , n3922 );
    not g1813 ( n3240 , n4358 );
    and g1814 ( n1764 , n3231 , n3653 );
    nor g1815 ( n4760 , n3519 , n5064 );
    nor g1816 ( n5186 , n2934 , n5107 );
    or g1817 ( n2171 , n2652 , n6100 );
    or g1818 ( n3513 , n6108 , n1977 );
    and g1819 ( n457 , n2190 , n1788 );
    nor g1820 ( n242 , n6010 , n5283 );
    and g1821 ( n1260 , n176 , n3333 );
    not g1822 ( n6144 , n4398 );
    not g1823 ( n920 , n2671 );
    not g1824 ( n900 , n1966 );
    not g1825 ( n1785 , n5106 );
    not g1826 ( n3615 , n1572 );
    not g1827 ( n1181 , n5624 );
    and g1828 ( n3043 , n1141 , n1180 );
    and g1829 ( n2160 , n1923 , n4892 );
    nor g1830 ( n4330 , n1820 , n4755 );
    not g1831 ( n2652 , n2554 );
    or g1832 ( n1660 , n289 , n96 );
    not g1833 ( n1648 , n1518 );
    nor g1834 ( n5572 , n720 , n3563 );
    or g1835 ( n1184 , n6177 , n3198 );
    nor g1836 ( n2181 , n2606 , n4837 );
    or g1837 ( n1673 , n3540 , n2147 );
    nor g1838 ( n5591 , n1381 , n3433 );
    or g1839 ( n1757 , n5094 , n3696 );
    or g1840 ( n2571 , n3340 , n5321 );
    not g1841 ( n2552 , n4260 );
    or g1842 ( n4556 , n4332 , n1370 );
    or g1843 ( n3404 , n2665 , n1338 );
    not g1844 ( n3764 , n2030 );
    nor g1845 ( n2976 , n4723 , n4002 );
    and g1846 ( n6258 , n5143 , n1664 );
    not g1847 ( n3972 , n445 );
    and g1848 ( n2735 , n4947 , n5292 );
    or g1849 ( n1005 , n5369 , n3661 );
    and g1850 ( n4803 , n1203 , n732 );
    nor g1851 ( n4730 , n2730 , n6233 );
    nor g1852 ( n620 , n4046 , n2786 );
    or g1853 ( n4927 , n3269 , n5364 );
    not g1854 ( n556 , n4432 );
    and g1855 ( n1845 , n5216 , n4752 );
    or g1856 ( n1629 , n2630 , n4463 );
    or g1857 ( n5402 , n1248 , n3675 );
    and g1858 ( n4620 , n3460 , n4528 );
    or g1859 ( n2918 , n736 , n1662 );
    nor g1860 ( n2392 , n1536 , n5266 );
    or g1861 ( n4875 , n5282 , n774 );
    and g1862 ( n5059 , n2083 , n3238 );
    or g1863 ( n4401 , n967 , n1493 );
    not g1864 ( n3791 , n2162 );
    nor g1865 ( n539 , n2505 , n1892 );
    not g1866 ( n4533 , n224 );
    not g1867 ( n4827 , n4427 );
    or g1868 ( n2474 , n1143 , n930 );
    or g1869 ( n6193 , n3063 , n3767 );
    and g1870 ( n762 , n3965 , n3074 );
    or g1871 ( n2995 , n2360 , n2166 );
    and g1872 ( n4911 , n2787 , n5878 );
    not g1873 ( n2891 , n6295 );
    nor g1874 ( n4424 , n1780 , n3302 );
    and g1875 ( n190 , n2071 , n6180 );
    nor g1876 ( n819 , n1256 , n3301 );
    not g1877 ( n6288 , n5883 );
    not g1878 ( n5138 , n3786 );
    and g1879 ( n3442 , n2236 , n3780 );
    and g1880 ( n1299 , n3963 , n4044 );
    or g1881 ( n2097 , n2129 , n4548 );
    or g1882 ( n2263 , n5666 , n21 );
    not g1883 ( n4376 , n2790 );
    not g1884 ( n1505 , n5773 );
    or g1885 ( n4625 , n1554 , n4197 );
    not g1886 ( n481 , n3155 );
    nor g1887 ( n4661 , n2420 , n635 );
    or g1888 ( n3460 , n742 , n1466 );
    not g1889 ( n5525 , n4268 );
    or g1890 ( n555 , n6066 , n5207 );
    nor g1891 ( n633 , n4898 , n2939 );
    not g1892 ( n2054 , n1514 );
    not g1893 ( n1990 , n4547 );
    and g1894 ( n5266 , n1289 , n4954 );
    not g1895 ( n4059 , n1728 );
    buf g1896 ( n3660 , n1550 );
    not g1897 ( n2154 , n865 );
    not g1898 ( n3940 , n3451 );
    not g1899 ( n4574 , n5155 );
    not g1900 ( n2682 , n2694 );
    nor g1901 ( n3785 , n1633 , n4828 );
    and g1902 ( n3869 , n844 , n4823 );
    or g1903 ( n4630 , n3427 , n449 );
    or g1904 ( n3412 , n4002 , n5250 );
    not g1905 ( n0 , n5480 );
    or g1906 ( n3631 , n4299 , n661 );
    not g1907 ( n1023 , n4009 );
    or g1908 ( n3550 , n2482 , n6229 );
    and g1909 ( n2842 , n4842 , n0 );
    not g1910 ( n2975 , n3117 );
    or g1911 ( n4221 , n1585 , n5657 );
    not g1912 ( n91 , n1604 );
    and g1913 ( n2619 , n3294 , n944 );
    and g1914 ( n4472 , n585 , n3514 );
    and g1915 ( n5564 , n3964 , n4383 );
    and g1916 ( n2901 , n102 , n3689 );
    not g1917 ( n2833 , n1483 );
    not g1918 ( n4825 , n2269 );
    not g1919 ( n2851 , n4358 );
    or g1920 ( n829 , n2854 , n5212 );
    not g1921 ( n6020 , n4487 );
    or g1922 ( n5217 , n3530 , n3516 );
    nor g1923 ( n343 , n232 , n3018 );
    or g1924 ( n5442 , n1167 , n6057 );
    not g1925 ( n69 , n3596 );
    nor g1926 ( n4344 , n988 , n4302 );
    not g1927 ( n4499 , n4571 );
    nor g1928 ( n4388 , n4338 , n980 );
    not g1929 ( n6249 , n5248 );
    or g1930 ( n292 , n5078 , n1973 );
    and g1931 ( n1735 , n983 , n6059 );
    or g1932 ( n941 , n1900 , n2807 );
    and g1933 ( n3633 , n2341 , n4104 );
    or g1934 ( n3455 , n4892 , n2422 );
    or g1935 ( n3634 , n5975 , n5886 );
    nor g1936 ( n2692 , n3861 , n2679 );
    nor g1937 ( n5541 , n2978 , n991 );
    or g1938 ( n893 , n5600 , n4822 );
    not g1939 ( n3683 , n3077 );
    or g1940 ( n2442 , n4616 , n3231 );
    and g1941 ( n5775 , n2747 , n3907 );
    or g1942 ( n6218 , n2617 , n6039 );
    and g1943 ( n1509 , n1677 , n4625 );
    not g1944 ( n1277 , n38 );
    and g1945 ( n3326 , n1416 , n3102 );
    and g1946 ( n772 , n2713 , n2845 );
    nor g1947 ( n315 , n2843 , n5278 );
    or g1948 ( n848 , n2237 , n6275 );
    or g1949 ( n5814 , n604 , n2584 );
    not g1950 ( n5690 , n1615 );
    and g1951 ( n2919 , n4290 , n5819 );
    not g1952 ( n2126 , n2638 );
    or g1953 ( n525 , n2139 , n5926 );
    not g1954 ( n3629 , n4251 );
    and g1955 ( n5043 , n2691 , n583 );
    or g1956 ( n2472 , n1727 , n4193 );
    and g1957 ( n3205 , n549 , n5332 );
    and g1958 ( n3948 , n4796 , n5450 );
    not g1959 ( n2562 , n3971 );
    nor g1960 ( n3346 , n3222 , n5976 );
    or g1961 ( n4690 , n702 , n2525 );
    nor g1962 ( n4831 , n2851 , n5897 );
    not g1963 ( n2874 , n2465 );
    or g1964 ( n3106 , n6174 , n2550 );
    or g1965 ( n5457 , n5862 , n4559 );
    and g1966 ( n2149 , n764 , n1214 );
    or g1967 ( n4486 , n5264 , n3563 );
    nor g1968 ( n2678 , n4339 , n101 );
    and g1969 ( n1430 , n5791 , n2701 );
    nor g1970 ( n5199 , n2656 , n3909 );
    not g1971 ( n4671 , n6105 );
    and g1972 ( n261 , n1296 , n2560 );
    not g1973 ( n6116 , n3991 );
    not g1974 ( n3565 , n3023 );
    not g1975 ( n6059 , n5952 );
    or g1976 ( n6019 , n547 , n3751 );
    nor g1977 ( n1867 , n5084 , n4412 );
    and g1978 ( n522 , n3254 , n5702 );
    or g1979 ( n2814 , n4906 , n3998 );
    nor g1980 ( n3261 , n4058 , n2413 );
    not g1981 ( n4965 , n4159 );
    not g1982 ( n788 , n3091 );
    not g1983 ( n4218 , n5904 );
    or g1984 ( n2401 , n4467 , n4346 );
    not g1985 ( n814 , n2729 );
    and g1986 ( n5128 , n682 , n3755 );
    and g1987 ( n3957 , n5036 , n3776 );
    and g1988 ( n5851 , n2118 , n3518 );
    or g1989 ( n4127 , n5489 , n2992 );
    not g1990 ( n1 , n2710 );
    or g1991 ( n5494 , n3702 , n2277 );
    nor g1992 ( n5841 , n3569 , n6030 );
    or g1993 ( n319 , n3233 , n947 );
    nor g1994 ( n4138 , n3353 , n344 );
    or g1995 ( n5421 , n3208 , n3445 );
    not g1996 ( n2391 , n1958 );
    not g1997 ( n3414 , n1909 );
    not g1998 ( n5475 , n963 );
    nor g1999 ( n5597 , n3164 , n1894 );
    nor g2000 ( n1027 , n971 , n5256 );
    or g2001 ( n1779 , n2385 , n6061 );
    and g2002 ( n3389 , n1928 , n1728 );
    not g2003 ( n4843 , n1196 );
    nor g2004 ( n2544 , n4093 , n3002 );
    or g2005 ( n40 , n2799 , n2935 );
    not g2006 ( n6224 , n4334 );
    or g2007 ( n3703 , n5208 , n2038 );
    nor g2008 ( n3917 , n5081 , n3442 );
    not g2009 ( n2448 , n5691 );
    or g2010 ( n4458 , n6092 , n3819 );
    not g2011 ( n3325 , n5557 );
    and g2012 ( n2611 , n1479 , n5961 );
    or g2013 ( n4389 , n6266 , n63 );
    and g2014 ( n364 , n5395 , n4757 );
    or g2015 ( n3351 , n4933 , n2795 );
    not g2016 ( n5204 , n1595 );
    or g2017 ( n928 , n6064 , n4941 );
    nor g2018 ( n4880 , n5249 , n4029 );
    not g2019 ( n461 , n1162 );
    or g2020 ( n1893 , n5786 , n4265 );
    not g2021 ( n3665 , n4312 );
    not g2022 ( n6079 , n1601 );
    not g2023 ( n4461 , n5208 );
    and g2024 ( n4287 , n3613 , n1750 );
    or g2025 ( n1275 , n4556 , n3576 );
    or g2026 ( n5872 , n207 , n4373 );
    or g2027 ( n663 , n5095 , n6206 );
    and g2028 ( n5819 , n4955 , n702 );
    or g2029 ( n1402 , n1410 , n4072 );
    or g2030 ( n5126 , n3744 , n5118 );
    nor g2031 ( n5811 , n4632 , n2258 );
    nor g2032 ( n2839 , n2804 , n1849 );
    or g2033 ( n1579 , n2234 , n1074 );
    and g2034 ( n2256 , n4770 , n4668 );
    or g2035 ( n4528 , n2210 , n592 );
    nor g2036 ( n4645 , n1335 , n4731 );
    not g2037 ( n5697 , n1114 );
    or g2038 ( n2587 , n5920 , n2248 );
    and g2039 ( n6078 , n3574 , n436 );
    or g2040 ( n1351 , n6172 , n4455 );
    or g2041 ( n1716 , n5436 , n5740 );
    and g2042 ( n4835 , n2825 , n2752 );
    not g2043 ( n3559 , n180 );
    not g2044 ( n1313 , n3761 );
    nor g2045 ( n2921 , n5137 , n5343 );
    and g2046 ( n3733 , n5398 , n152 );
    and g2047 ( n4631 , n4326 , n2950 );
    or g2048 ( n3585 , n293 , n338 );
    nor g2049 ( n685 , n184 , n5586 );
    not g2050 ( n5262 , n5515 );
    and g2051 ( n6234 , n5191 , n1362 );
    or g2052 ( n4443 , n5082 , n5448 );
    nor g2053 ( n4179 , n430 , n48 );
    and g2054 ( n4550 , n4304 , n2899 );
    not g2055 ( n4413 , n5858 );
    nor g2056 ( n4279 , n5860 , n5161 );
    nor g2057 ( n1010 , n5830 , n5069 );
    nor g2058 ( n5643 , n2937 , n493 );
    or g2059 ( n4979 , n5484 , n1579 );
    nor g2060 ( n3899 , n2734 , n3446 );
    or g2061 ( n710 , n2372 , n579 );
    nor g2062 ( n1715 , n3055 , n3625 );
    nor g2063 ( n6107 , n378 , n1334 );
    or g2064 ( n3203 , n5065 , n3082 );
    nor g2065 ( n2447 , n4395 , n5445 );
    nor g2066 ( n4284 , n4370 , n3338 );
    and g2067 ( n918 , n4571 , n469 );
    not g2068 ( n1251 , n4461 );
    nor g2069 ( n4485 , n6247 , n4091 );
    nor g2070 ( n2286 , n5989 , n1100 );
    not g2071 ( n4557 , n6251 );
    or g2072 ( n3918 , n4750 , n1121 );
    and g2073 ( n1983 , n2811 , n2163 );
    not g2074 ( n6245 , n3034 );
    or g2075 ( n958 , n3332 , n3380 );
    and g2076 ( n5746 , n5560 , n846 );
    or g2077 ( n4699 , n1124 , n1739 );
    or g2078 ( n6085 , n2206 , n2729 );
    or g2079 ( n6235 , n3240 , n5010 );
    not g2080 ( n978 , n5052 );
    or g2081 ( n715 , n2218 , n6141 );
    or g2082 ( n3708 , n787 , n2900 );
    or g2083 ( n1237 , n3918 , n879 );
    or g2084 ( n1363 , n4941 , n955 );
    or g2085 ( n2850 , n5869 , n303 );
    or g2086 ( n5409 , n5848 , n5440 );
    or g2087 ( n5722 , n5071 , n3839 );
    or g2088 ( n2222 , n460 , n5214 );
    or g2089 ( n400 , n5190 , n1091 );
    nor g2090 ( n2477 , n286 , n620 );
    not g2091 ( n2770 , n3220 );
    not g2092 ( n2008 , n5906 );
    not g2093 ( n3834 , n4925 );
    not g2094 ( n1169 , n3021 );
    not g2095 ( n1599 , n2022 );
    and g2096 ( n4588 , n1985 , n347 );
    or g2097 ( n2258 , n2063 , n1286 );
    or g2098 ( n2669 , n3545 , n6220 );
    and g2099 ( n5076 , n5438 , n1520 );
    not g2100 ( n6223 , n1670 );
    nor g2101 ( n6139 , n4164 , n220 );
    or g2102 ( n4183 , n1039 , n1663 );
    not g2103 ( n3275 , n5230 );
    and g2104 ( n1462 , n4501 , n4612 );
    nor g2105 ( n5201 , n3262 , n4530 );
    and g2106 ( n4532 , n3856 , n979 );
    nor g2107 ( n5344 , n4582 , n5562 );
    or g2108 ( n465 , n2585 , n4740 );
    or g2109 ( n3238 , n1808 , n1143 );
    and g2110 ( n2212 , n3645 , n5292 );
    or g2111 ( n5578 , n5451 , n2285 );
    and g2112 ( n4644 , n2602 , n5909 );
    and g2113 ( n3443 , n3109 , n3459 );
    nor g2114 ( n6292 , n3644 , n3079 );
    or g2115 ( n5522 , n4238 , n3706 );
    or g2116 ( n2504 , n5094 , n5779 );
    and g2117 ( n3645 , n1824 , n1903 );
    and g2118 ( n1214 , n5963 , n5566 );
    not g2119 ( n1829 , n459 );
    nor g2120 ( n4718 , n5659 , n3435 );
    or g2121 ( n5153 , n1804 , n1969 );
    and g2122 ( n5025 , n537 , n2997 );
    and g2123 ( n70 , n5095 , n4448 );
    and g2124 ( n413 , n1658 , n844 );
    not g2125 ( n5559 , n4539 );
    not g2126 ( n3988 , n758 );
    and g2127 ( n5532 , n3391 , n5506 );
    and g2128 ( n1176 , n2587 , n300 );
    or g2129 ( n3494 , n2448 , n266 );
    or g2130 ( n1879 , n4630 , n34 );
    not g2131 ( n1567 , n858 );
    nor g2132 ( n3173 , n3665 , n4787 );
    or g2133 ( n3116 , n4598 , n5978 );
    not g2134 ( n3110 , n2988 );
    and g2135 ( n4447 , n3067 , n6249 );
    or g2136 ( n3763 , n4508 , n1995 );
    not g2137 ( n627 , n125 );
    not g2138 ( n5955 , n3444 );
    or g2139 ( n2353 , n156 , n1430 );
    not g2140 ( n1399 , n4631 );
    not g2141 ( n4824 , n3815 );
    and g2142 ( n5316 , n5816 , n2943 );
    and g2143 ( n3560 , n507 , n972 );
    not g2144 ( n2679 , n4208 );
    not g2145 ( n5524 , n35 );
    not g2146 ( n974 , n109 );
    not g2147 ( n5508 , n351 );
    not g2148 ( n776 , n592 );
    nor g2149 ( n2933 , n1883 , n6280 );
    or g2150 ( n2590 , n1234 , n4863 );
    nor g2151 ( n3525 , n4050 , n158 );
    nor g2152 ( n1940 , n6235 , n1390 );
    nor g2153 ( n2323 , n5460 , n2272 );
    not g2154 ( n4341 , n4599 );
    and g2155 ( n3411 , n3431 , n138 );
    nor g2156 ( n6191 , n740 , n5124 );
    nor g2157 ( n3789 , n1087 , n3782 );
    or g2158 ( n57 , n4331 , n1525 );
    and g2159 ( n1058 , n1436 , n602 );
    or g2160 ( n2100 , n1329 , n703 );
    or g2161 ( n3985 , n2356 , n1129 );
    and g2162 ( n6302 , n5682 , n5583 );
    or g2163 ( n4321 , n1015 , n4175 );
    or g2164 ( n5520 , n4984 , n1531 );
    not g2165 ( n367 , n3941 );
    or g2166 ( n2830 , n3361 , n3367 );
    and g2167 ( n483 , n1034 , n5768 );
    or g2168 ( n1807 , n2039 , n3445 );
    or g2169 ( n2821 , n5412 , n6033 );
    not g2170 ( n775 , n4723 );
    not g2171 ( n1533 , n428 );
    and g2172 ( n1544 , n4247 , n5205 );
    not g2173 ( n5681 , n1172 );
    and g2174 ( n2000 , n3298 , n4539 );
    and g2175 ( n1912 , n1868 , n2344 );
    not g2176 ( n4337 , n3573 );
    or g2177 ( n983 , n5453 , n4638 );
    or g2178 ( n4830 , n1058 , n868 );
    and g2179 ( n5419 , n2166 , n5611 );
    and g2180 ( n1655 , n3135 , n696 );
    or g2181 ( n2957 , n853 , n1916 );
    not g2182 ( n4172 , n1247 );
    and g2183 ( n4240 , n4125 , n3167 );
    not g2184 ( n6158 , n4751 );
    and g2185 ( n4539 , n1293 , n4928 );
    and g2186 ( n2328 , n3322 , n2176 );
    and g2187 ( n4716 , n1111 , n4321 );
    or g2188 ( n2233 , n6052 , n5665 );
    or g2189 ( n4500 , n3553 , n510 );
    not g2190 ( n3534 , n5501 );
    and g2191 ( n2003 , n5465 , n5177 );
    or g2192 ( n4702 , n4964 , n453 );
    or g2193 ( n913 , n2085 , n4953 );
    or g2194 ( n1730 , n3001 , n2419 );
    or g2195 ( n5824 , n4686 , n5414 );
    or g2196 ( n5112 , n59 , n978 );
    not g2197 ( n6275 , n4853 );
    and g2198 ( n1205 , n3209 , n4508 );
    and g2199 ( n5308 , n3781 , n2650 );
    nor g2200 ( n329 , n649 , n4686 );
    nor g2201 ( n728 , n3400 , n3027 );
    nor g2202 ( n3280 , n3158 , n1553 );
    or g2203 ( n1042 , n2319 , n3851 );
    not g2204 ( n1895 , n1224 );
    or g2205 ( n374 , n4347 , n5455 );
    or g2206 ( n3854 , n4210 , n77 );
    nor g2207 ( n3265 , n1687 , n4521 );
    or g2208 ( n202 , n3403 , n2351 );
    nor g2209 ( n3827 , n2535 , n3128 );
    and g2210 ( n3034 , n4469 , n4246 );
    nor g2211 ( n5856 , n1914 , n3487 );
    or g2212 ( n5936 , n4346 , n1831 );
    or g2213 ( n3472 , n1654 , n4901 );
    or g2214 ( n5359 , n4021 , n5525 );
    nor g2215 ( n4680 , n1976 , n5919 );
    or g2216 ( n5243 , n1002 , n4078 );
    nor g2217 ( n4088 , n605 , n1015 );
    or g2218 ( n718 , n304 , n664 );
    or g2219 ( n684 , n348 , n4335 );
    not g2220 ( n1472 , n5363 );
    or g2221 ( n2473 , n3349 , n921 );
    not g2222 ( n350 , n4930 );
    nor g2223 ( n2121 , n1508 , n5729 );
    or g2224 ( n3847 , n2352 , n482 );
    not g2225 ( n3104 , n5752 );
    and g2226 ( n2772 , n6297 , n231 );
    not g2227 ( n5695 , n851 );
    nor g2228 ( n5253 , n4278 , n3735 );
    not g2229 ( n807 , n4569 );
    not g2230 ( n751 , n1397 );
    not g2231 ( n642 , n216 );
    and g2232 ( n4196 , n1919 , n1213 );
    and g2233 ( n2122 , n738 , n4370 );
    nor g2234 ( n5431 , n327 , n4099 );
    not g2235 ( n5254 , n3596 );
    or g2236 ( n1124 , n3666 , n4357 );
    or g2237 ( n5626 , n2169 , n666 );
    not g2238 ( n5890 , n1391 );
    or g2239 ( n3314 , n4209 , n5446 );
    and g2240 ( n3056 , n690 , n750 );
    not g2241 ( n491 , n5901 );
    not g2242 ( n1258 , n2975 );
    or g2243 ( n2691 , n1903 , n735 );
    or g2244 ( n4732 , n5801 , n5109 );
    not g2245 ( n3807 , n4599 );
    and g2246 ( n806 , n2317 , n1012 );
    and g2247 ( n1851 , n5068 , n750 );
    or g2248 ( n4285 , n1974 , n3045 );
    or g2249 ( n6133 , n3962 , n632 );
    not g2250 ( n4102 , n3417 );
    not g2251 ( n1800 , n1340 );
    or g2252 ( n4677 , n6246 , n84 );
    nor g2253 ( n4859 , n1295 , n4318 );
    not g2254 ( n682 , n5910 );
    or g2255 ( n4066 , n4197 , n4782 );
    and g2256 ( n2475 , n769 , n1262 );
    not g2257 ( n846 , n4347 );
    not g2258 ( n2410 , n5413 );
    not g2259 ( n4890 , n1845 );
    not g2260 ( n2681 , n3410 );
    or g2261 ( n1556 , n5703 , n539 );
    or g2262 ( n2533 , n1193 , n5057 );
    not g2263 ( n390 , n2111 );
    and g2264 ( n662 , n5761 , n683 );
    or g2265 ( n2333 , n4233 , n3357 );
    nor g2266 ( n450 , n5104 , n4701 );
    not g2267 ( n4590 , n6034 );
    nor g2268 ( n1071 , n3499 , n5544 );
    or g2269 ( n2855 , n5753 , n4522 );
    and g2270 ( n4618 , n3694 , n5878 );
    not g2271 ( n1186 , n1714 );
    nor g2272 ( n5635 , n1701 , n1383 );
    nor g2273 ( n2382 , n937 , n1902 );
    nor g2274 ( n5338 , n2363 , n5737 );
    or g2275 ( n4116 , n3714 , n343 );
    or g2276 ( n3804 , n3686 , n4301 );
    nor g2277 ( n247 , n4443 , n1408 );
    and g2278 ( n2072 , n3137 , n3322 );
    nor g2279 ( n653 , n927 , n3737 );
    not g2280 ( n3593 , n3494 );
    nor g2281 ( n3342 , n4108 , n1229 );
    nor g2282 ( n1692 , n1255 , n1637 );
    and g2283 ( n899 , n2865 , n2615 );
    or g2284 ( n6187 , n2698 , n274 );
    not g2285 ( n910 , n3322 );
    and g2286 ( n1308 , n3978 , n1258 );
    not g2287 ( n3339 , n137 );
    not g2288 ( n4505 , n1187 );
    not g2289 ( n999 , n3826 );
    nor g2290 ( n1746 , n5097 , n3420 );
    not g2291 ( n463 , n890 );
    or g2292 ( n1606 , n1221 , n4880 );
    nor g2293 ( n6042 , n5918 , n5487 );
    and g2294 ( n5604 , n155 , n4793 );
    nor g2295 ( n3574 , n5652 , n4216 );
    and g2296 ( n1641 , n3650 , n1906 );
    and g2297 ( n6094 , n3343 , n941 );
    not g2298 ( n5391 , n3756 );
    and g2299 ( n3087 , n3207 , n5441 );
    and g2300 ( n4385 , n3196 , n2361 );
    or g2301 ( n1015 , n373 , n2909 );
    not g2302 ( n1635 , n213 );
    and g2303 ( n6163 , n5337 , n4378 );
    or g2304 ( n4725 , n6147 , n1120 );
    not g2305 ( n1378 , n1935 );
    not g2306 ( n6090 , n366 );
    not g2307 ( n5714 , n3472 );
    nor g2308 ( n5941 , n4169 , n1166 );
    not g2309 ( n1397 , n4992 );
    or g2310 ( n2801 , n179 , n3897 );
    and g2311 ( n2355 , n2790 , n5995 );
    nor g2312 ( n3136 , n4589 , n1991 );
    or g2313 ( n4418 , n5314 , n3243 );
    and g2314 ( n5315 , n2682 , n4952 );
    nor g2315 ( n966 , n1888 , n6216 );
    or g2316 ( n1880 , n3486 , n397 );
    not g2317 ( n4106 , n3077 );
    and g2318 ( n5976 , n2315 , n5385 );
    and g2319 ( n5356 , n4464 , n1904 );
    or g2320 ( n5236 , n4654 , n5958 );
    nor g2321 ( n3176 , n3628 , n1517 );
    and g2322 ( n1546 , n5911 , n2434 );
    nor g2323 ( n294 , n159 , n5500 );
    nor g2324 ( n3515 , n1218 , n2950 );
    not g2325 ( n5077 , n37 );
    or g2326 ( n2282 , n1808 , n4168 );
    nor g2327 ( n5070 , n6231 , n5151 );
    not g2328 ( n1304 , n6241 );
    or g2329 ( n56 , n1013 , n2378 );
    or g2330 ( n727 , n4229 , n5767 );
    or g2331 ( n4783 , n1304 , n115 );
    nor g2332 ( n474 , n4260 , n678 );
    and g2333 ( n1314 , n5074 , n4331 );
    and g2334 ( n1870 , n1829 , n2836 );
    or g2335 ( n1639 , n533 , n418 );
    nor g2336 ( n123 , n4775 , n4576 );
    or g2337 ( n5650 , n3425 , n2901 );
    not g2338 ( n3345 , n591 );
    or g2339 ( n5044 , n152 , n1228 );
    not g2340 ( n3654 , n585 );
    not g2341 ( n1633 , n2250 );
    or g2342 ( n5241 , n6082 , n6193 );
    and g2343 ( n2694 , n2813 , n3237 );
    not g2344 ( n1664 , n4921 );
    nor g2345 ( n3591 , n1593 , n2818 );
    or g2346 ( n3908 , n287 , n1206 );
    or g2347 ( n5145 , n4578 , n4411 );
    and g2348 ( n4578 , n4970 , n2022 );
    or g2349 ( n2774 , n5295 , n382 );
    or g2350 ( n651 , n2466 , n5987 );
    or g2351 ( n4449 , n5972 , n1884 );
    and g2352 ( n703 , n4221 , n5807 );
    and g2353 ( n979 , n4459 , n1262 );
    not g2354 ( n3568 , n3836 );
    nor g2355 ( n4553 , n3142 , n1734 );
    and g2356 ( n4967 , n5834 , n2051 );
    or g2357 ( n3700 , n3575 , n328 );
    and g2358 ( n3387 , n217 , n1708 );
    or g2359 ( n3747 , n2189 , n2637 );
    not g2360 ( n5502 , n5930 );
    or g2361 ( n2853 , n5972 , n5735 );
    or g2362 ( n3752 , n3955 , n4155 );
    or g2363 ( n741 , n805 , n489 );
    nor g2364 ( n2743 , n1643 , n871 );
    or g2365 ( n4393 , n28 , n1851 );
    nor g2366 ( n4099 , n5363 , n2126 );
    and g2367 ( n1687 , n2803 , n714 );
    or g2368 ( n839 , n5234 , n5025 );
    or g2369 ( n3430 , n340 , n5145 );
    nor g2370 ( n3635 , n4720 , n2586 );
    or g2371 ( n3810 , n3498 , n5195 );
    or g2372 ( n2013 , n1085 , n5110 );
    or g2373 ( n2261 , n863 , n1350 );
    and g2374 ( n5950 , n2002 , n2327 );
    not g2375 ( n5948 , n1049 );
    nor g2376 ( n6280 , n856 , n5345 );
    or g2377 ( n2538 , n683 , n3546 );
    not g2378 ( n3480 , n4570 );
    or g2379 ( n972 , n3716 , n551 );
    or g2380 ( n3735 , n40 , n3359 );
    and g2381 ( n4362 , n2105 , n799 );
    or g2382 ( n3941 , n5907 , n2486 );
    not g2383 ( n3533 , n3582 );
    not g2384 ( n2218 , n798 );
    nor g2385 ( n5486 , n3155 , n5793 );
    not g2386 ( n3959 , n2546 );
    not g2387 ( n488 , n5559 );
    or g2388 ( n1032 , n1971 , n618 );
    nor g2389 ( n3603 , n3879 , n344 );
    nor g2390 ( n597 , n1587 , n3852 );
    not g2391 ( n4913 , n2528 );
    not g2392 ( n1459 , n1593 );
    or g2393 ( n2034 , n1744 , n5978 );
    not g2394 ( n5803 , n885 );
    not g2395 ( n738 , n5506 );
    or g2396 ( n1017 , n1824 , n324 );
    and g2397 ( n2969 , n5876 , n5938 );
    nor g2398 ( n4093 , n1125 , n3922 );
    or g2399 ( n4579 , n2680 , n1089 );
    or g2400 ( n6291 , n3932 , n4497 );
    or g2401 ( n3982 , n3227 , n1796 );
    or g2402 ( n874 , n948 , n5993 );
    or g2403 ( n1479 , n2832 , n3999 );
    or g2404 ( n4201 , n1671 , n1271 );
    nor g2405 ( n4188 , n5291 , n2212 );
    or g2406 ( n3636 , n731 , n1632 );
    and g2407 ( n5577 , n1846 , n5681 );
    nor g2408 ( n4329 , n2261 , n2867 );
    nor g2409 ( n950 , n5514 , n3251 );
    or g2410 ( n2737 , n4245 , n5649 );
    not g2411 ( n4763 , n4098 );
    not g2412 ( n2166 , n3910 );
    nor g2413 ( n3872 , n4442 , n543 );
    and g2414 ( n2177 , n5282 , n4615 );
    not g2415 ( n2905 , n1770 );
    or g2416 ( n5724 , n3015 , n2073 );
    or g2417 ( n1929 , n2594 , n3352 );
    and g2418 ( n2510 , n5226 , n240 );
    not g2419 ( n3797 , n4336 );
    not g2420 ( n3503 , n910 );
    or g2421 ( n197 , n4391 , n3477 );
    or g2422 ( n842 , n1690 , n2815 );
    nor g2423 ( n2852 , n2309 , n3663 );
    nor g2424 ( n2362 , n2668 , n4597 );
    nor g2425 ( n5794 , n5992 , n2923 );
    and g2426 ( n303 , n4333 , n221 );
    and g2427 ( n3364 , n790 , n1264 );
    nor g2428 ( n4673 , n2709 , n3652 );
    nor g2429 ( n2237 , n1465 , n2721 );
    or g2430 ( n5109 , n1238 , n1953 );
    or g2431 ( n4966 , n5984 , n841 );
    or g2432 ( n5664 , n4583 , n833 );
    not g2433 ( n1771 , n4278 );
    not g2434 ( n3861 , n6213 );
    or g2435 ( n397 , n5959 , n5067 );
    or g2436 ( n2813 , n4037 , n592 );
    not g2437 ( n1681 , n400 );
    not g2438 ( n4466 , n5205 );
    or g2439 ( n2200 , n883 , n1663 );
    nor g2440 ( n2493 , n1501 , n2144 );
    or g2441 ( n2439 , n4981 , n1368 );
    not g2442 ( n4675 , n2621 );
    or g2443 ( n3927 , n6010 , n503 );
    or g2444 ( n5644 , n1376 , n88 );
    and g2445 ( n1269 , n5341 , n4789 );
    not g2446 ( n4324 , n5496 );
    not g2447 ( n454 , n1910 );
    or g2448 ( n4001 , n5247 , n4663 );
    not g2449 ( n5975 , n1582 );
    or g2450 ( n1451 , n2148 , n614 );
    not g2451 ( n5501 , n5215 );
    or g2452 ( n3863 , n2824 , n4645 );
    or g2453 ( n5542 , n5858 , n1757 );
    or g2454 ( n3407 , n5009 , n2729 );
    nor g2455 ( n5793 , n286 , n2040 );
    not g2456 ( n3273 , n4833 );
    or g2457 ( n1688 , n350 , n6045 );
    or g2458 ( n1528 , n1911 , n1570 );
    and g2459 ( n6171 , n5318 , n3834 );
    or g2460 ( n580 , n3304 , n959 );
    not g2461 ( n427 , n1989 );
    nor g2462 ( n1035 , n2697 , n4507 );
    nor g2463 ( n3623 , n20 , n4557 );
    or g2464 ( n6148 , n1513 , n1093 );
    or g2465 ( n1706 , n146 , n4142 );
    and g2466 ( n1431 , n1375 , n5758 );
    and g2467 ( n4292 , n2893 , n5097 );
    or g2468 ( n43 , n5775 , n3177 );
    and g2469 ( n1476 , n4190 , n4853 );
    or g2470 ( n6222 , n2937 , n2026 );
    nor g2471 ( n881 , n5562 , n4360 );
    not g2472 ( n4473 , n2078 );
    not g2473 ( n6267 , n1102 );
    not g2474 ( n439 , n5728 );
    not g2475 ( n5588 , n5969 );
    and g2476 ( n6069 , n1617 , n3858 );
    nor g2477 ( n2388 , n4613 , n3295 );
    or g2478 ( n2631 , n531 , n2653 );
    not g2479 ( n2136 , n4355 );
    nor g2480 ( n186 , n2764 , n5988 );
    or g2481 ( n4903 , n5168 , n1112 );
    or g2482 ( n3843 , n1054 , n5242 );
    and g2483 ( n592 , n4567 , n5088 );
    not g2484 ( n1425 , n864 );
    not g2485 ( n2795 , n2321 );
    nor g2486 ( n199 , n353 , n1844 );
    or g2487 ( n1370 , n1813 , n5654 );
    not g2488 ( n5462 , n1111 );
    or g2489 ( n4274 , n1472 , n4366 );
    not g2490 ( n4048 , n5005 );
    not g2491 ( n2487 , n864 );
    nor g2492 ( n1473 , n3424 , n5754 );
    or g2493 ( n1029 , n1255 , n3723 );
    nor g2494 ( n26 , n578 , n939 );
    and g2495 ( n962 , n2131 , n1624 );
    or g2496 ( n2205 , n1038 , n1260 );
    not g2497 ( n3101 , n5103 );
    or g2498 ( n4506 , n6218 , n4903 );
    and g2499 ( n2537 , n3740 , n1161 );
    not g2500 ( n948 , n1770 );
    or g2501 ( n269 , n3135 , n1470 );
    and g2502 ( n1931 , n554 , n5127 );
    not g2503 ( n5645 , n3734 );
    nor g2504 ( n4969 , n824 , n2984 );
    or g2505 ( n4474 , n2578 , n3896 );
    not g2506 ( n5859 , n1571 );
    nor g2507 ( n3096 , n3763 , n2354 );
    or g2508 ( n4605 , n5580 , n1872 );
    or g2509 ( n1862 , n1874 , n1053 );
    not g2510 ( n4006 , n1355 );
    nor g2511 ( n3616 , n997 , n6159 );
    or g2512 ( n5007 , n3914 , n4074 );
    not g2513 ( n4746 , n1191 );
    not g2514 ( n883 , n4995 );
    not g2515 ( n4757 , n1774 );
    nor g2516 ( n4915 , n3995 , n4707 );
    nor g2517 ( n497 , n5011 , n3641 );
    and g2518 ( n4315 , n1711 , n2660 );
    not g2519 ( n1562 , n4533 );
    not g2520 ( n4470 , n5998 );
    and g2521 ( n6073 , n4945 , n814 );
    and g2522 ( n4340 , n4516 , n2532 );
    and g2523 ( n5197 , n2852 , n4421 );
    and g2524 ( n5246 , n695 , n2570 );
    or g2525 ( n1056 , n499 , n1200 );
    or g2526 ( n6047 , n3755 , n4932 );
    nor g2527 ( n812 , n278 , n4872 );
    or g2528 ( n203 , n5588 , n3847 );
    not g2529 ( n4212 , n3019 );
    or g2530 ( n251 , n3481 , n5284 );
    or g2531 ( n1317 , n4450 , n2230 );
    or g2532 ( n568 , n3647 , n3326 );
    not g2533 ( n3499 , n1241 );
    not g2534 ( n368 , n3535 );
    not g2535 ( n720 , n4726 );
    and g2536 ( n5927 , n4200 , n4491 );
    and g2537 ( n4909 , n5951 , n4910 );
    not g2538 ( n1115 , n5252 );
    or g2539 ( n3870 , n3795 , n1081 );
    not g2540 ( n3129 , n3061 );
    nor g2541 ( n5763 , n1032 , n5560 );
    or g2542 ( n2922 , n2132 , n3591 );
    or g2543 ( n167 , n4567 , n2855 );
    not g2544 ( n5877 , n2132 );
    and g2545 ( n2453 , n2204 , n3551 );
    or g2546 ( n5767 , n3827 , n3853 );
    or g2547 ( n3648 , n3763 , n4024 );
    or g2548 ( n3206 , n3993 , n5 );
    and g2549 ( n183 , n3216 , n233 );
    nor g2550 ( n1616 , n5573 , n5784 );
    nor g2551 ( n1590 , n2067 , n333 );
    or g2552 ( n1150 , n5967 , n2492 );
    not g2553 ( n5926 , n4929 );
    or g2554 ( n4912 , n5817 , n2880 );
    not g2555 ( n284 , n5985 );
    not g2556 ( n2698 , n146 );
    and g2557 ( n6077 , n5738 , n1582 );
    nor g2558 ( n1901 , n3780 , n2305 );
    nor g2559 ( n5550 , n253 , n1674 );
    or g2560 ( n3775 , n2070 , n3212 );
    not g2561 ( n5141 , n4303 );
    or g2562 ( n276 , n3646 , n2942 );
    or g2563 ( n4426 , n5745 , n1442 );
    not g2564 ( n689 , n2440 );
    nor g2565 ( n970 , n2389 , n961 );
    or g2566 ( n2305 , n5953 , n1043 );
    not g2567 ( n1882 , n798 );
    or g2568 ( n3435 , n3497 , n4309 );
    nor g2569 ( n6297 , n3417 , n4685 );
    and g2570 ( n1246 , n3035 , n3058 );
    or g2571 ( n753 , n1778 , n544 );
    not g2572 ( n3926 , n1743 );
    or g2573 ( n878 , n1863 , n97 );
    nor g2574 ( n2065 , n687 , n2401 );
    or g2575 ( n3632 , n4425 , n2113 );
    not g2576 ( n1382 , n3645 );
    not g2577 ( n4259 , n1216 );
    not g2578 ( n3219 , n101 );
    not g2579 ( n4288 , n4998 );
    nor g2580 ( n5937 , n3409 , n2749 );
    nor g2581 ( n4867 , n3279 , n6244 );
    and g2582 ( n5693 , n1546 , n2143 );
    nor g2583 ( n5406 , n3568 , n1575 );
    nor g2584 ( n4691 , n2789 , n2151 );
    or g2585 ( n4368 , n4850 , n2874 );
    or g2586 ( n1713 , n5176 , n631 );
    nor g2587 ( n4917 , n4152 , n3595 );
    nor g2588 ( n2865 , n5602 , n5136 );
    or g2589 ( n2397 , n4657 , n4627 );
    or g2590 ( n5049 , n2712 , n111 );
    or g2591 ( n5548 , n3542 , n6001 );
    not g2592 ( n5745 , n6201 );
    nor g2593 ( n5286 , n407 , n5603 );
    or g2594 ( n1839 , n1894 , n1018 );
    not g2595 ( n4670 , n6239 );
    not g2596 ( n3485 , n687 );
    not g2597 ( n3514 , n5711 );
    or g2598 ( n870 , n2399 , n4048 );
    nor g2599 ( n4325 , n1976 , n75 );
    nor g2600 ( n4055 , n6142 , n4802 );
    not g2601 ( n2815 , n1381 );
    not g2602 ( n2740 , n4605 );
    and g2603 ( n191 , n880 , n2630 );
    or g2604 ( n4462 , n1312 , n911 );
    nor g2605 ( n2736 , n2254 , n3961 );
    nor g2606 ( n3865 , n234 , n3076 );
    not g2607 ( n2847 , n1521 );
    not g2608 ( n3324 , n4495 );
    and g2609 ( n643 , n770 , n1497 );
    or g2610 ( n5515 , n1156 , n4181 );
    and g2611 ( n6212 , n4137 , n1046 );
    or g2612 ( n5087 , n147 , n1080 );
    not g2613 ( n4788 , n4490 );
    not g2614 ( n2216 , n2157 );
    or g2615 ( n3496 , n94 , n3192 );
    or g2616 ( n3504 , n4016 , n1445 );
    or g2617 ( n2450 , n5028 , n5693 );
    and g2618 ( n2025 , n3916 , n3022 );
    nor g2619 ( n4177 , n6011 , n5824 );
    and g2620 ( n798 , n486 , n3559 );
    not g2621 ( n4165 , n1226 );
    nor g2622 ( n3353 , n4677 , n4758 );
    and g2623 ( n2574 , n504 , n4911 );
    or g2624 ( n5164 , n5076 , n5838 );
    and g2625 ( n2515 , n3773 , n3606 );
    or g2626 ( n4547 , n1091 , n4028 );
    and g2627 ( n3191 , n4203 , n122 );
    not g2628 ( n3299 , n3895 );
    not g2629 ( n5636 , n1816 );
    nor g2630 ( n1145 , n623 , n1259 );
    nor g2631 ( n63 , n2228 , n3977 );
    nor g2632 ( n4198 , n4604 , n2423 );
    and g2633 ( n5628 , n5062 , n1760 );
    and g2634 ( n3483 , n5748 , n6195 );
    not g2635 ( n3372 , n657 );
    not g2636 ( n3124 , n3379 );
    not g2637 ( n2299 , n606 );
    not g2638 ( n5416 , n6198 );
    not g2639 ( n172 , n1563 );
    and g2640 ( n2372 , n5422 , n726 );
    or g2641 ( n1812 , n2808 , n3762 );
    nor g2642 ( n2844 , n2604 , n1398 );
    or g2643 ( n3445 , n4502 , n3924 );
    or g2644 ( n5991 , n152 , n2941 );
    not g2645 ( n787 , n5354 );
    or g2646 ( n6209 , n2495 , n3806 );
    nor g2647 ( n295 , n3853 , n4228 );
    not g2648 ( n3146 , n938 );
    or g2649 ( n6070 , n3146 , n2964 );
    nor g2650 ( n1160 , n2332 , n6169 );
    or g2651 ( n3329 , n251 , n3865 );
    nor g2652 ( n3970 , n321 , n4719 );
    nor g2653 ( n699 , n457 , n4521 );
    or g2654 ( n171 , n1556 , n5835 );
    not g2655 ( n1068 , n5700 );
    nor g2656 ( n5806 , n135 , n1418 );
    or g2657 ( n1426 , n831 , n5798 );
    or g2658 ( n1856 , n3335 , n1502 );
    or g2659 ( n5123 , n4577 , n82 );
    nor g2660 ( n1804 , n5192 , n1807 );
    not g2661 ( n6211 , n4971 );
    or g2662 ( n1209 , n2869 , n1859 );
    not g2663 ( n2418 , n784 );
    not g2664 ( n4987 , n4744 );
    not g2665 ( n4375 , n3214 );
    nor g2666 ( n6161 , n4894 , n440 );
    nor g2667 ( n4109 , n2580 , n236 );
    and g2668 ( n2761 , n1046 , n5258 );
    or g2669 ( n1928 , n4868 , n3996 );
    nor g2670 ( n2575 , n943 , n5282 );
    or g2671 ( n2117 , n6213 , n1723 );
    not g2672 ( n2277 , n4821 );
    and g2673 ( n862 , n1560 , n6111 );
    not g2674 ( n4657 , n4565 );
    nor g2675 ( n5427 , n1096 , n302 );
    not g2676 ( n734 , n1890 );
    or g2677 ( n3652 , n5778 , n3670 );
    and g2678 ( n2860 , n3118 , n1360 );
    not g2679 ( n4968 , n1996 );
    or g2680 ( n3704 , n4415 , n5996 );
    or g2681 ( n1141 , n4906 , n5604 );
    and g2682 ( n1130 , n5020 , n2660 );
    nor g2683 ( n3816 , n3162 , n6067 );
    or g2684 ( n6117 , n1282 , n5590 );
    not g2685 ( n6127 , n6154 );
    and g2686 ( n2561 , n759 , n5048 );
    or g2687 ( n3167 , n900 , n3753 );
    and g2688 ( n3468 , n624 , n4514 );
    not g2689 ( n177 , n4202 );
    or g2690 ( n5487 , n4642 , n6081 );
    nor g2691 ( n222 , n2537 , n6063 );
    not g2692 ( n4674 , n3689 );
    not g2693 ( n5611 , n1986 );
    or g2694 ( n2346 , n331 , n4226 );
    not g2695 ( n2555 , n443 );
    not g2696 ( n3964 , n2205 );
    or g2697 ( n4787 , n5692 , n1254 );
    not g2698 ( n811 , n1928 );
    not g2699 ( n3032 , n5670 );
    or g2700 ( n3165 , n5643 , n2021 );
    not g2701 ( n5641 , n1169 );
    or g2702 ( n5748 , n5683 , n6042 );
    not g2703 ( n4776 , n2199 );
    nor g2704 ( n4560 , n529 , n6018 );
    or g2705 ( n2195 , n4700 , n4368 );
    not g2706 ( n90 , n3043 );
    nor g2707 ( n511 , n4467 , n5936 );
    or g2708 ( n5447 , n5543 , n1332 );
    not g2709 ( n4818 , n813 );
    nor g2710 ( n3721 , n5127 , n5802 );
    or g2711 ( n4810 , n572 , n3050 );
    not g2712 ( n1033 , n3906 );
    and g2713 ( n3913 , n2408 , n5211 );
    and g2714 ( n1346 , n851 , n567 );
    and g2715 ( n6226 , n6253 , n4380 );
    nor g2716 ( n781 , n5351 , n6274 );
    or g2717 ( n1650 , n1897 , n3903 );
    not g2718 ( n908 , n5188 );
    nor g2719 ( n4322 , n3681 , n5095 );
    or g2720 ( n664 , n5809 , n4328 );
    and g2721 ( n229 , n1382 , n5461 );
    or g2722 ( n4509 , n1549 , n3490 );
    or g2723 ( n869 , n6053 , n5314 );
    nor g2724 ( n1884 , n1688 , n2727 );
    or g2725 ( n2001 , n5859 , n5325 );
    not g2726 ( n5616 , n4045 );
    or g2727 ( n2517 , n1838 , n162 );
    or g2728 ( n4491 , n3953 , n4313 );
    and g2729 ( n4882 , n1533 , n1319 );
    or g2730 ( n671 , n5407 , n3972 );
    or g2731 ( n1406 , n411 , n3329 );
    or g2732 ( n4943 , n952 , n1645 );
    or g2733 ( n391 , n519 , n1235 );
    or g2734 ( n2315 , n4575 , n3846 );
    or g2735 ( n3115 , n3743 , n4474 );
    and g2736 ( n4422 , n570 , n4947 );
    nor g2737 ( n1535 , n5624 , n1164 );
    not g2738 ( n4721 , n1669 );
    or g2739 ( n33 , n6062 , n2186 );
    or g2740 ( n4420 , n3202 , n710 );
    or g2741 ( n4029 , n4260 , n5898 );
    not g2742 ( n2557 , n5796 );
    nor g2743 ( n1658 , n3690 , n3327 );
    nor g2744 ( n2485 , n1309 , n5796 );
    not g2745 ( n3798 , n1776 );
    nor g2746 ( n805 , n2299 , n5859 );
    not g2747 ( n1697 , n5136 );
    and g2748 ( n5491 , n828 , n4614 );
    nor g2749 ( n1072 , n5813 , n4647 );
    not g2750 ( n85 , n1509 );
    not g2751 ( n2191 , n2000 );
    or g2752 ( n5959 , n1220 , n2703 );
    and g2753 ( n3583 , n5976 , n55 );
    and g2754 ( n565 , n6145 , n1085 );
    and g2755 ( n2265 , n3269 , n1643 );
    not g2756 ( n6219 , n4777 );
    not g2757 ( n1076 , n1464 );
    or g2758 ( n1806 , n213 , n708 );
    not g2759 ( n3330 , n3509 );
    nor g2760 ( n5272 , n3667 , n5800 );
    not g2761 ( n1731 , n4057 );
    not g2762 ( n4782 , n2087 );
    not g2763 ( n2045 , n3731 );
    not g2764 ( n5558 , n3633 );
    and g2765 ( n5627 , n1858 , n2081 );
    nor g2766 ( n423 , n1943 , n4377 );
    or g2767 ( n4453 , n677 , n1475 );
    not g2768 ( n665 , n1433 );
    and g2769 ( n3778 , n4342 , n6211 );
    or g2770 ( n690 , n2082 , n5350 );
    or g2771 ( n3675 , n4579 , n4095 );
    nor g2772 ( n5776 , n5964 , n4664 );
    or g2773 ( n1520 , n4747 , n5042 );
    nor g2774 ( n149 , n1547 , n5981 );
    nor g2775 ( n3595 , n2243 , n1283 );
    or g2776 ( n589 , n5940 , n441 );
    not g2777 ( n2757 , n462 );
    nor g2778 ( n487 , n4392 , n3802 );
    not g2779 ( n2486 , n3140 );
    or g2780 ( n5674 , n2216 , n5232 );
    and g2781 ( n4998 , n5554 , n758 );
    or g2782 ( n1842 , n4331 , n2318 );
    and g2783 ( n5073 , n4147 , n1611 );
    not g2784 ( n1926 , n2706 );
    not g2785 ( n3920 , n6157 );
    or g2786 ( n5030 , n407 , n1625 );
    or g2787 ( n1506 , n5595 , n4624 );
    or g2788 ( n5179 , n1240 , n4307 );
    nor g2789 ( n636 , n3971 , n4315 );
    and g2790 ( n4298 , n4811 , n6222 );
    or g2791 ( n4133 , n5157 , n4055 );
    or g2792 ( n1294 , n2010 , n1148 );
    or g2793 ( n5656 , n3501 , n2759 );
    not g2794 ( n1485 , n1451 );
    not g2795 ( n3130 , n2969 );
    or g2796 ( n5514 , n2308 , n10 );
    nor g2797 ( n4685 , n2849 , n5737 );
    not g2798 ( n4030 , n3042 );
    or g2799 ( n5949 , n5521 , n4432 );
    or g2800 ( n5932 , n3107 , n5273 );
    and g2801 ( n370 , n1264 , n1825 );
    or g2802 ( n2141 , n1738 , n4407 );
    nor g2803 ( n2494 , n5701 , n404 );
    or g2804 ( n108 , n4175 , n903 );
    nor g2805 ( n1848 , n1608 , n400 );
    nor g2806 ( n2368 , n3648 , n881 );
    not g2807 ( n965 , n5842 );
    not g2808 ( n4983 , n3195 );
    and g2809 ( n15 , n4431 , n1462 );
    or g2810 ( n5417 , n4016 , n1307 );
    and g2811 ( n2959 , n4503 , n5970 );
    and g2812 ( n797 , n5153 , n5396 );
    or g2813 ( n3521 , n1865 , n2632 );
    not g2814 ( n5935 , n1488 );
    or g2815 ( n2109 , n6119 , n6008 );
    not g2816 ( n2666 , n1533 );
    or g2817 ( n4734 , n5200 , n1294 );
    or g2818 ( n2229 , n3680 , n2403 );
    nor g2819 ( n4525 , n5883 , n3143 );
    buf g2820 ( n1421 , n5509 );
    or g2821 ( n6276 , n1555 , n1292 );
    not g2822 ( n1868 , n763 );
    and g2823 ( n3190 , n4401 , n4590 );
    not g2824 ( n3408 , n5769 );
    not g2825 ( n2220 , n1131 );
    and g2826 ( n3333 , n4989 , n717 );
    not g2827 ( n4242 , n1612 );
    or g2828 ( n4190 , n6088 , n3121 );
    or g2829 ( n5373 , n2396 , n5620 );
    not g2830 ( n6003 , n1356 );
    nor g2831 ( n1236 , n4933 , n2685 );
    not g2832 ( n5045 , n3955 );
    or g2833 ( n1097 , n1562 , n5653 );
    and g2834 ( n850 , n3778 , n1342 );
    nor g2835 ( n3470 , n2400 , n1275 );
    not g2836 ( n217 , n2765 );
    and g2837 ( n1554 , n3558 , n2483 );
    and g2838 ( n4134 , n4025 , n3683 );
    and g2839 ( n1011 , n5546 , n4493 );
    or g2840 ( n5327 , n1790 , n5265 );
    nor g2841 ( n5622 , n1888 , n3683 );
    or g2842 ( n6251 , n4676 , n4729 );
    and g2843 ( n6271 , n4963 , n6221 );
    or g2844 ( n3713 , n3249 , n4573 );
    or g2845 ( n3989 , n792 , n379 );
    or g2846 ( n2518 , n2608 , n4971 );
    and g2847 ( n1666 , n6069 , n3276 );
    or g2848 ( n266 , n3345 , n1815 );
    or g2849 ( n2379 , n2261 , n2868 );
    nor g2850 ( n5483 , n6182 , n3522 );
    or g2851 ( n5561 , n3344 , n5713 );
    not g2852 ( n1992 , n6066 );
    or g2853 ( n404 , n3141 , n391 );
    and g2854 ( n1004 , n4817 , n1595 );
    not g2855 ( n5040 , n5945 );
    and g2856 ( n3943 , n120 , n1711 );
    not g2857 ( n5203 , n1993 );
    not g2858 ( n5477 , n2242 );
    not g2859 ( n478 , n5393 );
    and g2860 ( n1147 , n4133 , n3157 );
    not g2861 ( n4313 , n1417 );
    not g2862 ( n1080 , n2916 );
    and g2863 ( n4076 , n2745 , n322 );
    and g2864 ( n2732 , n4697 , n4898 );
    and g2865 ( n3803 , n5672 , n3640 );
    or g2866 ( n5912 , n5974 , n2877 );
    not g2867 ( n5188 , n4835 );
    not g2868 ( n1708 , n5962 );
    and g2869 ( n3322 , n4889 , n2434 );
    not g2870 ( n10 , n904 );
    and g2871 ( n1671 , n6207 , n180 );
    buf g2872 ( n584 , n5509 );
    or g2873 ( n3678 , n3906 , n5315 );
    or g2874 ( n3771 , n4431 , n74 );
    not g2875 ( n3933 , n3181 );
    nor g2876 ( n401 , n1603 , n2875 );
    and g2877 ( n3060 , n1225 , n5991 );
    or g2878 ( n446 , n1621 , n1544 );
    not g2879 ( n5563 , n3977 );
    not g2880 ( n5545 , n529 );
    or g2881 ( n5709 , n3421 , n500 );
    or g2882 ( n3971 , n1016 , n4119 );
    not g2883 ( n2416 , n4162 );
    or g2884 ( n1333 , n3721 , n2515 );
    nor g2885 ( n3866 , n1052 , n2714 );
    not g2886 ( n5538 , n6090 );
    not g2887 ( n3730 , n2563 );
    nor g2888 ( n578 , n3578 , n4302 );
    nor g2889 ( n4070 , n1020 , n2902 );
    not g2890 ( n5468 , n587 );
    nor g2891 ( n1908 , n51 , n5012 );
    or g2892 ( n4255 , n6087 , n996 );
    nor g2893 ( n1372 , n4159 , n637 );
    not g2894 ( n5366 , n5031 );
    not g2895 ( n5476 , n4788 );
    nor g2896 ( n4689 , n1237 , n5569 );
    or g2897 ( n1753 , n686 , n5092 );
    and g2898 ( n2546 , n2386 , n3048 );
    or g2899 ( n3478 , n3417 , n1006 );
    not g2900 ( n4676 , n3859 );
    nor g2901 ( n3067 , n2142 , n2596 );
    and g2902 ( n3543 , n2652 , n3681 );
    not g2903 ( n447 , n3396 );
    not g2904 ( n2014 , n2760 );
    and g2905 ( n2883 , n3325 , n3723 );
    not g2906 ( n472 , n1267 );
    or g2907 ( n6071 , n303 , n2046 );
    nor g2908 ( n3889 , n6031 , n5659 );
    not g2909 ( n3243 , n426 );
    not g2910 ( n3765 , n3771 );
    and g2911 ( n3237 , n5568 , n5285 );
    not g2912 ( n4519 , n3608 );
    or g2913 ( n1024 , n2124 , n3610 );
    or g2914 ( n5720 , n3174 , n2122 );
    nor g2915 ( n405 , n520 , n4363 );
    not g2916 ( n2483 , n2836 );
    and g2917 ( n615 , n53 , n5396 );
    or g2918 ( n2812 , n114 , n5790 );
    or g2919 ( n3571 , n4113 , n1491 );
    not g2920 ( n4656 , n3700 );
    or g2921 ( n4253 , n3348 , n3161 );
    not g2922 ( n4752 , n4737 );
    nor g2923 ( n3086 , n4440 , n5210 );
    or g2924 ( n2248 , n4961 , n2357 );
    nor g2925 ( n4791 , n977 , n1618 );
    not g2926 ( n155 , n3919 );
    nor g2927 ( n1055 , n1953 , n4603 );
    and g2928 ( n4623 , n3038 , n19 );
    nor g2929 ( n27 , n4436 , n3556 );
    not g2930 ( n2503 , n6096 );
    or g2931 ( n756 , n4058 , n4015 );
    not g2932 ( n3160 , n4413 );
    not g2933 ( n731 , n6143 );
    or g2934 ( n1344 , n1720 , n170 );
    not g2935 ( n5493 , n1509 );
    and g2936 ( n2633 , n5592 , n3079 );
    or g2937 ( n1455 , n2954 , n1982 );
    or g2938 ( n4335 , n586 , n3824 );
    not g2939 ( n5974 , n660 );
    or g2940 ( n1541 , n1891 , n5291 );
    not g2941 ( n4614 , n5857 );
    or g2942 ( n6266 , n5696 , n1414 );
    not g2943 ( n1802 , n3307 );
    nor g2944 ( n5335 , n2539 , n5175 );
    nor g2945 ( n2489 , n2582 , n2694 );
    nor g2946 ( n2558 , n3180 , n1049 );
    or g2947 ( n1138 , n4338 , n1577 );
    or g2948 ( n906 , n3999 , n4585 );
    not g2949 ( n313 , n4081 );
    not g2950 ( n5292 , n2577 );
    not g2951 ( n6035 , n1220 );
    not g2952 ( n513 , n1512 );
    not g2953 ( n159 , n2986 );
    or g2954 ( n4290 , n4810 , n3919 );
    and g2955 ( n1070 , n2007 , n4495 );
    not g2956 ( n3836 , n6181 );
    and g2957 ( n2111 , n1278 , n4614 );
    and g2958 ( n4710 , n543 , n4809 );
    or g2959 ( n6182 , n6299 , n6055 );
    nor g2960 ( n6199 , n4168 , n1313 );
    nor g2961 ( n6044 , n1797 , n5762 );
    not g2962 ( n3507 , n2846 );
    or g2963 ( n3792 , n268 , n3769 );
    not g2964 ( n4653 , n4381 );
    nor g2965 ( n1642 , n5333 , n2938 );
    and g2966 ( n3720 , n6283 , n5555 );
    not g2967 ( n2600 , n3849 );
    or g2968 ( n3731 , n1888 , n534 );
    not g2969 ( n3754 , n5276 );
    or g2970 ( n3321 , n4626 , n2074 );
    not g2971 ( n1118 , n5757 );
    not g2972 ( n6238 , n918 );
    buf g2973 ( n2120 , n4422 );
    not g2974 ( n2781 , n831 );
    not g2975 ( n2675 , n1420 );
    and g2976 ( n2276 , n627 , n1267 );
    not g2977 ( n3502 , n5995 );
    or g2978 ( n1653 , n4699 , n153 );
    not g2979 ( n3063 , n4550 );
    nor g2980 ( n5833 , n3447 , n1846 );
    not g2981 ( n23 , n3133 );
    not g2982 ( n4149 , n1548 );
    not g2983 ( n3990 , n5309 );
    or g2984 ( n5411 , n871 , n1856 );
    nor g2985 ( n2459 , n1821 , n2616 );
    not g2986 ( n4044 , n5506 );
    not g2987 ( n5103 , n5634 );
    or g2988 ( n2411 , n6121 , n5408 );
    not g2989 ( n949 , n2763 );
    not g2990 ( n6111 , n1854 );
    not g2991 ( n1050 , n4644 );
    or g2992 ( n6076 , n3338 , n817 );
    or g2993 ( n4232 , n3270 , n2452 );
    not g2994 ( n5160 , n5391 );
    or g2995 ( n4366 , n784 , n5018 );
    nor g2996 ( n2156 , n5049 , n2447 );
    and g2997 ( n4696 , n727 , n231 );
    not g2998 ( n2635 , n3299 );
    or g2999 ( n14 , n4899 , n1209 );
    or g3000 ( n1969 , n2624 , n3622 );
    and g3001 ( n4440 , n1196 , n2458 );
    nor g3002 ( n1331 , n4786 , n1167 );
    nor g3003 ( n4973 , n2989 , n5429 );
    not g3004 ( n5275 , n2072 );
    not g3005 ( n2020 , n4060 );
    nor g3006 ( n3696 , n621 , n3590 );
    nor g3007 ( n5198 , n512 , n4199 );
    nor g3008 ( n5341 , n4562 , n924 );
    and g3009 ( n1036 , n753 , n5412 );
    or g3010 ( n4963 , n3102 , n5679 );
    or g3011 ( n2230 , n309 , n2892 );
    not g3012 ( n2224 , n345 );
    and g3013 ( n1598 , n6212 , n1967 );
    not g3014 ( n3846 , n327 );
    or g3015 ( n3547 , n6150 , n4523 );
    or g3016 ( n5379 , n4287 , n302 );
    or g3017 ( n1219 , n556 , n2138 );
    and g3018 ( n3701 , n5791 , n849 );
    not g3019 ( n61 , n1870 );
    and g3020 ( n3582 , n4315 , n5339 );
    nor g3021 ( n973 , n6017 , n5844 );
    nor g3022 ( n4724 , n5694 , n3244 );
    not g3023 ( n3171 , n3871 );
    or g3024 ( n5066 , n5741 , n5626 );
    nor g3025 ( n1614 , n4058 , n2259 );
    not g3026 ( n5789 , n1142 );
    or g3027 ( n596 , n3586 , n3356 );
    or g3028 ( n4384 , n5810 , n2642 );
    nor g3029 ( n2426 , n637 , n5872 );
    or g3030 ( n2334 , n2876 , n5304 );
    or g3031 ( n2155 , n3733 , n1291 );
    not g3032 ( n5370 , n1021 );
    or g3033 ( n4211 , n4746 , n5478 );
    not g3034 ( n6262 , n5893 );
    not g3035 ( n2075 , n1446 );
    not g3036 ( n5346 , n4406 );
    not g3037 ( n5565 , n455 );
    or g3038 ( n4857 , n1123 , n119 );
    not g3039 ( n1123 , n6113 );
    not g3040 ( n4563 , n5963 );
    and g3041 ( n5560 , n5686 , n6167 );
    and g3042 ( n1810 , n4480 , n1703 );
    and g3043 ( n1743 , n1035 , n2120 );
    and g3044 ( n4944 , n3016 , n178 );
    not g3045 ( n1941 , n2759 );
    or g3046 ( n6058 , n1540 , n2106 );
    not g3047 ( n2219 , n3632 );
    not g3048 ( n3305 , n3761 );
    and g3049 ( n5221 , n2481 , n3859 );
    or g3050 ( n815 , n5852 , n701 );
    and g3051 ( n4848 , n5699 , n1187 );
    or g3052 ( n3178 , n2076 , n171 );
    or g3053 ( n5016 , n834 , n1109 );
    and g3054 ( n4071 , n2381 , n5700 );
    and g3055 ( n986 , n217 , n1434 );
    or g3056 ( n2749 , n4294 , n5051 );
    or g3057 ( n2576 , n319 , n1719 );
    not g3058 ( n1228 , n3030 );
    not g3059 ( n3189 , n212 );
    or g3060 ( n5015 , n523 , n5016 );
    not g3061 ( n6010 , n37 );
    not g3062 ( n2340 , n6181 );
    or g3063 ( n3380 , n5420 , n3302 );
    not g3064 ( n2897 , n5433 );
    not g3065 ( n4051 , n5438 );
    or g3066 ( n6287 , n3672 , n4622 );
    not g3067 ( n2547 , n4418 );
    not g3068 ( n1336 , n4451 );
    not g3069 ( n2007 , n3577 );
    or g3070 ( n5088 , n1668 , n5536 );
    nor g3071 ( n5987 , n2405 , n234 );
    not g3072 ( n2863 , n3733 );
    and g3073 ( n5531 , n275 , n4334 );
    or g3074 ( n467 , n471 , n130 );
    and g3075 ( n695 , n5825 , n1980 );
    and g3076 ( n5065 , n4708 , n5022 );
    and g3077 ( n5397 , n3411 , n5475 );
    or g3078 ( n5971 , n5322 , n1335 );
    not g3079 ( n3300 , n1216 );
    not g3080 ( n2236 , n2174 );
    or g3081 ( n5679 , n535 , n1940 );
    and g3082 ( n6014 , n3376 , n3258 );
    nor g3083 ( n3085 , n4716 , n3854 );
    not g3084 ( n3965 , n127 );
    or g3085 ( n3978 , n6102 , n3334 );
    nor g3086 ( n163 , n2666 , n2323 );
    or g3087 ( n326 , n4037 , n5536 );
    nor g3088 ( n5966 , n2528 , n2715 );
    or g3089 ( n622 , n4027 , n2536 );
    not g3090 ( n5579 , n2980 );
    nor g3091 ( n2974 , n3632 , n4013 );
    not g3092 ( n4747 , n2806 );
    not g3093 ( n494 , n3364 );
    nor g3094 ( n223 , n266 , n2364 );
    or g3095 ( n3464 , n978 , n1584 );
    nor g3096 ( n4354 , n4615 , n1515 );
    not g3097 ( n5809 , n1423 );
    nor g3098 ( n976 , n2808 , n1474 );
    nor g3099 ( n2549 , n966 , n1303 );
    not g3100 ( n3046 , n1266 );
    and g3101 ( n2522 , n1107 , n2533 );
    nor g3102 ( n4986 , n3061 , n1714 );
    not g3103 ( n1841 , n1187 );
    and g3104 ( n3357 , n5155 , n2103 );
    not g3105 ( n3057 , n521 );
    not g3106 ( n4202 , n532 );
    and g3107 ( n4513 , n3284 , n4458 );
    nor g3108 ( n4596 , n2566 , n2971 );
    not g3109 ( n1385 , n2595 );
    or g3110 ( n5553 , n3210 , n5594 );
    or g3111 ( n5999 , n5747 , n1310 );
    or g3112 ( n3286 , n2908 , n552 );
    not g3113 ( n4770 , n4065 );
    or g3114 ( n3490 , n278 , n4798 );
    or g3115 ( n3961 , n3880 , n4438 );
    not g3116 ( n1738 , n5014 );
    not g3117 ( n4047 , n3394 );
    and g3118 ( n4408 , n4323 , n5702 );
    or g3119 ( n4036 , n1939 , n193 );
    and g3120 ( n2076 , n6218 , n593 );
    nor g3121 ( n1064 , n636 , n342 );
    and g3122 ( n4916 , n2139 , n3829 );
    nor g3123 ( n1031 , n3044 , n6125 );
    not g3124 ( n2089 , n4163 );
    not g3125 ( n3208 , n3131 );
    nor g3126 ( n2254 , n5685 , n2257 );
    or g3127 ( n3878 , n3619 , n1451 );
    and g3128 ( n6072 , n2968 , n5576 );
    or g3129 ( n2947 , n4760 , n4728 );
    or g3130 ( n1511 , n5493 , n3800 );
    not g3131 ( n5378 , n1915 );
    nor g3132 ( n3454 , n4108 , n47 );
    or g3133 ( n1502 , n2520 , n5453 );
    not g3134 ( n4832 , n5122 );
    and g3135 ( n5445 , n6250 , n1635 );
    or g3136 ( n3218 , n6093 , n5736 );
    or g3137 ( n1109 , n5362 , n5425 );
    or g3138 ( n5485 , n4756 , n5325 );
    nor g3139 ( n2568 , n3975 , n5338 );
    or g3140 ( n5686 , n1413 , n4456 );
    or g3141 ( n5855 , n1739 , n2822 );
    nor g3142 ( n4694 , n1123 , n4453 );
    nor g3143 ( n3794 , n4203 , n6247 );
    not g3144 ( n3912 , n3333 );
    not g3145 ( n5117 , n1594 );
    not g3146 ( n5768 , n3037 );
    or g3147 ( n3688 , n6184 , n272 );
    or g3148 ( n817 , n4563 , n3375 );
    or g3149 ( n1469 , n3752 , n4066 );
    and g3150 ( n411 , n2615 , n1413 );
    and g3151 ( n971 , n5209 , n2271 );
    or g3152 ( n3584 , n1023 , n3481 );
    not g3153 ( n821 , n5848 );
    or g3154 ( n2981 , n3451 , n4763 );
    not g3155 ( n4176 , n4570 );
    or g3156 ( n1302 , n6030 , n5397 );
    not g3157 ( n1503 , n1028 );
    not g3158 ( n1327 , n5490 );
    nor g3159 ( n6036 , n1905 , n2008 );
    not g3160 ( n2133 , n3963 );
    or g3161 ( n2243 , n3514 , n1675 );
    and g3162 ( n5791 , n4915 , n5150 );
    not g3163 ( n2455 , n985 );
    not g3164 ( n5887 , n918 );
    or g3165 ( n783 , n3580 , n953 );
    and g3166 ( n6067 , n3223 , n1954 );
    nor g3167 ( n5831 , n5602 , n4090 );
    nor g3168 ( n380 , n1000 , n1062 );
    nor g3169 ( n1088 , n505 , n4715 );
    not g3170 ( n98 , n1684 );
    not g3171 ( n5509 , n2970 );
    or g3172 ( n2463 , n1334 , n5092 );
    or g3173 ( n2354 , n1315 , n6098 );
    and g3174 ( n1584 , n1559 , n1582 );
    nor g3175 ( n5862 , n3140 , n895 );
    not g3176 ( n1066 , n2997 );
    nor g3177 ( n4226 , n1614 , n4846 );
    not g3178 ( n2689 , n2162 );
    or g3179 ( n3098 , n1326 , n368 );
    not g3180 ( n220 , n4332 );
    not g3181 ( n1821 , n2925 );
    not g3182 ( n1640 , n6 );
    or g3183 ( n5274 , n5328 , n408 );
    not g3184 ( n5115 , n2435 );
    and g3185 ( n3689 , n1482 , n3324 );
    or g3186 ( n2553 , n4348 , n2648 );
    or g3187 ( n1153 , n2 , n4485 );
    or g3188 ( n2936 , n1925 , n2870 );
    nor g3189 ( n1003 , n1935 , n6148 );
    not g3190 ( n6207 , n6053 );
    not g3191 ( n6176 , n2264 );
    nor g3192 ( n62 , n6012 , n3905 );
    or g3193 ( n507 , n3046 , n964 );
    not g3194 ( n5752 , n2930 );
    not g3195 ( n2724 , n4202 );
    or g3196 ( n5864 , n2316 , n294 );
    not g3197 ( n2656 , n1294 );
    not g3198 ( n4219 , n1122 );
    and g3199 ( n2094 , n3323 , n3289 );
    not g3200 ( n4148 , n541 );
    not g3201 ( n1361 , n5837 );
    not g3202 ( n3386 , n1378 );
    nor g3203 ( n6136 , n721 , n3288 );
    not g3204 ( n2176 , n1267 );
    not g3205 ( n546 , n2160 );
    and g3206 ( n1131 , n2343 , n2577 );
    or g3207 ( n1090 , n2583 , n6047 );
    nor g3208 ( n4785 , n4348 , n4600 );
    not g3209 ( n1475 , n914 );
    nor g3210 ( n3857 , n4242 , n5815 );
    and g3211 ( n3935 , n1564 , n4277 );
    nor g3212 ( n5265 , n3980 , n1995 );
    not g3213 ( n2090 , n410 );
    and g3214 ( n1876 , n3983 , n5237 );
    and g3215 ( n5244 , n5884 , n1008 );
    and g3216 ( n2811 , n6110 , n3849 );
    and g3217 ( n5163 , n5417 , n413 );
    nor g3218 ( n1747 , n6300 , n4053 );
    nor g3219 ( n4600 , n6208 , n5799 );
    nor g3220 ( n3469 , n1220 , n3577 );
    not g3221 ( n4479 , n3744 );
    not g3222 ( n87 , n4047 );
    and g3223 ( n732 , n559 , n3951 );
    not g3224 ( n158 , n5717 );
    nor g3225 ( n1611 , n6234 , n1071 );
    and g3226 ( n543 , n2005 , n2126 );
    and g3227 ( n2058 , n3125 , n6035 );
    nor g3228 ( n6065 , n2305 , n5875 );
    or g3229 ( n3900 , n25 , n645 );
    or g3230 ( n1695 , n762 , n3599 );
    or g3231 ( n5838 , n4243 , n3898 );
    not g3232 ( n834 , n5129 );
    not g3233 ( n2992 , n2770 );
    not g3234 ( n4889 , n2741 );
    or g3235 ( n1364 , n5892 , n2295 );
    or g3236 ( n2614 , n6002 , n4655 );
    not g3237 ( n887 , n5714 );
    or g3238 ( n3998 , n4499 , n5008 );
    not g3239 ( n5092 , n4620 );
    and g3240 ( n1739 , n1591 , n4873 );
    nor g3241 ( n4475 , n583 , n5687 );
    nor g3242 ( n1778 , n4353 , n4805 );
    nor g3243 ( n2609 , n552 , n5854 );
    or g3244 ( n3557 , n941 , n2148 );
    and g3245 ( n1624 , n3561 , n5634 );
    not g3246 ( n1894 , n796 );
    or g3247 ( n5547 , n259 , n2947 );
    nor g3248 ( n6254 , n4512 , n1896 );
    not g3249 ( n2199 , n3196 );
    not g3250 ( n4993 , n5699 );
    and g3251 ( n5623 , n288 , n986 );
    not g3252 ( n4650 , n3613 );
    nor g3253 ( n672 , n3972 , n964 );
    nor g3254 ( n575 , n437 , n3727 );
    nor g3255 ( n2371 , n792 , n5027 );
    not g3256 ( n281 , n1743 );
    or g3257 ( n4160 , n6075 , n3020 );
    nor g3258 ( n1365 , n1563 , n6170 );
    or g3259 ( n4792 , n2029 , n5915 );
    or g3260 ( n1119 , n5770 , n2092 );
    and g3261 ( n5151 , n3114 , n5627 );
    or g3262 ( n5216 , n2764 , n2654 );
    not g3263 ( n2144 , n4168 );
    or g3264 ( n5075 , n2910 , n3581 );
    not g3265 ( n2303 , n2231 );
    and g3266 ( n4155 , n3572 , n4248 );
    or g3267 ( n1095 , n5556 , n1059 );
    not g3268 ( n1767 , n4159 );
    or g3269 ( n1073 , n1817 , n2541 );
    nor g3270 ( n519 , n3492 , n5494 );
    nor g3271 ( n5660 , n6107 , n2168 );
    and g3272 ( n5700 , n3073 , n3209 );
    not g3273 ( n178 , n1092 );
    not g3274 ( n902 , n3019 );
    nor g3275 ( n4090 , n3911 , n3502 );
    nor g3276 ( n5762 , n2168 , n1718 );
    nor g3277 ( n4249 , n5205 , n1061 );
    or g3278 ( n4627 , n1893 , n3292 );
    nor g3279 ( n1911 , n5852 , n1999 );
    not g3280 ( n5671 , n4578 );
    nor g3281 ( n1452 , n2154 , n5843 );
    or g3282 ( n4871 , n4300 , n3112 );
    or g3283 ( n5863 , n4588 , n4374 );
    and g3284 ( n6002 , n1737 , n4674 );
    not g3285 ( n3015 , n2285 );
    nor g3286 ( n6101 , n1329 , n5227 );
    not g3287 ( n586 , n6069 );
    or g3288 ( n5594 , n2382 , n3925 );
    not g3289 ( n2478 , n3241 );
    not g3290 ( n2980 , n4039 );
    not g3291 ( n5861 , n3695 );
    nor g3292 ( n4261 , n4400 , n1027 );
    nor g3293 ( n5600 , n1171 , n541 );
    or g3294 ( n1038 , n5688 , n2872 );
    nor g3295 ( n5369 , n2496 , n3996 );
    or g3296 ( n2019 , n2604 , n1962 );
    not g3297 ( n4872 , n5418 );
    or g3298 ( n1190 , n4340 , n6083 );
    and g3299 ( n538 , n1491 , n3401 );
    and g3300 ( n1984 , n2167 , n4030 );
    not g3301 ( n3212 , n1025 );
    and g3302 ( n3891 , n2032 , n3225 );
    not g3303 ( n3934 , n562 );
    not g3304 ( n4191 , n4477 );
    not g3305 ( n1849 , n297 );
    and g3306 ( n4492 , n3303 , n1667 );
    or g3307 ( n5147 , n2409 , n2754 );
    or g3308 ( n4312 , n2152 , n1848 );
    not g3309 ( n1162 , n5663 );
    not g3310 ( n1963 , n5264 );
    nor g3311 ( n2516 , n5937 , n1753 );
    nor g3312 ( n1030 , n5061 , n2109 );
    nor g3313 ( n371 , n4987 , n4625 );
    nor g3314 ( n6151 , n484 , n1713 );
    nor g3315 ( n3397 , n106 , n2772 );
    or g3316 ( n4302 , n2127 , n2755 );
    and g3317 ( n3302 , n3433 , n4450 );
    and g3318 ( n3195 , n2667 , n2562 );
    or g3319 ( n5805 , n1432 , n1537 );
    or g3320 ( n2785 , n2444 , n3116 );
    nor g3321 ( n1510 , n777 , n3758 );
    not g3322 ( n3296 , n4550 );
    or g3323 ( n2023 , n5045 , n5722 );
    nor g3324 ( n5528 , n4618 , n697 );
    not g3325 ( n6173 , n2798 );
    and g3326 ( n1838 , n5947 , n5711 );
    and g3327 ( n3267 , n4003 , n5106 );
    or g3328 ( n4161 , n1695 , n3162 );
    nor g3329 ( n5009 , n5324 , n5905 );
    or g3330 ( n3137 , n1302 , n1232 );
    and g3331 ( n3604 , n2279 , n6070 );
    nor g3332 ( n5304 , n6158 , n4557 );
    nor g3333 ( n603 , n3822 , n3506 );
    or g3334 ( n4768 , n3030 , n2839 );
    or g3335 ( n4220 , n5367 , n6040 );
    and g3336 ( n6150 , n1698 , n5634 );
    or g3337 ( n4091 , n2269 , n2362 );
    nor g3338 ( n3134 , n4150 , n5619 );
    nor g3339 ( n6296 , n60 , n716 );
    nor g3340 ( n3252 , n2322 , n4531 );
    nor g3341 ( n926 , n2108 , n3178 );
    nor g3342 ( n2260 , n4773 , n477 );
    nor g3343 ( n448 , n2823 , n2831 );
    and g3344 ( n4510 , n1528 , n1515 );
    nor g3345 ( n4184 , n126 , n3538 );
    or g3346 ( n218 , n994 , n2769 );
    not g3347 ( n4361 , n5915 );
    nor g3348 ( n2898 , n5310 , n2830 );
    or g3349 ( n2169 , n5258 , n5190 );
    nor g3350 ( n102 , n5817 , n5760 );
    not g3351 ( n4708 , n1810 );
    nor g3352 ( n3148 , n5248 , n4590 );
    or g3353 ( n4206 , n2942 , n1288 );
    not g3354 ( n4083 , n3458 );
    or g3355 ( n5796 , n3402 , n1587 );
    not g3356 ( n4700 , n5437 );
    nor g3357 ( n3541 , n3660 , n1673 );
    not g3358 ( n6157 , n3841 );
    not g3359 ( n2565 , n6273 );
    or g3360 ( n302 , n3998 , n2537 );
    or g3361 ( n5010 , n3461 , n1050 );
    or g3362 ( n328 , n2448 , n2438 );
    and g3363 ( n1094 , n289 , n2841 );
    and g3364 ( n1287 , n4263 , n3893 );
    nor g3365 ( n3158 , n4119 , n3943 );
    not g3366 ( n917 , n483 );
    or g3367 ( n4289 , n2712 , n1885 );
    nor g3368 ( n2686 , n297 , n4683 );
    nor g3369 ( n1468 , n3229 , n4158 );
    and g3370 ( n2232 , n3813 , n5512 );
    or g3371 ( n5770 , n5966 , n2031 );
    or g3372 ( n1496 , n2799 , n783 );
    or g3373 ( n5701 , n499 , n5588 );
    not g3374 ( n4589 , n2860 );
    not g3375 ( n3065 , n4267 );
    not g3376 ( n1675 , n216 );
    not g3377 ( n1489 , n1679 );
    or g3378 ( n2373 , n417 , n5380 );
    or g3379 ( n4204 , n2875 , n4160 );
    or g3380 ( n3831 , n4743 , n656 );
    nor g3381 ( n669 , n2560 , n2909 );
    not g3382 ( n4606 , n2336 );
    nor g3383 ( n1353 , n1965 , n3557 );
    or g3384 ( n4349 , n5141 , n3947 );
    or g3385 ( n4356 , n232 , n2195 );
    or g3386 ( n2223 , n1811 , n720 );
    not g3387 ( n2202 , n2010 );
    nor g3388 ( n262 , n4774 , n655 );
    or g3389 ( n3712 , n4353 , n3520 );
    nor g3390 ( n2082 , n2406 , n5999 );
    not g3391 ( n4637 , n837 );
    or g3392 ( n4114 , n1705 , n173 );
    not g3393 ( n2771 , n1873 );
    not g3394 ( n1885 , n5948 );
    or g3395 ( n4537 , n4373 , n3393 );
    or g3396 ( n2011 , n2688 , n3537 );
    or g3397 ( n1674 , n1730 , n1793 );
    and g3398 ( n5703 , n5585 , n4447 );
    or g3399 ( n4223 , n3597 , n1455 );
    nor g3400 ( n3312 , n2268 , n3659 );
    not g3401 ( n2859 , n4156 );
    and g3402 ( n1019 , n5671 , n5492 );
    nor g3403 ( n632 , n4641 , n2141 );
    or g3404 ( n6270 , n1131 , n722 );
    or g3405 ( n5637 , n2119 , n1402 );
    not g3406 ( n3436 , n5986 );
    or g3407 ( n5313 , n3837 , n4530 );
    or g3408 ( n6278 , n1039 , n1083 );
    or g3409 ( n3814 , n612 , n4285 );
    nor g3410 ( n2275 , n1886 , n5217 );
    nor g3411 ( n449 , n305 , n2639 );
    not g3412 ( n174 , n3531 );
    or g3413 ( n4540 , n5821 , n3844 );
    not g3414 ( n3786 , n1287 );
    and g3415 ( n2174 , n3775 , n3672 );
    not g3416 ( n1878 , n536 );
    and g3417 ( n4974 , n5306 , n1478 );
    or g3418 ( n4123 , n1900 , n4447 );
    or g3419 ( n764 , n5416 , n2397 );
    nor g3420 ( n3498 , n1269 , n5109 );
    nor g3421 ( n704 , n1974 , n17 );
    or g3422 ( n2114 , n1306 , n1748 );
    not g3423 ( n4390 , n4120 );
    not g3424 ( n3382 , n6198 );
    or g3425 ( n5326 , n2673 , n1239 );
    not g3426 ( n3904 , n692 );
    and g3427 ( n5915 , n5116 , n4804 );
    not g3428 ( n2715 , n2003 );
    and g3429 ( n5884 , n3582 , n3809 );
    not g3430 ( n2211 , n2118 );
    or g3431 ( n54 , n2088 , n975 );
    and g3432 ( n6264 , n139 , n4561 );
    nor g3433 ( n1756 , n2474 , n179 );
    and g3434 ( n3809 , n915 , n4136 );
    or g3435 ( n3055 , n1588 , n4814 );
    not g3436 ( n610 , n3127 );
    nor g3437 ( n58 , n5195 , n1055 );
    and g3438 ( n5913 , n1242 , n2783 );
    not g3439 ( n5900 , n3817 );
    and g3440 ( n5827 , n2488 , n1996 );
    not g3441 ( n3187 , n2365 );
    nor g3442 ( n2062 , n3316 , n1366 );
    nor g3443 ( n1914 , n3155 , n7 );
    or g3444 ( n2451 , n3717 , n3911 );
    or g3445 ( n2507 , n3678 , n653 );
    nor g3446 ( n5820 , n103 , n3250 );
    not g3447 ( n5110 , n1104 );
    not g3448 ( n2908 , n1446 );
    nor g3449 ( n7 , n2545 , n286 );
    nor g3450 ( n117 , n670 , n4031 );
    or g3451 ( n1423 , n161 , n4968 );
    or g3452 ( n1261 , n2697 , n3637 );
    and g3453 ( n5048 , n399 , n2719 );
    not g3454 ( n2107 , n1422 );
    not g3455 ( n1547 , n5558 );
    or g3456 ( n2396 , n3673 , n4801 );
    or g3457 ( n4959 , n2493 , n3017 );
    nor g3458 ( n280 , n5901 , n628 );
    not g3459 ( n5920 , n5390 );
    or g3460 ( n2559 , n498 , n6028 );
    or g3461 ( n5741 , n4743 , n3061 );
    and g3462 ( n2403 , n6020 , n4094 );
    not g3463 ( n1565 , n4771 );
    or g3464 ( n1514 , n1999 , n1861 );
    or g3465 ( n3282 , n513 , n3713 );
    not g3466 ( n6141 , n2794 );
    and g3467 ( n3373 , n3390 , n2462 );
    and g3468 ( n78 , n1919 , n2217 );
    not g3469 ( n1264 , n577 );
    nor g3470 ( n4235 , n5182 , n3920 );
    nor g3471 ( n230 , n4167 , n6152 );
    not g3472 ( n5849 , n2557 );
    not g3473 ( n1051 , n5817 );
    not g3474 ( n3801 , n2611 );
    nor g3475 ( n804 , n1349 , n2783 );
    or g3476 ( n2179 , n3160 , n6029 );
    nor g3477 ( n3229 , n1371 , n3980 );
    or g3478 ( n885 , n2022 , n5545 );
    and g3479 ( n5150 , n1102 , n5058 );
    or g3480 ( n1587 , n3472 , n2769 );
    and g3481 ( n993 , n5044 , n5398 );
    nor g3482 ( n5908 , n3728 , n3515 );
    nor g3483 ( n3495 , n423 , n5595 );
    and g3484 ( n562 , n845 , n4772 );
    and g3485 ( n2074 , n2501 , n5000 );
    and g3486 ( n206 , n12 , n1656 );
    not g3487 ( n780 , n782 );
    nor g3488 ( n4095 , n1461 , n332 );
    or g3489 ( n453 , n5006 , n3944 );
    nor g3490 ( n841 , n4664 , n625 );
    not g3491 ( n3796 , n4746 );
    not g3492 ( n5261 , n4742 );
    nor g3493 ( n5271 , n1853 , n4059 );
    nor g3494 ( n1823 , n3360 , n1429 );
    or g3495 ( n5716 , n495 , n2247 );
    not g3496 ( n6050 , n190 );
    and g3497 ( n3439 , n1070 , n6035 );
    or g3498 ( n2225 , n723 , n154 );
    not g3499 ( n2147 , n4852 );
    or g3500 ( n5854 , n4484 , n5239 );
    and g3501 ( n1212 , n1759 , n1114 );
    and g3502 ( n1273 , n4572 , n2704 );
    nor g3503 ( n600 , n5059 , n5003 );
    or g3504 ( n3348 , n2949 , n4518 );
    or g3505 ( n1750 , n3194 , n5481 );
    nor g3506 ( n4942 , n4757 , n4556 );
    nor g3507 ( n6215 , n5374 , n222 );
    or g3508 ( n4493 , n800 , n4023 );
    not g3509 ( n307 , n1497 );
    or g3510 ( n1226 , n862 , n1725 );
    and g3511 ( n6220 , n355 , n1547 );
    not g3512 ( n3179 , n4493 );
    nor g3513 ( n1165 , n426 , n5141 );
    and g3514 ( n5910 , n5759 , n1668 );
    nor g3515 ( n1026 , n1861 , n5398 );
    not g3516 ( n4110 , n4705 );
    not g3517 ( n5423 , n2320 );
    and g3518 ( n235 , n2437 , n6022 );
    nor g3519 ( n6185 , n4507 , n5485 );
    and g3520 ( n5784 , n2888 , n1273 );
    or g3521 ( n3016 , n787 , n5308 );
    or g3522 ( n4515 , n1205 , n5201 );
    not g3523 ( n2625 , n2178 );
    or g3524 ( n4189 , n4330 , n2933 );
    nor g3525 ( n1539 , n3293 , n4241 );
    and g3526 ( n1980 , n3842 , n6127 );
    and g3527 ( n4409 , n4836 , n6138 );
    or g3528 ( n694 , n463 , n4166 );
    or g3529 ( n2926 , n4273 , n3280 );
    or g3530 ( n3328 , n1179 , n6227 );
    nor g3531 ( n1710 , n5378 , n2283 );
    not g3532 ( n2339 , n3100 );
    or g3533 ( n5785 , n4498 , n5734 );
    not g3534 ( n3524 , n2473 );
    or g3535 ( n66 , n3152 , n2797 );
    nor g3536 ( n4041 , n5166 , n3236 );
    or g3537 ( n6160 , n1859 , n4280 );
    not g3538 ( n786 , n184 );
    or g3539 ( n921 , n3728 , n1931 );
    and g3540 ( n3808 , n2927 , n2224 );
    or g3541 ( n5259 , n4289 , n6232 );
    or g3542 ( n4808 , n21 , n2359 );
    nor g3543 ( n1987 , n1576 , n4329 );
    nor g3544 ( n1352 , n3826 , n2602 );
    and g3545 ( n1360 , n3902 , n5366 );
    and g3546 ( n630 , n3539 , n3883 );
    or g3547 ( n5425 , n1217 , n1789 );
    nor g3548 ( n6202 , n3457 , n3168 );
    or g3549 ( n4237 , n3354 , n6024 );
    not g3550 ( n1465 , n880 );
    not g3551 ( n5465 , n4743 );
    or g3552 ( n723 , n237 , n866 );
    not g3553 ( n4145 , n3809 );
    nor g3554 ( n2398 , n5389 , n3864 );
    and g3555 ( n2460 , n4923 , n3894 );
    nor g3556 ( n498 , n1636 , n6278 );
    and g3557 ( n4801 , n2848 , n3742 );
    not g3558 ( n3966 , n1654 );
    or g3559 ( n460 , n4698 , n633 );
    or g3560 ( n1563 , n1946 , n2617 );
    or g3561 ( n5142 , n5368 , n5185 );
    not g3562 ( n1049 , n4408 );
    nor g3563 ( n1881 , n1023 , n1136 );
    and g3564 ( n2514 , n4975 , n1728 );
    not g3565 ( n2296 , n1761 );
    nor g3566 ( n2274 , n3484 , n1130 );
    not g3567 ( n2673 , n2804 );
    nor g3568 ( n2731 , n56 , n5586 );
    not g3569 ( n3742 , n3756 );
    or g3570 ( n3581 , n4515 , n5556 );
    or g3571 ( n2043 , n5225 , n2348 );
    or g3572 ( n5006 , n5360 , n5301 );
    and g3573 ( n1939 , n1337 , n1797 );
    not g3574 ( n5072 , n1240 );
    and g3575 ( n2016 , n5507 , n3255 );
    nor g3576 ( n2040 , n936 , n4035 );
    not g3577 ( n3446 , n3038 );
    nor g3578 ( n5278 , n4503 , n4717 );
    not g3579 ( n6303 , n1912 );
    and g3580 ( n2998 , n5529 , n216 );
    or g3581 ( n1086 , n2530 , n3183 );
    not g3582 ( n4733 , n5716 );
    not g3583 ( n140 , n2689 );
    nor g3584 ( n3506 , n3783 , n778 );
    or g3585 ( n4722 , n339 , n4542 );
    and g3586 ( n2035 , n1386 , n3965 );
    nor g3587 ( n3142 , n4248 , n1311 );
    not g3588 ( n5340 , n5202 );
    and g3589 ( n5332 , n671 , n513 );
    nor g3590 ( n4386 , n5925 , n2475 );
    not g3591 ( n1815 , n364 );
    or g3592 ( n1155 , n329 , n766 );
    or g3593 ( n4543 , n3066 , n709 );
    nor g3594 ( n5218 , n4897 , n6015 );
    not g3595 ( n4855 , n3745 );
    and g3596 ( n2364 , n970 , n5280 );
    or g3597 ( n3217 , n1097 , n2627 );
    and g3598 ( n1604 , n6137 , n6168 );
    nor g3599 ( n2629 , n2129 , n4471 );
    nor g3600 ( n5618 , n587 , n5223 );
    not g3601 ( n3005 , n2503 );
    not g3602 ( n4419 , n4894 );
    not g3603 ( n1787 , n6000 );
    or g3604 ( n3555 , n5532 , n5979 );
    and g3605 ( n436 , n5581 , n2546 );
    not g3606 ( n1816 , n2471 );
    and g3607 ( n2228 , n565 , n865 );
    or g3608 ( n5337 , n811 , n2739 );
    nor g3609 ( n4564 , n6085 , n5187 );
    not g3610 ( n84 , n4333 );
    or g3611 ( n293 , n3222 , n2246 );
    and g3612 ( n4572 , n3823 , n4207 );
    not g3613 ( n4809 , n4922 );
    and g3614 ( n831 , n2645 , n2060 );
    not g3615 ( n4545 , n906 );
    or g3616 ( n3576 , n4254 , n550 );
    or g3617 ( n5408 , n4092 , n376 );
    or g3618 ( n3628 , n2400 , n443 );
    nor g3619 ( n45 , n599 , n5473 );
    nor g3620 ( n3066 , n2027 , n3932 );
    nor g3621 ( n5069 , n2519 , n2477 );
    and g3622 ( n3617 , n2601 , n5807 );
    nor g3623 ( n3440 , n5506 , n5102 );
    nor g3624 ( n749 , n3452 , n2723 );
    not g3625 ( n1001 , n2189 );
    or g3626 ( n5782 , n4866 , n2233 );
    not g3627 ( n916 , n4541 );
    nor g3628 ( n4581 , n594 , n1651 );
    nor g3629 ( n5306 , n3700 , n2540 );
    not g3630 ( n179 , n998 );
    or g3631 ( n332 , n5303 , n2921 );
    and g3632 ( n3745 , n1304 , n1151 );
    or g3633 ( n5051 , n1723 , n1466 );
    nor g3634 ( n5380 , n5238 , n712 );
    not g3635 ( n5580 , n506 );
    nor g3636 ( n5189 , n4663 , n3674 );
    not g3637 ( n3207 , n5864 );
    or g3638 ( n4162 , n3577 , n4319 );
    and g3639 ( n3049 , n885 , n4970 );
    nor g3640 ( n82 , n5967 , n2398 );
    or g3641 ( n5858 , n785 , n5708 );
    or g3642 ( n5621 , n254 , n2325 );
    nor g3643 ( n1101 , n5645 , n4423 );
    or g3644 ( n6188 , n4957 , n2358 );
    not g3645 ( n5673 , n1704 );
    and g3646 ( n4698 , n2063 , n3809 );
    not g3647 ( n2196 , n913 );
    and g3648 ( n6030 , n3431 , n4816 );
    nor g3649 ( n5682 , n5524 , n2342 );
    or g3650 ( n614 , n2819 , n5319 );
    not g3651 ( n5990 , n2905 );
    or g3652 ( n6000 , n2551 , n3084 );
    not g3653 ( n3044 , n2228 );
    nor g3654 ( n1448 , n5575 , n4900 );
    not g3655 ( n6096 , n4848 );
    or g3656 ( n2297 , n5780 , n4298 );
    not g3657 ( n3400 , n177 );
    and g3658 ( n5539 , n4316 , n121 );
    not g3659 ( n35 , n4781 );
    or g3660 ( n3155 , n6129 , n1665 );
    or g3661 ( n1825 , n4599 , n4224 );
    nor g3662 ( n3336 , n2478 , n1934 );
    not g3663 ( n2456 , n610 );
    nor g3664 ( n4350 , n2791 , n4532 );
    not g3665 ( n681 , n1505 );
    not g3666 ( n1504 , n842 );
    nor g3667 ( n330 , n4142 , n1044 );
    and g3668 ( n526 , n3858 , n4751 );
    nor g3669 ( n406 , n1019 , n5126 );
    and g3670 ( n2421 , n1119 , n31 );
    and g3671 ( n2962 , n5890 , n357 );
    or g3672 ( n5039 , n4569 , n4138 );
    nor g3673 ( n3758 , n18 , n2705 );
    or g3674 ( n3658 , n6103 , n3201 );
    nor g3675 ( n4282 , n5277 , n81 );
    or g3676 ( n2630 , n1413 , n4376 );
    or g3677 ( n3241 , n3061 , n1952 );
    nor g3678 ( n3828 , n4804 , n421 );
    nor g3679 ( n4692 , n3486 , n6212 );
    not g3680 ( n5148 , n126 );
    not g3681 ( n232 , n3660 );
    and g3682 ( n1180 , n4397 , n4918 );
    not g3683 ( n1946 , n6050 );
    and g3684 ( n1817 , n5170 , n5772 );
    nor g3685 ( n258 , n461 , n412 );
    nor g3686 ( n752 , n5298 , n487 );
    nor g3687 ( n1429 , n1958 , n1522 );
    or g3688 ( n4504 , n4291 , n2818 );
    not g3689 ( n4988 , n316 );
    not g3690 ( n4755 , n4940 );
    nor g3691 ( n5497 , n2757 , n2903 );
    and g3692 ( n5946 , n395 , n4194 );
    or g3693 ( n3947 , n4082 , n3039 );
    not g3694 ( n5903 , n5357 );
    not g3695 ( n6012 , n1516 );
    nor g3696 ( n823 , n5551 , n3624 );
    and g3697 ( n476 , n1989 , n5353 );
    and g3698 ( n1762 , n5129 , n662 );
    or g3699 ( n872 , n1450 , n3899 );
    nor g3700 ( n4920 , n4553 , n5731 );
    nor g3701 ( n238 , n5091 , n2147 );
    not g3702 ( n1575 , n3651 );
    and g3703 ( n1225 , n1379 , n2192 );
    or g3704 ( n2497 , n5488 , n2035 );
    or g3705 ( n492 , n5389 , n3877 );
    and g3706 ( n4397 , n1139 , n2830 );
    not g3707 ( n4921 , n5627 );
    and g3708 ( n1712 , n2662 , n1635 );
    not g3709 ( n938 , n3679 );
    or g3710 ( n1250 , n1706 , n3263 );
    nor g3711 ( n3384 , n1949 , n4529 );
    nor g3712 ( n5371 , n1340 , n6006 );
    nor g3713 ( n1744 , n4676 , n5043 );
    or g3714 ( n2096 , n1124 , n1310 );
    nor g3715 ( n162 , n5990 , n5130 );
    or g3716 ( n5317 , n5173 , n4475 );
    or g3717 ( n4971 , n6197 , n3860 );
    nor g3718 ( n3108 , n2378 , n2889 );
    nor g3719 ( n5053 , n30 , n4789 );
    and g3720 ( n1262 , n5213 , n5096 );
    not g3721 ( n3987 , n4965 );
    not g3722 ( n6109 , n3606 );
    and g3723 ( n3260 , n3379 , n5990 );
    nor g3724 ( n4542 , n1002 , n2467 );
    not g3725 ( n2593 , n5436 );
    or g3726 ( n2742 , n5238 , n5001 );
    or g3727 ( n213 , n5812 , n1913 );
    or g3728 ( n4187 , n2647 , n4484 );
    or g3729 ( n4446 , n5849 , n4393 );
    or g3730 ( n4948 , n1461 , n5833 );
    nor g3731 ( n595 , n4010 , n5528 );
    nor g3732 ( n4769 , n6079 , n4669 );
    or g3733 ( n4010 , n5081 , n3642 );
    nor g3734 ( n4750 , n2826 , n5865 );
    or g3735 ( n3149 , n1083 , n1204 );
    not g3736 ( n2234 , n2503 );
    not g3737 ( n2281 , n638 );
    nor g3738 ( n2165 , n1413 , n3717 );
    nor g3739 ( n3637 , n461 , n1253 );
    or g3740 ( n1305 , n2883 , n1230 );
    or g3741 ( n2709 , n2117 , n718 );
    not g3742 ( n4989 , n4767 );
    or g3743 ( n2495 , n3320 , n2106 );
    nor g3744 ( n2531 , n2771 , n3439 );
    or g3745 ( n5537 , n2287 , n724 );
    and g3746 ( n980 , n72 , n4720 );
    nor g3747 ( n198 , n459 , n1537 );
    not g3748 ( n3107 , n5961 );
    not g3749 ( n421 , n5973 );
    and g3750 ( n4382 , n315 , n5970 );
    and g3751 ( n1615 , n3443 , n3980 );
    not g3752 ( n3031 , n4668 );
    or g3753 ( n927 , n2360 , n5631 );
    and g3754 ( n38 , n1992 , n5387 );
    not g3755 ( n2148 , n4047 );
    not g3756 ( n6008 , n5111 );
    nor g3757 ( n2982 , n176 , n4660 );
    nor g3758 ( n4395 , n3407 , n1806 );
    and g3759 ( n3000 , n3379 , n1675 );
    or g3760 ( n440 , n3419 , n6209 );
    nor g3761 ( n5220 , n4335 , n5331 );
    and g3762 ( n3716 , n4928 , n4534 );
    or g3763 ( n3486 , n4771 , n4231 );
    and g3764 ( n1920 , n2825 , n4092 );
    or g3765 ( n5764 , n2523 , n5171 );
    not g3766 ( n6227 , n4555 );
    not g3767 ( n3270 , n4306 );
    not g3768 ( n1120 , n4810 );
    nor g3769 ( n4802 , n2634 , n2459 );
    or g3770 ( n5441 , n616 , n476 );
    or g3771 ( n4124 , n1634 , n5944 );
    and g3772 ( n1910 , n5618 , n3079 );
    nor g3773 ( n2304 , n4974 , n5874 );
    buf g3774 ( n4800 , n1857 );
    nor g3775 ( n968 , n2919 , n595 );
    not g3776 ( n335 , n2574 );
    not g3777 ( n4236 , n3796 );
    and g3778 ( n955 , n3207 , n1722 );
    and g3779 ( n2112 , n5591 , n2081 );
    nor g3780 ( n1284 , n2691 , n1752 );
    or g3781 ( n2010 , n1972 , n823 );
    nor g3782 ( n6172 , n5662 , n259 );
    not g3783 ( n338 , n6277 );
    or g3784 ( n1480 , n189 , n5388 );
    or g3785 ( n5567 , n4445 , n5255 );
    or g3786 ( n3698 , n2449 , n5500 );
    not g3787 ( n5479 , n4533 );
    or g3788 ( n5587 , n4180 , n2098 );
    not g3789 ( n135 , n5581 );
    not g3790 ( n5543 , n2993 );
    or g3791 ( n4065 , n1562 , n925 );
    and g3792 ( n1497 , n5431 , n4809 );
    or g3793 ( n1182 , n3985 , n4934 );
    not g3794 ( n5807 , n5534 );
    or g3795 ( n5303 , n1076 , n5126 );
    nor g3796 ( n3522 , n5166 , n641 );
    nor g3797 ( n4684 , n749 , n1358 );
    not g3798 ( n2583 , n3480 );
    and g3799 ( n5868 , n1268 , n2196 );
    nor g3800 ( n3707 , n1750 , n2181 );
    or g3801 ( n1037 , n4364 , n5927 );
    not g3802 ( n2462 , n4608 );
    nor g3803 ( n4126 , n4569 , n3603 );
    or g3804 ( n1974 , n5106 , n6034 );
    nor g3805 ( n5951 , n843 , n3040 );
    not g3806 ( n3024 , n99 );
    and g3807 ( n3739 , n2011 , n6046 );
    and g3808 ( n930 , n2014 , n1045 );
    and g3809 ( n5576 , n5311 , n4378 );
    not g3810 ( n4678 , n2967 );
    and g3811 ( n1679 , n4943 , n3512 );
    not g3812 ( n4406 , n2045 );
    or g3813 ( n2312 , n71 , n4722 );
    and g3814 ( n5170 , n5683 , n6195 );
    not g3815 ( n1463 , n2724 );
    and g3816 ( n2857 , n3823 , n1044 );
    or g3817 ( n6281 , n1841 , n4042 );
    not g3818 ( n2794 , n2097 );
    and g3819 ( n1899 , n3862 , n4067 );
    not g3820 ( n1976 , n4524 );
    nor g3821 ( n2240 , n899 , n5777 );
    or g3822 ( n896 , n3270 , n3616 );
    or g3823 ( n4991 , n6207 , n2738 );
    or g3824 ( n53 , n1969 , n4382 );
    not g3825 ( n381 , n1755 );
    nor g3826 ( n5361 , n1616 , n5658 );
    nor g3827 ( n537 , n3127 , n2445 );
    not g3828 ( n2071 , n4916 );
    not g3829 ( n3815 , n3524 );
    not g3830 ( n5952 , n4380 );
    nor g3831 ( n2345 , n5122 , n5695 );
    nor g3832 ( n143 , n5235 , n2665 );
    and g3833 ( n1256 , n2133 , n5288 );
    or g3834 ( n1240 , n917 , n3002 );
    not g3835 ( n5715 , n5789 );
    and g3836 ( n42 , n6298 , n3325 );
    nor g3837 ( n1233 , n3429 , n608 );
    nor g3838 ( n1775 , n609 , n4381 );
    or g3839 ( n621 , n2931 , n891 );
    and g3840 ( n1157 , n4215 , n3364 );
    not g3841 ( n4367 , n5377 );
    not g3842 ( n2543 , n717 );
    not g3843 ( n5965 , n2045 );
    or g3844 ( n6206 , n1200 , n6204 );
    and g3845 ( n484 , n4842 , n2922 );
    and g3846 ( n4297 , n1177 , n5928 );
    or g3847 ( n4068 , n3472 , n2394 );
    or g3848 ( n5609 , n4843 , n4169 );
    nor g3849 ( n2788 , n3829 , n1154 );
    not g3850 ( n1494 , n3716 );
    nor g3851 ( n2971 , n107 , n2379 );
    or g3852 ( n3013 , n590 , n1553 );
    or g3853 ( n3949 , n3818 , n1377 );
    or g3854 ( n3249 , n3890 , n4405 );
    and g3855 ( n637 , n285 , n1090 );
    not g3856 ( n301 , n196 );
    nor g3857 ( n309 , n1381 , n444 );
    not g3858 ( n3618 , n3891 );
    nor g3859 ( n5047 , n3929 , n6266 );
    not g3860 ( n6189 , n148 );
    and g3861 ( n5655 , n5381 , n4104 );
    nor g3862 ( n389 , n4561 , n3774 );
    or g3863 ( n4496 , n5796 , n3979 );
    and g3864 ( n4512 , n2432 , n4106 );
    not g3865 ( n531 , n1413 );
    nor g3866 ( n4559 , n2243 , n2330 );
    and g3867 ( n4529 , n4896 , n366 );
    or g3868 ( n3337 , n3536 , n323 );
    and g3869 ( n1140 , n742 , n4032 );
    nor g3870 ( n2167 , n5632 , n2896 );
    not g3871 ( n2506 , n6210 );
    not g3872 ( n912 , n2614 );
    not g3873 ( n577 , n5269 );
    not g3874 ( n1108 , n5333 );
    nor g3875 ( n2581 , n95 , n4051 );
    nor g3876 ( n1852 , n5995 , n491 );
    and g3877 ( n1737 , n4511 , n556 );
    nor g3878 ( n5815 , n5173 , n2479 );
    not g3879 ( n6217 , n1598 );
    nor g3880 ( n4939 , n1106 , n723 );
    or g3881 ( n4060 , n4613 , n273 );
    nor g3882 ( n5754 , n2850 , n5895 );
    nor g3883 ( n4262 , n2289 , n6037 );
    not g3884 ( n138 , n2621 );
    nor g3885 ( n4371 , n4477 , n5159 );
    nor g3886 ( n2424 , n3345 , n3468 );
    not g3887 ( n5750 , n3926 );
    not g3888 ( n4283 , n350 );
    and g3889 ( n154 , n2708 , n4516 );
    or g3890 ( n5633 , n150 , n5724 );
    or g3891 ( n5582 , n4742 , n5004 );
    or g3892 ( n654 , n5152 , n4568 );
    not g3893 ( n3975 , n5746 );
    or g3894 ( n170 , n5888 , n1814 );
    nor g3895 ( n1254 , n2349 , n2576 );
    nor g3896 ( n4020 , n4399 , n1093 );
    nor g3897 ( n2920 , n3007 , n3095 );
    nor g3898 ( n2464 , n2149 , n2989 );
    not g3899 ( n1824 , n5521 );
    or g3900 ( n6286 , n118 , n2636 );
    and g3901 ( n5570 , n4879 , n4962 );
    or g3902 ( n3994 , n129 , n2984 );
    or g3903 ( n923 , n5874 , n3026 );
    or g3904 ( n4147 , n3568 , n4143 );
    not g3905 ( n5105 , n1568 );
    or g3906 ( n4972 , n1515 , n4741 );
    not g3907 ( n744 , n1360 );
    and g3908 ( n2806 , n2455 , n1409 );
    nor g3909 ( n5876 , n5177 , n6199 );
    or g3910 ( n4530 , n1068 , n1684 );
    and g3911 ( n4602 , n1385 , n2256 );
    not g3912 ( n3784 , n1094 );
    or g3913 ( n5740 , n3221 , n728 );
    and g3914 ( n5264 , n92 , n689 );
    or g3915 ( n3944 , n2335 , n4815 );
    and g3916 ( n3466 , n5744 , n4419 );
    and g3917 ( n6016 , n256 , n660 );
    or g3918 ( n4643 , n2456 , n3072 );
    and g3919 ( n2070 , n2145 , n5624 );
    nor g3920 ( n3184 , n3343 , n87 );
    not g3921 ( n3482 , n4339 );
    not g3922 ( n579 , n6226 );
    not g3923 ( n5489 , n2848 );
    not g3924 ( n395 , n5128 );
    not g3925 ( n4314 , n3199 );
    and g3926 ( n4267 , n3110 , n2419 );
    nor g3927 ( n838 , n4112 , n3285 );
    not g3928 ( n3242 , n792 );
    not g3929 ( n987 , n310 );
    nor g3930 ( n3561 , n2644 , n201 );
    or g3931 ( n31 , n5365 , n4222 );
    not g3932 ( n2175 , n3792 );
    not g3933 ( n1959 , n1605 );
    or g3934 ( n5289 , n3676 , n3014 );
    or g3935 ( n2623 , n3741 , n1476 );
    not g3936 ( n4239 , n2117 );
    nor g3937 ( n5608 , n4639 , n4173 );
    not g3938 ( n1389 , n337 );
    nor g3939 ( n5382 , n76 , n2623 );
    nor g3940 ( n5446 , n4718 , n2613 );
    not g3941 ( n2245 , n1576 );
    not g3942 ( n1689 , n2200 );
    not g3943 ( n236 , n5090 );
    nor g3944 ( n79 , n4700 , n4500 );
    nor g3945 ( n3138 , n1202 , n2414 );
    or g3946 ( n4480 , n6168 , n427 );
    and g3947 ( n1844 , n4755 , n3164 );
    or g3948 ( n415 , n3267 , n1127 );
    or g3949 ( n3052 , n5106 , n6249 );
    and g3950 ( n2914 , n711 , n490 );
    not g3951 ( n5886 , n758 );
    not g3952 ( n3304 , n4291 );
    nor g3953 ( n1950 , n2473 , n2792 );
    not g3954 ( n2624 , n5538 );
    and g3955 ( n4633 , n2962 , n5411 );
    or g3956 ( n393 , n2549 , n2253 );
    not g3957 ( n2805 , n5048 );
    or g3958 ( n5482 , n5901 , n2676 );
    and g3959 ( n5825 , n5336 , n2734 );
    and g3960 ( n4790 , n2124 , n5857 );
    not g3961 ( n5534 , n1951 );
    not g3962 ( n2973 , n2243 );
    or g3963 ( n1334 , n239 , n3987 );
    and g3964 ( n813 , n956 , n1052 );
    nor g3965 ( n6104 , n927 , n5149 );
    or g3966 ( n2752 , n5135 , n1116 );
    not g3967 ( n895 , n3421 );
    or g3968 ( n803 , n1318 , n3936 );
    and g3969 ( n3287 , n4849 , n1586 );
    and g3970 ( n1998 , n5788 , n4002 );
    or g3971 ( n5630 , n5399 , n2928 );
    or g3972 ( n1374 , n3887 , n3098 );
    not g3973 ( n4514 , n1370 );
    or g3974 ( n1481 , n159 , n1632 );
    or g3975 ( n3221 , n2589 , n202 );
    not g3976 ( n305 , n5773 );
    not g3977 ( n5328 , n3560 );
    or g3978 ( n3223 , n5305 , n5263 );
    not g3979 ( n4548 , n452 );
    or g3980 ( n2967 , n5882 , n84 );
    or g3981 ( n4304 , n4790 , n1681 );
    and g3982 ( n2929 , n3170 , n5365 );
    not g3983 ( n1945 , n5285 );
    not g3984 ( n981 , n2604 );
    nor g3985 ( n5451 , n1108 , n5178 );
    not g3986 ( n5797 , n2281 );
    and g3987 ( n4853 , n2190 , n2803 );
    and g3988 ( n2077 , n2125 , n2202 );
    or g3989 ( n1803 , n1599 , n4924 );
    or g3990 ( n2143 , n4675 , n576 );
    and g3991 ( n6013 , n6192 , n1664 );
    not g3992 ( n3233 , n521 );
    or g3993 ( n5452 , n3259 , n3601 );
    not g3994 ( n4749 , n523 );
    not g3995 ( n1060 , n1774 );
    or g3996 ( n5687 , n122 , n4271 );
    and g3997 ( n2907 , n2233 , n1181 );
    not g3998 ( n3303 , n1727 );
    not g3999 ( n3021 , n2425 );
    and g4000 ( n5575 , n464 , n1930 );
    not g4001 ( n1270 , n2584 );
    or g4002 ( n4775 , n5881 , n2509 );
    or g4003 ( n2720 , n2884 , n29 );
    not g4004 ( n2880 , n4656 );
    not g4005 ( n4271 , n5707 );
    not g4006 ( n4039 , n3366 );
    not g4007 ( n708 , n1566 );
    nor g4008 ( n5632 , n1262 , n5042 );
    and g4009 ( n1191 , n2418 , n2032 );
    or g4010 ( n1466 , n2210 , n3463 );
    or g4011 ( n3856 , n2453 , n1795 );
    not g4012 ( n3078 , n4447 );
    nor g4013 ( n482 , n5858 , n4086 );
    not g4014 ( n5533 , n196 );
    and g4015 ( n1114 , n3434 , n1849 );
    or g4016 ( n3045 , n2282 , n5030 );
    or g4017 ( n1583 , n3952 , n580 );
    not g4018 ( n2607 , n3374 );
    or g4019 ( n1358 , n5206 , n2659 );
    or g4020 ( n1602 , n5176 , n5755 );
    not g4021 ( n41 , n439 );
    or g4022 ( n2400 , n4562 , n2262 );
    nor g4023 ( n3569 , n5276 , n4982 );
    not g4024 ( n148 , n4194 );
    or g4025 ( n2528 , n2884 , n2804 );
    and g4026 ( n1786 , n3182 , n1438 );
    nor g4027 ( n5149 , n4 , n3910 );
    not g4028 ( n1007 , n3780 );
    or g4029 ( n6247 , n3191 , n2394 );
    and g4030 ( n3458 , n4437 , n2327 );
    nor g4031 ( n1112 , n2781 , n1763 );
    nor g4032 ( n2461 , n4098 , n1981 );
    and g4033 ( n1770 , n2223 , n2882 );
    not g4034 ( n5350 , n1906 );
    or g4035 ( n210 , n1942 , n2940 );
    nor g4036 ( n5403 , n3507 , n2650 );
    not g4037 ( n6181 , n4422 );
    not g4038 ( n4552 , n4023 );
    or g4039 ( n4814 , n3585 , n5241 );
    not g4040 ( n5930 , n3588 );
    or g4041 ( n5540 , n5023 , n6238 );
    and g4042 ( n1393 , n2543 , n4117 );
    or g4043 ( n4402 , n2410 , n870 );
    or g4044 ( n1833 , n5286 , n5609 );
    or g4045 ( n2620 , n3246 , n4831 );
    or g4046 ( n4611 , n946 , n1715 );
    nor g4047 ( n1938 , n189 , n5198 );
    not g4048 ( n4021 , n2232 );
    not g4049 ( n288 , n49 );
    nor g4050 ( n5988 , n2313 , n1490 );
    and g4051 ( n4026 , n3204 , n1836 );
    not g4052 ( n3492 , n6165 );
    and g4053 ( n4342 , n4277 , n3560 );
    or g4054 ( n2875 , n4737 , n2001 );
    not g4055 ( n3511 , n1324 );
    and g4056 ( n3453 , n2232 , n1342 );
    and g4057 ( n1836 , n538 , n5842 );
    nor g4058 ( n3825 , n1048 , n5543 );
    nor g4059 ( n1129 , n4470 , n5590 );
    and g4060 ( n3356 , n5893 , n5701 );
    not g4061 ( n2649 , n5850 );
    nor g4062 ( n1558 , n2711 , n5279 );
    not g4063 ( n6301 , n4954 );
    or g4064 ( n4396 , n2236 , n1801 );
    or g4065 ( n5448 , n1749 , n112 );
    nor g4066 ( n3727 , n3031 , n3185 );
    or g4067 ( n3409 , n5541 , n5637 );
    or g4068 ( n1295 , n1402 , n5060 );
    not g4069 ( n2802 , n2831 );
    and g4070 ( n5161 , n4430 , n3300 );
    not g4071 ( n3755 , n3290 );
    or g4072 ( n5850 , n228 , n3439 );
    and g4073 ( n331 , n2796 , n4979 );
    not g4074 ( n2428 , n500 );
    or g4075 ( n3145 , n5199 , n699 );
    or g4076 ( n4591 , n1724 , n4171 );
    or g4077 ( n5751 , n4033 , n4185 );
    and g4078 ( n2053 , n3658 , n3323 );
    not g4079 ( n259 , n1813 );
    or g4080 ( n5067 , n1025 , n3814 );
    not g4081 ( n5610 , n5150 );
    or g4082 ( n6098 , n1726 , n5006 );
    and g4083 ( n1178 , n2248 , n5014 );
    not g4084 ( n5008 , n140 );
    not g4085 ( n1436 , n3567 );
    nor g4086 ( n1585 , n466 , n3792 );
    and g4087 ( n5242 , n3159 , n3100 );
    not g4088 ( n2640 , n2213 );
    and g4089 ( n3038 , n1157 , n5215 );
    not g4090 ( n1046 , n824 );
    or g4091 ( n4982 , n5157 , n1596 );
    and g4092 ( n1907 , n4890 , n452 );
    not g4093 ( n3244 , n1564 );
    not g4094 ( n2846 , n1898 );
    not g4095 ( n4128 , n3260 );
    or g4096 ( n5084 , n5925 , n768 );
    not g4097 ( n5696 , n2340 );
    not g4098 ( n6121 , n3921 );
    not g4099 ( n5892 , n4214 );
    or g4100 ( n1377 , n5021 , n2974 );
    not g4101 ( n1652 , n2758 );
    not g4102 ( n224 , n4804 );
    and g4103 ( n1464 , n131 , n384 );
    not g4104 ( n4248 , n6118 );
    and g4105 ( n312 , n5928 , n782 );
    not g4106 ( n4869 , n1273 );
    nor g4107 ( n733 , n4699 , n4689 );
    and g4108 ( n1268 , n3893 , n3861 );
    and g4109 ( n1396 , n4493 , n2873 );
    and g4110 ( n5668 , n835 , n356 );
    nor g4111 ( n1107 , n4721 , n5486 );
    not g4112 ( n2454 , n1211 );
    and g4113 ( n3374 , n2778 , n200 );
    or g4114 ( n3194 , n4128 , n4488 );
    or g4115 ( n2713 , n201 , n2370 );
    or g4116 ( n193 , n489 , n719 );
    not g4117 ( n499 , n5873 );
    nor g4118 ( n5835 , n5516 , n66 );
    or g4119 ( n5657 , n1149 , n2831 );
    not g4120 ( n2617 , n1871 );
    and g4121 ( n253 , n3052 , n4003 );
    or g4122 ( n6061 , n73 , n5329 );
    not g4123 ( n4858 , n6003 );
    or g4124 ( n1028 , n1347 , n3794 );
    and g4125 ( n1622 , n4848 , n1461 );
    not g4126 ( n735 , n648 );
    or g4127 ( n120 , n4735 , n3784 );
    nor g4128 ( n3456 , n4305 , n2308 );
    nor g4129 ( n2183 , n3860 , n4428 );
    not g4130 ( n5698 , n882 );
    or g4131 ( n1197 , n3787 , n3770 );
    or g4132 ( n1782 , n234 , n4920 );
    and g4133 ( n2383 , n3732 , n4144 );
    or g4134 ( n3310 , n157 , n4990 );
    not g4135 ( n1244 , n4568 );
    not g4136 ( n4962 , n6200 );
    or g4137 ( n3254 , n4069 , n3781 );
    or g4138 ( n2018 , n1978 , n3042 );
    not g4139 ( n826 , n488 );
    and g4140 ( n5228 , n6288 , n4866 );
    or g4141 ( n458 , n4011 , n1182 );
    and g4142 ( n1495 , n2115 , n5623 );
    not g4143 ( n3540 , n172 );
    not g4144 ( n52 , n2093 );
    and g4145 ( n2088 , n1308 , n1737 );
    or g4146 ( n3923 , n4327 , n2173 );
    or g4147 ( n4873 , n5324 , n5853 );
    not g4148 ( n1515 , n4050 );
    or g4149 ( n903 , n5076 , n431 );
    or g4150 ( n4544 , n1327 , n923 );
    or g4151 ( n3936 , n3083 , n5224 );
    and g4152 ( n736 , n5969 , n1978 );
    not g4153 ( n2560 , n2075 );
    nor g4154 ( n2536 , n6119 , n1184 );
    and g4155 ( n4428 , n1904 , n3633 );
    nor g4156 ( n136 , n4370 , n3963 );
    not g4157 ( n4850 , n3458 );
    or g4158 ( n6261 , n3490 , n6191 );
    not g4159 ( n5167 , n6002 );
    and g4160 ( n1444 , n1183 , n5512 );
    or g4161 ( n3012 , n4286 , n5707 );
    and g4162 ( n6 , n2344 , n5466 );
    and g4163 ( n2878 , n668 , n1164 );
    not g4164 ( n6273 , n305 );
    not g4165 ( n3939 , n3084 );
    nor g4166 ( n4243 , n5638 , n2530 );
    or g4167 ( n4863 , n5079 , n2812 );
    and g4168 ( n2941 , n2050 , n2720 );
    nor g4169 ( n1596 , n6142 , n3120 );
    or g4170 ( n3334 , n5769 , n4182 );
    and g4171 ( n2135 , n2107 , n4445 );
    or g4172 ( n2645 , n2247 , n751 );
    or g4173 ( n828 , n1091 , n2500 );
    nor g4174 ( n1508 , n2278 , n6085 );
    not g4175 ( n3651 , n3929 );
    nor g4176 ( n4404 , n4429 , n934 );
    not g4177 ( n1400 , n3429 );
    and g4178 ( n2441 , n2693 , n1906 );
    not g4179 ( n3410 , n4087 );
    not g4180 ( n2052 , n2355 );
    or g4181 ( n4192 , n1186 , n5725 );
    nor g4182 ( n3211 , n2543 , n2982 );
    and g4183 ( n4847 , n1509 , n5851 );
    not g4184 ( n2124 , n5190 );
    nor g4185 ( n1403 , n3095 , n1908 );
    or g4186 ( n5629 , n266 , n2293 );
    and g4187 ( n4728 , n5483 , n5096 );
    nor g4188 ( n5727 , n3847 , n4946 );
    or g4189 ( n5790 , n4894 , n6279 );
    or g4190 ( n4667 , n5488 , n5019 );
    not g4191 ( n2605 , n2276 );
    or g4192 ( n5348 , n4220 , n1437 );
    nor g4193 ( n4025 , n1820 , n1844 );
    nor g4194 ( n5944 , n6072 , n2033 );
    not g4195 ( n4501 , n2963 );
    nor g4196 ( n2186 , n3033 , n5219 );
    not g4197 ( n3715 , n2691 );
    and g4198 ( n4323 , n4797 , n480 );
    not g4199 ( n4089 , n2332 );
    not g4200 ( n2207 , n1678 );
    not g4201 ( n3661 , n5037 );
    or g4202 ( n175 , n5852 , n6183 );
    not g4203 ( n1701 , n2048 );
    or g4204 ( n612 , n240 , n3644 );
    or g4205 ( n6095 , n2600 , n1199 );
    not g4206 ( n3122 , n4134 );
    not g4207 ( n4450 , n1690 );
    nor g4208 ( n1523 , n4319 , n2081 );
    or g4209 ( n385 , n5637 , n2484 );
    not g4210 ( n4469 , n3885 );
    and g4211 ( n4953 , n4341 , n5907 );
    and g4212 ( n5011 , n1751 , n5540 );
    nor g4213 ( n1137 , n5602 , n4981 );
    not g4214 ( n2061 , n2506 );
    nor g4215 ( n1925 , n2563 , n2428 );
    and g4216 ( n1122 , n998 , n4276 );
    and g4217 ( n2017 , n2990 , n4727 );
    nor g4218 ( n5612 , n5049 , n4269 );
    and g4219 ( n1863 , n1574 , n5375 );
    and g4220 ( n4117 , n989 , n967 );
    or g4221 ( n4258 , n430 , n2346 );
    and g4222 ( n601 , n6251 , n526 );
    or g4223 ( n2628 , n1052 , n3381 );
    not g4224 ( n6274 , n3778 );
    or g4225 ( n675 , n4994 , n1916 );
    not g4226 ( n3928 , n1175 );
    nor g4227 ( n1395 , n400 , n1278 );
    or g4228 ( n3554 , n4935 , n916 );
    not g4229 ( n5885 , n815 );
    or g4230 ( n5470 , n1699 , n389 );
    not g4231 ( n5996 , n1459 );
    or g4232 ( n2481 , n4598 , n2612 );
    not g4233 ( n185 , n2282 );
    or g4234 ( n1592 , n5913 , n3450 );
    not g4235 ( n5585 , n3190 );
    or g4236 ( n1702 , n1827 , n4703 );
    and g4237 ( n3112 , n3321 , n4930 );
    and g4238 ( n2264 , n1365 , n2270 );
    not g4239 ( n1832 , n4882 );
    or g4240 ( n455 , n3990 , n6238 );
    nor g4241 ( n6229 , n5961 , n3768 );
    nor g4242 ( n2307 , n4723 , n6131 );
    not g4243 ( n1135 , n581 );
    nor g4244 ( n1577 , n4119 , n5698 );
    not g4245 ( n2431 , n873 );
    nor g4246 ( n5911 , n1590 , n754 );
    and g4247 ( n5523 , n4195 , n6225 );
    nor g4248 ( n719 , n1109 , n1907 );
    or g4249 ( n5552 , n1747 , n40 );
    not g4250 ( n2399 , n383 );
    or g4251 ( n1892 , n3078 , n2057 );
    not g4252 ( n2705 , n4365 );
    or g4253 ( n1454 , n4978 , n1176 );
    not g4254 ( n1319 , n5965 );
    and g4255 ( n4263 , n6120 , n80 );
    and g4256 ( n4380 , n2220 , n3501 );
    nor g4257 ( n5080 , n3671 , n553 );
    not g4258 ( n609 , n494 );
    not g4259 ( n2521 , n374 );
    not g4260 ( n2498 , n2036 );
    or g4261 ( n3331 , n5114 , n5185 );
    or g4262 ( n4209 , n5399 , n872 );
    or g4263 ( n3842 , n1213 , n924 );
    not g4264 ( n3491 , n3519 );
    not g4265 ( n4400 , n929 );
    and g4266 ( n4108 , n4792 , n1409 );
    not g4267 ( n3355 , n1180 );
    or g4268 ( n1320 , n368 , n2427 );
    or g4269 ( n1161 , n2234 , n5231 );
    not g4270 ( n1843 , n1544 );
    or g4271 ( n567 , n4451 , n3166 );
    and g4272 ( n4898 , n5548 , n1397 );
    and g4273 ( n506 , n3432 , n4524 );
    and g4274 ( n109 , n5543 , n3037 );
    or g4275 ( n3232 , n5809 , n3693 );
    or g4276 ( n1921 , n6217 , n3766 );
    or g4277 ( n311 , n199 , n3601 );
    and g4278 ( n107 , n920 , n301 );
    nor g4279 ( n299 , n4010 , n5154 );
    not g4280 ( n5120 , n1471 );
    nor g4281 ( n4024 , n5138 , n2114 );
    not g4282 ( n647 , n5610 );
    or g4283 ( n1234 , n2554 , n459 );
    not g4284 ( n124 , n3380 );
    and g4285 ( n2890 , n4552 , n4534 );
    and g4286 ( n1340 , n2919 , n2264 );
    and g4287 ( n4291 , n2562 , n3150 );
    nor g4288 ( n1098 , n3911 , n2015 );
    or g4289 ( n5002 , n13 , n4812 );
    nor g4290 ( n2539 , n2310 , n3791 );
    or g4291 ( n130 , n5594 , n1305 );
    or g4292 ( n5144 , n3670 , n6215 );
    nor g4293 ( n1482 , n861 , n1523 );
    not g4294 ( n4508 , n300 );
    not g4295 ( n2956 , n147 );
    and g4296 ( n1159 , n765 , n2740 );
    or g4297 ( n3114 , n905 , n1641 );
    not g4298 ( n133 , n628 );
    or g4299 ( n1404 , n3225 , n248 );
    nor g4300 ( n5527 , n2437 , n2671 );
    nor g4301 ( n131 , n4604 , n6243 );
    or g4302 ( n1680 , n3092 , n1299 );
    not g4303 ( n3619 , n147 );
    not g4304 ( n2660 , n882 );
    nor g4305 ( n279 , n2301 , n2882 );
    not g4306 ( n3320 , n963 );
    nor g4307 ( n2779 , n4019 , n5372 );
    not g4308 ( n4241 , n617 );
    or g4309 ( n588 , n2582 , n3925 );
    or g4310 ( n2079 , n2371 , n1236 );
    nor g4311 ( n5846 , n4973 , n2337 );
    or g4312 ( n4152 , n3654 , n2517 );
    not g4313 ( n3535 , n2939 );
    or g4314 ( n2755 , n2934 , n116 );
    not g4315 ( n1164 , n6052 );
    and g4316 ( n1289 , n1394 , n5409 );
    nor g4317 ( n8 , n2056 , n2043 );
    or g4318 ( n517 , n1838 , n5457 );
    or g4319 ( n840 , n822 , n2967 );
    and g4320 ( n650 , n4282 , n4772 );
    or g4321 ( n4062 , n3341 , n2496 );
    or g4322 ( n982 , n2058 , n515 );
    or g4323 ( n5733 , n2993 , n1972 );
    not g4324 ( n3819 , n3712 );
    and g4325 ( n3627 , n5006 , n5444 );
    nor g4326 ( n5124 , n2193 , n1740 );
    or g4327 ( n20 , n2757 , n3104 );
    not g4328 ( n1188 , n1941 );
    and g4329 ( n4651 , n5651 , n2954 );
    or g4330 ( n3376 , n11 , n2044 );
    not g4331 ( n298 , n3957 );
    not g4332 ( n1830 , n2070 );
    nor g4333 ( n5331 , n3566 , n2659 );
    not g4334 ( n2889 , n3464 );
    and g4335 ( n2535 , n1683 , n4327 );
    not g4336 ( n5307 , n432 );
    not g4337 ( n2650 , n887 );
    or g4338 ( n234 , n2747 , n2526 );
    not g4339 ( n5357 , n4948 );
    and g4340 ( n99 , n277 , n997 );
    or g4341 ( n2716 , n2899 , n2886 );
    not g4342 ( n4583 , n4562 );
    not g4343 ( n3220 , n5444 );
    or g4344 ( n1609 , n4354 , n2464 );
    or g4345 ( n2128 , n5179 , n5598 );
    and g4346 ( n2661 , n3271 , n3319 );
    nor g4347 ( n4603 , n1295 , n2292 );
    or g4348 ( n4844 , n5867 , n4865 );
    or g4349 ( n2376 , n597 , n4543 );
    or g4350 ( n5667 , n4601 , n2959 );
    or g4351 ( n3570 , n112 , n4813 );
    nor g4352 ( n3876 , n2146 , n1094 );
    not g4353 ( n942 , n4849 );
    not g4354 ( n5022 , n6217 );
    and g4355 ( n1934 , n4224 , n3129 );
    nor g4356 ( n3072 , n1738 , n14 );
    nor g4357 ( n996 , n4385 , n1097 );
    or g4358 ( n5659 , n3234 , n3119 );
    or g4359 ( n5401 , n689 , n922 );
    or g4360 ( n707 , n1619 , n1344 );
    or g4361 ( n1343 , n5726 , n2527 );
    not g4362 ( n3463 , n5868 );
    nor g4363 ( n359 , n1529 , n3570 );
    not g4364 ( n1493 , n1041 );
    not g4365 ( n150 , n6092 );
    not g4366 ( n1303 , n6248 );
    or g4367 ( n2259 , n2345 , n1347 );
    or g4368 ( n5895 , n524 , n3145 );
    and g4369 ( n4567 , n5845 , n3363 );
    and g4370 ( n706 , n1941 , n2343 );
    not g4371 ( n2344 , n6089 );
    nor g4372 ( n1312 , n351 , n1458 );
    not g4373 ( n2157 , n546 );
    not g4374 ( n1919 , n5997 );
    or g4375 ( n3530 , n2473 , n5313 );
    and g4376 ( n5652 , n4652 , n1196 );
    not g4377 ( n479 , n2554 );
    and g4378 ( n2818 , n980 , n3150 );
    not g4379 ( n1608 , n4584 );
    nor g4380 ( n2152 , n5190 , n5178 );
    or g4381 ( n451 , n5907 , n6272 );
    not g4382 ( n5035 , n5896 );
    nor g4383 ( n3974 , n2801 , n5245 );
    or g4384 ( n3995 , n3838 , n5050 );
    and g4385 ( n503 , n5283 , n4479 );
    or g4386 ( n1949 , n3182 , n5249 );
    nor g4387 ( n4412 , n4664 , n187 );
    not g4388 ( n3624 , n5749 );
    not g4389 ( n2843 , n1195 );
    nor g4390 ( n3902 , n6038 , n3645 );
    or g4391 ( n2824 , n3945 , n6163 );
    nor g4392 ( n4961 , n2216 , n1907 );
    not g4393 ( n5801 , n4196 );
    or g4394 ( n1961 , n3347 , n818 );
    or g4395 ( n2653 , n1137 , n6077 );
    or g4396 ( n2711 , n5091 , n5684 );
    nor g4397 ( n244 , n3701 , n4546 );
    and g4398 ( n3433 , n444 , n4347 );
    or g4399 ( n5871 , n6027 , n5194 );
    and g4400 ( n1859 , n6098 , n4631 );
    not g4401 ( n5981 , n1564 );
    not g4402 ( n2210 , n5538 );
    not g4403 ( n859 , n2925 );
    and g4404 ( n3073 , n2907 , n6288 );
    or g4405 ( n1745 , n4394 , n2779 );
    not g4406 ( n5398 , n4403 );
    and g4407 ( n4804 , n1822 , n129 );
    and g4408 ( n3196 , n4071 , n2633 );
    not g4409 ( n4807 , n4519 );
    or g4410 ( n4276 , n548 , n4768 );
    nor g4411 ( n4022 , n3130 , n2775 );
    or g4412 ( n1749 , n3226 , n5142 );
    or g4413 ( n1683 , n2816 , n1870 );
    and g4414 ( n4952 , n3614 , n388 );
    or g4415 ( n1288 , n4481 , n1713 );
    not g4416 ( n5536 , n3893 );
    not g4417 ( n2217 , n2534 );
    not g4418 ( n1203 , n3000 );
    not g4419 ( n318 , n3509 );
    or g4420 ( n2817 , n642 , n4667 );
    or g4421 ( n3120 , n3317 , n2516 );
    and g4422 ( n1532 , n761 , n2542 );
    nor g4423 ( n1887 , n356 , n342 );
    nor g4424 ( n5598 , n1330 , n2903 );
    or g4425 ( n5607 , n151 , n3901 );
    and g4426 ( n6092 , n6223 , n1248 );
    not g4427 ( n4067 , n4615 );
    and g4428 ( n4731 , n5542 , n5172 );
    not g4429 ( n6018 , n18 );
    or g4430 ( n5804 , n225 , n5621 );
    or g4431 ( n2831 , n2410 , n4914 );
    nor g4432 ( n4641 , n1886 , n1957 );
    not g4433 ( n3781 , n3852 );
    not g4434 ( n5393 , n5798 );
    and g4435 ( n5136 , n4981 , n4723 );
    and g4436 ( n4503 , n3878 , n929 );
    nor g4437 ( n3011 , n1545 , n3628 );
    nor g4438 ( n83 , n3578 , n4492 );
    not g4439 ( n1085 , n4983 );
    nor g4440 ( n5139 , n3335 , n5552 );
    or g4441 ( n1559 , n4414 , n6094 );
    and g4442 ( n964 , n2123 , n1705 );
    not g4443 ( n799 , n4164 );
    not g4444 ( n2395 , n3984 );
    or g4445 ( n2564 , n4888 , n1396 );
    not g4446 ( n3702 , n1984 );
    or g4447 ( n2601 , n5657 , n2725 );
    or g4448 ( n1492 , n6074 , n1212 );
    and g4449 ( n3859 , n4053 , n200 );
    not g4450 ( n352 , n3122 );
    or g4451 ( n2829 , n121 , n3821 );
    not g4452 ( n1967 , n103 );
    or g4453 ( n2488 , n3166 , n5749 );
    not g4454 ( n2532 , n6004 );
    nor g4455 ( n3986 , n4867 , n3810 );
    or g4456 ( n1286 , n6231 , n6278 );
    and g4457 ( n5215 , n4651 , n5625 );
    or g4458 ( n3744 , n2840 , n3976 );
    nor g4459 ( n5526 , n5589 , n3445 );
    nor g4460 ( n2158 , n103 , n1936 );
    not g4461 ( n1617 , n4417 );
    or g4462 ( n3385 , n2069 , n4959 );
    not g4463 ( n5358 , n3699 );
    nor g4464 ( n2037 , n5654 , n1060 );
    not g4465 ( n5830 , n2533 );
    or g4466 ( n4907 , n555 , n4205 );
    nor g4467 ( n1519 , n4490 , n5630 );
    not g4468 ( n2990 , n3548 );
    or g4469 ( n2390 , n5364 , n5458 );
    or g4470 ( n1955 , n4960 , n2314 );
    nor g4471 ( n1517 , n4707 , n4682 );
    nor g4472 ( n5648 , n5666 , n3173 );
    nor g4473 ( n1719 , n4020 , n533 );
    or g4474 ( n3882 , n4353 , n1367 );
    not g4475 ( n3597 , n5354 );
    and g4476 ( n11 , n4194 , n5514 );
    or g4477 ( n1498 , n4339 , n211 );
    and g4478 ( n5436 , n5288 , n2440 );
    nor g4479 ( n2823 , n5763 , n1263 );
    and g4480 ( n5086 , n617 , n2519 );
    nor g4481 ( n5071 , n126 , n821 );
    not g4482 ( n6131 , n679 );
    or g4483 ( n5195 , n3607 , n4588 );
    or g4484 ( n3724 , n1113 , n5373 );
    nor g4485 ( n1077 , n1776 , n5846 );
    and g4486 ( n536 , n2054 , n3111 );
    and g4487 ( n2636 , n1038 , n521 );
    or g4488 ( n2598 , n4881 , n1351 );
    not g4489 ( n5336 , n5408 );
    or g4490 ( n1873 , n1220 , n945 );
    not g4491 ( n582 , n2016 );
    nor g4492 ( n5958 , n1549 , n2009 );
    nor g4493 ( n4300 , n1471 , n4637 );
    or g4494 ( n4975 , n6068 , n5399 );
    or g4495 ( n5729 , n2227 , n6073 );
    or g4496 ( n1059 , n100 , n1011 );
    nor g4497 ( n3236 , n3096 , n4056 );
    or g4498 ( n1350 , n4997 , n5981 );
    not g4499 ( n4016 , n36 );
    or g4500 ( n5013 , n830 , n3620 );
    nor g4501 ( n2203 , n4448 , n471 );
    nor g4502 ( n361 , n4098 , n225 );
    and g4503 ( n2242 , n3012 , n4876 );
    nor g4504 ( n3737 , n5013 , n3311 );
    nor g4505 ( n5206 , n868 , n5356 );
    or g4506 ( n3054 , n3175 , n5221 );
    or g4507 ( n5055 , n99 , n2619 );
    or g4508 ( n5653 , n623 , n1281 );
    and g4509 ( n4870 , n3196 , n1440 );
    and g4510 ( n5945 , n609 , n3389 );
    not g4511 ( n1342 , n5418 );
    or g4512 ( n2024 , n3948 , n1672 );
    nor g4513 ( n283 , n794 , n3487 );
    nor g4514 ( n2298 , n2172 , n4775 );
    not g4515 ( n1158 , n2840 );
    or g4516 ( n3888 , n819 , n6262 );
    or g4517 ( n2854 , n4186 , n5361 );
    nor g4518 ( n894 , n1645 , n5880 );
    and g4519 ( n3231 , n4709 , n2321 );
    and g4520 ( n6277 , n5257 , n4514 );
    not g4521 ( n2643 , n4362 );
    nor g4522 ( n1736 , n4658 , n852 );
    not g4523 ( n3477 , n1057 );
    not g4524 ( n3022 , n3281 );
    and g4525 ( n4326 , n3572 , n5148 );
    nor g4526 ( n961 , n4550 , n2293 );
    not g4527 ( n4745 , n2453 );
    or g4528 ( n3428 , n4586 , n5158 );
    or g4529 ( n2683 , n1075 , n149 );
    and g4530 ( n585 , n3527 , n1327 );
    not g4531 ( n3135 , n240 );
    or g4532 ( n398 , n2777 , n235 );
    and g4533 ( n1791 , n4361 , n5063 );
    or g4534 ( n2621 , n4100 , n210 );
    not g4535 ( n4005 , n480 );
    nor g4536 ( n4865 , n4271 , n44 );
    and g4537 ( n3378 , n2101 , n2428 );
    and g4538 ( n2394 , n2128 , n3330 );
    or g4539 ( n1022 , n2378 , n4460 );
    not g4540 ( n4430 , n4790 );
    or g4541 ( n1527 , n4403 , n3564 );
    and g4542 ( n4107 , n1495 , n4468 );
    or g4543 ( n5651 , n1290 , n5997 );
    or g4544 ( n3068 , n5134 , n1832 );
    not g4545 ( n1696 , n2676 );
    and g4546 ( n644 , n2728 , n2347 );
    and g4547 ( n1837 , n5677 , n5927 );
    or g4548 ( n1677 , n4021 , n1355 );
    or g4549 ( n5414 , n2489 , n3958 );
    nor g4550 ( n1694 , n5899 , n1496 );
    not g4551 ( n6015 , n944 );
    or g4552 ( n5232 , n1440 , n2374 );
    and g4553 ( n4427 , n1036 , n2266 );
    and g4554 ( n6138 , n6080 , n2567 );
    and g4555 ( n5747 , n3572 , n1425 );
    or g4556 ( n4741 , n3169 , n3688 );
    nor g4557 ( n16 , n327 , n3032 );
    or g4558 ( n5898 , n3106 , n5615 );
    or g4559 ( n4040 , n5678 , n3998 );
    and g4560 ( n1777 , n3428 , n2455 );
    not g4561 ( n3119 , n4147 );
    nor g4562 ( n1450 , n301 , n6041 );
    or g4563 ( n1759 , n6073 , n4564 );
    nor g4564 ( n3886 , n4115 , n4716 );
    and g4565 ( n3092 , n4191 , n4044 );
    not g4566 ( n2816 , n2255 );
    not g4567 ( n1170 , n4196 );
    or g4568 ( n1065 , n2678 , n60 );
    not g4569 ( n2150 , n376 );
    not g4570 ( n702 , n3084 );
    and g4571 ( n141 , n3937 , n4305 );
    and g4572 ( n3035 , n4926 , n1258 );
    or g4573 ( n2792 , n4539 , n3837 );
    not g4574 ( n1540 , n644 );
    nor g4575 ( n3839 , n2871 , n6146 );
    not g4576 ( n2634 , n3167 );
    or g4577 ( n2269 , n2625 , n182 );
    not g4578 ( n39 , n3285 );
    not g4579 ( n3193 , n2588 );
    and g4580 ( n3612 , n3043 , n2814 );
    nor g4581 ( n5551 , n4332 , n1813 );
    or g4582 ( n1143 , n2804 , n4743 );
    not g4583 ( n425 , n5723 );
    nor g4584 ( n748 , n78 , n5617 );
    or g4585 ( n4429 , n4502 , n1463 );
    not g4586 ( n4695 , n1091 );
    not g4587 ( n3643 , n2221 );
    nor g4588 ( n282 , n271 , n110 );
    nor g4589 ( n3434 , n548 , n2003 );
    and g4590 ( n3010 , n4320 , n5196 );
    or g4591 ( n5957 , n837 , n4104 );
    nor g4592 ( n3500 , n4050 , n2965 );
    and g4593 ( n5919 , n1339 , n1269 );
    and g4594 ( n5488 , n5891 , n1770 );
    nor g4595 ( n1580 , n3140 , n2733 );
    or g4596 ( n5504 , n4253 , n1742 );
    or g4597 ( n2188 , n1349 , n5913 );
    nor g4598 ( n348 , n4425 , n1655 );
    and g4599 ( n5155 , n2385 , n755 );
    and g4600 ( n5467 , n2740 , n1427 );
    not g4601 ( n1271 , n869 );
    and g4602 ( n5387 , n2013 , n3466 );
    or g4603 ( n1025 , n4866 , n6052 );
    not g4604 ( n2505 , n786 );
    or g4605 ( n2828 , n3336 , n4979 );
    and g4606 ( n5813 , n61 , n1234 );
    not g4607 ( n118 , n2153 );
    not g4608 ( n6027 , n4805 );
    and g4609 ( n3548 , n2787 , n6301 );
    not g4610 ( n4761 , n212 );
    or g4611 ( n5125 , n2785 , n771 );
    and g4612 ( n5193 , n2985 , n6118 );
    not g4613 ( n3080 , n5228 );
    and g4614 ( n1227 , n1787 , n1318 );
    nor g4615 ( n2204 , n4454 , n2759 );
    and g4616 ( n2361 , n6046 , n2299 );
    not g4617 ( n825 , n5032 );
    not g4618 ( n3079 , n3829 );
    not g4619 ( n606 , n452 );
    not g4620 ( n3589 , n5750 );
    or g4621 ( n264 , n6186 , n263 );
    not g4622 ( n3058 , n1588 );
    and g4623 ( n3756 , n5423 , n6223 );
    not g4624 ( n1318 , n4735 );
    nor g4625 ( n697 , n4979 , n3552 );
    nor g4626 ( n3537 , n2160 , n4738 );
    or g4627 ( n1935 , n3413 , n1103 );
    nor g4628 ( n3562 , n1294 , n5108 );
    and g4629 ( n3852 , n3426 , n318 );
    nor g4630 ( n6260 , n1004 , n3342 );
    not g4631 ( n658 , n4595 );
    not g4632 ( n2078 , n1457 );
    or g4633 ( n2793 , n4674 , n4252 );
    not g4634 ( n1516 , n2305 );
    nor g4635 ( n1957 , n5463 , n5863 );
    or g4636 ( n2189 , n1714 , n5490 );
    not g4637 ( n1045 , n5177 );
    and g4638 ( n5003 , n5243 , n2969 );
    and g4639 ( n3896 , n5156 , n6201 );
    and g4640 ( n6233 , n4428 , n2229 );
    not g4641 ( n3103 , n1690 );
    not g4642 ( n721 , n5596 );
    and g4643 ( n5765 , n195 , n352 );
    and g4644 ( n617 , n5209 , n2533 );
    not g4645 ( n6167 , n3687 );
    not g4646 ( n5517 , n4776 );
    not g4647 ( n5510 , n4752 );
    or g4648 ( n583 , n2735 , n2212 );
    not g4649 ( n3497 , n4297 );
    nor g4650 ( n2987 , n4777 , n5366 );
    nor g4651 ( n635 , n1885 , n1921 );
    and g4652 ( n4626 , n501 , n2572 );
    nor g4653 ( n502 , n2349 , n5415 );
    not g4654 ( n1293 , n1964 );
    or g4655 ( n4573 , n2320 , n6179 );
    or g4656 ( n5874 , n2829 , n1467 );
    and g4657 ( n784 , n919 , n4771 );
    not g4658 ( n1726 , n890 );
    nor g4659 ( n4642 , n4254 , n684 );
    nor g4660 ( n5360 , n366 , n3987 );
    or g4661 ( n1301 , n1419 , n5712 );
    not g4662 ( n304 , n6277 );
    or g4663 ( n1347 , n1898 , n443 );
    nor g4664 ( n5180 , n165 , n3808 );
    nor g4665 ( n3358 , n3767 , n5083 );
    or g4666 ( n5984 , n5597 , n1922 );
    nor g4667 ( n1253 , n540 , n5642 );
    or g4668 ( n6024 , n1173 , n415 );
    and g4669 ( n3929 , n619 , n3372 );
    nor g4670 ( n1174 , n1889 , n5229 );
    or g4671 ( n4851 , n2196 , n3924 );
    nor g4672 ( n1913 , n2649 , n5017 );
    nor g4673 ( n5033 , n3813 , n3490 );
    and g4674 ( n2056 , n838 , n2377 );
    or g4675 ( n3036 , n889 , n1793 );
    not g4676 ( n2526 , n810 );
    or g4677 ( n4908 , n3355 , n62 );
    and g4678 ( n4995 , n3224 , n951 );
    not g4679 ( n6159 , n4110 );
    nor g4680 ( n4118 , n1215 , n2843 );
    or g4681 ( n2048 , n1052 , n801 );
    and g4682 ( n5839 , n5513 , n5665 );
    not g4683 ( n602 , n4336 );
    or g4684 ( n250 , n5931 , n2529 );
    nor g4685 ( n5321 , n6235 , n976 );
    not g4686 ( n4686 , n5262 );
    or g4687 ( n4924 , n4560 , n2844 );
    not g4688 ( n5226 , n4425 );
    and g4689 ( n5159 , n4726 , n5288 );
    or g4690 ( n3811 , n4083 , n3634 );
    or g4691 ( n4784 , n3278 , n2041 );
    and g4692 ( n5678 , n4184 , n3904 );
    not g4693 ( n527 , n3748 );
    or g4694 ( n3608 , n2508 , n5525 );
    not g4695 ( n2021 , n4811 );
    nor g4696 ( n3528 , n626 , n2379 );
    nor g4697 ( n1551 , n142 , n5980 );
    and g4698 ( n429 , n1566 , n2227 );
    or g4699 ( n745 , n5110 , n741 );
    not g4700 ( n372 , n3188 );
    and g4701 ( n3413 , n4657 , n4486 );
    and g4702 ( n4516 , n1594 , n6105 );
    or g4703 ( n2701 , n2444 , n4766 );
    and g4704 ( n4845 , n3389 , n6203 );
    or g4705 ( n3599 , n3848 , n3306 );
    and g4706 ( n4379 , n4259 , n5190 );
    and g4707 ( n300 , n3080 , n2107 );
    or g4708 ( n176 , n6227 , n568 );
    not g4709 ( n3449 , n3347 );
    nor g4710 ( n4019 , n3355 , n6065 );
    or g4711 ( n114 , n2744 , n1255 );
    not g4712 ( n4178 , n3226 );
    or g4713 ( n5247 , n4111 , n5290 );
    and g4714 ( n3640 , n4198 , n3797 );
    not g4715 ( n3172 , n4071 );
    or g4716 ( n3976 , n5233 , n4891 );
    nor g4717 ( n6243 , n1512 , n4905 );
    not g4718 ( n877 , n4580 );
    or g4719 ( n5869 , n5077 , n3093 );
    not g4720 ( n4061 , n1890 );
    or g4721 ( n1435 , n1154 , n2222 );
    or g4722 ( n4320 , n3363 , n10 );
    not g4723 ( n2139 , n612 );
    not g4724 ( n137 , n191 );
    and g4725 ( n254 , n2217 , n4451 );
    or g4726 ( n714 , n3687 , n3433 );
    or g4727 ( n221 , n3654 , n4610 );
    nor g4728 ( n6039 , n5496 , n6008 );
    or g4729 ( n4779 , n3000 , n363 );
    or g4730 ( n2138 , n334 , n3997 );
    not g4731 ( n2085 , n1001 );
    or g4732 ( n5734 , n2449 , n902 );
    or g4733 ( n5078 , n3447 , n933 );
    or g4734 ( n2458 , n4364 , n3636 );
    nor g4735 ( n1127 , n4241 , n2838 );
    or g4736 ( n5118 , n4721 , n4213 );
    and g4737 ( n3906 , n3933 , n3614 );
    not g4738 ( n1537 , n3543 );
    not g4739 ( n3131 , n1949 );
    or g4740 ( n969 , n4175 , n5164 );
    nor g4741 ( n1700 , n2979 , n1701 );
    not g4742 ( n3128 , n5616 );
    not g4743 ( n5208 , n4510 );
    and g4744 ( n2363 , n820 , n2150 );
    or g4745 ( n2699 , n5263 , n3476 );
    nor g4746 ( n2983 , n5856 , n5256 );
    not g4747 ( n1536 , n2787 );
    not g4748 ( n1526 , n581 );
    or g4749 ( n3025 , n658 , n2392 );
    or g4750 ( n4799 , n4789 , n1272 );
    not g4751 ( n6113 , n3286 );
    not g4752 ( n1956 , n3513 );
    and g4753 ( n5606 , n1095 , n3871 );
    and g4754 ( n2756 , n4634 , n2111 );
    and g4755 ( n4293 , n5855 , n562 );
    not g4756 ( n1362 , n2751 );
    and g4757 ( n898 , n4948 , n4848 );
    or g4758 ( n1241 , n2890 , n3179 );
    not g4759 ( n5744 , n314 );
    and g4760 ( n4078 , n4152 , n650 );
    or g4761 ( n6250 , n429 , n2662 );
    or g4762 ( n2928 , n4235 , n473 );
    nor g4763 ( n214 , n5533 , n2932 );
    not g4764 ( n3779 , n1337 );
    not g4765 ( n3549 , n1371 );
    not g4766 ( n1173 , n5706 );
    nor g4767 ( n2314 , n2607 , n1558 );
    not g4768 ( n944 , n560 );
    nor g4769 ( n414 , n3349 , n1115 );
    not g4770 ( n4146 , n3815 );
    and g4771 ( n5723 , n1809 , n6111 );
    and g4772 ( n750 , n2559 , n457 );
    nor g4773 ( n5458 , n281 , n2450 );
    and g4774 ( n2677 , n6071 , n168 );
    not g4775 ( n2930 , n526 );
    or g4776 ( n277 , n781 , n3168 );
    and g4777 ( n2221 , n218 , n3009 );
    or g4778 ( n1662 , n4483 , n739 );
    not g4779 ( n5732 , n399 );
    not g4780 ( n2916 , n734 );
    not g4781 ( n32 , n5872 );
    not g4782 ( n2326 , n6192 );
    and g4783 ( n1196 , n2214 , n5808 );
    or g4784 ( n607 , n5802 , n6160 );
    and g4785 ( n2520 , n3151 , n2120 );
    and g4786 ( n1307 , n791 , n2111 );
    and g4787 ( n1709 , n2140 , n5188 );
    and g4788 ( n670 , n2162 , n1384 );
    or g4789 ( n3014 , n361 , n5253 );
    or g4790 ( n3983 , n4434 , n1038 );
    and g4791 ( n1594 , n2800 , n6120 );
    and g4792 ( n2972 , n1261 , n2453 );
    not g4793 ( n1207 , n3608 );
    or g4794 ( n5713 , n5820 , n5612 );
    or g4795 ( n5394 , n444 , n1650 );
    or g4796 ( n2977 , n5784 , n4966 );
    nor g4797 ( n1322 , n2390 , n5828 );
    not g4798 ( n5027 , n2289 );
    not g4799 ( n5649 , n3754 );
    nor g4800 ( n5964 , n623 , n3875 );
    not g4801 ( n5566 , n3307 );
    nor g4802 ( n2540 , n243 , n430 );
    nor g4803 ( n5554 , n4356 , n3424 );
    or g4804 ( n132 , n4850 , n3917 );
    nor g4805 ( n5592 , n696 , n4375 );
    or g4806 ( n3826 , n4303 , n369 );
    and g4807 ( n4524 , n2469 , n5307 );
    not g4808 ( n5599 , n2349 );
    not g4809 ( n6200 , n2194 );
    not g4810 ( n5386 , n3055 );
    or g4811 ( n1531 , n1165 , n901 );
    or g4812 ( n5001 , n2415 , n1403 );
    not g4813 ( n5288 , n5906 );
    and g4814 ( n4345 , n3218 , n3950 );
    nor g4815 ( n2940 , n2093 , n5226 );
    and g4816 ( n6242 , n5837 , n5785 );
    not g4817 ( n2512 , n2279 );
    or g4818 ( n4840 , n4177 , n1155 );
    and g4819 ( n2658 , n3047 , n1265 );
    and g4820 ( n2465 , n5839 , n1181 );
    not g4821 ( n5095 , n2744 );
    not g4822 ( n911 , n2552 );
    or g4823 ( n608 , n1251 , n5078 );
    or g4824 ( n5586 , n2565 , n1772 );
    not g4825 ( n379 , n1244 );
    not g4826 ( n86 , n6303 );
    not g4827 ( n212 , n899 );
    or g4828 ( n4996 , n4590 , n265 );
    and g4829 ( n5329 , n3454 , n3583 );
    nor g4830 ( n89 , n3690 , n2899 );
    and g4831 ( n2763 , n4351 , n2160 );
    nor g4832 ( n402 , n5028 , n2435 );
    not g4833 ( n613 , n5548 );
    and g4834 ( n6225 , n1541 , n6219 );
    or g4835 ( n1552 , n6150 , n962 );
    not g4836 ( n3806 , n5750 );
    or g4837 ( n6134 , n2428 , n3555 );
    not g4838 ( n2244 , n3233 );
    not g4839 ( n278 , n3606 );
    not g4840 ( n2882 , n1905 );
    nor g4841 ( n667 , n1485 , n4377 );
    and g4842 ( n3088 , n5946 , n1602 );
    not g4843 ( n4874 , n411 );
    or g4844 ( n5449 , n594 , n4517 );
    nor g4845 ( n3118 , n3726 , n6121 );
    not g4846 ( n5412 , n369 );
    and g4847 ( n5480 , n3331 , n6123 );
    nor g4848 ( n4624 , n201 , n4527 );
    nor g4849 ( n855 , n1546 , n2499 );
    or g4850 ( n5334 , n2145 , n4679 );
    nor g4851 ( n1720 , n2534 , n1981 );
    or g4852 ( n4417 , n3835 , n1125 );
    nor g4853 ( n48 , n1613 , n182 );
    not g4854 ( n4742 , n1036 );
    not g4855 ( n4756 , n2276 );
    and g4856 ( n1727 , n2018 , n5945 );
    or g4857 ( n4377 , n2644 , n1361 );
    and g4858 ( n287 , n1391 , n695 );
    or g4859 ( n3245 , n3250 , n4018 );
    nor g4860 ( n4931 , n327 , n4687 );
    not g4861 ( n4919 , n1861 );
    and g4862 ( n3671 , n4144 , n3328 );
    not g4863 ( n1357 , n977 );
    or g4864 ( n3937 , n3810 , n3099 );
    nor g4865 ( n5943 , n2490 , n1902 );
    and g4866 ( n1102 , n3684 , n2832 );
    or g4867 ( n4042 , n1426 , n2689 );
    not g4868 ( n2924 , n3884 );
    and g4869 ( n4954 , n5908 , n5323 );
    nor g4870 ( n3291 , n1389 , n2906 );
    or g4871 ( n4862 , n4870 , n2011 );
    not g4872 ( n1643 , n91 );
    nor g4873 ( n2912 , n3062 , n123 );
    or g4874 ( n3892 , n133 , n5822 );
    and g4875 ( n1267 , n3065 , n1696 );
    and g4876 ( n3942 , n4052 , n4602 );
    not g4877 ( n5688 , n2524 );
    and g4878 ( n192 , n1386 , n1057 );
    and g4879 ( n5893 , n3047 , n4636 );
    not g4880 ( n4246 , n4130 );
    nor g4881 ( n6040 , n5358 , n2992 );
    or g4882 ( n3276 , n1216 , n427 );
    not g4883 ( n4207 , n432 );
    or g4884 ( n4094 , n3444 , n4988 );
    not g4885 ( n1864 , n2914 );
    nor g4886 ( n5083 , n3156 , n54 );
    and g4887 ( n4842 , n416 , n806 );
    and g4888 ( n4484 , n3461 , n4697 );
    or g4889 ( n1266 , n4888 , n4023 );
    or g4890 ( n3081 , n2039 , n2316 );
    or g4891 ( n5270 , n2419 , n1963 );
    not g4892 ( n2747 , n3209 );
    nor g4893 ( n1682 , n4665 , n312 );
    not g4894 ( n2835 , n5640 );
    or g4895 ( n1013 , n4916 , n9 );
    nor g4896 ( n1962 , n2425 , n1899 );
    nor g4897 ( n3246 , n587 , n5877 );
    nor g4898 ( n6125 , n2456 , n2881 );
    or g4899 ( n4558 , n3802 , n2590 );
    nor g4900 ( n5899 , n4547 , n1192 );
    or g4901 ( n2646 , n2466 , n893 );
    and g4902 ( n417 , n3584 , n2860 );
    not g4903 ( n559 , n4472 );
    not g4904 ( n4003 , n2142 );
    not g4905 ( n1428 , n2104 );
    nor g4906 ( n2443 , n3037 , n3624 );
    or g4907 ( n520 , n4887 , n3358 );
    and g4908 ( n518 , n1575 , n2372 );
    and g4909 ( n3780 , n1823 , n4494 );
    and g4910 ( n5544 , n3010 , n4146 );
    not g4911 ( n2500 , n4584 );
    or g4912 ( n2953 , n5139 , n3676 );
    or g4913 ( n119 , n1475 , n1279 );
    not g4914 ( n2417 , n3436 );
    not g4915 ( n1348 , n4310 );
    and g4916 ( n1564 , n2674 , n6211 );
    nor g4917 ( n822 , n5654 , n4734 );
    not g4918 ( n3672 , n1958 );
    nor g4919 ( n81 , n5490 , n3807 );
    nor g4920 ( n5368 , n4727 , n5540 );
    nor g4921 ( n5642 , n2835 , n1938 );
    nor g4922 ( n325 , n111 , n4421 );
    and g4923 ( n6239 , n117 , n4165 );
    and g4924 ( n3647 , n2430 , n5884 );
    nor g4925 ( n514 , n4238 , n2130 );
    not g4926 ( n1780 , n842 );
    nor g4927 ( n5983 , n4186 , n3134 );
    and g4928 ( n2706 , n5163 , n4369 );
    nor g4929 ( n4069 , n3366 , n2182 );
    nor g4930 ( n2690 , n367 , n5298 );
    not g4931 ( n759 , n2467 );
    not g4932 ( n3363 , n6224 );
    and g4933 ( n3670 , n3475 , n1128 );
    and g4934 ( n4483 , n5026 , n4268 );
    nor g4935 ( n4780 , n3489 , n2585 );
    not g4936 ( n5998 , n5819 );
    not g4937 ( n1827 , n1809 );
    or g4938 ( n1619 , n3451 , n4058 );
    or g4939 ( n1717 , n5836 , n1405 );
    or g4940 ( n501 , n6053 , n4418 );
    or g4941 ( n2438 , n4429 , n946 );
    and g4942 ( n5302 , n3843 , n986 );
    not g4943 ( n4885 , n4626 );
    or g4944 ( n768 , n2833 , n5227 );
    and g4945 ( n901 , n5582 , n3931 );
    or g4946 ( n4318 , n5051 , n1835 );
    and g4947 ( n4893 , n1473 , n2465 );
    or g4948 ( n1394 , n1218 , n2927 );
    or g4949 ( n5154 , n4769 , n2 );
    nor g4950 ( n4008 , n2004 , n4337 );
    not g4951 ( n5130 , n2973 );
    or g4952 ( n5639 , n3992 , n2853 );
    nor g4953 ( n3674 , n2918 , n4153 );
    or g4954 ( n2293 , n2569 , n1222 );
    nor g4955 ( n2290 , n6256 , n3416 );
    nor g4956 ( n5719 , n4433 , n5268 );
    nor g4957 ( n3790 , n2569 , n1126 );
    not g4958 ( n1649 , n5965 );
    and g4959 ( n3567 , n5141 , n5426 );
    nor g4960 ( n4013 , n190 , n4449 );
    not g4961 ( n3258 , n3510 );
    or g4962 ( n1898 , n1783 , n3597 );
    not g4963 ( n2585 , n1888 );
    or g4964 ( n248 , n16 , n832 );
    and g4965 ( n2734 , n2461 , n2413 );
    not g4966 ( n4829 , n4448 );
    not g4967 ( n1521 , n1428 );
    nor g4968 ( n3566 , n4997 , n4830 );
    not g4969 ( n2935 , n5825 );
    not g4970 ( n408 , n1207 );
    not g4971 ( n2985 , n2335 );
    or g4972 ( n6081 , n1592 , n5571 );
    and g4973 ( n5707 , n1192 , n2500 );
    nor g4974 ( n1646 , n4537 , n2304 );
    not g4975 ( n4854 , n2649 );
    nor g4976 ( n1110 , n5391 , n5348 );
    or g4977 ( n286 , n2497 , n5287 );
    not g4978 ( n2491 , n4117 );
    not g4979 ( n71 , n3474 );
    or g4980 ( n3508 , n1790 , n5494 );
    or g4981 ( n4839 , n2859 , n5601 );
    nor g4982 ( n2068 , n5861 , n4127 );
    nor g4983 ( n2278 , n3589 , n6140 );
    and g4984 ( n2246 , n5385 , n4575 );
    not g4985 ( n1128 , n4754 );
    not g4986 ( n5111 , n4356 );
    not g4987 ( n4431 , n1980 );
    and g4988 ( n257 , n3710 , n3939 );
    and g4989 ( n3343 , n4123 , n681 );
    and g4990 ( n2739 , n566 , n1114 );
    or g4991 ( n1734 , n239 , n1684 );
    or g4992 ( n5239 , n4520 , n2183 );
    not g4993 ( n5097 , n1924 );
    not g4994 ( n5810 , n2735 );
    not g4995 ( n3909 , n4678 );
    and g4996 ( n1477 , n5891 , n3260 );
    or g4997 ( n3694 , n1384 , n898 );
    or g4998 ( n1883 , n6267 , n4661 );
    not g4999 ( n5323 , n5127 );
    not g5000 ( n5041 , n3835 );
    buf g5001 ( n3849 , n2016 );
    or g5002 ( n1684 , n2097 , n5489 );
    not g5003 ( n701 , n5628 );
    or g5004 ( n3766 , n5477 , n2334 );
    not g5005 ( n4222 , n4334 );
    not g5006 ( n5706 , n5256 );
    not g5007 ( n3699 , n5193 );
    not g5008 ( n4900 , n2559 );
    not g5009 ( n168 , n3744 );
    not g5010 ( n2404 , n1302 );
    nor g5011 ( n3383 , n3907 , n3962 );
    or g5012 ( n1449 , n1731 , n6163 );
    or g5013 ( n4465 , n1280 , n1031 );
    or g5014 ( n4936 , n5926 , n4916 );
    or g5015 ( n5737 , n1761 , n2736 );
    or g5016 ( n1272 , n2963 , n3908 );
    and g5017 ( n356 , n6185 , n2120 );
    nor g5018 ( n496 , n2672 , n3961 );
    not g5019 ( n1330 , n5986 );
    nor g5020 ( n5061 , n1439 , n470 );
    or g5021 ( n5902 , n954 , n5056 );
    or g5022 ( n1315 , n1372 , n6060 );
    not g5023 ( n3431 , n1420 );
    or g5024 ( n2597 , n5086 , n1173 );
    not g5025 ( n2877 , n4625 );
    and g5026 ( n4000 , n3217 , n1791 );
    and g5027 ( n347 , n6230 , n1313 );
    and g5028 ( n4208 , n1580 , n4341 );
    or g5029 ( n5400 , n5479 , n3617 );
    nor g5030 ( n5546 , n1082 , n5313 );
    not g5031 ( n4498 , n3448 );
    not g5032 ( n1152 , n3171 );
    or g5033 ( n67 , n821 , n3075 );
    and g5034 ( n2657 , n6226 , n744 );
    not g5035 ( n5970 , n5864 );
    and g5036 ( n4203 , n1765 , n5986 );
    not g5037 ( n2695 , n5900 );
    nor g5038 ( n793 , n3320 , n1499 );
    and g5039 ( n4714 , n4178 , n3660 );
    not g5040 ( n6248 , n3162 );
    or g5041 ( n6178 , n830 , n4673 );
    nor g5042 ( n5923 , n2696 , n664 );
    or g5043 ( n1041 , n5450 , n573 );
    nor g5044 ( n3897 , n4218 , n600 );
    nor g5045 ( n853 , n4536 , n2768 );
    or g5046 ( n5870 , n5499 , n2963 );
    or g5047 ( n2786 , n936 , n2944 );
    nor g5048 ( n2966 , n618 , n4635 );
    not g5049 ( n2888 , n4086 );
    or g5050 ( n2676 , n628 , n3001 );
    and g5051 ( n2102 , n446 , n6214 );
    or g5052 ( n12 , n137 , n6205 );
    not g5053 ( n4964 , n4467 );
    nor g5054 ( n1699 , n4212 , n5163 );
    nor g5055 ( n3536 , n387 , n3286 );
    or g5056 ( n3365 , n4735 , n2551 );
    or g5057 ( n2917 , n1850 , n3 );
    nor g5058 ( n1230 , n5421 , n3309 );
    nor g5059 ( n3592 , n3575 , n4611 );
    or g5060 ( n5354 , n1654 , n3940 );
    not g5061 ( n3361 , n1189 );
    or g5062 ( n4569 , n5736 , n1961 );
    not g5063 ( n994 , n2400 );
    and g5064 ( n2826 , n451 , n3802 );
    nor g5065 ( n2778 , n4454 , n2987 );
    or g5066 ( n564 , n2360 , n5611 );
    not g5067 ( n1626 , n2980 );
    or g5068 ( n2722 , n5668 , n3119 );
    or g5069 ( n4442 , n5670 , n5363 );
    nor g5070 ( n2896 , n6210 , n3920 );
    nor g5071 ( n2226 , n867 , n5135 );
    or g5072 ( n3552 , n4909 , n5330 );
    and g5073 ( n2668 , n1379 , n2564 );
    nor g5074 ( n2476 , n1972 , n799 );
    nor g5075 ( n4227 , n5277 , n1186 );
    nor g5076 ( n5223 , n2132 , n4856 );
    and g5077 ( n2719 , n2235 , n2144 );
    or g5078 ( n2215 , n390 , n5629 );
    or g5079 ( n5349 , n2808 , n6136 );
    not g5080 ( n4613 , n410 );
    not g5081 ( n2306 , n1767 );
    or g5082 ( n1748 , n1568 , n3812 );
    nor g5083 ( n3132 , n4729 , n2460 );
    or g5084 ( n4477 , n5102 , n1905 );
    or g5085 ( n3027 , n530 , n5039 );
    not g5086 ( n6122 , n2884 );
    not g5087 ( n1924 , n1707 );
    not g5088 ( n2081 , n5829 );
    or g5089 ( n4546 , n5732 , n292 );
    not g5090 ( n4932 , n113 );
    not g5091 ( n1044 , n6154 );
    not g5092 ( n5881 , n4703 );
    not g5093 ( n5704 , n2819 );
    nor g5094 ( n1858 , n4495 , n1504 );
    or g5095 ( n3650 , n1519 , n6015 );
    and g5096 ( n219 , n3035 , n3978 );
    nor g5097 ( n2009 , n1056 , n5034 );
    or g5098 ( n5181 , n6263 , n2657 );
    not g5099 ( n6001 , n6053 );
    not g5100 ( n960 , n5843 );
    and g5101 ( n4520 , n2087 , n4487 );
    not g5102 ( n4392 , n3174 );
    nor g5103 ( n3590 , n2390 , n827 );
    and g5104 ( n5209 , n2137 , n5281 );
    and g5105 ( n5882 , n2817 , n3378 );
    not g5106 ( n3992 , n3644 );
    nor g5107 ( n3880 , n1591 , n2096 );
    not g5108 ( n5939 , n57 );
    and g5109 ( n4639 , n5806 , n4952 );
    and g5110 ( n2279 , n3019 , n410 );
    or g5111 ( n1461 , n778 , n468 );
    nor g5112 ( n4950 , n2919 , n299 );
    or g5113 ( n4077 , n948 , n3526 );
    or g5114 ( n2480 , n2826 , n2061 );
    or g5115 ( n6192 , n4538 , n5746 );
    nor g5116 ( n3467 , n5117 , n5553 );
    not g5117 ( n384 , n3089 );
    and g5118 ( n3848 , n2188 , n1649 );
    and g5119 ( n1359 , n3483 , n5000 );
    or g5120 ( n2791 , n1257 , n205 );
    or g5121 ( n6244 , n3604 , n4732 );
    and g5122 ( n6155 , n507 , n4933 );
    or g5123 ( n2178 , n5134 , n3004 );
    nor g5124 ( n1291 , n1527 , n1551 );
    nor g5125 ( n5994 , n3030 , n6122 );
    and g5126 ( n5364 , n1047 , n5578 );
    or g5127 ( n3820 , n4694 , n3337 );
    nor g5128 ( n3018 , n5011 , n2116 );
    nor g5129 ( n757 , n2809 , n3313 );
    or g5130 ( n5169 , n3991 , n2275 );
    and g5131 ( n2978 , n5087 , n1191 );
    or g5132 ( n344 , n3213 , n6112 );
    not g5133 ( n6088 , n1431 );
    nor g5134 ( n4171 , n5830 , n646 );
    or g5135 ( n4933 , n3349 , n3989 );
    nor g5136 ( n5676 , n897 , n1572 );
    or g5137 ( n2206 , n2184 , n655 );
    or g5138 ( n3609 , n5074 , n3404 );
    nor g5139 ( n4457 , n4276 , n4064 );
    not g5140 ( n4821 , n4108 );
    or g5141 ( n2257 , n2480 , n2096 );
    not g5142 ( n1379 , n2288 );
    or g5143 ( n2060 , n442 , n1439 );
    not g5144 ( n5495 , n1227 );
    or g5145 ( n4655 , n3541 , n2717 );
    and g5146 ( n3968 , n2437 , n1721 );
    not g5147 ( n2923 , n3993 );
    not g5148 ( n6263 , n4532 );
    and g5149 ( n5129 , n2347 , n3466 );
    and g5150 ( n2827 , n445 , n4905 );
    nor g5151 ( n3292 , n5084 , n5776 );
    not g5152 ( n3837 , n5721 );
    not g5153 ( n145 , n4869 );
    nor g5154 ( n3427 , n6123 , n3988 );
    or g5155 ( n3812 , n4157 , n6009 );
    nor g5156 ( n2119 , n5280 , n5787 );
    or g5157 ( n5853 , n1346 , n2480 );
    and g5158 ( n2579 , n4156 , n4208 );
    or g5159 ( n5658 , n4150 , n4167 );
    not g5160 ( n3028 , n23 );
    not g5161 ( n4317 , n2720 );
    not g5162 ( n1215 , n2250 );
    not g5163 ( n6183 , n3969 );
    nor g5164 ( n2405 , n1422 , n2776 );
    or g5165 ( n5743 , n3129 , n2784 );
    not g5166 ( n2057 , n2219 );
    nor g5167 ( n4082 , n5426 , n5412 );
    and g5168 ( n2251 , n1411 , n3888 );
    nor g5169 ( n3620 , n2709 , n1128 );
    not g5170 ( n2938 , n4339 );
    not g5171 ( n2409 , n3012 );
    and g5172 ( n4096 , n478 , n4479 );
    not g5173 ( n2780 , n1104 );
    not g5174 ( n2444 , n2417 );
    nor g5175 ( n2272 , n5165 , n2322 );
    or g5176 ( n2466 , n3589 , n4402 );
    not g5177 ( n4648 , n495 );
    nor g5178 ( n2041 , n5890 , n5320 );
    or g5179 ( n4764 , n588 , n2622 );
    or g5180 ( n255 , n2931 , n2399 );
    and g5181 ( n3100 , n5565 , n4885 );
    and g5182 ( n3605 , n5549 , n1673 );
    nor g5183 ( n252 , n143 , n3508 );
    or g5184 ( n4594 , n1155 , n5924 );
    not g5185 ( n4970 , n777 );
    not g5186 ( n310 , n5524 );
    not g5187 ( n6145 , n5485 );
    and g5188 ( n2834 , n4144 , n5260 );
    not g5189 ( n2106 , n5115 );
    and g5190 ( n4951 , n1300 , n4526 );
    nor g5191 ( n6074 , n548 , n2673 );
    or g5192 ( n3216 , n318 , n1587 );
    not g5193 ( n810 , n3962 );
    not g5194 ( n2899 , n6175 );
    not g5195 ( n5568 , n1786 );
    and g5196 ( n532 , n352 , n2130 );
    nor g5197 ( n3388 , n93 , n1465 );
    and g5198 ( n2849 , n496 , n2150 );
    nor g5199 ( n4681 , n5593 , n927 );
    and g5200 ( n4849 , n5048 , n4352 );
    and g5201 ( n975 , n4852 , n3632 );
    not g5202 ( n4984 , n5314 );
    or g5203 ( n3741 , n5497 , n3623 );
    or g5204 ( n5156 , n776 , n1373 );
    or g5205 ( n611 , n4028 , n3551 );
    and g5206 ( n951 , n1457 , n5850 );
    not g5207 ( n4166 , n4952 );
    nor g5208 ( n2292 , n3230 , n164 );
    not g5209 ( n2342 , n565 );
    or g5210 ( n2864 , n1746 , n1480 );
    or g5211 ( n557 , n1893 , n1867 );
    not g5212 ( n693 , n5104 );
    not g5213 ( n1105 , n2090 );
    or g5214 ( n6142 , n1607 , n5015 );
    not g5215 ( n2513 , n1931 );
    not g5216 ( n184 , n1946 );
    nor g5217 ( n5922 , n1626 , n5352 );
    or g5218 ( n4957 , n5848 , n4467 );
    and g5219 ( n4703 , n335 , n2017 );
    nor g5220 ( n5469 , n1570 , n5885 );
    or g5221 ( n1686 , n3064 , n3386 );
    and g5222 ( n1446 , n2307 , n3502 );
    and g5223 ( n3907 , n6116 , n1787 );
    or g5224 ( n4200 , n1741 , n2696 );
    not g5225 ( n3777 , n2273 );
    or g5226 ( n5799 , n704 , n3792 );
    and g5227 ( n3051 , n5181 , n4835 );
    nor g5228 ( n5826 , n4245 , n3253 );
    or g5229 ( n3475 , n5372 , n3612 );
    nor g5230 ( n466 , n2676 , n729 );
    and g5231 ( n1964 , n2224 , n3955 );
    nor g5232 ( n1936 , n4231 , n1046 );
    not g5233 ( n5074 , n3993 );
    not g5234 ( n3677 , n3484 );
    nor g5235 ( n1784 , n285 , n2911 );
    or g5236 ( n5463 , n4273 , n630 );
    or g5237 ( n3465 , n5523 , n4967 );
    not g5238 ( n3999 , n4281 );
    and g5239 ( n6105 , n3362 , n1997 );
    and g5240 ( n2104 , n4931 , n2994 );
    not g5241 ( n919 , n2638 );
    or g5242 ( n553 , n2834 , n4546 );
    nor g5243 ( n2380 , n5316 , n4417 );
    nor g5244 ( n4662 , n696 , n3992 );
    not g5245 ( n6004 , n1945 );
    or g5246 ( n4834 , n2610 , n1583 );
    and g5247 ( n4727 , n3473 , n3242 );
    not g5248 ( n4286 , n4312 );
    not g5249 ( n2608 , n507 );
    nor g5250 ( n3377 , n5376 , n6013 );
    not g5251 ( n4456 , n5602 );
    not g5252 ( n2365 , n1008 );
    and g5253 ( n649 , n2858 , n5193 );
    and g5254 ( n2961 , n602 , n4353 );
    and g5255 ( n914 , n5244 , n5950 );
    nor g5256 ( n2201 , n2289 , n800 );
    or g5257 ( n1208 , n2007 , n4017 );
    and g5258 ( n1057 , n1309 , n1788 );
    or g5259 ( n5250 , n2595 , n545 );
    or g5260 ( n3062 , n1099 , n4038 );
    and g5261 ( n3996 , n4317 , n3227 );
    or g5262 ( n3090 , n3940 , n5289 );
    and g5263 ( n4269 , n1069 , n206 );
    not g5264 ( n6214 , n3053 );
    not g5265 ( n5385 , n747 );
    not g5266 ( n4007 , n20 );
    and g5267 ( n241 , n4574 , n5385 );
    or g5268 ( n5194 , n5718 , n1210 );
    or g5269 ( n1793 , n2956 , n5319 );
    not g5270 ( n1571 , n1109 );
    or g5271 ( n1970 , n1764 , n888 );
    not g5272 ( n3799 , n1834 );
    or g5273 ( n2499 , n255 , n3806 );
    and g5274 ( n3185 , n4000 , n4710 );
    nor g5275 ( n34 , n4288 , n2209 );
    or g5276 ( n3253 , n104 , n5494 );
    or g5277 ( n3956 , n3221 , n928 );
    nor g5278 ( n5057 , n5903 , n3287 );
    or g5279 ( n1953 , n4172 , n4429 );
    nor g5280 ( n6126 , n381 , n4121 );
    nor g5281 ( n2906 , n3011 , n2312 );
    not g5282 ( n4444 , n1032 );
    or g5283 ( n5405 , n813 , n615 );
    not g5284 ( n6149 , n6197 );
    and g5285 ( n1200 , n3259 , n4246 );
    or g5286 ( n5453 , n2468 , n5406 );
    not g5287 ( n4073 , n5417 );
    not g5288 ( n909 , n2763 );
    not g5289 ( n5137 , n2695 );
    not g5290 ( n1550 , n2948 );
    not g5291 ( n1231 , n183 );
    or g5292 ( n2989 , n69 , n5971 );
    or g5293 ( n4037 , n3028 , n2624 );
    nor g5294 ( n5152 , n5252 , n5519 );
    and g5295 ( n4999 , n5607 , n1307 );
    and g5296 ( n3625 , n4258 , n1478 );
    or g5297 ( n4476 , n3635 , n3682 );
    not g5298 ( n111 , n5599 );
    nor g5299 ( n50 , n5919 , n5109 );
    not g5300 ( n2140 , n386 );
    or g5301 ( n4819 , n3265 , n3145 );
    nor g5302 ( n2359 , n2746 , n5146 );
    and g5303 ( n2963 , n6127 , n4562 );
    and g5304 ( n2777 , n1928 , n5697 );
    and g5305 ( n1667 , n6072 , n1630 );
    or g5306 ( n2789 , n2267 , n5695 );
    and g5307 ( n4910 , n3132 , n2200 );
    nor g5308 ( n3340 , n1621 , n4247 );
    and g5309 ( n1278 , n611 , n1608 );
    or g5310 ( n1814 , n2360 , n3418 );
    or g5311 ( n5214 , n568 , n2620 );
    and g5312 ( n5432 , n3241 , n3305 );
    or g5313 ( n4729 , n5043 , n3377 );
    or g5314 ( n5404 , n2570 , n876 );
    not g5315 ( n4197 , n3813 );
    or g5316 ( n1995 , n1781 , n949 );
    or g5317 ( n827 , n5157 , n640 );
    not g5318 ( n1525 , n3053 );
    or g5319 ( n1380 , n5475 , n3600 );
    nor g5320 ( n680 , n2182 , n5922 );
    or g5321 ( n574 , n6032 , n380 );
    or g5322 ( n4739 , n3204 , n1742 );
    or g5323 ( n1916 , n1935 , n4255 );
    not g5324 ( n2573 , n4310 );
    or g5325 ( n420 , n5292 , n264 );
    nor g5326 ( n2357 , n909 , n3957 );
    or g5327 ( n3424 , n1866 , n1647 );
    or g5328 ( n4580 , n854 , n4548 );
    not g5329 ( n105 , n522 );
    or g5330 ( n267 , n414 , n6014 );
    not g5331 ( n3818 , n5450 );
    or g5332 ( n1524 , n1536 , n4499 );
    not g5333 ( n3607 , n41 );
    or g5334 ( n3659 , n2583 , n6153 );
    not g5335 ( n4522 , n4263 );
    not g5336 ( n1631 , n2446 );
    or g5337 ( n4075 , n6 , n6265 );
    or g5338 ( n121 , n2692 , n1733 );
    or g5339 ( n2659 , n1393 , n1661 );
    and g5340 ( n4351 , n6105 , n854 );
    and g5341 ( n47 , n3517 , n4602 );
    or g5342 ( n4992 , n4049 , n837 );
    not g5343 ( n1795 , n6253 );
    or g5344 ( n1206 , n3765 , n1322 );
    nor g5345 ( n5924 , n5824 , n3668 );
    or g5346 ( n5310 , n4319 , n1729 );
    or g5347 ( n6204 , n2203 , n1077 );
    not g5348 ( n889 , n3334 );
    not g5349 ( n2871 , n5678 );
    nor g5350 ( n5034 , n3123 , n166 );
    and g5351 ( n3953 , n3449 , n6048 );
    and g5352 ( n4140 , n6245 , n3453 );
    nor g5353 ( n6230 , n5277 , n779 );
    nor g5354 ( n4902 , n736 , n4006 );
    or g5355 ( n28 , n3630 , n1710 );
    nor g5356 ( n1698 , n2845 , n1717 );
    or g5357 ( n4549 , n4939 , n3639 );
    not g5358 ( n1401 , n3205 );
    not g5359 ( n2311 , n582 );
    nor g5360 ( n2268 , n2282 , n5432 );
    nor g5361 ( n5933 , n2958 , n3234 );
    not g5362 ( n5969 , n419 );
    and g5363 ( n2423 , n6027 , n3089 );
    not g5364 ( n2799 , n2311 );
    and g5365 ( n410 , n634 , n1290 );
    not g5366 ( n5000 , n1297 );
    not g5367 ( n3776 , n2655 );
    or g5368 ( n5098 , n52 , n2066 );
    not g5369 ( n1601 , n6247 );
    not g5370 ( n6118 , n4957 );
    or g5371 ( n5769 , n374 , n5029 );
    nor g5372 ( n3295 , n2091 , n6043 );
    and g5373 ( n5691 , n3041 , n1144 );
    not g5374 ( n3398 , n5090 );
    not g5375 ( n5131 , n3715 );
    and g5376 ( n929 , n3036 , n789 );
    not g5377 ( n1154 , n2436 );
    and g5378 ( n990 , n5449 , n4106 );
    and g5379 ( n6252 , n1812 , n5646 );
    not g5380 ( n1316 , n3535 );
    not g5381 ( n3074 , n4488 );
    not g5382 ( n5362 , n2157 );
    or g5383 ( n2415 , n401 , n2375 );
    nor g5384 ( n6268 , n114 , n4174 );
    not g5385 ( n5779 , n621 );
    and g5386 ( n4301 , n502 , n1548 );
    and g5387 ( n201 , n3521 , n3190 );
    not g5388 ( n5114 , n4714 );
    nor g5389 ( n2313 , n6268 , n911 );
    or g5390 ( n4199 , n1171 , n5841 );
    or g5391 ( n4032 , n731 , n4325 );
    nor g5392 ( n743 , n4162 , n842 );
    not g5393 ( n2412 , n4589 );
    or g5394 ( n2250 , n4886 , n5430 );
    or g5395 ( n4079 , n6054 , n932 );
    or g5396 ( n5056 , n535 , n2571 );
    nor g5397 ( n4647 , n639 , n6240 );
    not g5398 ( n3307 , n1680 );
    and g5399 ( n2810 , n1574 , n3718 );
    or g5400 ( n4280 , n1964 , n3247 );
    or g5401 ( n5834 , n5480 , n5347 );
    or g5402 ( n2684 , n5932 , n3153 );
    or g5403 ( n5222 , n1354 , n4129 );
    or g5404 ( n5788 , n280 , n5297 );
    and g5405 ( n1075 , n3870 , n2674 );
    not g5406 ( n2308 , n2929 );
    or g5407 ( n4980 , n2331 , n43 );
    and g5408 ( n1424 , n896 , n5884 );
    not g5409 ( n2934 , n1895 );
    or g5410 ( n851 , n4451 , n974 );
    or g5411 ( n5225 , n804 , n5383 );
    and g5412 ( n1474 , n5574 , n4636 );
    and g5413 ( n2162 , n5723 , n4911 );
    or g5414 ( n5962 , n1910 , n190 );
    not g5415 ( n5795 , n1802 );
    or g5416 ( n1902 , n2679 , n2687 );
    not g5417 ( n4772 , n1201 );
    or g5418 ( n1440 , n877 , n5570 );
    not g5419 ( n2586 , n4119 );
    not g5420 ( n934 , n4072 );
    not g5421 ( n1349 , n3414 );
    not g5422 ( n1831 , n5233 );
    and g5423 ( n3392 , n5693 , n6058 );
    or g5424 ( n2095 , n2914 , n6257 );
    nor g5425 ( n2887 , n4045 , n4857 );
    nor g5426 ( n5296 , n1903 , n556 );
    and g5427 ( n1915 , n6276 , n5064 );
    not g5428 ( n4452 , n638 );
    nor g5429 ( n3938 , n1776 , n3736 );
    not g5430 ( n5282 , n2714 );
    not g5431 ( n5918 , n1631 );
    or g5432 ( n3835 , n1 , n4139 );
    and g5433 ( n4693 , n3165 , n2722 );
    or g5434 ( n2837 , n4213 , n2718 );
    nor g5435 ( n73 , n755 , n3512 );
    or g5436 ( n3162 , n4670 , n2319 );
    or g5437 ( n767 , n2859 , n514 );
    not g5438 ( n3050 , n4396 );
    or g5439 ( n4941 , n5914 , n135 );
    not g5440 ( n3143 , n2408 );
    or g5441 ( n5889 , n3160 , n6182 );
    or g5442 ( n164 , n1927 , n5302 );
    not g5443 ( n4004 , n365 );
    not g5444 ( n5325 , n1762 );
    not g5445 ( n3850 , n1246 );
    and g5446 ( n3429 , n4219 , n730 );
    or g5447 ( n3641 , n1673 , n208 );
    or g5448 ( n2511 , n5064 , n1819 );
    and g5449 ( n763 , n4207 , n146 );
    not g5450 ( n6021 , n407 );
    not g5451 ( n6137 , n4379 );
    nor g5452 ( n5847 , n5386 , n3700 );
    or g5453 ( n485 , n1565 , n5561 );
    and g5454 ( n1488 , n5982 , n1438 );
    and g5455 ( n1993 , n5002 , n972 );
    not g5456 ( n854 , n5510 );
    and g5457 ( n4194 , n167 , n5196 );
    not g5458 ( n4150 , n5356 );
    nor g5459 ( n2479 , n5687 , n4958 );
    nor g5460 ( n4946 , n5832 , n1740 );
    nor g5461 ( n857 , n2841 , n3939 );
    and g5462 ( n5603 , n4244 , n3685 );
    or g5463 ( n3247 , n2426 , n354 );
    not g5464 ( n2055 , n2199 );
    not g5465 ( n2994 , n747 );
    not g5466 ( n1657 , n2752 );
    or g5467 ( n4463 , n836 , n4877 );
    or g5468 ( n4017 , n4416 , n6258 );
    not g5469 ( n4541 , n4167 );
    or g5470 ( n5175 , n1937 , n1226 );
    or g5471 ( n2927 , n3955 , n5148 );
    or g5472 ( n3977 , n4704 , n4628 );
    and g5473 ( n6195 , n1702 , n4827 );
    not g5474 ( n1529 , n4727 );
    nor g5475 ( n4797 , n3402 , n5967 );
    nor g5476 ( n3979 , n5445 , n5125 );
    not g5477 ( n5625 , n4170 );
    not g5478 ( n1605 , n4305 );
    or g5479 ( n5905 , n4691 , n2932 );
    nor g5480 ( n4438 , n4847 , n3853 );
    not g5481 ( n4536 , n4733 );
    not g5482 ( n5640 , n3651 );
    or g5483 ( n3405 , n4777 , n6190 );
    or g5484 ( n3638 , n5785 , n4999 );
    not g5485 ( n3881 , n2104 );
    or g5486 ( n5749 , n4332 , n3692 );
    nor g5487 ( n2680 , n4604 , n6027 );
    and g5488 ( n729 , n4666 , n3579 );
    nor g5489 ( n5410 , n3146 , n991 );
    and g5490 ( n599 , n5550 , n394 );
    and g5491 ( n998 , n4062 , n4919 );
    or g5492 ( n5042 , n5685 , n2061 );
    not g5493 ( n5238 , n2175 );
    not g5494 ( n2387 , n192 );
    or g5495 ( n5251 , n4637 , n4264 );
    nor g5496 ( n1718 , n2463 , n4080 );
    nor g5497 ( n6124 , n2047 , n5660 );
    and g5498 ( n1704 , n386 , n5215 );
    nor g5499 ( n3833 , n1122 , n3291 );
    or g5500 ( n5399 , n4381 , n1659 );
    or g5501 ( n2616 , n4426 , n3169 );
    or g5502 ( n3417 , n3332 , n3975 );
    and g5503 ( n3298 , n1241 , n3756 );
    or g5504 ( n2913 , n5469 , n1827 );
    or g5505 ( n2708 , n3106 , n4103 );
    nor g5506 ( n4112 , n3299 , n246 );
    or g5507 ( n4084 , n1316 , n4730 );
    or g5508 ( n4762 , n1703 , n3725 );
    and g5509 ( n1387 , n4126 , n2104 );
    nor g5510 ( n4489 , n2851 , n2866 );
    not g5511 ( n2039 , n4441 );
    nor g5512 ( n5942 , n5662 , n2037 );
    or g5513 ( n5068 , n5218 , n5350 );
    or g5514 ( n1610 , n3832 , n6188 );
    and g5515 ( n3209 , n6285 , n2431 );
    nor g5516 ( n1944 , n4365 , n5803 );
    or g5517 ( n4072 , n4680 , n4250 );
    or g5518 ( n1043 , n6147 , n3361 );
    nor g5519 ( n434 , n6161 , n6085 );
    not g5520 ( n6120 , n694 );
    and g5521 ( n5107 , n3350 , n4592 );
    not g5522 ( n5484 , n4352 );
    or g5523 ( n2446 , n6086 , n2561 );
    not g5524 ( n5020 , n980 );
    nor g5525 ( n3311 , n3464 , n458 );
    or g5526 ( n3471 , n1001 , n779 );
    not g5527 ( n2385 , n4043 );
    and g5528 ( n339 , n2555 , n5460 );
    or g5529 ( n2861 , n4597 , n5661 );
    nor g5530 ( n5726 , n3037 , n6054 );
    not g5531 ( n5953 , n5309 );
    not g5532 ( n5249 , n6004 );
    not g5533 ( n2703 , n2416 );
    not g5534 ( n3512 , n6017 );
    nor g5535 ( n245 , n5177 , n2069 );
    not g5536 ( n231 , n6088 );
    nor g5537 ( n5507 , n360 , n2029 );
    or g5538 ( n1798 , n5508 , n5803 );
    not g5539 ( n2800 , n2191 );
    or g5540 ( n3594 , n168 , n5077 );
    not g5541 ( n1637 , n5557 );
    and g5542 ( n2316 , n3122 , n1633 );
    not g5543 ( n5418 , n4744 );
    not g5544 ( n2582 , n3764 );
    not g5545 ( n4441 , n4828 );
    or g5546 ( n365 , n1918 , n4026 );
    nor g5547 ( n3257 , n3087 , n1363 );
    not g5548 ( n5808 , n5601 );
    nor g5549 ( n3251 , n5128 , n6151 );
    or g5550 ( n5294 , n1829 , n2816 );
    or g5551 ( n5518 , n2036 , n4841 );
    and g5552 ( n1769 , n3712 , n3882 );
    nor g5553 ( n816 , n5344 , n3648 );
    and g5554 ( n2321 , n2827 , n384 );
    not g5555 ( n428 , n2783 );
    and g5556 ( n3954 , n3567 , n4984 );
    and g5557 ( n1979 , n3274 , n2052 );
    not g5558 ( n4738 , n2055 );
    nor g5559 ( n4632 , n873 , n435 );
    or g5560 ( n3481 , n1136 , n2328 );
    not g5561 ( n4372 , n650 );
    or g5562 ( n1930 , n4525 , n1805 );
    or g5563 ( n459 , n687 , n1432 );
    not g5564 ( n3749 , n6269 );
    not g5565 ( n2103 , n1443 );
    or g5566 ( n3653 , n812 , n5328 );
    and g5567 ( n1612 , n4876 , n5022 );
    and g5568 ( n5986 , n1057 , n1679 );
    or g5569 ( n3228 , n4773 , n5887 );
    nor g5570 ( n4154 , n2198 , n2342 );
    and g5571 ( n3991 , n2431 , n6128 );
    and g5572 ( n1192 , n1498 , n1108 );
    and g5573 ( n5122 , n1336 , n1048 );
    not g5574 ( n2253 , n5498 );
    not g5575 ( n4170 , n1462 );
    not g5576 ( n1247 , n4270 );
    not g5577 ( n3269 , n711 );
    not g5578 ( n5339 , n4720 );
    not g5579 ( n3402 , n483 );
    and g5580 ( n1809 , n4314 , n1036 );
    and g5581 ( n5224 , n968 , n3458 );
    or g5582 ( n4310 , n4119 , n6290 );
    not g5583 ( n3262 , n2885 );
    and g5584 ( n144 , n2255 , n1831 );
    or g5585 ( n666 , n290 , n5270 );
    nor g5586 ( n3029 , n4389 , n2134 );
    not g5587 ( n333 , n2741 );
    not g5588 ( n2036 , n1019 );
    nor g5589 ( n5474 , n3935 , n2288 );
    not g5590 ( n4794 , n779 );
    and g5591 ( n3226 , n2573 , n4083 );
    and g5592 ( n3 , n5400 , n1388 );
    nor g5593 ( n1766 , n25 , n133 );
    not g5594 ( n5802 , n1218 );
    not g5595 ( n2712 , n3840 );
    not g5596 ( n4507 , n865 );
    and g5597 ( n1300 , n3453 , n3895 );
    nor g5598 ( n1891 , n2577 , n5521 );
    not g5599 ( n2730 , n4898 );
    nor g5600 ( n5187 , n4257 , n5229 );
    not g5601 ( n2984 , n2005 );
    or g5602 ( n3009 , n4882 , n3801 );
    not g5603 ( n515 , n22 );
    not g5604 ( n4608 , n1951 );
    nor g5605 ( n2589 , n3437 , n4394 );
    or g5606 ( n5063 , n4889 , n4065 );
    nor g5607 ( n3139 , n388 , n4225 );
    not g5608 ( n1195 , n1807 );
    or g5609 ( n6190 , n4188 , n3504 );
    not g5610 ( n2291 , n3912 );
    not g5611 ( n2030 , n2546 );
    or g5612 ( n3222 , n4043 , n6017 );
    not g5613 ( n1607 , n6200 );
    nor g5614 ( n226 , n6302 , n2025 );
    not g5615 ( n5730 , n4245 );
    or g5616 ( n789 , n2956 , n2706 );
    or g5617 ( n4748 , n2864 , n4420 );
    and g5618 ( n5052 , n5089 , n65 );
    and g5619 ( n3323 , n2504 , n3968 );
    nor g5620 ( n5569 , n64 , n4389 );
    nor g5621 ( n1139 , n3184 , n1901 );
    nor g5622 ( n2881 , n2141 , n725 );
    not g5623 ( n1328 , n2961 );
    or g5624 ( n5963 , n3799 , n1160 );
    not g5625 ( n2566 , n2245 );
    nor g5626 ( n1991 , n2595 , n5608 );
    nor g5627 ( n5245 , n5273 , n3085 );
    and g5628 ( n2848 , n798 , n3776 );
    nor g5629 ( n5434 , n4845 , n2472 );
    or g5630 ( n833 , n924 , n5384 );
    not g5631 ( n4439 , n850 );
    nor g5632 ( n291 , n5220 , n6081 );
    not g5633 ( n6032 , n4413 );
    not g5634 ( n2845 , n1451 );
    not g5635 ( n3071 , n1588 );
    or g5636 ( n5529 , n874 , n450 );
    not g5637 ( n1054 , n1270 );
    not g5638 ( n360 , n3583 );
    not g5639 ( n2098 , n4995 );
    or g5640 ( n1242 , n5403 , n5771 );
    or g5641 ( n3711 , n6122 , n1492 );
    not g5642 ( n868 , n2542 );
    or g5643 ( n5456 , n6018 , n5405 );
    nor g5644 ( n2006 , n5314 , n3826 );
    and g5645 ( n4086 , n3771 , n5625 );
    and g5646 ( n2151 , n4968 , n1336 );
    nor g5647 ( n5192 , n4886 , n990 );
    or g5648 ( n2185 , n3395 , n1408 );
    not g5649 ( n1415 , n4555 );
    not g5650 ( n5460 , n3684 );
    not g5651 ( n6168 , n5860 );
    or g5652 ( n3774 , n6193 , n902 );
    nor g5653 ( n1811 , n2440 , n6282 );
    nor g5654 ( n6194 , n4432 , n3372 );
    not g5655 ( n4270 , n347 );
    not g5656 ( n4789 , n4142 );
    or g5657 ( n5283 , n1669 , n478 );
    or g5658 ( n2550 , n1786 , n2180 );
    not g5659 ( n3447 , n2695 );
    not g5660 ( n4311 , n5636 );
    or g5661 ( n1185 , n6169 , n2187 );
    or g5662 ( n4018 , n2761 , n3373 );
    not g5663 ( n5977 , n5425 );
    or g5664 ( n1296 , n5237 , n4367 );
    and g5665 ( n5230 , n5656 , n3482 );
    not g5666 ( n638 , n695 );
    not g5667 ( n416 , n5523 );
    not g5668 ( n2758 , n3830 );
    or g5669 ( n3915 , n2367 , n2606 );
    not g5670 ( n573 , n1942 );
    or g5671 ( n1187 , n2065 , n511 );
    and g5672 ( n717 , n516 , n5226 );
    or g5673 ( n5367 , n2885 , n1950 );
    and g5674 ( n605 , n3256 , n3110 );
    and g5675 ( n5699 , n5393 , n1019 );
    or g5676 ( n4652 , n2458 , n5941 );
    not g5677 ( n591 , n2643 );
    not g5678 ( n5680 , n5907 );
    not g5679 ( n5231 , n1799 );
    nor g5680 ( n3197 , n692 , n4964 );
    or g5681 ( n5968 , n2043 , n4189 );
    or g5682 ( n5694 , n355 , n5646 );
    and g5683 ( n1500 , n5310 , n3689 );
    nor g5684 ( n4455 , n2599 , n737 );
    or g5685 ( n5684 , n6264 , n3108 );
    and g5686 ( n4688 , n1758 , n6143 );
    or g5687 ( n2819 , n1730 , n3267 );
    nor g5688 ( n1801 , n2874 , n1866 );
    nor g5689 ( n2080 , n1194 , n2880 );
    or g5690 ( n4629 , n715 , n3172 );
    and g5691 ( n711 , n5491 , n4259 );
    or g5692 ( n2687 , n1949 , n3393 );
    not g5693 ( n6272 , n2733 );
    or g5694 ( n3706 , n2250 , n1466 );
    and g5695 ( n3157 , n1743 , n402 );
    or g5696 ( n1923 , n1314 , n6021 );
    not g5697 ( n4928 , n165 );
    and g5698 ( n2885 , n6171 , n3499 );
    nor g5699 ( n6083 , n4671 , n852 );
    nor g5700 ( n3981 , n1352 , n5989 );
    and g5701 ( n1079 , n2698 , n30 );
    or g5702 ( n3729 , n3218 , n5119 );
    or g5703 ( n2567 , n3990 , n4725 );
    or g5704 ( n1093 , n2918 , n3285 );
    and g5705 ( n5772 , n4409 , n4256 );
    nor g5706 ( n4765 , n6159 , n5055 );
    or g5707 ( n504 , n1622 , n1384 );
    or g5708 ( n1405 , n4073 , n219 );
    not g5709 ( n5276 , n3411 );
    or g5710 ( n1973 , n5003 , n2353 );
    or g5711 ( n2187 , n4780 , n575 );
    or g5712 ( n1499 , n3981 , n4862 );
    or g5713 ( n4488 , n3731 , n3835 );
    nor g5714 ( n860 , n3133 , n797 );
    nor g5715 ( n2198 , n3171 , n5775 );
    nor g5716 ( n6026 , n1048 , n109 );
    nor g5717 ( n2910 , n5180 , n3530 );
    not g5718 ( n3181 , n639 );
    or g5719 ( n5774 , n1785 , n1639 );
    not g5720 ( n2327 , n2841 );
    not g5721 ( n1871 , n4820 );
    and g5722 ( n3539 , n1837 , n3777 );
    or g5723 ( n204 , n6219 , n6270 );
    nor g5724 ( n6237 , n3621 , n3398 );
    not g5725 ( n6087 , n1791 );
    nor g5726 ( n907 , n1807 , n27 );
    or g5727 ( n3657 , n6035 , n5650 );
    not g5728 ( n2063 , n3677 );
    or g5729 ( n4137 , n5258 , n5353 );
    not g5730 ( n3117 , n5310 );
    or g5731 ( n1543 , n3866 , n2979 );
    not g5732 ( n270 , n4256 );
    nor g5733 ( n1828 , n1972 , n1412 );
    nor g5734 ( n3663 , n1576 , n3478 );
    and g5735 ( n438 , n1510 , n5545 );
    not g5736 ( n1257 , n4651 );
    or g5737 ( n2073 , n1878 , n409 );
    and g5738 ( n1383 , n1484 , n5717 );
    not g5739 ( n80 , n4037 );
    and g5740 ( n1484 , n1648 , n94 );
    not g5741 ( n5466 , n594 );
    and g5742 ( n5269 , n3471 , n3129 );
    not g5743 ( n2569 , n938 );
    nor g5744 ( n5840 , n1806 , n4387 );
    and g5745 ( n3853 , n5851 , n4439 );
    and g5746 ( n2949 , n3533 , n4504 );
    nor g5747 ( n1555 , n1443 , n4043 );
    and g5748 ( n2414 , n1540 , n4675 );
    and g5749 ( n6130 , n4486 , n4075 );
    or g5750 ( n407 , n3993 , n3053 );
    not g5751 ( n4586 , n3583 );
    or g5752 ( n6135 , n6300 , n1250 );
    or g5753 ( n5443 , n785 , n3413 );
    or g5754 ( n661 , n3691 , n282 );
    or g5755 ( n3040 , n2625 , n6079 );
    not g5756 ( n2655 , n3640 );
    not g5757 ( n2194 , n3362 );
    not g5758 ( n383 , n490 );
    not g5759 ( n3871 , n1066 );
    not g5760 ( n260 , n6096 );
    nor g5761 ( n2350 , n3457 , n5046 );
    not g5762 ( n5413 , n91 );
    and g5763 ( n2484 , n4211 , n4266 );
    or g5764 ( n4945 , n1000 , n5917 );
    nor g5765 ( n5894 , n3845 , n1983 );
    and g5766 ( n3064 , n6101 , n1526 );
    nor g5767 ( n493 , n6106 , n3986 );
    nor g5768 ( n5615 , n1363 , n5667 );
    not g5769 ( n3255 , n5534 );
    nor g5770 ( n5318 , n2004 , n2123 );
    not g5771 ( n5351 , n6109 );
    nor g5772 ( n4646 , n906 , n291 );
    nor g5773 ( n2164 , n1777 , n5320 );
    and g5774 ( n5082 , n1756 , n5037 );
    nor g5775 ( n2197 , n768 , n1956 );
    nor g5776 ( n5024 , n4279 , n2338 );
    and g5777 ( n3042 , n5443 , n1680 );
    or g5778 ( n6153 , n2092 , n2911 );
    nor g5779 ( n3370 , n5233 , n3485 );
    or g5780 ( n5896 , n76 , n1679 );
    not g5781 ( n388 , n3959 );
    not g5782 ( n1457 , n4607 );
    or g5783 ( n2932 , n2454 , n5182 );
    or g5784 ( n1534 , n1689 , n6251 );
    or g5785 ( n2358 , n869 , n1880 );
    nor g5786 ( n5210 , n1098 , n5609 );
    and g5787 ( n4565 , n990 , n1581 );
    or g5788 ( n4836 , n3931 , n2339 );
    not g5789 ( n1707 , n2112 );
    or g5790 ( n5113 , n2954 , n3966 );
    not g5791 ( n6208 , n2675 );
    not g5792 ( n3230 , n3101 );
    or g5793 ( n678 , n5414 , n6078 );
    and g5794 ( n2108 , n1030 , n593 );
    not g5795 ( n6068 , n1988 );
    buf g5796 ( n2360 , n913 );
    or g5797 ( n1772 , n2207 , n1892 );
    not g5798 ( n2790 , n2451 );
    and g5799 ( n1082 , n379 , n4552 );
    not g5800 ( n6048 , n3881 );
    or g5801 ( n5675 , n5482 , n4834 );
    or g5802 ( n1177 , n3803 , n3398 );
    or g5803 ( n1392 , n3548 , n1233 );
    nor g5804 ( n761 , n2028 , n1847 );
    or g5805 ( n533 , n2205 , n5345 );
    nor g5806 ( n1020 , n257 , n4912 );
    or g5807 ( n2862 , n5886 , n1833 );
    nor g5808 ( n4478 , n3889 , n2613 );
    not g5809 ( n3484 , n4504 );
    nor g5810 ( n6216 , n931 , n6265 );
    and g5811 ( n758 , n5281 , n5773 );
    or g5812 ( n115 , n3097 , n3277 );
    or g5813 ( n1877 , n5879 , n2801 );
    nor g5814 ( n2192 , n6155 , n5186 );
    not g5815 ( n3545 , n3532 );
    and g5816 ( n4697 , n2064 , n6214 );
    and g5817 ( n4930 , n5655 , n5120 );
    nor g5818 ( n2457 , n4370 , n6036 );
    not g5819 ( n3457 , n4110 );
    nor g5820 ( n659 , n4270 , n1040 );
    nor g5821 ( n2775 , n5330 , n2991 );
    or g5822 ( n4264 , n613 , n4489 );
    and g5823 ( n5135 , n3873 , n220 );
    or g5824 ( n5050 , n71 , n5130 );
    not g5825 ( n181 , n5181 );
    or g5826 ( n922 , n4716 , n995 );
    or g5827 ( n3517 , n6104 , n4173 );
    and g5828 ( n4481 , n2842 , n2750 );
    not g5829 ( n5353 , n4937 );
    not g5830 ( n2067 , n627 );
    and g5831 ( n1434 , n6225 , n2767 );
    or g5832 ( n3868 , n1642 , n2972 );
    or g5833 ( n5207 , n3215 , n5459 );
    not g5834 ( n1581 , n3489 );
    not g5835 ( n2700 , n899 );
    and g5836 ( n4923 , n1836 , n4995 );
    nor g5837 ( n3210 , n4371 , n5421 );
    nor g5838 ( n4535 , n5857 , n4695 );
    and g5839 ( n6114 , n536 , n4403 );
    not g5840 ( n5134 , n2719 );
    or g5841 ( n5860 , n4823 , n6175 );
    or g5842 ( n5389 , n5579 , n3344 );
    nor g5843 ( n6284 , n1538 , n5439 );
    or g5844 ( n3610 , n4535 , n4621 );
    and g5845 ( n5736 , n1926 , n3071 );
    or g5846 ( n456 , n3772 , n5066 );
    not g5847 ( n1665 , n4849 );
    not g5848 ( n2970 , n5113 );
    not g5849 ( n5780 , n2722 );
    and g5850 ( n2012 , n2239 , n3013 );
    not g5851 ( n5940 , n4319 );
    and g5852 ( n1282 , n6007 , n2391 );
    nor g5853 ( n2955 , n982 , n4650 );
    nor g5854 ( n396 , n3452 , n829 );
    not g5855 ( n5297 , n679 );
    and g5856 ( n1438 , n4818 , n5508 );
    or g5857 ( n725 , n11 , n3088 );
    not g5858 ( n1846 , n6086 );
    nor g5859 ( n4460 , n49 , n1073 );
    or g5860 ( n3423 , n5826 , n252 );
    not g5861 ( n1900 , n5704 );
    or g5862 ( n5473 , n5864 , n4400 );
    not g5863 ( n2050 , n2031 );
    not g5864 ( n3102 , n4697 );
    or g5865 ( n925 , n125 , n1567 );
    nor g5866 ( n3309 , n5652 , n2670 );
    not g5867 ( n4868 , n1453 );
    and g5868 ( n1213 , n4606 , n3966 );
    or g5869 ( n2750 , n1512 , n672 );
    or g5870 ( n646 , n5303 , n3886 );
    not g5871 ( n3596 , n1978 );
    or g5872 ( n100 , n987 , n1205 );
    and g5873 ( n5571 , n2263 , n6069 );
    or g5874 ( n4433 , n381 , n1301 );
    and g5875 ( n558 , n1815 , n6277 );
    and g5876 ( n4135 , n1225 , n5434 );
    not g5877 ( n992 , n5757 );
    not g5878 ( n2091 , n1144 );
    or g5879 ( n1453 , n152 , n2528 );
    or g5880 ( n3234 , n1920 , n3051 );
    nor g5881 ( n1835 , n5103 , n5240 );
    nor g5882 ( n5980 , n6106 , n58 );
    not g5883 ( n1290 , n1619 );
    and g5884 ( n189 , n3584 , n2112 );
    not g5885 ( n2270 , n2975 );
    or g5886 ( n774 , n5921 , n1609 );
    not g5887 ( n3033 , n1924 );
    or g5888 ( n2170 , n2955 , n5379 );
    nor g5889 ( n4097 , n1726 , n4899 );
    not g5890 ( n790 , n2826 );
    or g5891 ( n616 , n4231 , n5258 );
    or g5892 ( n2592 , n6081 , n2684 );
    not g5893 ( n3768 , n2640 );
    or g5894 ( n1855 , n506 , n1814 );
    not g5895 ( n205 , n908 );
    nor g5896 ( n5054 , n3140 , n6084 );
    and g5897 ( n4174 , n3144 , n3325 );
    not g5898 ( n1628 , n4439 );
    or g5899 ( n849 , n706 , n3928 );
    nor g5900 ( n1456 , n3084 , n1530 );
    and g5901 ( n2320 , n3834 , n4888 );
    nor g5902 ( n3686 , n4584 , n2618 );
    not g5903 ( n686 , n3167 );
    or g5904 ( n1685 , n2780 , n4036 );
    not g5905 ( n4113 , n2244 );
    or g5906 ( n5844 , n894 , n2387 );
    nor g5907 ( n2492 , n5389 , n2156 );
    nor g5908 ( n4294 , n2470 , n3230 );
    not g5909 ( n3705 , n4331 );
    not g5910 ( n4758 , n4998 );
    nor g5911 ( n1994 , n5293 , n207 );
    not g5912 ( n6082 , n160 );
    nor g5913 ( n215 , n5408 , n2962 );
    or g5914 ( n1978 , n2563 , n5720 );
    or g5915 ( n1982 , n522 , n4844 );
    not g5916 ( n462 , n1489 );
    and g5917 ( n4811 , n5073 , n4297 );
    nor g5918 ( n2952 , n349 , n4478 );
    not g5919 ( n1561 , n1760 );
    or g5920 ( n5038 , n5062 , n3863 );
    and g5921 ( n2580 , n676 , n4146 );
    not g5922 ( n1087 , n3073 );
    or g5923 ( n1518 , n2714 , n4050 );
    and g5924 ( n2903 , n3319 , n5316 );
    not g5925 ( n5663 , n1360 );
    not g5926 ( n6093 , n3953 );
    or g5927 ( n4795 , n660 , n4987 );
    or g5928 ( n409 , n5860 , n2879 );
    or g5929 ( n3163 , n3847 , n2936 );
    not g5930 ( n890 , n3699 );
    and g5931 ( n3980 , n5105 , n4838 );
    not g5932 ( n72 , n1016 );
    or g5933 ( n96 , n857 , n4765 );
    or g5934 ( n2797 , n454 , n1892 );
    and g5935 ( n3039 , n5349 , n4644 );
    nor g5936 ( n378 , n1518 , n3862 );
    or g5937 ( n4706 , n2144 , n5764 );
    or g5938 ( n5738 , n4414 , n1879 );
    nor g5939 ( n1447 , n3915 , n4650 );
    or g5940 ( n4035 , n6275 , n4696 );
    not g5941 ( n1376 , n3231 );
    and g5942 ( n4985 , n4063 , n5837 );
    or g5943 ( n437 , n2702 , n953 );
    and g5944 ( n6056 , n4306 , n4504 );
    and g5945 ( n1578 , n4586 , n2333 );
    or g5946 ( n6025 , n2586 , n839 );
    and g5947 ( n6290 , n1711 , n3365 );
    nor g5948 ( n5343 , n2446 , n4646 );
    nor g5949 ( n1441 , n2502 , n4948 );
    nor g5950 ( n3855 , n1909 , n2592 );
    or g5951 ( n4374 , n50 , n1132 );
    not g5952 ( n435 , n120 );
    or g5953 ( n4056 , n2025 , n1454 );
    and g5954 ( n1410 , n3777 , n1792 );
    or g5955 ( n5433 , n824 , n3186 );
    and g5956 ( n1416 , n914 , n6221 );
    or g5957 ( n4659 , n185 , n2760 );
    or g5958 ( n2302 , n5466 , n5968 );
    or g5959 ( n274 , n5053 , n2663 );
    or g5960 ( n3375 , n279 , n227 );
    or g5961 ( n1865 , n2057 , n270 );
    or g5962 ( n932 , n6139 , n3592 );
    and g5963 ( n3006 , n4648 , n1621 );
    or g5964 ( n4894 , n2436 , n2132 );
    nor g5965 ( n4938 , n2027 , n424 );
    or g5966 ( n3294 , n349 , n1557 );
    nor g5967 ( n2086 , n4125 , n4672 );
    nor g5968 ( n1274 , n2935 , n2208 );
    or g5969 ( n21 , n5147 , n2334 );
    nor g5970 ( n3425 , n861 , n2007 );
    and g5971 ( n5234 , n2660 , n4735 );
    or g5972 ( n5595 , n6242 , n667 );
    not g5973 ( n1636 , n6056 );
    or g5974 ( n6055 , n1578 , n2197 );
    or g5975 ( n5613 , n4049 , n5120 );
    or g5976 ( n5822 , n596 , n969 );
    not g5977 ( n4111 , n169 );
    and g5978 ( n5800 , n1979 , n3189 );
    nor g5979 ( n1014 , n6038 , n6194 );
    nor g5980 ( n1773 , n2122 , n1299 );
    nor g5981 ( n3714 , n4338 , n72 );
    and g5982 ( n5435 , n918 , n6228 );
    nor g5983 ( n2283 , n3438 , n3268 );
    not g5984 ( n6203 , n1988 );
    or g5985 ( n3125 , n1070 , n317 );
    not g5986 ( n6106 , n4176 );
    not g5987 ( n1586 , n4803 );
    and g5988 ( n2335 , n1425 , n4346 );
    or g5989 ( n4585 , n2136 , n2805 );
    not g5990 ( n5171 , n2239 );
    not g5991 ( n3235 , n4220 );
    or g5992 ( n2879 , n5495 , n5675 );
    not g5993 ( n4307 , n197 );
    not g5994 ( n4295 , n6184 );
    nor g5995 ( n13 , n5576 , n3608 );
    not g5996 ( n2807 , n3190 );
    not g5997 ( n4658 , n4351 );
    nor g5998 ( n4033 , n2836 , n479 );
    and g5999 ( n1311 , n5936 , n1425 );
    nor g6000 ( n4 , n3418 , n1159 );
    nor g6001 ( n3341 , n152 , n2884 );
    nor g6002 ( n1121 , n2480 , n3841 );
    and g6003 ( n4672 , n4985 , n4620 );
    or g6004 ( n1078 , n6158 , n883 );
    not g6005 ( n377 , n4725 );
    not g6006 ( n3967 , n25 );
    or g6007 ( n3642 , n1524 , n5023 );
    or g6008 ( n3676 , n1709 , n2407 );
    nor g6009 ( n5300 , n4097 , n3297 );
    nor g6010 ( n2084 , n3969 , n5628 );
    not g6011 ( n795 , n3411 );
    and g6012 ( n366 , n4295 , n1648 );
    or g6013 ( n5320 , n1199 , n5658 );
    not g6014 ( n742 , n4839 );
    nor g6015 ( n4459 , n6299 , n1826 );
    or g6016 ( n1947 , n413 , n5785 );
    not g6017 ( n1204 , n2674 );
    not g6018 ( n5023 , n5723 );
    or g6019 ( n2241 , n2318 , n954 );
    and g6020 ( n648 , n1873 , n5461 );
    and g6021 ( n6255 , n1060 , n1443 );
    nor g6022 ( n652 , n2969 , n1389 );
    not g6023 ( n3510 , n3524 );
    nor g6024 ( n5669 , n2599 , n4446 );
    or g6025 ( n2965 , n2913 , n2924 );
    nor g6026 ( n5165 , n1395 , n4289 );
    or g6027 ( n655 , n528 , n4350 );
    not g6028 ( n5873 , n3750 );
    not g6029 ( n5938 , n1501 );
    or g6030 ( n1222 , n4061 , n2847 );
    nor g6031 ( n4822 , n5920 , n1782 );
    or g6032 ( n2525 , n3581 , n5169 );
    or g6033 ( n876 , n5042 , n6049 );
    not g6034 ( n5280 , n3193 );
    or g6035 ( n5934 , n4755 , n2977 );
    not g6036 ( n1408 , n5549 );
    and g6037 ( n4411 , n1063 , n438 );
    or g6038 ( n6213 , n5709 , n5532 );
    or g6039 ( n1761 , n191 , n3149 );
    not g6040 ( n4435 , n2390 );
    and g6041 ( n5287 , n3741 , n192 );
    not g6042 ( n1211 , n4059 );
    or g6043 ( n2422 , n5794 , n6271 );
    not g6044 ( n2667 , n5234 );
    not g6045 ( n1981 , n4832 );
    and g6046 ( n1569 , n1321 , n2471 );
    or g6047 ( n3883 , n4432 , n2531 );
    not g6048 ( n1000 , n1462 );
    not g6049 ( n1104 , n780 );
    or g6050 ( n2118 , n4971 , n4428 );
    nor g6051 ( n3004 , n1586 , n1477 );
    nor g6052 ( n4141 , n6048 , n2458 );
    not g6053 ( n412 , n3921 );
    not g6054 ( n4434 , n1491 );
    and g6055 ( n2467 , n4803 , n509 );
    not g6056 ( n5133 , n3613 );
    not g6057 ( n129 , n3486 );
    not g6058 ( n1281 , n788 );
    not g6059 ( n5424 , n22 );
endmodule
