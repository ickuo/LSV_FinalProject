module top( n3 , n6 , n13 , n25 , n27 , n32 , n40 , n41 , n44 , 
n51 , n55 , n57 , n58 , n60 , n62 , n64 , n80 , n83 , n86 , 
n93 , n95 , n103 , n104 , n110 , n116 , n129 , n130 , n131 , n133 , 
n136 , n140 , n144 , n157 , n164 , n167 , n172 , n175 , n181 , n182 , 
n183 , n196 , n205 , n210 , n213 , n216 , n225 , n229 , n234 , n236 , 
n257 , n260 , n266 , n272 , n274 , n275 , n276 , n281 , n286 , n289 , 
n293 , n297 , n299 , n315 , n318 , n325 , n332 , n334 , n340 , n344 , 
n357 , n362 , n365 , n375 , n397 , n402 , n404 , n406 , n414 , n418 , 
n427 , n432 , n433 , n434 , n439 , n441 , n442 , n445 , n447 , n450 , 
n455 , n463 , n466 , n470 , n471 , n476 , n484 , n488 , n490 , n492 , 
n494 , n502 , n509 , n511 , n512 , n520 , n521 );
    input n25 , n27 , n40 , n41 , n60 , n80 , n93 , n95 , n104 , 
n116 , n131 , n133 , n140 , n144 , n157 , n167 , n172 , n175 , n181 , 
n182 , n183 , n205 , n210 , n216 , n225 , n260 , n266 , n275 , n281 , 
n286 , n293 , n297 , n299 , n315 , n318 , n325 , n344 , n362 , n402 , 
n418 , n427 , n432 , n433 , n439 , n441 , n442 , n445 , n447 , n463 , 
n466 , n470 , n476 , n484 , n490 , n492 , n494 , n502 , n509 , n521 ;
    output n3 , n6 , n13 , n32 , n44 , n51 , n55 , n57 , n58 , 
n62 , n64 , n83 , n86 , n103 , n110 , n129 , n130 , n136 , n164 , 
n196 , n213 , n229 , n234 , n236 , n257 , n272 , n274 , n276 , n289 , 
n332 , n334 , n340 , n357 , n365 , n375 , n397 , n404 , n406 , n414 , 
n434 , n450 , n455 , n471 , n488 , n511 , n512 , n520 ;
    wire n0 , n1 , n2 , n4 , n5 , n7 , n8 , n9 , n10 , 
n11 , n12 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , 
n22 , n23 , n24 , n26 , n28 , n29 , n30 , n31 , n33 , n34 , 
n35 , n36 , n37 , n38 , n39 , n42 , n43 , n45 , n46 , n47 , 
n48 , n49 , n50 , n52 , n53 , n54 , n56 , n59 , n61 , n63 , 
n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , 
n75 , n76 , n77 , n78 , n79 , n81 , n82 , n84 , n85 , n87 , 
n88 , n89 , n90 , n91 , n92 , n94 , n96 , n97 , n98 , n99 , 
n100 , n101 , n102 , n105 , n106 , n107 , n108 , n109 , n111 , n112 , 
n113 , n114 , n115 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , 
n124 , n125 , n126 , n127 , n128 , n132 , n134 , n135 , n137 , n138 , 
n139 , n141 , n142 , n143 , n145 , n146 , n147 , n148 , n149 , n150 , 
n151 , n152 , n153 , n154 , n155 , n156 , n158 , n159 , n160 , n161 , 
n162 , n163 , n165 , n166 , n168 , n169 , n170 , n171 , n173 , n174 , 
n176 , n177 , n178 , n179 , n180 , n184 , n185 , n186 , n187 , n188 , 
n189 , n190 , n191 , n192 , n193 , n194 , n195 , n197 , n198 , n199 , 
n200 , n201 , n202 , n203 , n204 , n206 , n207 , n208 , n209 , n211 , 
n212 , n214 , n215 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , 
n224 , n226 , n227 , n228 , n230 , n231 , n232 , n233 , n235 , n237 , 
n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , 
n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n258 , 
n259 , n261 , n262 , n263 , n264 , n265 , n267 , n268 , n269 , n270 , 
n271 , n273 , n277 , n278 , n279 , n280 , n282 , n283 , n284 , n285 , 
n287 , n288 , n290 , n291 , n292 , n294 , n295 , n296 , n298 , n300 , 
n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , 
n311 , n312 , n313 , n314 , n316 , n317 , n319 , n320 , n321 , n322 , 
n323 , n324 , n326 , n327 , n328 , n329 , n330 , n331 , n333 , n335 , 
n336 , n337 , n338 , n339 , n341 , n342 , n343 , n345 , n346 , n347 , 
n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n358 , 
n359 , n360 , n361 , n363 , n364 , n366 , n367 , n368 , n369 , n370 , 
n371 , n372 , n373 , n374 , n376 , n377 , n378 , n379 , n380 , n381 , 
n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , 
n392 , n393 , n394 , n395 , n396 , n398 , n399 , n400 , n401 , n403 , 
n405 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n415 , n416 , 
n417 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n428 , 
n429 , n430 , n431 , n435 , n436 , n437 , n438 , n440 , n443 , n444 , 
n446 , n448 , n449 , n451 , n452 , n453 , n454 , n456 , n457 , n458 , 
n459 , n460 , n461 , n462 , n464 , n465 , n467 , n468 , n469 , n472 , 
n473 , n474 , n475 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , 
n485 , n486 , n487 , n489 , n491 , n493 , n495 , n496 , n497 , n498 , 
n499 , n500 , n501 , n503 , n504 , n505 , n506 , n507 , n508 , n510 , 
n513 , n514 , n515 , n516 , n517 , n518 , n519 , n522 , n523 , n524 , 
n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , 
n535 , n536 , n537 ;
    xnor g0 ( n389 , n93 , n133 );
    not g1 ( n351 , n482 );
    xnor g2 ( n124 , n232 , n40 );
    and g3 ( n143 , n260 , n447 );
    xnor g4 ( n16 , n378 , n151 );
    and g5 ( n535 , n476 , n183 );
    and g6 ( n139 , n447 , n402 );
    not g7 ( n276 , n144 );
    and g8 ( n251 , n259 , n531 );
    nor g9 ( n156 , n518 , n383 );
    nor g10 ( n117 , n249 , n534 );
    or g11 ( n98 , n227 , n235 );
    and g12 ( n285 , n176 , n338 );
    xnor g13 ( n446 , n338 , n176 );
    nor g14 ( n312 , n447 , n166 );
    xnor g15 ( n272 , n270 , n361 );
    not g16 ( n146 , n175 );
    not g17 ( n471 , n534 );
    or g18 ( n77 , n393 , n312 );
    nor g19 ( n26 , n132 , n85 );
    not g20 ( n248 , n484 );
    xnor g21 ( n187 , n222 , n502 );
    not g22 ( n336 , n168 );
    not g23 ( n300 , n152 );
    and g24 ( n527 , n155 , n138 );
    or g25 ( n219 , n164 , n176 );
    not g26 ( n134 , n2 );
    or g27 ( n488 , n74 , n37 );
    and g28 ( n67 , n345 , n349 );
    not g29 ( n290 , n172 );
    and g30 ( n499 , n268 , n517 );
    or g31 ( n102 , n447 , n342 );
    and g32 ( n192 , n290 , n350 );
    not g33 ( n37 , n66 );
    not g34 ( n135 , n447 );
    xnor g35 ( n237 , n108 , n389 );
    buf g36 ( n86 , n0 );
    not g37 ( n14 , n516 );
    not g38 ( n378 , n267 );
    not g39 ( n491 , n24 );
    or g40 ( n320 , n241 , n39 );
    not g41 ( n368 , n80 );
    not g42 ( n105 , n56 );
    xnor g43 ( n533 , n468 , n523 );
    or g44 ( n347 , n113 , n152 );
    xnor g45 ( n166 , n215 , n492 );
    or g46 ( n152 , n206 , n505 );
    and g47 ( n241 , n95 , n447 );
    or g48 ( n340 , n477 , n36 );
    nor g49 ( n74 , n465 , n194 );
    or g50 ( n416 , n276 , n458 );
    xnor g51 ( n57 , n231 , n400 );
    or g52 ( n309 , n305 , n385 );
    nor g53 ( n384 , n183 , n476 );
    and g54 ( n515 , n222 , n343 );
    not g55 ( n481 , n124 );
    nor g56 ( n437 , n447 , n237 );
    and g57 ( n12 , n125 , n153 );
    or g58 ( n343 , n60 , n502 );
    xnor g59 ( n55 , n524 , n49 );
    xnor g60 ( n240 , n59 , n86 );
    and g61 ( n345 , n469 , n447 );
    not g62 ( n404 , n144 );
    or g63 ( n9 , n498 , n392 );
    and g64 ( n159 , n367 , n394 );
    nor g65 ( n269 , n503 , n516 );
    or g66 ( n267 , n180 , n264 );
    not g67 ( n501 , n252 );
    xnor g68 ( n204 , n425 , n218 );
    nor g69 ( n20 , n144 , n447 );
    xor g70 ( n323 , n526 , n133 );
    or g71 ( n360 , n37 , n294 );
    not g72 ( n397 , n328 );
    nor g73 ( n217 , n534 , n165 );
    and g74 ( n352 , n486 , n219 );
    and g75 ( n200 , n439 , n447 );
    and g76 ( n82 , n281 , n447 );
    not g77 ( n21 , n318 );
    xnor g78 ( n262 , n50 , n207 );
    nor g79 ( n218 , n217 , n36 );
    xor g80 ( n252 , n417 , n442 );
    nor g81 ( n53 , n121 , n221 );
    or g82 ( n295 , n118 , n336 );
    or g83 ( n500 , n444 , n8 );
    not g84 ( n189 , n275 );
    or g85 ( n465 , n139 , n20 );
    xnor g86 ( n88 , n38 , n502 );
    or g87 ( n339 , n468 , n523 );
    or g88 ( n451 , n242 , n31 );
    or g89 ( n230 , n30 , n515 );
    or g90 ( n495 , n487 , n464 );
    or g91 ( n115 , n88 , n329 );
    or g92 ( n274 , n506 , n518 );
    not g93 ( n169 , n507 );
    not g94 ( n304 , n396 );
    or g95 ( n50 , n395 , n35 );
    or g96 ( n319 , n46 , n87 );
    xnor g97 ( n390 , n178 , n344 );
    and g98 ( n393 , n140 , n447 );
    nor g99 ( n380 , n149 , n517 );
    not g100 ( n305 , n286 );
    not g101 ( n113 , n267 );
    xnor g102 ( n120 , n211 , n476 );
    and g103 ( n507 , n263 , n228 );
    xnor g104 ( n209 , n385 , n286 );
    or g105 ( n63 , n482 , n50 );
    not g106 ( n202 , n55 );
    and g107 ( n430 , n163 , n360 );
    or g108 ( n222 , n245 , n73 );
    not g109 ( n106 , n490 );
    or g110 ( n155 , n46 , n7 );
    and g111 ( n426 , n532 , n347 );
    or g112 ( n440 , n525 , n76 );
    or g113 ( n403 , n296 , n251 );
    or g114 ( n520 , n247 , n123 );
    not g115 ( n45 , n465 );
    or g116 ( n511 , n376 , n308 );
    and g117 ( n529 , n122 , n337 );
    not g118 ( n282 , n306 );
    and g119 ( n242 , n181 , n490 );
    or g120 ( n314 , n462 , n530 );
    and g121 ( n48 , n522 , n443 );
    or g122 ( n153 , n131 , n293 );
    xnor g123 ( n94 , n353 , n15 );
    and g124 ( n35 , n324 , n359 );
    not g125 ( n477 , n351 );
    or g126 ( n454 , n161 , n239 );
    nor g127 ( n73 , n192 , n353 );
    nor g128 ( n421 , n201 , n97 );
    or g129 ( n44 , n224 , n184 );
    not g130 ( n422 , n436 );
    and g131 ( n493 , n67 , n503 );
    and g132 ( n158 , n209 , n387 );
    and g133 ( n448 , n199 , n443 );
    or g134 ( n215 , n535 , n372 );
    and g135 ( n288 , n416 , n450 );
    not g136 ( n311 , n482 );
    xnor g137 ( n38 , n327 , n299 );
    not g138 ( n341 , n375 );
    and g139 ( n420 , n63 , n168 );
    nor g140 ( n510 , n266 , n132 );
    not g141 ( n114 , n320 );
    not g142 ( n193 , n325 );
    or g143 ( n142 , n429 , n437 );
    and g144 ( n268 , n75 , n212 );
    nor g145 ( n407 , n447 , n262 );
    and g146 ( n239 , n89 , n265 );
    or g147 ( n307 , n128 , n56 );
    and g148 ( n398 , n430 , n507 );
    and g149 ( n126 , n445 , n144 );
    or g150 ( n163 , n489 , n317 );
    buf g151 ( n434 , 1'b0 );
    not g152 ( n3 , n501 );
    and g153 ( n29 , n94 , n42 );
    xnor g154 ( n208 , n481 , n324 );
    or g155 ( n179 , n449 , n71 );
    not g156 ( n503 , n77 );
    xnor g157 ( n22 , n321 , n318 );
    not g158 ( n101 , n315 );
    or g159 ( n327 , n377 , n12 );
    or g160 ( n108 , n137 , n189 );
    or g161 ( n28 , n148 , n24 );
    not g162 ( n524 , n534 );
    nor g163 ( n211 , n85 , n510 );
    not g164 ( n474 , n203 );
    not g165 ( n387 , n447 );
    or g166 ( n321 , n368 , n52 );
    and g167 ( n513 , n300 , n378 );
    not g168 ( n425 , n396 );
    or g169 ( n415 , n193 , n54 );
    and g170 ( n254 , n316 , n447 );
    and g171 ( n278 , n148 , n447 );
    and g172 ( n431 , n5 , n1 );
    or g173 ( n263 , n447 , n223 );
    xnor g174 ( n196 , n438 , n86 );
    and g175 ( n475 , n54 , n193 );
    or g176 ( n486 , n386 , n177 );
    and g177 ( n417 , n299 , n327 );
    or g178 ( n91 , n45 , n194 );
    or g179 ( n409 , n42 , n288 );
    not g180 ( n436 , n4 );
    xnor g181 ( n6 , n24 , n214 );
    xnor g182 ( n234 , n425 , n279 );
    nor g183 ( n271 , n27 , n266 );
    not g184 ( n145 , n144 );
    not g185 ( n291 , n124 );
    not g186 ( n277 , n470 );
    or g187 ( n122 , n364 , n147 );
    and g188 ( n356 , n367 , n10 );
    not g189 ( n292 , n301 );
    xnor g190 ( n64 , n255 , n162 );
    not g191 ( n405 , n118 );
    nor g192 ( n435 , n135 , n499 );
    or g193 ( n358 , n315 , n422 );
    not g194 ( n349 , n478 );
    not g195 ( n90 , n491 );
    not g196 ( n270 , n77 );
    and g197 ( n326 , n68 , n179 );
    not g198 ( n449 , n266 );
    and g199 ( n245 , n172 , n509 );
    or g200 ( n337 , n101 , n19 );
    or g201 ( n125 , n242 , n33 );
    or g202 ( n414 , n254 , n280 );
    not g203 ( n382 , n447 );
    not g204 ( n443 , n447 );
    not g205 ( n505 , n356 );
    not g206 ( n413 , n11 );
    xnor g207 ( n226 , n326 , n183 );
    or g208 ( n141 , n277 , n202 );
    xnor g209 ( n154 , n104 , n315 );
    xor g210 ( n43 , n309 , n116 );
    and g211 ( n284 , n99 , n10 );
    not g212 ( n255 , n114 );
    or g213 ( n265 , n133 , n184 );
    and g214 ( n482 , n232 , n40 );
    xnor g215 ( n406 , n23 , n508 );
    xnor g216 ( n0 , n220 , n293 );
    nor g217 ( n253 , n172 , n4 );
    not g218 ( n366 , n485 );
    nor g219 ( n34 , n447 , n371 );
    or g220 ( n58 , n493 , n500 );
    or g221 ( n10 , n143 , n310 );
    or g222 ( n52 , n84 , n453 );
    and g223 ( n335 , n157 , n447 );
    not g224 ( n42 , n534 );
    not g225 ( n532 , n376 );
    not g226 ( n394 , n10 );
    not g227 ( n396 , n291 );
    nor g228 ( n514 , n447 , n307 );
    not g229 ( n164 , n292 );
    not g230 ( n174 , n215 );
    or g231 ( n357 , n117 , n283 );
    or g232 ( n68 , n271 , n529 );
    and g233 ( n232 , n126 , n210 );
    not g234 ( n212 , n92 );
    xnor g235 ( n32 , n151 , n426 );
    or g236 ( n330 , n21 , n321 );
    nor g237 ( n224 , n463 , n47 );
    not g238 ( n526 , n170 );
    not g239 ( n467 , n521 );
    or g240 ( n459 , n496 , n127 );
    or g241 ( n11 , n46 , n528 );
    not g242 ( n338 , n331 );
    and g243 ( n30 , n502 , n60 );
    nor g244 ( n75 , n516 , n28 );
    not g245 ( n128 , n507 );
    nor g246 ( n15 , n245 , n192 );
    and g247 ( n261 , n171 , n267 );
    not g248 ( n469 , n148 );
    not g249 ( n170 , n536 );
    or g250 ( n24 , n335 , n48 );
    not g251 ( n350 , n509 );
    or g252 ( n151 , n82 , n158 );
    nor g253 ( n17 , n447 , n208 );
    or g254 ( n359 , n397 , n320 );
    and g255 ( n201 , n428 , n90 );
    not g256 ( n355 , n47 );
    nor g257 ( n313 , n447 , n388 );
    not g258 ( n331 , n301 );
    and g259 ( n487 , n173 , n150 );
    xnor g260 ( n369 , n252 , n419 );
    or g261 ( n176 , n277 , n341 );
    and g262 ( n231 , n373 , n404 );
    and g263 ( n310 , n22 , n127 );
    or g264 ( n69 , n471 , n94 );
    not g265 ( n496 , n362 );
    nor g266 ( n537 , n93 , n133 );
    or g267 ( n78 , n86 , n59 );
    not g268 ( n346 , n93 );
    or g269 ( n149 , n199 , n366 );
    or g270 ( n329 , n253 , n314 );
    and g271 ( n353 , n96 , n415 );
    xnor g272 ( n13 , n319 , n369 );
    not g273 ( n71 , n27 );
    xnor g274 ( n365 , n477 , n472 );
    nor g275 ( n361 , n278 , n448 );
    not g276 ( n190 , n344 );
    or g277 ( n100 , n408 , n160 );
    and g278 ( n429 , n432 , n447 );
    not g279 ( n328 , n291 );
    nor g280 ( n464 , n489 , n412 );
    and g281 ( n423 , n390 , n531 );
    not g282 ( n19 , n104 );
    nor g283 ( n162 , n247 , n17 );
    or g284 ( n8 , n354 , n250 );
    and g285 ( n408 , n392 , n450 );
    not g286 ( n236 , n479 );
    and g287 ( n287 , n495 , n72 );
    not g288 ( n84 , n466 );
    and g289 ( n247 , n398 , n447 );
    xnor g290 ( n62 , n3 , n120 );
    and g291 ( n111 , n128 , n65 );
    nor g292 ( n171 , n300 , n186 );
    and g293 ( n303 , n523 , n397 );
    nor g294 ( n283 , n2 , n416 );
    or g295 ( n453 , n190 , n178 );
    and g296 ( n370 , n454 , n358 );
    nor g297 ( n456 , n447 , n43 );
    and g298 ( n462 , n422 , n172 );
    and g299 ( n81 , n433 , n447 );
    xnor g300 ( n334 , n145 , n333 );
    not g301 ( n199 , n420 );
    not g302 ( n188 , n25 );
    xnor g303 ( n227 , n79 , n521 );
    or g304 ( n1 , n480 , n18 );
    xnor g305 ( n110 , n486 , n446 );
    or g306 ( n508 , n16 , n426 );
    buf g307 ( n534 , n107 );
    not g308 ( n92 , n270 );
    and g309 ( n97 , n268 , n447 );
    and g310 ( n367 , n371 , n379 );
    and g311 ( n147 , n119 , n410 );
    xnor g312 ( n472 , n230 , n61 );
    or g313 ( n289 , n345 , n195 );
    or g314 ( n497 , n29 , n483 );
    not g315 ( n379 , n447 );
    and g316 ( n316 , n499 , n394 );
    or g317 ( n391 , n467 , n248 );
    or g318 ( n516 , n457 , n423 );
    not g319 ( n478 , n14 );
    and g320 ( n264 , n461 , n135 );
    and g321 ( n118 , n114 , n398 );
    xor g322 ( n136 , n238 , n348 );
    xnor g323 ( n56 , n458 , n495 );
    not g324 ( n306 , n79 );
    not g325 ( n273 , n203 );
    or g326 ( n72 , n65 , n169 );
    nor g327 ( n214 , n493 , n428 );
    xnor g328 ( n322 , n504 , n205 );
    not g329 ( n512 , n445 );
    xnor g330 ( n388 , n226 , n476 );
    and g331 ( n233 , n420 , n379 );
    or g332 ( n195 , n191 , n407 );
    xnor g333 ( n51 , n221 , n323 );
    not g334 ( n489 , n142 );
    and g335 ( n160 , n9 , n231 );
    not g336 ( n460 , n492 );
    xnor g337 ( n455 , n141 , n240 );
    not g338 ( n7 , n57 );
    not g339 ( n138 , n170 );
    nor g340 ( n372 , n384 , n326 );
    not g341 ( n203 , n2 );
    or g342 ( n221 , n137 , n83 );
    and g343 ( n457 , n297 , n447 );
    not g344 ( n130 , n311 );
    xnor g345 ( n392 , n391 , n411 );
    and g346 ( n180 , n216 , n447 );
    not g347 ( n373 , n333 );
    nor g348 ( n197 , n382 , n66 );
    and g349 ( n518 , n413 , n47 );
    or g350 ( n213 , n130 , n204 );
    xnor g351 ( n107 , n126 , n210 );
    xnor g352 ( n374 , n330 , n418 );
    and g353 ( n371 , n380 , n90 );
    and g354 ( n377 , n293 , n131 );
    or g355 ( n96 , n475 , n391 );
    xnor g356 ( n70 , n27 , n266 );
    xnor g357 ( n438 , n239 , n315 );
    xor g358 ( n235 , n138 , n494 );
    xnor g359 ( n375 , n497 , n533 );
    xnor g360 ( n2 , n144 , n445 );
    or g361 ( n228 , n302 , n379 );
    not g362 ( n244 , n370 );
    and g363 ( n296 , n225 , n447 );
    not g364 ( n184 , n221 );
    or g365 ( n238 , n399 , n424 );
    xnor g366 ( n523 , n187 , n60 );
    not g367 ( n150 , n431 );
    not g368 ( n79 , n355 );
    xnor g369 ( n522 , n453 , n466 );
    and g370 ( n424 , n374 , n382 );
    and g371 ( n483 , n100 , n69 );
    not g372 ( n517 , n403 );
    or g373 ( n89 , n479 , n53 );
    or g374 ( n185 , n198 , n330 );
    xor g375 ( n109 , n518 , n155 );
    or g376 ( n410 , n346 , n121 );
    and g377 ( n395 , n255 , n304 );
    not g378 ( n246 , n182 );
    not g379 ( n83 , n282 );
    and g380 ( n376 , n186 , n113 );
    and g381 ( n381 , n497 , n339 );
    and g382 ( n399 , n167 , n447 );
    not g383 ( n127 , n447 );
    not g384 ( n480 , n41 );
    or g385 ( n308 , n513 , n261 );
    or g386 ( n178 , n460 , n174 );
    xnor g387 ( n49 , n94 , n100 );
    xnor g388 ( n229 , n403 , n421 );
    nor g389 ( n161 , n101 , n86 );
    and g390 ( n354 , n519 , n212 );
    not g391 ( n4 , n0 );
    not g392 ( n137 , n463 );
    xnor g393 ( n243 , n529 , n70 );
    xnor g394 ( n461 , n185 , n182 );
    and g395 ( n412 , n431 , n91 );
    not g396 ( n452 , n475 );
    not g397 ( n536 , n479 );
    or g398 ( n504 , n303 , n381 );
    nor g399 ( n364 , n104 , n315 );
    nor g400 ( n383 , n236 , n155 );
    and g401 ( n506 , n11 , n306 );
    xnor g402 ( n333 , n484 , n521 );
    xor g403 ( n530 , n252 , n205 );
    and g404 ( n428 , n233 , n485 );
    and g405 ( n194 , n102 , n459 );
    or g406 ( n119 , n537 , n108 );
    not g407 ( n468 , n124 );
    not g408 ( n206 , n238 );
    and g409 ( n36 , n409 , n481 );
    not g410 ( n458 , n534 );
    xnor g411 ( n401 , n294 , n363 );
    xnor g412 ( n479 , n298 , n451 );
    not g413 ( n87 , n365 );
    and g414 ( n386 , n59 , n86 );
    not g415 ( n301 , n38 );
    or g416 ( n324 , n111 , n287 );
    and g417 ( n444 , n269 , n233 );
    xnor g418 ( n257 , n26 , n266 );
    or g419 ( n59 , n527 , n156 );
    nor g420 ( n76 , n447 , n105 );
    or g421 ( n298 , n146 , n188 );
    and g422 ( n485 , n478 , n77 );
    not g423 ( n498 , n273 );
    xnor g424 ( n342 , n275 , n463 );
    nor g425 ( n249 , n445 , n145 );
    xnor g426 ( n400 , n498 , n392 );
    not g427 ( n54 , n494 );
    xnor g428 ( n61 , n322 , n427 );
    and g429 ( n473 , n194 , n465 );
    and g430 ( n85 , n244 , n164 );
    xor g431 ( n207 , n311 , n336 );
    nor g432 ( n33 , n31 , n298 );
    and g433 ( n31 , n106 , n112 );
    and g434 ( n132 , n370 , n38 );
    not g435 ( n18 , n447 );
    not g436 ( n302 , n441 );
    or g437 ( n419 , n285 , n352 );
    xnor g438 ( n223 , n147 , n154 );
    and g439 ( n256 , n440 , n169 );
    xnor g440 ( n47 , n175 , n25 );
    not g441 ( n65 , n534 );
    nor g442 ( n258 , n447 , n91 );
    not g443 ( n528 , n334 );
    nor g444 ( n250 , n366 , n233 );
    nor g445 ( n525 , n18 , n430 );
    xnor g446 ( n220 , n125 , n131 );
    or g447 ( n5 , n447 , n165 );
    not g448 ( n165 , n134 );
    or g449 ( n168 , n81 , n313 );
    and g450 ( n317 , n150 , n473 );
    and g451 ( n177 , n78 , n141 );
    not g452 ( n198 , n418 );
    xnor g453 ( n259 , n52 , n80 );
    xnor g454 ( n279 , n524 , n288 );
    not g455 ( n450 , n474 );
    not g456 ( n66 , n473 );
    not g457 ( n112 , n181 );
    or g458 ( n123 , n514 , n256 );
    not g459 ( n121 , n133 );
    or g460 ( n280 , n159 , n284 );
    not g461 ( n531 , n447 );
    or g462 ( n348 , n356 , n254 );
    or g463 ( n99 , n34 , n435 );
    not g464 ( n173 , n91 );
    nor g465 ( n519 , n349 , n345 );
    and g466 ( n186 , n254 , n206 );
    xnor g467 ( n103 , n526 , n109 );
    nor g468 ( n332 , n98 , n115 );
    or g469 ( n148 , n405 , n168 );
    not g470 ( n294 , n431 );
    nor g471 ( n191 , n387 , n295 );
    nor g472 ( n39 , n447 , n243 );
    xnor g473 ( n129 , n142 , n401 );
    not g474 ( n46 , n470 );
    and g475 ( n411 , n415 , n452 );
    or g476 ( n363 , n197 , n258 );
    or g477 ( n23 , n200 , n456 );
    or g478 ( n385 , n246 , n185 );
endmodule
