module top( n55 , n94 , n249 , n280 , n550 , n563 , n593 , n637 , n1171 , 
n1227 , n1234 , n1507 , n1548 , n1579 , n1624 , n1643 , n1872 , n1970 , n1971 , 
n2199 , n2407 , n2492 , n2769 , n3186 , n3789 , n3940 , n3997 , n4059 , n4140 , 
n4147 , n4197 , n4278 , n4301 , n4309 , n4535 , n4660 , n5250 , n5432 , n5605 , 
n5813 , n5816 , n5896 , n5964 , n6212 , n6358 , n6502 , n6818 , n6963 , n6968 , 
n7106 , n7305 , n7356 , n7362 , n7458 , n7839 , n7946 , n8220 , n8494 , n8627 , 
n9144 , n9147 , n9177 , n9285 , n9309 , n9604 , n9641 , n9996 , n10196 , n10598 , 
n10625 , n11134 , n11297 , n11416 , n11457 , n11508 , n11588 , n11787 , n12133 , n12421 , 
n12725 , n13134 , n13295 , n13454 , n13613 , n13820 , n13989 , n14042 , n14180 , n14186 , 
n14308 , n14344 , n14471 , n14707 , n15027 , n15046 , n15070 , n15710 , n15851 , n16058 , 
n16560 , n16598 , n16780 , n16999 , n17120 , n17193 , n17358 , n17421 , n17489 , n17516 , 
n17744 , n17774 , n17776 , n18212 , n18236 , n18405 , n18683 , n18866 , n18953 , n19080 , 
n19221 , n19367 , n19580 , n19744 , n19747 , n19754 , n20078 , n20140 , n20260 , n20288 , 
n20363 , n20662 , n20672 , n20921 , n20949 , n21548 , n21703 , n21958 , n22361 , n23017 , 
n23032 , n23150 , n23161 , n23871 , n23880 , n23895 , n23981 , n24622 , n24626 , n24868 , 
n25069 , n25123 , n25303 , n25407 , n25549 , n25588 , n25636 , n25936 , n27028 , n27239 , 
n27268 , n27311 , n27400 , n27663 , n27666 , n27884 , n27892 , n27942 , n27990 , n28064 , 
n28239 , n28500 , n28518 , n28523 , n28755 , n29027 , n29147 , n29214 , n29640 , n29719 , 
n29808 , n29816 , n30030 , n30071 , n30175 , n30892 , n31222 , n31241 , n31263 , n31478 , 
n31827 , n31920 , n32088 , n32277 , n32698 , n33134 , n33257 , n33699 , n33981 , n33999 , 
n34021 , n34053 , n34136 , n34267 , n34292 , n34561 , n34565 , n34573 , n34590 , n34653 , 
n34686 , n34788 , n34955 , n34963 , n34997 , n35104 , n35301 , n35411 , n35732 , n36117 , 
n36230 , n36514 , n36687 , n36693 , n36903 , n37434 , n37890 , n38016 , n38157 , n38217 , 
n38527 , n38813 , n38819 , n38879 , n38894 , n38920 , n39213 , n39266 , n39309 , n39450 , 
n39536 , n40152 , n40220 , n40560 , n40586 , n40907 , n40979 , n41277 , n41315 , n41487 , 
n41534 , n41700 , n41767 , n42232 , n42248 , n42278 , n42523 );
    input n55 , n249 , n280 , n563 , n637 , n1171 , n1234 , n1507 , n1643 , 
n1971 , n2199 , n2769 , n3186 , n3940 , n3997 , n4140 , n4147 , n4278 , n4309 , 
n5250 , n5605 , n5816 , n5896 , n5964 , n6212 , n6502 , n6818 , n6968 , n7106 , 
n7305 , n7356 , n7362 , n7946 , n8494 , n8627 , n9147 , n9285 , n9604 , n9641 , 
n10598 , n11297 , n11787 , n12421 , n12725 , n13454 , n13613 , n13989 , n14042 , n14180 , 
n14186 , n14471 , n14707 , n15070 , n16058 , n16598 , n16780 , n17120 , n17193 , n17489 , 
n17516 , n17744 , n17774 , n18212 , n18683 , n18866 , n18953 , n19221 , n19367 , n19580 , 
n19747 , n20140 , n20363 , n20949 , n22361 , n23032 , n23150 , n23871 , n23981 , n24622 , 
n24868 , n25069 , n25123 , n25588 , n25936 , n27892 , n27942 , n28518 , n28755 , n29640 , 
n29719 , n29808 , n29816 , n30892 , n31222 , n31827 , n32277 , n33981 , n34021 , n34053 , 
n34136 , n34292 , n34565 , n34590 , n34653 , n34686 , n34788 , n35104 , n35301 , n35411 , 
n36117 , n36230 , n38016 , n38157 , n38217 , n38819 , n38879 , n38894 , n38920 , n39266 , 
n39309 , n39450 , n40152 , n40586 , n40907 , n40979 , n41277 , n41534 , n42248 ;
    output n94 , n550 , n593 , n1227 , n1548 , n1579 , n1624 , n1872 , n1970 , 
n2407 , n2492 , n3789 , n4059 , n4197 , n4301 , n4535 , n4660 , n5432 , n5813 , 
n6358 , n6963 , n7458 , n7839 , n8220 , n9144 , n9177 , n9309 , n9996 , n10196 , 
n10625 , n11134 , n11416 , n11457 , n11508 , n11588 , n12133 , n13134 , n13295 , n13820 , 
n14308 , n14344 , n15027 , n15046 , n15710 , n15851 , n16560 , n16999 , n17358 , n17421 , 
n17776 , n18236 , n18405 , n19080 , n19744 , n19754 , n20078 , n20260 , n20288 , n20662 , 
n20672 , n20921 , n21548 , n21703 , n21958 , n23017 , n23161 , n23880 , n23895 , n24626 , 
n25303 , n25407 , n25549 , n25636 , n27028 , n27239 , n27268 , n27311 , n27400 , n27663 , 
n27666 , n27884 , n27990 , n28064 , n28239 , n28500 , n28523 , n29027 , n29147 , n29214 , 
n30030 , n30071 , n30175 , n31241 , n31263 , n31478 , n31920 , n32088 , n32698 , n33134 , 
n33257 , n33699 , n33999 , n34267 , n34561 , n34573 , n34955 , n34963 , n34997 , n35732 , 
n36514 , n36687 , n36693 , n36903 , n37434 , n37890 , n38527 , n38813 , n39213 , n39536 , 
n40220 , n40560 , n41315 , n41487 , n41700 , n41767 , n42232 , n42278 , n42523 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , 
n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , 
n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , 
n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , 
n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , 
n49 , n50 , n51 , n52 , n53 , n54 , n56 , n57 , n58 , n59 , 
n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
n90 , n91 , n92 , n93 , n95 , n96 , n97 , n98 , n99 , n100 , 
n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n250 , n251 , 
n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , 
n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , 
n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n281 , n282 , 
n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , 
n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , 
n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , 
n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , 
n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , 
n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , 
n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , 
n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , 
n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , 
n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , 
n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , 
n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , 
n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , 
n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , 
n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , 
n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , 
n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , 
n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , 
n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , 
n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , 
n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , 
n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , 
n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , 
n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , 
n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , 
n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , 
n543 , n544 , n545 , n546 , n547 , n548 , n549 , n551 , n552 , n553 , 
n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n564 , 
n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , 
n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n594 , n595 , 
n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , 
n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , 
n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , 
n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , 
n636 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , 
n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , 
n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , 
n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , 
n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , 
n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , 
n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , 
n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , 
n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , 
n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , 
n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , 
n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , 
n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , 
n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , 
n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , 
n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , 
n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , 
n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , 
n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , 
n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , 
n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , 
n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , 
n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , 
n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , 
n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , 
n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , 
n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , 
n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , 
n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , 
n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , 
n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , 
n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , 
n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , 
n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , 
n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , 
n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , 
n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , 
n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , 
n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , 
n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , 
n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , 
n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , 
n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , 
n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , 
n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , 
n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , 
n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , 
n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , 
n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , 
n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , 
n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , 
n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , 
n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , 
n1167 , n1168 , n1169 , n1170 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , 
n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , 
n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , 
n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , 
n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , 
n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1228 , 
n1229 , n1230 , n1231 , n1232 , n1233 , n1235 , n1236 , n1237 , n1238 , n1239 , 
n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1508 , n1509 , n1510 , 
n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , 
n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , 
n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , 
n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1549 , n1550 , n1551 , 
n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , 
n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , 
n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1580 , n1581 , n1582 , 
n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , 
n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , 
n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , 
n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , 
n1623 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , 
n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1644 , 
n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , 
n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , 
n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , 
n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , 
n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , 
n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , 
n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , 
n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , 
n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , 
n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , 
n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , 
n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , 
n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , 
n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , 
n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , 
n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , 
n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , 
n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , 
n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , 
n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , 
n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , 
n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , 
n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1873 , n1874 , n1875 , 
n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , 
n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , 
n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , 
n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , 
n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , 
n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , 
n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , 
n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , 
n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , 
n1966 , n1967 , n1968 , n1969 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , 
n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , 
n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , 
n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , 
n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , 
n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , 
n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , 
n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , 
n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , 
n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , 
n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , 
n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , 
n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , 
n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , 
n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , 
n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , 
n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , 
n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , 
n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , 
n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , 
n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , 
n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , 
n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , 
n2198 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , 
n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , 
n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , 
n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , 
n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , 
n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , 
n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , 
n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , 
n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , 
n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , 
n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , 
n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , 
n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , 
n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , 
n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , 
n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , 
n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , 
n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , 
n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , 
n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , 
n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2408 , n2409 , 
n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
n2490 , n2491 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , 
n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , 
n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , 
n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , 
n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , 
n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , 
n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , 
n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , 
n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , 
n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , 
n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , 
n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , 
n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , 
n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , 
n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , 
n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , 
n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , 
n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , 
n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , 
n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , 
n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , 
n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , 
n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , 
n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , 
n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , 
n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , 
n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2770 , n2771 , 
n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , 
n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , 
n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , 
n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , 
n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , 
n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , 
n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , 
n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , 
n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , 
n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , 
n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , 
n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , 
n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , 
n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , 
n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , 
n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , 
n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , 
n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , 
n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , 
n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , 
n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , 
n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , 
n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , 
n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , 
n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , 
n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , 
n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , 
n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , 
n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , 
n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , 
n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , 
n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , 
n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , 
n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , 
n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , 
n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , 
n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , 
n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , 
n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , 
n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , 
n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , 
n3182 , n3183 , n3184 , n3185 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , 
n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , 
n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , 
n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , 
n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , 
n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , 
n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , 
n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , 
n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , 
n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , 
n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , 
n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , 
n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , 
n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , 
n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , 
n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , 
n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , 
n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , 
n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , 
n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , 
n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , 
n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , 
n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , 
n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , 
n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , 
n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , 
n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , 
n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , 
n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , 
n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , 
n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , 
n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , 
n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , 
n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , 
n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , 
n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , 
n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , 
n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , 
n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , 
n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , 
n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , 
n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , 
n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , 
n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , 
n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , 
n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , 
n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , 
n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , 
n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , 
n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , 
n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , 
n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , 
n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , 
n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , 
n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , 
n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , 
n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , 
n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , 
n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , 
n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , 
n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3790 , n3791 , n3792 , n3793 , 
n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , 
n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , 
n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , 
n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , 
n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , 
n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , 
n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , 
n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , 
n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , 
n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , 
n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , 
n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , 
n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , 
n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , 
n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3941 , n3942 , n3943 , n3944 , 
n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , 
n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , 
n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , 
n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , 
n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , 
n3995 , n3996 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , 
n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , 
n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , 
n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , 
n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , 
n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , 
n4056 , n4057 , n4058 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , 
n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , 
n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , 
n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , 
n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , 
n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , 
n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , 
n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , 
n4137 , n4138 , n4139 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4148 , 
n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , 
n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , 
n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , 
n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , 
n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4198 , n4199 , 
n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , 
n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , 
n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , 
n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , 
n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , 
n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , 
n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , 
n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4279 , n4280 , 
n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , 
n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , 
n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4310 , n4311 , n4312 , 
n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , 
n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , 
n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , 
n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , 
n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , 
n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , 
n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , 
n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , 
n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , 
n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , 
n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , 
n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , 
n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , 
n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , 
n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , 
n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , 
n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , 
n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , 
n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , 
n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , 
n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , 
n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , 
n4533 , n4534 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , 
n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , 
n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , 
n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , 
n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , 
n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , 
n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , 
n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , 
n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , 
n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , 
n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , 
n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , 
n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4661 , n4662 , n4663 , n4664 , 
n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , 
n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , 
n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , 
n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , 
n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , 
n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , 
n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , 
n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , 
n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , 
n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , 
n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , 
n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , 
n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , 
n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , 
n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , 
n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , 
n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , 
n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , 
n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , 
n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , 
n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , 
n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , 
n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , 
n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , 
n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , 
n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , 
n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , 
n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , 
n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , 
n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , 
n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , 
n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , 
n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , 
n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , 
n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , 
n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , 
n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , 
n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , 
n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , 
n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , 
n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , 
n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , 
n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , 
n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , 
n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , 
n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , 
n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , 
n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , 
n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , 
n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , 
n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , 
n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , 
n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , 
n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , 
n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , 
n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , 
n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , 
n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , 
n5245 , n5246 , n5247 , n5248 , n5249 , n5251 , n5252 , n5253 , n5254 , n5255 , 
n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , 
n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , 
n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , 
n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , 
n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , 
n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , 
n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , 
n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , 
n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , 
n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , 
n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , 
n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , 
n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , 
n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , 
n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , 
n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , 
n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , 
n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5433 , n5434 , n5435 , n5436 , 
n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , 
n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , 
n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , 
n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , 
n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , 
n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , 
n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , 
n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , 
n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , 
n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , 
n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , 
n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , 
n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , 
n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , 
n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , 
n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , 
n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5606 , n5607 , 
n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , 
n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , 
n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , 
n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , 
n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , 
n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , 
n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , 
n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , 
n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , 
n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , 
n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , 
n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , 
n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , 
n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , 
n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , 
n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , 
n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , 
n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , 
n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , 
n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , 
n5808 , n5809 , n5810 , n5811 , n5812 , n5814 , n5815 , n5817 , n5818 , n5819 , 
n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , 
n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , 
n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , 
n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , 
n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , 
n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , 
n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , 
n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5897 , n5898 , n5899 , n5900 , 
n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , 
n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , 
n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , 
n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , 
n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , 
n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , 
n5961 , n5962 , n5963 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , 
n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , 
n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , 
n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , 
n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , 
n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , 
n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , 
n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , 
n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , 
n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , 
n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , 
n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , 
n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , 
n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , 
n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , 
n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , 
n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , 
n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , 
n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , 
n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , 
n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , 
n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , 
n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , 
n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , 
n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , 
n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , 
n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , 
n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , 
n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , 
n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , 
n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , 
n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , 
n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , 
n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , 
n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , 
n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , 
n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , 
n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , 
n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , 
n6353 , n6354 , n6355 , n6356 , n6357 , n6359 , n6360 , n6361 , n6362 , n6363 , 
n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , 
n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , 
n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , 
n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , 
n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , 
n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , 
n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , 
n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , 
n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , 
n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , 
n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , 
n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , 
n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , 
n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6503 , n6504 , 
n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , 
n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , 
n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , 
n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , 
n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , 
n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , 
n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , 
n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , 
n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , 
n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , 
n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , 
n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , 
n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , 
n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , 
n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , 
n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , 
n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , 
n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , 
n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , 
n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , 
n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , 
n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , 
n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , 
n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , 
n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , 
n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , 
n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , 
n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , 
n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , 
n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , 
n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , 
n6815 , n6816 , n6817 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , 
n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , 
n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , 
n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , 
n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , 
n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , 
n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , 
n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , 
n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , 
n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , 
n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , 
n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , 
n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , 
n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , 
n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6964 , n6965 , n6966 , 
n6967 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , 
n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , 
n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , 
n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , 
n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , 
n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , 
n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , 
n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , 
n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , 
n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , 
n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , 
n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , 
n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , 
n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7107 , n7108 , 
n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , 
n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , 
n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , 
n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , 
n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , 
n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , 
n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , 
n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , 
n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , 
n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , 
n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , 
n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , 
n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , 
n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , 
n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , 
n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , 
n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , 
n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , 
n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , 
n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7306 , n7307 , n7308 , n7309 , 
n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , 
n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , 
n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , 
n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , 
n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7357 , n7358 , n7359 , n7360 , 
n7361 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , 
n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , 
n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , 
n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , 
n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , 
n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , 
n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , 
n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , 
n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , 
n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7459 , n7460 , n7461 , n7462 , 
n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , 
n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , 
n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , 
n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , 
n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , 
n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , 
n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , 
n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , 
n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , 
n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , 
n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , 
n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , 
n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , 
n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , 
n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , 
n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , 
n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , 
n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , 
n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , 
n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , 
n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , 
n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , 
n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , 
n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , 
n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , 
n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , 
n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , 
n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , 
n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , 
n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , 
n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , 
n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , 
n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , 
n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , 
n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , 
n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , 
n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , 
n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7840 , n7841 , n7842 , n7843 , 
n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , 
n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , 
n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , 
n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , 
n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , 
n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , 
n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , 
n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , 
n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , 
n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , 
n7944 , n7945 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , 
n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , 
n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , 
n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , 
n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , 
n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , 
n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , 
n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , 
n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , 
n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , 
n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , 
n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , 
n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , 
n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , 
n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , 
n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , 
n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , 
n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , 
n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , 
n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , 
n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , 
n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , 
n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , 
n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , 
n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , 
n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , 
n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , 
n8215 , n8216 , n8217 , n8218 , n8219 , n8221 , n8222 , n8223 , n8224 , n8225 , 
n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , 
n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , 
n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , 
n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , 
n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , 
n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , 
n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , 
n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , 
n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , 
n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , 
n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , 
n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , 
n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , 
n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , 
n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , 
n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , 
n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , 
n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , 
n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , 
n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , 
n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , 
n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , 
n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , 
n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , 
n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , 
n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , 
n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8495 , n8496 , 
n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , 
n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , 
n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , 
n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , 
n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , 
n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , 
n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , 
n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , 
n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , 
n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , 
n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , 
n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , 
n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , 
n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , 
n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , 
n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , 
n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , 
n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , 
n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , 
n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , 
n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , 
n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , 
n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , 
n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , 
n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , 
n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , 
n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , 
n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , 
n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , 
n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , 
n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , 
n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , 
n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , 
n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , 
n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , 
n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , 
n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , 
n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , 
n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , 
n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , 
n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , 
n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , 
n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , 
n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , 
n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , 
n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , 
n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , 
n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , 
n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , 
n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , 
n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , 
n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , 
n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , 
n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , 
n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , 
n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , 
n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , 
n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , 
n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , 
n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , 
n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , 
n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , 
n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , 
n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , 
n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9145 , n9146 , n9148 , n9149 , 
n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , 
n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , 
n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9178 , n9179 , n9180 , 
n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , 
n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , 
n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , 
n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , 
n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , 
n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , 
n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , 
n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , 
n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , 
n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , 
n9281 , n9282 , n9283 , n9284 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , 
n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , 
n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9310 , n9311 , n9312 , 
n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , 
n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , 
n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , 
n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , 
n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , 
n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , 
n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , 
n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , 
n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , 
n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , 
n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , 
n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , 
n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , 
n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , 
n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , 
n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , 
n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , 
n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , 
n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , 
n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , 
n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , 
n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , 
n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , 
n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , 
n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , 
n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , 
n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , 
n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , 
n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , 
n9603 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , 
n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , 
n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , 
n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9642 , n9643 , n9644 , 
n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , 
n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , 
n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , 
n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , 
n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , 
n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , 
n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , 
n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , 
n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , 
n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , 
n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , 
n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , 
n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , 
n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , 
n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , 
n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , 
n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , 
n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , 
n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , 
n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , 
n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , 
n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , 
n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , 
n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , 
n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , 
n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , 
n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , 
n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , 
n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , 
n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , 
n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , 
n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , 
n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , 
n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , 
n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , 
n9995 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , 
n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , 
n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , 
n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , 
n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , 
n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , 
n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , 
n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , 
n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , 
n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , 
n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , 
n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , 
n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , 
n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , 
n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , 
n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , 
n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , 
n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , 
n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , 
n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , 
n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , 
n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , 
n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , 
n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , 
n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , 
n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , 
n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , 
n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , 
n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , 
n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , 
n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , 
n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , 
n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , 
n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , 
n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , 
n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , 
n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , 
n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , 
n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , 
n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , 
n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , 
n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , 
n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , 
n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , 
n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , 
n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , 
n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , 
n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , 
n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , 
n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , 
n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , 
n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , 
n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , 
n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , 
n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , 
n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , 
n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , 
n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , 
n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , 
n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , 
n10597 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , 
n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , 
n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10626 , n10627 , n10628 , 
n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , 
n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , 
n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , 
n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , 
n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , 
n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , 
n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , 
n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , 
n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , 
n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , 
n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , 
n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , 
n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , 
n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , 
n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , 
n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , 
n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , 
n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , 
n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , 
n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , 
n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , 
n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , 
n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , 
n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , 
n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , 
n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , 
n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , 
n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , 
n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , 
n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , 
n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , 
n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , 
n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , 
n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , 
n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , 
n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , 
n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , 
n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , 
n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , 
n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , 
n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , 
n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , 
n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , 
n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , 
n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , 
n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , 
n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , 
n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , 
n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , 
n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , 
n11129 , n11130 , n11131 , n11132 , n11133 , n11135 , n11136 , n11137 , n11138 , n11139 , 
n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , 
n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , 
n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , 
n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , 
n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , 
n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , 
n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , 
n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , 
n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , 
n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , 
n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , 
n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , 
n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , 
n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , 
n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , 
n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11298 , n11299 , n11300 , 
n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , 
n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , 
n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , 
n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , 
n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , 
n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , 
n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , 
n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , 
n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , 
n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , 
n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , 
n11411 , n11412 , n11413 , n11414 , n11415 , n11417 , n11418 , n11419 , n11420 , n11421 , 
n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , 
n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , 
n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , 
n11452 , n11453 , n11454 , n11455 , n11456 , n11458 , n11459 , n11460 , n11461 , n11462 , 
n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , 
n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , 
n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , 
n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , 
n11503 , n11504 , n11505 , n11506 , n11507 , n11509 , n11510 , n11511 , n11512 , n11513 , 
n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , 
n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , 
n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , 
n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , 
n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , 
n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , 
n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , 
n11584 , n11585 , n11586 , n11587 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , 
n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , 
n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , 
n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , 
n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , 
n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , 
n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , 
n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , 
n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , 
n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , 
n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , 
n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , 
n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , 
n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , 
n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , 
n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , 
n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , 
n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , 
n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , 
n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , 
n11785 , n11786 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , 
n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , 
n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , 
n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , 
n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , 
n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , 
n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , 
n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , 
n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , 
n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , 
n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , 
n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , 
n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , 
n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , 
n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , 
n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , 
n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , 
n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , 
n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , 
n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , 
n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , 
n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , 
n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , 
n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , 
n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , 
n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , 
n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , 
n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , 
n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , 
n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , 
n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , 
n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , 
n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , 
n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , 
n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12134 , n12135 , n12136 , 
n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , 
n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , 
n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , 
n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , 
n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , 
n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , 
n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , 
n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , 
n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , 
n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , 
n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , 
n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , 
n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , 
n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , 
n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , 
n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , 
n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , 
n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , 
n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , 
n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , 
n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , 
n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , 
n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , 
n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , 
n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , 
n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , 
n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , 
n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , 
n12417 , n12418 , n12419 , n12420 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , 
n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , 
n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , 
n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , 
n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , 
n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , 
n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , 
n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , 
n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , 
n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , 
n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , 
n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , 
n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , 
n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , 
n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , 
n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , 
n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , 
n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , 
n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , 
n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , 
n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , 
n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , 
n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , 
n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , 
n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , 
n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , 
n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , 
n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , 
n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , 
n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , 
n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12726 , n12727 , n12728 , 
n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , 
n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , 
n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , 
n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , 
n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , 
n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , 
n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , 
n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , 
n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , 
n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , 
n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , 
n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , 
n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , 
n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , 
n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , 
n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , 
n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , 
n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , 
n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , 
n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , 
n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , 
n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , 
n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , 
n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , 
n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , 
n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , 
n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , 
n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , 
n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , 
n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , 
n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , 
n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , 
n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , 
n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , 
n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , 
n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , 
n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , 
n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , 
n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , 
n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , 
n13129 , n13130 , n13131 , n13132 , n13133 , n13135 , n13136 , n13137 , n13138 , n13139 , 
n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , 
n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , 
n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , 
n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , 
n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , 
n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , 
n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , 
n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , 
n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , 
n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , 
n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , 
n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , 
n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , 
n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , 
n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , 
n13290 , n13291 , n13292 , n13293 , n13294 , n13296 , n13297 , n13298 , n13299 , n13300 , 
n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , 
n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , 
n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , 
n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , 
n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , 
n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , 
n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , 
n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , 
n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , 
n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , 
n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , 
n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , 
n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , 
n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , 
n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , 
n13451 , n13452 , n13453 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , 
n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , 
n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , 
n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , 
n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , 
n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , 
n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , 
n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , 
n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , 
n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , 
n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , 
n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , 
n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , 
n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , 
n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , 
n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , 
n13612 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , 
n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , 
n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , 
n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , 
n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , 
n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , 
n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , 
n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , 
n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , 
n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , 
n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , 
n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , 
n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , 
n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , 
n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , 
n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , 
n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , 
n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , 
n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , 
n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , 
n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13821 , n13822 , n13823 , 
n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , 
n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , 
n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , 
n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , 
n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , 
n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , 
n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , 
n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , 
n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , 
n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , 
n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , 
n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , 
n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , 
n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , 
n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , 
n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , 
n13984 , n13985 , n13986 , n13987 , n13988 , n13990 , n13991 , n13992 , n13993 , n13994 , 
n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , 
n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , 
n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , 
n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , 
n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14043 , n14044 , n14045 , 
n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , 
n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , 
n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , 
n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , 
n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , 
n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , 
n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , 
n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , 
n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , 
n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , 
n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , 
n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , 
n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , 
n14176 , n14177 , n14178 , n14179 , n14181 , n14182 , n14183 , n14184 , n14185 , n14187 , 
n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , 
n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , 
n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , 
n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , 
n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , 
n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , 
n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , 
n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , 
n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , 
n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , 
n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , 
n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , 
n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , 
n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , 
n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , 
n14339 , n14340 , n14341 , n14342 , n14343 , n14345 , n14346 , n14347 , n14348 , n14349 , 
n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , 
n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , 
n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , 
n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , 
n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , 
n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , 
n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , 
n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , 
n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , 
n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , 
n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , 
n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , 
n14470 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , 
n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , 
n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , 
n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , 
n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , 
n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , 
n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , 
n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , 
n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , 
n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , 
n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , 
n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , 
n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , 
n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , 
n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , 
n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , 
n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , 
n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , 
n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , 
n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , 
n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , 
n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , 
n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , 
n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14708 , n14709 , n14710 , n14711 , 
n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , 
n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , 
n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , 
n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , 
n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , 
n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , 
n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , 
n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , 
n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , 
n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , 
n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , 
n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , 
n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , 
n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , 
n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , 
n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , 
n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , 
n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , 
n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , 
n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , 
n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , 
n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , 
n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , 
n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , 
n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , 
n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , 
n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , 
n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , 
n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , 
n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , 
n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , 
n15022 , n15023 , n15024 , n15025 , n15026 , n15028 , n15029 , n15030 , n15031 , n15032 , 
n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , 
n15043 , n15044 , n15045 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , 
n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , 
n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15071 , n15072 , n15073 , n15074 , 
n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , 
n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , 
n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , 
n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , 
n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , 
n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , 
n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , 
n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , 
n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , 
n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , 
n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , 
n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , 
n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , 
n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , 
n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , 
n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , 
n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , 
n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , 
n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , 
n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , 
n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , 
n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , 
n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , 
n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , 
n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , 
n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , 
n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , 
n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , 
n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , 
n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , 
n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , 
n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , 
n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , 
n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , 
n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , 
n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , 
n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , 
n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , 
n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , 
n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , 
n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , 
n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , 
n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , 
n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , 
n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , 
n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , 
n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , 
n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , 
n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , 
n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , 
n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , 
n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , 
n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , 
n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , 
n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , 
n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , 
n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , 
n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , 
n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , 
n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , 
n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , 
n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , 
n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , 
n15705 , n15706 , n15707 , n15708 , n15709 , n15711 , n15712 , n15713 , n15714 , n15715 , 
n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , 
n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , 
n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , 
n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , 
n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , 
n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , 
n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , 
n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , 
n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , 
n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , 
n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , 
n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , 
n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , 
n15846 , n15847 , n15848 , n15849 , n15850 , n15852 , n15853 , n15854 , n15855 , n15856 , 
n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , 
n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , 
n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , 
n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , 
n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , 
n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , 
n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , 
n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , 
n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , 
n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , 
n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , 
n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , 
n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , 
n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , 
n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , 
n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , 
n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , 
n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , 
n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , 
n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , 
n16057 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , 
n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , 
n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , 
n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , 
n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , 
n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , 
n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , 
n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , 
n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , 
n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , 
n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , 
n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , 
n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , 
n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , 
n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , 
n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , 
n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , 
n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , 
n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , 
n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , 
n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , 
n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , 
n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , 
n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , 
n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , 
n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , 
n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , 
n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , 
n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , 
n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , 
n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , 
n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , 
n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , 
n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , 
n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , 
n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , 
n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , 
n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , 
n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , 
n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , 
n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , 
n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , 
n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , 
n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , 
n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , 
n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , 
n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , 
n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , 
n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , 
n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , 
n16558 , n16559 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , 
n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , 
n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , 
n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16599 , 
n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , 
n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , 
n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , 
n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , 
n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , 
n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , 
n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , 
n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , 
n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , 
n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , 
n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , 
n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , 
n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , 
n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , 
n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , 
n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , 
n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , 
n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , 
n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , 
n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , 
n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , 
n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , 
n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , 
n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , 
n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , 
n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , 
n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , 
n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , 
n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , 
n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , 
n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , 
n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , 
n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , 
n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , 
n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , 
n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , 
n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , 
n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , 
n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , 
n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n17000 , n17001 , 
n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , 
n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , 
n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , 
n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , 
n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , 
n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , 
n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , 
n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , 
n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , 
n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , 
n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , 
n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17121 , n17122 , 
n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , 
n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , 
n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , 
n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , 
n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , 
n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , 
n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , 
n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , 
n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , 
n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , 
n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , 
n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , 
n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , 
n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , 
n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , 
n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , 
n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , 
n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , 
n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , 
n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , 
n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , 
n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , 
n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , 
n17354 , n17355 , n17356 , n17357 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , 
n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , 
n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , 
n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , 
n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , 
n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , 
n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17422 , n17423 , n17424 , n17425 , 
n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , 
n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , 
n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , 
n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , 
n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , 
n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , 
n17486 , n17487 , n17488 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , 
n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , 
n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17517 , 
n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , 
n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , 
n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , 
n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , 
n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , 
n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , 
n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , 
n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , 
n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , 
n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , 
n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , 
n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , 
n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , 
n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , 
n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , 
n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , 
n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , 
n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , 
n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , 
n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , 
n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , 
n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , 
n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17745 , n17746 , n17747 , n17748 , 
n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , 
n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , 
n17769 , n17770 , n17771 , n17772 , n17773 , n17775 , n17777 , n17778 , n17779 , n17780 , 
n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , 
n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , 
n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , 
n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , 
n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , 
n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , 
n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , 
n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , 
n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , 
n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , 
n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , 
n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , 
n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , 
n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , 
n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , 
n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , 
n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , 
n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , 
n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , 
n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , 
n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , 
n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , 
n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , 
n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , 
n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , 
n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , 
n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , 
n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , 
n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , 
n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , 
n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , 
n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , 
n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , 
n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , 
n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , 
n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , 
n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , 
n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , 
n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , 
n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , 
n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , 
n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , 
n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , 
n18211 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , 
n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , 
n18232 , n18233 , n18234 , n18235 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , 
n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , 
n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , 
n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , 
n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , 
n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , 
n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , 
n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , 
n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , 
n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , 
n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , 
n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , 
n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , 
n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , 
n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , 
n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , 
n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , 
n18403 , n18404 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , 
n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , 
n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , 
n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , 
n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , 
n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , 
n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , 
n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , 
n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , 
n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , 
n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , 
n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , 
n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , 
n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , 
n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , 
n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , 
n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , 
n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , 
n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , 
n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , 
n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , 
n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , 
n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , 
n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , 
n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , 
n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , 
n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , 
n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18684 , 
n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , 
n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , 
n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , 
n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , 
n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , 
n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , 
n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , 
n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , 
n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , 
n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , 
n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , 
n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , 
n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , 
n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , 
n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , 
n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , 
n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , 
n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , 
n18865 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , 
n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , 
n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , 
n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , 
n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , 
n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , 
n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , 
n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , 
n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18954 , n18955 , n18956 , 
n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , 
n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , 
n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , 
n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , 
n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , 
n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , 
n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , 
n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , 
n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , 
n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , 
n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , 
n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , 
n19077 , n19078 , n19079 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , 
n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , 
n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , 
n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , 
n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , 
n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , 
n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , 
n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , 
n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , 
n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , 
n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , 
n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , 
n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , 
n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , 
n19218 , n19219 , n19220 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , 
n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , 
n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , 
n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , 
n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , 
n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , 
n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , 
n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , 
n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , 
n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , 
n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , 
n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , 
n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , 
n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , 
n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19368 , n19369 , 
n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , 
n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , 
n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , 
n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , 
n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , 
n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , 
n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , 
n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , 
n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , 
n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , 
n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , 
n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , 
n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , 
n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , 
n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , 
n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , 
n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , 
n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , 
n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , 
n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , 
n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , 
n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , 
n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , 
n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , 
n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , 
n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , 
n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , 
n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , 
n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , 
n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , 
n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , 
n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , 
n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , 
n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , 
n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , 
n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , 
n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , 
n19741 , n19742 , n19743 , n19745 , n19746 , n19748 , n19749 , n19750 , n19751 , n19752 , 
n19753 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , 
n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , 
n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , 
n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , 
n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , 
n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , 
n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , 
n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , 
n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , 
n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , 
n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , 
n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , 
n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , 
n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , 
n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , 
n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , 
n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , 
n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , 
n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , 
n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , 
n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , 
n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , 
n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , 
n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , 
n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , 
n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , 
n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , 
n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , 
n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , 
n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , 
n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , 
n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , 
n20074 , n20075 , n20076 , n20077 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , 
n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , 
n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , 
n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , 
n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , 
n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , 
n20135 , n20136 , n20137 , n20138 , n20139 , n20141 , n20142 , n20143 , n20144 , n20145 , 
n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , 
n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , 
n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , 
n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , 
n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , 
n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , 
n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , 
n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , 
n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , 
n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , 
n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , 
n20256 , n20257 , n20258 , n20259 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , 
n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , 
n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , 
n20287 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , 
n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , 
n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , 
n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , 
n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , 
n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , 
n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , 
n20358 , n20359 , n20360 , n20361 , n20362 , n20364 , n20365 , n20366 , n20367 , n20368 , 
n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , 
n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , 
n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , 
n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , 
n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , 
n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , 
n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , 
n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , 
n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , 
n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , 
n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , 
n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , 
n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , 
n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , 
n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , 
n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , 
n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , 
n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , 
n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , 
n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , 
n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , 
n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , 
n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , 
n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , 
n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , 
n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , 
n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , 
n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , 
n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , 
n20659 , n20660 , n20661 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , 
n20670 , n20671 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , 
n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , 
n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , 
n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , 
n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , 
n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , 
n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , 
n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , 
n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , 
n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , 
n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , 
n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , 
n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , 
n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , 
n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , 
n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , 
n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , 
n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , 
n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , 
n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , 
n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , 
n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , 
n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , 
n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , 
n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , 
n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , 
n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , 
n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20950 , n20951 , n20952 , 
n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , 
n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , 
n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , 
n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , 
n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , 
n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , 
n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , 
n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , 
n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , 
n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , 
n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , 
n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , 
n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , 
n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , 
n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , 
n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , 
n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , 
n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , 
n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , 
n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , 
n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , 
n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , 
n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , 
n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , 
n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , 
n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , 
n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , 
n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , 
n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , 
n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , 
n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , 
n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , 
n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , 
n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , 
n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , 
n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , 
n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , 
n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , 
n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , 
n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , 
n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , 
n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , 
n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , 
n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , 
n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , 
n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , 
n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , 
n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , 
n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , 
n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , 
n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , 
n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , 
n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , 
n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , 
n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , 
n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , 
n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , 
n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , 
n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , 
n21543 , n21544 , n21545 , n21546 , n21547 , n21549 , n21550 , n21551 , n21552 , n21553 , 
n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , 
n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , 
n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , 
n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , 
n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , 
n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , 
n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , 
n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , 
n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , 
n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , 
n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , 
n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , 
n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , 
n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , 
n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21704 , 
n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , 
n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , 
n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , 
n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , 
n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , 
n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , 
n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , 
n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , 
n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , 
n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , 
n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , 
n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , 
n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , 
n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , 
n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , 
n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , 
n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , 
n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , 
n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , 
n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , 
n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , 
n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , 
n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , 
n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , 
n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , 
n21955 , n21956 , n21957 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , 
n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , 
n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , 
n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , 
n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , 
n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , 
n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , 
n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , 
n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , 
n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , 
n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , 
n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , 
n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , 
n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , 
n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , 
n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , 
n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , 
n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , 
n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , 
n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , 
n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , 
n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , 
n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , 
n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , 
n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , 
n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , 
n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , 
n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , 
n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , 
n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , 
n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , 
n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , 
n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , 
n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , 
n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , 
n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , 
n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , 
n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , 
n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , 
n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , 
n22356 , n22357 , n22358 , n22359 , n22360 , n22362 , n22363 , n22364 , n22365 , n22366 , 
n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , 
n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , 
n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , 
n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , 
n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , 
n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , 
n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , 
n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , 
n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , 
n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , 
n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , 
n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , 
n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , 
n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , 
n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , 
n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , 
n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , 
n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , 
n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , 
n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , 
n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , 
n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , 
n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , 
n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , 
n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , 
n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , 
n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , 
n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , 
n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , 
n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , 
n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , 
n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , 
n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , 
n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , 
n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , 
n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , 
n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , 
n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , 
n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , 
n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , 
n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , 
n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , 
n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , 
n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , 
n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , 
n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , 
n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , 
n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , 
n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , 
n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , 
n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , 
n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , 
n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , 
n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , 
n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , 
n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , 
n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , 
n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , 
n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , 
n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , 
n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , 
n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , 
n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , 
n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , 
n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , 
n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , 
n23028 , n23029 , n23030 , n23031 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , 
n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , 
n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , 
n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , 
n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , 
n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , 
n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , 
n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , 
n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , 
n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , 
n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , 
n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , 
n23149 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , 
n23160 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , 
n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , 
n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , 
n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , 
n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , 
n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , 
n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , 
n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , 
n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , 
n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , 
n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , 
n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , 
n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , 
n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , 
n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , 
n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , 
n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , 
n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , 
n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , 
n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , 
n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , 
n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , 
n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , 
n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , 
n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , 
n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , 
n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , 
n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , 
n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , 
n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , 
n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , 
n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , 
n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , 
n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , 
n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , 
n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , 
n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , 
n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , 
n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , 
n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , 
n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , 
n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , 
n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , 
n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , 
n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , 
n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , 
n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , 
n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , 
n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , 
n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , 
n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , 
n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , 
n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , 
n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , 
n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , 
n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , 
n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , 
n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , 
n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , 
n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , 
n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , 
n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , 
n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , 
n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , 
n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , 
n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , 
n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , 
n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , 
n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , 
n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , 
n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , 
n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23881 , n23882 , 
n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , 
n23893 , n23894 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , 
n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , 
n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , 
n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , 
n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , 
n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , 
n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , 
n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , 
n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23982 , n23983 , n23984 , 
n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , 
n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , 
n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , 
n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , 
n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , 
n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , 
n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , 
n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , 
n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , 
n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , 
n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , 
n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , 
n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , 
n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , 
n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , 
n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , 
n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , 
n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , 
n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , 
n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , 
n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , 
n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , 
n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , 
n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , 
n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , 
n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , 
n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , 
n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , 
n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , 
n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , 
n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , 
n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , 
n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , 
n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , 
n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , 
n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , 
n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , 
n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , 
n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , 
n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , 
n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , 
n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , 
n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , 
n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , 
n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , 
n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , 
n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , 
n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , 
n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , 
n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , 
n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , 
n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , 
n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , 
n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , 
n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , 
n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , 
n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , 
n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , 
n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , 
n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , 
n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , 
n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , 
n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , 
n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24623 , n24624 , n24625 , 
n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , 
n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , 
n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , 
n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , 
n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , 
n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , 
n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , 
n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , 
n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , 
n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , 
n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , 
n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , 
n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , 
n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , 
n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , 
n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , 
n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , 
n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , 
n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , 
n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , 
n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , 
n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , 
n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , 
n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , 
n24867 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , 
n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , 
n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , 
n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , 
n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , 
n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , 
n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , 
n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , 
n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , 
n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , 
n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , 
n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , 
n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , 
n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , 
n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , 
n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , 
n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , 
n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , 
n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , 
n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , 
n25068 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , 
n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , 
n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , 
n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , 
n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , 
n25119 , n25120 , n25121 , n25122 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , 
n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , 
n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , 
n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , 
n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , 
n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , 
n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , 
n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , 
n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , 
n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , 
n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , 
n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , 
n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , 
n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , 
n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , 
n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , 
n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , 
n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , 
n25300 , n25301 , n25302 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , 
n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , 
n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , 
n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , 
n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , 
n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , 
n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , 
n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , 
n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , 
n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , 
n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25408 , n25409 , n25410 , n25411 , 
n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , 
n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , 
n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , 
n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , 
n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , 
n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , 
n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , 
n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , 
n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , 
n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , 
n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , 
n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , 
n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , 
n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25550 , n25551 , n25552 , 
n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , 
n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , 
n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , 
n25583 , n25584 , n25585 , n25586 , n25587 , n25589 , n25590 , n25591 , n25592 , n25593 , 
n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , 
n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , 
n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , 
n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , 
n25634 , n25635 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , 
n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , 
n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , 
n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , 
n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , 
n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , 
n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , 
n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , 
n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , 
n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , 
n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , 
n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , 
n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , 
n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , 
n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , 
n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , 
n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , 
n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , 
n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , 
n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , 
n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , 
n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , 
n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , 
n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , 
n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , 
n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , 
n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , 
n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , 
n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , 
n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , 
n25935 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , 
n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , 
n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , 
n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , 
n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , 
n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , 
n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , 
n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , 
n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , 
n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , 
n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , 
n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , 
n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , 
n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , 
n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , 
n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , 
n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , 
n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , 
n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , 
n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , 
n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , 
n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , 
n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , 
n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , 
n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , 
n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , 
n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , 
n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , 
n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , 
n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , 
n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , 
n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , 
n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , 
n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , 
n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , 
n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , 
n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , 
n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , 
n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , 
n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , 
n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , 
n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , 
n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , 
n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , 
n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , 
n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , 
n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , 
n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , 
n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , 
n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , 
n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , 
n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , 
n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , 
n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , 
n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , 
n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , 
n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , 
n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , 
n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , 
n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , 
n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , 
n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , 
n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , 
n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , 
n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , 
n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , 
n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , 
n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , 
n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , 
n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , 
n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , 
n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , 
n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , 
n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , 
n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , 
n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , 
n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , 
n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , 
n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , 
n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , 
n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , 
n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , 
n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , 
n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , 
n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , 
n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , 
n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , 
n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , 
n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , 
n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , 
n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , 
n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , 
n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , 
n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , 
n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , 
n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , 
n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , 
n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , 
n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , 
n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , 
n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , 
n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , 
n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , 
n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , 
n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , 
n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , 
n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , 
n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , 
n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , 
n27026 , n27027 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , 
n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , 
n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , 
n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , 
n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , 
n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , 
n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , 
n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , 
n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , 
n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , 
n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , 
n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , 
n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , 
n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , 
n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , 
n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , 
n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , 
n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , 
n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , 
n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , 
n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , 
n27237 , n27238 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , 
n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , 
n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , 
n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , 
n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , 
n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , 
n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , 
n27309 , n27310 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , 
n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , 
n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , 
n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , 
n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , 
n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , 
n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , 
n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , 
n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , 
n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , 
n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , 
n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , 
n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , 
n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , 
n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , 
n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , 
n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , 
n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , 
n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , 
n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , 
n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , 
n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , 
n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , 
n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , 
n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , 
n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , 
n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , 
n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , 
n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , 
n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , 
n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , 
n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , 
n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , 
n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , 
n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , 
n27661 , n27662 , n27664 , n27665 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , 
n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , 
n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , 
n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , 
n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , 
n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , 
n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , 
n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , 
n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , 
n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , 
n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , 
n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , 
n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , 
n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , 
n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , 
n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , 
n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , 
n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , 
n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , 
n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , 
n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , 
n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , 
n27883 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27893 , n27894 , 
n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , 
n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , 
n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , 
n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , 
n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27943 , n27944 , n27945 , 
n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , 
n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , 
n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , 
n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , 
n27986 , n27987 , n27988 , n27989 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , 
n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , 
n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , 
n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , 
n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , 
n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , 
n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , 
n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28065 , n28066 , n28067 , 
n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , 
n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , 
n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , 
n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , 
n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , 
n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , 
n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , 
n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , 
n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , 
n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , 
n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , 
n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , 
n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , 
n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , 
n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , 
n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , 
n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , 
n28238 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , 
n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , 
n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , 
n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , 
n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , 
n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , 
n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , 
n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , 
n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , 
n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , 
n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , 
n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , 
n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , 
n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , 
n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , 
n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , 
n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , 
n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , 
n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , 
n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , 
n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , 
n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , 
n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , 
n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , 
n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , 
n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , 
n28499 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , 
n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28519 , n28520 , 
n28521 , n28522 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , 
n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , 
n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , 
n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , 
n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , 
n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , 
n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , 
n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , 
n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , 
n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , 
n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , 
n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , 
n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , 
n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , 
n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , 
n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , 
n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , 
n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , 
n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , 
n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , 
n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , 
n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , 
n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , 
n28752 , n28753 , n28754 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , 
n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , 
n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , 
n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , 
n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , 
n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , 
n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , 
n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , 
n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , 
n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , 
n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , 
n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , 
n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , 
n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , 
n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , 
n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , 
n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , 
n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , 
n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , 
n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , 
n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , 
n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , 
n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , 
n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , 
n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , 
n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , 
n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , 
n29023 , n29024 , n29025 , n29026 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , 
n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , 
n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , 
n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , 
n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , 
n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , 
n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , 
n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , 
n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , 
n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , 
n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , 
n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , 
n29144 , n29145 , n29146 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , 
n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , 
n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , 
n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , 
n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , 
n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , 
n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29215 , 
n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , 
n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , 
n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , 
n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , 
n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , 
n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , 
n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , 
n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , 
n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , 
n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , 
n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , 
n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , 
n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , 
n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , 
n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , 
n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , 
n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , 
n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , 
n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , 
n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , 
n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , 
n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , 
n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , 
n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , 
n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , 
n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , 
n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , 
n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , 
n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , 
n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , 
n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , 
n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , 
n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , 
n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , 
n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , 
n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , 
n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , 
n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , 
n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , 
n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , 
n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , 
n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , 
n29636 , n29637 , n29638 , n29639 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , 
n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , 
n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , 
n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , 
n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , 
n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , 
n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , 
n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , 
n29717 , n29718 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , 
n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , 
n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , 
n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , 
n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , 
n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , 
n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , 
n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , 
n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , 
n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29817 , n29818 , n29819 , 
n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , 
n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , 
n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , 
n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , 
n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , 
n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , 
n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , 
n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , 
n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , 
n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , 
n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , 
n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , 
n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , 
n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , 
n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , 
n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , 
n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , 
n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , 
n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , 
n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , 
n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , 
n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , 
n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , 
n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , 
n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , 
n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , 
n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , 
n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , 
n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , 
n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , 
n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , 
n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , 
n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , 
n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , 
n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , 
n30172 , n30173 , n30174 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , 
n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , 
n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , 
n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , 
n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , 
n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , 
n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , 
n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , 
n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , 
n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , 
n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , 
n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , 
n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , 
n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , 
n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , 
n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , 
n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , 
n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , 
n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , 
n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , 
n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , 
n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , 
n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , 
n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , 
n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , 
n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , 
n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , 
n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , 
n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , 
n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , 
n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , 
n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , 
n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , 
n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , 
n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , 
n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , 
n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , 
n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , 
n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , 
n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , 
n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , 
n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , 
n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , 
n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , 
n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , 
n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , 
n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , 
n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , 
n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , 
n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , 
n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , 
n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , 
n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , 
n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , 
n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , 
n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , 
n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , 
n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , 
n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , 
n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , 
n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , 
n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , 
n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , 
n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , 
n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , 
n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , 
n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , 
n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , 
n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , 
n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , 
n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , 
n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30893 , 
n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , 
n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , 
n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , 
n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , 
n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , 
n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , 
n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , 
n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , 
n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , 
n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , 
n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , 
n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , 
n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , 
n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , 
n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , 
n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , 
n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , 
n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , 
n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , 
n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , 
n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , 
n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , 
n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , 
n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , 
n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , 
n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , 
n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , 
n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , 
n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , 
n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , 
n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , 
n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , 
n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31223 , n31224 , 
n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , 
n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31242 , n31243 , n31244 , n31245 , 
n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , 
n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31264 , n31265 , n31266 , 
n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , 
n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , 
n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , 
n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , 
n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , 
n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , 
n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , 
n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , 
n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , 
n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , 
n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , 
n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , 
n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , 
n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , 
n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , 
n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , 
n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , 
n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , 
n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , 
n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , 
n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , 
n31477 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , 
n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , 
n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , 
n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , 
n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , 
n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , 
n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , 
n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , 
n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , 
n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , 
n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , 
n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , 
n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , 
n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , 
n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , 
n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , 
n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , 
n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , 
n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , 
n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , 
n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , 
n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , 
n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , 
n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , 
n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , 
n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , 
n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , 
n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , 
n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , 
n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , 
n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , 
n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , 
n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , 
n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , 
n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31828 , 
n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , 
n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , 
n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , 
n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , 
n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , 
n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , 
n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , 
n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , 
n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , 
n31919 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , 
n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , 
n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , 
n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , 
n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , 
n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , 
n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , 
n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , 
n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , 
n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , 
n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , 
n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , 
n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , 
n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , 
n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , 
n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , 
n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32089 , n32090 , 
n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , 
n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , 
n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , 
n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , 
n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , 
n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , 
n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , 
n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , 
n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , 
n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , 
n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , 
n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , 
n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , 
n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , 
n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , 
n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , 
n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , 
n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , 
n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32278 , n32279 , n32280 , n32281 , 
n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , 
n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , 
n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , 
n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , 
n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , 
n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , 
n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , 
n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , 
n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , 
n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , 
n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , 
n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , 
n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , 
n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , 
n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , 
n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , 
n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , 
n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , 
n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , 
n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , 
n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , 
n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , 
n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , 
n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , 
n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , 
n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , 
n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , 
n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , 
n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , 
n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , 
n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , 
n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , 
n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , 
n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , 
n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , 
n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , 
n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , 
n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , 
n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , 
n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , 
n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , 
n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32699 , n32700 , n32701 , n32702 , 
n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , 
n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , 
n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , 
n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , 
n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , 
n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , 
n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , 
n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , 
n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , 
n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , 
n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , 
n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , 
n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , 
n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , 
n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , 
n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , 
n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , 
n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , 
n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , 
n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , 
n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , 
n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , 
n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , 
n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , 
n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , 
n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , 
n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , 
n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , 
n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , 
n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , 
n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , 
n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , 
n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , 
n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , 
n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , 
n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , 
n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , 
n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , 
n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , 
n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , 
n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , 
n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , 
n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , 
n33133 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , 
n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , 
n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , 
n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , 
n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , 
n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , 
n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , 
n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , 
n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , 
n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , 
n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , 
n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , 
n33254 , n33255 , n33256 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , 
n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , 
n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , 
n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , 
n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , 
n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , 
n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , 
n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , 
n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , 
n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , 
n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , 
n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , 
n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , 
n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , 
n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , 
n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , 
n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , 
n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , 
n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , 
n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , 
n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , 
n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , 
n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , 
n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , 
n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , 
n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , 
n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , 
n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , 
n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , 
n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , 
n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , 
n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , 
n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , 
n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , 
n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , 
n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , 
n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , 
n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , 
n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , 
n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , 
n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , 
n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , 
n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , 
n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , 
n33695 , n33696 , n33697 , n33698 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , 
n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , 
n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , 
n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , 
n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , 
n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , 
n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , 
n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , 
n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , 
n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , 
n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , 
n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , 
n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , 
n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , 
n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , 
n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , 
n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , 
n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , 
n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , 
n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , 
n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , 
n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , 
n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , 
n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , 
n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , 
n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , 
n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , 
n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , 
n33976 , n33977 , n33978 , n33979 , n33980 , n33982 , n33983 , n33984 , n33985 , n33986 , 
n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , 
n33997 , n33998 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , 
n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , 
n34018 , n34019 , n34020 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , 
n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , 
n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , 
n34049 , n34050 , n34051 , n34052 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , 
n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , 
n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , 
n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , 
n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , 
n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , 
n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , 
n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , 
n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34137 , n34138 , n34139 , n34140 , 
n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , 
n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , 
n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , 
n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , 
n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , 
n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , 
n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , 
n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , 
n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , 
n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , 
n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , 
n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , 
n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34268 , n34269 , n34270 , n34271 , 
n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , 
n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , 
n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , 
n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , 
n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , 
n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , 
n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , 
n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , 
n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , 
n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , 
n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , 
n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , 
n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , 
n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , 
n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , 
n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , 
n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , 
n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , 
n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , 
n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , 
n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , 
n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , 
n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , 
n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , 
n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , 
n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , 
n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , 
n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , 
n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34562 , n34563 , 
n34564 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34574 , n34575 , 
n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , 
n34586 , n34587 , n34588 , n34589 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , 
n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , 
n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , 
n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , 
n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , 
n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , 
n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34654 , n34655 , n34656 , n34657 , 
n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , 
n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , 
n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34687 , n34688 , 
n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , 
n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , 
n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , 
n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , 
n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , 
n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , 
n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , 
n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , 
n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , 
n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34789 , 
n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , 
n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , 
n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , 
n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , 
n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , 
n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , 
n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , 
n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , 
n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , 
n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , 
n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , 
n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , 
n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , 
n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , 
n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , 
n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , 
n34950 , n34951 , n34952 , n34953 , n34954 , n34956 , n34957 , n34958 , n34959 , n34960 , 
n34961 , n34962 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , 
n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , 
n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , 
n34992 , n34993 , n34994 , n34995 , n34996 , n34998 , n34999 , n35000 , n35001 , n35002 , 
n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , 
n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , 
n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , 
n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , 
n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , 
n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , 
n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , 
n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , 
n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , 
n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , 
n35103 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , 
n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , 
n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , 
n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , 
n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , 
n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , 
n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , 
n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , 
n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , 
n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , 
n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , 
n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , 
n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , 
n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , 
n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , 
n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , 
n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , 
n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , 
n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , 
n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35302 , n35303 , n35304 , 
n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , 
n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , 
n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , 
n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , 
n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , 
n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , 
n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , 
n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , 
n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , 
n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , 
n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35412 , n35413 , n35414 , n35415 , 
n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , 
n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , 
n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , 
n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , 
n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , 
n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , 
n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , 
n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , 
n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , 
n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , 
n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , 
n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , 
n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , 
n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , 
n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , 
n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , 
n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , 
n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , 
n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , 
n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , 
n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , 
n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , 
n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , 
n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , 
n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , 
n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , 
n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , 
n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , 
n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , 
n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , 
n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , 
n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35733 , n35734 , n35735 , n35736 , 
n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , 
n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , 
n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , 
n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , 
n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , 
n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , 
n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , 
n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , 
n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , 
n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , 
n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , 
n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , 
n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , 
n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , 
n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , 
n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , 
n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , 
n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , 
n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , 
n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , 
n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , 
n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , 
n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , 
n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , 
n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , 
n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , 
n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , 
n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , 
n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , 
n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , 
n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , 
n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , 
n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , 
n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , 
n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , 
n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , 
n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , 
n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , 
n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , 
n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , 
n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , 
n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , 
n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , 
n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , 
n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , 
n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , 
n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , 
n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , 
n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , 
n36228 , n36229 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , 
n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , 
n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , 
n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , 
n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , 
n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , 
n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , 
n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , 
n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , 
n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , 
n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , 
n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , 
n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , 
n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , 
n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , 
n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , 
n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , 
n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , 
n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , 
n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , 
n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , 
n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , 
n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , 
n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , 
n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , 
n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , 
n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , 
n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , 
n36509 , n36510 , n36511 , n36512 , n36513 , n36515 , n36516 , n36517 , n36518 , n36519 , 
n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , 
n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , 
n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , 
n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , 
n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , 
n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , 
n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , 
n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , 
n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , 
n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , 
n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , 
n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , 
n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , 
n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , 
n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , 
n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , 
n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36688 , n36689 , n36690 , 
n36691 , n36692 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , 
n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , 
n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , 
n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , 
n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , 
n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , 
n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , 
n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , 
n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , 
n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , 
n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , 
n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , 
n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , 
n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , 
n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , 
n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , 
n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , 
n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , 
n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , 
n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , 
n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , 
n36902 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , 
n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , 
n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , 
n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , 
n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , 
n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , 
n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , 
n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , 
n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , 
n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , 
n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , 
n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , 
n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , 
n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , 
n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , 
n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , 
n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , 
n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , 
n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , 
n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , 
n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , 
n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , 
n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , 
n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , 
n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , 
n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , 
n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , 
n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , 
n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , 
n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , 
n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , 
n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , 
n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , 
n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , 
n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , 
n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , 
n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , 
n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , 
n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , 
n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , 
n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , 
n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , 
n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , 
n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , 
n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , 
n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , 
n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , 
n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , 
n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , 
n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , 
n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , 
n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , 
n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , 
n37433 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , 
n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , 
n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , 
n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , 
n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , 
n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , 
n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , 
n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , 
n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , 
n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , 
n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , 
n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , 
n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , 
n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , 
n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , 
n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , 
n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , 
n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , 
n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , 
n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , 
n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , 
n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , 
n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , 
n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , 
n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , 
n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , 
n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , 
n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , 
n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , 
n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , 
n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , 
n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , 
n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , 
n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , 
n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , 
n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , 
n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , 
n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , 
n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , 
n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , 
n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , 
n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , 
n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , 
n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , 
n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , 
n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37891 , n37892 , n37893 , n37894 , 
n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , 
n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , 
n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , 
n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , 
n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , 
n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , 
n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , 
n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , 
n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , 
n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , 
n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , 
n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , 
n38015 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , 
n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , 
n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , 
n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , 
n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , 
n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , 
n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , 
n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , 
n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , 
n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , 
n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , 
n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , 
n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , 
n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , 
n38156 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , 
n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , 
n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , 
n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , 
n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , 
n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , 
n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , 
n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , 
n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , 
n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , 
n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , 
n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , 
n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , 
n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , 
n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , 
n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , 
n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , 
n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , 
n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , 
n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , 
n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , 
n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , 
n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , 
n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , 
n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , 
n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , 
n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , 
n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , 
n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , 
n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , 
n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , 
n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , 
n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , 
n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , 
n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , 
n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , 
n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38528 , 
n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , 
n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , 
n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , 
n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , 
n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , 
n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , 
n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , 
n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , 
n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , 
n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , 
n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , 
n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , 
n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , 
n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , 
n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , 
n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , 
n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , 
n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , 
n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , 
n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , 
n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , 
n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , 
n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , 
n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , 
n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , 
n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , 
n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , 
n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , 
n38809 , n38810 , n38811 , n38812 , n38814 , n38815 , n38816 , n38817 , n38818 , n38820 , 
n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , 
n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , 
n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , 
n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , 
n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , 
n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38880 , n38881 , 
n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , 
n38892 , n38893 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , 
n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , 
n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38921 , n38922 , n38923 , 
n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , 
n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , 
n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , 
n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , 
n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , 
n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , 
n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , 
n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , 
n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , 
n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , 
n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , 
n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , 
n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , 
n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , 
n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , 
n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , 
n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , 
n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , 
n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , 
n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , 
n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , 
n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , 
n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , 
n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , 
n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , 
n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , 
n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , 
n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , 
n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39214 , 
n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , 
n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , 
n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , 
n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , 
n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , 
n39265 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , 
n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , 
n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , 
n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , 
n39306 , n39307 , n39308 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , 
n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , 
n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , 
n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , 
n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , 
n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , 
n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , 
n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , 
n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , 
n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , 
n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , 
n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , 
n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , 
n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , 
n39447 , n39448 , n39449 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , 
n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , 
n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , 
n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , 
n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , 
n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , 
n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , 
n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , 
n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39537 , n39538 , 
n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , 
n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , 
n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , 
n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , 
n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , 
n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , 
n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , 
n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , 
n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , 
n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , 
n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , 
n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , 
n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , 
n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , 
n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , 
n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , 
n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , 
n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , 
n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , 
n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , 
n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , 
n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , 
n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , 
n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , 
n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , 
n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , 
n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , 
n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , 
n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , 
n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , 
n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , 
n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , 
n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , 
n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , 
n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , 
n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , 
n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , 
n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , 
n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , 
n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , 
n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , 
n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , 
n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , 
n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , 
n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , 
n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , 
n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , 
n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , 
n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , 
n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , 
n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , 
n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , 
n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , 
n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , 
n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , 
n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , 
n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , 
n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , 
n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , 
n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , 
n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , 
n40149 , n40150 , n40151 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , 
n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , 
n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , 
n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , 
n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , 
n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , 
n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , 
n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , 
n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , 
n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , 
n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , 
n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , 
n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , 
n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , 
n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , 
n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , 
n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , 
n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , 
n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , 
n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , 
n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , 
n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , 
n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , 
n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , 
n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , 
n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , 
n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , 
n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , 
n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , 
n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , 
n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , 
n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , 
n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , 
n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , 
n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , 
n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , 
n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , 
n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , 
n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , 
n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , 
n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40561 , 
n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , 
n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , 
n40582 , n40583 , n40584 , n40585 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , 
n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , 
n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , 
n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , 
n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , 
n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , 
n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , 
n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , 
n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , 
n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , 
n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , 
n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , 
n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , 
n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , 
n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , 
n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , 
n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , 
n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , 
n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , 
n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , 
n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , 
n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , 
n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , 
n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , 
n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , 
n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , 
n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , 
n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , 
n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , 
n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , 
n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , 
n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , 
n40903 , n40904 , n40905 , n40906 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , 
n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , 
n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , 
n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , 
n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , 
n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , 
n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , 
n40974 , n40975 , n40976 , n40977 , n40978 , n40980 , n40981 , n40982 , n40983 , n40984 , 
n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , 
n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , 
n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , 
n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , 
n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , 
n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , 
n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , 
n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , 
n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , 
n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , 
n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , 
n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , 
n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , 
n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , 
n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , 
n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , 
n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , 
n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , 
n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , 
n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , 
n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , 
n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , 
n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , 
n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , 
n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , 
n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , 
n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , 
n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , 
n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , 
n41275 , n41276 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , 
n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , 
n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , 
n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41316 , 
n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , 
n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , 
n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , 
n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , 
n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , 
n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , 
n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , 
n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , 
n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , 
n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , 
n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , 
n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , 
n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , 
n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , 
n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , 
n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , 
n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , 
n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , 
n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , 
n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , 
n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , 
n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41535 , n41536 , n41537 , n41538 , 
n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , 
n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , 
n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , 
n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , 
n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , 
n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , 
n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , 
n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , 
n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , 
n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , 
n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , 
n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , 
n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , 
n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , 
n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , 
n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , 
n41699 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , 
n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , 
n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , 
n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , 
n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , 
n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , 
n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41768 , n41769 , n41770 , 
n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , 
n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , 
n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , 
n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , 
n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , 
n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , 
n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , 
n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , 
n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , 
n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , 
n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , 
n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , 
n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , 
n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , 
n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , 
n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , 
n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , 
n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , 
n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , 
n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , 
n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , 
n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , 
n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , 
n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , 
n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , 
n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , 
n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , 
n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , 
n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , 
n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , 
n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , 
n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , 
n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , 
n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , 
n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , 
n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , 
n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , 
n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , 
n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , 
n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , 
n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , 
n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , 
n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , 
n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , 
n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , 
n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , 
n42231 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , 
n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42249 , n42250 , n42251 , n42252 , 
n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , 
n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , 
n42273 , n42274 , n42275 , n42276 , n42277 , n42279 , n42280 , n42281 , n42282 , n42283 , 
n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , 
n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , 
n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , 
n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , 
n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , 
n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , 
n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , 
n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , 
n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , 
n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , 
n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , 
n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , 
n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , 
n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , 
n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , 
n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , 
n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , 
n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , 
n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , 
n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , 
n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , 
n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , 
n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , 
n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42524 , 
n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , 
n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , 
n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , 
n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , 
n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , 
n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , 
n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , 
n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , 
n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , 
n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , 
n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , 
n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , 
n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , 
n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , 
n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , 
n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , 
n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , 
n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , 
n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , 
n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , 
n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , 
n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , 
n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , 
n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , 
n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , 
n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , 
n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , 
n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , 
n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , 
n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , 
n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , 
n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , 
n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , 
n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , 
n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , 
n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , 
n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , 
n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , 
n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , 
n42915 , n42916 , n42917 , n42918 ;
    and g0 ( n29522 , n36744 , n39284 );
    or g1 ( n40908 , n20893 , n1027 );
    or g2 ( n12450 , n6628 , n8053 );
    or g3 ( n24494 , n24480 , n4669 );
    or g4 ( n20307 , n18172 , n21670 );
    not g5 ( n29803 , n41253 );
    or g6 ( n1942 , n14707 , n28987 );
    or g7 ( n23969 , n2167 , n1223 );
    nor g8 ( n3863 , n34292 , n41823 );
    and g9 ( n40226 , n22229 , n6128 );
    nor g10 ( n40763 , n27344 , n7892 );
    nor g11 ( n39910 , n16620 , n13448 );
    or g12 ( n35596 , n8087 , n30380 );
    or g13 ( n21320 , n30237 , n31760 );
    or g14 ( n5716 , n40455 , n24017 );
    nor g15 ( n6791 , n1507 , n8143 );
    nor g16 ( n22562 , n17744 , n17388 );
    nor g17 ( n37177 , n2918 , n41041 );
    nor g18 ( n29848 , n15070 , n10155 );
    not g19 ( n13830 , n28843 );
    or g20 ( n17064 , n35466 , n27345 );
    not g21 ( n3955 , n37968 );
    and g22 ( n33776 , n20024 , n4690 );
    and g23 ( n28889 , n3296 , n1686 );
    or g24 ( n35775 , n41941 , n24340 );
    not g25 ( n21459 , n17722 );
    and g26 ( n1479 , n16323 , n20297 );
    nor g27 ( n11862 , n34049 , n6609 );
    not g28 ( n40861 , n34654 );
    xnor g29 ( n16419 , n10535 , n1300 );
    nor g30 ( n15737 , n36117 , n1948 );
    and g31 ( n38554 , n21756 , n20886 );
    or g32 ( n31667 , n10504 , n26453 );
    and g33 ( n8202 , n42674 , n6993 );
    or g34 ( n26678 , n28461 , n30976 );
    or g35 ( n6724 , n31318 , n40629 );
    and g36 ( n15578 , n23823 , n23410 );
    not g37 ( n21796 , n34957 );
    or g38 ( n42213 , n11092 , n20503 );
    or g39 ( n8866 , n14324 , n36461 );
    or g40 ( n42364 , n122 , n21494 );
    or g41 ( n30590 , n26226 , n8462 );
    or g42 ( n320 , n22440 , n4321 );
    and g43 ( n32200 , n26759 , n22952 );
    nor g44 ( n42134 , n18034 , n25380 );
    or g45 ( n997 , n6306 , n31671 );
    not g46 ( n40772 , n37760 );
    nor g47 ( n5791 , n26323 , n34282 );
    or g48 ( n4300 , n3660 , n31044 );
    not g49 ( n4746 , n28325 );
    xnor g50 ( n33430 , n37309 , n34849 );
    or g51 ( n3297 , n8494 , n10333 );
    or g52 ( n18361 , n11120 , n29939 );
    or g53 ( n23449 , n40670 , n15573 );
    and g54 ( n12061 , n11512 , n39833 );
    and g55 ( n7087 , n38287 , n24100 );
    or g56 ( n26754 , n5356 , n925 );
    not g57 ( n42642 , n40704 );
    xnor g58 ( n16257 , n7282 , n1972 );
    not g59 ( n38269 , n11525 );
    xnor g60 ( n34624 , n16143 , n41158 );
    not g61 ( n42166 , n23648 );
    not g62 ( n3109 , n7463 );
    nor g63 ( n36639 , n19856 , n38606 );
    xnor g64 ( n17884 , n31269 , n4525 );
    nor g65 ( n22529 , n7987 , n19066 );
    not g66 ( n9313 , n42257 );
    nor g67 ( n34365 , n26776 , n27954 );
    xnor g68 ( n3405 , n38789 , n29348 );
    or g69 ( n26483 , n2388 , n27962 );
    or g70 ( n29379 , n35712 , n12249 );
    or g71 ( n10231 , n9472 , n5850 );
    not g72 ( n29332 , n37653 );
    or g73 ( n20868 , n6273 , n20494 );
    and g74 ( n41877 , n41640 , n14771 );
    or g75 ( n10963 , n12947 , n32858 );
    nor g76 ( n32876 , n18866 , n26491 );
    xnor g77 ( n38332 , n20972 , n30386 );
    or g78 ( n17184 , n33981 , n20239 );
    or g79 ( n10054 , n4913 , n21558 );
    or g80 ( n5078 , n33134 , n15832 );
    nor g81 ( n37389 , n6179 , n1265 );
    not g82 ( n18921 , n36484 );
    not g83 ( n10527 , n9512 );
    or g84 ( n9036 , n23246 , n13495 );
    xnor g85 ( n3535 , n7717 , n25983 );
    or g86 ( n12678 , n19271 , n23610 );
    not g87 ( n18244 , n40141 );
    or g88 ( n29518 , n11976 , n482 );
    xnor g89 ( n21382 , n15591 , n25945 );
    and g90 ( n4611 , n20791 , n27460 );
    xnor g91 ( n17439 , n31956 , n36971 );
    not g92 ( n13586 , n38916 );
    not g93 ( n13979 , n41939 );
    and g94 ( n29300 , n42103 , n590 );
    or g95 ( n22738 , n41982 , n27485 );
    xnor g96 ( n210 , n2659 , n36198 );
    nor g97 ( n41397 , n32913 , n16204 );
    nor g98 ( n17416 , n5896 , n19163 );
    not g99 ( n34841 , n41945 );
    or g100 ( n3200 , n26927 , n8549 );
    or g101 ( n28215 , n37647 , n30779 );
    or g102 ( n16913 , n34505 , n3728 );
    or g103 ( n6287 , n37438 , n25541 );
    or g104 ( n12283 , n30600 , n32800 );
    or g105 ( n22682 , n5124 , n22104 );
    or g106 ( n6587 , n9135 , n15369 );
    and g107 ( n23848 , n11698 , n14799 );
    xnor g108 ( n30602 , n29185 , n9866 );
    and g109 ( n814 , n9458 , n21842 );
    or g110 ( n20368 , n23818 , n8710 );
    and g111 ( n31828 , n38707 , n34780 );
    or g112 ( n40172 , n39266 , n14726 );
    or g113 ( n20891 , n34358 , n19129 );
    and g114 ( n9462 , n22712 , n5346 );
    or g115 ( n23343 , n26927 , n39859 );
    or g116 ( n31732 , n37169 , n31860 );
    and g117 ( n9276 , n17112 , n20454 );
    or g118 ( n29830 , n4153 , n15236 );
    not g119 ( n15421 , n26817 );
    or g120 ( n995 , n42813 , n38481 );
    nor g121 ( n32959 , n29866 , n38700 );
    nor g122 ( n22455 , n1847 , n21076 );
    or g123 ( n13036 , n41205 , n30646 );
    and g124 ( n32521 , n26735 , n3058 );
    not g125 ( n20224 , n18915 );
    not g126 ( n15818 , n10025 );
    not g127 ( n34840 , n5496 );
    nor g128 ( n30304 , n5640 , n16888 );
    xnor g129 ( n37599 , n31436 , n38157 );
    and g130 ( n16809 , n25070 , n42091 );
    or g131 ( n10116 , n8646 , n30074 );
    or g132 ( n27181 , n29135 , n22898 );
    or g133 ( n27291 , n24203 , n5420 );
    or g134 ( n30765 , n14236 , n37950 );
    or g135 ( n17129 , n18611 , n39930 );
    and g136 ( n35478 , n14352 , n14841 );
    not g137 ( n30084 , n19658 );
    xnor g138 ( n24726 , n378 , n19446 );
    or g139 ( n18278 , n34941 , n42706 );
    nor g140 ( n34127 , n33981 , n23881 );
    or g141 ( n15668 , n8183 , n4449 );
    not g142 ( n40067 , n17441 );
    and g143 ( n16119 , n7325 , n21594 );
    or g144 ( n28000 , n3223 , n18712 );
    nor g145 ( n35660 , n4736 , n11413 );
    or g146 ( n4196 , n5605 , n4006 );
    not g147 ( n31421 , n19108 );
    xnor g148 ( n37823 , n18689 , n26956 );
    or g149 ( n33319 , n5910 , n28086 );
    xnor g150 ( n16263 , n41013 , n30090 );
    or g151 ( n11447 , n31286 , n4654 );
    and g152 ( n5677 , n10708 , n32641 );
    xnor g153 ( n13722 , n32178 , n12650 );
    not g154 ( n24665 , n30959 );
    or g155 ( n13738 , n8003 , n24371 );
    or g156 ( n41979 , n10284 , n7977 );
    or g157 ( n28136 , n6578 , n8362 );
    and g158 ( n31907 , n22366 , n20029 );
    and g159 ( n27819 , n38349 , n29642 );
    and g160 ( n39121 , n40009 , n39957 );
    not g161 ( n41047 , n2326 );
    or g162 ( n10509 , n36553 , n30780 );
    or g163 ( n4037 , n40349 , n24471 );
    or g164 ( n5734 , n42391 , n15541 );
    xnor g165 ( n36177 , n17430 , n270 );
    or g166 ( n16423 , n18865 , n9640 );
    and g167 ( n9341 , n12539 , n26506 );
    or g168 ( n26842 , n12286 , n11218 );
    nor g169 ( n25262 , n3769 , n27203 );
    or g170 ( n5776 , n29587 , n42132 );
    or g171 ( n16202 , n27517 , n20145 );
    nor g172 ( n17649 , n39266 , n9709 );
    or g173 ( n10015 , n23498 , n41981 );
    not g174 ( n39839 , n30555 );
    xnor g175 ( n39188 , n4094 , n8494 );
    or g176 ( n21827 , n15282 , n17940 );
    and g177 ( n14346 , n8879 , n28162 );
    and g178 ( n12128 , n1491 , n15168 );
    and g179 ( n37711 , n7072 , n38655 );
    and g180 ( n2016 , n23525 , n17699 );
    not g181 ( n31048 , n6984 );
    or g182 ( n32148 , n4131 , n22319 );
    xnor g183 ( n16904 , n29300 , n38157 );
    xnor g184 ( n5613 , n36009 , n35754 );
    and g185 ( n34448 , n2790 , n30695 );
    xnor g186 ( n1097 , n8250 , n31402 );
    nor g187 ( n13465 , n39025 , n24097 );
    and g188 ( n29314 , n24086 , n1222 );
    not g189 ( n18916 , n5947 );
    or g190 ( n7271 , n5279 , n24479 );
    or g191 ( n15024 , n29857 , n39731 );
    xnor g192 ( n23861 , n41013 , n8363 );
    not g193 ( n10434 , n27555 );
    or g194 ( n21406 , n16598 , n13416 );
    not g195 ( n18510 , n35158 );
    or g196 ( n28519 , n33964 , n39839 );
    xnor g197 ( n4287 , n15437 , n2440 );
    or g198 ( n19467 , n29542 , n29884 );
    not g199 ( n164 , n37193 );
    not g200 ( n4329 , n11081 );
    and g201 ( n4735 , n42685 , n37048 );
    and g202 ( n14368 , n7484 , n28902 );
    or g203 ( n35640 , n14945 , n6878 );
    and g204 ( n65 , n40546 , n16883 );
    not g205 ( n30622 , n2400 );
    or g206 ( n21849 , n30590 , n6826 );
    nor g207 ( n8373 , n29423 , n23005 );
    or g208 ( n15201 , n8374 , n10996 );
    xnor g209 ( n12378 , n10644 , n7277 );
    or g210 ( n1111 , n36186 , n33289 );
    or g211 ( n35442 , n36272 , n37361 );
    and g212 ( n38487 , n12148 , n12737 );
    not g213 ( n24505 , n402 );
    not g214 ( n36423 , n31626 );
    or g215 ( n38161 , n14057 , n21906 );
    and g216 ( n4145 , n38324 , n33165 );
    nor g217 ( n13839 , n21249 , n39824 );
    or g218 ( n10 , n20564 , n31021 );
    and g219 ( n12791 , n7638 , n7998 );
    nor g220 ( n4097 , n4601 , n37530 );
    nor g221 ( n20256 , n24045 , n38541 );
    not g222 ( n12836 , n14870 );
    or g223 ( n42210 , n27762 , n42058 );
    or g224 ( n4068 , n14450 , n39635 );
    not g225 ( n25751 , n23209 );
    not g226 ( n41545 , n13753 );
    xnor g227 ( n17631 , n20206 , n16139 );
    or g228 ( n14509 , n26808 , n14501 );
    not g229 ( n11832 , n36274 );
    or g230 ( n20318 , n28725 , n21446 );
    and g231 ( n40354 , n34126 , n30972 );
    and g232 ( n42351 , n27262 , n19231 );
    not g233 ( n17216 , n12934 );
    or g234 ( n29687 , n30174 , n8567 );
    not g235 ( n13997 , n42089 );
    and g236 ( n2124 , n3737 , n26315 );
    nor g237 ( n11258 , n13604 , n15746 );
    not g238 ( n38679 , n21998 );
    xnor g239 ( n23121 , n8924 , n14471 );
    or g240 ( n29164 , n35269 , n37411 );
    or g241 ( n37739 , n15384 , n13807 );
    xnor g242 ( n19203 , n35154 , n35571 );
    and g243 ( n23409 , n10224 , n15066 );
    or g244 ( n36054 , n9317 , n40305 );
    or g245 ( n29662 , n42575 , n29334 );
    or g246 ( n18653 , n36130 , n35382 );
    or g247 ( n6021 , n9462 , n7401 );
    or g248 ( n9257 , n2508 , n29203 );
    or g249 ( n30162 , n35033 , n15095 );
    xnor g250 ( n30579 , n23941 , n388 );
    and g251 ( n28441 , n29826 , n31176 );
    xnor g252 ( n27763 , n1216 , n28421 );
    or g253 ( n33783 , n10610 , n40956 );
    nor g254 ( n15071 , n29812 , n37924 );
    not g255 ( n6574 , n27425 );
    and g256 ( n32495 , n22327 , n12438 );
    xnor g257 ( n8976 , n40813 , n3043 );
    and g258 ( n29547 , n40026 , n18327 );
    nor g259 ( n16429 , n19211 , n35475 );
    or g260 ( n32096 , n33492 , n8460 );
    or g261 ( n14227 , n4043 , n4200 );
    or g262 ( n4472 , n16051 , n41359 );
    nor g263 ( n30893 , n33240 , n28350 );
    or g264 ( n35950 , n34772 , n20578 );
    and g265 ( n8997 , n25467 , n2691 );
    and g266 ( n17194 , n4840 , n38206 );
    xnor g267 ( n26898 , n39760 , n7869 );
    or g268 ( n34034 , n7947 , n32605 );
    or g269 ( n16355 , n24326 , n25451 );
    nor g270 ( n22734 , n22726 , n32691 );
    or g271 ( n36297 , n9141 , n32091 );
    or g272 ( n20104 , n398 , n2623 );
    and g273 ( n32545 , n39329 , n3272 );
    and g274 ( n16248 , n7641 , n34823 );
    or g275 ( n1298 , n27924 , n8143 );
    not g276 ( n25950 , n12253 );
    or g277 ( n28267 , n10460 , n28275 );
    or g278 ( n15627 , n16624 , n25142 );
    nor g279 ( n10051 , n24086 , n1222 );
    or g280 ( n37512 , n10496 , n17069 );
    and g281 ( n41516 , n12815 , n30562 );
    xnor g282 ( n35329 , n9900 , n30008 );
    and g283 ( n9941 , n7855 , n32960 );
    or g284 ( n19924 , n28484 , n25626 );
    not g285 ( n158 , n32807 );
    not g286 ( n25899 , n6402 );
    not g287 ( n10088 , n22954 );
    not g288 ( n6970 , n8706 );
    not g289 ( n21186 , n2957 );
    and g290 ( n4499 , n2550 , n42892 );
    or g291 ( n24091 , n41218 , n4202 );
    nor g292 ( n30402 , n16489 , n38006 );
    or g293 ( n14397 , n33981 , n37742 );
    xnor g294 ( n18939 , n38685 , n30232 );
    or g295 ( n14513 , n12180 , n24783 );
    and g296 ( n38401 , n37514 , n37958 );
    nor g297 ( n24848 , n8193 , n18418 );
    or g298 ( n21147 , n32481 , n17956 );
    xnor g299 ( n8717 , n3817 , n26841 );
    not g300 ( n22095 , n37991 );
    not g301 ( n28034 , n18728 );
    or g302 ( n21601 , n23621 , n12011 );
    or g303 ( n28852 , n20658 , n13958 );
    or g304 ( n14816 , n16052 , n26753 );
    or g305 ( n24890 , n25721 , n28363 );
    xnor g306 ( n25371 , n23706 , n16245 );
    or g307 ( n42581 , n33973 , n36198 );
    xnor g308 ( n38391 , n71 , n34475 );
    nor g309 ( n1247 , n25348 , n6521 );
    or g310 ( n12391 , n5910 , n42841 );
    or g311 ( n31401 , n40876 , n14738 );
    not g312 ( n6247 , n2513 );
    or g313 ( n29676 , n42893 , n39975 );
    or g314 ( n28618 , n7356 , n17464 );
    or g315 ( n3951 , n16907 , n17191 );
    and g316 ( n6446 , n33070 , n31152 );
    nor g317 ( n13520 , n11847 , n41438 );
    not g318 ( n11677 , n21183 );
    xnor g319 ( n20987 , n26579 , n6570 );
    or g320 ( n3293 , n739 , n31890 );
    or g321 ( n3547 , n17970 , n5185 );
    or g322 ( n16716 , n11575 , n7883 );
    not g323 ( n14490 , n28667 );
    and g324 ( n25040 , n40771 , n22995 );
    xnor g325 ( n37789 , n6371 , n14471 );
    and g326 ( n41373 , n11966 , n5486 );
    not g327 ( n36387 , n1088 );
    nor g328 ( n5308 , n28502 , n24215 );
    xnor g329 ( n34887 , n6625 , n23933 );
    or g330 ( n36985 , n10926 , n37106 );
    and g331 ( n35109 , n26831 , n9585 );
    xnor g332 ( n33302 , n8694 , n17407 );
    or g333 ( n27844 , n9135 , n24515 );
    or g334 ( n7627 , n22649 , n37721 );
    not g335 ( n8534 , n15509 );
    or g336 ( n36421 , n228 , n9299 );
    or g337 ( n6465 , n3848 , n14036 );
    or g338 ( n28095 , n29743 , n25234 );
    nor g339 ( n16229 , n14782 , n21498 );
    or g340 ( n10441 , n33203 , n25704 );
    nor g341 ( n14458 , n35597 , n29861 );
    or g342 ( n13156 , n18411 , n6221 );
    or g343 ( n3507 , n20145 , n7239 );
    and g344 ( n27274 , n30980 , n21862 );
    and g345 ( n12955 , n18995 , n9520 );
    not g346 ( n31033 , n31588 );
    not g347 ( n36890 , n17602 );
    and g348 ( n31807 , n27493 , n38385 );
    and g349 ( n24190 , n32788 , n40690 );
    xnor g350 ( n21937 , n42715 , n8146 );
    xnor g351 ( n33106 , n28987 , n14707 );
    or g352 ( n39797 , n23683 , n19096 );
    not g353 ( n2488 , n21246 );
    and g354 ( n27449 , n20623 , n17937 );
    or g355 ( n38536 , n42447 , n35398 );
    and g356 ( n7042 , n22636 , n11015 );
    or g357 ( n7133 , n28160 , n29211 );
    or g358 ( n20665 , n21361 , n30265 );
    or g359 ( n27990 , n41863 , n41520 );
    and g360 ( n35700 , n9362 , n24490 );
    or g361 ( n9933 , n538 , n29957 );
    or g362 ( n38382 , n34231 , n11961 );
    and g363 ( n12012 , n29561 , n31312 );
    not g364 ( n39813 , n39477 );
    and g365 ( n3238 , n41773 , n4568 );
    nor g366 ( n42906 , n37667 , n3094 );
    or g367 ( n26030 , n10146 , n42804 );
    not g368 ( n30336 , n7407 );
    or g369 ( n18048 , n29489 , n4792 );
    or g370 ( n3820 , n37868 , n19563 );
    or g371 ( n12356 , n27420 , n20675 );
    or g372 ( n37828 , n18314 , n36428 );
    not g373 ( n42553 , n6699 );
    or g374 ( n37441 , n12642 , n16534 );
    not g375 ( n27722 , n41992 );
    or g376 ( n26747 , n39699 , n2144 );
    or g377 ( n28868 , n34458 , n29298 );
    or g378 ( n8957 , n17482 , n7848 );
    xnor g379 ( n905 , n21476 , n25011 );
    or g380 ( n36617 , n10646 , n12449 );
    or g381 ( n15636 , n42859 , n40315 );
    and g382 ( n2224 , n31293 , n1434 );
    or g383 ( n15322 , n19523 , n37641 );
    and g384 ( n3790 , n17384 , n34627 );
    xnor g385 ( n24814 , n39432 , n23807 );
    and g386 ( n32091 , n1731 , n11717 );
    or g387 ( n22586 , n20031 , n30564 );
    nor g388 ( n9653 , n34292 , n11683 );
    or g389 ( n18820 , n24818 , n10936 );
    or g390 ( n37927 , n20988 , n28870 );
    or g391 ( n32654 , n9567 , n25504 );
    not g392 ( n12700 , n29949 );
    or g393 ( n36489 , n13059 , n734 );
    not g394 ( n42473 , n1171 );
    or g395 ( n14258 , n42099 , n32859 );
    or g396 ( n5521 , n192 , n26976 );
    not g397 ( n40358 , n12599 );
    or g398 ( n30718 , n5329 , n26111 );
    xnor g399 ( n31698 , n38371 , n27926 );
    and g400 ( n2234 , n42200 , n8258 );
    not g401 ( n25308 , n6809 );
    not g402 ( n7084 , n2329 );
    or g403 ( n1513 , n15750 , n36647 );
    not g404 ( n36798 , n14321 );
    not g405 ( n13205 , n24281 );
    not g406 ( n34267 , n4999 );
    xnor g407 ( n23873 , n26579 , n7203 );
    and g408 ( n37139 , n16894 , n9791 );
    nor g409 ( n19510 , n36117 , n20494 );
    or g410 ( n3843 , n16611 , n35797 );
    nor g411 ( n17941 , n16598 , n35818 );
    not g412 ( n23472 , n20393 );
    and g413 ( n9986 , n37979 , n39482 );
    nor g414 ( n31606 , n11784 , n34557 );
    not g415 ( n26352 , n18635 );
    or g416 ( n30215 , n30357 , n1082 );
    or g417 ( n19012 , n25271 , n19188 );
    nor g418 ( n42776 , n13604 , n5198 );
    or g419 ( n26811 , n35287 , n36621 );
    or g420 ( n28233 , n19185 , n14755 );
    and g421 ( n36718 , n36059 , n11430 );
    not g422 ( n15143 , n18605 );
    and g423 ( n2801 , n130 , n11758 );
    or g424 ( n17773 , n8564 , n6268 );
    or g425 ( n25290 , n5564 , n19382 );
    or g426 ( n39315 , n10060 , n24247 );
    or g427 ( n6142 , n32135 , n27516 );
    nor g428 ( n13019 , n24731 , n41402 );
    nor g429 ( n23764 , n32152 , n39754 );
    not g430 ( n5206 , n19340 );
    not g431 ( n9958 , n12006 );
    or g432 ( n26983 , n15007 , n39707 );
    xnor g433 ( n15347 , n10527 , n3046 );
    and g434 ( n4565 , n7924 , n11874 );
    and g435 ( n17442 , n12475 , n2911 );
    or g436 ( n18050 , n17798 , n21848 );
    and g437 ( n31779 , n6974 , n16217 );
    xnor g438 ( n2963 , n36009 , n4366 );
    not g439 ( n24939 , n22176 );
    not g440 ( n33775 , n2892 );
    and g441 ( n9908 , n3482 , n23499 );
    and g442 ( n18935 , n34377 , n41018 );
    and g443 ( n36305 , n38106 , n41435 );
    or g444 ( n5315 , n36602 , n36962 );
    xnor g445 ( n16860 , n2462 , n27975 );
    nor g446 ( n34182 , n38058 , n29434 );
    or g447 ( n7033 , n17665 , n41144 );
    xnor g448 ( n7014 , n30271 , n41099 );
    or g449 ( n14799 , n34099 , n42827 );
    not g450 ( n18275 , n30684 );
    or g451 ( n17051 , n39251 , n19698 );
    and g452 ( n26353 , n4771 , n20979 );
    or g453 ( n16710 , n19766 , n10365 );
    or g454 ( n13873 , n37392 , n19009 );
    or g455 ( n9683 , n14671 , n37591 );
    or g456 ( n17208 , n35301 , n36796 );
    and g457 ( n24020 , n34071 , n5015 );
    or g458 ( n28480 , n8539 , n11514 );
    or g459 ( n21418 , n28709 , n1712 );
    not g460 ( n495 , n29444 );
    and g461 ( n6838 , n25992 , n31133 );
    and g462 ( n18243 , n39891 , n31790 );
    not g463 ( n18311 , n17835 );
    and g464 ( n11068 , n25761 , n28011 );
    or g465 ( n36871 , n21574 , n15472 );
    or g466 ( n4032 , n39839 , n22115 );
    not g467 ( n38321 , n9777 );
    xnor g468 ( n5593 , n35867 , n8798 );
    xnor g469 ( n19322 , n2862 , n23993 );
    and g470 ( n40675 , n25484 , n41051 );
    or g471 ( n7246 , n29738 , n31271 );
    not g472 ( n5914 , n12251 );
    not g473 ( n24894 , n23921 );
    and g474 ( n21547 , n3310 , n5418 );
    nor g475 ( n5980 , n9576 , n24542 );
    xnor g476 ( n33846 , n39640 , n28453 );
    not g477 ( n41969 , n33889 );
    or g478 ( n42680 , n9292 , n27429 );
    or g479 ( n24869 , n39981 , n5242 );
    not g480 ( n9292 , n7762 );
    and g481 ( n8608 , n21052 , n23611 );
    or g482 ( n19412 , n33411 , n6392 );
    not g483 ( n29782 , n13373 );
    or g484 ( n42215 , n2124 , n22920 );
    xnor g485 ( n31512 , n9079 , n18731 );
    or g486 ( n18993 , n2492 , n9443 );
    and g487 ( n13012 , n4916 , n1766 );
    nor g488 ( n9416 , n35886 , n15060 );
    nor g489 ( n26010 , n39897 , n13485 );
    xnor g490 ( n20894 , n35553 , n4694 );
    nor g491 ( n482 , n17431 , n22594 );
    xnor g492 ( n22830 , n807 , n33357 );
    or g493 ( n7100 , n14484 , n2646 );
    or g494 ( n30278 , n14039 , n41616 );
    or g495 ( n38686 , n23759 , n4559 );
    or g496 ( n17531 , n4717 , n2335 );
    not g497 ( n31542 , n9691 );
    or g498 ( n6910 , n27444 , n14944 );
    or g499 ( n35060 , n6589 , n31945 );
    or g500 ( n26859 , n11340 , n8019 );
    nor g501 ( n32650 , n26058 , n9234 );
    or g502 ( n17309 , n18004 , n5813 );
    nor g503 ( n29941 , n24972 , n30590 );
    or g504 ( n20291 , n20294 , n15990 );
    or g505 ( n10370 , n16052 , n540 );
    not g506 ( n39059 , n205 );
    and g507 ( n24229 , n11371 , n5638 );
    and g508 ( n22640 , n10753 , n26694 );
    and g509 ( n23795 , n28449 , n29683 );
    or g510 ( n36545 , n23921 , n11914 );
    and g511 ( n6153 , n14101 , n41248 );
    or g512 ( n33812 , n25376 , n1292 );
    or g513 ( n13940 , n36245 , n5048 );
    or g514 ( n34286 , n36799 , n25178 );
    xnor g515 ( n39372 , n30512 , n36959 );
    and g516 ( n23953 , n21540 , n34112 );
    xnor g517 ( n15343 , n22799 , n16594 );
    xnor g518 ( n16297 , n31107 , n23998 );
    not g519 ( n26367 , n33595 );
    or g520 ( n40309 , n7839 , n33746 );
    and g521 ( n1122 , n8337 , n4858 );
    or g522 ( n10422 , n27627 , n1144 );
    and g523 ( n20835 , n18391 , n37240 );
    or g524 ( n30196 , n13646 , n12710 );
    or g525 ( n806 , n7488 , n14441 );
    nor g526 ( n30329 , n24591 , n24649 );
    and g527 ( n10310 , n12314 , n37650 );
    or g528 ( n14464 , n8721 , n24757 );
    or g529 ( n4079 , n15981 , n5657 );
    or g530 ( n16900 , n29938 , n27039 );
    and g531 ( n13730 , n20989 , n4497 );
    not g532 ( n21336 , n16965 );
    or g533 ( n27254 , n181 , n35337 );
    and g534 ( n42616 , n6401 , n38278 );
    xnor g535 ( n19740 , n18625 , n19143 );
    xnor g536 ( n35869 , n42064 , n18055 );
    or g537 ( n19814 , n4018 , n27529 );
    or g538 ( n8993 , n6478 , n29199 );
    xnor g539 ( n40887 , n19785 , n2048 );
    and g540 ( n24330 , n24368 , n37295 );
    or g541 ( n37091 , n33197 , n6316 );
    or g542 ( n9580 , n6954 , n5904 );
    or g543 ( n26300 , n32856 , n4669 );
    and g544 ( n9457 , n24968 , n10367 );
    and g545 ( n23815 , n42916 , n7054 );
    not g546 ( n28060 , n15151 );
    or g547 ( n12556 , n36815 , n35631 );
    and g548 ( n17134 , n14587 , n13031 );
    and g549 ( n18651 , n29493 , n11861 );
    or g550 ( n20398 , n7295 , n10811 );
    or g551 ( n1156 , n17515 , n2337 );
    or g552 ( n30420 , n37520 , n29719 );
    nor g553 ( n8875 , n23971 , n22735 );
    not g554 ( n36394 , n34414 );
    and g555 ( n20957 , n23945 , n27339 );
    and g556 ( n27700 , n40263 , n28978 );
    and g557 ( n34692 , n8301 , n25559 );
    not g558 ( n16939 , n13454 );
    xnor g559 ( n21254 , n12226 , n23821 );
    nor g560 ( n2202 , n9281 , n35020 );
    nor g561 ( n16381 , n28313 , n2322 );
    and g562 ( n37600 , n7796 , n28446 );
    or g563 ( n10803 , n15232 , n32025 );
    xnor g564 ( n35161 , n36712 , n37234 );
    and g565 ( n26070 , n21051 , n21549 );
    not g566 ( n28850 , n3361 );
    or g567 ( n36331 , n15569 , n7351 );
    not g568 ( n10414 , n26268 );
    and g569 ( n13191 , n6104 , n6008 );
    or g570 ( n3008 , n27703 , n19132 );
    xnor g571 ( n38760 , n35727 , n29012 );
    and g572 ( n2831 , n8849 , n22475 );
    not g573 ( n1572 , n41623 );
    nor g574 ( n40795 , n20067 , n39083 );
    nor g575 ( n3307 , n28787 , n12277 );
    not g576 ( n17703 , n2846 );
    not g577 ( n34445 , n6198 );
    or g578 ( n34020 , n18916 , n1144 );
    nor g579 ( n15631 , n30262 , n431 );
    or g580 ( n11000 , n35454 , n14728 );
    xnor g581 ( n37127 , n9133 , n8511 );
    or g582 ( n14670 , n26122 , n7445 );
    not g583 ( n27931 , n34043 );
    or g584 ( n2494 , n32433 , n31629 );
    and g585 ( n31469 , n6059 , n412 );
    and g586 ( n11647 , n27461 , n24334 );
    nor g587 ( n29210 , n1978 , n31332 );
    not g588 ( n9855 , n23716 );
    nor g589 ( n13239 , n14707 , n4650 );
    not g590 ( n19527 , n4956 );
    or g591 ( n9017 , n9473 , n30034 );
    or g592 ( n5029 , n16575 , n24793 );
    xnor g593 ( n32847 , n41013 , n20302 );
    or g594 ( n6134 , n14452 , n6125 );
    or g595 ( n12525 , n40350 , n6255 );
    and g596 ( n24450 , n9803 , n17816 );
    or g597 ( n35953 , n27108 , n37584 );
    or g598 ( n13177 , n2193 , n29852 );
    or g599 ( n27557 , n38976 , n21628 );
    or g600 ( n10471 , n12722 , n33970 );
    or g601 ( n22705 , n41380 , n42327 );
    or g602 ( n5453 , n19124 , n32060 );
    and g603 ( n19053 , n24099 , n42805 );
    or g604 ( n13196 , n5829 , n3290 );
    and g605 ( n24569 , n605 , n41341 );
    or g606 ( n33315 , n65 , n959 );
    or g607 ( n21241 , n4561 , n34036 );
    or g608 ( n20709 , n3464 , n27683 );
    or g609 ( n12517 , n10057 , n32364 );
    nor g610 ( n2332 , n30604 , n305 );
    and g611 ( n15955 , n20582 , n19012 );
    or g612 ( n12613 , n30507 , n31334 );
    xnor g613 ( n42199 , n24943 , n29067 );
    or g614 ( n19626 , n10425 , n20694 );
    and g615 ( n8526 , n38596 , n7755 );
    or g616 ( n34629 , n28438 , n7863 );
    and g617 ( n15215 , n32414 , n10469 );
    or g618 ( n29991 , n6120 , n16466 );
    and g619 ( n22032 , n6301 , n19042 );
    not g620 ( n26242 , n2562 );
    and g621 ( n7882 , n20479 , n14123 );
    and g622 ( n3726 , n9178 , n29472 );
    and g623 ( n1065 , n24754 , n32973 );
    and g624 ( n13480 , n8860 , n20843 );
    or g625 ( n15197 , n20258 , n40419 );
    or g626 ( n35147 , n16564 , n21390 );
    nor g627 ( n18239 , n16598 , n28786 );
    and g628 ( n1679 , n39987 , n22737 );
    nor g629 ( n14532 , n10735 , n11348 );
    or g630 ( n3908 , n24745 , n4631 );
    or g631 ( n18268 , n38124 , n16575 );
    xnor g632 ( n18500 , n34731 , n27546 );
    and g633 ( n41853 , n23047 , n14571 );
    not g634 ( n13354 , n31104 );
    xnor g635 ( n24461 , n27560 , n34386 );
    nor g636 ( n6267 , n34444 , n12818 );
    and g637 ( n642 , n40307 , n2693 );
    or g638 ( n22446 , n22619 , n13904 );
    or g639 ( n27591 , n23758 , n5200 );
    and g640 ( n41888 , n18129 , n21360 );
    and g641 ( n13003 , n7171 , n2636 );
    xnor g642 ( n26759 , n40757 , n20750 );
    or g643 ( n22045 , n11321 , n2671 );
    xnor g644 ( n25378 , n12524 , n36328 );
    not g645 ( n14810 , n31336 );
    or g646 ( n3397 , n14506 , n24965 );
    or g647 ( n30187 , n9187 , n1163 );
    not g648 ( n37061 , n12124 );
    nor g649 ( n38723 , n2199 , n30884 );
    nor g650 ( n32835 , n36117 , n35339 );
    or g651 ( n19752 , n17573 , n35346 );
    or g652 ( n5527 , n18244 , n9551 );
    and g653 ( n20148 , n10522 , n6951 );
    xnor g654 ( n41500 , n34562 , n36802 );
    or g655 ( n30762 , n4084 , n1160 );
    or g656 ( n7091 , n38149 , n37675 );
    and g657 ( n15000 , n31187 , n42317 );
    and g658 ( n26066 , n36003 , n39097 );
    or g659 ( n32994 , n26196 , n4264 );
    and g660 ( n35465 , n37765 , n33953 );
    not g661 ( n5174 , n39436 );
    or g662 ( n36246 , n30530 , n16369 );
    not g663 ( n30041 , n7024 );
    or g664 ( n30195 , n8004 , n19383 );
    nor g665 ( n34231 , n17193 , n1518 );
    or g666 ( n1662 , n34594 , n17735 );
    nor g667 ( n35372 , n24629 , n14843 );
    and g668 ( n4775 , n1315 , n9226 );
    xnor g669 ( n18814 , n42200 , n8258 );
    or g670 ( n41268 , n30318 , n26845 );
    xnor g671 ( n19491 , n15325 , n38756 );
    xnor g672 ( n27259 , n9453 , n9815 );
    not g673 ( n13409 , n6502 );
    or g674 ( n30021 , n12286 , n23802 );
    and g675 ( n17815 , n19330 , n23987 );
    xnor g676 ( n5464 , n35477 , n31006 );
    xnor g677 ( n36439 , n17285 , n38880 );
    xnor g678 ( n10881 , n12487 , n13783 );
    nor g679 ( n2854 , n28489 , n37292 );
    and g680 ( n23582 , n8818 , n23370 );
    or g681 ( n25225 , n7410 , n10780 );
    not g682 ( n42484 , n18328 );
    not g683 ( n16258 , n34658 );
    or g684 ( n33326 , n31187 , n38142 );
    and g685 ( n26858 , n784 , n745 );
    or g686 ( n8887 , n14471 , n35928 );
    or g687 ( n7054 , n7028 , n12408 );
    xnor g688 ( n31746 , n28313 , n29756 );
    xnor g689 ( n33496 , n2868 , n30404 );
    or g690 ( n28834 , n35483 , n30800 );
    or g691 ( n22420 , n9468 , n37247 );
    not g692 ( n18007 , n35063 );
    or g693 ( n2029 , n36932 , n35495 );
    and g694 ( n20021 , n33331 , n883 );
    or g695 ( n2954 , n40702 , n13774 );
    and g696 ( n16798 , n41889 , n24074 );
    or g697 ( n30109 , n13275 , n4716 );
    or g698 ( n7115 , n40676 , n29930 );
    or g699 ( n633 , n14877 , n20078 );
    nor g700 ( n38453 , n23266 , n41615 );
    xnor g701 ( n10327 , n32779 , n20207 );
    and g702 ( n924 , n38393 , n3324 );
    xnor g703 ( n11252 , n18689 , n8420 );
    and g704 ( n42424 , n26375 , n31581 );
    or g705 ( n9869 , n33611 , n11714 );
    nor g706 ( n21751 , n29427 , n40634 );
    or g707 ( n21943 , n33683 , n2542 );
    xnor g708 ( n24419 , n41013 , n12994 );
    or g709 ( n11100 , n33449 , n27818 );
    and g710 ( n42159 , n6620 , n24398 );
    or g711 ( n11392 , n14481 , n21821 );
    and g712 ( n19169 , n15840 , n6936 );
    or g713 ( n16492 , n6415 , n12858 );
    and g714 ( n2825 , n40615 , n9070 );
    and g715 ( n34229 , n5669 , n30727 );
    or g716 ( n20697 , n20797 , n3957 );
    and g717 ( n19674 , n5144 , n10901 );
    or g718 ( n22251 , n7948 , n30446 );
    nor g719 ( n7848 , n38922 , n488 );
    not g720 ( n42915 , n6402 );
    xnor g721 ( n13964 , n30315 , n25941 );
    not g722 ( n31917 , n32009 );
    xnor g723 ( n26503 , n784 , n24497 );
    not g724 ( n26847 , n1823 );
    and g725 ( n40434 , n39921 , n19938 );
    nor g726 ( n840 , n18866 , n16508 );
    or g727 ( n26781 , n972 , n11003 );
    nor g728 ( n40164 , n32374 , n25301 );
    and g729 ( n14218 , n17192 , n9491 );
    and g730 ( n42025 , n23260 , n38652 );
    nor g731 ( n32046 , n16598 , n7009 );
    or g732 ( n10596 , n41580 , n29024 );
    or g733 ( n35028 , n31452 , n38320 );
    nor g734 ( n25416 , n13336 , n33653 );
    nor g735 ( n17547 , n36961 , n33069 );
    nor g736 ( n11911 , n10434 , n18269 );
    xnor g737 ( n40205 , n29323 , n2020 );
    or g738 ( n36773 , n30865 , n6527 );
    nor g739 ( n11987 , n17120 , n13744 );
    or g740 ( n14630 , n42896 , n1852 );
    xnor g741 ( n35576 , n9142 , n12818 );
    or g742 ( n2737 , n8739 , n22767 );
    not g743 ( n41187 , n26764 );
    not g744 ( n6962 , n26358 );
    and g745 ( n503 , n26043 , n35117 );
    not g746 ( n9060 , n37552 );
    nor g747 ( n32627 , n4795 , n10406 );
    or g748 ( n30102 , n12620 , n17903 );
    nor g749 ( n17382 , n28026 , n38812 );
    and g750 ( n5889 , n12957 , n42149 );
    nor g751 ( n42905 , n20879 , n24958 );
    and g752 ( n25937 , n5652 , n41504 );
    not g753 ( n41972 , n28357 );
    or g754 ( n8775 , n16706 , n23211 );
    not g755 ( n41998 , n39065 );
    and g756 ( n16299 , n19107 , n14505 );
    or g757 ( n32459 , n16052 , n33987 );
    not g758 ( n6604 , n3144 );
    or g759 ( n35926 , n41338 , n31671 );
    and g760 ( n33295 , n23497 , n7576 );
    or g761 ( n12269 , n15429 , n39651 );
    xnor g762 ( n36931 , n22650 , n12213 );
    not g763 ( n2507 , n22863 );
    xnor g764 ( n41399 , n2461 , n36855 );
    or g765 ( n24346 , n5575 , n12129 );
    xnor g766 ( n41685 , n415 , n30272 );
    not g767 ( n33297 , n25994 );
    not g768 ( n37709 , n32573 );
    or g769 ( n5087 , n32808 , n31361 );
    or g770 ( n35760 , n41345 , n834 );
    and g771 ( n27485 , n96 , n12478 );
    not g772 ( n11663 , n19235 );
    or g773 ( n10726 , n23598 , n5167 );
    or g774 ( n13035 , n36296 , n5131 );
    and g775 ( n33813 , n7976 , n26829 );
    not g776 ( n25710 , n37196 );
    xnor g777 ( n2958 , n41843 , n27795 );
    not g778 ( n28319 , n21675 );
    or g779 ( n30827 , n21472 , n34308 );
    and g780 ( n4745 , n40777 , n28906 );
    and g781 ( n4421 , n1935 , n11002 );
    and g782 ( n388 , n26485 , n34464 );
    or g783 ( n5886 , n9518 , n41079 );
    or g784 ( n8570 , n28442 , n12206 );
    nor g785 ( n14560 , n5768 , n30355 );
    xnor g786 ( n25521 , n9412 , n27193 );
    and g787 ( n27406 , n3216 , n29179 );
    or g788 ( n602 , n36790 , n19497 );
    nor g789 ( n37373 , n10117 , n20815 );
    or g790 ( n14282 , n26845 , n13883 );
    nor g791 ( n28510 , n4345 , n33582 );
    not g792 ( n34960 , n29117 );
    nor g793 ( n39346 , n27286 , n16042 );
    xnor g794 ( n18454 , n27396 , n28737 );
    and g795 ( n33025 , n23304 , n16484 );
    not g796 ( n9512 , n5912 );
    and g797 ( n28666 , n27961 , n2780 );
    or g798 ( n32784 , n21204 , n10512 );
    or g799 ( n4349 , n40253 , n16597 );
    or g800 ( n25967 , n19438 , n38175 );
    or g801 ( n15871 , n5881 , n41371 );
    nor g802 ( n38359 , n13550 , n22059 );
    not g803 ( n34751 , n10759 );
    xnor g804 ( n4920 , n24218 , n32149 );
    or g805 ( n24304 , n14855 , n29062 );
    or g806 ( n17597 , n9160 , n25567 );
    or g807 ( n15336 , n35692 , n9375 );
    or g808 ( n4184 , n355 , n27036 );
    and g809 ( n9703 , n30370 , n40847 );
    or g810 ( n21519 , n27047 , n24592 );
    and g811 ( n40254 , n22576 , n24694 );
    and g812 ( n4866 , n10982 , n17755 );
    not g813 ( n2800 , n128 );
    or g814 ( n23356 , n36077 , n27849 );
    or g815 ( n16217 , n3097 , n19762 );
    xnor g816 ( n19772 , n40337 , n34289 );
    or g817 ( n16743 , n23901 , n38358 );
    xnor g818 ( n33851 , n542 , n9089 );
    or g819 ( n25176 , n29135 , n17472 );
    not g820 ( n26906 , n7862 );
    not g821 ( n25142 , n2018 );
    and g822 ( n40231 , n25165 , n6725 );
    and g823 ( n39155 , n25538 , n11292 );
    or g824 ( n42836 , n961 , n29703 );
    and g825 ( n28486 , n22970 , n20228 );
    or g826 ( n41589 , n28245 , n33022 );
    nor g827 ( n37333 , n34628 , n34908 );
    or g828 ( n8269 , n12232 , n21452 );
    and g829 ( n33428 , n18799 , n19598 );
    or g830 ( n12723 , n16052 , n19644 );
    or g831 ( n20927 , n39862 , n2247 );
    or g832 ( n27408 , n2068 , n24816 );
    or g833 ( n29464 , n34436 , n34069 );
    and g834 ( n34140 , n16454 , n23832 );
    not g835 ( n42220 , n3178 );
    not g836 ( n15354 , n2101 );
    not g837 ( n2069 , n15449 );
    not g838 ( n26810 , n2611 );
    nor g839 ( n25881 , n4253 , n33202 );
    and g840 ( n28578 , n32297 , n2252 );
    and g841 ( n4292 , n29036 , n39510 );
    not g842 ( n13433 , n34417 );
    nor g843 ( n40551 , n15070 , n42509 );
    and g844 ( n33963 , n29352 , n16867 );
    not g845 ( n15426 , n9637 );
    not g846 ( n35455 , n38862 );
    or g847 ( n28807 , n35263 , n37633 );
    and g848 ( n23127 , n30270 , n6645 );
    xnor g849 ( n41390 , n18702 , n16060 );
    or g850 ( n33490 , n21527 , n42694 );
    not g851 ( n22089 , n33632 );
    nor g852 ( n16485 , n36117 , n22131 );
    not g853 ( n25729 , n29963 );
    and g854 ( n35438 , n39874 , n3942 );
    or g855 ( n41932 , n5564 , n8188 );
    and g856 ( n3506 , n28218 , n36825 );
    or g857 ( n8999 , n9687 , n18314 );
    not g858 ( n25368 , n26824 );
    not g859 ( n17436 , n21293 );
    or g860 ( n25508 , n12549 , n11116 );
    not g861 ( n11843 , n16595 );
    not g862 ( n42895 , n38598 );
    and g863 ( n9338 , n13479 , n496 );
    and g864 ( n33422 , n14096 , n12436 );
    not g865 ( n20777 , n8202 );
    not g866 ( n32744 , n41206 );
    and g867 ( n19362 , n11880 , n173 );
    xnor g868 ( n14456 , n31107 , n27803 );
    and g869 ( n37042 , n40256 , n38553 );
    or g870 ( n4299 , n19983 , n31475 );
    or g871 ( n40050 , n36003 , n39097 );
    or g872 ( n27404 , n18918 , n9974 );
    or g873 ( n41810 , n41499 , n32980 );
    and g874 ( n33423 , n24950 , n14538 );
    not g875 ( n33667 , n29975 );
    not g876 ( n16465 , n29131 );
    and g877 ( n29558 , n3201 , n16262 );
    or g878 ( n14540 , n36071 , n16679 );
    nor g879 ( n35797 , n18395 , n37506 );
    nor g880 ( n41779 , n27745 , n7994 );
    xnor g881 ( n32447 , n2637 , n39812 );
    or g882 ( n32373 , n14707 , n13599 );
    or g883 ( n18151 , n2012 , n24006 );
    or g884 ( n7154 , n41859 , n26081 );
    or g885 ( n4722 , n40500 , n14294 );
    or g886 ( n1315 , n5577 , n32179 );
    not g887 ( n4102 , n40725 );
    or g888 ( n6457 , n8460 , n2064 );
    or g889 ( n24021 , n4862 , n24254 );
    not g890 ( n10332 , n38918 );
    not g891 ( n18785 , n29066 );
    or g892 ( n16461 , n32809 , n29939 );
    or g893 ( n11969 , n22859 , n33640 );
    or g894 ( n29765 , n35497 , n2876 );
    or g895 ( n22414 , n29091 , n5026 );
    or g896 ( n22737 , n3317 , n38135 );
    or g897 ( n30576 , n6180 , n15428 );
    nor g898 ( n39594 , n23325 , n25970 );
    xnor g899 ( n12115 , n35293 , n3592 );
    not g900 ( n20408 , n37477 );
    xnor g901 ( n29243 , n11614 , n2516 );
    not g902 ( n27924 , n16397 );
    and g903 ( n161 , n15551 , n3904 );
    and g904 ( n36724 , n25420 , n16931 );
    or g905 ( n1034 , n35148 , n7299 );
    or g906 ( n19954 , n38662 , n10232 );
    not g907 ( n24327 , n20425 );
    and g908 ( n30207 , n9307 , n33961 );
    or g909 ( n12629 , n19869 , n36817 );
    and g910 ( n16362 , n10800 , n23155 );
    nor g911 ( n16927 , n7100 , n15110 );
    nor g912 ( n35232 , n23345 , n7304 );
    or g913 ( n29491 , n39365 , n3677 );
    or g914 ( n34617 , n27180 , n28014 );
    or g915 ( n15849 , n7889 , n29551 );
    or g916 ( n13104 , n12392 , n24508 );
    not g917 ( n6762 , n36132 );
    nor g918 ( n39394 , n3883 , n36359 );
    not g919 ( n26845 , n17527 );
    and g920 ( n35503 , n25633 , n38369 );
    not g921 ( n5053 , n22681 );
    or g922 ( n22672 , n19494 , n18687 );
    or g923 ( n3181 , n927 , n39153 );
    or g924 ( n19972 , n42054 , n14716 );
    or g925 ( n20036 , n25279 , n41094 );
    nor g926 ( n35664 , n9233 , n41619 );
    or g927 ( n193 , n18775 , n19957 );
    nor g928 ( n2502 , n16812 , n3031 );
    not g929 ( n3113 , n33292 );
    or g930 ( n25533 , n3925 , n37245 );
    or g931 ( n38410 , n30001 , n3030 );
    nor g932 ( n3991 , n31882 , n728 );
    nor g933 ( n24438 , n18550 , n11673 );
    not g934 ( n23115 , n13746 );
    nor g935 ( n6509 , n5896 , n7649 );
    or g936 ( n28187 , n40295 , n19456 );
    not g937 ( n27476 , n14180 );
    not g938 ( n13984 , n40753 );
    nor g939 ( n9591 , n17272 , n42631 );
    or g940 ( n16727 , n32100 , n22501 );
    or g941 ( n10905 , n37450 , n3287 );
    not g942 ( n37255 , n3832 );
    or g943 ( n11757 , n25600 , n20756 );
    not g944 ( n11477 , n9917 );
    or g945 ( n3345 , n41534 , n33946 );
    or g946 ( n41770 , n16738 , n12802 );
    or g947 ( n8771 , n17091 , n21738 );
    or g948 ( n15115 , n12105 , n11163 );
    and g949 ( n42411 , n25270 , n10301 );
    or g950 ( n30416 , n10324 , n20174 );
    or g951 ( n22063 , n38453 , n15186 );
    and g952 ( n13926 , n10494 , n6530 );
    nor g953 ( n21732 , n15823 , n1817 );
    not g954 ( n40742 , n19741 );
    or g955 ( n21356 , n35069 , n14104 );
    and g956 ( n8763 , n20783 , n32075 );
    nor g957 ( n37334 , n9741 , n8257 );
    nor g958 ( n573 , n14268 , n13893 );
    xnor g959 ( n34592 , n24668 , n26676 );
    and g960 ( n15522 , n3379 , n11173 );
    or g961 ( n6833 , n13094 , n38327 );
    or g962 ( n24792 , n19707 , n16636 );
    or g963 ( n1937 , n32386 , n17174 );
    xnor g964 ( n28529 , n26579 , n25943 );
    or g965 ( n1165 , n15908 , n24254 );
    and g966 ( n2508 , n37551 , n3208 );
    not g967 ( n12651 , n27478 );
    and g968 ( n7868 , n26918 , n37865 );
    and g969 ( n37615 , n6624 , n18419 );
    or g970 ( n26414 , n24618 , n28253 );
    or g971 ( n16153 , n26944 , n21063 );
    not g972 ( n26406 , n6379 );
    or g973 ( n5352 , n28488 , n38793 );
    nor g974 ( n35469 , n348 , n15389 );
    not g975 ( n23349 , n38769 );
    and g976 ( n25488 , n29365 , n36333 );
    or g977 ( n35031 , n39539 , n39448 );
    or g978 ( n17795 , n24656 , n6622 );
    not g979 ( n12241 , n24712 );
    or g980 ( n32301 , n27840 , n29445 );
    or g981 ( n251 , n3583 , n37864 );
    or g982 ( n35675 , n25359 , n36848 );
    or g983 ( n30048 , n2042 , n24724 );
    or g984 ( n41221 , n17109 , n10992 );
    or g985 ( n12005 , n28143 , n38639 );
    or g986 ( n42410 , n18891 , n33583 );
    and g987 ( n38816 , n8869 , n29556 );
    xnor g988 ( n16936 , n4896 , n41997 );
    not g989 ( n20204 , n26268 );
    or g990 ( n42802 , n24180 , n14462 );
    not g991 ( n20557 , n6379 );
    or g992 ( n7323 , n23031 , n1502 );
    and g993 ( n18169 , n41850 , n17537 );
    or g994 ( n41141 , n35450 , n41287 );
    or g995 ( n19758 , n32089 , n5348 );
    or g996 ( n36845 , n6512 , n22154 );
    nor g997 ( n33209 , n19378 , n1514 );
    and g998 ( n31443 , n10843 , n8677 );
    or g999 ( n4942 , n10306 , n9130 );
    nor g1000 ( n11822 , n5144 , n1585 );
    and g1001 ( n26244 , n11287 , n14208 );
    or g1002 ( n22963 , n40703 , n11494 );
    or g1003 ( n21429 , n39596 , n4669 );
    not g1004 ( n13046 , n366 );
    not g1005 ( n29382 , n14888 );
    not g1006 ( n39723 , n7950 );
    or g1007 ( n18909 , n28392 , n8265 );
    or g1008 ( n6213 , n31823 , n37645 );
    or g1009 ( n42013 , n17853 , n16232 );
    xnor g1010 ( n828 , n14637 , n2229 );
    xnor g1011 ( n32544 , n13683 , n27112 );
    or g1012 ( n23958 , n31265 , n36032 );
    or g1013 ( n32932 , n24223 , n41849 );
    not g1014 ( n41127 , n23701 );
    and g1015 ( n2175 , n30465 , n1962 );
    and g1016 ( n31019 , n40418 , n2999 );
    and g1017 ( n40855 , n10842 , n21087 );
    or g1018 ( n29401 , n19987 , n31426 );
    nor g1019 ( n16294 , n31542 , n22652 );
    or g1020 ( n39976 , n8981 , n26740 );
    nor g1021 ( n10181 , n35301 , n16550 );
    not g1022 ( n22147 , n37698 );
    and g1023 ( n15948 , n39224 , n24906 );
    not g1024 ( n29593 , n41758 );
    or g1025 ( n12173 , n991 , n17100 );
    and g1026 ( n33482 , n20279 , n10340 );
    or g1027 ( n4615 , n26585 , n39098 );
    nor g1028 ( n24294 , n19522 , n12729 );
    and g1029 ( n5602 , n32630 , n5412 );
    nor g1030 ( n39906 , n16885 , n24528 );
    not g1031 ( n31503 , n36942 );
    nor g1032 ( n3729 , n22519 , n15973 );
    or g1033 ( n21115 , n37111 , n19475 );
    not g1034 ( n13216 , n28707 );
    nor g1035 ( n9812 , n6059 , n412 );
    or g1036 ( n42137 , n23153 , n35267 );
    xnor g1037 ( n1813 , n784 , n25614 );
    or g1038 ( n41582 , n15933 , n19778 );
    not g1039 ( n13711 , n38319 );
    or g1040 ( n8403 , n5964 , n36946 );
    not g1041 ( n8658 , n15956 );
    or g1042 ( n21256 , n40497 , n6397 );
    or g1043 ( n35020 , n25201 , n28249 );
    or g1044 ( n4367 , n30616 , n18173 );
    or g1045 ( n27441 , n35006 , n32792 );
    nor g1046 ( n6139 , n40532 , n24608 );
    nor g1047 ( n9523 , n22387 , n42173 );
    and g1048 ( n8707 , n33689 , n31380 );
    xnor g1049 ( n13269 , n842 , n7040 );
    nor g1050 ( n14090 , n14707 , n20936 );
    or g1051 ( n27866 , n39365 , n4156 );
    xnor g1052 ( n37038 , n14746 , n23955 );
    nor g1053 ( n21544 , n41856 , n24973 );
    not g1054 ( n16039 , n31775 );
    not g1055 ( n1703 , n26738 );
    or g1056 ( n32753 , n175 , n24565 );
    xnor g1057 ( n39301 , n21681 , n20745 );
    or g1058 ( n19094 , n1472 , n10111 );
    and g1059 ( n39055 , n3515 , n9854 );
    xnor g1060 ( n29631 , n37807 , n31968 );
    and g1061 ( n8988 , n30409 , n24947 );
    and g1062 ( n31292 , n42235 , n23416 );
    not g1063 ( n40337 , n28632 );
    or g1064 ( n14197 , n38048 , n17428 );
    and g1065 ( n12409 , n24808 , n32219 );
    and g1066 ( n13599 , n41257 , n24558 );
    or g1067 ( n10131 , n38340 , n1742 );
    or g1068 ( n28302 , n13005 , n41215 );
    not g1069 ( n19470 , n26477 );
    nor g1070 ( n38414 , n5001 , n15192 );
    and g1071 ( n15307 , n608 , n6935 );
    nor g1072 ( n943 , n19725 , n18325 );
    or g1073 ( n39738 , n6340 , n20403 );
    xnor g1074 ( n6444 , n18530 , n40303 );
    or g1075 ( n34476 , n4217 , n33041 );
    and g1076 ( n13194 , n28657 , n41716 );
    not g1077 ( n28160 , n20046 );
    and g1078 ( n21923 , n16834 , n17235 );
    not g1079 ( n16852 , n954 );
    and g1080 ( n42068 , n31797 , n16348 );
    and g1081 ( n8722 , n18489 , n8165 );
    not g1082 ( n9660 , n34443 );
    or g1083 ( n26827 , n11471 , n15854 );
    not g1084 ( n35221 , n4122 );
    not g1085 ( n1568 , n4147 );
    or g1086 ( n21800 , n33684 , n11755 );
    and g1087 ( n1934 , n36185 , n17116 );
    not g1088 ( n14172 , n37635 );
    or g1089 ( n7518 , n19898 , n6787 );
    not g1090 ( n22088 , n38454 );
    xnor g1091 ( n10098 , n37464 , n22630 );
    or g1092 ( n19850 , n9539 , n361 );
    nor g1093 ( n3698 , n23026 , n26288 );
    xnor g1094 ( n42181 , n18874 , n23590 );
    or g1095 ( n21737 , n5541 , n19762 );
    or g1096 ( n38285 , n22142 , n11031 );
    xnor g1097 ( n29232 , n34105 , n25200 );
    nor g1098 ( n36637 , n2249 , n2149 );
    not g1099 ( n15616 , n14580 );
    and g1100 ( n21319 , n2414 , n33192 );
    or g1101 ( n3384 , n17717 , n36606 );
    and g1102 ( n41985 , n17369 , n27248 );
    or g1103 ( n41453 , n10115 , n32752 );
    and g1104 ( n8675 , n19177 , n8717 );
    or g1105 ( n7380 , n31514 , n36314 );
    or g1106 ( n39606 , n35447 , n35521 );
    or g1107 ( n34812 , n18866 , n40241 );
    not g1108 ( n14642 , n17426 );
    and g1109 ( n11192 , n12861 , n28199 );
    not g1110 ( n8370 , n42877 );
    or g1111 ( n19541 , n36364 , n39193 );
    or g1112 ( n4800 , n1663 , n36653 );
    and g1113 ( n42246 , n5769 , n8239 );
    not g1114 ( n18875 , n12294 );
    or g1115 ( n15514 , n23562 , n13486 );
    or g1116 ( n41292 , n10045 , n2020 );
    not g1117 ( n781 , n21746 );
    or g1118 ( n36326 , n10651 , n1995 );
    or g1119 ( n25326 , n13843 , n37495 );
    or g1120 ( n34756 , n26789 , n11727 );
    and g1121 ( n16232 , n42114 , n6698 );
    and g1122 ( n37425 , n11842 , n28455 );
    not g1123 ( n22100 , n15356 );
    not g1124 ( n8821 , n41022 );
    or g1125 ( n35421 , n41728 , n12821 );
    nor g1126 ( n33236 , n38806 , n23141 );
    not g1127 ( n12161 , n38898 );
    or g1128 ( n13233 , n35302 , n31430 );
    or g1129 ( n31787 , n30171 , n32956 );
    not g1130 ( n10986 , n6704 );
    nor g1131 ( n39464 , n13420 , n25297 );
    or g1132 ( n19444 , n33691 , n41237 );
    or g1133 ( n30903 , n20412 , n36722 );
    and g1134 ( n31081 , n1501 , n19551 );
    xnor g1135 ( n422 , n36645 , n29632 );
    nor g1136 ( n8184 , n9350 , n20379 );
    xnor g1137 ( n29189 , n14594 , n15452 );
    or g1138 ( n17417 , n17063 , n2136 );
    xnor g1139 ( n11615 , n8612 , n11179 );
    or g1140 ( n14795 , n94 , n24300 );
    and g1141 ( n5356 , n21973 , n2733 );
    xnor g1142 ( n34275 , n11927 , n30156 );
    or g1143 ( n29697 , n22991 , n23984 );
    or g1144 ( n28720 , n14707 , n41318 );
    or g1145 ( n38065 , n8546 , n7617 );
    xnor g1146 ( n15199 , n40454 , n42037 );
    and g1147 ( n12236 , n33602 , n35680 );
    not g1148 ( n10383 , n11285 );
    nor g1149 ( n34108 , n30685 , n10925 );
    or g1150 ( n2945 , n15651 , n10722 );
    and g1151 ( n24011 , n39164 , n25189 );
    and g1152 ( n30119 , n38094 , n23573 );
    xnor g1153 ( n13031 , n726 , n42538 );
    xnor g1154 ( n532 , n6625 , n20936 );
    or g1155 ( n30341 , n6538 , n37321 );
    or g1156 ( n1621 , n17783 , n12388 );
    nor g1157 ( n32313 , n32331 , n6476 );
    nor g1158 ( n19683 , n37582 , n26386 );
    xnor g1159 ( n5372 , n41480 , n16941 );
    or g1160 ( n16731 , n30643 , n41275 );
    or g1161 ( n6938 , n11904 , n29850 );
    or g1162 ( n38903 , n5341 , n33914 );
    not g1163 ( n37222 , n22558 );
    or g1164 ( n10105 , n29058 , n25021 );
    or g1165 ( n17533 , n20482 , n39262 );
    or g1166 ( n24275 , n17216 , n38472 );
    or g1167 ( n40530 , n759 , n35193 );
    or g1168 ( n34425 , n32277 , n13375 );
    nor g1169 ( n20065 , n12105 , n6505 );
    xnor g1170 ( n3696 , n15145 , n39369 );
    or g1171 ( n25147 , n3738 , n13873 );
    not g1172 ( n22622 , n11861 );
    or g1173 ( n9715 , n2701 , n1168 );
    or g1174 ( n1618 , n14905 , n765 );
    not g1175 ( n35614 , n33991 );
    or g1176 ( n42834 , n24657 , n4838 );
    not g1177 ( n10967 , n35814 );
    nor g1178 ( n25904 , n19807 , n35427 );
    or g1179 ( n25999 , n23657 , n20038 );
    or g1180 ( n24829 , n33042 , n39696 );
    or g1181 ( n35152 , n35787 , n5258 );
    or g1182 ( n1795 , n22711 , n41337 );
    or g1183 ( n37431 , n4535 , n19733 );
    or g1184 ( n13459 , n6943 , n24452 );
    and g1185 ( n32564 , n13323 , n31589 );
    or g1186 ( n9022 , n32102 , n40419 );
    and g1187 ( n10790 , n17210 , n36097 );
    nor g1188 ( n5951 , n295 , n30173 );
    or g1189 ( n40533 , n8545 , n3728 );
    and g1190 ( n8289 , n29960 , n34645 );
    and g1191 ( n26999 , n32199 , n350 );
    or g1192 ( n38377 , n17259 , n6512 );
    and g1193 ( n33700 , n8915 , n14830 );
    or g1194 ( n40502 , n4492 , n28297 );
    or g1195 ( n21901 , n28840 , n14685 );
    xnor g1196 ( n14302 , n25619 , n2584 );
    or g1197 ( n25195 , n5941 , n33353 );
    xnor g1198 ( n15947 , n29740 , n12435 );
    or g1199 ( n19466 , n29531 , n28028 );
    not g1200 ( n40617 , n26613 );
    xnor g1201 ( n31215 , n29501 , n10031 );
    or g1202 ( n25923 , n4541 , n36292 );
    and g1203 ( n34460 , n35225 , n12329 );
    or g1204 ( n36358 , n25222 , n28822 );
    nor g1205 ( n42582 , n38696 , n1818 );
    and g1206 ( n32396 , n14293 , n23188 );
    or g1207 ( n2191 , n22133 , n2078 );
    or g1208 ( n12239 , n8844 , n20296 );
    or g1209 ( n1517 , n24226 , n1949 );
    and g1210 ( n14362 , n10139 , n35063 );
    nor g1211 ( n37110 , n33386 , n39440 );
    not g1212 ( n30068 , n25700 );
    or g1213 ( n3304 , n32534 , n28505 );
    or g1214 ( n40693 , n24243 , n1122 );
    not g1215 ( n2626 , n34729 );
    and g1216 ( n40367 , n8812 , n20192 );
    or g1217 ( n35590 , n37101 , n31231 );
    and g1218 ( n5358 , n37860 , n21883 );
    or g1219 ( n3832 , n32600 , n22495 );
    and g1220 ( n22024 , n5733 , n37453 );
    or g1221 ( n28579 , n31662 , n24623 );
    or g1222 ( n31143 , n18916 , n39216 );
    or g1223 ( n11387 , n33343 , n34069 );
    or g1224 ( n14597 , n444 , n12153 );
    not g1225 ( n10153 , n13716 );
    nor g1226 ( n17151 , n31379 , n39675 );
    and g1227 ( n28629 , n42013 , n31407 );
    or g1228 ( n18906 , n41381 , n12471 );
    or g1229 ( n39892 , n7030 , n29593 );
    and g1230 ( n6333 , n21895 , n12647 );
    or g1231 ( n34441 , n41923 , n15248 );
    or g1232 ( n1442 , n6578 , n9365 );
    not g1233 ( n40352 , n20392 );
    and g1234 ( n4338 , n20863 , n26278 );
    or g1235 ( n28287 , n33755 , n24157 );
    or g1236 ( n13682 , n12280 , n20349 );
    nor g1237 ( n42712 , n5175 , n10445 );
    xnor g1238 ( n29869 , n5144 , n36741 );
    not g1239 ( n27742 , n39442 );
    or g1240 ( n34412 , n41356 , n36533 );
    or g1241 ( n42639 , n2763 , n28646 );
    not g1242 ( n27035 , n21197 );
    and g1243 ( n3316 , n8152 , n885 );
    or g1244 ( n17677 , n13837 , n7730 );
    nor g1245 ( n4004 , n29824 , n9943 );
    or g1246 ( n2441 , n35479 , n14526 );
    not g1247 ( n30262 , n34173 );
    or g1248 ( n8596 , n16598 , n2394 );
    or g1249 ( n15260 , n8530 , n1970 );
    or g1250 ( n38240 , n41388 , n17576 );
    and g1251 ( n20161 , n6323 , n24311 );
    nor g1252 ( n4161 , n35255 , n9128 );
    nor g1253 ( n18809 , n28022 , n24774 );
    not g1254 ( n33026 , n26056 );
    xnor g1255 ( n10613 , n542 , n21084 );
    nor g1256 ( n36951 , n30005 , n16263 );
    or g1257 ( n14424 , n42769 , n6068 );
    not g1258 ( n42455 , n21151 );
    not g1259 ( n9752 , n231 );
    or g1260 ( n28353 , n32644 , n15366 );
    xnor g1261 ( n358 , n31581 , n26375 );
    or g1262 ( n40779 , n8775 , n29440 );
    or g1263 ( n12735 , n5449 , n21268 );
    or g1264 ( n39627 , n14529 , n21111 );
    or g1265 ( n12141 , n9417 , n1200 );
    or g1266 ( n22741 , n24745 , n4321 );
    and g1267 ( n26111 , n6149 , n18802 );
    not g1268 ( n22177 , n22555 );
    and g1269 ( n5707 , n17064 , n41476 );
    and g1270 ( n35981 , n29399 , n24469 );
    and g1271 ( n23936 , n36638 , n32932 );
    not g1272 ( n5375 , n41854 );
    not g1273 ( n14549 , n29821 );
    not g1274 ( n27086 , n19435 );
    or g1275 ( n14869 , n39825 , n2786 );
    xnor g1276 ( n30205 , n30752 , n22924 );
    and g1277 ( n34495 , n28858 , n41953 );
    nor g1278 ( n2043 , n708 , n24038 );
    or g1279 ( n12406 , n17851 , n16447 );
    nor g1280 ( n817 , n35789 , n30631 );
    nor g1281 ( n34150 , n14485 , n15195 );
    nor g1282 ( n36606 , n25588 , n5377 );
    or g1283 ( n38780 , n42857 , n2802 );
    and g1284 ( n34712 , n2282 , n8958 );
    or g1285 ( n1445 , n34561 , n41678 );
    and g1286 ( n17515 , n276 , n18227 );
    and g1287 ( n14276 , n11271 , n2073 );
    and g1288 ( n35339 , n21492 , n14736 );
    or g1289 ( n28751 , n3420 , n37703 );
    or g1290 ( n2428 , n4812 , n5122 );
    or g1291 ( n21087 , n18937 , n19960 );
    xnor g1292 ( n77 , n40 , n4735 );
    or g1293 ( n8350 , n9676 , n11581 );
    nor g1294 ( n39038 , n3540 , n23465 );
    and g1295 ( n39977 , n30006 , n22047 );
    nor g1296 ( n29936 , n34416 , n27354 );
    and g1297 ( n41521 , n41677 , n41814 );
    or g1298 ( n32429 , n37214 , n37605 );
    not g1299 ( n20096 , n33430 );
    nor g1300 ( n17948 , n14707 , n40043 );
    or g1301 ( n40711 , n27666 , n21547 );
    nor g1302 ( n12350 , n33418 , n36937 );
    and g1303 ( n1852 , n8136 , n10381 );
    or g1304 ( n15141 , n27690 , n2276 );
    and g1305 ( n15184 , n29087 , n15859 );
    xnor g1306 ( n39692 , n31099 , n37978 );
    not g1307 ( n13111 , n22378 );
    and g1308 ( n15905 , n3435 , n1079 );
    not g1309 ( n36345 , n31522 );
    xnor g1310 ( n34349 , n11426 , n39173 );
    and g1311 ( n36411 , n38749 , n8317 );
    not g1312 ( n24608 , n42395 );
    or g1313 ( n24568 , n19580 , n2813 );
    not g1314 ( n17655 , n24766 );
    nor g1315 ( n35773 , n4546 , n11405 );
    nor g1316 ( n28611 , n14471 , n4666 );
    or g1317 ( n27811 , n37129 , n11607 );
    not g1318 ( n11629 , n12308 );
    or g1319 ( n15345 , n16973 , n41145 );
    and g1320 ( n4193 , n18500 , n36900 );
    or g1321 ( n31381 , n8228 , n2095 );
    not g1322 ( n19582 , n30826 );
    nor g1323 ( n11849 , n35790 , n39821 );
    or g1324 ( n2498 , n40995 , n13145 );
    not g1325 ( n39544 , n13042 );
    or g1326 ( n20797 , n18212 , n29640 );
    or g1327 ( n13922 , n28832 , n11947 );
    and g1328 ( n13251 , n35230 , n12600 );
    xnor g1329 ( n6657 , n30615 , n37612 );
    or g1330 ( n30811 , n18622 , n28418 );
    nor g1331 ( n9649 , n27961 , n31546 );
    not g1332 ( n17426 , n28411 );
    not g1333 ( n33250 , n17101 );
    or g1334 ( n25979 , n27232 , n1177 );
    or g1335 ( n16681 , n36583 , n25215 );
    and g1336 ( n9233 , n20387 , n18553 );
    xnor g1337 ( n1954 , n3994 , n25588 );
    or g1338 ( n41658 , n37362 , n26435 );
    or g1339 ( n42212 , n8969 , n25621 );
    and g1340 ( n2977 , n7162 , n25272 );
    not g1341 ( n35861 , n39057 );
    or g1342 ( n9560 , n40703 , n11200 );
    and g1343 ( n10890 , n21644 , n703 );
    not g1344 ( n24053 , n15396 );
    and g1345 ( n15211 , n1382 , n19800 );
    or g1346 ( n29001 , n18093 , n24782 );
    nor g1347 ( n36893 , n29859 , n17574 );
    nor g1348 ( n40138 , n34565 , n37724 );
    or g1349 ( n27073 , n29857 , n15498 );
    or g1350 ( n15520 , n9417 , n37947 );
    nor g1351 ( n40039 , n1507 , n6949 );
    nor g1352 ( n27584 , n28872 , n28937 );
    and g1353 ( n457 , n26751 , n10959 );
    or g1354 ( n39235 , n22 , n12220 );
    or g1355 ( n1403 , n15388 , n6925 );
    or g1356 ( n6251 , n13598 , n27666 );
    or g1357 ( n17897 , n39385 , n38982 );
    not g1358 ( n12896 , n16285 );
    and g1359 ( n10743 , n6210 , n14974 );
    or g1360 ( n41618 , n26492 , n35179 );
    or g1361 ( n29795 , n14920 , n41124 );
    not g1362 ( n38388 , n7008 );
    nor g1363 ( n35549 , n28431 , n4482 );
    and g1364 ( n29076 , n35162 , n7192 );
    not g1365 ( n3954 , n22187 );
    or g1366 ( n34614 , n20921 , n11805 );
    and g1367 ( n8052 , n21214 , n36173 );
    xnor g1368 ( n17549 , n11633 , n20565 );
    not g1369 ( n21381 , n40299 );
    and g1370 ( n36955 , n42541 , n33587 );
    not g1371 ( n2042 , n22022 );
    not g1372 ( n5347 , n26022 );
    or g1373 ( n33891 , n14673 , n11253 );
    or g1374 ( n24406 , n14240 , n3828 );
    or g1375 ( n20798 , n20244 , n31346 );
    not g1376 ( n16204 , n27950 );
    or g1377 ( n34396 , n6708 , n24104 );
    or g1378 ( n23083 , n30275 , n1405 );
    and g1379 ( n14442 , n720 , n31360 );
    and g1380 ( n9801 , n40364 , n30096 );
    not g1381 ( n2794 , n38985 );
    and g1382 ( n25161 , n26734 , n25260 );
    nor g1383 ( n8732 , n36667 , n3267 );
    and g1384 ( n5831 , n33614 , n596 );
    xnor g1385 ( n26899 , n36712 , n339 );
    or g1386 ( n30955 , n32288 , n37131 );
    or g1387 ( n15612 , n22926 , n19781 );
    nor g1388 ( n24054 , n5964 , n17432 );
    xnor g1389 ( n23242 , n36094 , n28275 );
    and g1390 ( n2436 , n38330 , n28091 );
    or g1391 ( n8030 , n19523 , n36244 );
    xnor g1392 ( n38943 , n3970 , n39878 );
    and g1393 ( n10242 , n20500 , n38875 );
    or g1394 ( n17080 , n21895 , n12647 );
    not g1395 ( n38926 , n39323 );
    or g1396 ( n13755 , n39823 , n18075 );
    or g1397 ( n15319 , n5091 , n14945 );
    or g1398 ( n9957 , n30683 , n17383 );
    or g1399 ( n5117 , n12383 , n513 );
    nor g1400 ( n12710 , n14746 , n15893 );
    not g1401 ( n30638 , n10010 );
    or g1402 ( n39592 , n20697 , n25458 );
    or g1403 ( n24571 , n8031 , n29273 );
    or g1404 ( n23853 , n28647 , n5035 );
    or g1405 ( n41423 , n3432 , n10866 );
    not g1406 ( n22855 , n11058 );
    or g1407 ( n25467 , n37161 , n2213 );
    or g1408 ( n587 , n18072 , n15451 );
    xnor g1409 ( n7300 , n11436 , n40335 );
    or g1410 ( n24874 , n644 , n18591 );
    xnor g1411 ( n10418 , n42666 , n38367 );
    or g1412 ( n9628 , n35386 , n20590 );
    or g1413 ( n278 , n33911 , n42368 );
    or g1414 ( n15337 , n15934 , n19894 );
    not g1415 ( n31227 , n13470 );
    not g1416 ( n7975 , n928 );
    nor g1417 ( n16103 , n974 , n4633 );
    xnor g1418 ( n17949 , n12506 , n23622 );
    nor g1419 ( n12784 , n38146 , n40990 );
    xnor g1420 ( n11815 , n3500 , n38310 );
    or g1421 ( n12301 , n25965 , n35740 );
    and g1422 ( n37894 , n27855 , n31855 );
    or g1423 ( n16572 , n7314 , n2644 );
    and g1424 ( n30017 , n6768 , n1366 );
    nor g1425 ( n27626 , n19164 , n2436 );
    or g1426 ( n6630 , n19954 , n1340 );
    xnor g1427 ( n18986 , n4620 , n41235 );
    or g1428 ( n34295 , n14074 , n35907 );
    or g1429 ( n29277 , n11567 , n25413 );
    and g1430 ( n22924 , n24036 , n39504 );
    xnor g1431 ( n41041 , n22296 , n23102 );
    or g1432 ( n18745 , n37292 , n10967 );
    not g1433 ( n2451 , n18138 );
    and g1434 ( n13635 , n40900 , n17041 );
    and g1435 ( n40450 , n30766 , n9450 );
    or g1436 ( n10114 , n12851 , n42539 );
    not g1437 ( n3146 , n36372 );
    nor g1438 ( n36280 , n36117 , n36883 );
    or g1439 ( n20801 , n26238 , n6512 );
    not g1440 ( n11449 , n41208 );
    and g1441 ( n281 , n18256 , n1907 );
    not g1442 ( n38064 , n27408 );
    or g1443 ( n16988 , n12489 , n35772 );
    or g1444 ( n4325 , n9318 , n17062 );
    and g1445 ( n18842 , n21213 , n2782 );
    not g1446 ( n15590 , n24856 );
    nor g1447 ( n42206 , n21115 , n19692 );
    or g1448 ( n31340 , n33361 , n37871 );
    or g1449 ( n31408 , n33392 , n38408 );
    nor g1450 ( n15210 , n41970 , n32769 );
    nor g1451 ( n29099 , n15860 , n6718 );
    and g1452 ( n33910 , n6587 , n17140 );
    not g1453 ( n30508 , n23191 );
    or g1454 ( n9853 , n11097 , n7071 );
    not g1455 ( n5722 , n15565 );
    or g1456 ( n36438 , n31090 , n31950 );
    and g1457 ( n1061 , n21680 , n8110 );
    not g1458 ( n14925 , n36114 );
    not g1459 ( n12871 , n40630 );
    or g1460 ( n16024 , n6063 , n8395 );
    or g1461 ( n26657 , n7139 , n10975 );
    or g1462 ( n20550 , n17193 , n26197 );
    and g1463 ( n19000 , n13311 , n28365 );
    or g1464 ( n24298 , n36470 , n11026 );
    not g1465 ( n5193 , n19692 );
    nor g1466 ( n15428 , n1507 , n23974 );
    xnor g1467 ( n19373 , n9155 , n7893 );
    and g1468 ( n9075 , n3597 , n1428 );
    or g1469 ( n24361 , n40449 , n3311 );
    and g1470 ( n2672 , n9268 , n31377 );
    not g1471 ( n40468 , n14081 );
    or g1472 ( n30829 , n6598 , n16682 );
    not g1473 ( n23921 , n23500 );
    not g1474 ( n27284 , n18870 );
    or g1475 ( n39031 , n7864 , n21378 );
    or g1476 ( n17621 , n19535 , n3031 );
    or g1477 ( n17996 , n14420 , n25390 );
    nor g1478 ( n13077 , n14707 , n8772 );
    or g1479 ( n28334 , n17293 , n40712 );
    or g1480 ( n39434 , n36880 , n1113 );
    not g1481 ( n773 , n4802 );
    not g1482 ( n41577 , n38929 );
    or g1483 ( n20599 , n41601 , n3353 );
    xnor g1484 ( n32604 , n20331 , n10965 );
    not g1485 ( n18235 , n19178 );
    xnor g1486 ( n7316 , n14642 , n16856 );
    or g1487 ( n27681 , n17313 , n9285 );
    and g1488 ( n39250 , n1506 , n27677 );
    not g1489 ( n7511 , n33915 );
    not g1490 ( n42667 , n26137 );
    or g1491 ( n41524 , n33747 , n38107 );
    and g1492 ( n36376 , n5086 , n39238 );
    not g1493 ( n1316 , n38898 );
    or g1494 ( n31717 , n22892 , n4589 );
    or g1495 ( n16265 , n5597 , n6719 );
    and g1496 ( n2537 , n42761 , n36170 );
    and g1497 ( n23993 , n19872 , n3025 );
    not g1498 ( n8270 , n29494 );
    or g1499 ( n16645 , n38592 , n5456 );
    and g1500 ( n16879 , n7915 , n5410 );
    or g1501 ( n33895 , n25317 , n6438 );
    and g1502 ( n7752 , n9950 , n1916 );
    or g1503 ( n12911 , n35377 , n28361 );
    xnor g1504 ( n33921 , n37153 , n28937 );
    and g1505 ( n6536 , n38028 , n20959 );
    xnor g1506 ( n36579 , n11436 , n17657 );
    or g1507 ( n31646 , n38909 , n36687 );
    not g1508 ( n27758 , n6790 );
    or g1509 ( n37511 , n23971 , n13781 );
    nor g1510 ( n22240 , n7356 , n28750 );
    or g1511 ( n19299 , n15149 , n31250 );
    nor g1512 ( n26730 , n33134 , n42538 );
    or g1513 ( n8197 , n29879 , n11301 );
    or g1514 ( n31384 , n21118 , n30978 );
    or g1515 ( n34213 , n22623 , n37347 );
    or g1516 ( n9552 , n14455 , n32097 );
    or g1517 ( n2852 , n30658 , n904 );
    or g1518 ( n21231 , n11640 , n38600 );
    or g1519 ( n38203 , n36569 , n21231 );
    and g1520 ( n750 , n365 , n3604 );
    and g1521 ( n39137 , n10683 , n40958 );
    or g1522 ( n27940 , n13117 , n7169 );
    or g1523 ( n42819 , n20092 , n24399 );
    xnor g1524 ( n27740 , n41515 , n8216 );
    not g1525 ( n13651 , n1941 );
    not g1526 ( n12821 , n6913 );
    or g1527 ( n10425 , n35193 , n36742 );
    and g1528 ( n34646 , n23469 , n29680 );
    or g1529 ( n2594 , n4670 , n37955 );
    or g1530 ( n9077 , n42558 , n16325 );
    or g1531 ( n16269 , n12112 , n17720 );
    or g1532 ( n33483 , n10160 , n13952 );
    or g1533 ( n11175 , n37340 , n41649 );
    or g1534 ( n15037 , n21338 , n14489 );
    or g1535 ( n16854 , n17292 , n9740 );
    xnor g1536 ( n4024 , n105 , n22640 );
    or g1537 ( n20491 , n15253 , n34955 );
    and g1538 ( n19664 , n8203 , n21737 );
    or g1539 ( n32562 , n42867 , n34949 );
    or g1540 ( n615 , n40476 , n12559 );
    nor g1541 ( n28520 , n26053 , n15193 );
    or g1542 ( n35793 , n32213 , n579 );
    nor g1543 ( n220 , n36697 , n37305 );
    and g1544 ( n36568 , n15910 , n16596 );
    and g1545 ( n6229 , n18678 , n14138 );
    nor g1546 ( n20268 , n4546 , n17367 );
    xnor g1547 ( n16525 , n18859 , n10249 );
    nor g1548 ( n39759 , n5494 , n2019 );
    nor g1549 ( n25494 , n11460 , n40643 );
    not g1550 ( n16703 , n37833 );
    xnor g1551 ( n38946 , n41218 , n4866 );
    not g1552 ( n4157 , n8382 );
    nor g1553 ( n27601 , n42780 , n39720 );
    and g1554 ( n5670 , n26622 , n14744 );
    and g1555 ( n15688 , n32889 , n19234 );
    nor g1556 ( n21338 , n14193 , n13020 );
    or g1557 ( n14862 , n31988 , n11931 );
    or g1558 ( n23245 , n34965 , n5124 );
    and g1559 ( n33741 , n9127 , n42821 );
    not g1560 ( n16534 , n17490 );
    not g1561 ( n20900 , n33702 );
    and g1562 ( n9987 , n40630 , n27830 );
    and g1563 ( n15967 , n22514 , n15586 );
    and g1564 ( n1203 , n15975 , n13772 );
    xnor g1565 ( n13574 , n618 , n1076 );
    not g1566 ( n32783 , n20485 );
    not g1567 ( n31940 , n25411 );
    or g1568 ( n15595 , n14500 , n33859 );
    and g1569 ( n24162 , n7607 , n34005 );
    or g1570 ( n26485 , n6872 , n41981 );
    nor g1571 ( n3870 , n3944 , n18295 );
    and g1572 ( n36407 , n25593 , n5251 );
    or g1573 ( n5208 , n14487 , n31198 );
    and g1574 ( n12449 , n15665 , n13976 );
    or g1575 ( n33871 , n32759 , n38981 );
    xnor g1576 ( n42472 , n31539 , n16832 );
    xnor g1577 ( n24573 , n12161 , n41405 );
    and g1578 ( n3627 , n640 , n40633 );
    or g1579 ( n41378 , n39828 , n40004 );
    and g1580 ( n36182 , n10157 , n27307 );
    or g1581 ( n557 , n34708 , n22353 );
    and g1582 ( n16159 , n17481 , n26633 );
    or g1583 ( n2414 , n11324 , n35732 );
    or g1584 ( n40463 , n30895 , n39810 );
    xnor g1585 ( n20573 , n12836 , n23233 );
    or g1586 ( n18577 , n34832 , n22156 );
    and g1587 ( n4850 , n27200 , n39835 );
    or g1588 ( n12918 , n22666 , n11134 );
    or g1589 ( n19999 , n7541 , n29545 );
    or g1590 ( n34950 , n3108 , n10363 );
    not g1591 ( n20811 , n26902 );
    xnor g1592 ( n30778 , n38081 , n35807 );
    nor g1593 ( n42677 , n13118 , n28828 );
    and g1594 ( n34428 , n15630 , n14015 );
    or g1595 ( n20108 , n26765 , n33785 );
    or g1596 ( n21144 , n17120 , n19004 );
    or g1597 ( n1700 , n12024 , n16882 );
    or g1598 ( n21832 , n38841 , n40882 );
    xnor g1599 ( n25459 , n12358 , n25229 );
    not g1600 ( n22482 , n8232 );
    xnor g1601 ( n25065 , n40176 , n35306 );
    not g1602 ( n23930 , n9923 );
    not g1603 ( n10152 , n17441 );
    xnor g1604 ( n35734 , n42739 , n22511 );
    not g1605 ( n16633 , n9441 );
    nor g1606 ( n34988 , n8935 , n32004 );
    or g1607 ( n42482 , n33995 , n6102 );
    nor g1608 ( n24933 , n5291 , n4592 );
    and g1609 ( n3654 , n36745 , n15450 );
    xnor g1610 ( n33944 , n28225 , n33922 );
    and g1611 ( n11863 , n34883 , n22668 );
    or g1612 ( n16779 , n14776 , n13407 );
    or g1613 ( n11354 , n13767 , n20796 );
    or g1614 ( n3332 , n21534 , n26202 );
    not g1615 ( n28415 , n16699 );
    or g1616 ( n716 , n34616 , n28791 );
    and g1617 ( n36420 , n22107 , n18899 );
    or g1618 ( n31824 , n40323 , n42214 );
    or g1619 ( n3699 , n31566 , n36983 );
    xnor g1620 ( n9815 , n3713 , n2793 );
    and g1621 ( n41980 , n33725 , n32101 );
    and g1622 ( n29755 , n21827 , n13027 );
    or g1623 ( n32622 , n29418 , n32410 );
    xnor g1624 ( n39410 , n36628 , n27203 );
    or g1625 ( n11213 , n34565 , n37073 );
    not g1626 ( n8591 , n13111 );
    and g1627 ( n41346 , n41838 , n39476 );
    xnor g1628 ( n26538 , n40232 , n5896 );
    nor g1629 ( n33572 , n31916 , n36255 );
    xnor g1630 ( n20715 , n27035 , n40139 );
    and g1631 ( n10654 , n14138 , n26441 );
    xnor g1632 ( n21669 , n30832 , n6837 );
    not g1633 ( n8108 , n31729 );
    xnor g1634 ( n15311 , n7922 , n23337 );
    nor g1635 ( n38115 , n39367 , n9399 );
    not g1636 ( n3976 , n520 );
    and g1637 ( n38279 , n7550 , n37410 );
    or g1638 ( n29415 , n35133 , n753 );
    or g1639 ( n2431 , n41655 , n20648 );
    or g1640 ( n12681 , n28352 , n31170 );
    and g1641 ( n6148 , n3963 , n3060 );
    nor g1642 ( n1902 , n22089 , n18078 );
    nor g1643 ( n6764 , n35965 , n25107 );
    xnor g1644 ( n41559 , n32470 , n29162 );
    nor g1645 ( n7696 , n1015 , n35934 );
    nor g1646 ( n34546 , n25296 , n19032 );
    xnor g1647 ( n28251 , n11436 , n18908 );
    nor g1648 ( n18403 , n14226 , n1934 );
    or g1649 ( n12534 , n10274 , n42015 );
    or g1650 ( n12985 , n30508 , n4350 );
    nor g1651 ( n12127 , n24156 , n24363 );
    not g1652 ( n20920 , n20553 );
    and g1653 ( n8844 , n20119 , n11946 );
    not g1654 ( n4231 , n30869 );
    and g1655 ( n23313 , n27757 , n41648 );
    and g1656 ( n782 , n25088 , n21790 );
    and g1657 ( n38034 , n37726 , n21147 );
    not g1658 ( n36569 , n19334 );
    or g1659 ( n33533 , n10903 , n3978 );
    not g1660 ( n13394 , n30930 );
    or g1661 ( n28162 , n38621 , n26353 );
    not g1662 ( n7313 , n32861 );
    xnor g1663 ( n24918 , n12207 , n35123 );
    or g1664 ( n27943 , n1032 , n31580 );
    nor g1665 ( n12568 , n38964 , n21421 );
    not g1666 ( n14831 , n8879 );
    or g1667 ( n42750 , n27558 , n27660 );
    xnor g1668 ( n16162 , n36998 , n13416 );
    not g1669 ( n5389 , n7359 );
    not g1670 ( n42534 , n13152 );
    not g1671 ( n19753 , n18584 );
    nor g1672 ( n9484 , n16039 , n9727 );
    or g1673 ( n12720 , n37664 , n7768 );
    and g1674 ( n24618 , n14835 , n12801 );
    nor g1675 ( n25391 , n3795 , n12620 );
    not g1676 ( n40128 , n39742 );
    nor g1677 ( n39122 , n5768 , n8516 );
    xnor g1678 ( n21504 , n8591 , n8451 );
    or g1679 ( n2663 , n24749 , n31326 );
    xnor g1680 ( n26507 , n32297 , n41509 );
    or g1681 ( n38787 , n38678 , n19744 );
    xnor g1682 ( n6486 , n41901 , n39007 );
    or g1683 ( n36505 , n40947 , n33289 );
    or g1684 ( n28822 , n36235 , n28308 );
    or g1685 ( n24744 , n27294 , n35277 );
    nor g1686 ( n24350 , n23585 , n957 );
    not g1687 ( n9168 , n26538 );
    nor g1688 ( n41902 , n15050 , n40474 );
    not g1689 ( n15611 , n28821 );
    or g1690 ( n29221 , n41721 , n37633 );
    xnor g1691 ( n26335 , n11131 , n4973 );
    xnor g1692 ( n17455 , n11670 , n4140 );
    and g1693 ( n8485 , n2326 , n34211 );
    and g1694 ( n35756 , n28939 , n6321 );
    nor g1695 ( n28127 , n14471 , n24260 );
    nor g1696 ( n2909 , n14707 , n31961 );
    and g1697 ( n31762 , n5045 , n21946 );
    and g1698 ( n37510 , n9946 , n34756 );
    or g1699 ( n34366 , n34391 , n32780 );
    not g1700 ( n6781 , n30627 );
    nor g1701 ( n16336 , n26454 , n8484 );
    and g1702 ( n21555 , n26009 , n37343 );
    xnor g1703 ( n14375 , n15972 , n10035 );
    or g1704 ( n20342 , n42855 , n32256 );
    or g1705 ( n13901 , n2434 , n24547 );
    and g1706 ( n26731 , n33925 , n13935 );
    not g1707 ( n6636 , n37094 );
    and g1708 ( n12258 , n36505 , n30187 );
    or g1709 ( n36166 , n33334 , n40702 );
    and g1710 ( n13992 , n31729 , n15059 );
    xnor g1711 ( n35264 , n22243 , n9547 );
    not g1712 ( n34050 , n4990 );
    and g1713 ( n9253 , n22685 , n25757 );
    not g1714 ( n25172 , n30405 );
    not g1715 ( n28318 , n34163 );
    not g1716 ( n33224 , n22845 );
    xnor g1717 ( n22354 , n32517 , n16974 );
    or g1718 ( n38598 , n32825 , n6227 );
    or g1719 ( n2094 , n26845 , n35533 );
    and g1720 ( n22531 , n39872 , n1634 );
    or g1721 ( n26499 , n24755 , n4660 );
    or g1722 ( n22690 , n41040 , n33954 );
    not g1723 ( n27734 , n27964 );
    not g1724 ( n27925 , n17342 );
    or g1725 ( n41076 , n14945 , n31006 );
    or g1726 ( n35661 , n27919 , n31950 );
    xnor g1727 ( n12274 , n16546 , n34686 );
    xnor g1728 ( n41837 , n18990 , n16966 );
    or g1729 ( n29916 , n41466 , n5110 );
    not g1730 ( n39962 , n13696 );
    or g1731 ( n29633 , n28805 , n14776 );
    xnor g1732 ( n8724 , n41718 , n34430 );
    xnor g1733 ( n6338 , n12024 , n39056 );
    or g1734 ( n37102 , n18230 , n26404 );
    and g1735 ( n9750 , n8261 , n22887 );
    and g1736 ( n21050 , n25867 , n32282 );
    or g1737 ( n29297 , n32321 , n10898 );
    not g1738 ( n38060 , n13167 );
    or g1739 ( n30617 , n1999 , n29286 );
    or g1740 ( n24181 , n17014 , n35742 );
    xnor g1741 ( n16105 , n7836 , n15746 );
    not g1742 ( n39551 , n39011 );
    not g1743 ( n31346 , n38289 );
    xnor g1744 ( n530 , n105 , n41556 );
    xnor g1745 ( n19725 , n39531 , n18421 );
    or g1746 ( n8528 , n26474 , n3423 );
    nor g1747 ( n27523 , n4388 , n13814 );
    xnor g1748 ( n13858 , n29452 , n583 );
    nor g1749 ( n29849 , n13272 , n28394 );
    or g1750 ( n5617 , n40661 , n23133 );
    or g1751 ( n42348 , n26879 , n37982 );
    or g1752 ( n20414 , n8847 , n38237 );
    or g1753 ( n23352 , n38022 , n22949 );
    not g1754 ( n25042 , n37306 );
    or g1755 ( n14288 , n32053 , n21409 );
    or g1756 ( n36442 , n313 , n25690 );
    xnor g1757 ( n32772 , n36106 , n3614 );
    and g1758 ( n16536 , n39717 , n7762 );
    or g1759 ( n8965 , n31830 , n20250 );
    xnor g1760 ( n37063 , n36009 , n33235 );
    and g1761 ( n6848 , n26805 , n42145 );
    and g1762 ( n33275 , n24798 , n906 );
    nor g1763 ( n4608 , n38157 , n19927 );
    nor g1764 ( n40423 , n18909 , n15099 );
    or g1765 ( n4858 , n28647 , n32991 );
    or g1766 ( n28106 , n17105 , n23328 );
    or g1767 ( n4944 , n38879 , n16529 );
    or g1768 ( n1596 , n31634 , n3439 );
    and g1769 ( n6187 , n26125 , n25183 );
    or g1770 ( n26970 , n440 , n25771 );
    not g1771 ( n33774 , n40297 );
    or g1772 ( n5723 , n25526 , n23779 );
    not g1773 ( n29053 , n38504 );
    xnor g1774 ( n19392 , n23902 , n33066 );
    not g1775 ( n25863 , n22526 );
    or g1776 ( n6748 , n4552 , n34542 );
    nor g1777 ( n41499 , n41119 , n13841 );
    and g1778 ( n13238 , n28557 , n20872 );
    xnor g1779 ( n17868 , n14242 , n16748 );
    or g1780 ( n32049 , n6618 , n5328 );
    or g1781 ( n34467 , n7139 , n38518 );
    or g1782 ( n15120 , n8952 , n33488 );
    or g1783 ( n32696 , n37698 , n30045 );
    and g1784 ( n21157 , n21684 , n10105 );
    and g1785 ( n12972 , n25098 , n12023 );
    xnor g1786 ( n22052 , n7503 , n28941 );
    or g1787 ( n695 , n1062 , n27278 );
    and g1788 ( n39332 , n865 , n29623 );
    or g1789 ( n41748 , n40554 , n10529 );
    not g1790 ( n26122 , n2062 );
    and g1791 ( n7111 , n4143 , n2500 );
    nor g1792 ( n23916 , n36112 , n7283 );
    xnor g1793 ( n41683 , n13172 , n7356 );
    and g1794 ( n16851 , n25644 , n32500 );
    xnor g1795 ( n28201 , n32253 , n34023 );
    nor g1796 ( n20742 , n38761 , n13854 );
    xnor g1797 ( n23324 , n29854 , n39967 );
    and g1798 ( n12461 , n7967 , n19920 );
    or g1799 ( n8060 , n40144 , n8442 );
    nor g1800 ( n21778 , n13160 , n15211 );
    or g1801 ( n4524 , n41997 , n15780 );
    xnor g1802 ( n38454 , n784 , n36517 );
    nor g1803 ( n23531 , n19833 , n30500 );
    or g1804 ( n32140 , n37211 , n31999 );
    or g1805 ( n9689 , n2145 , n35574 );
    xnor g1806 ( n27629 , n17891 , n14471 );
    or g1807 ( n25864 , n16431 , n33643 );
    or g1808 ( n24532 , n36815 , n20939 );
    nor g1809 ( n1854 , n29640 , n13318 );
    or g1810 ( n5971 , n37231 , n17709 );
    xnor g1811 ( n18850 , n21973 , n2258 );
    and g1812 ( n3714 , n16051 , n41359 );
    xnor g1813 ( n26146 , n3053 , n7087 );
    or g1814 ( n6186 , n37725 , n41224 );
    xnor g1815 ( n28810 , n32178 , n869 );
    and g1816 ( n36833 , n38640 , n13671 );
    or g1817 ( n24544 , n17984 , n9936 );
    xnor g1818 ( n9014 , n15896 , n36989 );
    or g1819 ( n11083 , n14707 , n14601 );
    and g1820 ( n32818 , n8525 , n534 );
    and g1821 ( n1139 , n24944 , n26842 );
    or g1822 ( n13458 , n39529 , n3034 );
    or g1823 ( n36878 , n1043 , n33330 );
    and g1824 ( n28200 , n20762 , n27469 );
    and g1825 ( n1096 , n26086 , n42555 );
    nor g1826 ( n12685 , n35406 , n18154 );
    or g1827 ( n7976 , n17721 , n33775 );
    not g1828 ( n26627 , n32824 );
    not g1829 ( n27151 , n10891 );
    or g1830 ( n9153 , n9609 , n31503 );
    or g1831 ( n26164 , n35267 , n25089 );
    not g1832 ( n34391 , n20190 );
    or g1833 ( n27293 , n25526 , n14142 );
    nor g1834 ( n36481 , n16780 , n36528 );
    not g1835 ( n19469 , n32716 );
    and g1836 ( n15776 , n11801 , n23428 );
    not g1837 ( n16143 , n26902 );
    and g1838 ( n19442 , n20708 , n33895 );
    or g1839 ( n29736 , n19221 , n26000 );
    and g1840 ( n34131 , n30689 , n26537 );
    or g1841 ( n31047 , n5106 , n31733 );
    and g1842 ( n23888 , n27774 , n36666 );
    or g1843 ( n12131 , n38806 , n38143 );
    xnor g1844 ( n35688 , n18227 , n276 );
    and g1845 ( n22528 , n3987 , n39162 );
    or g1846 ( n10162 , n19994 , n14235 );
    xnor g1847 ( n13118 , n4334 , n38799 );
    not g1848 ( n35356 , n20608 );
    nor g1849 ( n18324 , n34565 , n12676 );
    not g1850 ( n27334 , n4109 );
    or g1851 ( n14783 , n33955 , n28500 );
    or g1852 ( n31567 , n37493 , n34594 );
    or g1853 ( n15603 , n4870 , n7944 );
    xnor g1854 ( n9076 , n23619 , n22761 );
    not g1855 ( n30234 , n26762 );
    and g1856 ( n38822 , n1544 , n3241 );
    or g1857 ( n533 , n20174 , n29604 );
    nor g1858 ( n2660 , n23712 , n7080 );
    or g1859 ( n34852 , n18379 , n40561 );
    or g1860 ( n24124 , n39539 , n9163 );
    nor g1861 ( n22183 , n14091 , n4169 );
    xnor g1862 ( n33512 , n2956 , n33232 );
    not g1863 ( n1201 , n40532 );
    and g1864 ( n20855 , n38365 , n31576 );
    and g1865 ( n8996 , n21241 , n694 );
    or g1866 ( n18632 , n10672 , n19442 );
    nor g1867 ( n10964 , n41352 , n7471 );
    and g1868 ( n41411 , n10746 , n35329 );
    not g1869 ( n33072 , n30776 );
    xnor g1870 ( n1430 , n17377 , n30777 );
    xnor g1871 ( n30415 , n31989 , n5365 );
    not g1872 ( n25016 , n12077 );
    not g1873 ( n5163 , n27860 );
    and g1874 ( n41327 , n22895 , n38370 );
    and g1875 ( n1535 , n24067 , n34668 );
    not g1876 ( n37119 , n29987 );
    or g1877 ( n29920 , n12722 , n41254 );
    or g1878 ( n42294 , n39799 , n13941 );
    nor g1879 ( n5877 , n18866 , n15832 );
    or g1880 ( n9391 , n19753 , n31325 );
    or g1881 ( n6347 , n16479 , n35624 );
    xnor g1882 ( n8358 , n29823 , n4876 );
    and g1883 ( n14321 , n27009 , n6412 );
    and g1884 ( n10899 , n16810 , n24838 );
    or g1885 ( n2627 , n33427 , n32180 );
    or g1886 ( n37476 , n28492 , n13215 );
    and g1887 ( n8344 , n23220 , n22817 );
    not g1888 ( n25474 , n10362 );
    not g1889 ( n19194 , n1490 );
    and g1890 ( n9749 , n16355 , n36366 );
    or g1891 ( n4638 , n41609 , n26416 );
    or g1892 ( n19515 , n19623 , n35370 );
    and g1893 ( n3072 , n41392 , n7110 );
    or g1894 ( n8714 , n4839 , n26806 );
    or g1895 ( n4845 , n28475 , n6325 );
    and g1896 ( n7820 , n18917 , n34283 );
    or g1897 ( n35235 , n28725 , n4580 );
    or g1898 ( n10494 , n7839 , n39902 );
    or g1899 ( n39142 , n42026 , n20684 );
    and g1900 ( n6496 , n9403 , n33848 );
    not g1901 ( n35745 , n20425 );
    and g1902 ( n21628 , n19174 , n3895 );
    or g1903 ( n40181 , n26353 , n42694 );
    or g1904 ( n35053 , n37119 , n5983 );
    xnor g1905 ( n12506 , n36998 , n35818 );
    not g1906 ( n12024 , n31352 );
    xnor g1907 ( n12590 , n14364 , n418 );
    or g1908 ( n4860 , n5348 , n39342 );
    or g1909 ( n182 , n33328 , n15455 );
    nor g1910 ( n38508 , n21724 , n36202 );
    and g1911 ( n41644 , n27076 , n23058 );
    not g1912 ( n38371 , n9331 );
    and g1913 ( n40576 , n18382 , n25805 );
    or g1914 ( n1121 , n4791 , n25142 );
    nor g1915 ( n9125 , n4064 , n40205 );
    or g1916 ( n23415 , n17120 , n27110 );
    or g1917 ( n19274 , n16235 , n27034 );
    or g1918 ( n9309 , n40100 , n4665 );
    not g1919 ( n20190 , n4886 );
    or g1920 ( n6129 , n23509 , n8464 );
    xnor g1921 ( n15447 , n27789 , n26549 );
    or g1922 ( n7022 , n12397 , n7873 );
    or g1923 ( n14903 , n16711 , n12152 );
    or g1924 ( n6801 , n24448 , n42372 );
    or g1925 ( n38834 , n9979 , n11714 );
    or g1926 ( n2340 , n20207 , n14057 );
    nor g1927 ( n23226 , n17120 , n15795 );
    xnor g1928 ( n36208 , n40 , n33705 );
    or g1929 ( n23702 , n14608 , n30140 );
    or g1930 ( n19764 , n39933 , n16988 );
    nor g1931 ( n18023 , n20811 , n18121 );
    nor g1932 ( n42708 , n12327 , n22285 );
    and g1933 ( n7167 , n6251 , n1007 );
    or g1934 ( n14729 , n42231 , n2555 );
    nor g1935 ( n41350 , n17179 , n18920 );
    nor g1936 ( n24867 , n28836 , n9118 );
    nor g1937 ( n25938 , n33790 , n34944 );
    or g1938 ( n40341 , n36806 , n6234 );
    and g1939 ( n3859 , n14185 , n14098 );
    not g1940 ( n25188 , n22647 );
    or g1941 ( n13772 , n14756 , n36565 );
    and g1942 ( n40668 , n12664 , n26304 );
    not g1943 ( n23489 , n26925 );
    nor g1944 ( n34424 , n37616 , n30061 );
    not g1945 ( n10439 , n6826 );
    or g1946 ( n627 , n35301 , n9632 );
    and g1947 ( n5991 , n7509 , n5537 );
    or g1948 ( n4275 , n34130 , n7619 );
    and g1949 ( n26035 , n13350 , n11792 );
    or g1950 ( n31154 , n34315 , n30071 );
    or g1951 ( n17374 , n30197 , n3295 );
    or g1952 ( n14764 , n18663 , n1013 );
    xnor g1953 ( n34035 , n11799 , n13480 );
    or g1954 ( n8323 , n18348 , n33446 );
    or g1955 ( n7138 , n11404 , n40879 );
    or g1956 ( n11486 , n9727 , n22715 );
    nor g1957 ( n22129 , n14471 , n20985 );
    or g1958 ( n3123 , n16564 , n16591 );
    or g1959 ( n11560 , n20449 , n9862 );
    nor g1960 ( n34529 , n18530 , n9965 );
    xnor g1961 ( n8416 , n24265 , n40951 );
    or g1962 ( n10896 , n16195 , n5057 );
    xnor g1963 ( n16377 , n14557 , n36117 );
    or g1964 ( n19901 , n9748 , n30216 );
    not g1965 ( n6503 , n39764 );
    or g1966 ( n20774 , n1374 , n37890 );
    xnor g1967 ( n40962 , n42064 , n17473 );
    or g1968 ( n36100 , n34994 , n6669 );
    not g1969 ( n33261 , n30571 );
    or g1970 ( n39979 , n4565 , n11613 );
    not g1971 ( n34945 , n4822 );
    or g1972 ( n37612 , n18664 , n15387 );
    and g1973 ( n869 , n42818 , n28550 );
    not g1974 ( n40686 , n4999 );
    nor g1975 ( n20510 , n39266 , n39196 );
    or g1976 ( n412 , n15877 , n16341 );
    not g1977 ( n21174 , n40851 );
    or g1978 ( n29729 , n27374 , n19842 );
    or g1979 ( n14355 , n27311 , n11978 );
    not g1980 ( n15730 , n42743 );
    or g1981 ( n33758 , n19196 , n21094 );
    or g1982 ( n30702 , n20404 , n36235 );
    and g1983 ( n13450 , n42739 , n22511 );
    or g1984 ( n31802 , n2885 , n26296 );
    or g1985 ( n16992 , n29697 , n30308 );
    or g1986 ( n31118 , n13418 , n32432 );
    and g1987 ( n37014 , n41408 , n31548 );
    or g1988 ( n27054 , n14223 , n9508 );
    xnor g1989 ( n30065 , n34628 , n42307 );
    or g1990 ( n19912 , n3372 , n17931 );
    nor g1991 ( n39724 , n23325 , n19376 );
    nor g1992 ( n37864 , n33367 , n10495 );
    nor g1993 ( n17212 , n38806 , n32172 );
    or g1994 ( n7078 , n33624 , n4928 );
    not g1995 ( n21296 , n30560 );
    and g1996 ( n26189 , n27399 , n2544 );
    nor g1997 ( n33677 , n4869 , n36659 );
    or g1998 ( n31116 , n328 , n40048 );
    or g1999 ( n42400 , n13371 , n4092 );
    not g2000 ( n28667 , n14206 );
    not g2001 ( n41260 , n23483 );
    xnor g2002 ( n15567 , n13444 , n20722 );
    xnor g2003 ( n3038 , n8489 , n21274 );
    not g2004 ( n25438 , n37615 );
    and g2005 ( n3867 , n1193 , n10968 );
    nor g2006 ( n37869 , n5926 , n29627 );
    or g2007 ( n7186 , n32892 , n37524 );
    or g2008 ( n22526 , n17608 , n18715 );
    not g2009 ( n21899 , n3069 );
    or g2010 ( n34482 , n26512 , n24786 );
    not g2011 ( n18333 , n5846 );
    xnor g2012 ( n25258 , n31989 , n19659 );
    nor g2013 ( n25350 , n2806 , n35953 );
    not g2014 ( n16870 , n20564 );
    xnor g2015 ( n29501 , n34731 , n31979 );
    nor g2016 ( n35584 , n22482 , n27017 );
    not g2017 ( n14265 , n35833 );
    or g2018 ( n546 , n35317 , n28813 );
    xnor g2019 ( n14714 , n13597 , n2865 );
    or g2020 ( n20653 , n23198 , n41913 );
    nor g2021 ( n13937 , n41745 , n17648 );
    or g2022 ( n1333 , n9634 , n1564 );
    or g2023 ( n1562 , n36980 , n17389 );
    or g2024 ( n17822 , n15505 , n42664 );
    xnor g2025 ( n29469 , n11584 , n5267 );
    and g2026 ( n1626 , n5630 , n42203 );
    or g2027 ( n20081 , n10574 , n28419 );
    or g2028 ( n19696 , n10459 , n29258 );
    not g2029 ( n33301 , n35666 );
    or g2030 ( n12966 , n26372 , n40323 );
    or g2031 ( n15859 , n22181 , n26943 );
    or g2032 ( n25618 , n933 , n16614 );
    or g2033 ( n21043 , n35526 , n12968 );
    nor g2034 ( n35847 , n38189 , n18527 );
    or g2035 ( n38890 , n41110 , n41147 );
    or g2036 ( n6414 , n18242 , n16470 );
    not g2037 ( n18928 , n32814 );
    or g2038 ( n10140 , n24114 , n10296 );
    or g2039 ( n29096 , n35301 , n17990 );
    or g2040 ( n32677 , n37348 , n18316 );
    or g2041 ( n3355 , n27449 , n21175 );
    xnor g2042 ( n2283 , n42833 , n1727 );
    and g2043 ( n40480 , n39525 , n42756 );
    or g2044 ( n25866 , n32709 , n18435 );
    nor g2045 ( n11770 , n37086 , n34529 );
    xnor g2046 ( n22342 , n27691 , n19221 );
    nor g2047 ( n5004 , n15608 , n20384 );
    not g2048 ( n6479 , n8117 );
    nor g2049 ( n23246 , n7510 , n242 );
    and g2050 ( n30544 , n4881 , n13076 );
    xnor g2051 ( n10519 , n29740 , n31098 );
    and g2052 ( n21037 , n13118 , n28828 );
    not g2053 ( n37539 , n27308 );
    and g2054 ( n19672 , n10093 , n36361 );
    and g2055 ( n16792 , n11985 , n30433 );
    and g2056 ( n28533 , n34721 , n18092 );
    or g2057 ( n2207 , n31542 , n42105 );
    xnor g2058 ( n21905 , n36394 , n36425 );
    or g2059 ( n1354 , n24790 , n24077 );
    not g2060 ( n3387 , n34053 );
    and g2061 ( n29831 , n8325 , n28460 );
    xnor g2062 ( n25584 , n174 , n25743 );
    and g2063 ( n19750 , n24628 , n22008 );
    or g2064 ( n7162 , n39977 , n28963 );
    not g2065 ( n11847 , n32938 );
    xnor g2066 ( n32764 , n26082 , n41851 );
    and g2067 ( n31975 , n40258 , n34357 );
    or g2068 ( n34714 , n7612 , n4158 );
    not g2069 ( n4750 , n31746 );
    and g2070 ( n39794 , n12936 , n34784 );
    or g2071 ( n27888 , n19744 , n22448 );
    not g2072 ( n36087 , n18637 );
    or g2073 ( n3533 , n24879 , n33248 );
    or g2074 ( n28259 , n16916 , n33806 );
    and g2075 ( n11105 , n4597 , n507 );
    nor g2076 ( n6808 , n14117 , n30554 );
    xnor g2077 ( n27492 , n10043 , n13927 );
    or g2078 ( n1102 , n38346 , n15006 );
    and g2079 ( n8980 , n16177 , n30541 );
    not g2080 ( n11279 , n13902 );
    or g2081 ( n35619 , n30294 , n2565 );
    not g2082 ( n22634 , n26673 );
    and g2083 ( n4098 , n1333 , n12267 );
    or g2084 ( n12974 , n33981 , n34359 );
    or g2085 ( n4398 , n10953 , n11028 );
    or g2086 ( n40134 , n26789 , n15960 );
    nor g2087 ( n31511 , n25461 , n36800 );
    or g2088 ( n1991 , n26387 , n35610 );
    or g2089 ( n10150 , n4552 , n8115 );
    and g2090 ( n40571 , n9623 , n20221 );
    or g2091 ( n7686 , n9184 , n3468 );
    and g2092 ( n41858 , n19946 , n16196 );
    not g2093 ( n2803 , n3945 );
    and g2094 ( n19720 , n7656 , n14106 );
    and g2095 ( n32259 , n42146 , n424 );
    or g2096 ( n40395 , n27879 , n36839 );
    or g2097 ( n11013 , n41519 , n34666 );
    xnor g2098 ( n17431 , n36046 , n2448 );
    or g2099 ( n3566 , n14622 , n38185 );
    not g2100 ( n16264 , n36298 );
    nor g2101 ( n21773 , n18335 , n9725 );
    or g2102 ( n7005 , n819 , n35638 );
    or g2103 ( n3513 , n4414 , n3031 );
    not g2104 ( n13866 , n29117 );
    not g2105 ( n25041 , n34686 );
    xnor g2106 ( n39610 , n11449 , n37984 );
    xnor g2107 ( n24591 , n34352 , n28594 );
    nor g2108 ( n25754 , n11063 , n489 );
    or g2109 ( n12595 , n38704 , n33024 );
    and g2110 ( n20069 , n37227 , n30050 );
    or g2111 ( n37113 , n33776 , n20446 );
    not g2112 ( n38810 , n1804 );
    and g2113 ( n33047 , n15756 , n24174 );
    or g2114 ( n39281 , n15461 , n28312 );
    not g2115 ( n10926 , n27570 );
    not g2116 ( n2616 , n19448 );
    or g2117 ( n31653 , n27323 , n2296 );
    xnor g2118 ( n39809 , n7683 , n5964 );
    not g2119 ( n15717 , n20980 );
    xnor g2120 ( n38917 , n14953 , n39904 );
    or g2121 ( n26866 , n38879 , n25833 );
    and g2122 ( n11273 , n2403 , n23804 );
    or g2123 ( n4434 , n26164 , n9947 );
    xnor g2124 ( n39841 , n20904 , n15596 );
    or g2125 ( n20316 , n12641 , n12244 );
    or g2126 ( n22341 , n19361 , n10802 );
    or g2127 ( n1563 , n12938 , n13238 );
    or g2128 ( n36005 , n3325 , n41413 );
    nor g2129 ( n40634 , n36998 , n21057 );
    or g2130 ( n33153 , n997 , n24374 );
    xnor g2131 ( n11690 , n12007 , n29778 );
    xnor g2132 ( n14782 , n8255 , n41312 );
    xnor g2133 ( n35768 , n27598 , n27130 );
    xnor g2134 ( n27399 , n40886 , n13569 );
    xnor g2135 ( n32262 , n19822 , n37424 );
    or g2136 ( n13608 , n17193 , n37064 );
    not g2137 ( n38899 , n27148 );
    xnor g2138 ( n6353 , n29855 , n38380 );
    or g2139 ( n22315 , n11048 , n1688 );
    xnor g2140 ( n23388 , n14243 , n18451 );
    not g2141 ( n26058 , n5675 );
    or g2142 ( n29620 , n12820 , n33363 );
    not g2143 ( n13677 , n28347 );
    not g2144 ( n24538 , n18730 );
    not g2145 ( n27439 , n30902 );
    not g2146 ( n32893 , n40332 );
    or g2147 ( n11664 , n34561 , n33228 );
    or g2148 ( n7781 , n11495 , n3636 );
    or g2149 ( n2011 , n40259 , n11215 );
    or g2150 ( n1559 , n35915 , n12090 );
    and g2151 ( n7771 , n16405 , n15117 );
    and g2152 ( n20683 , n20385 , n17480 );
    or g2153 ( n33097 , n16839 , n25206 );
    and g2154 ( n31232 , n30146 , n22843 );
    or g2155 ( n35176 , n37207 , n26119 );
    or g2156 ( n40415 , n35294 , n8685 );
    and g2157 ( n33523 , n41636 , n6449 );
    and g2158 ( n32988 , n14509 , n35917 );
    and g2159 ( n24194 , n42602 , n33894 );
    or g2160 ( n12441 , n32479 , n29292 );
    xnor g2161 ( n35849 , n24002 , n16681 );
    xnor g2162 ( n24136 , n18192 , n36849 );
    not g2163 ( n19296 , n8059 );
    not g2164 ( n10475 , n2217 );
    or g2165 ( n37783 , n26052 , n36962 );
    not g2166 ( n41819 , n15396 );
    and g2167 ( n41546 , n23811 , n25921 );
    and g2168 ( n22606 , n41234 , n32234 );
    nor g2169 ( n18707 , n34704 , n29653 );
    and g2170 ( n13188 , n15150 , n27305 );
    and g2171 ( n12627 , n30135 , n33169 );
    xnor g2172 ( n36267 , n6625 , n4987 );
    or g2173 ( n29470 , n15504 , n7016 );
    or g2174 ( n15047 , n36296 , n27945 );
    or g2175 ( n11274 , n29027 , n7094 );
    not g2176 ( n10353 , n6715 );
    and g2177 ( n35094 , n25340 , n39179 );
    or g2178 ( n33579 , n3910 , n36393 );
    or g2179 ( n38699 , n6211 , n32145 );
    or g2180 ( n15938 , n4699 , n1326 );
    or g2181 ( n9623 , n3223 , n32942 );
    and g2182 ( n11583 , n34489 , n12340 );
    and g2183 ( n17166 , n17616 , n42601 );
    and g2184 ( n7751 , n13875 , n24912 );
    xnor g2185 ( n38299 , n23608 , n16707 );
    and g2186 ( n5252 , n8058 , n9605 );
    or g2187 ( n1372 , n37496 , n1013 );
    or g2188 ( n12436 , n1889 , n988 );
    and g2189 ( n16325 , n25955 , n12941 );
    and g2190 ( n18230 , n36886 , n29578 );
    or g2191 ( n838 , n24894 , n38647 );
    or g2192 ( n11710 , n6380 , n25504 );
    and g2193 ( n24899 , n18216 , n9960 );
    xnor g2194 ( n16486 , n36998 , n32919 );
    or g2195 ( n37274 , n2759 , n14487 );
    and g2196 ( n34285 , n22556 , n1973 );
    and g2197 ( n31756 , n3016 , n17878 );
    or g2198 ( n39428 , n3583 , n33378 );
    not g2199 ( n30531 , n38300 );
    xnor g2200 ( n39390 , n18880 , n5952 );
    not g2201 ( n16253 , n1 );
    not g2202 ( n26580 , n21763 );
    or g2203 ( n18161 , n20835 , n24982 );
    nor g2204 ( n14237 , n29395 , n25851 );
    and g2205 ( n240 , n17834 , n13440 );
    or g2206 ( n6778 , n38430 , n7030 );
    nor g2207 ( n10234 , n38955 , n32460 );
    or g2208 ( n41522 , n30407 , n16368 );
    nor g2209 ( n25496 , n4271 , n41985 );
    or g2210 ( n13152 , n39095 , n28901 );
    xnor g2211 ( n8036 , n1841 , n14829 );
    or g2212 ( n33942 , n38996 , n2649 );
    xnor g2213 ( n25190 , n29905 , n20715 );
    or g2214 ( n893 , n39625 , n39408 );
    and g2215 ( n4665 , n14803 , n32838 );
    or g2216 ( n16348 , n29543 , n36256 );
    nor g2217 ( n8419 , n4375 , n12464 );
    and g2218 ( n40689 , n22661 , n28284 );
    or g2219 ( n37001 , n41762 , n36687 );
    xnor g2220 ( n18774 , n4118 , n9094 );
    xnor g2221 ( n21368 , n16320 , n7293 );
    nor g2222 ( n1632 , n33303 , n28106 );
    and g2223 ( n14232 , n11474 , n22857 );
    or g2224 ( n9334 , n16371 , n8728 );
    or g2225 ( n5325 , n1806 , n33698 );
    or g2226 ( n40780 , n6170 , n39459 );
    or g2227 ( n28244 , n32191 , n25728 );
    or g2228 ( n14135 , n18335 , n15143 );
    or g2229 ( n15605 , n21155 , n11423 );
    or g2230 ( n14453 , n7275 , n22885 );
    and g2231 ( n24357 , n1048 , n39136 );
    and g2232 ( n30599 , n19441 , n32840 );
    nor g2233 ( n18167 , n19459 , n27252 );
    xnor g2234 ( n3752 , n22899 , n33410 );
    xnor g2235 ( n22474 , n11434 , n20337 );
    not g2236 ( n29084 , n24479 );
    and g2237 ( n39446 , n8477 , n35851 );
    or g2238 ( n19985 , n6333 , n40259 );
    xnor g2239 ( n53 , n41039 , n33981 );
    not g2240 ( n1419 , n20714 );
    or g2241 ( n18154 , n11573 , n29744 );
    and g2242 ( n41963 , n5815 , n11313 );
    or g2243 ( n4573 , n10836 , n7085 );
    not g2244 ( n2210 , n27655 );
    not g2245 ( n9617 , n20766 );
    xnor g2246 ( n34304 , n41013 , n225 );
    or g2247 ( n39119 , n42447 , n15121 );
    not g2248 ( n23681 , n25025 );
    not g2249 ( n35521 , n23970 );
    not g2250 ( n18146 , n19952 );
    and g2251 ( n29104 , n33215 , n41518 );
    nor g2252 ( n12003 , n11799 , n22517 );
    and g2253 ( n41129 , n37490 , n40969 );
    not g2254 ( n29667 , n25247 );
    and g2255 ( n3679 , n5946 , n11442 );
    or g2256 ( n7554 , n28568 , n34496 );
    xnor g2257 ( n17285 , n27874 , n19986 );
    or g2258 ( n2747 , n5228 , n17026 );
    or g2259 ( n26768 , n26354 , n18668 );
    and g2260 ( n38544 , n20445 , n8443 );
    or g2261 ( n41043 , n14945 , n12744 );
    xnor g2262 ( n22827 , n2753 , n932 );
    or g2263 ( n23379 , n23784 , n3933 );
    nor g2264 ( n40837 , n16598 , n39958 );
    or g2265 ( n10949 , n27871 , n3728 );
    and g2266 ( n25300 , n33490 , n19256 );
    nor g2267 ( n20993 , n30146 , n22843 );
    and g2268 ( n36143 , n40737 , n10588 );
    or g2269 ( n17894 , n29789 , n19958 );
    xnor g2270 ( n12952 , n24442 , n11052 );
    xnor g2271 ( n1431 , n26406 , n31680 );
    not g2272 ( n7363 , n15864 );
    xnor g2273 ( n16185 , n11436 , n2470 );
    xnor g2274 ( n10367 , n36009 , n6949 );
    or g2275 ( n23488 , n19884 , n17606 );
    and g2276 ( n4495 , n31149 , n34928 );
    xnor g2277 ( n26347 , n9079 , n24480 );
    or g2278 ( n22391 , n4099 , n42161 );
    and g2279 ( n18337 , n40159 , n41610 );
    nor g2280 ( n28419 , n37494 , n14184 );
    or g2281 ( n9605 , n8941 , n840 );
    or g2282 ( n9450 , n41560 , n10999 );
    or g2283 ( n26454 , n7847 , n24107 );
    or g2284 ( n7929 , n20754 , n30878 );
    and g2285 ( n26675 , n31034 , n7499 );
    xnor g2286 ( n24332 , n2232 , n6217 );
    or g2287 ( n39618 , n40827 , n12153 );
    and g2288 ( n34048 , n26487 , n522 );
    or g2289 ( n4723 , n25142 , n38233 );
    not g2290 ( n39174 , n366 );
    or g2291 ( n37676 , n12540 , n34278 );
    not g2292 ( n31733 , n39793 );
    and g2293 ( n37718 , n28169 , n14066 );
    and g2294 ( n36651 , n22559 , n22289 );
    or g2295 ( n38961 , n33755 , n16914 );
    or g2296 ( n39074 , n40194 , n42912 );
    or g2297 ( n19101 , n24143 , n18070 );
    and g2298 ( n18541 , n13086 , n41409 );
    nor g2299 ( n29170 , n16237 , n14182 );
    and g2300 ( n41954 , n10131 , n9776 );
    not g2301 ( n37804 , n41206 );
    and g2302 ( n3788 , n17395 , n41083 );
    nor g2303 ( n20781 , n33981 , n12545 );
    and g2304 ( n36184 , n9916 , n5843 );
    and g2305 ( n31748 , n35971 , n15804 );
    or g2306 ( n40738 , n15470 , n31919 );
    xnor g2307 ( n21681 , n32794 , n29069 );
    and g2308 ( n37305 , n16561 , n15240 );
    or g2309 ( n16400 , n37119 , n21976 );
    and g2310 ( n60 , n981 , n35754 );
    and g2311 ( n42497 , n14288 , n14781 );
    not g2312 ( n21765 , n16699 );
    or g2313 ( n14514 , n31097 , n17247 );
    not g2314 ( n14198 , n1561 );
    and g2315 ( n30680 , n36060 , n1675 );
    or g2316 ( n40149 , n3754 , n27540 );
    and g2317 ( n26985 , n26053 , n15193 );
    or g2318 ( n36775 , n7864 , n704 );
    or g2319 ( n31406 , n9451 , n32210 );
    nor g2320 ( n30921 , n5642 , n35602 );
    or g2321 ( n24334 , n8848 , n28371 );
    or g2322 ( n4570 , n1292 , n22436 );
    not g2323 ( n42657 , n36066 );
    xnor g2324 ( n37401 , n16525 , n1563 );
    xnor g2325 ( n14418 , n31989 , n18770 );
    or g2326 ( n16944 , n2155 , n35879 );
    or g2327 ( n411 , n3494 , n18213 );
    nor g2328 ( n27842 , n12016 , n11598 );
    or g2329 ( n18848 , n36976 , n20036 );
    xnor g2330 ( n23298 , n35727 , n12601 );
    xnor g2331 ( n2091 , n24332 , n11334 );
    not g2332 ( n21424 , n32825 );
    not g2333 ( n21297 , n106 );
    and g2334 ( n290 , n17471 , n24865 );
    or g2335 ( n548 , n35879 , n36279 );
    xnor g2336 ( n36028 , n34479 , n22587 );
    or g2337 ( n16173 , n3801 , n10068 );
    not g2338 ( n9240 , n13720 );
    not g2339 ( n39392 , n20889 );
    or g2340 ( n2450 , n27327 , n34267 );
    or g2341 ( n29399 , n14867 , n8745 );
    xnor g2342 ( n37 , n14596 , n16256 );
    not g2343 ( n15301 , n23001 );
    not g2344 ( n26888 , n17406 );
    not g2345 ( n10314 , n5271 );
    nor g2346 ( n24967 , n19221 , n196 );
    or g2347 ( n5483 , n32239 , n19027 );
    nor g2348 ( n3157 , n40347 , n27954 );
    or g2349 ( n38990 , n35034 , n12279 );
    nor g2350 ( n27124 , n773 , n27740 );
    or g2351 ( n33714 , n35093 , n2463 );
    or g2352 ( n289 , n42383 , n35749 );
    or g2353 ( n27475 , n4549 , n42544 );
    and g2354 ( n10488 , n26950 , n31867 );
    nor g2355 ( n16902 , n4447 , n37699 );
    or g2356 ( n9669 , n17361 , n793 );
    and g2357 ( n8621 , n22702 , n29171 );
    or g2358 ( n2604 , n13098 , n116 );
    not g2359 ( n19770 , n33793 );
    or g2360 ( n1571 , n21091 , n32676 );
    nor g2361 ( n41520 , n21571 , n39368 );
    or g2362 ( n29478 , n31326 , n29370 );
    or g2363 ( n38095 , n21604 , n9673 );
    not g2364 ( n18395 , n22777 );
    not g2365 ( n10903 , n40301 );
    xnor g2366 ( n13010 , n10526 , n18177 );
    xnor g2367 ( n1804 , n22263 , n20242 );
    xnor g2368 ( n7190 , n11434 , n31530 );
    or g2369 ( n27600 , n2000 , n26927 );
    and g2370 ( n34179 , n25028 , n14536 );
    xnor g2371 ( n8354 , n751 , n40760 );
    or g2372 ( n35408 , n1987 , n14306 );
    not g2373 ( n20274 , n28653 );
    not g2374 ( n9200 , n5351 );
    xnor g2375 ( n1912 , n13444 , n2454 );
    nor g2376 ( n29326 , n18401 , n27135 );
    or g2377 ( n38452 , n33981 , n17620 );
    xnor g2378 ( n23177 , n22556 , n1973 );
    nor g2379 ( n16753 , n25447 , n22205 );
    nor g2380 ( n38663 , n9843 , n30018 );
    and g2381 ( n33539 , n22374 , n16360 );
    and g2382 ( n4510 , n18322 , n23175 );
    not g2383 ( n17299 , n19407 );
    or g2384 ( n22838 , n39047 , n7728 );
    or g2385 ( n42788 , n15569 , n33271 );
    not g2386 ( n40127 , n23504 );
    or g2387 ( n25313 , n20852 , n27450 );
    or g2388 ( n30808 , n36974 , n19290 );
    and g2389 ( n32762 , n22572 , n38482 );
    not g2390 ( n17984 , n22310 );
    or g2391 ( n42807 , n8024 , n22823 );
    xnor g2392 ( n4104 , n12836 , n31482 );
    xnor g2393 ( n41285 , n28614 , n40102 );
    or g2394 ( n28895 , n7061 , n8626 );
    or g2395 ( n5010 , n8301 , n25559 );
    nor g2396 ( n19603 , n22458 , n13284 );
    and g2397 ( n38547 , n42438 , n32903 );
    or g2398 ( n42053 , n40978 , n38833 );
    or g2399 ( n32909 , n8004 , n41902 );
    or g2400 ( n10972 , n2156 , n11373 );
    or g2401 ( n25369 , n10879 , n5124 );
    and g2402 ( n32973 , n42129 , n15016 );
    not g2403 ( n3334 , n19248 );
    or g2404 ( n7982 , n12059 , n27974 );
    and g2405 ( n26093 , n4696 , n10214 );
    and g2406 ( n39905 , n2274 , n11587 );
    not g2407 ( n4345 , n8949 );
    or g2408 ( n41606 , n12966 , n18249 );
    not g2409 ( n35766 , n34014 );
    not g2410 ( n38325 , n14058 );
    nor g2411 ( n21129 , n25384 , n9976 );
    not g2412 ( n28634 , n32476 );
    or g2413 ( n21463 , n1588 , n229 );
    and g2414 ( n14236 , n42587 , n261 );
    or g2415 ( n6926 , n34843 , n30992 );
    or g2416 ( n26047 , n9376 , n13285 );
    or g2417 ( n12384 , n4115 , n30222 );
    xnor g2418 ( n22038 , n13509 , n39266 );
    xnor g2419 ( n16158 , n38173 , n18593 );
    or g2420 ( n33340 , n19811 , n5889 );
    and g2421 ( n41431 , n37370 , n2886 );
    not g2422 ( n15169 , n33731 );
    not g2423 ( n19067 , n41357 );
    nor g2424 ( n42901 , n35439 , n14789 );
    nor g2425 ( n18664 , n42340 , n24271 );
    nor g2426 ( n1038 , n7461 , n3733 );
    or g2427 ( n33045 , n7839 , n12665 );
    xnor g2428 ( n144 , n33184 , n42902 );
    or g2429 ( n15273 , n22122 , n17199 );
    not g2430 ( n37643 , n19651 );
    xnor g2431 ( n27287 , n27423 , n32626 );
    and g2432 ( n24783 , n15221 , n13270 );
    or g2433 ( n1471 , n17120 , n10168 );
    and g2434 ( n3270 , n42587 , n23829 );
    or g2435 ( n24051 , n12499 , n35068 );
    xnor g2436 ( n37644 , n21877 , n15973 );
    and g2437 ( n15519 , n9705 , n29491 );
    or g2438 ( n30624 , n18837 , n13566 );
    not g2439 ( n17481 , n26877 );
    or g2440 ( n29072 , n2609 , n6516 );
    or g2441 ( n15656 , n32683 , n5369 );
    or g2442 ( n10495 , n31405 , n12062 );
    nor g2443 ( n22221 , n16952 , n35306 );
    or g2444 ( n5118 , n23990 , n42017 );
    or g2445 ( n36118 , n6734 , n13176 );
    or g2446 ( n37443 , n38416 , n32771 );
    or g2447 ( n31588 , n4557 , n10080 );
    or g2448 ( n29797 , n28524 , n34569 );
    nor g2449 ( n1569 , n12155 , n20104 );
    or g2450 ( n26775 , n19891 , n25393 );
    and g2451 ( n38061 , n926 , n16085 );
    or g2452 ( n30480 , n10598 , n8178 );
    xnor g2453 ( n42728 , n16742 , n38492 );
    or g2454 ( n24796 , n6053 , n19890 );
    nor g2455 ( n6387 , n36918 , n27559 );
    and g2456 ( n30428 , n36622 , n42879 );
    not g2457 ( n19804 , n37526 );
    xnor g2458 ( n42002 , n6625 , n15313 );
    nor g2459 ( n13163 , n36093 , n31587 );
    not g2460 ( n32558 , n21975 );
    xnor g2461 ( n33458 , n5144 , n23224 );
    and g2462 ( n23632 , n10470 , n32438 );
    not g2463 ( n11614 , n26620 );
    or g2464 ( n8134 , n18441 , n2034 );
    not g2465 ( n27572 , n38263 );
    xnor g2466 ( n7497 , n1664 , n25356 );
    not g2467 ( n11136 , n22816 );
    or g2468 ( n32511 , n40269 , n40325 );
    or g2469 ( n9531 , n32605 , n42295 );
    xnor g2470 ( n4482 , n11380 , n20760 );
    or g2471 ( n34025 , n3920 , n19637 );
    or g2472 ( n3284 , n9961 , n22983 );
    or g2473 ( n17811 , n9785 , n38183 );
    or g2474 ( n39109 , n39133 , n3276 );
    and g2475 ( n25516 , n26373 , n42632 );
    and g2476 ( n33103 , n34417 , n16835 );
    and g2477 ( n29607 , n822 , n10868 );
    or g2478 ( n13385 , n37402 , n17104 );
    and g2479 ( n23522 , n24065 , n21541 );
    or g2480 ( n39321 , n34809 , n35253 );
    or g2481 ( n35067 , n39939 , n4301 );
    or g2482 ( n26527 , n38556 , n36040 );
    or g2483 ( n41017 , n981 , n38130 );
    or g2484 ( n24057 , n28458 , n32359 );
    nor g2485 ( n35226 , n8904 , n911 );
    not g2486 ( n37868 , n25592 );
    or g2487 ( n17231 , n3071 , n3410 );
    nor g2488 ( n26161 , n39449 , n122 );
    or g2489 ( n6167 , n20503 , n39299 );
    not g2490 ( n30075 , n37576 );
    or g2491 ( n619 , n268 , n10786 );
    and g2492 ( n29730 , n3400 , n25332 );
    or g2493 ( n7458 , n13475 , n38025 );
    or g2494 ( n33552 , n23350 , n41259 );
    or g2495 ( n27362 , n30212 , n19890 );
    or g2496 ( n2927 , n31288 , n38211 );
    nor g2497 ( n35319 , n39927 , n1418 );
    or g2498 ( n29154 , n23517 , n8116 );
    or g2499 ( n29694 , n7540 , n27351 );
    nor g2500 ( n34733 , n24064 , n6838 );
    nor g2501 ( n30190 , n4040 , n37535 );
    nor g2502 ( n30999 , n654 , n15022 );
    or g2503 ( n32431 , n36954 , n35608 );
    or g2504 ( n1465 , n20296 , n4884 );
    xnor g2505 ( n37452 , n29740 , n2811 );
    or g2506 ( n41095 , n38879 , n27675 );
    or g2507 ( n30951 , n34687 , n28345 );
    and g2508 ( n8128 , n7858 , n22939 );
    and g2509 ( n5092 , n249 , n1433 );
    not g2510 ( n10072 , n7125 );
    not g2511 ( n33706 , n34933 );
    or g2512 ( n40376 , n7376 , n1207 );
    not g2513 ( n20706 , n29899 );
    or g2514 ( n27604 , n7188 , n15406 );
    and g2515 ( n42561 , n16720 , n19939 );
    or g2516 ( n37386 , n21703 , n6990 );
    and g2517 ( n13662 , n3820 , n8357 );
    not g2518 ( n22175 , n21306 );
    xnor g2519 ( n16847 , n16745 , n2649 );
    or g2520 ( n10735 , n22491 , n37598 );
    or g2521 ( n18124 , n35261 , n24327 );
    not g2522 ( n20980 , n2093 );
    and g2523 ( n31382 , n24853 , n20736 );
    nor g2524 ( n30437 , n33617 , n6035 );
    or g2525 ( n8211 , n16680 , n6216 );
    not g2526 ( n20972 , n2857 );
    and g2527 ( n4631 , n10541 , n2447 );
    or g2528 ( n1810 , n33815 , n27548 );
    or g2529 ( n18636 , n32245 , n30032 );
    or g2530 ( n2941 , n28778 , n23081 );
    or g2531 ( n13789 , n34475 , n10698 );
    nor g2532 ( n18157 , n18212 , n14905 );
    or g2533 ( n27571 , n17153 , n41767 );
    not g2534 ( n27718 , n10208 );
    nor g2535 ( n38113 , n1941 , n25692 );
    not g2536 ( n23170 , n13301 );
    xnor g2537 ( n23581 , n22776 , n5605 );
    or g2538 ( n35785 , n4700 , n4108 );
    and g2539 ( n38740 , n25465 , n7556 );
    and g2540 ( n22914 , n30760 , n42605 );
    xnor g2541 ( n18967 , n15823 , n20196 );
    not g2542 ( n2705 , n25916 );
    or g2543 ( n16413 , n14299 , n25251 );
    or g2544 ( n22237 , n18608 , n30669 );
    nor g2545 ( n19913 , n19602 , n14836 );
    or g2546 ( n4691 , n36295 , n22395 );
    or g2547 ( n12357 , n20092 , n33014 );
    not g2548 ( n12158 , n2735 );
    not g2549 ( n12431 , n19033 );
    or g2550 ( n11357 , n6628 , n20476 );
    or g2551 ( n15034 , n16191 , n6415 );
    xnor g2552 ( n24258 , n25042 , n16912 );
    not g2553 ( n25064 , n41700 );
    xnor g2554 ( n23482 , n39532 , n10804 );
    not g2555 ( n2372 , n30738 );
    or g2556 ( n19801 , n16590 , n17339 );
    not g2557 ( n37919 , n18429 );
    not g2558 ( n18090 , n25853 );
    xnor g2559 ( n37295 , n34235 , n20748 );
    or g2560 ( n12714 , n18847 , n29322 );
    or g2561 ( n31631 , n34994 , n5653 );
    xnor g2562 ( n6934 , n29740 , n29842 );
    nor g2563 ( n18015 , n29717 , n38435 );
    and g2564 ( n24812 , n25871 , n17007 );
    not g2565 ( n14806 , n5147 );
    not g2566 ( n28447 , n19364 );
    and g2567 ( n41639 , n32275 , n31455 );
    xnor g2568 ( n18220 , n19547 , n28989 );
    not g2569 ( n13707 , n39366 );
    nor g2570 ( n22358 , n11646 , n2925 );
    xnor g2571 ( n17762 , n37083 , n36417 );
    not g2572 ( n17909 , n22954 );
    nor g2573 ( n36264 , n6558 , n13930 );
    and g2574 ( n29290 , n34616 , n28791 );
    not g2575 ( n27477 , n28326 );
    nor g2576 ( n22732 , n17744 , n1334 );
    not g2577 ( n14776 , n15439 );
    not g2578 ( n39082 , n9116 );
    xnor g2579 ( n40064 , n38685 , n6464 );
    not g2580 ( n9460 , n402 );
    xnor g2581 ( n12816 , n38101 , n12865 );
    or g2582 ( n12422 , n12677 , n9160 );
    or g2583 ( n9788 , n19811 , n33903 );
    or g2584 ( n2709 , n23381 , n10857 );
    not g2585 ( n42648 , n39087 );
    and g2586 ( n27548 , n22215 , n5300 );
    not g2587 ( n8345 , n31189 );
    or g2588 ( n4383 , n27918 , n3036 );
    not g2589 ( n9155 , n41603 );
    or g2590 ( n5737 , n17144 , n19111 );
    or g2591 ( n6071 , n37008 , n29525 );
    and g2592 ( n14019 , n25898 , n8072 );
    or g2593 ( n16353 , n23809 , n15335 );
    not g2594 ( n6544 , n1883 );
    xnor g2595 ( n32517 , n26579 , n7256 );
    and g2596 ( n4781 , n14786 , n34355 );
    xnor g2597 ( n36224 , n16573 , n41258 );
    or g2598 ( n2729 , n39149 , n2149 );
    or g2599 ( n33610 , n2510 , n40556 );
    or g2600 ( n93 , n16996 , n13145 );
    not g2601 ( n40086 , n21710 );
    nor g2602 ( n17832 , n6038 , n5988 );
    and g2603 ( n10008 , n23851 , n29374 );
    nor g2604 ( n19863 , n1371 , n2428 );
    not g2605 ( n9264 , n32094 );
    and g2606 ( n34511 , n15515 , n19959 );
    or g2607 ( n28762 , n23739 , n31914 );
    and g2608 ( n3767 , n34065 , n15067 );
    or g2609 ( n1482 , n21752 , n33923 );
    nor g2610 ( n3469 , n36345 , n35993 );
    nor g2611 ( n42600 , n30818 , n15607 );
    and g2612 ( n42374 , n23902 , n34380 );
    or g2613 ( n31191 , n14707 , n20831 );
    not g2614 ( n36880 , n25649 );
    nor g2615 ( n20611 , n3893 , n35728 );
    or g2616 ( n23441 , n6362 , n27042 );
    and g2617 ( n10837 , n37272 , n21518 );
    or g2618 ( n29086 , n10771 , n27176 );
    not g2619 ( n13701 , n40674 );
    or g2620 ( n33117 , n33556 , n239 );
    or g2621 ( n12593 , n27798 , n7837 );
    xnor g2622 ( n29450 , n14758 , n34495 );
    not g2623 ( n17070 , n7785 );
    nor g2624 ( n33615 , n35310 , n4630 );
    not g2625 ( n13981 , n12144 );
    or g2626 ( n8931 , n41699 , n12915 );
    not g2627 ( n32367 , n29660 );
    not g2628 ( n35274 , n40781 );
    and g2629 ( n42131 , n25884 , n6784 );
    xnor g2630 ( n32528 , n2182 , n4550 );
    nor g2631 ( n8752 , n27786 , n23138 );
    or g2632 ( n34753 , n19769 , n27107 );
    and g2633 ( n22833 , n14876 , n20284 );
    nor g2634 ( n38017 , n31096 , n31570 );
    not g2635 ( n32485 , n4208 );
    and g2636 ( n18542 , n27597 , n3365 );
    or g2637 ( n16468 , n41534 , n26281 );
    or g2638 ( n39654 , n26707 , n11001 );
    or g2639 ( n25117 , n28205 , n20867 );
    and g2640 ( n9574 , n16435 , n14533 );
    and g2641 ( n25356 , n2605 , n3827 );
    or g2642 ( n25495 , n13367 , n15963 );
    or g2643 ( n873 , n12392 , n18156 );
    or g2644 ( n41693 , n25078 , n35616 );
    or g2645 ( n37196 , n17360 , n18352 );
    not g2646 ( n21888 , n20553 );
    and g2647 ( n39589 , n11277 , n42807 );
    or g2648 ( n5184 , n5643 , n28208 );
    or g2649 ( n33004 , n14471 , n17891 );
    not g2650 ( n2009 , n4023 );
    xnor g2651 ( n23549 , n16693 , n1177 );
    and g2652 ( n36405 , n5030 , n30196 );
    nor g2653 ( n18627 , n24898 , n10249 );
    nor g2654 ( n8755 , n16730 , n4483 );
    nor g2655 ( n30525 , n41534 , n36494 );
    or g2656 ( n25049 , n16586 , n27122 );
    not g2657 ( n21918 , n24737 );
    xnor g2658 ( n38450 , n28299 , n29873 );
    or g2659 ( n2201 , n31452 , n36707 );
    not g2660 ( n24825 , n40387 );
    not g2661 ( n19365 , n35291 );
    or g2662 ( n36276 , n40645 , n3009 );
    and g2663 ( n41586 , n41256 , n5544 );
    nor g2664 ( n8362 , n12261 , n16555 );
    or g2665 ( n40758 , n40437 , n10491 );
    not g2666 ( n11640 , n21870 );
    not g2667 ( n17724 , n9671 );
    and g2668 ( n13980 , n31236 , n40905 );
    nor g2669 ( n25087 , n40298 , n14882 );
    or g2670 ( n31507 , n20684 , n11752 );
    and g2671 ( n24638 , n11840 , n9688 );
    or g2672 ( n8481 , n10562 , n12484 );
    not g2673 ( n39140 , n16041 );
    or g2674 ( n18992 , n36037 , n9617 );
    or g2675 ( n35425 , n21312 , n27039 );
    xnor g2676 ( n15340 , n17154 , n19944 );
    or g2677 ( n5756 , n37368 , n24254 );
    not g2678 ( n18051 , n27766 );
    and g2679 ( n25001 , n30539 , n14938 );
    or g2680 ( n3969 , n9971 , n42379 );
    or g2681 ( n30387 , n5716 , n28249 );
    or g2682 ( n24946 , n18475 , n27910 );
    or g2683 ( n5359 , n33464 , n1892 );
    or g2684 ( n5003 , n1689 , n34999 );
    xnor g2685 ( n41241 , n22888 , n10531 );
    not g2686 ( n14692 , n30651 );
    or g2687 ( n16555 , n35438 , n10077 );
    or g2688 ( n30633 , n3562 , n33775 );
    and g2689 ( n8038 , n7890 , n9679 );
    and g2690 ( n25133 , n32924 , n16448 );
    nor g2691 ( n23296 , n2199 , n18426 );
    and g2692 ( n15167 , n14333 , n8838 );
    or g2693 ( n26254 , n7710 , n3715 );
    nor g2694 ( n12191 , n32336 , n21008 );
    or g2695 ( n16475 , n10569 , n12345 );
    xnor g2696 ( n19499 , n16745 , n13130 );
    or g2697 ( n34897 , n22589 , n37787 );
    xnor g2698 ( n17343 , n2130 , n21761 );
    or g2699 ( n1323 , n3764 , n23521 );
    nor g2700 ( n32362 , n32407 , n18051 );
    or g2701 ( n19761 , n11146 , n4474 );
    not g2702 ( n34195 , n19002 );
    nor g2703 ( n13438 , n18866 , n19450 );
    or g2704 ( n40614 , n32008 , n28921 );
    or g2705 ( n16347 , n42490 , n22518 );
    xnor g2706 ( n37489 , n34731 , n9936 );
    and g2707 ( n10998 , n14772 , n9112 );
    nor g2708 ( n5465 , n1186 , n42462 );
    xnor g2709 ( n14797 , n3435 , n1079 );
    not g2710 ( n40457 , n21595 );
    or g2711 ( n3647 , n2008 , n41577 );
    or g2712 ( n37532 , n33755 , n3971 );
    xnor g2713 ( n4168 , n17225 , n17126 );
    or g2714 ( n18615 , n24771 , n28046 );
    nor g2715 ( n5115 , n6548 , n38344 );
    not g2716 ( n29711 , n4432 );
    or g2717 ( n33868 , n15952 , n33655 );
    xnor g2718 ( n31877 , n15842 , n15448 );
    and g2719 ( n5195 , n41946 , n27199 );
    nor g2720 ( n28856 , n39060 , n37875 );
    xnor g2721 ( n14989 , n42064 , n4599 );
    and g2722 ( n33543 , n14605 , n17652 );
    nor g2723 ( n2882 , n5810 , n11610 );
    or g2724 ( n5209 , n34637 , n23659 );
    or g2725 ( n4849 , n15681 , n5437 );
    or g2726 ( n18198 , n32100 , n34679 );
    and g2727 ( n2583 , n37738 , n1851 );
    or g2728 ( n16580 , n14707 , n3910 );
    and g2729 ( n31629 , n3665 , n23524 );
    nor g2730 ( n32749 , n40108 , n5955 );
    nor g2731 ( n16971 , n11679 , n34789 );
    or g2732 ( n334 , n27388 , n32991 );
    nor g2733 ( n10961 , n4290 , n3344 );
    and g2734 ( n14733 , n3765 , n33131 );
    or g2735 ( n18388 , n15852 , n32194 );
    or g2736 ( n1236 , n37938 , n2994 );
    or g2737 ( n26356 , n13149 , n33085 );
    nor g2738 ( n24515 , n23868 , n38797 );
    not g2739 ( n35887 , n30684 );
    and g2740 ( n28921 , n30495 , n25763 );
    not g2741 ( n4435 , n36704 );
    not g2742 ( n37306 , n21515 );
    or g2743 ( n29029 , n36979 , n2939 );
    nor g2744 ( n27976 , n29567 , n2458 );
    not g2745 ( n37806 , n4206 );
    xnor g2746 ( n33509 , n842 , n4964 );
    not g2747 ( n35231 , n41641 );
    or g2748 ( n200 , n22543 , n20296 );
    and g2749 ( n35303 , n6758 , n35785 );
    not g2750 ( n34997 , n27188 );
    and g2751 ( n17502 , n1878 , n4426 );
    or g2752 ( n2374 , n14192 , n8360 );
    or g2753 ( n34696 , n12456 , n40471 );
    or g2754 ( n28587 , n14287 , n28924 );
    and g2755 ( n41387 , n14150 , n10948 );
    nor g2756 ( n28805 , n36595 , n23668 );
    and g2757 ( n26079 , n6167 , n18226 );
    or g2758 ( n33201 , n22037 , n9548 );
    xnor g2759 ( n22918 , n42064 , n24194 );
    nor g2760 ( n17072 , n35039 , n27413 );
    not g2761 ( n24574 , n13219 );
    or g2762 ( n11836 , n1902 , n26482 );
    xnor g2763 ( n9371 , n17137 , n34965 );
    and g2764 ( n32 , n11171 , n19426 );
    or g2765 ( n41436 , n27923 , n12051 );
    or g2766 ( n40165 , n11374 , n6716 );
    or g2767 ( n37670 , n14591 , n10784 );
    or g2768 ( n8839 , n8786 , n15511 );
    or g2769 ( n14230 , n7172 , n23924 );
    not g2770 ( n37633 , n26655 );
    or g2771 ( n34306 , n42904 , n33264 );
    or g2772 ( n29225 , n16893 , n6883 );
    not g2773 ( n37098 , n35522 );
    not g2774 ( n18677 , n17378 );
    nor g2775 ( n20241 , n29004 , n32899 );
    xnor g2776 ( n32328 , n41013 , n20100 );
    or g2777 ( n36935 , n19366 , n6946 );
    xnor g2778 ( n30410 , n14601 , n14707 );
    and g2779 ( n19965 , n27093 , n4957 );
    and g2780 ( n23500 , n7671 , n8930 );
    not g2781 ( n12591 , n41186 );
    not g2782 ( n36046 , n13054 );
    or g2783 ( n34758 , n39330 , n4028 );
    xnor g2784 ( n9307 , n34352 , n41887 );
    nor g2785 ( n15341 , n7621 , n11688 );
    and g2786 ( n23586 , n37046 , n18195 );
    not g2787 ( n8825 , n33106 );
    or g2788 ( n14423 , n27643 , n26740 );
    and g2789 ( n37186 , n6964 , n33000 );
    and g2790 ( n11860 , n14400 , n5593 );
    xnor g2791 ( n34783 , n33917 , n15918 );
    or g2792 ( n16155 , n40108 , n28488 );
    or g2793 ( n9310 , n26287 , n8700 );
    nor g2794 ( n910 , n30066 , n32828 );
    or g2795 ( n20675 , n31265 , n13303 );
    nor g2796 ( n15333 , n23260 , n38652 );
    not g2797 ( n25777 , n14394 );
    not g2798 ( n33621 , n1252 );
    nor g2799 ( n31789 , n22695 , n13084 );
    not g2800 ( n18550 , n42554 );
    nor g2801 ( n6264 , n13659 , n24141 );
    or g2802 ( n40646 , n25573 , n25852 );
    and g2803 ( n22010 , n15994 , n24985 );
    and g2804 ( n18197 , n5191 , n42788 );
    or g2805 ( n21810 , n746 , n27712 );
    or g2806 ( n19098 , n30652 , n17008 );
    nor g2807 ( n16093 , n27627 , n25488 );
    or g2808 ( n11720 , n30674 , n10172 );
    or g2809 ( n18503 , n23242 , n11537 );
    not g2810 ( n12210 , n23168 );
    not g2811 ( n39757 , n28595 );
    or g2812 ( n40084 , n15384 , n28421 );
    or g2813 ( n24850 , n3165 , n39558 );
    xnor g2814 ( n1935 , n35938 , n8155 );
    xnor g2815 ( n38972 , n36009 , n9798 );
    xnor g2816 ( n2947 , n17563 , n24782 );
    or g2817 ( n12862 , n39207 , n729 );
    and g2818 ( n5071 , n17378 , n39675 );
    or g2819 ( n35905 , n3593 , n360 );
    not g2820 ( n20727 , n29169 );
    xnor g2821 ( n36800 , n2205 , n35149 );
    xnor g2822 ( n7454 , n8428 , n2264 );
    or g2823 ( n38116 , n5132 , n39168 );
    or g2824 ( n33240 , n1068 , n4553 );
    or g2825 ( n34600 , n555 , n36393 );
    xnor g2826 ( n37464 , n12524 , n2380 );
    xnor g2827 ( n36749 , n4304 , n7665 );
    and g2828 ( n31095 , n41044 , n19408 );
    or g2829 ( n23845 , n4193 , n39085 );
    and g2830 ( n593 , n20282 , n36637 );
    xnor g2831 ( n9530 , n19231 , n27262 );
    or g2832 ( n39212 , n10835 , n18575 );
    xnor g2833 ( n1232 , n15467 , n28651 );
    or g2834 ( n36048 , n1096 , n35569 );
    or g2835 ( n34851 , n5701 , n40116 );
    xnor g2836 ( n26581 , n37309 , n29172 );
    or g2837 ( n4384 , n20092 , n32169 );
    and g2838 ( n30113 , n7929 , n16524 );
    and g2839 ( n31370 , n18410 , n36489 );
    nor g2840 ( n6655 , n15403 , n7031 );
    not g2841 ( n29110 , n34450 );
    or g2842 ( n565 , n27311 , n31720 );
    xnor g2843 ( n3799 , n41747 , n18400 );
    and g2844 ( n37072 , n28338 , n1869 );
    and g2845 ( n14618 , n12444 , n2810 );
    or g2846 ( n18384 , n10180 , n27179 );
    not g2847 ( n2758 , n11619 );
    or g2848 ( n32279 , n7339 , n14982 );
    or g2849 ( n37472 , n13629 , n11708 );
    not g2850 ( n10600 , n4806 );
    not g2851 ( n13918 , n18941 );
    and g2852 ( n18837 , n14816 , n8343 );
    or g2853 ( n13206 , n40728 , n2545 );
    not g2854 ( n6257 , n23586 );
    or g2855 ( n28278 , n13868 , n35682 );
    nor g2856 ( n19894 , n26341 , n35527 );
    xnor g2857 ( n206 , n23918 , n858 );
    not g2858 ( n15315 , n7798 );
    and g2859 ( n39939 , n18684 , n18768 );
    and g2860 ( n15082 , n2081 , n21226 );
    nor g2861 ( n10077 , n27733 , n17317 );
    or g2862 ( n39937 , n25779 , n14622 );
    nor g2863 ( n28524 , n34582 , n28054 );
    or g2864 ( n32836 , n19183 , n9692 );
    nor g2865 ( n14755 , n8194 , n33427 );
    or g2866 ( n14536 , n24621 , n35090 );
    or g2867 ( n32307 , n39292 , n15333 );
    nor g2868 ( n27411 , n28170 , n34156 );
    and g2869 ( n23148 , n42282 , n38728 );
    or g2870 ( n4476 , n39752 , n36944 );
    xnor g2871 ( n16051 , n7961 , n39266 );
    not g2872 ( n32589 , n6790 );
    or g2873 ( n17470 , n1321 , n22984 );
    nor g2874 ( n10512 , n13921 , n41097 );
    xnor g2875 ( n4443 , n40 , n41032 );
    or g2876 ( n11916 , n35772 , n14093 );
    xnor g2877 ( n18626 , n21415 , n23077 );
    nor g2878 ( n36301 , n1339 , n20408 );
    or g2879 ( n29398 , n6254 , n3715 );
    not g2880 ( n21286 , n42338 );
    or g2881 ( n31594 , n1720 , n14398 );
    xnor g2882 ( n7782 , n25884 , n21947 );
    nor g2883 ( n10546 , n21351 , n1166 );
    or g2884 ( n13876 , n9461 , n15564 );
    or g2885 ( n15259 , n35333 , n5244 );
    or g2886 ( n19520 , n657 , n15780 );
    or g2887 ( n10382 , n12522 , n25305 );
    xnor g2888 ( n10464 , n34564 , n27620 );
    and g2889 ( n22956 , n39599 , n24069 );
    and g2890 ( n42414 , n7234 , n15119 );
    and g2891 ( n323 , n27386 , n34598 );
    or g2892 ( n1514 , n3106 , n15134 );
    not g2893 ( n35557 , n1593 );
    and g2894 ( n23423 , n11214 , n41330 );
    nor g2895 ( n10341 , n5401 , n42169 );
    nor g2896 ( n2288 , n36486 , n2793 );
    not g2897 ( n16121 , n5855 );
    or g2898 ( n3244 , n32685 , n19627 );
    nor g2899 ( n2142 , n22109 , n15751 );
    or g2900 ( n24655 , n17797 , n33020 );
    or g2901 ( n25366 , n26681 , n38176 );
    and g2902 ( n6483 , n10281 , n39649 );
    not g2903 ( n17015 , n5875 );
    or g2904 ( n9519 , n37520 , n9641 );
    or g2905 ( n28094 , n32277 , n21002 );
    and g2906 ( n9524 , n37596 , n22198 );
    nor g2907 ( n13067 , n8400 , n8672 );
    and g2908 ( n25077 , n4253 , n33202 );
    and g2909 ( n37438 , n23345 , n7304 );
    xnor g2910 ( n35246 , n4341 , n6073 );
    not g2911 ( n6675 , n14585 );
    or g2912 ( n9786 , n7039 , n10184 );
    or g2913 ( n8882 , n4538 , n18399 );
    or g2914 ( n34820 , n19879 , n27683 );
    or g2915 ( n18887 , n24153 , n31556 );
    or g2916 ( n24089 , n9177 , n23602 );
    and g2917 ( n15409 , n6940 , n11736 );
    or g2918 ( n30650 , n21025 , n40473 );
    nor g2919 ( n18420 , n4677 , n11017 );
    nor g2920 ( n28393 , n2455 , n27115 );
    and g2921 ( n37408 , n12870 , n33932 );
    nor g2922 ( n35143 , n14707 , n6126 );
    xnor g2923 ( n12047 , n2161 , n5595 );
    not g2924 ( n12305 , n28114 );
    and g2925 ( n11208 , n17743 , n1596 );
    and g2926 ( n16060 , n34507 , n37602 );
    not g2927 ( n26927 , n32271 );
    nor g2928 ( n5692 , n18395 , n32873 );
    or g2929 ( n37350 , n24625 , n19707 );
    nor g2930 ( n19559 , n22072 , n33428 );
    and g2931 ( n6492 , n37000 , n13705 );
    and g2932 ( n42510 , n27073 , n16153 );
    or g2933 ( n4116 , n11033 , n42405 );
    or g2934 ( n2397 , n31168 , n33330 );
    or g2935 ( n9534 , n30235 , n30092 );
    not g2936 ( n3136 , n23165 );
    nor g2937 ( n35296 , n6175 , n39116 );
    nor g2938 ( n14610 , n36117 , n1738 );
    nor g2939 ( n23939 , n38406 , n3344 );
    and g2940 ( n15722 , n39331 , n33846 );
    nor g2941 ( n35346 , n15070 , n28130 );
    nor g2942 ( n42378 , n11847 , n12607 );
    and g2943 ( n14917 , n11300 , n5873 );
    or g2944 ( n42717 , n32245 , n22149 );
    and g2945 ( n3240 , n14878 , n17271 );
    or g2946 ( n13510 , n25505 , n23109 );
    not g2947 ( n26596 , n6456 );
    or g2948 ( n39631 , n14317 , n12867 );
    or g2949 ( n3197 , n40170 , n7414 );
    xnor g2950 ( n8222 , n443 , n31082 );
    xnor g2951 ( n26651 , n25655 , n13522 );
    or g2952 ( n21988 , n5896 , n20100 );
    or g2953 ( n35248 , n35473 , n34648 );
    or g2954 ( n1593 , n15937 , n16814 );
    nor g2955 ( n22154 , n37695 , n23303 );
    nor g2956 ( n444 , n3633 , n1250 );
    nor g2957 ( n23163 , n35678 , n37340 );
    or g2958 ( n30100 , n30737 , n39022 );
    and g2959 ( n29919 , n13405 , n24118 );
    or g2960 ( n33183 , n14493 , n19480 );
    or g2961 ( n3887 , n25451 , n29320 );
    not g2962 ( n21029 , n32520 );
    not g2963 ( n41718 , n10748 );
    or g2964 ( n4189 , n42896 , n1649 );
    or g2965 ( n41959 , n18178 , n5496 );
    or g2966 ( n33717 , n36419 , n10125 );
    or g2967 ( n28391 , n2581 , n10329 );
    or g2968 ( n29009 , n6503 , n2752 );
    or g2969 ( n14736 , n15604 , n36225 );
    or g2970 ( n13056 , n17304 , n34278 );
    or g2971 ( n39873 , n8010 , n22068 );
    nor g2972 ( n8378 , n14377 , n22336 );
    or g2973 ( n17604 , n19809 , n40389 );
    nor g2974 ( n3932 , n23941 , n16631 );
    or g2975 ( n33586 , n40038 , n10364 );
    or g2976 ( n28175 , n30417 , n21856 );
    and g2977 ( n23607 , n21943 , n39698 );
    or g2978 ( n29582 , n25681 , n33788 );
    and g2979 ( n11326 , n34572 , n13996 );
    not g2980 ( n14855 , n27222 );
    or g2981 ( n42024 , n24154 , n2114 );
    not g2982 ( n14457 , n30344 );
    not g2983 ( n8638 , n18953 );
    xnor g2984 ( n34889 , n258 , n14147 );
    or g2985 ( n18226 , n35614 , n36874 );
    nor g2986 ( n3700 , n4416 , n12633 );
    and g2987 ( n15918 , n34983 , n34046 );
    and g2988 ( n19911 , n39035 , n1128 );
    or g2989 ( n25399 , n19694 , n22892 );
    or g2990 ( n11341 , n18775 , n14449 );
    and g2991 ( n12352 , n26429 , n39480 );
    not g2992 ( n152 , n15533 );
    not g2993 ( n17532 , n24511 );
    xnor g2994 ( n16884 , n26579 , n7783 );
    not g2995 ( n5583 , n35493 );
    nor g2996 ( n21269 , n1338 , n19294 );
    or g2997 ( n12133 , n16292 , n21839 );
    not g2998 ( n38266 , n40674 );
    or g2999 ( n27909 , n4895 , n29787 );
    and g3000 ( n19548 , n35862 , n36885 );
    not g3001 ( n5679 , n22426 );
    or g3002 ( n42249 , n33981 , n27237 );
    and g3003 ( n18872 , n3983 , n30003 );
    and g3004 ( n24153 , n25746 , n18569 );
    not g3005 ( n22346 , n28956 );
    or g3006 ( n35693 , n27916 , n35081 );
    not g3007 ( n17880 , n928 );
    or g3008 ( n37369 , n5311 , n4570 );
    not g3009 ( n25733 , n4025 );
    and g3010 ( n21692 , n18039 , n25240 );
    or g3011 ( n18012 , n13179 , n20124 );
    or g3012 ( n27544 , n15282 , n11435 );
    and g3013 ( n41905 , n37686 , n1565 );
    not g3014 ( n17159 , n40499 );
    and g3015 ( n13065 , n33389 , n32511 );
    or g3016 ( n5668 , n27092 , n30777 );
    and g3017 ( n24895 , n32529 , n28157 );
    nor g3018 ( n25113 , n18131 , n40286 );
    or g3019 ( n32363 , n41699 , n29755 );
    xnor g3020 ( n4 , n21381 , n27071 );
    xnor g3021 ( n18225 , n260 , n13382 );
    and g3022 ( n34135 , n18280 , n32491 );
    not g3023 ( n9711 , n26005 );
    xnor g3024 ( n41781 , n20245 , n9238 );
    nor g3025 ( n776 , n16489 , n19009 );
    or g3026 ( n1476 , n38463 , n29100 );
    not g3027 ( n17293 , n42248 );
    and g3028 ( n24197 , n9624 , n20417 );
    not g3029 ( n20072 , n7574 );
    nor g3030 ( n1462 , n22534 , n5114 );
    nor g3031 ( n35426 , n3581 , n7616 );
    not g3032 ( n22950 , n1142 );
    not g3033 ( n9708 , n38097 );
    or g3034 ( n26936 , n3934 , n18313 );
    or g3035 ( n24824 , n18621 , n5183 );
    and g3036 ( n26387 , n30100 , n13743 );
    not g3037 ( n28897 , n23308 );
    not g3038 ( n2562 , n13857 );
    or g3039 ( n266 , n25656 , n4717 );
    or g3040 ( n18766 , n6440 , n14540 );
    or g3041 ( n29624 , n19221 , n27691 );
    or g3042 ( n7140 , n33640 , n34276 );
    not g3043 ( n36119 , n25853 );
    not g3044 ( n33190 , n38504 );
    and g3045 ( n701 , n21505 , n9592 );
    not g3046 ( n13913 , n25265 );
    or g3047 ( n28797 , n5170 , n36568 );
    and g3048 ( n4562 , n33620 , n10255 );
    nor g3049 ( n8302 , n27572 , n40126 );
    xnor g3050 ( n28769 , n39475 , n10439 );
    or g3051 ( n1919 , n29106 , n34267 );
    nor g3052 ( n20755 , n38430 , n21781 );
    or g3053 ( n24982 , n41601 , n8440 );
    xnor g3054 ( n3825 , n34562 , n23555 );
    not g3055 ( n24466 , n2892 );
    or g3056 ( n30507 , n19159 , n738 );
    not g3057 ( n4327 , n41950 );
    and g3058 ( n8572 , n42334 , n22958 );
    not g3059 ( n17243 , n22292 );
    and g3060 ( n12592 , n3283 , n24169 );
    not g3061 ( n37175 , n23170 );
    or g3062 ( n31752 , n16095 , n21703 );
    not g3063 ( n17429 , n2063 );
    or g3064 ( n12275 , n13974 , n5006 );
    and g3065 ( n34171 , n3484 , n14401 );
    or g3066 ( n36818 , n22579 , n14780 );
    xnor g3067 ( n27880 , n30594 , n13611 );
    not g3068 ( n38006 , n31825 );
    and g3069 ( n34110 , n12946 , n41070 );
    and g3070 ( n1994 , n22041 , n30551 );
    not g3071 ( n1015 , n665 );
    and g3072 ( n5035 , n21461 , n16179 );
    not g3073 ( n24131 , n6562 );
    and g3074 ( n5884 , n37302 , n7520 );
    and g3075 ( n40643 , n38026 , n36588 );
    not g3076 ( n2298 , n30014 );
    not g3077 ( n13444 , n35301 );
    or g3078 ( n7880 , n15147 , n11357 );
    or g3079 ( n6405 , n26520 , n42888 );
    not g3080 ( n22820 , n26902 );
    xnor g3081 ( n20061 , n3455 , n13601 );
    or g3082 ( n39510 , n36899 , n16928 );
    xnor g3083 ( n37366 , n20958 , n21531 );
    or g3084 ( n10302 , n38022 , n5620 );
    and g3085 ( n5122 , n41362 , n22874 );
    not g3086 ( n22495 , n210 );
    and g3087 ( n34222 , n26766 , n13896 );
    or g3088 ( n8170 , n1404 , n1263 );
    and g3089 ( n29583 , n4205 , n300 );
    and g3090 ( n6097 , n11748 , n39214 );
    nor g3091 ( n9327 , n22580 , n20346 );
    or g3092 ( n21449 , n14723 , n32715 );
    or g3093 ( n41557 , n9505 , n769 );
    and g3094 ( n38853 , n34968 , n25287 );
    or g3095 ( n2050 , n18072 , n14436 );
    and g3096 ( n10900 , n39950 , n31505 );
    nor g3097 ( n15701 , n35132 , n38514 );
    not g3098 ( n42152 , n26332 );
    and g3099 ( n28400 , n29223 , n14663 );
    and g3100 ( n18471 , n41060 , n3682 );
    not g3101 ( n33330 , n24531 );
    not g3102 ( n39402 , n15840 );
    and g3103 ( n8309 , n41925 , n27544 );
    and g3104 ( n22862 , n33875 , n40518 );
    xnor g3105 ( n6469 , n39455 , n34292 );
    xnor g3106 ( n4090 , n2385 , n22674 );
    or g3107 ( n7539 , n508 , n40157 );
    not g3108 ( n22428 , n19514 );
    or g3109 ( n33112 , n40966 , n22834 );
    nor g3110 ( n6555 , n26058 , n20412 );
    nor g3111 ( n42427 , n34292 , n13606 );
    nor g3112 ( n11998 , n7811 , n31767 );
    or g3113 ( n27013 , n14797 , n17104 );
    or g3114 ( n15898 , n41532 , n41877 );
    and g3115 ( n4486 , n41884 , n74 );
    or g3116 ( n6428 , n32957 , n20395 );
    or g3117 ( n10074 , n41266 , n27992 );
    or g3118 ( n21110 , n17740 , n21850 );
    xnor g3119 ( n40649 , n40 , n12756 );
    and g3120 ( n36284 , n35723 , n3391 );
    or g3121 ( n25891 , n20427 , n7558 );
    not g3122 ( n35608 , n41807 );
    xnor g3123 ( n25020 , n25619 , n30587 );
    not g3124 ( n35105 , n33170 );
    or g3125 ( n26857 , n24362 , n20473 );
    and g3126 ( n19476 , n39692 , n16685 );
    and g3127 ( n39747 , n26016 , n4992 );
    and g3128 ( n26578 , n34890 , n17103 );
    or g3129 ( n33388 , n35963 , n22985 );
    and g3130 ( n8066 , n17715 , n41202 );
    not g3131 ( n21400 , n30184 );
    or g3132 ( n21683 , n5048 , n29186 );
    and g3133 ( n4830 , n26980 , n26368 );
    or g3134 ( n5996 , n40335 , n21372 );
    not g3135 ( n3322 , n11352 );
    or g3136 ( n36044 , n16452 , n21268 );
    and g3137 ( n30142 , n25855 , n24047 );
    nor g3138 ( n14615 , n5896 , n14766 );
    nor g3139 ( n25929 , n1506 , n27677 );
    or g3140 ( n15247 , n33330 , n24563 );
    not g3141 ( n5341 , n37088 );
    and g3142 ( n39944 , n30808 , n4975 );
    or g3143 ( n37686 , n34258 , n8473 );
    or g3144 ( n16365 , n32916 , n8114 );
    or g3145 ( n15635 , n21703 , n21314 );
    and g3146 ( n39660 , n11377 , n20620 );
    or g3147 ( n9332 , n25573 , n31770 );
    xnor g3148 ( n10254 , n20872 , n28557 );
    not g3149 ( n24551 , n26120 );
    and g3150 ( n12081 , n38577 , n30000 );
    or g3151 ( n33771 , n1441 , n21496 );
    or g3152 ( n24080 , n4535 , n12690 );
    or g3153 ( n41269 , n27798 , n34243 );
    xnor g3154 ( n33168 , n28884 , n21527 );
    not g3155 ( n28489 , n10072 );
    and g3156 ( n25393 , n4571 , n17580 );
    or g3157 ( n11948 , n19503 , n8616 );
    and g3158 ( n26301 , n28747 , n18717 );
    or g3159 ( n25296 , n11952 , n31446 );
    or g3160 ( n23161 , n19786 , n10730 );
    and g3161 ( n42539 , n10942 , n20849 );
    xnor g3162 ( n13813 , n33570 , n31163 );
    and g3163 ( n34283 , n35936 , n40959 );
    or g3164 ( n33962 , n8819 , n14511 );
    not g3165 ( n14682 , n7892 );
    nor g3166 ( n29462 , n39339 , n17789 );
    or g3167 ( n29179 , n3362 , n22831 );
    or g3168 ( n20213 , n7235 , n5918 );
    and g3169 ( n25446 , n39135 , n40828 );
    and g3170 ( n11592 , n3007 , n14391 );
    or g3171 ( n18650 , n18652 , n31618 );
    xnor g3172 ( n7371 , n23025 , n32756 );
    not g3173 ( n2529 , n36953 );
    and g3174 ( n24560 , n7605 , n17391 );
    and g3175 ( n37058 , n8400 , n8672 );
    not g3176 ( n38935 , n32813 );
    and g3177 ( n6209 , n32152 , n39754 );
    nor g3178 ( n442 , n38035 , n10473 );
    or g3179 ( n28068 , n14407 , n26615 );
    not g3180 ( n23891 , n10525 );
    not g3181 ( n15131 , n32533 );
    or g3182 ( n41815 , n35089 , n33034 );
    or g3183 ( n42139 , n2223 , n12056 );
    not g3184 ( n29058 , n4517 );
    nor g3185 ( n18797 , n1336 , n4592 );
    or g3186 ( n14522 , n18424 , n5277 );
    and g3187 ( n31098 , n19250 , n2236 );
    or g3188 ( n21719 , n36117 , n7827 );
    and g3189 ( n38994 , n40797 , n16254 );
    or g3190 ( n18610 , n2789 , n5903 );
    or g3191 ( n29537 , n13178 , n15807 );
    not g3192 ( n41352 , n23455 );
    or g3193 ( n27144 , n31950 , n4600 );
    and g3194 ( n1583 , n8517 , n1018 );
    or g3195 ( n22996 , n19452 , n40019 );
    or g3196 ( n29793 , n11328 , n12672 );
    or g3197 ( n15923 , n18798 , n30799 );
    or g3198 ( n19775 , n9137 , n586 );
    or g3199 ( n30727 , n8602 , n32698 );
    or g3200 ( n6314 , n16186 , n30567 );
    and g3201 ( n5678 , n21127 , n3268 );
    xnor g3202 ( n25601 , n11436 , n26244 );
    and g3203 ( n26460 , n15543 , n3493 );
    or g3204 ( n40440 , n40253 , n11645 );
    xnor g3205 ( n32660 , n34352 , n17385 );
    and g3206 ( n30199 , n15644 , n42559 );
    and g3207 ( n18367 , n24645 , n23885 );
    and g3208 ( n21410 , n35242 , n11589 );
    nor g3209 ( n42887 , n9295 , n28469 );
    and g3210 ( n25732 , n31018 , n31880 );
    or g3211 ( n3730 , n7694 , n29060 );
    nor g3212 ( n42306 , n28563 , n19474 );
    and g3213 ( n28495 , n16425 , n14282 );
    not g3214 ( n26992 , n36298 );
    and g3215 ( n21524 , n29807 , n41251 );
    or g3216 ( n36525 , n8339 , n37553 );
    or g3217 ( n18582 , n14048 , n32139 );
    nor g3218 ( n36433 , n40929 , n26580 );
    nor g3219 ( n26001 , n1507 , n37585 );
    or g3220 ( n21355 , n34391 , n8831 );
    not g3221 ( n7949 , n9899 );
    nor g3222 ( n9509 , n1507 , n6400 );
    or g3223 ( n23766 , n26712 , n14895 );
    nor g3224 ( n11446 , n33215 , n41518 );
    and g3225 ( n5271 , n33793 , n20177 );
    and g3226 ( n12044 , n31202 , n39349 );
    xnor g3227 ( n34341 , n15467 , n18292 );
    and g3228 ( n25536 , n29587 , n42132 );
    not g3229 ( n38957 , n26201 );
    or g3230 ( n23416 , n10598 , n1138 );
    nor g3231 ( n18182 , n25688 , n20845 );
    and g3232 ( n5148 , n14311 , n15161 );
    not g3233 ( n13809 , n2242 );
    and g3234 ( n6646 , n8017 , n14429 );
    not g3235 ( n14440 , n28537 );
    and g3236 ( n17624 , n23513 , n36324 );
    nor g3237 ( n33354 , n8494 , n15012 );
    or g3238 ( n9978 , n29964 , n26823 );
    and g3239 ( n1312 , n38746 , n28838 );
    nor g3240 ( n5750 , n33838 , n30371 );
    or g3241 ( n36884 , n39904 , n37263 );
    xnor g3242 ( n27574 , n21534 , n7061 );
    xnor g3243 ( n27596 , n42118 , n7493 );
    and g3244 ( n3091 , n20433 , n7018 );
    nor g3245 ( n21242 , n36047 , n11342 );
    not g3246 ( n4355 , n18429 );
    nor g3247 ( n1020 , n16598 , n4338 );
    or g3248 ( n17993 , n32874 , n39663 );
    or g3249 ( n21131 , n13885 , n28002 );
    or g3250 ( n17945 , n15206 , n4052 );
    or g3251 ( n29734 , n6415 , n3799 );
    or g3252 ( n35863 , n40995 , n15925 );
    xnor g3253 ( n32502 , n40336 , n39486 );
    not g3254 ( n2313 , n38569 );
    and g3255 ( n6825 , n20057 , n8308 );
    not g3256 ( n25392 , n40895 );
    or g3257 ( n38873 , n39589 , n11165 );
    or g3258 ( n17085 , n8645 , n12553 );
    or g3259 ( n4720 , n41433 , n21546 );
    or g3260 ( n5412 , n29224 , n19026 );
    or g3261 ( n42837 , n12184 , n16498 );
    xnor g3262 ( n17255 , n4937 , n40080 );
    or g3263 ( n15151 , n36630 , n42251 );
    or g3264 ( n22284 , n20174 , n16314 );
    and g3265 ( n2844 , n8824 , n6304 );
    or g3266 ( n19427 , n10674 , n18712 );
    or g3267 ( n7974 , n10674 , n39294 );
    nor g3268 ( n39681 , n17744 , n2333 );
    nor g3269 ( n7595 , n3769 , n41723 );
    or g3270 ( n5702 , n42779 , n21942 );
    and g3271 ( n38169 , n26042 , n791 );
    nor g3272 ( n1497 , n1315 , n9226 );
    xnor g3273 ( n10235 , n18530 , n5790 );
    nor g3274 ( n28020 , n1847 , n12540 );
    not g3275 ( n36221 , n40373 );
    or g3276 ( n37838 , n24537 , n36408 );
    not g3277 ( n31498 , n10565 );
    or g3278 ( n13589 , n23509 , n22051 );
    nor g3279 ( n26003 , n39412 , n34743 );
    and g3280 ( n3046 , n18124 , n34220 );
    xnor g3281 ( n3004 , n14506 , n10467 );
    nor g3282 ( n5854 , n2199 , n40231 );
    or g3283 ( n15494 , n33154 , n40952 );
    nor g3284 ( n39776 , n30856 , n23909 );
    or g3285 ( n28085 , n40867 , n11210 );
    not g3286 ( n37647 , n22953 );
    not g3287 ( n8547 , n40041 );
    or g3288 ( n23903 , n20680 , n3715 );
    or g3289 ( n11182 , n14707 , n2330 );
    and g3290 ( n1115 , n322 , n33941 );
    not g3291 ( n28692 , n16673 );
    not g3292 ( n27298 , n14082 );
    nor g3293 ( n33142 , n17120 , n24299 );
    xnor g3294 ( n21982 , n21332 , n12219 );
    xnor g3295 ( n8159 , n31479 , n20987 );
    or g3296 ( n5014 , n7196 , n24162 );
    or g3297 ( n27314 , n37009 , n25002 );
    not g3298 ( n2753 , n5522 );
    not g3299 ( n18914 , n25607 );
    and g3300 ( n25115 , n35595 , n29003 );
    and g3301 ( n1158 , n6201 , n22733 );
    or g3302 ( n42397 , n31869 , n3728 );
    xnor g3303 ( n15055 , n15495 , n38717 );
    or g3304 ( n20466 , n38887 , n16394 );
    or g3305 ( n31359 , n27802 , n8555 );
    or g3306 ( n1154 , n29098 , n28262 );
    and g3307 ( n25886 , n40762 , n25074 );
    or g3308 ( n3470 , n29803 , n40593 );
    or g3309 ( n17046 , n35286 , n20716 );
    xnor g3310 ( n9449 , n25701 , n2039 );
    or g3311 ( n13166 , n1387 , n31979 );
    xnor g3312 ( n21502 , n23761 , n18173 );
    or g3313 ( n41834 , n10067 , n18861 );
    and g3314 ( n34384 , n29353 , n25255 );
    not g3315 ( n917 , n9382 );
    not g3316 ( n38938 , n40265 );
    and g3317 ( n41892 , n12596 , n39577 );
    or g3318 ( n25255 , n15675 , n14669 );
    not g3319 ( n37392 , n17834 );
    and g3320 ( n18271 , n27647 , n37782 );
    and g3321 ( n32150 , n30149 , n28497 );
    or g3322 ( n42341 , n22617 , n3538 );
    nor g3323 ( n3516 , n11268 , n13916 );
    not g3324 ( n21675 , n4208 );
    or g3325 ( n24130 , n4842 , n28078 );
    or g3326 ( n5693 , n4982 , n37633 );
    or g3327 ( n3827 , n13701 , n34984 );
    not g3328 ( n30840 , n17636 );
    not g3329 ( n10941 , n8833 );
    xnor g3330 ( n33019 , n34562 , n23698 );
    not g3331 ( n3795 , n13523 );
    or g3332 ( n11997 , n16897 , n944 );
    and g3333 ( n19224 , n7691 , n12404 );
    and g3334 ( n28959 , n8494 , n9404 );
    nor g3335 ( n30924 , n32720 , n24863 );
    xnor g3336 ( n36950 , n17561 , n37106 );
    nor g3337 ( n37134 , n33617 , n21531 );
    or g3338 ( n20910 , n23238 , n37942 );
    or g3339 ( n3283 , n18798 , n39749 );
    not g3340 ( n26309 , n241 );
    or g3341 ( n31863 , n3156 , n37058 );
    or g3342 ( n13805 , n14085 , n34470 );
    or g3343 ( n36777 , n38670 , n12198 );
    or g3344 ( n5346 , n13657 , n20750 );
    or g3345 ( n41367 , n27626 , n25545 );
    or g3346 ( n33273 , n36901 , n20145 );
    or g3347 ( n7738 , n36401 , n25343 );
    and g3348 ( n16287 , n39685 , n7470 );
    and g3349 ( n1273 , n37319 , n21945 );
    or g3350 ( n15939 , n36914 , n10179 );
    nor g3351 ( n15188 , n22040 , n36199 );
    or g3352 ( n17619 , n16736 , n18756 );
    or g3353 ( n20289 , n22447 , n19600 );
    and g3354 ( n19765 , n25870 , n21699 );
    xnor g3355 ( n25879 , n38749 , n27132 );
    or g3356 ( n33460 , n26935 , n8803 );
    and g3357 ( n17726 , n35935 , n17458 );
    not g3358 ( n33556 , n41321 );
    or g3359 ( n13382 , n10199 , n3924 );
    or g3360 ( n31174 , n39617 , n27039 );
    xnor g3361 ( n23351 , n19052 , n3330 );
    and g3362 ( n4532 , n5084 , n31650 );
    xnor g3363 ( n16528 , n37899 , n37565 );
    or g3364 ( n318 , n141 , n30243 );
    or g3365 ( n2208 , n1815 , n13437 );
    xnor g3366 ( n38774 , n12146 , n35815 );
    xnor g3367 ( n41489 , n26776 , n38879 );
    or g3368 ( n34746 , n28771 , n19288 );
    or g3369 ( n38226 , n20511 , n9405 );
    not g3370 ( n20851 , n33639 );
    not g3371 ( n1406 , n14351 );
    nor g3372 ( n16694 , n8547 , n24423 );
    not g3373 ( n41669 , n30993 );
    xnor g3374 ( n22702 , n105 , n17844 );
    and g3375 ( n3706 , n20371 , n15816 );
    or g3376 ( n1715 , n24261 , n38211 );
    or g3377 ( n14926 , n16897 , n28765 );
    or g3378 ( n38230 , n14112 , n27145 );
    xnor g3379 ( n30343 , n11633 , n35019 );
    or g3380 ( n36307 , n12663 , n37134 );
    or g3381 ( n34387 , n19471 , n39956 );
    not g3382 ( n35386 , n8202 );
    not g3383 ( n34922 , n36843 );
    nor g3384 ( n4991 , n6364 , n16162 );
    or g3385 ( n6343 , n15426 , n40665 );
    and g3386 ( n5472 , n19697 , n14818 );
    and g3387 ( n17798 , n23383 , n7967 );
    and g3388 ( n10542 , n6551 , n6556 );
    not g3389 ( n29623 , n39841 );
    or g3390 ( n17412 , n42874 , n425 );
    nor g3391 ( n28955 , n41699 , n10180 );
    nor g3392 ( n3912 , n7763 , n28809 );
    or g3393 ( n32619 , n4046 , n27127 );
    and g3394 ( n6726 , n3168 , n32049 );
    not g3395 ( n15813 , n40997 );
    or g3396 ( n11681 , n14083 , n6959 );
    xnor g3397 ( n27076 , n11436 , n8374 );
    or g3398 ( n1741 , n17877 , n26157 );
    or g3399 ( n11335 , n33013 , n14567 );
    xnor g3400 ( n3193 , n26691 , n15963 );
    and g3401 ( n39479 , n10228 , n24913 );
    and g3402 ( n23420 , n23367 , n27979 );
    and g3403 ( n34217 , n7480 , n2580 );
    nor g3404 ( n19103 , n26447 , n9739 );
    not g3405 ( n27446 , n25570 );
    and g3406 ( n30914 , n7105 , n37929 );
    or g3407 ( n34297 , n25483 , n16971 );
    or g3408 ( n37660 , n33328 , n10670 );
    nor g3409 ( n5713 , n41699 , n14317 );
    or g3410 ( n25322 , n2095 , n18065 );
    xnor g3411 ( n686 , n7489 , n17503 );
    and g3412 ( n23498 , n23836 , n38070 );
    not g3413 ( n9775 , n10614 );
    or g3414 ( n11422 , n30691 , n824 );
    or g3415 ( n26039 , n17135 , n37120 );
    or g3416 ( n23630 , n9823 , n35531 );
    and g3417 ( n25289 , n31099 , n12819 );
    or g3418 ( n37962 , n11571 , n1023 );
    or g3419 ( n34252 , n41260 , n16806 );
    nor g3420 ( n7288 , n31074 , n7014 );
    not g3421 ( n38801 , n25647 );
    or g3422 ( n35597 , n14374 , n11732 );
    and g3423 ( n3992 , n23086 , n4731 );
    nor g3424 ( n33712 , n8494 , n22480 );
    not g3425 ( n21268 , n9874 );
    or g3426 ( n16518 , n4312 , n20296 );
    or g3427 ( n6800 , n38333 , n23949 );
    and g3428 ( n3811 , n42120 , n32945 );
    or g3429 ( n11421 , n2556 , n42722 );
    not g3430 ( n33639 , n5337 );
    and g3431 ( n8619 , n8868 , n6816 );
    nor g3432 ( n4575 , n3453 , n17571 );
    xnor g3433 ( n10304 , n36539 , n31760 );
    or g3434 ( n6495 , n4842 , n21722 );
    xnor g3435 ( n39180 , n9886 , n25403 );
    and g3436 ( n10623 , n38302 , n22978 );
    and g3437 ( n40759 , n15209 , n34104 );
    or g3438 ( n40282 , n41773 , n13163 );
    and g3439 ( n14895 , n35343 , n20435 );
    or g3440 ( n23275 , n8978 , n10892 );
    and g3441 ( n27062 , n18940 , n27032 );
    and g3442 ( n30976 , n29123 , n22305 );
    not g3443 ( n22812 , n3101 );
    not g3444 ( n22837 , n31155 );
    and g3445 ( n26204 , n18903 , n29483 );
    or g3446 ( n16071 , n16926 , n19179 );
    or g3447 ( n20926 , n17073 , n40062 );
    not g3448 ( n14622 , n27506 );
    nor g3449 ( n12757 , n751 , n21563 );
    or g3450 ( n5733 , n18139 , n33775 );
    xnor g3451 ( n35599 , n36009 , n11857 );
    not g3452 ( n39903 , n18934 );
    or g3453 ( n9791 , n1577 , n8914 );
    xnor g3454 ( n1858 , n32178 , n38795 );
    and g3455 ( n30666 , n17261 , n22643 );
    xnor g3456 ( n31376 , n4501 , n42105 );
    not g3457 ( n28320 , n40833 );
    nor g3458 ( n41930 , n24356 , n11685 );
    or g3459 ( n33425 , n39946 , n39533 );
    nor g3460 ( n5525 , n726 , n20594 );
    or g3461 ( n17518 , n15914 , n32489 );
    and g3462 ( n31753 , n9305 , n6724 );
    and g3463 ( n40665 , n13561 , n2397 );
    nor g3464 ( n16881 , n25729 , n9325 );
    or g3465 ( n36260 , n3502 , n31168 );
    xnor g3466 ( n5111 , n24912 , n13875 );
    not g3467 ( n623 , n31528 );
    not g3468 ( n21090 , n3446 );
    or g3469 ( n3216 , n5896 , n27367 );
    nor g3470 ( n9553 , n26446 , n15968 );
    and g3471 ( n32971 , n28250 , n29725 );
    not g3472 ( n29429 , n10554 );
    xnor g3473 ( n29783 , n24943 , n41284 );
    or g3474 ( n14328 , n8413 , n22201 );
    or g3475 ( n41825 , n13571 , n35586 );
    or g3476 ( n19908 , n1500 , n4567 );
    not g3477 ( n15118 , n13714 );
    or g3478 ( n4878 , n6174 , n41355 );
    nor g3479 ( n41768 , n16726 , n18892 );
    or g3480 ( n2932 , n33030 , n10874 );
    and g3481 ( n40184 , n33938 , n16326 );
    xnor g3482 ( n1311 , n1113 , n8494 );
    nor g3483 ( n10217 , n4820 , n33 );
    or g3484 ( n7177 , n35847 , n5261 );
    and g3485 ( n1335 , n11609 , n38970 );
    and g3486 ( n28111 , n12516 , n33969 );
    or g3487 ( n27615 , n4335 , n7050 );
    nor g3488 ( n8761 , n42298 , n12151 );
    and g3489 ( n39844 , n35894 , n16450 );
    and g3490 ( n2153 , n23529 , n401 );
    or g3491 ( n6237 , n22201 , n1718 );
    xnor g3492 ( n39669 , n28443 , n23498 );
    or g3493 ( n12438 , n19811 , n9075 );
    or g3494 ( n5160 , n7850 , n3487 );
    or g3495 ( n31545 , n14724 , n5419 );
    nor g3496 ( n11746 , n36806 , n23779 );
    and g3497 ( n4144 , n16478 , n23371 );
    not g3498 ( n34634 , n16264 );
    or g3499 ( n14285 , n14471 , n1309 );
    nor g3500 ( n23623 , n24190 , n9883 );
    or g3501 ( n20340 , n33216 , n37100 );
    or g3502 ( n8854 , n14504 , n12739 );
    or g3503 ( n34154 , n18120 , n10020 );
    or g3504 ( n2642 , n7775 , n1735 );
    or g3505 ( n3493 , n32277 , n451 );
    nor g3506 ( n16502 , n8812 , n20192 );
    or g3507 ( n37078 , n30204 , n42657 );
    nor g3508 ( n9134 , n27801 , n20610 );
    or g3509 ( n30556 , n27153 , n17055 );
    and g3510 ( n29495 , n28864 , n36493 );
    or g3511 ( n35669 , n38149 , n34567 );
    and g3512 ( n30908 , n39748 , n25663 );
    not g3513 ( n9151 , n5915 );
    or g3514 ( n35440 , n25501 , n5978 );
    not g3515 ( n17036 , n14632 );
    or g3516 ( n10541 , n3632 , n18102 );
    and g3517 ( n18756 , n28652 , n16277 );
    and g3518 ( n30086 , n11744 , n15456 );
    or g3519 ( n30661 , n35572 , n24752 );
    or g3520 ( n20235 , n5859 , n17641 );
    nor g3521 ( n34189 , n34565 , n9207 );
    xor g3522 ( n35051 , n10747 , n37158 );
    not g3523 ( n11595 , n37306 );
    xnor g3524 ( n34973 , n4558 , n17488 );
    or g3525 ( n23278 , n35281 , n25996 );
    and g3526 ( n38524 , n41773 , n41039 );
    not g3527 ( n11368 , n875 );
    and g3528 ( n27459 , n40941 , n3594 );
    and g3529 ( n33912 , n39703 , n9153 );
    or g3530 ( n20034 , n4717 , n24299 );
    not g3531 ( n16566 , n21439 );
    and g3532 ( n24215 , n11772 , n1040 );
    or g3533 ( n5870 , n18737 , n13703 );
    or g3534 ( n34347 , n28468 , n1661 );
    or g3535 ( n28190 , n17968 , n28887 );
    not g3536 ( n7448 , n19026 );
    xnor g3537 ( n36898 , n15480 , n19979 );
    xnor g3538 ( n35575 , n11855 , n18394 );
    or g3539 ( n8684 , n36558 , n26495 );
    or g3540 ( n34717 , n16780 , n8945 );
    or g3541 ( n18655 , n4335 , n5059 );
    or g3542 ( n34597 , n35267 , n7447 );
    not g3543 ( n4905 , n7014 );
    or g3544 ( n33381 , n8584 , n15895 );
    or g3545 ( n38139 , n34720 , n17827 );
    nor g3546 ( n25444 , n10565 , n37610 );
    nor g3547 ( n4332 , n30568 , n1587 );
    nor g3548 ( n30357 , n545 , n6029 );
    xnor g3549 ( n19037 , n16215 , n41762 );
    not g3550 ( n33632 , n5186 );
    and g3551 ( n30728 , n15064 , n38424 );
    or g3552 ( n16449 , n42405 , n16499 );
    or g3553 ( n42785 , n1651 , n14851 );
    or g3554 ( n38432 , n26933 , n39131 );
    nor g3555 ( n27277 , n42556 , n26275 );
    or g3556 ( n1604 , n22004 , n29884 );
    xnor g3557 ( n29436 , n9020 , n36179 );
    or g3558 ( n11748 , n7560 , n2982 );
    or g3559 ( n31160 , n35719 , n39869 );
    not g3560 ( n33951 , n7824 );
    not g3561 ( n3735 , n10072 );
    and g3562 ( n37558 , n17266 , n11873 );
    nor g3563 ( n903 , n35590 , n25449 );
    not g3564 ( n39365 , n21178 );
    and g3565 ( n5586 , n380 , n42350 );
    not g3566 ( n4040 , n16127 );
    not g3567 ( n37561 , n4159 );
    or g3568 ( n13270 , n34779 , n31234 );
    or g3569 ( n2930 , n5232 , n39580 );
    or g3570 ( n27409 , n32800 , n29772 );
    xnor g3571 ( n19305 , n18840 , n22050 );
    nor g3572 ( n10204 , n1197 , n19969 );
    nor g3573 ( n27788 , n16965 , n29444 );
    nor g3574 ( n35610 , n4140 , n13051 );
    xnor g3575 ( n41027 , n17315 , n37151 );
    nor g3576 ( n21611 , n40982 , n36516 );
    xnor g3577 ( n5417 , n31290 , n3267 );
    or g3578 ( n17479 , n14407 , n40017 );
    xnor g3579 ( n1826 , n105 , n31399 );
    or g3580 ( n17400 , n18618 , n33600 );
    xnor g3581 ( n31896 , n21973 , n42867 );
    or g3582 ( n9081 , n14707 , n6550 );
    and g3583 ( n7994 , n10309 , n39668 );
    or g3584 ( n11240 , n41086 , n5035 );
    and g3585 ( n21847 , n19024 , n35842 );
    nor g3586 ( n42227 , n28075 , n39519 );
    not g3587 ( n15842 , n16699 );
    nor g3588 ( n35492 , n28917 , n5812 );
    or g3589 ( n13326 , n42327 , n8402 );
    not g3590 ( n28335 , n2298 );
    xnor g3591 ( n4848 , n16532 , n31771 );
    and g3592 ( n17407 , n1125 , n30256 );
    or g3593 ( n8533 , n29280 , n11986 );
    or g3594 ( n39938 , n5192 , n7199 );
    or g3595 ( n66 , n11513 , n24408 );
    or g3596 ( n26531 , n34565 , n8494 );
    xnor g3597 ( n13022 , n35015 , n4938 );
    or g3598 ( n3268 , n11327 , n15257 );
    xnor g3599 ( n6787 , n41145 , n16973 );
    xnor g3600 ( n19141 , n25057 , n35434 );
    and g3601 ( n35518 , n13292 , n19956 );
    and g3602 ( n21123 , n13595 , n17184 );
    nor g3603 ( n22850 , n5413 , n39974 );
    nor g3604 ( n23954 , n23657 , n5368 );
    or g3605 ( n21169 , n11196 , n2802 );
    not g3606 ( n24062 , n9754 );
    not g3607 ( n12939 , n35305 );
    nor g3608 ( n3590 , n11345 , n39336 );
    nor g3609 ( n35730 , n14815 , n17115 );
    or g3610 ( n14428 , n16996 , n20431 );
    or g3611 ( n11623 , n29031 , n38669 );
    or g3612 ( n12444 , n42446 , n8813 );
    or g3613 ( n11315 , n4657 , n25704 );
    or g3614 ( n24936 , n34132 , n28461 );
    xnor g3615 ( n28323 , n32042 , n10161 );
    nor g3616 ( n183 , n36307 , n31224 );
    not g3617 ( n37777 , n9657 );
    nor g3618 ( n15351 , n26069 , n7655 );
    not g3619 ( n9796 , n21480 );
    xnor g3620 ( n38162 , n12919 , n30289 );
    or g3621 ( n29654 , n7111 , n37346 );
    and g3622 ( n25840 , n7588 , n12274 );
    or g3623 ( n622 , n30585 , n11310 );
    or g3624 ( n12737 , n12872 , n42419 );
    or g3625 ( n40744 , n29058 , n21243 );
    or g3626 ( n17213 , n21359 , n462 );
    or g3627 ( n34934 , n20163 , n34421 );
    or g3628 ( n19062 , n37131 , n38113 );
    and g3629 ( n26185 , n42607 , n23433 );
    nor g3630 ( n38360 , n41773 , n15701 );
    or g3631 ( n12701 , n34202 , n38713 );
    not g3632 ( n12392 , n2486 );
    nor g3633 ( n10086 , n37356 , n5231 );
    and g3634 ( n31727 , n41872 , n5604 );
    and g3635 ( n41089 , n11875 , n32281 );
    not g3636 ( n8953 , n30911 );
    or g3637 ( n10959 , n34793 , n20652 );
    nor g3638 ( n37217 , n562 , n10638 );
    nor g3639 ( n10082 , n5531 , n39058 );
    and g3640 ( n33445 , n17324 , n138 );
    xnor g3641 ( n12960 , n15467 , n34738 );
    and g3642 ( n7979 , n39877 , n8807 );
    nor g3643 ( n11735 , n27206 , n40359 );
    or g3644 ( n37870 , n4028 , n13830 );
    or g3645 ( n28001 , n23598 , n828 );
    nor g3646 ( n30963 , n31837 , n19347 );
    and g3647 ( n17244 , n8300 , n38936 );
    xnor g3648 ( n25605 , n5144 , n8703 );
    or g3649 ( n25511 , n41547 , n3551 );
    xnor g3650 ( n3124 , n33253 , n29021 );
    and g3651 ( n3931 , n41970 , n32769 );
    and g3652 ( n19097 , n14542 , n12747 );
    or g3653 ( n23594 , n6295 , n21860 );
    and g3654 ( n31584 , n42679 , n15824 );
    or g3655 ( n21635 , n18866 , n27904 );
    not g3656 ( n21966 , n34062 );
    not g3657 ( n6813 , n26275 );
    or g3658 ( n22801 , n30489 , n2095 );
    or g3659 ( n146 , n37015 , n37250 );
    and g3660 ( n15731 , n20313 , n2347 );
    or g3661 ( n34191 , n41679 , n31156 );
    and g3662 ( n6971 , n20970 , n28147 );
    xnor g3663 ( n11130 , n1768 , n41351 );
    or g3664 ( n28004 , n42610 , n39954 );
    not g3665 ( n7984 , n5478 );
    xnor g3666 ( n4272 , n14399 , n37310 );
    or g3667 ( n29805 , n11766 , n33780 );
    not g3668 ( n42479 , n33803 );
    and g3669 ( n32137 , n25972 , n33533 );
    or g3670 ( n38396 , n19425 , n39911 );
    or g3671 ( n40148 , n33464 , n25888 );
    or g3672 ( n1833 , n16564 , n41088 );
    nor g3673 ( n3021 , n24373 , n7914 );
    not g3674 ( n31570 , n24088 );
    or g3675 ( n39156 , n25557 , n16687 );
    not g3676 ( n29534 , n1485 );
    xnor g3677 ( n31938 , n11436 , n21091 );
    or g3678 ( n10847 , n7215 , n34677 );
    and g3679 ( n6282 , n9272 , n9070 );
    xnor g3680 ( n37487 , n28231 , n10304 );
    xnor g3681 ( n26271 , n3146 , n31759 );
    nor g3682 ( n16678 , n39935 , n15140 );
    xnor g3683 ( n35499 , n2503 , n72 );
    not g3684 ( n12414 , n20113 );
    and g3685 ( n29564 , n23251 , n38850 );
    or g3686 ( n21996 , n2367 , n15371 );
    xnor g3687 ( n31024 , n36973 , n2867 );
    or g3688 ( n28977 , n7756 , n28889 );
    or g3689 ( n23914 , n23378 , n29077 );
    not g3690 ( n18638 , n6887 );
    not g3691 ( n31617 , n39446 );
    or g3692 ( n38596 , n30908 , n30358 );
    not g3693 ( n15388 , n32887 );
    not g3694 ( n31999 , n42425 );
    nor g3695 ( n10599 , n30145 , n13882 );
    or g3696 ( n29471 , n1900 , n17416 );
    xnor g3697 ( n17673 , n14594 , n21076 );
    not g3698 ( n24218 , n11409 );
    xnor g3699 ( n2888 , n1224 , n7714 );
    xnor g3700 ( n26362 , n21133 , n21833 );
    or g3701 ( n7529 , n4470 , n40144 );
    xnor g3702 ( n18365 , n31989 , n26491 );
    and g3703 ( n18782 , n14037 , n8570 );
    and g3704 ( n15897 , n2360 , n42741 );
    or g3705 ( n14914 , n2972 , n7354 );
    or g3706 ( n20931 , n39954 , n17190 );
    or g3707 ( n36746 , n22730 , n21526 );
    and g3708 ( n24400 , n16919 , n3965 );
    or g3709 ( n6996 , n11152 , n21172 );
    or g3710 ( n33489 , n25964 , n3917 );
    not g3711 ( n41337 , n26366 );
    or g3712 ( n38528 , n37771 , n24598 );
    or g3713 ( n25082 , n30822 , n14873 );
    and g3714 ( n25499 , n6314 , n39925 );
    xnor g3715 ( n26440 , n11426 , n11620 );
    or g3716 ( n18845 , n31918 , n39761 );
    nor g3717 ( n16456 , n1507 , n11218 );
    not g3718 ( n34987 , n23469 );
    and g3719 ( n28625 , n29940 , n27528 );
    and g3720 ( n33196 , n13853 , n42608 );
    nor g3721 ( n28996 , n16811 , n18238 );
    or g3722 ( n24269 , n23637 , n16313 );
    nor g3723 ( n11005 , n26794 , n4704 );
    xnor g3724 ( n32899 , n29740 , n23453 );
    or g3725 ( n8639 , n9955 , n31627 );
    or g3726 ( n1901 , n1656 , n28684 );
    nor g3727 ( n41156 , n12230 , n20353 );
    or g3728 ( n10036 , n29800 , n25303 );
    or g3729 ( n19721 , n42792 , n30305 );
    nor g3730 ( n40952 , n39412 , n4323 );
    nor g3731 ( n26889 , n28593 , n3709 );
    or g3732 ( n38546 , n17224 , n5261 );
    and g3733 ( n7873 , n13431 , n9689 );
    or g3734 ( n9520 , n10511 , n32340 );
    and g3735 ( n14240 , n16551 , n5838 );
    or g3736 ( n25901 , n3417 , n20503 );
    not g3737 ( n23164 , n14274 );
    not g3738 ( n11766 , n37815 );
    or g3739 ( n27095 , n30068 , n15038 );
    or g3740 ( n39856 , n3392 , n41526 );
    or g3741 ( n925 , n18495 , n29986 );
    or g3742 ( n13086 , n24530 , n19540 );
    nor g3743 ( n21342 , n22207 , n26798 );
    or g3744 ( n21040 , n41307 , n37674 );
    or g3745 ( n37936 , n4926 , n25480 );
    nor g3746 ( n34749 , n25826 , n11620 );
    or g3747 ( n17364 , n28024 , n3190 );
    or g3748 ( n23020 , n41225 , n38626 );
    and g3749 ( n32830 , n31445 , n42336 );
    and g3750 ( n19935 , n1384 , n35052 );
    or g3751 ( n24648 , n3526 , n18459 );
    or g3752 ( n25257 , n39165 , n28080 );
    or g3753 ( n42496 , n35337 , n25900 );
    not g3754 ( n33740 , n19776 );
    not g3755 ( n27958 , n33091 );
    nor g3756 ( n9764 , n12894 , n26271 );
    or g3757 ( n27497 , n35156 , n32582 );
    or g3758 ( n36605 , n644 , n7237 );
    or g3759 ( n31173 , n2586 , n22718 );
    and g3760 ( n38622 , n9029 , n23391 );
    or g3761 ( n6219 , n5197 , n17856 );
    nor g3762 ( n3130 , n24442 , n41858 );
    or g3763 ( n22854 , n19307 , n38562 );
    nor g3764 ( n4219 , n12921 , n11990 );
    not g3765 ( n34030 , n4208 );
    or g3766 ( n1304 , n4271 , n38845 );
    or g3767 ( n11124 , n39521 , n11960 );
    or g3768 ( n26429 , n23082 , n36802 );
    not g3769 ( n14434 , n29389 );
    and g3770 ( n940 , n29503 , n10995 );
    and g3771 ( n24582 , n38634 , n26282 );
    or g3772 ( n34798 , n7414 , n9399 );
    xnor g3773 ( n15258 , n22899 , n25127 );
    xnor g3774 ( n25639 , n6760 , n33728 );
    and g3775 ( n11362 , n16173 , n13079 );
    not g3776 ( n1075 , n12734 );
    or g3777 ( n35783 , n22161 , n32885 );
    xnor g3778 ( n35961 , n5759 , n2180 );
    and g3779 ( n40714 , n12611 , n3495 );
    or g3780 ( n40260 , n22570 , n39517 );
    xnor g3781 ( n23034 , n18625 , n36765 );
    or g3782 ( n13372 , n17610 , n30517 );
    nor g3783 ( n35365 , n20167 , n28953 );
    not g3784 ( n10375 , n21354 );
    xnor g3785 ( n29160 , n9775 , n2316 );
    not g3786 ( n29412 , n24724 );
    not g3787 ( n3431 , n18350 );
    and g3788 ( n38530 , n38686 , n32763 );
    or g3789 ( n38522 , n11899 , n26285 );
    nor g3790 ( n19117 , n14471 , n10075 );
    and g3791 ( n27691 , n30636 , n19758 );
    or g3792 ( n1347 , n3738 , n4461 );
    nor g3793 ( n25073 , n34292 , n24581 );
    or g3794 ( n29602 , n7230 , n20644 );
    or g3795 ( n13434 , n26895 , n2773 );
    or g3796 ( n30277 , n94 , n38783 );
    nor g3797 ( n38347 , n25727 , n13021 );
    not g3798 ( n33628 , n3560 );
    not g3799 ( n21925 , n15784 );
    not g3800 ( n38395 , n10661 );
    or g3801 ( n35650 , n31061 , n3408 );
    xnor g3802 ( n5332 , n22263 , n17506 );
    or g3803 ( n25396 , n27098 , n9282 );
    or g3804 ( n3169 , n9508 , n15085 );
    not g3805 ( n26591 , n1977 );
    xnor g3806 ( n24553 , n3713 , n35032 );
    not g3807 ( n11410 , n33626 );
    or g3808 ( n18531 , n29857 , n27580 );
    or g3809 ( n1163 , n15987 , n433 );
    xnor g3810 ( n19703 , n37153 , n17135 );
    nor g3811 ( n39983 , n20707 , n12744 );
    or g3812 ( n19717 , n14557 , n13687 );
    xnor g3813 ( n12881 , n36667 , n16578 );
    xnor g3814 ( n19197 , n28156 , n30944 );
    or g3815 ( n39629 , n8993 , n27603 );
    and g3816 ( n41456 , n1005 , n13184 );
    xnor g3817 ( n28631 , n35322 , n8980 );
    and g3818 ( n22618 , n25185 , n2641 );
    or g3819 ( n22768 , n16256 , n21942 );
    and g3820 ( n21473 , n9295 , n28469 );
    or g3821 ( n27003 , n39213 , n33440 );
    xnor g3822 ( n23839 , n11436 , n20018 );
    not g3823 ( n3442 , n12069 );
    or g3824 ( n10668 , n33951 , n32681 );
    nor g3825 ( n33333 , n36158 , n11576 );
    or g3826 ( n27853 , n24924 , n41954 );
    not g3827 ( n27053 , n30809 );
    xnor g3828 ( n6177 , n22546 , n25654 );
    not g3829 ( n17152 , n35060 );
    or g3830 ( n26107 , n33167 , n28021 );
    or g3831 ( n30535 , n21703 , n6037 );
    or g3832 ( n32655 , n32070 , n19312 );
    and g3833 ( n18166 , n40203 , n20303 );
    xnor g3834 ( n19624 , n14242 , n34473 );
    or g3835 ( n41482 , n18877 , n38996 );
    or g3836 ( n41535 , n35915 , n8503 );
    or g3837 ( n38605 , n42405 , n6665 );
    or g3838 ( n32678 , n31542 , n37809 );
    not g3839 ( n31677 , n24846 );
    not g3840 ( n34008 , n21379 );
    and g3841 ( n39528 , n23839 , n6200 );
    or g3842 ( n20607 , n29219 , n18406 );
    and g3843 ( n16683 , n39060 , n37875 );
    not g3844 ( n16511 , n22669 );
    not g3845 ( n17252 , n22533 );
    and g3846 ( n40144 , n11910 , n5621 );
    or g3847 ( n30148 , n18866 , n6053 );
    or g3848 ( n25177 , n35258 , n21023 );
    not g3849 ( n15293 , n5388 );
    or g3850 ( n34453 , n32092 , n6615 );
    not g3851 ( n6178 , n18122 );
    or g3852 ( n37826 , n10677 , n24732 );
    or g3853 ( n32115 , n38879 , n659 );
    not g3854 ( n13489 , n29958 );
    or g3855 ( n9144 , n1358 , n19805 );
    or g3856 ( n7183 , n39977 , n14579 );
    xnor g3857 ( n21077 , n34731 , n42321 );
    xnor g3858 ( n42480 , n15972 , n16497 );
    not g3859 ( n35307 , n21515 );
    and g3860 ( n20378 , n26955 , n20155 );
    xnor g3861 ( n17333 , n32470 , n4160 );
    or g3862 ( n25330 , n16505 , n37642 );
    and g3863 ( n20089 , n37130 , n12254 );
    or g3864 ( n12091 , n15375 , n17012 );
    or g3865 ( n20320 , n31443 , n30616 );
    not g3866 ( n29330 , n25768 );
    nor g3867 ( n35085 , n35927 , n4148 );
    or g3868 ( n37416 , n38173 , n13587 );
    or g3869 ( n29671 , n14286 , n3543 );
    or g3870 ( n18489 , n18326 , n29915 );
    nor g3871 ( n3848 , n14707 , n16784 );
    xnor g3872 ( n24572 , n35525 , n32440 );
    or g3873 ( n40188 , n4745 , n22808 );
    or g3874 ( n28354 , n9253 , n28861 );
    or g3875 ( n37668 , n27793 , n17900 );
    or g3876 ( n20944 , n3867 , n38196 );
    not g3877 ( n14468 , n9182 );
    or g3878 ( n38368 , n14707 , n23744 );
    and g3879 ( n19405 , n18678 , n5945 );
    not g3880 ( n24243 , n24372 );
    or g3881 ( n6245 , n7742 , n4669 );
    nor g3882 ( n41169 , n21769 , n4614 );
    nor g3883 ( n24217 , n19547 , n9009 );
    and g3884 ( n9790 , n20211 , n9069 );
    nor g3885 ( n37852 , n40228 , n10244 );
    not g3886 ( n16160 , n26565 );
    nor g3887 ( n25236 , n27281 , n12042 );
    not g3888 ( n13974 , n27837 );
    xnor g3889 ( n34968 , n14932 , n12415 );
    and g3890 ( n19727 , n20871 , n17741 );
    not g3891 ( n38174 , n38043 );
    or g3892 ( n6725 , n41961 , n41732 );
    xnor g3893 ( n7357 , n28851 , n40603 );
    nor g3894 ( n26790 , n8122 , n36384 );
    xnor g3895 ( n37130 , n41013 , n4101 );
    or g3896 ( n34563 , n14647 , n1893 );
    or g3897 ( n17803 , n26179 , n14489 );
    and g3898 ( n12415 , n28012 , n7402 );
    not g3899 ( n28745 , n570 );
    and g3900 ( n11048 , n35240 , n3527 );
    or g3901 ( n41142 , n19929 , n19660 );
    and g3902 ( n22294 , n21459 , n15752 );
    and g3903 ( n8324 , n1179 , n41796 );
    or g3904 ( n28988 , n16673 , n23378 );
    xnor g3905 ( n4519 , n40337 , n9263 );
    not g3906 ( n4872 , n36132 );
    or g3907 ( n20011 , n35483 , n13862 );
    and g3908 ( n21216 , n36212 , n16015 );
    and g3909 ( n38763 , n30858 , n34451 );
    and g3910 ( n21221 , n22613 , n37345 );
    nor g3911 ( n26760 , n30558 , n1411 );
    or g3912 ( n42 , n29346 , n41107 );
    nor g3913 ( n30835 , n16598 , n36862 );
    not g3914 ( n15564 , n22574 );
    xnor g3915 ( n34975 , n41218 , n38348 );
    xnor g3916 ( n31355 , n17673 , n9685 );
    and g3917 ( n17045 , n35084 , n35926 );
    and g3918 ( n14680 , n6064 , n38210 );
    or g3919 ( n15469 , n14595 , n15040 );
    xnor g3920 ( n29604 , n37876 , n19684 );
    or g3921 ( n30174 , n20941 , n42544 );
    xnor g3922 ( n33595 , n20487 , n12075 );
    or g3923 ( n4153 , n17109 , n42135 );
    or g3924 ( n15736 , n12943 , n12598 );
    or g3925 ( n26137 , n1246 , n16764 );
    not g3926 ( n21700 , n1787 );
    or g3927 ( n42178 , n24022 , n2647 );
    xnor g3928 ( n35342 , n12086 , n17615 );
    or g3929 ( n42661 , n29609 , n23374 );
    and g3930 ( n19036 , n31148 , n42576 );
    or g3931 ( n39069 , n33708 , n32165 );
    and g3932 ( n42824 , n40864 , n27479 );
    not g3933 ( n23736 , n40297 );
    nor g3934 ( n38435 , n16057 , n6441 );
    or g3935 ( n2383 , n41601 , n8032 );
    and g3936 ( n40916 , n32431 , n34152 );
    and g3937 ( n28675 , n13740 , n38478 );
    nor g3938 ( n26360 , n33570 , n42406 );
    or g3939 ( n39085 , n29336 , n38423 );
    xnor g3940 ( n3052 , n25673 , n34300 );
    and g3941 ( n42518 , n28332 , n7392 );
    nor g3942 ( n32718 , n5144 , n27043 );
    or g3943 ( n1976 , n27924 , n816 );
    and g3944 ( n12375 , n38502 , n23142 );
    not g3945 ( n5411 , n2413 );
    and g3946 ( n180 , n3990 , n33861 );
    and g3947 ( n41533 , n25296 , n19032 );
    or g3948 ( n31745 , n30919 , n40138 );
    and g3949 ( n42223 , n34795 , n17760 );
    or g3950 ( n26067 , n35534 , n12725 );
    or g3951 ( n3669 , n38273 , n32410 );
    or g3952 ( n31977 , n25715 , n26050 );
    nor g3953 ( n22098 , n34292 , n32185 );
    or g3954 ( n30804 , n15010 , n22199 );
    xnor g3955 ( n40895 , n36998 , n20939 );
    or g3956 ( n19889 , n30349 , n3715 );
    not g3957 ( n18466 , n19607 );
    or g3958 ( n37473 , n31370 , n35216 );
    not g3959 ( n4074 , n34726 );
    or g3960 ( n36385 , n9151 , n38690 );
    and g3961 ( n24739 , n13838 , n10781 );
    not g3962 ( n27895 , n7561 );
    and g3963 ( n2658 , n9190 , n35929 );
    not g3964 ( n991 , n14224 );
    nor g3965 ( n9349 , n9035 , n7493 );
    and g3966 ( n35418 , n4790 , n14185 );
    or g3967 ( n15395 , n27989 , n33243 );
    or g3968 ( n37650 , n31261 , n25674 );
    not g3969 ( n1404 , n29892 );
    or g3970 ( n24859 , n38996 , n13003 );
    and g3971 ( n6930 , n8642 , n26441 );
    and g3972 ( n32668 , n3450 , n26464 );
    or g3973 ( n7919 , n23655 , n40178 );
    or g3974 ( n17791 , n28143 , n17165 );
    not g3975 ( n16967 , n4886 );
    or g3976 ( n6697 , n30091 , n22320 );
    or g3977 ( n19246 , n33903 , n41207 );
    not g3978 ( n23923 , n8009 );
    or g3979 ( n38803 , n34703 , n19848 );
    or g3980 ( n14148 , n344 , n16558 );
    nor g3981 ( n38896 , n42572 , n25460 );
    and g3982 ( n25968 , n7736 , n31017 );
    or g3983 ( n21497 , n19774 , n42625 );
    xnor g3984 ( n25572 , n35471 , n36368 );
    or g3985 ( n42892 , n40148 , n15599 );
    or g3986 ( n9379 , n11617 , n33101 );
    or g3987 ( n11565 , n31963 , n1289 );
    and g3988 ( n28885 , n9611 , n39860 );
    or g3989 ( n1099 , n14481 , n35384 );
    xnor g3990 ( n25414 , n28443 , n27306 );
    or g3991 ( n16934 , n1484 , n29309 );
    or g3992 ( n23985 , n25907 , n3267 );
    nor g3993 ( n15092 , n15070 , n24400 );
    or g3994 ( n11064 , n13282 , n30028 );
    or g3995 ( n38627 , n4022 , n17987 );
    not g3996 ( n24250 , n3970 );
    and g3997 ( n29615 , n41749 , n18559 );
    and g3998 ( n3525 , n29446 , n33503 );
    or g3999 ( n13829 , n28013 , n6976 );
    not g4000 ( n15054 , n33435 );
    and g4001 ( n29957 , n42436 , n17143 );
    or g4002 ( n14437 , n40271 , n19346 );
    not g4003 ( n14181 , n36384 );
    xnor g4004 ( n40581 , n32427 , n36610 );
    or g4005 ( n14977 , n37255 , n5987 );
    and g4006 ( n32060 , n25688 , n20845 );
    or g4007 ( n36025 , n39929 , n13468 );
    or g4008 ( n28990 , n9417 , n7019 );
    or g4009 ( n16120 , n4470 , n474 );
    nor g4010 ( n32195 , n16660 , n12198 );
    or g4011 ( n21672 , n39118 , n9632 );
    nor g4012 ( n36258 , n6539 , n2978 );
    or g4013 ( n22697 , n26904 , n36407 );
    or g4014 ( n9758 , n8626 , n673 );
    xnor g4015 ( n7796 , n29796 , n775 );
    or g4016 ( n27541 , n39746 , n10491 );
    or g4017 ( n13214 , n18775 , n13061 );
    xnor g4018 ( n2082 , n21003 , n13763 );
    and g4019 ( n15044 , n3070 , n30661 );
    or g4020 ( n26593 , n4948 , n19340 );
    and g4021 ( n6216 , n39418 , n24039 );
    not g4022 ( n13887 , n42049 );
    nor g4023 ( n35076 , n2688 , n22789 );
    or g4024 ( n15491 , n2505 , n21584 );
    or g4025 ( n42095 , n1233 , n30435 );
    and g4026 ( n16006 , n24302 , n8858 );
    or g4027 ( n34765 , n24547 , n9 );
    xnor g4028 ( n4657 , n14330 , n28493 );
    and g4029 ( n6588 , n41921 , n36270 );
    xnor g4030 ( n36677 , n37235 , n30173 );
    or g4031 ( n9229 , n16530 , n14790 );
    not g4032 ( n19020 , n38486 );
    xnor g4033 ( n9004 , n27658 , n799 );
    and g4034 ( n41939 , n40640 , n23222 );
    or g4035 ( n6155 , n36807 , n28262 );
    not g4036 ( n12233 , n8266 );
    and g4037 ( n30799 , n29070 , n9227 );
    xnor g4038 ( n19039 , n36998 , n21103 );
    not g4039 ( n21457 , n27895 );
    not g4040 ( n6011 , n30877 );
    nor g4041 ( n37099 , n33026 , n20369 );
    not g4042 ( n13455 , n31432 );
    not g4043 ( n9654 , n32273 );
    and g4044 ( n35739 , n26246 , n24741 );
    and g4045 ( n7749 , n19200 , n16413 );
    xnor g4046 ( n34892 , n119 , n27194 );
    not g4047 ( n32600 , n4591 );
    or g4048 ( n26136 , n22247 , n35798 );
    or g4049 ( n42768 , n27311 , n15278 );
    and g4050 ( n29596 , n41380 , n13924 );
    or g4051 ( n37398 , n7683 , n35834 );
    and g4052 ( n39570 , n5920 , n37318 );
    and g4053 ( n6098 , n4430 , n35424 );
    or g4054 ( n6953 , n11050 , n41350 );
    not g4055 ( n21402 , n42283 );
    or g4056 ( n12111 , n6423 , n11362 );
    not g4057 ( n17827 , n23595 );
    not g4058 ( n22387 , n36137 );
    not g4059 ( n42343 , n41755 );
    xnor g4060 ( n17530 , n9050 , n36406 );
    xnor g4061 ( n18934 , n14969 , n10976 );
    or g4062 ( n29626 , n5605 , n42875 );
    nor g4063 ( n10672 , n14471 , n13446 );
    and g4064 ( n7483 , n6010 , n7631 );
    and g4065 ( n33316 , n15490 , n34895 );
    and g4066 ( n10928 , n19541 , n11396 );
    and g4067 ( n14598 , n20602 , n28379 );
    and g4068 ( n3560 , n11944 , n25358 );
    or g4069 ( n31182 , n17255 , n19209 );
    nor g4070 ( n17972 , n14338 , n33666 );
    xnor g4071 ( n2462 , n36998 , n39958 );
    nor g4072 ( n15276 , n26446 , n17149 );
    not g4073 ( n23823 , n20737 );
    or g4074 ( n1851 , n31374 , n31146 );
    not g4075 ( n7986 , n15196 );
    and g4076 ( n38153 , n21610 , n2985 );
    or g4077 ( n26291 , n24898 , n11068 );
    and g4078 ( n35818 , n28671 , n39868 );
    or g4079 ( n35991 , n11231 , n28894 );
    and g4080 ( n37954 , n8478 , n38498 );
    not g4081 ( n31791 , n13106 );
    and g4082 ( n1327 , n39498 , n42656 );
    and g4083 ( n41509 , n14446 , n14849 );
    and g4084 ( n6365 , n15648 , n2871 );
    and g4085 ( n19668 , n29206 , n2741 );
    not g4086 ( n28258 , n33240 );
    and g4087 ( n4740 , n41013 , n5731 );
    nor g4088 ( n22013 , n23868 , n20748 );
    and g4089 ( n12672 , n23712 , n7080 );
    or g4090 ( n18076 , n2066 , n31469 );
    and g4091 ( n37505 , n14284 , n34680 );
    and g4092 ( n23959 , n212 , n40873 );
    or g4093 ( n15146 , n3357 , n37906 );
    and g4094 ( n21031 , n33201 , n13982 );
    and g4095 ( n11818 , n26649 , n5659 );
    or g4096 ( n38460 , n31517 , n41632 );
    or g4097 ( n28146 , n31649 , n42165 );
    and g4098 ( n3417 , n15853 , n17202 );
    or g4099 ( n16686 , n16545 , n14622 );
    not g4100 ( n19618 , n25013 );
    nor g4101 ( n31750 , n35301 , n21906 );
    or g4102 ( n37714 , n30369 , n19117 );
    nor g4103 ( n20259 , n31791 , n23313 );
    nor g4104 ( n2151 , n33973 , n232 );
    and g4105 ( n38773 , n2566 , n39777 );
    xnor g4106 ( n247 , n28612 , n2153 );
    not g4107 ( n5696 , n35932 );
    not g4108 ( n5634 , n36718 );
    nor g4109 ( n8568 , n5367 , n36971 );
    or g4110 ( n13499 , n425 , n31301 );
    and g4111 ( n9127 , n33988 , n434 );
    not g4112 ( n11785 , n12634 );
    or g4113 ( n2879 , n37980 , n32424 );
    or g4114 ( n15189 , n41386 , n35866 );
    not g4115 ( n34440 , n1862 );
    or g4116 ( n35496 , n13616 , n2063 );
    and g4117 ( n33040 , n28664 , n31204 );
    or g4118 ( n34573 , n5092 , n7952 );
    nor g4119 ( n28472 , n6011 , n42177 );
    xnor g4120 ( n26355 , n36998 , n34228 );
    or g4121 ( n24685 , n2720 , n13825 );
    nor g4122 ( n17361 , n1153 , n38994 );
    or g4123 ( n29723 , n24103 , n6367 );
    xnor g4124 ( n28126 , n39178 , n5426 );
    or g4125 ( n954 , n17478 , n14149 );
    xnor g4126 ( n1303 , n2263 , n11381 );
    not g4127 ( n20461 , n35279 );
    not g4128 ( n1255 , n8663 );
    and g4129 ( n6299 , n5732 , n20441 );
    not g4130 ( n30864 , n24000 );
    not g4131 ( n22268 , n34789 );
    or g4132 ( n35725 , n20703 , n18364 );
    not g4133 ( n7648 , n4391 );
    or g4134 ( n26779 , n10953 , n13877 );
    or g4135 ( n34220 , n27015 , n25343 );
    or g4136 ( n38625 , n11794 , n10560 );
    not g4137 ( n37694 , n13009 );
    nor g4138 ( n36283 , n17120 , n21820 );
    or g4139 ( n25825 , n18844 , n32180 );
    nor g4140 ( n11762 , n28698 , n29800 );
    and g4141 ( n34422 , n11187 , n3393 );
    nor g4142 ( n39608 , n12156 , n7013 );
    not g4143 ( n30830 , n35394 );
    or g4144 ( n3282 , n30282 , n38006 );
    not g4145 ( n19086 , n8240 );
    and g4146 ( n30881 , n20376 , n21619 );
    nor g4147 ( n17968 , n19990 , n27520 );
    and g4148 ( n21873 , n6538 , n37321 );
    nor g4149 ( n12205 , n8589 , n35076 );
    or g4150 ( n25205 , n35868 , n32130 );
    and g4151 ( n38406 , n473 , n41772 );
    or g4152 ( n3279 , n23790 , n20520 );
    nor g4153 ( n34850 , n23535 , n32038 );
    not g4154 ( n29030 , n4122 );
    xnor g4155 ( n2242 , n323 , n38879 );
    not g4156 ( n4919 , n15224 );
    and g4157 ( n36549 , n12312 , n20044 );
    and g4158 ( n22818 , n14929 , n19887 );
    and g4159 ( n5658 , n12932 , n37080 );
    not g4160 ( n15178 , n32147 );
    and g4161 ( n28425 , n21326 , n14257 );
    or g4162 ( n17290 , n8126 , n17017 );
    nor g4163 ( n38808 , n4743 , n8920 );
    or g4164 ( n1423 , n3856 , n17706 );
    or g4165 ( n15181 , n5408 , n15931 );
    not g4166 ( n30014 , n39145 );
    xnor g4167 ( n15523 , n38260 , n16213 );
    or g4168 ( n8956 , n28745 , n10907 );
    not g4169 ( n11524 , n22339 );
    and g4170 ( n7773 , n28730 , n24524 );
    or g4171 ( n42784 , n28689 , n6690 );
    or g4172 ( n34991 , n10499 , n26147 );
    nor g4173 ( n6987 , n5905 , n26261 );
    xnor g4174 ( n25324 , n20451 , n34565 );
    or g4175 ( n9230 , n19848 , n23406 );
    and g4176 ( n31967 , n33767 , n12715 );
    and g4177 ( n2116 , n39486 , n40336 );
    and g4178 ( n8808 , n523 , n30946 );
    or g4179 ( n29863 , n16067 , n32180 );
    and g4180 ( n9839 , n2508 , n29203 );
    and g4181 ( n18974 , n31808 , n29605 );
    and g4182 ( n3775 , n18297 , n18416 );
    not g4183 ( n39364 , n5016 );
    and g4184 ( n41813 , n29392 , n42236 );
    nor g4185 ( n13112 , n5896 , n24326 );
    nor g4186 ( n26592 , n42553 , n15009 );
    not g4187 ( n14974 , n32958 );
    and g4188 ( n3291 , n19028 , n15453 );
    nor g4189 ( n6976 , n19221 , n23756 );
    and g4190 ( n31669 , n15070 , n32293 );
    and g4191 ( n32566 , n15961 , n11992 );
    nor g4192 ( n16488 , n2199 , n28200 );
    or g4193 ( n2536 , n37112 , n292 );
    or g4194 ( n12644 , n881 , n33217 );
    or g4195 ( n37226 , n40389 , n31747 );
    not g4196 ( n21973 , n24610 );
    or g4197 ( n15704 , n24307 , n11603 );
    not g4198 ( n13720 , n1287 );
    and g4199 ( n35631 , n13047 , n26333 );
    not g4200 ( n9508 , n24747 );
    not g4201 ( n21515 , n34021 );
    or g4202 ( n7233 , n7708 , n40787 );
    and g4203 ( n2815 , n29424 , n39305 );
    and g4204 ( n42855 , n7246 , n18125 );
    and g4205 ( n24635 , n30179 , n42402 );
    or g4206 ( n19500 , n15070 , n32151 );
    and g4207 ( n38904 , n10164 , n39657 );
    xnor g4208 ( n23656 , n27713 , n42889 );
    and g4209 ( n7048 , n11687 , n1328 );
    nor g4210 ( n36299 , n2199 , n216 );
    not g4211 ( n23934 , n2302 );
    nor g4212 ( n10400 , n16598 , n5218 );
    not g4213 ( n18348 , n31757 );
    xnor g4214 ( n33278 , n39640 , n40495 );
    or g4215 ( n28671 , n9824 , n27868 );
    and g4216 ( n7549 , n34768 , n35794 );
    not g4217 ( n38555 , n36953 );
    xnor g4218 ( n20770 , n5144 , n15550 );
    nor g4219 ( n6493 , n6179 , n17190 );
    or g4220 ( n3105 , n20710 , n31156 );
    or g4221 ( n26487 , n3812 , n22288 );
    and g4222 ( n36995 , n3061 , n3624 );
    nor g4223 ( n9185 , n14813 , n27080 );
    not g4224 ( n15621 , n14865 );
    or g4225 ( n30987 , n16339 , n40371 );
    and g4226 ( n11378 , n28071 , n29376 );
    or g4227 ( n28679 , n21357 , n18473 );
    or g4228 ( n19646 , n16617 , n12139 );
    nor g4229 ( n27377 , n25539 , n33242 );
    or g4230 ( n41198 , n35294 , n28604 );
    nor g4231 ( n28532 , n11663 , n15258 );
    and g4232 ( n29712 , n27608 , n9498 );
    or g4233 ( n32076 , n13918 , n35410 );
    or g4234 ( n7163 , n26928 , n26640 );
    or g4235 ( n39234 , n14350 , n42569 );
    not g4236 ( n8615 , n32620 );
    or g4237 ( n30175 , n10266 , n9428 );
    or g4238 ( n4423 , n20729 , n2184 );
    or g4239 ( n3734 , n25349 , n37900 );
    not g4240 ( n13784 , n39176 );
    or g4241 ( n40594 , n9377 , n12992 );
    or g4242 ( n37456 , n33365 , n9670 );
    not g4243 ( n42557 , n22680 );
    and g4244 ( n338 , n12513 , n8598 );
    nor g4245 ( n2812 , n2370 , n20185 );
    not g4246 ( n21987 , n11414 );
    nor g4247 ( n26939 , n5001 , n10879 );
    and g4248 ( n13375 , n2421 , n3175 );
    nor g4249 ( n40685 , n4154 , n15307 );
    and g4250 ( n564 , n28192 , n40963 );
    xnor g4251 ( n9985 , n16693 , n25702 );
    xnor g4252 ( n35487 , n18954 , n14450 );
    not g4253 ( n6809 , n15441 );
    xnor g4254 ( n8257 , n31989 , n29693 );
    or g4255 ( n26188 , n27124 , n31156 );
    and g4256 ( n26795 , n11227 , n17820 );
    or g4257 ( n1983 , n20089 , n20050 );
    and g4258 ( n18731 , n40328 , n35435 );
    or g4259 ( n35920 , n550 , n7453 );
    and g4260 ( n31773 , n4647 , n4005 );
    or g4261 ( n9922 , n4660 , n13926 );
    or g4262 ( n8161 , n22417 , n9779 );
    and g4263 ( n36076 , n6334 , n10372 );
    or g4264 ( n26863 , n11066 , n17249 );
    and g4265 ( n25902 , n4386 , n28498 );
    not g4266 ( n39452 , n4122 );
    not g4267 ( n21992 , n8673 );
    or g4268 ( n15949 , n17036 , n7287 );
    or g4269 ( n22101 , n23012 , n35028 );
    not g4270 ( n16049 , n2114 );
    not g4271 ( n18584 , n4587 );
    not g4272 ( n40874 , n15605 );
    or g4273 ( n34912 , n17256 , n4850 );
    xnor g4274 ( n33678 , n32351 , n15013 );
    not g4275 ( n6423 , n29987 );
    or g4276 ( n25048 , n18009 , n35120 );
    not g4277 ( n29028 , n19257 );
    or g4278 ( n34663 , n20418 , n9216 );
    nor g4279 ( n32639 , n26178 , n10315 );
    nor g4280 ( n10066 , n28649 , n10452 );
    xnor g4281 ( n16619 , n14502 , n42857 );
    and g4282 ( n41942 , n32713 , n32373 );
    or g4283 ( n20704 , n2526 , n41977 );
    nor g4284 ( n42778 , n5302 , n11797 );
    and g4285 ( n6905 , n30855 , n8982 );
    or g4286 ( n7292 , n16910 , n15917 );
    or g4287 ( n36989 , n19149 , n36343 );
    and g4288 ( n27933 , n20679 , n27054 );
    not g4289 ( n2149 , n3151 );
    xnor g4290 ( n33990 , n24978 , n9209 );
    and g4291 ( n34248 , n29553 , n18241 );
    and g4292 ( n2732 , n26254 , n38513 );
    nor g4293 ( n33762 , n8515 , n33415 );
    xnor g4294 ( n39701 , n30022 , n9724 );
    or g4295 ( n6214 , n12051 , n7985 );
    not g4296 ( n3536 , n10725 );
    or g4297 ( n11933 , n6978 , n24037 );
    not g4298 ( n42544 , n32273 );
    not g4299 ( n40476 , n19667 );
    or g4300 ( n36927 , n31372 , n1493 );
    and g4301 ( n3215 , n33341 , n23598 );
    xnor g4302 ( n33203 , n42480 , n23072 );
    or g4303 ( n11275 , n39206 , n12947 );
    xnor g4304 ( n42827 , n2183 , n38034 );
    or g4305 ( n4876 , n6764 , n3480 );
    xnor g4306 ( n9071 , n11785 , n10007 );
    or g4307 ( n33138 , n26961 , n30112 );
    not g4308 ( n26663 , n35916 );
    or g4309 ( n17419 , n7346 , n42447 );
    or g4310 ( n9267 , n3909 , n13400 );
    not g4311 ( n30496 , n32905 );
    and g4312 ( n35375 , n35502 , n32292 );
    and g4313 ( n20407 , n20043 , n7596 );
    or g4314 ( n40745 , n32263 , n4584 );
    or g4315 ( n17978 , n40710 , n9515 );
    and g4316 ( n418 , n1773 , n33756 );
    xnor g4317 ( n1059 , n39721 , n3127 );
    or g4318 ( n41763 , n20851 , n30010 );
    not g4319 ( n20067 , n38263 );
    not g4320 ( n41147 , n11264 );
    or g4321 ( n39597 , n27924 , n25446 );
    not g4322 ( n5046 , n10709 );
    or g4323 ( n28951 , n8723 , n29508 );
    or g4324 ( n8316 , n26789 , n19224 );
    or g4325 ( n31445 , n36223 , n25858 );
    and g4326 ( n11286 , n13822 , n19577 );
    or g4327 ( n14021 , n12058 , n38363 );
    and g4328 ( n26895 , n10117 , n20815 );
    not g4329 ( n11216 , n10039 );
    not g4330 ( n30271 , n16253 );
    xnor g4331 ( n31568 , n23964 , n19938 );
    nor g4332 ( n28813 , n36697 , n5044 );
    nor g4333 ( n28180 , n31084 , n7497 );
    or g4334 ( n29433 , n8790 , n10433 );
    and g4335 ( n4751 , n35363 , n42112 );
    not g4336 ( n4280 , n32273 );
    or g4337 ( n21262 , n33615 , n16281 );
    and g4338 ( n10645 , n4681 , n14229 );
    or g4339 ( n8921 , n28807 , n2084 );
    or g4340 ( n33443 , n9322 , n16144 );
    or g4341 ( n386 , n16736 , n7732 );
    not g4342 ( n34752 , n34082 );
    not g4343 ( n25858 , n42268 );
    xnor g4344 ( n28628 , n542 , n25966 );
    or g4345 ( n42555 , n24734 , n27327 );
    or g4346 ( n37349 , n37564 , n36619 );
    xnor g4347 ( n28548 , n29740 , n17057 );
    not g4348 ( n38168 , n30463 );
    xnor g4349 ( n3607 , n25552 , n32811 );
    and g4350 ( n32368 , n16245 , n23706 );
    or g4351 ( n25550 , n12915 , n10926 );
    or g4352 ( n18725 , n38517 , n39539 );
    or g4353 ( n13027 , n16276 , n36520 );
    nor g4354 ( n20535 , n15070 , n3874 );
    not g4355 ( n30089 , n11740 );
    not g4356 ( n3728 , n20131 );
    and g4357 ( n33055 , n3069 , n34242 );
    or g4358 ( n10911 , n31538 , n3077 );
    not g4359 ( n4370 , n21254 );
    and g4360 ( n2238 , n24647 , n42458 );
    or g4361 ( n8987 , n4798 , n21865 );
    or g4362 ( n36769 , n33901 , n13124 );
    xnor g4363 ( n33089 , n35381 , n8822 );
    nor g4364 ( n24160 , n38356 , n27112 );
    and g4365 ( n7041 , n18288 , n11811 );
    and g4366 ( n23733 , n6917 , n41559 );
    or g4367 ( n3777 , n33963 , n4625 );
    and g4368 ( n14563 , n22854 , n318 );
    and g4369 ( n15974 , n22796 , n41690 );
    not g4370 ( n41961 , n21029 );
    xnor g4371 ( n8423 , n33179 , n42902 );
    nor g4372 ( n13278 , n8018 , n41994 );
    and g4373 ( n9896 , n37113 , n40708 );
    nor g4374 ( n19074 , n9275 , n18501 );
    or g4375 ( n17480 , n17654 , n18659 );
    nor g4376 ( n5995 , n4977 , n32862 );
    or g4377 ( n12916 , n15342 , n38061 );
    not g4378 ( n12389 , n24273 );
    or g4379 ( n17141 , n15094 , n26740 );
    or g4380 ( n3354 , n35430 , n41904 );
    and g4381 ( n24693 , n13060 , n28929 );
    and g4382 ( n7040 , n14943 , n40935 );
    and g4383 ( n34605 , n23358 , n22165 );
    nor g4384 ( n35178 , n7511 , n15893 );
    or g4385 ( n38970 , n18930 , n4239 );
    and g4386 ( n19707 , n22507 , n37291 );
    and g4387 ( n33866 , n17813 , n4683 );
    xnor g4388 ( n2378 , n41718 , n7019 );
    xnor g4389 ( n23846 , n23322 , n3648 );
    and g4390 ( n18898 , n18878 , n19223 );
    xnor g4391 ( n32015 , n105 , n939 );
    or g4392 ( n9337 , n22288 , n25784 );
    not g4393 ( n34861 , n18211 );
    and g4394 ( n868 , n22838 , n20908 );
    xnor g4395 ( n32138 , n15591 , n610 );
    not g4396 ( n37695 , n16904 );
    xnor g4397 ( n17055 , n1765 , n5555 );
    or g4398 ( n39678 , n34961 , n41822 );
    or g4399 ( n11499 , n31772 , n12220 );
    not g4400 ( n1451 , n24191 );
    xnor g4401 ( n23336 , n26579 , n14745 );
    xnor g4402 ( n30870 , n7489 , n28750 );
    nor g4403 ( n42543 , n36218 , n8534 );
    or g4404 ( n28279 , n25948 , n30434 );
    not g4405 ( n37146 , n10072 );
    or g4406 ( n35612 , n2516 , n20383 );
    not g4407 ( n26617 , n30405 );
    and g4408 ( n28561 , n30457 , n23719 );
    not g4409 ( n35721 , n8410 );
    nor g4410 ( n19730 , n13444 , n31036 );
    xnor g4411 ( n35676 , n31607 , n32971 );
    or g4412 ( n25921 , n26698 , n38800 );
    xnor g4413 ( n42422 , n15119 , n7234 );
    nor g4414 ( n27522 , n1011 , n17031 );
    nor g4415 ( n25000 , n7444 , n14078 );
    xnor g4416 ( n16828 , n23304 , n7708 );
    or g4417 ( n37923 , n41040 , n7209 );
    and g4418 ( n33522 , n16516 , n38768 );
    or g4419 ( n7328 , n32311 , n33385 );
    and g4420 ( n24740 , n39711 , n2552 );
    or g4421 ( n20006 , n42491 , n18346 );
    or g4422 ( n13538 , n34952 , n35385 );
    not g4423 ( n40006 , n20714 );
    and g4424 ( n11711 , n13267 , n18801 );
    not g4425 ( n37269 , n5456 );
    or g4426 ( n39832 , n7391 , n38166 );
    not g4427 ( n36687 , n32596 );
    and g4428 ( n37856 , n24155 , n25695 );
    or g4429 ( n25804 , n23348 , n2502 );
    or g4430 ( n22163 , n20499 , n19847 );
    or g4431 ( n800 , n1815 , n8655 );
    and g4432 ( n13903 , n33200 , n20844 );
    or g4433 ( n37865 , n11295 , n22814 );
    nor g4434 ( n40718 , n22783 , n16302 );
    or g4435 ( n30783 , n14851 , n4593 );
    nor g4436 ( n22871 , n16907 , n4 );
    xnor g4437 ( n29675 , n14658 , n24563 );
    and g4438 ( n5459 , n5217 , n16301 );
    or g4439 ( n36838 , n32352 , n38184 );
    xnor g4440 ( n17995 , n34562 , n9802 );
    or g4441 ( n16637 , n2853 , n34560 );
    xnor g4442 ( n42421 , n3934 , n12482 );
    nor g4443 ( n20778 , n16774 , n34113 );
    or g4444 ( n6079 , n4277 , n28887 );
    and g4445 ( n36947 , n14638 , n8161 );
    not g4446 ( n13357 , n33909 );
    or g4447 ( n22337 , n8927 , n38283 );
    or g4448 ( n25375 , n19766 , n16017 );
    or g4449 ( n30370 , n13760 , n4116 );
    and g4450 ( n40304 , n11107 , n2656 );
    or g4451 ( n34741 , n41305 , n22797 );
    and g4452 ( n35317 , n32379 , n4082 );
    and g4453 ( n7715 , n32309 , n10921 );
    and g4454 ( n4995 , n8842 , n40980 );
    or g4455 ( n32732 , n35633 , n26104 );
    or g4456 ( n7195 , n3554 , n6358 );
    or g4457 ( n35765 , n32451 , n9015 );
    xnor g4458 ( n9644 , n2886 , n37370 );
    or g4459 ( n36959 , n22325 , n22944 );
    xnor g4460 ( n2541 , n22296 , n10727 );
    not g4461 ( n35963 , n40674 );
    or g4462 ( n23487 , n7843 , n23123 );
    or g4463 ( n19187 , n13553 , n32316 );
    or g4464 ( n25251 , n13486 , n16029 );
    nor g4465 ( n42387 , n3769 , n24468 );
    not g4466 ( n39828 , n36792 );
    not g4467 ( n37156 , n39887 );
    not g4468 ( n6984 , n29560 );
    xnor g4469 ( n13154 , n39962 , n24776 );
    and g4470 ( n2472 , n27030 , n39678 );
    or g4471 ( n16018 , n27490 , n29209 );
    not g4472 ( n38431 , n16075 );
    not g4473 ( n25136 , n14589 );
    or g4474 ( n29364 , n14232 , n4660 );
    nor g4475 ( n32471 , n16780 , n13340 );
    and g4476 ( n2686 , n42312 , n30142 );
    or g4477 ( n37866 , n38825 , n27806 );
    nor g4478 ( n17380 , n27398 , n40951 );
    and g4479 ( n4799 , n6948 , n7672 );
    and g4480 ( n25803 , n38277 , n41087 );
    or g4481 ( n25635 , n37031 , n5599 );
    and g4482 ( n4772 , n16546 , n26441 );
    or g4483 ( n33370 , n37977 , n30125 );
    or g4484 ( n23672 , n33544 , n5585 );
    and g4485 ( n6426 , n21826 , n17043 );
    and g4486 ( n3164 , n32043 , n25698 );
    xnor g4487 ( n28414 , n4712 , n26265 );
    or g4488 ( n33756 , n9766 , n33321 );
    or g4489 ( n37178 , n16897 , n9550 );
    or g4490 ( n11965 , n890 , n7753 );
    and g4491 ( n4884 , n21832 , n5886 );
    or g4492 ( n42713 , n30190 , n15186 );
    not g4493 ( n32657 , n38197 );
    and g4494 ( n10166 , n35293 , n3592 );
    xnor g4495 ( n39604 , n18840 , n32988 );
    not g4496 ( n16074 , n32236 );
    xnor g4497 ( n22756 , n27110 , n17120 );
    not g4498 ( n7561 , n13095 );
    not g4499 ( n3262 , n23733 );
    nor g4500 ( n15728 , n1450 , n25916 );
    or g4501 ( n23167 , n33883 , n34866 );
    or g4502 ( n35828 , n18937 , n20683 );
    xnor g4503 ( n15420 , n24943 , n41485 );
    and g4504 ( n17083 , n2709 , n6045 );
    nor g4505 ( n28005 , n34429 , n4598 );
    not g4506 ( n23624 , n37762 );
    or g4507 ( n20441 , n13317 , n31547 );
    or g4508 ( n31084 , n35864 , n26305 );
    and g4509 ( n27676 , n5807 , n7450 );
    or g4510 ( n3381 , n6503 , n15346 );
    or g4511 ( n24977 , n31323 , n10926 );
    nor g4512 ( n513 , n27519 , n23891 );
    nor g4513 ( n1050 , n33981 , n12698 );
    or g4514 ( n7081 , n26607 , n17496 );
    and g4515 ( n1663 , n3739 , n14369 );
    or g4516 ( n22408 , n40798 , n4477 );
    or g4517 ( n5867 , n19958 , n19070 );
    not g4518 ( n11047 , n27010 );
    or g4519 ( n12567 , n19065 , n15954 );
    xnor g4520 ( n27778 , n18678 , n32691 );
    nor g4521 ( n29525 , n2199 , n12546 );
    and g4522 ( n39908 , n7259 , n21901 );
    and g4523 ( n24383 , n19554 , n3600 );
    xnor g4524 ( n42281 , n22263 , n7442 );
    and g4525 ( n24647 , n14124 , n18469 );
    nor g4526 ( n40104 , n10922 , n42849 );
    and g4527 ( n10068 , n42176 , n20262 );
    or g4528 ( n7302 , n34594 , n27489 );
    not g4529 ( n14609 , n21092 );
    and g4530 ( n37179 , n19856 , n38606 );
    or g4531 ( n36183 , n20532 , n13820 );
    nor g4532 ( n19830 , n33981 , n35180 );
    and g4533 ( n23337 , n38877 , n1697 );
    not g4534 ( n5102 , n24830 );
    or g4535 ( n17451 , n23972 , n23272 );
    or g4536 ( n29698 , n25275 , n24583 );
    or g4537 ( n1481 , n34939 , n14745 );
    not g4538 ( n18449 , n38717 );
    and g4539 ( n21777 , n40309 , n10420 );
    or g4540 ( n39777 , n18058 , n17679 );
    or g4541 ( n40976 , n25102 , n33252 );
    and g4542 ( n5843 , n34205 , n21374 );
    xnor g4543 ( n255 , n30752 , n19284 );
    xnor g4544 ( n758 , n38629 , n11004 );
    nor g4545 ( n4913 , n35135 , n18187 );
    and g4546 ( n9975 , n19699 , n21744 );
    not g4547 ( n11026 , n17301 );
    not g4548 ( n20156 , n9210 );
    nor g4549 ( n24639 , n27909 , n34012 );
    and g4550 ( n11637 , n18989 , n4439 );
    nor g4551 ( n17817 , n12264 , n24582 );
    not g4552 ( n21303 , n27223 );
    xnor g4553 ( n31274 , n29129 , n17045 );
    xnor g4554 ( n26329 , n7197 , n30381 );
    nor g4555 ( n24835 , n36047 , n8733 );
    or g4556 ( n15570 , n42798 , n38697 );
    nor g4557 ( n39783 , n34245 , n25162 );
    or g4558 ( n14486 , n15565 , n40571 );
    or g4559 ( n25056 , n2511 , n17903 );
    xnor g4560 ( n42452 , n42572 , n13926 );
    not g4561 ( n30061 , n12892 );
    not g4562 ( n28205 , n29719 );
    nor g4563 ( n14548 , n3817 , n24251 );
    not g4564 ( n2673 , n29835 );
    not g4565 ( n29717 , n5259 );
    xnor g4566 ( n27049 , n31297 , n11502 );
    and g4567 ( n29542 , n33306 , n32300 );
    nor g4568 ( n29628 , n34778 , n17830 );
    or g4569 ( n28016 , n4855 , n19526 );
    not g4570 ( n39025 , n37357 );
    not g4571 ( n177 , n27570 );
    nor g4572 ( n884 , n5367 , n40480 );
    not g4573 ( n42388 , n37253 );
    or g4574 ( n19489 , n31472 , n19556 );
    and g4575 ( n38590 , n29592 , n33769 );
    xnor g4576 ( n10969 , n7980 , n41088 );
    not g4577 ( n42707 , n4012 );
    or g4578 ( n16875 , n31769 , n2190 );
    or g4579 ( n9583 , n1956 , n35443 );
    not g4580 ( n39676 , n39611 );
    xnor g4581 ( n34497 , n1443 , n11848 );
    or g4582 ( n11418 , n36002 , n33667 );
    or g4583 ( n41166 , n3372 , n21211 );
    and g4584 ( n39974 , n37795 , n25783 );
    and g4585 ( n7889 , n18850 , n830 );
    and g4586 ( n24712 , n24128 , n6642 );
    or g4587 ( n808 , n36184 , n935 );
    or g4588 ( n16747 , n22748 , n487 );
    or g4589 ( n6234 , n30143 , n11326 );
    or g4590 ( n5468 , n17545 , n26922 );
    or g4591 ( n35247 , n32410 , n31812 );
    nor g4592 ( n17896 , n34559 , n42288 );
    nor g4593 ( n37342 , n14471 , n31420 );
    not g4594 ( n2728 , n36695 );
    or g4595 ( n4202 , n34773 , n22206 );
    not g4596 ( n39803 , n28479 );
    and g4597 ( n2484 , n25641 , n15471 );
    xnor g4598 ( n10840 , n24546 , n10718 );
    nor g4599 ( n20198 , n32701 , n10632 );
    or g4600 ( n10031 , n15802 , n36726 );
    or g4601 ( n10820 , n13014 , n41079 );
    or g4602 ( n2289 , n4660 , n26841 );
    or g4603 ( n33169 , n39828 , n29241 );
    nor g4604 ( n23003 , n37006 , n40835 );
    or g4605 ( n16304 , n12456 , n42240 );
    xnor g4606 ( n9989 , n42560 , n28050 );
    or g4607 ( n4889 , n4089 , n20718 );
    and g4608 ( n41152 , n35900 , n15786 );
    xnor g4609 ( n10585 , n11595 , n29547 );
    xnor g4610 ( n14331 , n35938 , n23522 );
    or g4611 ( n40343 , n15505 , n2809 );
    or g4612 ( n1787 , n26460 , n23581 );
    and g4613 ( n24022 , n42709 , n27005 );
    not g4614 ( n22953 , n12465 );
    xnor g4615 ( n20234 , n23606 , n19546 );
    or g4616 ( n26701 , n31562 , n3964 );
    nor g4617 ( n7379 , n14349 , n32450 );
    xnor g4618 ( n25822 , n2632 , n23717 );
    and g4619 ( n9612 , n4664 , n30068 );
    and g4620 ( n28491 , n30568 , n1587 );
    or g4621 ( n11736 , n24621 , n39201 );
    not g4622 ( n31550 , n7822 );
    or g4623 ( n28286 , n2819 , n36203 );
    nor g4624 ( n1947 , n12754 , n13083 );
    or g4625 ( n26653 , n37271 , n6247 );
    or g4626 ( n20990 , n40612 , n28481 );
    or g4627 ( n42485 , n30754 , n31012 );
    or g4628 ( n5263 , n7037 , n26312 );
    not g4629 ( n19532 , n10537 );
    or g4630 ( n22394 , n15377 , n19279 );
    or g4631 ( n5239 , n41356 , n15144 );
    or g4632 ( n25644 , n16709 , n3128 );
    xnor g4633 ( n9242 , n36998 , n1139 );
    xnor g4634 ( n7858 , n6625 , n748 );
    nor g4635 ( n21290 , n7105 , n37929 );
    nor g4636 ( n20589 , n34816 , n9912 );
    or g4637 ( n10524 , n20141 , n40226 );
    not g4638 ( n19514 , n36762 );
    or g4639 ( n18554 , n5718 , n22182 );
    or g4640 ( n7480 , n3105 , n38892 );
    nor g4641 ( n6810 , n1826 , n36149 );
    or g4642 ( n31876 , n32217 , n4747 );
    or g4643 ( n24472 , n9699 , n6207 );
    and g4644 ( n7009 , n22962 , n20214 );
    not g4645 ( n27039 , n38918 );
    or g4646 ( n30528 , n38851 , n15740 );
    nor g4647 ( n12890 , n275 , n7877 );
    and g4648 ( n30713 , n11889 , n1860 );
    or g4649 ( n28865 , n5419 , n18060 );
    or g4650 ( n5920 , n35013 , n25382 );
    and g4651 ( n25546 , n29656 , n40392 );
    and g4652 ( n2807 , n24275 , n17765 );
    nor g4653 ( n27207 , n15884 , n10347 );
    or g4654 ( n11518 , n16850 , n40110 );
    or g4655 ( n13638 , n8857 , n41539 );
    or g4656 ( n7294 , n21721 , n2767 );
    and g4657 ( n35191 , n28637 , n14212 );
    or g4658 ( n6580 , n42308 , n40787 );
    or g4659 ( n38404 , n23374 , n39999 );
    nor g4660 ( n32169 , n8119 , n6061 );
    and g4661 ( n10161 , n3896 , n16098 );
    or g4662 ( n14785 , n24482 , n1763 );
    not g4663 ( n41112 , n41026 );
    or g4664 ( n26980 , n34292 , n41561 );
    or g4665 ( n9770 , n19183 , n23946 );
    xnor g4666 ( n3604 , n18558 , n8893 );
    or g4667 ( n11589 , n2297 , n38817 );
    or g4668 ( n9902 , n29490 , n27611 );
    nor g4669 ( n37107 , n35607 , n8414 );
    or g4670 ( n39333 , n40323 , n34980 );
    or g4671 ( n16250 , n34411 , n27119 );
    and g4672 ( n19269 , n22377 , n31526 );
    nor g4673 ( n38057 , n17147 , n20023 );
    or g4674 ( n31666 , n35714 , n21268 );
    nor g4675 ( n34081 , n13230 , n21305 );
    not g4676 ( n34994 , n16397 );
    or g4677 ( n26138 , n25762 , n14501 );
    not g4678 ( n28402 , n41578 );
    nor g4679 ( n26319 , n31931 , n8520 );
    or g4680 ( n2154 , n15446 , n22833 );
    and g4681 ( n19960 , n17450 , n29387 );
    or g4682 ( n1985 , n12227 , n2348 );
    or g4683 ( n40353 , n25540 , n13866 );
    and g4684 ( n41681 , n2169 , n31245 );
    nor g4685 ( n21822 , n18928 , n26546 );
    or g4686 ( n20389 , n21642 , n21021 );
    nor g4687 ( n20717 , n33602 , n35680 );
    or g4688 ( n40972 , n23211 , n25090 );
    not g4689 ( n31562 , n3938 );
    or g4690 ( n6757 , n38590 , n10181 );
    not g4691 ( n19431 , n20818 );
    or g4692 ( n8290 , n40916 , n31847 );
    not g4693 ( n42798 , n20322 );
    and g4694 ( n10212 , n28938 , n33505 );
    or g4695 ( n6967 , n29234 , n41981 );
    nor g4696 ( n30983 , n36823 , n26193 );
    and g4697 ( n35292 , n39630 , n9615 );
    nor g4698 ( n36176 , n6574 , n4326 );
    or g4699 ( n38315 , n4535 , n13569 );
    and g4700 ( n35572 , n42700 , n23470 );
    xnor g4701 ( n33420 , n31989 , n5216 );
    or g4702 ( n18059 , n8389 , n37156 );
    and g4703 ( n12619 , n33090 , n22101 );
    or g4704 ( n16767 , n36238 , n2143 );
    and g4705 ( n4874 , n10258 , n26528 );
    or g4706 ( n1876 , n41533 , n13297 );
    xnor g4707 ( n35095 , n41511 , n19022 );
    xor g4708 ( n34385 , n11488 , n33495 );
    not g4709 ( n3344 , n19571 );
    xnor g4710 ( n10083 , n31099 , n40504 );
    not g4711 ( n5826 , n13753 );
    nor g4712 ( n34378 , n9376 , n7708 );
    and g4713 ( n4255 , n30849 , n12185 );
    nor g4714 ( n33166 , n16747 , n23336 );
    or g4715 ( n41416 , n20468 , n1274 );
    and g4716 ( n21240 , n606 , n208 );
    and g4717 ( n21812 , n29125 , n29114 );
    and g4718 ( n19929 , n29371 , n14426 );
    and g4719 ( n8963 , n2390 , n13286 );
    and g4720 ( n39023 , n24938 , n11359 );
    or g4721 ( n27737 , n38463 , n11863 );
    or g4722 ( n8666 , n30853 , n19762 );
    not g4723 ( n12484 , n3178 );
    or g4724 ( n14753 , n35999 , n37103 );
    and g4725 ( n40784 , n21223 , n13056 );
    or g4726 ( n32468 , n8494 , n35378 );
    or g4727 ( n3358 , n5258 , n16948 );
    nor g4728 ( n1017 , n22100 , n5677 );
    nor g4729 ( n29659 , n32212 , n34390 );
    or g4730 ( n33073 , n26790 , n22797 );
    not g4731 ( n22112 , n668 );
    or g4732 ( n16135 , n11964 , n28331 );
    and g4733 ( n19864 , n24997 , n34898 );
    not g4734 ( n18649 , n4941 );
    not g4735 ( n15801 , n11561 );
    not g4736 ( n24424 , n3271 );
    not g4737 ( n8563 , n10408 );
    nor g4738 ( n23111 , n17393 , n5149 );
    not g4739 ( n99 , n29436 );
    or g4740 ( n11150 , n4462 , n28540 );
    or g4741 ( n22978 , n13108 , n36816 );
    and g4742 ( n7650 , n13796 , n26248 );
    or g4743 ( n9657 , n40599 , n41893 );
    nor g4744 ( n17785 , n11702 , n34448 );
    not g4745 ( n205 , n19412 );
    not g4746 ( n981 , n13105 );
    and g4747 ( n29008 , n12099 , n1000 );
    not g4748 ( n24411 , n1743 );
    nor g4749 ( n32666 , n16172 , n11828 );
    xnor g4750 ( n15782 , n11436 , n5532 );
    nor g4751 ( n42153 , n31542 , n22900 );
    or g4752 ( n20903 , n22035 , n28766 );
    or g4753 ( n5621 , n40215 , n34672 );
    or g4754 ( n11894 , n5472 , n10926 );
    xnor g4755 ( n5177 , n23947 , n15863 );
    not g4756 ( n41427 , n15441 );
    xnor g4757 ( n2350 , n37153 , n13752 );
    not g4758 ( n20728 , n23689 );
    and g4759 ( n24369 , n6190 , n25857 );
    or g4760 ( n29656 , n41654 , n7173 );
    and g4761 ( n15253 , n40370 , n12363 );
    not g4762 ( n22542 , n30410 );
    nor g4763 ( n15482 , n14091 , n27480 );
    or g4764 ( n36566 , n2844 , n33262 );
    not g4765 ( n1622 , n33130 );
    or g4766 ( n22662 , n40703 , n7279 );
    not g4767 ( n20138 , n19412 );
    or g4768 ( n30240 , n13701 , n27859 );
    not g4769 ( n35103 , n38355 );
    or g4770 ( n5450 , n14487 , n40423 );
    or g4771 ( n4595 , n15185 , n22188 );
    or g4772 ( n38583 , n27758 , n42384 );
    nor g4773 ( n30069 , n14214 , n25491 );
    or g4774 ( n35480 , n12168 , n18444 );
    xnor g4775 ( n42209 , n11633 , n6346 );
    and g4776 ( n41139 , n125 , n9758 );
    and g4777 ( n13598 , n42641 , n37472 );
    or g4778 ( n42607 , n6558 , n9941 );
    and g4779 ( n14345 , n6269 , n37228 );
    or g4780 ( n42711 , n31337 , n42128 );
    or g4781 ( n39998 , n32362 , n15888 );
    or g4782 ( n16459 , n24183 , n26761 );
    not g4783 ( n36811 , n18969 );
    or g4784 ( n39970 , n12456 , n13482 );
    or g4785 ( n23966 , n21151 , n7088 );
    not g4786 ( n7199 , n17269 );
    or g4787 ( n16313 , n18314 , n16190 );
    not g4788 ( n29394 , n20140 );
    or g4789 ( n40971 , n37195 , n37856 );
    or g4790 ( n9568 , n9894 , n16456 );
    or g4791 ( n26671 , n7951 , n18902 );
    xnor g4792 ( n7801 , n1219 , n17061 );
    not g4793 ( n8986 , n5521 );
    xnor g4794 ( n24239 , n12007 , n12379 );
    or g4795 ( n6305 , n26393 , n17888 );
    or g4796 ( n23592 , n4492 , n23771 );
    and g4797 ( n38659 , n23902 , n18383 );
    or g4798 ( n34800 , n1803 , n10008 );
    and g4799 ( n7609 , n32522 , n9630 );
    and g4800 ( n22123 , n9559 , n4396 );
    or g4801 ( n3069 , n41030 , n37762 );
    not g4802 ( n31055 , n23524 );
    or g4803 ( n16888 , n23790 , n33355 );
    and g4804 ( n1211 , n34614 , n3150 );
    xnor g4805 ( n17766 , n41067 , n40684 );
    xnor g4806 ( n34760 , n42042 , n29106 );
    and g4807 ( n10889 , n21766 , n34777 );
    and g4808 ( n2198 , n4061 , n31270 );
    or g4809 ( n14889 , n33721 , n25096 );
    nor g4810 ( n8680 , n5964 , n2155 );
    not g4811 ( n23139 , n7975 );
    and g4812 ( n12307 , n31246 , n28720 );
    xnor g4813 ( n33035 , n6112 , n20569 );
    and g4814 ( n14769 , n41446 , n2723 );
    and g4815 ( n26688 , n37441 , n5542 );
    or g4816 ( n12139 , n34584 , n40936 );
    or g4817 ( n11235 , n24243 , n9159 );
    and g4818 ( n15452 , n14661 , n1650 );
    or g4819 ( n382 , n27582 , n22767 );
    xnor g4820 ( n37522 , n28319 , n41750 );
    and g4821 ( n13633 , n14995 , n27710 );
    or g4822 ( n42358 , n15854 , n7809 );
    or g4823 ( n35593 , n16074 , n20861 );
    not g4824 ( n37436 , n41603 );
    not g4825 ( n6494 , n40000 );
    not g4826 ( n9336 , n15356 );
    or g4827 ( n14082 , n32473 , n16735 );
    or g4828 ( n36557 , n12369 , n42345 );
    not g4829 ( n15638 , n10289 );
    not g4830 ( n24254 , n30826 );
    not g4831 ( n5337 , n9774 );
    not g4832 ( n18698 , n27470 );
    and g4833 ( n30502 , n30424 , n14984 );
    or g4834 ( n30193 , n25204 , n12059 );
    or g4835 ( n17666 , n42515 , n20865 );
    or g4836 ( n15226 , n40015 , n34146 );
    or g4837 ( n36252 , n42453 , n14252 );
    not g4838 ( n30784 , n9621 );
    not g4839 ( n40638 , n7035 );
    and g4840 ( n3563 , n37268 , n24919 );
    and g4841 ( n7884 , n21944 , n25564 );
    xnor g4842 ( n14327 , n16895 , n3384 );
    not g4843 ( n41245 , n37408 );
    not g4844 ( n33867 , n20365 );
    or g4845 ( n12654 , n13050 , n16638 );
    and g4846 ( n22336 , n38515 , n22251 );
    or g4847 ( n28782 , n14471 , n27236 );
    and g4848 ( n37047 , n35903 , n39343 );
    and g4849 ( n35514 , n18759 , n2402 );
    or g4850 ( n21640 , n39672 , n40820 );
    nor g4851 ( n16043 , n17243 , n9165 );
    not g4852 ( n1980 , n8274 );
    not g4853 ( n23982 , n21431 );
    xnor g4854 ( n20945 , n21954 , n20106 );
    and g4855 ( n27380 , n21339 , n3766 );
    and g4856 ( n13199 , n10040 , n16621 );
    or g4857 ( n3593 , n40323 , n5011 );
    or g4858 ( n29025 , n38818 , n18700 );
    not g4859 ( n31861 , n8241 );
    and g4860 ( n8022 , n41634 , n39183 );
    xnor g4861 ( n31540 , n10011 , n13040 );
    or g4862 ( n20005 , n42337 , n7145 );
    not g4863 ( n37235 , n28404 );
    or g4864 ( n21316 , n4510 , n30616 );
    or g4865 ( n31117 , n29973 , n4255 );
    not g4866 ( n33114 , n32937 );
    and g4867 ( n16116 , n20074 , n1786 );
    and g4868 ( n18249 , n1782 , n4859 );
    xnor g4869 ( n3438 , n31107 , n10402 );
    xnor g4870 ( n32220 , n15591 , n1200 );
    not g4871 ( n8769 , n25126 );
    nor g4872 ( n2623 , n4561 , n41592 );
    or g4873 ( n12257 , n5693 , n33279 );
    nor g4874 ( n23775 , n5594 , n22790 );
    not g4875 ( n31124 , n20866 );
    or g4876 ( n17838 , n17927 , n33773 );
    xnor g4877 ( n12750 , n13984 , n24468 );
    or g4878 ( n9595 , n19123 , n7737 );
    nor g4879 ( n961 , n15070 , n23558 );
    nor g4880 ( n4539 , n3317 , n12718 );
    or g4881 ( n41613 , n8658 , n14001 );
    xnor g4882 ( n32186 , n33796 , n38276 );
    and g4883 ( n33922 , n21423 , n14337 );
    not g4884 ( n24297 , n39132 );
    or g4885 ( n9387 , n32011 , n22201 );
    xnor g4886 ( n2906 , n17198 , n8707 );
    xnor g4887 ( n27024 , n18702 , n40656 );
    xnor g4888 ( n35789 , n5367 , n32111 );
    nor g4889 ( n21075 , n6899 , n1822 );
    not g4890 ( n6236 , n1487 );
    nor g4891 ( n16096 , n2199 , n18042 );
    or g4892 ( n12445 , n2370 , n11629 );
    not g4893 ( n820 , n1578 );
    and g4894 ( n19980 , n24161 , n18619 );
    or g4895 ( n36650 , n33107 , n42414 );
    nor g4896 ( n29669 , n5896 , n34712 );
    or g4897 ( n9864 , n32355 , n32525 );
    not g4898 ( n12552 , n10305 );
    xnor g4899 ( n450 , n42064 , n40231 );
    and g4900 ( n12157 , n12240 , n9537 );
    xnor g4901 ( n7389 , n27767 , n8014 );
    nor g4902 ( n31797 , n28490 , n35804 );
    or g4903 ( n26926 , n36550 , n33330 );
    and g4904 ( n15942 , n15308 , n7923 );
    or g4905 ( n40125 , n34100 , n27664 );
    xnor g4906 ( n37875 , n28443 , n20194 );
    xnor g4907 ( n7680 , n41013 , n41909 );
    not g4908 ( n39590 , n34326 );
    or g4909 ( n5859 , n37154 , n38676 );
    not g4910 ( n1961 , n11640 );
    and g4911 ( n1229 , n11529 , n29941 );
    or g4912 ( n27982 , n19630 , n27071 );
    and g4913 ( n21016 , n8406 , n18551 );
    nor g4914 ( n7447 , n32305 , n41407 );
    not g4915 ( n17753 , n13306 );
    and g4916 ( n12037 , n18624 , n38220 );
    or g4917 ( n27118 , n6722 , n8467 );
    or g4918 ( n31311 , n26882 , n897 );
    and g4919 ( n27194 , n38329 , n24673 );
    and g4920 ( n435 , n29786 , n18030 );
    or g4921 ( n30781 , n16161 , n24563 );
    xnor g4922 ( n39579 , n3656 , n29338 );
    and g4923 ( n22875 , n5718 , n32018 );
    and g4924 ( n13985 , n29679 , n14028 );
    not g4925 ( n25742 , n21377 );
    nor g4926 ( n31066 , n24028 , n42117 );
    not g4927 ( n10504 , n8189 );
    or g4928 ( n35222 , n35286 , n12331 );
    or g4929 ( n31654 , n15340 , n42446 );
    or g4930 ( n3150 , n23158 , n10079 );
    nor g4931 ( n8503 , n9190 , n35929 );
    or g4932 ( n33305 , n15173 , n11962 );
    nor g4933 ( n20968 , n9490 , n8307 );
    or g4934 ( n24907 , n19254 , n21268 );
    or g4935 ( n13171 , n24475 , n31634 );
    and g4936 ( n1585 , n15505 , n27213 );
    or g4937 ( n21307 , n4839 , n2812 );
    xnor g4938 ( n21055 , n32779 , n13193 );
    or g4939 ( n3926 , n1735 , n25127 );
    or g4940 ( n33101 , n31227 , n20505 );
    not g4941 ( n13841 , n6730 );
    nor g4942 ( n10178 , n25153 , n30950 );
    or g4943 ( n30906 , n31265 , n23518 );
    nor g4944 ( n36247 , n23875 , n18592 );
    xnor g4945 ( n4143 , n13444 , n12341 );
    nor g4946 ( n22819 , n10460 , n375 );
    and g4947 ( n11200 , n40908 , n38087 );
    or g4948 ( n20747 , n730 , n37328 );
    or g4949 ( n5103 , n40478 , n12011 );
    nor g4950 ( n23027 , n5964 , n24322 );
    not g4951 ( n36937 , n7689 );
    not g4952 ( n3053 , n9512 );
    or g4953 ( n25012 , n1525 , n32752 );
    nor g4954 ( n12776 , n28698 , n12558 );
    and g4955 ( n10063 , n9422 , n8423 );
    not g4956 ( n34735 , n19952 );
    not g4957 ( n37149 , n26620 );
    xnor g4958 ( n29005 , n18093 , n22639 );
    xnor g4959 ( n28931 , n27343 , n3928 );
    or g4960 ( n19709 , n38879 , n19151 );
    not g4961 ( n29098 , n1879 );
    or g4962 ( n2075 , n4301 , n16538 );
    xnor g4963 ( n14739 , n16693 , n41777 );
    or g4964 ( n16685 , n2386 , n23620 );
    nor g4965 ( n19661 , n32670 , n5942 );
    or g4966 ( n27493 , n34766 , n34821 );
    xnor g4967 ( n20612 , n39944 , n37216 );
    not g4968 ( n31210 , n14659 );
    xnor g4969 ( n33426 , n9827 , n23457 );
    nor g4970 ( n29984 , n40846 , n21669 );
    not g4971 ( n12882 , n28658 );
    or g4972 ( n17825 , n16872 , n710 );
    not g4973 ( n38778 , n4096 );
    or g4974 ( n8195 , n17624 , n37633 );
    or g4975 ( n34771 , n12799 , n8792 );
    or g4976 ( n30654 , n4625 , n32237 );
    and g4977 ( n17500 , n30542 , n31862 );
    nor g4978 ( n23894 , n35471 , n25309 );
    and g4979 ( n23646 , n30944 , n28156 );
    and g4980 ( n8683 , n19137 , n21230 );
    or g4981 ( n15640 , n29717 , n36720 );
    not g4982 ( n26028 , n7920 );
    and g4983 ( n40241 , n21344 , n39261 );
    xnor g4984 ( n8279 , n25041 , n4333 );
    or g4985 ( n17329 , n12286 , n41858 );
    and g4986 ( n2386 , n10031 , n29501 );
    or g4987 ( n39265 , n39516 , n28405 );
    or g4988 ( n18175 , n15116 , n6177 );
    or g4989 ( n30161 , n14112 , n42248 );
    or g4990 ( n19464 , n36071 , n13725 );
    or g4991 ( n37166 , n14342 , n7142 );
    not g4992 ( n22715 , n10100 );
    not g4993 ( n2589 , n42027 );
    xnor g4994 ( n17912 , n23026 , n32040 );
    or g4995 ( n40960 , n11036 , n41649 );
    or g4996 ( n32426 , n29052 , n38993 );
    or g4997 ( n18549 , n33330 , n33977 );
    or g4998 ( n6224 , n34862 , n26727 );
    xnor g4999 ( n37635 , n15617 , n35473 );
    not g5000 ( n20193 , n35197 );
    or g5001 ( n26757 , n34411 , n24764 );
    nor g5002 ( n31716 , n2199 , n36073 );
    and g5003 ( n35369 , n25235 , n18529 );
    or g5004 ( n16823 , n35452 , n34217 );
    or g5005 ( n14319 , n24582 , n31918 );
    not g5006 ( n38814 , n11223 );
    not g5007 ( n36727 , n6818 );
    or g5008 ( n25759 , n23636 , n34821 );
    or g5009 ( n2719 , n41596 , n42152 );
    nor g5010 ( n42775 , n3795 , n33494 );
    xnor g5011 ( n26447 , n31290 , n1609 );
    not g5012 ( n29714 , n54 );
    or g5013 ( n19513 , n8579 , n26090 );
    or g5014 ( n14544 , n25770 , n19865 );
    or g5015 ( n23075 , n18718 , n30448 );
    not g5016 ( n935 , n27987 );
    or g5017 ( n25405 , n20705 , n26343 );
    not g5018 ( n13338 , n17234 );
    or g5019 ( n32152 , n38776 , n41514 );
    not g5020 ( n17779 , n14043 );
    or g5021 ( n7735 , n1369 , n38196 );
    and g5022 ( n30001 , n12202 , n38531 );
    or g5023 ( n26557 , n2296 , n7454 );
    or g5024 ( n17892 , n1456 , n21731 );
    not g5025 ( n28698 , n101 );
    nor g5026 ( n34547 , n42699 , n3919 );
    and g5027 ( n41088 , n7959 , n24667 );
    or g5028 ( n2200 , n34074 , n14053 );
    xnor g5029 ( n9877 , n13467 , n40578 );
    or g5030 ( n14006 , n3139 , n35187 );
    not g5031 ( n32154 , n8747 );
    or g5032 ( n33056 , n17771 , n24297 );
    not g5033 ( n17853 , n34788 );
    nor g5034 ( n28944 , n17052 , n4592 );
    and g5035 ( n30841 , n23671 , n37921 );
    or g5036 ( n31725 , n38942 , n23272 );
    nor g5037 ( n9064 , n21156 , n34035 );
    or g5038 ( n27614 , n39208 , n32694 );
    not g5039 ( n25570 , n4147 );
    and g5040 ( n26094 , n3633 , n1250 );
    and g5041 ( n8514 , n38978 , n30988 );
    or g5042 ( n24680 , n35489 , n21172 );
    not g5043 ( n678 , n8729 );
    nor g5044 ( n23039 , n16670 , n30177 );
    nor g5045 ( n20775 , n604 , n37731 );
    or g5046 ( n41575 , n4773 , n12484 );
    or g5047 ( n20371 , n41040 , n3627 );
    nor g5048 ( n2948 , n17376 , n9027 );
    xnor g5049 ( n15160 , n37939 , n33278 );
    nor g5050 ( n41588 , n38879 , n24723 );
    or g5051 ( n7550 , n33077 , n34428 );
    nor g5052 ( n15827 , n22458 , n33212 );
    and g5053 ( n33920 , n12479 , n17715 );
    or g5054 ( n7205 , n15922 , n5124 );
    nor g5055 ( n34528 , n51 , n18818 );
    or g5056 ( n35209 , n3240 , n244 );
    nor g5057 ( n22174 , n6145 , n3503 );
    or g5058 ( n21617 , n6348 , n26239 );
    or g5059 ( n41587 , n31347 , n32303 );
    or g5060 ( n39829 , n10648 , n39134 );
    not g5061 ( n22476 , n19878 );
    or g5062 ( n3327 , n32803 , n11761 );
    and g5063 ( n17317 , n24256 , n39130 );
    not g5064 ( n11485 , n7377 );
    and g5065 ( n27746 , n23650 , n9562 );
    or g5066 ( n26872 , n24477 , n22148 );
    xnor g5067 ( n29835 , n34337 , n17930 );
    or g5068 ( n15023 , n13446 , n16897 );
    xnor g5069 ( n9740 , n11855 , n12579 );
    not g5070 ( n26016 , n25193 );
    not g5071 ( n18468 , n22136 );
    or g5072 ( n27214 , n24626 , n10940 );
    or g5073 ( n14400 , n2664 , n13787 );
    or g5074 ( n20649 , n4609 , n32446 );
    not g5075 ( n23761 , n6065 );
    not g5076 ( n28031 , n21145 );
    nor g5077 ( n23114 , n22383 , n26906 );
    or g5078 ( n16048 , n2965 , n18869 );
    nor g5079 ( n26600 , n5834 , n16376 );
    and g5080 ( n9983 , n10510 , n35106 );
    or g5081 ( n553 , n41601 , n21806 );
    or g5082 ( n8224 , n11166 , n21784 );
    or g5083 ( n4526 , n5248 , n35358 );
    or g5084 ( n21794 , n33166 , n6004 );
    nor g5085 ( n5480 , n22300 , n28628 );
    and g5086 ( n36862 , n40124 , n19764 );
    nor g5087 ( n18207 , n38922 , n40527 );
    and g5088 ( n19029 , n6652 , n11045 );
    not g5089 ( n29414 , n14854 );
    or g5090 ( n21682 , n39195 , n37693 );
    xnor g5091 ( n23186 , n27142 , n36006 );
    or g5092 ( n19429 , n40256 , n38553 );
    not g5093 ( n14392 , n38626 );
    and g5094 ( n36883 , n31574 , n6689 );
    not g5095 ( n40301 , n26871 );
    and g5096 ( n17930 , n2100 , n9595 );
    or g5097 ( n14835 , n23444 , n4353 );
    and g5098 ( n2991 , n4685 , n15744 );
    xnor g5099 ( n23265 , n41024 , n21039 );
    and g5100 ( n29843 , n9852 , n28310 );
    or g5101 ( n20177 , n18235 , n40983 );
    or g5102 ( n39073 , n23292 , n575 );
    or g5103 ( n26191 , n15388 , n27231 );
    and g5104 ( n34672 , n10489 , n10808 );
    xnor g5105 ( n760 , n1622 , n11324 );
    not g5106 ( n22619 , n16076 );
    or g5107 ( n40708 , n25014 , n35745 );
    or g5108 ( n2360 , n232 , n7321 );
    and g5109 ( n33392 , n40650 , n29048 );
    or g5110 ( n6789 , n32368 , n11470 );
    and g5111 ( n10756 , n6640 , n21963 );
    and g5112 ( n9634 , n26126 , n41255 );
    xnor g5113 ( n10796 , n899 , n41825 );
    not g5114 ( n18757 , n1896 );
    or g5115 ( n13950 , n9264 , n26132 );
    xnor g5116 ( n30920 , n148 , n18037 );
    and g5117 ( n10586 , n42004 , n36711 );
    or g5118 ( n2978 , n10484 , n28030 );
    or g5119 ( n28770 , n33676 , n21367 );
    nor g5120 ( n2185 , n39573 , n13967 );
    xnor g5121 ( n12978 , n23231 , n41106 );
    xnor g5122 ( n6942 , n42118 , n14561 );
    and g5123 ( n36548 , n30219 , n28645 );
    not g5124 ( n36628 , n29475 );
    and g5125 ( n20970 , n31305 , n6341 );
    or g5126 ( n35200 , n32730 , n12150 );
    or g5127 ( n30632 , n13334 , n4402 );
    xnor g5128 ( n21153 , n34352 , n584 );
    not g5129 ( n17295 , n32365 );
    and g5130 ( n30812 , n12617 , n16886 );
    nor g5131 ( n22759 , n25348 , n17924 );
    or g5132 ( n21455 , n26432 , n27958 );
    or g5133 ( n37319 , n23876 , n25440 );
    xnor g5134 ( n16111 , n17264 , n39201 );
    xnor g5135 ( n12242 , n16874 , n6979 );
    or g5136 ( n25608 , n28955 , n17983 );
    or g5137 ( n10630 , n17120 , n1668 );
    not g5138 ( n22216 , n20081 );
    or g5139 ( n4714 , n14955 , n27110 );
    or g5140 ( n29899 , n21499 , n27201 );
    or g5141 ( n17197 , n27411 , n1289 );
    or g5142 ( n19316 , n13335 , n41569 );
    and g5143 ( n2190 , n29981 , n35593 );
    or g5144 ( n824 , n17286 , n33328 );
    or g5145 ( n12082 , n14945 , n35100 );
    nor g5146 ( n33611 , n5926 , n14607 );
    and g5147 ( n1666 , n37926 , n21005 );
    or g5148 ( n20355 , n14217 , n12482 );
    not g5149 ( n33164 , n20991 );
    nor g5150 ( n40111 , n23502 , n1694 );
    or g5151 ( n34033 , n15185 , n377 );
    or g5152 ( n15765 , n10434 , n33824 );
    or g5153 ( n3145 , n474 , n21023 );
    and g5154 ( n40071 , n4146 , n25534 );
    not g5155 ( n7577 , n9334 );
    or g5156 ( n34449 , n9544 , n38529 );
    and g5157 ( n38281 , n20607 , n19529 );
    xnor g5158 ( n42250 , n18530 , n3943 );
    xnor g5159 ( n40982 , n16473 , n14939 );
    or g5160 ( n20785 , n1110 , n13040 );
    nor g5161 ( n14417 , n25727 , n26601 );
    or g5162 ( n8557 , n14507 , n16512 );
    not g5163 ( n31580 , n15439 );
    and g5164 ( n36128 , n37140 , n7941 );
    or g5165 ( n31414 , n27192 , n22355 );
    or g5166 ( n19304 , n41833 , n4660 );
    xnor g5167 ( n22082 , n37437 , n33350 );
    or g5168 ( n26726 , n14120 , n16636 );
    and g5169 ( n11312 , n40460 , n15047 );
    and g5170 ( n33903 , n10824 , n23432 );
    not g5171 ( n31634 , n18637 );
    nor g5172 ( n41150 , n32047 , n39234 );
    xnor g5173 ( n38118 , n31928 , n40943 );
    and g5174 ( n41258 , n11124 , n14207 );
    xnor g5175 ( n19658 , n33794 , n6154 );
    or g5176 ( n34343 , n13724 , n41336 );
    or g5177 ( n14080 , n38356 , n42489 );
    nor g5178 ( n30646 , n36667 , n9541 );
    and g5179 ( n40175 , n39360 , n25740 );
    not g5180 ( n29239 , n25328 );
    and g5181 ( n42636 , n15002 , n6230 );
    or g5182 ( n30899 , n13390 , n29856 );
    or g5183 ( n41118 , n20411 , n7216 );
    and g5184 ( n28918 , n14174 , n39269 );
    not g5185 ( n34527 , n24747 );
    xnor g5186 ( n20489 , n28185 , n30283 );
    not g5187 ( n37538 , n20992 );
    and g5188 ( n40871 , n35334 , n20876 );
    not g5189 ( n30543 , n26989 );
    not g5190 ( n9325 , n22222 );
    or g5191 ( n34333 , n16897 , n9837 );
    not g5192 ( n17777 , n29647 );
    or g5193 ( n40782 , n20654 , n38196 );
    nor g5194 ( n40129 , n38168 , n10906 );
    or g5195 ( n38177 , n27145 , n15847 );
    or g5196 ( n40488 , n25350 , n2517 );
    xnor g5197 ( n162 , n2915 , n37482 );
    not g5198 ( n2721 , n29121 );
    or g5199 ( n39840 , n24812 , n11425 );
    and g5200 ( n29750 , n29265 , n21445 );
    not g5201 ( n20173 , n18787 );
    and g5202 ( n23751 , n9583 , n40657 );
    or g5203 ( n38394 , n20325 , n42419 );
    and g5204 ( n15481 , n21128 , n36836 );
    or g5205 ( n1109 , n18236 , n13199 );
    and g5206 ( n7092 , n12770 , n33251 );
    xnor g5207 ( n29472 , n34844 , n4887 );
    or g5208 ( n18136 , n2704 , n26807 );
    or g5209 ( n35047 , n20161 , n17912 );
    xnor g5210 ( n32283 , n23139 , n14547 );
    xnor g5211 ( n17610 , n16039 , n32295 );
    xnor g5212 ( n27286 , n27184 , n5364 );
    and g5213 ( n14999 , n37436 , n24188 );
    or g5214 ( n36556 , n36296 , n1418 );
    and g5215 ( n19188 , n26016 , n6217 );
    and g5216 ( n42370 , n36215 , n32065 );
    nor g5217 ( n9757 , n23824 , n6529 );
    xnor g5218 ( n1344 , n737 , n28739 );
    and g5219 ( n41284 , n35596 , n40580 );
    xnor g5220 ( n12025 , n31419 , n4909 );
    xnor g5221 ( n29814 , n5891 , n37305 );
    or g5222 ( n13308 , n26505 , n2597 );
    or g5223 ( n31082 , n20957 , n6533 );
    or g5224 ( n41746 , n32996 , n22631 );
    or g5225 ( n34409 , n34634 , n25814 );
    not g5226 ( n15602 , n23202 );
    not g5227 ( n24636 , n13511 );
    or g5228 ( n32630 , n27071 , n1970 );
    or g5229 ( n14076 , n3036 , n40011 );
    nor g5230 ( n18726 , n8453 , n2901 );
    and g5231 ( n18706 , n28437 , n37034 );
    or g5232 ( n35018 , n5585 , n35895 );
    nor g5233 ( n16340 , n10598 , n29165 );
    not g5234 ( n37605 , n2321 );
    xnor g5235 ( n6456 , n27722 , n5153 );
    not g5236 ( n28502 , n31775 );
    or g5237 ( n1801 , n27820 , n41684 );
    or g5238 ( n37141 , n12182 , n11629 );
    and g5239 ( n10638 , n37200 , n22367 );
    or g5240 ( n40921 , n39140 , n11037 );
    or g5241 ( n41313 , n405 , n24739 );
    or g5242 ( n40694 , n21721 , n40536 );
    or g5243 ( n19990 , n19486 , n1643 );
    not g5244 ( n25619 , n41534 );
    xnor g5245 ( n7625 , n18678 , n26386 );
    or g5246 ( n15788 , n23958 , n16792 );
    and g5247 ( n41062 , n35613 , n25859 );
    or g5248 ( n1321 , n5378 , n35695 );
    and g5249 ( n34632 , n16824 , n1150 );
    and g5250 ( n24926 , n40743 , n40971 );
    or g5251 ( n24036 , n9244 , n35167 );
    or g5252 ( n10842 , n3686 , n14407 );
    not g5253 ( n28325 , n39176 );
    or g5254 ( n39673 , n34796 , n2286 );
    nor g5255 ( n11021 , n16404 , n29253 );
    and g5256 ( n39947 , n18469 , n41883 );
    nor g5257 ( n38073 , n6426 , n5719 );
    and g5258 ( n34128 , n5865 , n19634 );
    xnor g5259 ( n14340 , n36524 , n15070 );
    and g5260 ( n39543 , n18159 , n13859 );
    xnor g5261 ( n33960 , n10558 , n23957 );
    or g5262 ( n9481 , n9245 , n30183 );
    and g5263 ( n28329 , n34521 , n36923 );
    or g5264 ( n6205 , n7463 , n23975 );
    xnor g5265 ( n32755 , n31541 , n38475 );
    not g5266 ( n24268 , n29481 );
    nor g5267 ( n22244 , n10985 , n22772 );
    nor g5268 ( n33469 , n18951 , n15011 );
    or g5269 ( n39019 , n33763 , n10206 );
    or g5270 ( n42377 , n30496 , n4017 );
    or g5271 ( n34794 , n6560 , n27816 );
    and g5272 ( n1300 , n37769 , n4344 );
    nor g5273 ( n20142 , n8656 , n9468 );
    not g5274 ( n30865 , n11145 );
    or g5275 ( n9773 , n32830 , n4717 );
    xnor g5276 ( n4181 , n4260 , n14007 );
    nor g5277 ( n39388 , n17193 , n32089 );
    or g5278 ( n36478 , n35963 , n15958 );
    and g5279 ( n24440 , n17094 , n11062 );
    xnor g5280 ( n41261 , n24588 , n36790 );
    nor g5281 ( n30912 , n40575 , n30724 );
    or g5282 ( n4433 , n21286 , n39702 );
    xnor g5283 ( n25320 , n10226 , n34552 );
    and g5284 ( n33448 , n2037 , n28609 );
    not g5285 ( n37153 , n38898 );
    xnor g5286 ( n16720 , n10084 , n13580 );
    or g5287 ( n11807 , n4070 , n12337 );
    or g5288 ( n14101 , n3552 , n10763 );
    or g5289 ( n32984 , n19212 , n10616 );
    xnor g5290 ( n21872 , n20673 , n28358 );
    and g5291 ( n6893 , n26026 , n16280 );
    or g5292 ( n40310 , n14568 , n12947 );
    nor g5293 ( n24594 , n12226 , n14711 );
    not g5294 ( n2257 , n22303 );
    nor g5295 ( n10359 , n455 , n17166 );
    not g5296 ( n22579 , n18493 );
    and g5297 ( n39788 , n28824 , n23283 );
    and g5298 ( n1405 , n3118 , n18229 );
    xnor g5299 ( n42342 , n36483 , n33982 );
    nor g5300 ( n33311 , n17120 , n5673 );
    or g5301 ( n11905 , n35483 , n30328 );
    not g5302 ( n6359 , n36723 );
    and g5303 ( n22985 , n15622 , n13925 );
    xnor g5304 ( n11063 , n40 , n38743 );
    nor g5305 ( n19102 , n4340 , n29488 );
    and g5306 ( n30053 , n34713 , n28077 );
    and g5307 ( n38475 , n29603 , n15300 );
    or g5308 ( n6605 , n41312 , n15342 );
    and g5309 ( n10880 , n23247 , n1571 );
    not g5310 ( n16587 , n7808 );
    or g5311 ( n42237 , n41089 , n13820 );
    or g5312 ( n42148 , n14379 , n7216 );
    or g5313 ( n32127 , n3424 , n26992 );
    or g5314 ( n17690 , n5364 , n39481 );
    or g5315 ( n6821 , n18934 , n4468 );
    not g5316 ( n29767 , n7271 );
    or g5317 ( n5296 , n12886 , n29214 );
    nor g5318 ( n16368 , n35839 , n2327 );
    nor g5319 ( n37361 , n20410 , n16980 );
    nor g5320 ( n38750 , n32570 , n786 );
    xnor g5321 ( n31275 , n30830 , n14184 );
    nor g5322 ( n3787 , n39568 , n29143 );
    not g5323 ( n27579 , n31028 );
    or g5324 ( n11386 , n3569 , n29058 );
    or g5325 ( n7509 , n24070 , n18103 );
    or g5326 ( n34913 , n3035 , n5757 );
    nor g5327 ( n32449 , n19024 , n35842 );
    or g5328 ( n8544 , n39489 , n41897 );
    or g5329 ( n16858 , n12845 , n12210 );
    xnor g5330 ( n12962 , n3769 , n23038 );
    or g5331 ( n34901 , n16736 , n27819 );
    xnor g5332 ( n37006 , n9619 , n27645 );
    or g5333 ( n12748 , n38257 , n22715 );
    or g5334 ( n25345 , n1348 , n36400 );
    not g5335 ( n33145 , n30987 );
    not g5336 ( n38696 , n37652 );
    xnor g5337 ( n7674 , n31092 , n19161 );
    or g5338 ( n24536 , n34499 , n14750 );
    and g5339 ( n33223 , n11547 , n4989 );
    or g5340 ( n11363 , n6586 , n10605 );
    and g5341 ( n8069 , n31456 , n41638 );
    and g5342 ( n40492 , n36710 , n28926 );
    or g5343 ( n34509 , n8581 , n34195 );
    not g5344 ( n24278 , n19407 );
    and g5345 ( n8567 , n3839 , n25274 );
    or g5346 ( n6741 , n3519 , n18083 );
    nor g5347 ( n10581 , n12543 , n39773 );
    or g5348 ( n30391 , n6774 , n1369 );
    nor g5349 ( n14018 , n5964 , n24300 );
    not g5350 ( n19702 , n25624 );
    not g5351 ( n29932 , n30959 );
    not g5352 ( n6842 , n26969 );
    nor g5353 ( n29153 , n36300 , n21271 );
    nor g5354 ( n13639 , n8008 , n12218 );
    and g5355 ( n26312 , n34325 , n24795 );
    not g5356 ( n24313 , n38410 );
    and g5357 ( n28775 , n41054 , n21627 );
    or g5358 ( n14136 , n28885 , n34278 );
    nor g5359 ( n30733 , n14476 , n11365 );
    or g5360 ( n28082 , n30730 , n10530 );
    xnor g5361 ( n16310 , n23944 , n15624 );
    not g5362 ( n4765 , n41559 );
    and g5363 ( n14547 , n21486 , n6487 );
    not g5364 ( n35711 , n12098 );
    or g5365 ( n19072 , n27193 , n34609 );
    and g5366 ( n26498 , n23021 , n19201 );
    or g5367 ( n33598 , n26098 , n416 );
    or g5368 ( n33344 , n33853 , n5585 );
    not g5369 ( n37899 , n32485 );
    or g5370 ( n18125 , n14061 , n7610 );
    and g5371 ( n8171 , n27324 , n26826 );
    or g5372 ( n18462 , n31707 , n22244 );
    or g5373 ( n28193 , n42496 , n21700 );
    xnor g5374 ( n2596 , n22263 , n37064 );
    or g5375 ( n13135 , n11768 , n7754 );
    or g5376 ( n1272 , n14420 , n22499 );
    and g5377 ( n34985 , n31203 , n40829 );
    not g5378 ( n13095 , n7109 );
    nor g5379 ( n24664 , n15572 , n26021 );
    not g5380 ( n28774 , n13300 );
    not g5381 ( n38486 , n4907 );
    and g5382 ( n41385 , n15548 , n37772 );
    not g5383 ( n5081 , n24491 );
    not g5384 ( n2661 , n8240 );
    not g5385 ( n7840 , n22426 );
    xnor g5386 ( n16514 , n11535 , n37550 );
    or g5387 ( n17125 , n20174 , n31878 );
    and g5388 ( n29024 , n22694 , n23110 );
    xnor g5389 ( n40751 , n17464 , n7356 );
    not g5390 ( n34678 , n9273 );
    xnor g5391 ( n14981 , n37083 , n9722 );
    or g5392 ( n16327 , n23757 , n35834 );
    and g5393 ( n15545 , n21185 , n17412 );
    or g5394 ( n1714 , n38149 , n14643 );
    nor g5395 ( n21570 , n10856 , n26441 );
    or g5396 ( n36133 , n15576 , n6066 );
    and g5397 ( n40931 , n23045 , n24763 );
    or g5398 ( n25913 , n21773 , n33182 );
    not g5399 ( n17727 , n7395 );
    or g5400 ( n34928 , n34994 , n28646 );
    or g5401 ( n7501 , n20975 , n2328 );
    nor g5402 ( n16993 , n12646 , n31406 );
    not g5403 ( n18933 , n39737 );
    or g5404 ( n20668 , n32064 , n40367 );
    and g5405 ( n33350 , n24370 , n20909 );
    or g5406 ( n859 , n7551 , n20813 );
    and g5407 ( n20663 , n17523 , n26263 );
    not g5408 ( n25370 , n13301 );
    xnor g5409 ( n11454 , n36009 , n24354 );
    not g5410 ( n26669 , n24221 );
    xnor g5411 ( n36072 , n42542 , n40632 );
    or g5412 ( n35917 , n42447 , n3768 );
    or g5413 ( n26262 , n5585 , n12330 );
    nor g5414 ( n32308 , n37707 , n7053 );
    or g5415 ( n34028 , n31671 , n30485 );
    or g5416 ( n13952 , n41439 , n35256 );
    nor g5417 ( n16577 , n59 , n13860 );
    or g5418 ( n35811 , n13495 , n27277 );
    and g5419 ( n36073 , n13610 , n6875 );
    nor g5420 ( n26002 , n8903 , n9171 );
    xnor g5421 ( n37277 , n19945 , n18306 );
    or g5422 ( n6935 , n12481 , n14621 );
    not g5423 ( n11747 , n32328 );
    and g5424 ( n36256 , n25031 , n7633 );
    and g5425 ( n33923 , n14890 , n27777 );
    or g5426 ( n40396 , n12547 , n15095 );
    xnor g5427 ( n31831 , n14239 , n13036 );
    xnor g5428 ( n6715 , n35727 , n23751 );
    not g5429 ( n30869 , n33811 );
    and g5430 ( n42225 , n8397 , n20414 );
    or g5431 ( n12488 , n34527 , n27105 );
    or g5432 ( n19233 , n22905 , n42783 );
    or g5433 ( n33782 , n14458 , n40702 );
    xnor g5434 ( n25347 , n14649 , n3167 );
    and g5435 ( n26588 , n20807 , n34656 );
    and g5436 ( n36757 , n37732 , n23837 );
    or g5437 ( n6530 , n15646 , n18126 );
    or g5438 ( n2220 , n4436 , n8658 );
    and g5439 ( n39772 , n23983 , n2211 );
    or g5440 ( n27774 , n24007 , n3856 );
    and g5441 ( n3424 , n7918 , n34442 );
    or g5442 ( n13119 , n29790 , n42122 );
    or g5443 ( n24325 , n9347 , n21970 );
    or g5444 ( n10823 , n5335 , n37633 );
    or g5445 ( n28833 , n17957 , n39066 );
    or g5446 ( n35776 , n898 , n15998 );
    or g5447 ( n29981 , n29593 , n35070 );
    nor g5448 ( n8109 , n23425 , n34745 );
    or g5449 ( n32366 , n38157 , n31436 );
    xnor g5450 ( n14249 , n1216 , n5079 );
    xnor g5451 ( n30787 , n42064 , n30886 );
    and g5452 ( n42265 , n36140 , n21376 );
    and g5453 ( n22218 , n25620 , n25887 );
    xnor g5454 ( n40240 , n26190 , n31959 );
    and g5455 ( n10354 , n15512 , n52 );
    or g5456 ( n29010 , n35386 , n14110 );
    or g5457 ( n10994 , n7839 , n31807 );
    xnor g5458 ( n13052 , n29347 , n36858 );
    or g5459 ( n8217 , n36930 , n14666 );
    and g5460 ( n36518 , n7348 , n15171 );
    or g5461 ( n5162 , n29533 , n25526 );
    or g5462 ( n13790 , n23374 , n40763 );
    not g5463 ( n9835 , n5540 );
    xnor g5464 ( n14034 , n27789 , n19421 );
    or g5465 ( n17236 , n35301 , n8545 );
    or g5466 ( n32391 , n21048 , n11004 );
    nor g5467 ( n41250 , n1507 , n3719 );
    not g5468 ( n13949 , n9471 );
    nor g5469 ( n9259 , n31724 , n36096 );
    xnor g5470 ( n8413 , n42863 , n40224 );
    or g5471 ( n11512 , n14129 , n26461 );
    not g5472 ( n8969 , n3186 );
    xnor g5473 ( n31018 , n12190 , n16067 );
    and g5474 ( n9865 , n230 , n28686 );
    or g5475 ( n20773 , n286 , n19559 );
    or g5476 ( n8100 , n25588 , n25943 );
    not g5477 ( n33307 , n30729 );
    and g5478 ( n26399 , n39734 , n10050 );
    xnor g5479 ( n9878 , n10535 , n28953 );
    and g5480 ( n14844 , n26039 , n33092 );
    xnor g5481 ( n2674 , n34352 , n24475 );
    xnor g5482 ( n17392 , n1301 , n11320 );
    not g5483 ( n33796 , n19508 );
    or g5484 ( n21062 , n12336 , n16487 );
    not g5485 ( n40178 , n25649 );
    not g5486 ( n22982 , n25361 );
    or g5487 ( n14023 , n37455 , n18499 );
    not g5488 ( n42070 , n4621 );
    or g5489 ( n36427 , n32087 , n13605 );
    not g5490 ( n30504 , n24587 );
    not g5491 ( n20761 , n8573 );
    or g5492 ( n14709 , n26710 , n12210 );
    xnor g5493 ( n1629 , n36628 , n36038 );
    nor g5494 ( n39665 , n25469 , n37831 );
    or g5495 ( n38965 , n32 , n946 );
    and g5496 ( n25449 , n7905 , n32115 );
    and g5497 ( n31873 , n12221 , n35157 );
    xnor g5498 ( n22274 , n7924 , n11874 );
    and g5499 ( n22569 , n28022 , n24774 );
    and g5500 ( n9632 , n2642 , n35513 );
    and g5501 ( n1418 , n3534 , n32777 );
    and g5502 ( n22249 , n20159 , n18047 );
    or g5503 ( n5255 , n6431 , n20137 );
    nor g5504 ( n29304 , n37017 , n11837 );
    or g5505 ( n8065 , n14414 , n11918 );
    not g5506 ( n42217 , n28591 );
    or g5507 ( n38472 , n36071 , n22605 );
    nor g5508 ( n7165 , n39266 , n34418 );
    and g5509 ( n3498 , n34870 , n28794 );
    or g5510 ( n7122 , n1311 , n2837 );
    or g5511 ( n2295 , n12275 , n6563 );
    not g5512 ( n1926 , n28729 );
    or g5513 ( n22600 , n39059 , n8798 );
    and g5514 ( n1906 , n40247 , n18505 );
    and g5515 ( n3198 , n37417 , n5502 );
    nor g5516 ( n10930 , n2199 , n2172 );
    or g5517 ( n17338 , n8542 , n14682 );
    or g5518 ( n24971 , n8623 , n32623 );
    xnor g5519 ( n26989 , n10716 , n40983 );
    nor g5520 ( n31409 , n11318 , n28284 );
    xnor g5521 ( n23678 , n898 , n16081 );
    not g5522 ( n38735 , n19324 );
    and g5523 ( n16028 , n42593 , n5043 );
    nor g5524 ( n20780 , n36886 , n29578 );
    and g5525 ( n31235 , n9866 , n29185 );
    or g5526 ( n23024 , n23046 , n6999 );
    xnor g5527 ( n41298 , n38667 , n37121 );
    or g5528 ( n23613 , n25371 , n15006 );
    or g5529 ( n380 , n2199 , n36491 );
    nor g5530 ( n17453 , n42515 , n39967 );
    and g5531 ( n40368 , n38914 , n20976 );
    nor g5532 ( n24233 , n37643 , n11433 );
    or g5533 ( n427 , n27695 , n33151 );
    and g5534 ( n30334 , n3762 , n34706 );
    and g5535 ( n30028 , n36448 , n28203 );
    not g5536 ( n4015 , n24577 );
    not g5537 ( n11057 , n9637 );
    xnor g5538 ( n15566 , n31989 , n36832 );
    and g5539 ( n2896 , n14921 , n15546 );
    nor g5540 ( n32699 , n14307 , n42238 );
    xnor g5541 ( n9478 , n20958 , n8234 );
    and g5542 ( n1407 , n31392 , n6428 );
    and g5543 ( n15031 , n39225 , n4472 );
    xnor g5544 ( n35381 , n36009 , n32221 );
    xnor g5545 ( n19441 , n34352 , n32237 );
    and g5546 ( n37513 , n42390 , n14919 );
    and g5547 ( n42082 , n5820 , n16077 );
    or g5548 ( n29837 , n3086 , n18308 );
    nor g5549 ( n3639 , n2375 , n20126 );
    nor g5550 ( n35927 , n33781 , n18734 );
    not g5551 ( n25291 , n40907 );
    not g5552 ( n31582 , n12180 );
    and g5553 ( n30655 , n10771 , n27176 );
    and g5554 ( n18501 , n20251 , n18580 );
    nor g5555 ( n11325 , n25817 , n2881 );
    or g5556 ( n40848 , n21075 , n6415 );
    or g5557 ( n38550 , n7802 , n30640 );
    not g5558 ( n1044 , n13979 );
    and g5559 ( n12850 , n4976 , n35520 );
    xnor g5560 ( n32694 , n28120 , n16319 );
    nor g5561 ( n26672 , n38879 , n37978 );
    and g5562 ( n20131 , n39945 , n38794 );
    not g5563 ( n36309 , n1516 );
    or g5564 ( n30609 , n11204 , n39350 );
    or g5565 ( n8748 , n38196 , n38756 );
    not g5566 ( n21439 , n22134 );
    nor g5567 ( n38638 , n20851 , n13569 );
    xnor g5568 ( n4127 , n32048 , n30155 );
    or g5569 ( n24486 , n40662 , n4023 );
    or g5570 ( n32177 , n12226 , n17061 );
    not g5571 ( n12669 , n19578 );
    not g5572 ( n36822 , n42653 );
    not g5573 ( n9940 , n7309 );
    and g5574 ( n13587 , n41423 , n40416 );
    xnor g5575 ( n1786 , n36009 , n4853 );
    or g5576 ( n16754 , n25399 , n18861 );
    or g5577 ( n25854 , n3396 , n1436 );
    not g5578 ( n6004 , n35356 );
    and g5579 ( n15958 , n39185 , n35909 );
    and g5580 ( n33964 , n11638 , n39387 );
    or g5581 ( n28018 , n20763 , n34184 );
    or g5582 ( n26233 , n18385 , n24899 );
    or g5583 ( n24084 , n19416 , n27934 );
    or g5584 ( n39630 , n41057 , n3275 );
    not g5585 ( n31431 , n24255 );
    xnor g5586 ( n15988 , n4712 , n22955 );
    or g5587 ( n12844 , n26116 , n6537 );
    or g5588 ( n20812 , n21705 , n7139 );
    or g5589 ( n3896 , n30446 , n12551 );
    or g5590 ( n15921 , n1581 , n32246 );
    or g5591 ( n5856 , n11431 , n41158 );
    not g5592 ( n31213 , n42861 );
    not g5593 ( n3077 , n34527 );
    nor g5594 ( n31141 , n5964 , n42504 );
    not g5595 ( n16234 , n3442 );
    xnor g5596 ( n4600 , n29293 , n31872 );
    nor g5597 ( n16513 , n11319 , n33497 );
    or g5598 ( n9437 , n15443 , n26927 );
    or g5599 ( n40683 , n27733 , n31828 );
    and g5600 ( n19010 , n25726 , n19317 );
    not g5601 ( n22785 , n12662 );
    and g5602 ( n13014 , n26020 , n14827 );
    and g5603 ( n30259 , n2377 , n15017 );
    or g5604 ( n16523 , n38879 , n26776 );
    not g5605 ( n12078 , n32564 );
    and g5606 ( n17002 , n2206 , n19816 );
    or g5607 ( n32690 , n14079 , n23767 );
    or g5608 ( n9915 , n15232 , n33658 );
    or g5609 ( n4234 , n28149 , n8294 );
    and g5610 ( n17829 , n39019 , n39437 );
    and g5611 ( n32700 , n26856 , n42209 );
    or g5612 ( n39441 , n15157 , n5785 );
    or g5613 ( n40460 , n3580 , n14665 );
    xnor g5614 ( n20357 , n26579 , n21538 );
    or g5615 ( n1161 , n33815 , n41331 );
    xnor g5616 ( n27825 , n21797 , n35975 );
    nor g5617 ( n6262 , n40476 , n7435 );
    nor g5618 ( n31784 , n12570 , n3148 );
    not g5619 ( n26430 , n9360 );
    and g5620 ( n3745 , n39276 , n17692 );
    xnor g5621 ( n39899 , n29476 , n34406 );
    nor g5622 ( n3977 , n21633 , n25311 );
    or g5623 ( n32491 , n20130 , n36460 );
    or g5624 ( n1538 , n38663 , n21268 );
    or g5625 ( n32349 , n36408 , n1261 );
    or g5626 ( n10283 , n5161 , n29732 );
    and g5627 ( n28025 , n18283 , n27409 );
    or g5628 ( n29341 , n34762 , n19141 );
    not g5629 ( n32194 , n11887 );
    and g5630 ( n20218 , n8134 , n42456 );
    or g5631 ( n39133 , n42549 , n41413 );
    or g5632 ( n27894 , n39672 , n2309 );
    nor g5633 ( n29555 , n5030 , n30196 );
    or g5634 ( n29908 , n34728 , n31614 );
    not g5635 ( n27116 , n31655 );
    xnor g5636 ( n29575 , n119 , n3424 );
    xnor g5637 ( n540 , n12825 , n40658 );
    or g5638 ( n23822 , n36052 , n16657 );
    or g5639 ( n9339 , n10606 , n37299 );
    xnor g5640 ( n2318 , n14953 , n15044 );
    xnor g5641 ( n24640 , n36628 , n32044 );
    or g5642 ( n24415 , n20932 , n11466 );
    or g5643 ( n851 , n32117 , n40323 );
    or g5644 ( n8819 , n21730 , n36203 );
    or g5645 ( n18711 , n25154 , n21064 );
    or g5646 ( n15666 , n38293 , n4658 );
    or g5647 ( n14867 , n38423 , n39404 );
    xnor g5648 ( n15597 , n19463 , n30470 );
    or g5649 ( n33200 , n8241 , n40354 );
    not g5650 ( n42179 , n11407 );
    nor g5651 ( n41724 , n25588 , n2124 );
    and g5652 ( n23511 , n3002 , n38838 );
    not g5653 ( n21138 , n26121 );
    or g5654 ( n29613 , n10953 , n23039 );
    xnor g5655 ( n4586 , n105 , n38160 );
    not g5656 ( n11516 , n10649 );
    xnor g5657 ( n18385 , n36625 , n11339 );
    and g5658 ( n2916 , n13259 , n854 );
    and g5659 ( n30307 , n37898 , n15411 );
    and g5660 ( n41827 , n4523 , n20187 );
    nor g5661 ( n29182 , n6465 , n17579 );
    or g5662 ( n13264 , n22191 , n17636 );
    or g5663 ( n20614 , n5881 , n7816 );
    not g5664 ( n39398 , n17601 );
    or g5665 ( n19220 , n25113 , n17445 );
    nor g5666 ( n15516 , n39774 , n38275 );
    not g5667 ( n32727 , n13009 );
    and g5668 ( n32085 , n5639 , n11361 );
    not g5669 ( n13243 , n12924 );
    nor g5670 ( n22071 , n13508 , n18286 );
    and g5671 ( n15624 , n13959 , n30279 );
    xnor g5672 ( n3864 , n34731 , n3562 );
    and g5673 ( n27410 , n12248 , n37374 );
    or g5674 ( n6461 , n32940 , n19701 );
    or g5675 ( n33701 , n35506 , n2833 );
    not g5676 ( n23505 , n12680 );
    or g5677 ( n3600 , n9937 , n11388 );
    and g5678 ( n42645 , n13728 , n727 );
    or g5679 ( n39582 , n24767 , n25933 );
    or g5680 ( n42523 , n34158 , n28420 );
    nor g5681 ( n18481 , n24726 , n2 );
    and g5682 ( n29693 , n15592 , n35351 );
    or g5683 ( n5499 , n31263 , n40859 );
    or g5684 ( n10855 , n42905 , n41413 );
    and g5685 ( n216 , n36764 , n17074 );
    not g5686 ( n26108 , n6888 );
    nor g5687 ( n10540 , n13155 , n4592 );
    or g5688 ( n6157 , n38222 , n34091 );
    xnor g5689 ( n4141 , n18702 , n25546 );
    nor g5690 ( n21330 , n25547 , n17425 );
    nor g5691 ( n25254 , n15985 , n9352 );
    not g5692 ( n38493 , n38391 );
    or g5693 ( n21317 , n37073 , n41197 );
    not g5694 ( n23574 , n19021 );
    or g5695 ( n6228 , n13470 , n42073 );
    and g5696 ( n19163 , n11244 , n23913 );
    xnor g5697 ( n25050 , n11436 , n38483 );
    or g5698 ( n8648 , n22535 , n12319 );
    or g5699 ( n29166 , n21337 , n37787 );
    and g5700 ( n29686 , n14131 , n24419 );
    and g5701 ( n27058 , n2923 , n35229 );
    xnor g5702 ( n25323 , n23511 , n19221 );
    not g5703 ( n41923 , n39392 );
    or g5704 ( n34386 , n36685 , n41622 );
    or g5705 ( n11009 , n6237 , n2728 );
    xnor g5706 ( n42441 , n10612 , n33700 );
    and g5707 ( n15743 , n28429 , n11493 );
    and g5708 ( n36716 , n30093 , n9816 );
    xnor g5709 ( n23405 , n3367 , n38770 );
    or g5710 ( n27852 , n34856 , n36261 );
    or g5711 ( n21015 , n25136 , n24467 );
    and g5712 ( n30224 , n20699 , n35295 );
    nor g5713 ( n17982 , n9030 , n29840 );
    not g5714 ( n42284 , n36371 );
    xnor g5715 ( n27519 , n6625 , n36459 );
    or g5716 ( n10174 , n32789 , n20032 );
    and g5717 ( n34819 , n32581 , n37845 );
    and g5718 ( n19406 , n226 , n38300 );
    and g5719 ( n12931 , n34266 , n20005 );
    nor g5720 ( n18871 , n16907 , n5767 );
    not g5721 ( n37044 , n13106 );
    nor g5722 ( n29661 , n6424 , n27491 );
    or g5723 ( n12124 , n9413 , n41898 );
    nor g5724 ( n6381 , n29296 , n27711 );
    nor g5725 ( n37634 , n3911 , n29764 );
    or g5726 ( n25568 , n17927 , n20784 );
    nor g5727 ( n21478 , n1457 , n11949 );
    nor g5728 ( n2203 , n2971 , n28492 );
    or g5729 ( n7171 , n31496 , n19512 );
    or g5730 ( n13508 , n35191 , n14167 );
    or g5731 ( n19923 , n19980 , n22549 );
    xnor g5732 ( n37115 , n18530 , n22564 );
    nor g5733 ( n33356 , n25602 , n10544 );
    or g5734 ( n6401 , n6874 , n23563 );
    not g5735 ( n8626 , n29731 );
    or g5736 ( n5740 , n256 , n23797 );
    and g5737 ( n24259 , n29142 , n1481 );
    and g5738 ( n27080 , n26072 , n21422 );
    not g5739 ( n28050 , n3378 );
    not g5740 ( n40298 , n9300 );
    or g5741 ( n23611 , n14506 , n41985 );
    or g5742 ( n42168 , n31513 , n9508 );
    or g5743 ( n14065 , n7166 , n34634 );
    or g5744 ( n26445 , n40467 , n19724 );
    and g5745 ( n26343 , n39021 , n34247 );
    or g5746 ( n28980 , n7196 , n15904 );
    or g5747 ( n40108 , n35534 , n35411 );
    or g5748 ( n25241 , n9747 , n15186 );
    or g5749 ( n10631 , n30945 , n16675 );
    nor g5750 ( n34001 , n21840 , n15638 );
    or g5751 ( n3826 , n30536 , n7468 );
    or g5752 ( n10021 , n26065 , n22707 );
    or g5753 ( n19439 , n37315 , n15475 );
    and g5754 ( n30978 , n19495 , n16021 );
    and g5755 ( n32957 , n16726 , n18892 );
    and g5756 ( n12970 , n15487 , n21250 );
    or g5757 ( n40179 , n21074 , n29138 );
    nor g5758 ( n23984 , n19298 , n24920 );
    and g5759 ( n42125 , n12654 , n2452 );
    xnor g5760 ( n12009 , n31973 , n942 );
    or g5761 ( n37132 , n39765 , n35037 );
    xnor g5762 ( n35011 , n25043 , n1164 );
    and g5763 ( n9549 , n26867 , n21901 );
    not g5764 ( n16910 , n37088 );
    or g5765 ( n38643 , n20030 , n6187 );
    or g5766 ( n36735 , n26917 , n3009 );
    or g5767 ( n2605 , n12345 , n33501 );
    nor g5768 ( n36873 , n736 , n33899 );
    or g5769 ( n6376 , n10506 , n23130 );
    and g5770 ( n10295 , n17868 , n31952 );
    not g5771 ( n20958 , n24876 );
    or g5772 ( n5987 , n42896 , n24877 );
    not g5773 ( n19866 , n39452 );
    nor g5774 ( n510 , n39927 , n27015 );
    or g5775 ( n7112 , n34793 , n13574 );
    nor g5776 ( n19987 , n38761 , n28651 );
    not g5777 ( n1607 , n5185 );
    not g5778 ( n32402 , n27338 );
    or g5779 ( n16763 , n17335 , n11237 );
    nor g5780 ( n15154 , n38879 , n18315 );
    nor g5781 ( n19518 , n3763 , n40414 );
    or g5782 ( n21889 , n36976 , n27021 );
    xnor g5783 ( n32930 , n13984 , n39039 );
    or g5784 ( n27999 , n13937 , n27738 );
    or g5785 ( n36907 , n37901 , n27179 );
    nor g5786 ( n5485 , n13399 , n37607 );
    nor g5787 ( n2904 , n10152 , n26407 );
    nor g5788 ( n32802 , n6663 , n22785 );
    not g5789 ( n15285 , n7702 );
    or g5790 ( n19208 , n11984 , n34470 );
    nor g5791 ( n31146 , n17647 , n36849 );
    and g5792 ( n30144 , n39424 , n7779 );
    and g5793 ( n36021 , n12292 , n24799 );
    or g5794 ( n25684 , n36490 , n12704 );
    and g5795 ( n38533 , n27633 , n6366 );
    not g5796 ( n35134 , n36630 );
    xnor g5797 ( n6952 , n25426 , n10586 );
    and g5798 ( n11218 , n3182 , n39867 );
    xnor g5799 ( n37100 , n8851 , n40334 );
    or g5800 ( n13663 , n12952 , n38448 );
    xnor g5801 ( n34143 , n32470 , n2617 );
    or g5802 ( n5098 , n18983 , n6372 );
    and g5803 ( n1286 , n15704 , n5579 );
    nor g5804 ( n32846 , n299 , n33918 );
    nor g5805 ( n7849 , n20894 , n9100 );
    and g5806 ( n18287 , n13008 , n19670 );
    or g5807 ( n34068 , n34994 , n22721 );
    nor g5808 ( n5387 , n38640 , n21460 );
    or g5809 ( n16200 , n31628 , n15525 );
    nor g5810 ( n12036 , n17393 , n30759 );
    or g5811 ( n42736 , n27924 , n6092 );
    or g5812 ( n4971 , n39788 , n34468 );
    or g5813 ( n16567 , n23331 , n23692 );
    xnor g5814 ( n39486 , n42064 , n30884 );
    nor g5815 ( n12184 , n39330 , n11200 );
    and g5816 ( n31244 , n42757 , n16579 );
    and g5817 ( n29770 , n9019 , n39049 );
    or g5818 ( n23720 , n12264 , n30620 );
    or g5819 ( n32703 , n946 , n10851 );
    or g5820 ( n14798 , n39954 , n30757 );
    or g5821 ( n19195 , n31808 , n29605 );
    xnor g5822 ( n16786 , n31353 , n10138 );
    and g5823 ( n22718 , n35168 , n22081 );
    or g5824 ( n21556 , n32952 , n33590 );
    not g5825 ( n4463 , n3458 );
    or g5826 ( n8091 , n5964 , n24926 );
    and g5827 ( n9692 , n39664 , n13096 );
    and g5828 ( n31552 , n25022 , n17470 );
    not g5829 ( n32676 , n19364 );
    or g5830 ( n30607 , n11344 , n26993 );
    not g5831 ( n14057 , n31294 );
    or g5832 ( n6535 , n30888 , n24992 );
    and g5833 ( n11731 , n35039 , n27413 );
    nor g5834 ( n17287 , n5896 , n12994 );
    not g5835 ( n39992 , n27342 );
    or g5836 ( n32383 , n20704 , n28897 );
    not g5837 ( n37212 , n10778 );
    or g5838 ( n39335 , n18263 , n5090 );
    or g5839 ( n6275 , n124 , n18622 );
    and g5840 ( n22222 , n30942 , n21298 );
    or g5841 ( n18786 , n9677 , n18797 );
    or g5842 ( n38979 , n873 , n17260 );
    and g5843 ( n18042 , n6395 , n40745 );
    xnor g5844 ( n22182 , n21484 , n7191 );
    nor g5845 ( n22617 , n41662 , n6765 );
    or g5846 ( n25746 , n10853 , n24301 );
    not g5847 ( n11533 , n36978 );
    or g5848 ( n28967 , n10646 , n19349 );
    or g5849 ( n23810 , n10242 , n22920 );
    nor g5850 ( n5136 , n34641 , n38666 );
    or g5851 ( n23759 , n36844 , n11114 );
    xnor g5852 ( n20421 , n36009 , n3719 );
    and g5853 ( n22145 , n11338 , n11742 );
    not g5854 ( n33826 , n26655 );
    not g5855 ( n32890 , n31281 );
    or g5856 ( n21606 , n28839 , n13512 );
    or g5857 ( n660 , n33774 , n24841 );
    or g5858 ( n12790 , n14690 , n2565 );
    or g5859 ( n23865 , n35679 , n32676 );
    not g5860 ( n32597 , n32105 );
    or g5861 ( n34681 , n39526 , n25742 );
    or g5862 ( n5192 , n10707 , n573 );
    and g5863 ( n33432 , n1953 , n32416 );
    not g5864 ( n22802 , n42172 );
    or g5865 ( n33832 , n5654 , n24405 );
    and g5866 ( n28545 , n4719 , n25008 );
    or g5867 ( n40040 , n14548 , n1256 );
    or g5868 ( n21543 , n40231 , n1326 );
    xnor g5869 ( n31204 , n35154 , n1261 );
    and g5870 ( n24564 , n30065 , n33103 );
    and g5871 ( n4209 , n3621 , n22163 );
    nor g5872 ( n21956 , n23377 , n31617 );
    and g5873 ( n12886 , n797 , n25023 );
    not g5874 ( n32874 , n37357 );
    or g5875 ( n10649 , n22837 , n493 );
    not g5876 ( n37509 , n24030 );
    not g5877 ( n10629 , n694 );
    and g5878 ( n799 , n36908 , n7107 );
    or g5879 ( n5225 , n31520 , n31156 );
    and g5880 ( n5277 , n35718 , n2528 );
    or g5881 ( n38109 , n39699 , n8070 );
    or g5882 ( n36449 , n38879 , n31322 );
    not g5883 ( n12218 , n3645 );
    or g5884 ( n29944 , n29906 , n10703 );
    or g5885 ( n42090 , n1913 , n37611 );
    or g5886 ( n12454 , n26947 , n37120 );
    or g5887 ( n6661 , n6673 , n24112 );
    or g5888 ( n8532 , n4157 , n33836 );
    and g5889 ( n3727 , n3475 , n28278 );
    or g5890 ( n26732 , n7265 , n9308 );
    and g5891 ( n23955 , n29460 , n12034 );
    or g5892 ( n14314 , n24393 , n29050 );
    not g5893 ( n9616 , n39082 );
    not g5894 ( n29219 , n34590 );
    or g5895 ( n10489 , n32513 , n22423 );
    nor g5896 ( n42359 , n13697 , n29902 );
    nor g5897 ( n17961 , n39712 , n20800 );
    and g5898 ( n4563 , n35440 , n13162 );
    or g5899 ( n25128 , n37337 , n32822 );
    xnor g5900 ( n32404 , n34731 , n3091 );
    and g5901 ( n12733 , n41719 , n15416 );
    and g5902 ( n17153 , n1221 , n22150 );
    or g5903 ( n15376 , n22333 , n17844 );
    nor g5904 ( n20332 , n14091 , n16006 );
    not g5905 ( n39257 , n40841 );
    or g5906 ( n20786 , n17120 , n31315 );
    or g5907 ( n3791 , n36117 , n37843 );
    xnor g5908 ( n40601 , n34352 , n18844 );
    nor g5909 ( n20568 , n37571 , n9985 );
    and g5910 ( n8409 , n38932 , n36525 );
    not g5911 ( n42852 , n19747 );
    nor g5912 ( n9868 , n2199 , n12560 );
    nor g5913 ( n19869 , n37241 , n34592 );
    or g5914 ( n37154 , n10598 , n32277 );
    or g5915 ( n1939 , n13830 , n38135 );
    nor g5916 ( n14708 , n15070 , n35673 );
    not g5917 ( n2633 , n29558 );
    or g5918 ( n29603 , n35269 , n23373 );
    nor g5919 ( n29589 , n33274 , n24116 );
    or g5920 ( n26938 , n10704 , n35944 );
    or g5921 ( n2847 , n4062 , n23694 );
    not g5922 ( n17256 , n13300 );
    or g5923 ( n31219 , n24781 , n5850 );
    or g5924 ( n35308 , n11920 , n40259 );
    and g5925 ( n38258 , n10556 , n23395 );
    not g5926 ( n1555 , n42331 );
    or g5927 ( n22685 , n24745 , n31081 );
    or g5928 ( n22293 , n34318 , n38423 );
    or g5929 ( n5835 , n26059 , n23210 );
    not g5930 ( n25425 , n41189 );
    or g5931 ( n3190 , n7725 , n8992 );
    or g5932 ( n15028 , n23055 , n36530 );
    nor g5933 ( n7231 , n32898 , n12754 );
    xnor g5934 ( n11982 , n37436 , n38994 );
    or g5935 ( n4415 , n40316 , n9194 );
    and g5936 ( n40724 , n36562 , n26049 );
    or g5937 ( n4346 , n3583 , n42228 );
    and g5938 ( n30997 , n9651 , n14968 );
    or g5939 ( n23587 , n1971 , n36158 );
    xnor g5940 ( n31945 , n26904 , n940 );
    or g5941 ( n4051 , n8626 , n1164 );
    nor g5942 ( n36760 , n17120 , n7921 );
    or g5943 ( n35488 , n41339 , n27226 );
    or g5944 ( n2866 , n5170 , n31466 );
    or g5945 ( n40085 , n12876 , n6992 );
    and g5946 ( n26025 , n8411 , n16206 );
    or g5947 ( n15412 , n7255 , n34658 );
    and g5948 ( n19087 , n28515 , n2913 );
    or g5949 ( n42412 , n10219 , n6042 );
    not g5950 ( n19497 , n31157 );
    xnor g5951 ( n2917 , n33958 , n21356 );
    or g5952 ( n22839 , n36858 , n19104 );
    or g5953 ( n539 , n23472 , n38740 );
    nor g5954 ( n25648 , n38157 , n38120 );
    not g5955 ( n9057 , n36895 );
    or g5956 ( n31796 , n14519 , n37344 );
    xnor g5957 ( n39189 , n35727 , n24369 );
    or g5958 ( n2790 , n20321 , n25303 );
    and g5959 ( n932 , n6641 , n32845 );
    xnor g5960 ( n34956 , n6104 , n6008 );
    xnor g5961 ( n15790 , n21957 , n19517 );
    xnor g5962 ( n16002 , n5234 , n25816 );
    or g5963 ( n6336 , n1167 , n29690 );
    or g5964 ( n22849 , n5585 , n39038 );
    xnor g5965 ( n1708 , n38398 , n40991 );
    and g5966 ( n5660 , n5468 , n25085 );
    or g5967 ( n22648 , n37334 , n25626 );
    or g5968 ( n34554 , n31153 , n171 );
    nor g5969 ( n4788 , n1507 , n14238 );
    and g5970 ( n32114 , n27651 , n37508 );
    nor g5971 ( n4862 , n9930 , n24291 );
    nor g5972 ( n22550 , n7858 , n22939 );
    xnor g5973 ( n17097 , n9250 , n42546 );
    not g5974 ( n10819 , n27892 );
    or g5975 ( n41832 , n4783 , n3530 );
    and g5976 ( n34829 , n28315 , n14430 );
    and g5977 ( n40232 , n40003 , n4785 );
    or g5978 ( n38523 , n42665 , n36235 );
    and g5979 ( n7542 , n34854 , n13071 );
    nor g5980 ( n18087 , n22387 , n33029 );
    xnor g5981 ( n1705 , n7450 , n5807 );
    or g5982 ( n39307 , n13176 , n38245 );
    nor g5983 ( n6012 , n23994 , n29569 );
    or g5984 ( n14833 , n35948 , n33926 );
    and g5985 ( n37223 , n36804 , n20895 );
    xnor g5986 ( n30708 , n34471 , n39086 );
    and g5987 ( n9114 , n41840 , n16126 );
    or g5988 ( n4507 , n5896 , n22618 );
    and g5989 ( n41605 , n33871 , n7233 );
    or g5990 ( n13241 , n36434 , n15093 );
    and g5991 ( n6025 , n725 , n39540 );
    not g5992 ( n13301 , n20140 );
    not g5993 ( n38142 , n12745 );
    or g5994 ( n41952 , n41026 , n14443 );
    or g5995 ( n33929 , n33328 , n22664 );
    nor g5996 ( n9658 , n29499 , n10055 );
    and g5997 ( n26203 , n26428 , n5970 );
    or g5998 ( n26966 , n7187 , n19702 );
    xnor g5999 ( n2533 , n642 , n33981 );
    not g6000 ( n26348 , n6448 );
    or g6001 ( n41267 , n18914 , n13883 );
    and g6002 ( n12913 , n16132 , n33764 );
    nor g6003 ( n18377 , n42627 , n31783 );
    and g6004 ( n5232 , n22408 , n25138 );
    or g6005 ( n10658 , n17118 , n17173 );
    not g6006 ( n26789 , n16664 );
    and g6007 ( n19135 , n39110 , n17995 );
    and g6008 ( n10197 , n4938 , n35015 );
    not g6009 ( n6558 , n36731 );
    or g6010 ( n25983 , n33825 , n1717 );
    or g6011 ( n42232 , n9579 , n30671 );
    and g6012 ( n20460 , n35945 , n1182 );
    or g6013 ( n26724 , n23043 , n15301 );
    or g6014 ( n17938 , n21290 , n2095 );
    and g6015 ( n2354 , n1124 , n6678 );
    or g6016 ( n26957 , n13182 , n39676 );
    or g6017 ( n3575 , n18243 , n7737 );
    or g6018 ( n23629 , n7360 , n28999 );
    not g6019 ( n40331 , n17737 );
    not g6020 ( n29856 , n17301 );
    nor g6021 ( n35782 , n29714 , n34874 );
    not g6022 ( n4084 , n32824 );
    nor g6023 ( n37693 , n21090 , n28529 );
    or g6024 ( n33390 , n23368 , n40450 );
    or g6025 ( n25141 , n41583 , n29986 );
    or g6026 ( n23721 , n3823 , n11768 );
    xnor g6027 ( n18596 , n21545 , n33981 );
    xnor g6028 ( n22368 , n29740 , n36244 );
    or g6029 ( n7059 , n9772 , n16159 );
    or g6030 ( n10071 , n25266 , n17249 );
    nor g6031 ( n23753 , n14052 , n23977 );
    or g6032 ( n38765 , n33218 , n27353 );
    not g6033 ( n42902 , n7548 );
    or g6034 ( n32790 , n19260 , n21933 );
    or g6035 ( n22808 , n32100 , n16408 );
    xnor g6036 ( n12207 , n27396 , n477 );
    or g6037 ( n6585 , n2972 , n375 );
    xnor g6038 ( n24030 , n23431 , n31168 );
    or g6039 ( n9221 , n31854 , n3646 );
    or g6040 ( n10977 , n36896 , n30839 );
    and g6041 ( n24305 , n15323 , n35290 );
    or g6042 ( n22917 , n29834 , n17079 );
    not g6043 ( n23261 , n22160 );
    not g6044 ( n14115 , n23873 );
    or g6045 ( n23791 , n36344 , n3062 );
    nor g6046 ( n35777 , n25723 , n18783 );
    and g6047 ( n17347 , n40201 , n40642 );
    or g6048 ( n30594 , n10462 , n12842 );
    not g6049 ( n23462 , n7508 );
    xnor g6050 ( n35937 , n37403 , n1281 );
    and g6051 ( n35429 , n3147 , n34621 );
    not g6052 ( n1030 , n41289 );
    xnor g6053 ( n41220 , n4218 , n2726 );
    or g6054 ( n36900 , n27502 , n35210 );
    xnor g6055 ( n27421 , n28648 , n39413 );
    or g6056 ( n5559 , n6512 , n27023 );
    or g6057 ( n35979 , n18650 , n30089 );
    and g6058 ( n30886 , n41744 , n26717 );
    or g6059 ( n23413 , n13122 , n19848 );
    not g6060 ( n25594 , n32371 );
    xnor g6061 ( n42435 , n11785 , n41227 );
    or g6062 ( n6594 , n25101 , n34570 );
    nor g6063 ( n29696 , n35509 , n17569 );
    xnor g6064 ( n14665 , n10723 , n221 );
    or g6065 ( n2602 , n11629 , n26945 );
    and g6066 ( n8966 , n7717 , n25983 );
    or g6067 ( n32270 , n1732 , n32689 );
    or g6068 ( n11945 , n29337 , n8378 );
    and g6069 ( n28511 , n27299 , n9081 );
    or g6070 ( n40613 , n38157 , n29300 );
    or g6071 ( n22322 , n17640 , n4723 );
    or g6072 ( n32466 , n31263 , n3256 );
    and g6073 ( n26229 , n41786 , n31528 );
    xnor g6074 ( n29559 , n31161 , n15865 );
    and g6075 ( n41158 , n8168 , n35110 );
    nor g6076 ( n34249 , n5349 , n29636 );
    or g6077 ( n14830 , n35483 , n23821 );
    and g6078 ( n4374 , n16459 , n37844 );
    nor g6079 ( n18507 , n38879 , n39570 );
    or g6080 ( n24945 , n35575 , n41696 );
    or g6081 ( n30098 , n6510 , n40965 );
    and g6082 ( n14983 , n31450 , n14512 );
    and g6083 ( n9187 , n6901 , n41078 );
    nor g6084 ( n9857 , n6565 , n13314 );
    or g6085 ( n42752 , n10326 , n39273 );
    not g6086 ( n17138 , n28431 );
    not g6087 ( n39158 , n29394 );
    and g6088 ( n10854 , n6455 , n21020 );
    xnor g6089 ( n1072 , n5660 , n25588 );
    and g6090 ( n35459 , n21411 , n6681 );
    not g6091 ( n31764 , n27744 );
    buf g6092 ( n24077 , n12006 );
    and g6093 ( n18522 , n23454 , n33879 );
    not g6094 ( n6077 , n9110 );
    and g6095 ( n36802 , n10893 , n27166 );
    nor g6096 ( n15355 , n19813 , n17401 );
    or g6097 ( n26608 , n34003 , n32936 );
    or g6098 ( n28818 , n20037 , n328 );
    nor g6099 ( n33408 , n38084 , n30283 );
    xnor g6100 ( n29724 , n37969 , n967 );
    nor g6101 ( n7525 , n27722 , n10533 );
    nor g6102 ( n28398 , n6278 , n27444 );
    or g6103 ( n18733 , n9594 , n42446 );
    or g6104 ( n14352 , n25360 , n29952 );
    or g6105 ( n27128 , n30382 , n792 );
    not g6106 ( n4676 , n16 );
    and g6107 ( n16293 , n19483 , n8285 );
    or g6108 ( n6334 , n21113 , n19788 );
    not g6109 ( n12286 , n21029 );
    or g6110 ( n38959 , n40914 , n25528 );
    xnor g6111 ( n7422 , n19183 , n15837 );
    or g6112 ( n38187 , n30400 , n14569 );
    or g6113 ( n27253 , n6023 , n31545 );
    or g6114 ( n36753 , n35320 , n18758 );
    or g6115 ( n7809 , n11765 , n18393 );
    or g6116 ( n30331 , n9164 , n36235 );
    or g6117 ( n39628 , n14145 , n21725 );
    or g6118 ( n24666 , n37859 , n36848 );
    or g6119 ( n34335 , n3093 , n27809 );
    or g6120 ( n31348 , n42553 , n16856 );
    not g6121 ( n8319 , n32442 );
    not g6122 ( n20556 , n6552 );
    xnor g6123 ( n28155 , n25525 , n8379 );
    or g6124 ( n38076 , n6754 , n23314 );
    and g6125 ( n26934 , n37265 , n42233 );
    not g6126 ( n14817 , n27216 );
    xnor g6127 ( n37413 , n35727 , n10075 );
    or g6128 ( n32441 , n20332 , n5908 );
    or g6129 ( n26530 , n22000 , n32540 );
    or g6130 ( n25022 , n33486 , n30071 );
    not g6131 ( n34817 , n20361 );
    or g6132 ( n15446 , n16032 , n38662 );
    or g6133 ( n25017 , n41526 , n40821 );
    and g6134 ( n28880 , n40925 , n13214 );
    nor g6135 ( n22405 , n2961 , n15568 );
    or g6136 ( n40528 , n4222 , n1688 );
    or g6137 ( n4170 , n35032 , n9040 );
    and g6138 ( n38754 , n7060 , n19926 );
    or g6139 ( n19016 , n34013 , n15531 );
    or g6140 ( n33831 , n7265 , n8297 );
    not g6141 ( n36078 , n5613 );
    and g6142 ( n37585 , n22658 , n9933 );
    and g6143 ( n15651 , n32134 , n25227 );
    or g6144 ( n40166 , n30132 , n5916 );
    or g6145 ( n38883 , n42195 , n25784 );
    not g6146 ( n31290 , n27419 );
    or g6147 ( n18258 , n12446 , n28986 );
    or g6148 ( n25638 , n2478 , n10520 );
    and g6149 ( n14745 , n34580 , n22280 );
    not g6150 ( n3433 , n26818 );
    nor g6151 ( n2395 , n12389 , n24123 );
    xnor g6152 ( n20522 , n28781 , n22227 );
    and g6153 ( n7181 , n26383 , n831 );
    or g6154 ( n36688 , n2355 , n18750 );
    nor g6155 ( n28779 , n21766 , n34777 );
    or g6156 ( n3401 , n11163 , n23857 );
    and g6157 ( n8034 , n22428 , n41412 );
    not g6158 ( n9331 , n38862 );
    and g6159 ( n31129 , n39838 , n37164 );
    or g6160 ( n26223 , n5722 , n27938 );
    or g6161 ( n36392 , n30037 , n15397 );
    xnor g6162 ( n39718 , n26210 , n15610 );
    or g6163 ( n19543 , n42838 , n17514 );
    or g6164 ( n34005 , n17256 , n19971 );
    or g6165 ( n11338 , n36408 , n27194 );
    nor g6166 ( n9141 , n13769 , n25651 );
    not g6167 ( n16897 , n26344 );
    and g6168 ( n17001 , n14231 , n5562 );
    or g6169 ( n3153 , n18343 , n31005 );
    or g6170 ( n7517 , n9752 , n37996 );
    or g6171 ( n13184 , n34960 , n13509 );
    not g6172 ( n11855 , n24687 );
    not g6173 ( n904 , n294 );
    xnor g6174 ( n40939 , n21973 , n35511 );
    xnor g6175 ( n8527 , n23135 , n21447 );
    xnor g6176 ( n8072 , n5144 , n42616 );
    xnor g6177 ( n34937 , n22820 , n40736 );
    and g6178 ( n37584 , n24567 , n2906 );
    or g6179 ( n42583 , n39078 , n33798 );
    not g6180 ( n13284 , n42719 );
    and g6181 ( n10792 , n28873 , n5366 );
    and g6182 ( n40326 , n20150 , n42141 );
    xnor g6183 ( n34725 , n20411 , n2143 );
    xnor g6184 ( n28995 , n19926 , n7060 );
    or g6185 ( n37046 , n4223 , n34384 );
    or g6186 ( n4038 , n16996 , n2897 );
    xnor g6187 ( n7245 , n21178 , n9896 );
    nor g6188 ( n15318 , n24289 , n41642 );
    or g6189 ( n4230 , n29451 , n14773 );
    not g6190 ( n20457 , n32361 );
    nor g6191 ( n10770 , n37452 , n21168 );
    or g6192 ( n6471 , n27663 , n42672 );
    or g6193 ( n42298 , n16836 , n5832 );
    xnor g6194 ( n13620 , n23804 , n2403 );
    or g6195 ( n25134 , n30446 , n10991 );
    or g6196 ( n39338 , n28611 , n8306 );
    and g6197 ( n17794 , n36164 , n13168 );
    xnor g6198 ( n10058 , n16883 , n40546 );
    not g6199 ( n12293 , n41541 );
    nor g6200 ( n845 , n27681 , n12537 );
    or g6201 ( n11788 , n8680 , n28209 );
    or g6202 ( n9440 , n25372 , n4270 );
    and g6203 ( n17934 , n41104 , n4285 );
    and g6204 ( n21695 , n24761 , n24014 );
    nor g6205 ( n21494 , n11469 , n18472 );
    or g6206 ( n13708 , n12530 , n12307 );
    or g6207 ( n13826 , n6810 , n25279 );
    nor g6208 ( n124 , n21972 , n18829 );
    nor g6209 ( n27903 , n41662 , n14623 );
    not g6210 ( n34921 , n29351 );
    or g6211 ( n16946 , n33174 , n7650 );
    xnor g6212 ( n24129 , n42064 , n14963 );
    and g6213 ( n2992 , n34509 , n27821 );
    not g6214 ( n3306 , n29225 );
    xnor g6215 ( n22246 , n12063 , n41410 );
    and g6216 ( n40527 , n6972 , n35097 );
    or g6217 ( n27832 , n28984 , n7289 );
    or g6218 ( n40620 , n13469 , n24592 );
    and g6219 ( n3548 , n27253 , n33045 );
    or g6220 ( n37391 , n35963 , n27121 );
    xnor g6221 ( n31457 , n33253 , n32587 );
    xnor g6222 ( n37050 , n26955 , n20155 );
    xnor g6223 ( n3483 , n36513 , n7706 );
    not g6224 ( n13939 , n6335 );
    or g6225 ( n25678 , n42870 , n34688 );
    nor g6226 ( n2819 , n31279 , n35468 );
    or g6227 ( n38145 , n5018 , n13698 );
    nor g6228 ( n24277 , n10211 , n18062 );
    and g6229 ( n18504 , n35724 , n11983 );
    and g6230 ( n3439 , n39890 , n8131 );
    nor g6231 ( n831 , n13697 , n30893 );
    not g6232 ( n41007 , n26669 );
    and g6233 ( n23977 , n36785 , n2558 );
    not g6234 ( n23378 , n28630 );
    or g6235 ( n1943 , n24894 , n5989 );
    not g6236 ( n10740 , n33839 );
    and g6237 ( n11749 , n23054 , n41687 );
    xnor g6238 ( n34103 , n10535 , n1407 );
    nor g6239 ( n21838 , n40962 , n35128 );
    xnor g6240 ( n16137 , n34875 , n4568 );
    and g6241 ( n24431 , n749 , n30783 );
    or g6242 ( n27262 , n37317 , n36242 );
    or g6243 ( n23755 , n40450 , n27312 );
    and g6244 ( n16166 , n11007 , n27382 );
    and g6245 ( n13560 , n15530 , n4263 );
    or g6246 ( n7051 , n37847 , n32121 );
    not g6247 ( n33733 , n21407 );
    and g6248 ( n22131 , n8939 , n13990 );
    and g6249 ( n25551 , n39290 , n31820 );
    and g6250 ( n9874 , n3428 , n21763 );
    not g6251 ( n7071 , n20398 );
    not g6252 ( n40173 , n28325 );
    not g6253 ( n17715 , n12275 );
    xnor g6254 ( n19465 , n19077 , n16950 );
    xnor g6255 ( n38542 , n33884 , n34537 );
    not g6256 ( n36532 , n36420 );
    nor g6257 ( n29419 , n4725 , n19369 );
    xnor g6258 ( n14209 , n32662 , n2199 );
    or g6259 ( n23952 , n24289 , n41215 );
    xnor g6260 ( n18998 , n28869 , n7356 );
    xnor g6261 ( n15886 , n16693 , n36716 );
    not g6262 ( n40540 , n26566 );
    or g6263 ( n31349 , n1507 , n27260 );
    and g6264 ( n17574 , n10438 , n37501 );
    and g6265 ( n31186 , n39259 , n21437 );
    or g6266 ( n18414 , n29303 , n27567 );
    or g6267 ( n17047 , n41170 , n29404 );
    xnor g6268 ( n12253 , n36899 , n18098 );
    not g6269 ( n8540 , n8025 );
    nor g6270 ( n16962 , n1971 , n28337 );
    not g6271 ( n26935 , n12318 );
    or g6272 ( n17763 , n34762 , n22550 );
    not g6273 ( n7321 , n4782 );
    not g6274 ( n10078 , n34030 );
    or g6275 ( n30261 , n35298 , n9967 );
    and g6276 ( n16740 , n7185 , n1230 );
    nor g6277 ( n10657 , n34292 , n15212 );
    or g6278 ( n39017 , n42507 , n31834 );
    nor g6279 ( n28708 , n15051 , n38037 );
    nor g6280 ( n41754 , n11566 , n28544 );
    or g6281 ( n39228 , n40129 , n16028 );
    nor g6282 ( n32712 , n35009 , n29585 );
    and g6283 ( n24119 , n6213 , n31285 );
    xnor g6284 ( n16131 , n29083 , n32717 );
    and g6285 ( n16643 , n9529 , n29263 );
    and g6286 ( n30569 , n13206 , n33749 );
    or g6287 ( n26598 , n41892 , n20711 );
    or g6288 ( n29951 , n19915 , n28028 );
    xnor g6289 ( n24645 , n42064 , n16227 );
    nor g6290 ( n25152 , n37582 , n7874 );
    not g6291 ( n9964 , n26655 );
    and g6292 ( n14669 , n5152 , n18046 );
    nor g6293 ( n10115 , n40768 , n24172 );
    not g6294 ( n38416 , n28057 );
    and g6295 ( n27705 , n8458 , n5382 );
    or g6296 ( n40880 , n20174 , n34497 );
    or g6297 ( n4268 , n21125 , n4512 );
    or g6298 ( n14881 , n23082 , n14711 );
    and g6299 ( n34269 , n21762 , n15386 );
    or g6300 ( n39148 , n6869 , n951 );
    not g6301 ( n35154 , n32119 );
    xnor g6302 ( n4054 , n18558 , n21546 );
    xnor g6303 ( n7311 , n26579 , n11229 );
    or g6304 ( n35168 , n40110 , n31529 );
    or g6305 ( n12597 , n2616 , n19798 );
    nor g6306 ( n33105 , n4140 , n2876 );
    not g6307 ( n42585 , n23273 );
    or g6308 ( n13403 , n10576 , n40200 );
    not g6309 ( n5905 , n24121 );
    or g6310 ( n33136 , n36585 , n40948 );
    or g6311 ( n42366 , n30857 , n38766 );
    or g6312 ( n17635 , n363 , n6189 );
    and g6313 ( n1972 , n14092 , n20266 );
    and g6314 ( n13361 , n4265 , n39071 );
    nor g6315 ( n1641 , n27593 , n22090 );
    nor g6316 ( n23262 , n14471 , n12619 );
    or g6317 ( n10138 , n13393 , n26788 );
    not g6318 ( n42076 , n20224 );
    xnor g6319 ( n28712 , n20245 , n13347 );
    not g6320 ( n32731 , n14962 );
    nor g6321 ( n18103 , n29057 , n5774 );
    or g6322 ( n3449 , n422 , n39924 );
    or g6323 ( n33155 , n36169 , n41767 );
    xnor g6324 ( n25595 , n17225 , n39940 );
    not g6325 ( n3543 , n26655 );
    and g6326 ( n27392 , n4234 , n18198 );
    and g6327 ( n28683 , n7063 , n11154 );
    not g6328 ( n17393 , n16623 );
    not g6329 ( n17108 , n19366 );
    not g6330 ( n6394 , n37746 );
    xnor g6331 ( n4620 , n34844 , n11577 );
    and g6332 ( n939 , n8252 , n6103 );
    and g6333 ( n11768 , n36735 , n30180 );
    or g6334 ( n7184 , n22401 , n27732 );
    not g6335 ( n13470 , n17107 );
    and g6336 ( n2765 , n17479 , n2798 );
    and g6337 ( n37204 , n5196 , n6343 );
    xnor g6338 ( n36804 , n32297 , n12507 );
    not g6339 ( n5367 , n39742 );
    or g6340 ( n42759 , n22993 , n36030 );
    or g6341 ( n37165 , n41922 , n33236 );
    or g6342 ( n874 , n8972 , n36947 );
    or g6343 ( n3592 , n18514 , n13658 );
    not g6344 ( n16410 , n13859 );
    or g6345 ( n11578 , n30691 , n7214 );
    or g6346 ( n23896 , n21732 , n2537 );
    and g6347 ( n11845 , n18791 , n1401 );
    and g6348 ( n29778 , n21990 , n31684 );
    or g6349 ( n7495 , n24223 , n13940 );
    nor g6350 ( n2228 , n1500 , n7653 );
    and g6351 ( n3606 , n29146 , n42053 );
    or g6352 ( n24651 , n5465 , n3308 );
    or g6353 ( n1634 , n33330 , n12766 );
    or g6354 ( n42112 , n6165 , n32894 );
    or g6355 ( n24649 , n19778 , n27448 );
    not g6356 ( n23535 , n32384 );
    or g6357 ( n22060 , n28281 , n7507 );
    and g6358 ( n12482 , n30426 , n1204 );
    not g6359 ( n22519 , n25308 );
    nor g6360 ( n3703 , n16728 , n17488 );
    xnor g6361 ( n6747 , n35727 , n23795 );
    not g6362 ( n27028 , n3416 );
    or g6363 ( n17689 , n14370 , n1043 );
    and g6364 ( n4650 , n30332 , n5924 );
    xnor g6365 ( n37597 , n566 , n18868 );
    and g6366 ( n8216 , n27067 , n30770 );
    or g6367 ( n11865 , n26845 , n24965 );
    and g6368 ( n34643 , n16233 , n25769 );
    or g6369 ( n24587 , n12716 , n1639 );
    and g6370 ( n24490 , n33905 , n41478 );
    and g6371 ( n14260 , n15415 , n24517 );
    nor g6372 ( n8682 , n23431 , n15897 );
    or g6373 ( n4457 , n4140 , n12982 );
    and g6374 ( n7972 , n26241 , n7328 );
    or g6375 ( n4663 , n41802 , n25806 );
    and g6376 ( n31771 , n8323 , n15223 );
    or g6377 ( n34666 , n22369 , n26147 );
    not g6378 ( n2858 , n6408 );
    not g6379 ( n22934 , n8465 );
    or g6380 ( n41733 , n19636 , n18722 );
    xnor g6381 ( n2891 , n12900 , n9570 );
    or g6382 ( n6681 , n14945 , n34392 );
    and g6383 ( n7551 , n18843 , n25347 );
    or g6384 ( n37164 , n4680 , n34955 );
    nor g6385 ( n23290 , n18320 , n13486 );
    or g6386 ( n26297 , n40870 , n20971 );
    and g6387 ( n19090 , n28358 , n20673 );
    or g6388 ( n28719 , n15332 , n42492 );
    and g6389 ( n16784 , n32891 , n39046 );
    not g6390 ( n27037 , n8588 );
    and g6391 ( n25778 , n3095 , n38460 );
    and g6392 ( n451 , n30374 , n8895 );
    or g6393 ( n4693 , n8535 , n32532 );
    or g6394 ( n204 , n34918 , n11379 );
    nor g6395 ( n23098 , n14707 , n41678 );
    nor g6396 ( n25991 , n25588 , n7783 );
    xnor g6397 ( n42796 , n37670 , n11350 );
    or g6398 ( n11427 , n2199 , n32662 );
    not g6399 ( n34866 , n12464 );
    and g6400 ( n14829 , n19657 , n39089 );
    and g6401 ( n28492 , n12922 , n7005 );
    or g6402 ( n40609 , n29717 , n28507 );
    or g6403 ( n41675 , n26354 , n8505 );
    or g6404 ( n34915 , n11551 , n19702 );
    xnor g6405 ( n8786 , n20366 , n5896 );
    or g6406 ( n40747 , n39624 , n40329 );
    xnor g6407 ( n8230 , n42064 , n28200 );
    or g6408 ( n23054 , n16388 , n41649 );
    or g6409 ( n37260 , n17976 , n35918 );
    or g6410 ( n27185 , n454 , n38412 );
    and g6411 ( n10009 , n8120 , n17270 );
    and g6412 ( n19445 , n29839 , n30900 );
    and g6413 ( n21754 , n35077 , n29662 );
    or g6414 ( n13975 , n9509 , n31948 );
    not g6415 ( n32453 , n17486 );
    or g6416 ( n31558 , n7595 , n18578 );
    xnor g6417 ( n12144 , n22915 , n37427 );
    or g6418 ( n7366 , n22056 , n32773 );
    and g6419 ( n10146 , n4188 , n11975 );
    and g6420 ( n28994 , n15615 , n26957 );
    and g6421 ( n24374 , n27117 , n4662 );
    nor g6422 ( n16321 , n16829 , n14517 );
    nor g6423 ( n28295 , n37241 , n15553 );
    nor g6424 ( n41394 , n3850 , n35576 );
    nor g6425 ( n40536 , n25340 , n39179 );
    or g6426 ( n22547 , n16738 , n34908 );
    nor g6427 ( n2334 , n6248 , n37744 );
    xnor g6428 ( n11458 , n18696 , n2280 );
    not g6429 ( n25624 , n24747 );
    and g6430 ( n32798 , n39244 , n26541 );
    or g6431 ( n33769 , n14794 , n21232 );
    xnor g6432 ( n30873 , n16693 , n4499 );
    not g6433 ( n36983 , n30959 );
    or g6434 ( n16261 , n29000 , n7321 );
    nor g6435 ( n41392 , n36977 , n3344 );
    not g6436 ( n31268 , n8342 );
    or g6437 ( n35088 , n5933 , n20495 );
    nor g6438 ( n46 , n2199 , n5863 );
    or g6439 ( n7465 , n18816 , n32317 );
    not g6440 ( n3824 , n19862 );
    xnor g6441 ( n35684 , n14338 , n40400 );
    or g6442 ( n19241 , n23068 , n30652 );
    or g6443 ( n34062 , n7000 , n33845 );
    xnor g6444 ( n13487 , n30264 , n41373 );
    and g6445 ( n22122 , n15372 , n19992 );
    xnor g6446 ( n29990 , n34056 , n14525 );
    or g6447 ( n8635 , n12028 , n27181 );
    and g6448 ( n41555 , n10043 , n13927 );
    and g6449 ( n17277 , n27929 , n12544 );
    or g6450 ( n7614 , n8980 , n31728 );
    not g6451 ( n10169 , n24647 );
    not g6452 ( n9247 , n8780 );
    or g6453 ( n28768 , n2183 , n2516 );
    and g6454 ( n22351 , n20569 , n6112 );
    nor g6455 ( n13150 , n4410 , n11504 );
    nor g6456 ( n31834 , n5826 , n7878 );
    not g6457 ( n31091 , n12465 );
    and g6458 ( n13468 , n11387 , n32911 );
    not g6459 ( n16682 , n13668 );
    nor g6460 ( n738 , n16482 , n15220 );
    or g6461 ( n13558 , n32311 , n12152 );
    and g6462 ( n42634 , n21580 , n39650 );
    or g6463 ( n29315 , n6130 , n9784 );
    xnor g6464 ( n23601 , n31363 , n5224 );
    or g6465 ( n18046 , n12424 , n26494 );
    not g6466 ( n7265 , n3457 );
    not g6467 ( n30117 , n19136 );
    nor g6468 ( n28746 , n15289 , n20227 );
    or g6469 ( n11873 , n16109 , n22186 );
    not g6470 ( n25573 , n13886 );
    or g6471 ( n22008 , n18353 , n27540 );
    or g6472 ( n35716 , n28784 , n8886 );
    or g6473 ( n16574 , n37044 , n10035 );
    nor g6474 ( n22765 , n19221 , n2694 );
    not g6475 ( n27333 , n30697 );
    and g6476 ( n41879 , n4674 , n14801 );
    nor g6477 ( n40611 , n29859 , n21265 );
    and g6478 ( n29934 , n21765 , n1951 );
    or g6479 ( n36680 , n1880 , n41270 );
    and g6480 ( n34209 , n15313 , n3344 );
    and g6481 ( n31561 , n22769 , n40747 );
    xnor g6482 ( n12468 , n542 , n38690 );
    nor g6483 ( n15584 , n26689 , n23077 );
    or g6484 ( n9762 , n33912 , n41079 );
    xnor g6485 ( n22269 , n8019 , n7564 );
    or g6486 ( n22477 , n32092 , n34742 );
    or g6487 ( n40215 , n15049 , n12220 );
    xnor g6488 ( n18392 , n28252 , n30169 );
    nor g6489 ( n14263 , n36758 , n12448 );
    or g6490 ( n16589 , n27001 , n37252 );
    not g6491 ( n6929 , n41321 );
    or g6492 ( n33156 , n31613 , n1597 );
    or g6493 ( n35579 , n39556 , n40857 );
    or g6494 ( n18497 , n20086 , n32585 );
    not g6495 ( n18697 , n34357 );
    xnor g6496 ( n25810 , n39094 , n32738 );
    and g6497 ( n42020 , n38885 , n23356 );
    not g6498 ( n11436 , n34565 );
    not g6499 ( n23667 , n32371 );
    xnor g6500 ( n38342 , n11436 , n30349 );
    or g6501 ( n17705 , n40637 , n1967 );
    xnor g6502 ( n19291 , n10226 , n20069 );
    nor g6503 ( n28688 , n41616 , n31669 );
    nor g6504 ( n7469 , n18067 , n5758 );
    not g6505 ( n32433 , n28248 );
    or g6506 ( n37614 , n14607 , n14569 );
    xnor g6507 ( n5215 , n30043 , n7639 );
    and g6508 ( n19915 , n32636 , n20149 );
    nor g6509 ( n35738 , n26621 , n22488 );
    not g6510 ( n19969 , n33854 );
    or g6511 ( n31031 , n13361 , n22929 );
    nor g6512 ( n38306 , n1683 , n26809 );
    or g6513 ( n20592 , n37193 , n34754 );
    nor g6514 ( n42487 , n38917 , n5736 );
    not g6515 ( n10023 , n17239 );
    xnor g6516 ( n26154 , n28489 , n16287 );
    or g6517 ( n672 , n21532 , n42544 );
    or g6518 ( n36191 , n23359 , n19267 );
    not g6519 ( n41896 , n26229 );
    not g6520 ( n38597 , n2743 );
    not g6521 ( n17613 , n32457 );
    or g6522 ( n32129 , n9880 , n28539 );
    not g6523 ( n17423 , n1534 );
    or g6524 ( n27995 , n1461 , n19041 );
    or g6525 ( n15975 , n23472 , n13277 );
    or g6526 ( n36512 , n4535 , n610 );
    nor g6527 ( n16286 , n42435 , n26821 );
    and g6528 ( n42476 , n17769 , n10809 );
    not g6529 ( n11993 , n33200 );
    or g6530 ( n41936 , n18914 , n32136 );
    or g6531 ( n28119 , n14622 , n13186 );
    xnor g6532 ( n2861 , n30853 , n41534 );
    or g6533 ( n36981 , n14308 , n35303 );
    nor g6534 ( n35330 , n28917 , n19445 );
    nor g6535 ( n6306 , n27117 , n4662 );
    not g6536 ( n14649 , n36012 );
    or g6537 ( n12826 , n20173 , n18532 );
    not g6538 ( n17260 , n3404 );
    and g6539 ( n24606 , n33037 , n15465 );
    or g6540 ( n34262 , n42306 , n21856 );
    or g6541 ( n14636 , n9809 , n809 );
    not g6542 ( n28427 , n18196 );
    not g6543 ( n6102 , n3179 );
    nor g6544 ( n40926 , n7421 , n8299 );
    and g6545 ( n11931 , n37700 , n29601 );
    xnor g6546 ( n5594 , n11436 , n23542 );
    not g6547 ( n3602 , n20363 );
    or g6548 ( n2598 , n2425 , n24179 );
    and g6549 ( n14142 , n21843 , n29951 );
    or g6550 ( n4678 , n37031 , n11734 );
    or g6551 ( n19384 , n14707 , n18756 );
    or g6552 ( n22048 , n18911 , n6247 );
    not g6553 ( n1987 , n38226 );
    nor g6554 ( n5141 , n14217 , n24693 );
    or g6555 ( n2898 , n41458 , n23760 );
    and g6556 ( n20630 , n38934 , n37390 );
    xnor g6557 ( n13877 , n11570 , n33329 );
    nor g6558 ( n4711 , n42326 , n40268 );
    not g6559 ( n24527 , n6379 );
    or g6560 ( n5080 , n5896 , n28078 );
    and g6561 ( n37252 , n2222 , n32493 );
    or g6562 ( n38471 , n13786 , n14851 );
    and g6563 ( n34909 , n22546 , n25654 );
    xnor g6564 ( n37124 , n17137 , n38797 );
    not g6565 ( n39367 , n4165 );
    or g6566 ( n28238 , n11208 , n37787 );
    not g6567 ( n22105 , n4653 );
    xnor g6568 ( n21867 , n20019 , n24744 );
    or g6569 ( n22779 , n5964 , n31051 );
    or g6570 ( n42293 , n35732 , n36219 );
    and g6571 ( n31579 , n41707 , n8918 );
    and g6572 ( n37013 , n22421 , n15886 );
    xnor g6573 ( n10565 , n34562 , n40277 );
    or g6574 ( n5155 , n13361 , n14897 );
    and g6575 ( n40951 , n19304 , n1887 );
    not g6576 ( n2214 , n33220 );
    not g6577 ( n2174 , n4822 );
    or g6578 ( n23166 , n31523 , n22177 );
    or g6579 ( n32704 , n25993 , n11194 );
    and g6580 ( n38840 , n15417 , n3999 );
    or g6581 ( n18407 , n8817 , n22797 );
    or g6582 ( n24144 , n25209 , n38438 );
    xnor g6583 ( n4187 , n8872 , n37866 );
    and g6584 ( n13835 , n40254 , n13129 );
    and g6585 ( n1574 , n10200 , n31292 );
    xnor g6586 ( n27297 , n2293 , n19749 );
    nor g6587 ( n33259 , n42373 , n33799 );
    or g6588 ( n4214 , n3477 , n25303 );
    xnor g6589 ( n42744 , n15972 , n19922 );
    or g6590 ( n38418 , n13188 , n12152 );
    nor g6591 ( n33456 , n6547 , n36040 );
    nor g6592 ( n12739 , n41293 , n33482 );
    and g6593 ( n26435 , n34783 , n7049 );
    and g6594 ( n26601 , n13164 , n27497 );
    or g6595 ( n27472 , n32397 , n33765 );
    or g6596 ( n10185 , n13280 , n14560 );
    or g6597 ( n8644 , n20233 , n33212 );
    or g6598 ( n24487 , n5559 , n8986 );
    nor g6599 ( n37243 , n15003 , n14761 );
    nor g6600 ( n34853 , n31099 , n12819 );
    and g6601 ( n16782 , n32853 , n10749 );
    or g6602 ( n275 , n27466 , n9947 );
    nor g6603 ( n41384 , n13207 , n8880 );
    or g6604 ( n6036 , n32697 , n7066 );
    not g6605 ( n33279 , n9705 );
    and g6606 ( n30519 , n14334 , n26709 );
    and g6607 ( n1409 , n35488 , n27896 );
    or g6608 ( n28304 , n31997 , n41062 );
    nor g6609 ( n7269 , n41545 , n41528 );
    or g6610 ( n16632 , n8610 , n14952 );
    nor g6611 ( n16140 , n1617 , n33864 );
    xnor g6612 ( n24118 , n14315 , n39821 );
    and g6613 ( n23174 , n9984 , n12117 );
    and g6614 ( n20373 , n23680 , n18804 );
    xnor g6615 ( n14022 , n20487 , n40917 );
    or g6616 ( n27864 , n14749 , n34289 );
    not g6617 ( n31389 , n37686 );
    and g6618 ( n24279 , n34137 , n34671 );
    or g6619 ( n30319 , n32174 , n24934 );
    or g6620 ( n3310 , n26555 , n1416 );
    or g6621 ( n37417 , n25742 , n41734 );
    or g6622 ( n29128 , n3337 , n32869 );
    nor g6623 ( n36799 , n32225 , n1802 );
    or g6624 ( n11479 , n29023 , n12896 );
    not g6625 ( n42425 , n2101 );
    or g6626 ( n35816 , n28727 , n35219 );
    not g6627 ( n10530 , n34383 );
    or g6628 ( n31053 , n27090 , n32733 );
    and g6629 ( n16877 , n7943 , n35214 );
    or g6630 ( n31713 , n27530 , n34682 );
    nor g6631 ( n8992 , n9729 , n18728 );
    nor g6632 ( n32642 , n35285 , n29939 );
    or g6633 ( n11209 , n38879 , n656 );
    and g6634 ( n34004 , n41557 , n16641 );
    and g6635 ( n42368 , n30076 , n19403 );
    and g6636 ( n13860 , n15469 , n36057 );
    and g6637 ( n18132 , n18518 , n35904 );
    and g6638 ( n24836 , n6899 , n1822 );
    not g6639 ( n22984 , n10262 );
    nor g6640 ( n2131 , n36297 , n25571 );
    xnor g6641 ( n42666 , n25041 , n42489 );
    or g6642 ( n11730 , n29903 , n37767 );
    not g6643 ( n27761 , n7069 );
    nor g6644 ( n6867 , n33669 , n14297 );
    or g6645 ( n34982 , n34998 , n13566 );
    not g6646 ( n14888 , n15978 );
    or g6647 ( n9675 , n8212 , n26551 );
    and g6648 ( n5017 , n26503 , n9440 );
    xnor g6649 ( n20940 , n4960 , n24911 );
    not g6650 ( n39517 , n30532 );
    and g6651 ( n6683 , n38609 , n1170 );
    and g6652 ( n29249 , n4322 , n22400 );
    or g6653 ( n2271 , n15935 , n22379 );
    and g6654 ( n27507 , n20464 , n30524 );
    or g6655 ( n37928 , n6929 , n1038 );
    or g6656 ( n31976 , n11629 , n33566 );
    or g6657 ( n28925 , n27902 , n24575 );
    or g6658 ( n39549 , n28633 , n25440 );
    xnor g6659 ( n1811 , n20208 , n33284 );
    not g6660 ( n811 , n25520 );
    xnor g6661 ( n30419 , n26997 , n28567 );
    xnor g6662 ( n19351 , n40391 , n4241 );
    or g6663 ( n7067 , n42393 , n1303 );
    not g6664 ( n28075 , n36546 );
    or g6665 ( n15909 , n13868 , n5215 );
    xnor g6666 ( n12114 , n11436 , n24 );
    nor g6667 ( n8715 , n27137 , n38001 );
    and g6668 ( n10087 , n4898 , n30366 );
    or g6669 ( n18657 , n9763 , n33366 );
    not g6670 ( n19323 , n4705 );
    not g6671 ( n12990 , n34481 );
    not g6672 ( n31767 , n22303 );
    nor g6673 ( n11140 , n22089 , n34135 );
    or g6674 ( n11298 , n11410 , n40538 );
    and g6675 ( n5023 , n9453 , n9815 );
    and g6676 ( n35044 , n30887 , n17928 );
    nor g6677 ( n28140 , n1971 , n16047 );
    not g6678 ( n15254 , n34601 );
    or g6679 ( n791 , n32893 , n38603 );
    not g6680 ( n22385 , n41525 );
    xnor g6681 ( n16422 , n31368 , n5911 );
    xnor g6682 ( n10308 , n17222 , n34565 );
    or g6683 ( n16886 , n31647 , n2095 );
    or g6684 ( n7437 , n17951 , n33182 );
    or g6685 ( n8229 , n5828 , n33233 );
    and g6686 ( n35463 , n15042 , n42415 );
    not g6687 ( n302 , n35307 );
    or g6688 ( n33165 , n7652 , n6791 );
    and g6689 ( n22928 , n35388 , n5309 );
    nor g6690 ( n23640 , n24549 , n41103 );
    nor g6691 ( n30669 , n35347 , n27538 );
    nor g6692 ( n34198 , n19045 , n7167 );
    and g6693 ( n29162 , n26462 , n1711 );
    or g6694 ( n4456 , n15385 , n17035 );
    or g6695 ( n18849 , n3931 , n9909 );
    and g6696 ( n29069 , n31196 , n42168 );
    and g6697 ( n38553 , n23587 , n8856 );
    and g6698 ( n1653 , n23124 , n16167 );
    or g6699 ( n27279 , n8469 , n30055 );
    xnor g6700 ( n31686 , n3413 , n13062 );
    not g6701 ( n25349 , n12625 );
    not g6702 ( n11067 , n38901 );
    and g6703 ( n14416 , n35853 , n32752 );
    xnor g6704 ( n20506 , n28614 , n3595 );
    and g6705 ( n19254 , n23167 , n38069 );
    or g6706 ( n6644 , n31263 , n12234 );
    and g6707 ( n13577 , n39784 , n34734 );
    nor g6708 ( n9172 , n23535 , n22815 );
    or g6709 ( n13969 , n37092 , n35155 );
    xnor g6710 ( n21787 , n17137 , n7473 );
    and g6711 ( n14711 , n35570 , n10300 );
    or g6712 ( n38501 , n4654 , n14749 );
    not g6713 ( n14395 , n30721 );
    or g6714 ( n31044 , n38227 , n25078 );
    and g6715 ( n16315 , n40188 , n17517 );
    or g6716 ( n42760 , n32276 , n34818 );
    and g6717 ( n42470 , n30120 , n2275 );
    not g6718 ( n35995 , n30105 );
    and g6719 ( n9753 , n15817 , n42181 );
    and g6720 ( n35706 , n17792 , n30127 );
    xnor g6721 ( n33418 , n36973 , n12915 );
    xnor g6722 ( n17181 , n5073 , n4700 );
    or g6723 ( n37935 , n31784 , n21268 );
    nor g6724 ( n34748 , n24442 , n13985 );
    and g6725 ( n12249 , n23629 , n5641 );
    or g6726 ( n19301 , n26927 , n38100 );
    xnor g6727 ( n20887 , n34698 , n32771 );
    and g6728 ( n8086 , n16176 , n6276 );
    nor g6729 ( n25965 , n13609 , n32755 );
    xnor g6730 ( n20882 , n9240 , n30312 );
    or g6731 ( n36464 , n644 , n18180 );
    or g6732 ( n30145 , n11866 , n8074 );
    or g6733 ( n40000 , n21994 , n26340 );
    and g6734 ( n26968 , n20272 , n26405 );
    not g6735 ( n5573 , n18979 );
    not g6736 ( n15269 , n25746 );
    not g6737 ( n32082 , n27514 );
    or g6738 ( n33861 , n26862 , n40276 );
    or g6739 ( n38616 , n34565 , n3316 );
    not g6740 ( n30902 , n11830 );
    and g6741 ( n37851 , n39356 , n34714 );
    xnor g6742 ( n26826 , n24265 , n14232 );
    and g6743 ( n41097 , n31621 , n41782 );
    or g6744 ( n15962 , n33072 , n21916 );
    or g6745 ( n9103 , n10169 , n40901 );
    and g6746 ( n28434 , n843 , n11681 );
    nor g6747 ( n29336 , n18500 , n36900 );
    or g6748 ( n31496 , n15186 , n32028 );
    xnor g6749 ( n35839 , n38251 , n7267 );
    xnor g6750 ( n31410 , n22152 , n15008 );
    and g6751 ( n11061 , n40666 , n77 );
    nor g6752 ( n6459 , n21705 , n21845 );
    or g6753 ( n28616 , n1180 , n11754 );
    or g6754 ( n27174 , n36641 , n572 );
    or g6755 ( n34145 , n36014 , n36134 );
    or g6756 ( n29953 , n19740 , n8312 );
    and g6757 ( n17678 , n8405 , n3358 );
    or g6758 ( n31036 , n38311 , n19589 );
    or g6759 ( n8522 , n2399 , n5038 );
    not g6760 ( n17038 , n35455 );
    or g6761 ( n28747 , n20724 , n21856 );
    or g6762 ( n20136 , n17838 , n6481 );
    or g6763 ( n22374 , n30693 , n39804 );
    or g6764 ( n35973 , n6905 , n11095 );
    and g6765 ( n1436 , n29466 , n12287 );
    or g6766 ( n26207 , n11568 , n21111 );
    or g6767 ( n41451 , n6636 , n34924 );
    and g6768 ( n36162 , n22534 , n5114 );
    nor g6769 ( n35080 , n24745 , n1857 );
    and g6770 ( n25464 , n35832 , n24962 );
    and g6771 ( n18313 , n18848 , n33393 );
    or g6772 ( n15699 , n9508 , n19284 );
    and g6773 ( n33494 , n368 , n11919 );
    nor g6774 ( n14690 , n14871 , n25949 );
    or g6775 ( n23687 , n11008 , n34587 );
    and g6776 ( n28348 , n2787 , n25962 );
    or g6777 ( n26458 , n14407 , n21939 );
    nor g6778 ( n16181 , n35172 , n19981 );
    and g6779 ( n6042 , n25554 , n30707 );
    or g6780 ( n35641 , n23563 , n28701 );
    nor g6781 ( n37837 , n12009 , n25555 );
    and g6782 ( n40401 , n23451 , n22434 );
    or g6783 ( n37148 , n15096 , n38217 );
    and g6784 ( n41223 , n5969 , n30776 );
    and g6785 ( n22389 , n19427 , n40734 );
    and g6786 ( n22997 , n20573 , n24829 );
    or g6787 ( n36503 , n6613 , n4625 );
    and g6788 ( n35270 , n22114 , n34802 );
    and g6789 ( n12545 , n8725 , n6616 );
    xnor g6790 ( n2455 , n40833 , n22125 );
    or g6791 ( n14452 , n22201 , n36418 );
    or g6792 ( n31187 , n37520 , n29816 );
    not g6793 ( n22520 , n6108 );
    not g6794 ( n6131 , n150 );
    or g6795 ( n17146 , n5543 , n26510 );
    not g6796 ( n38878 , n30462 );
    nor g6797 ( n40115 , n42069 , n13697 );
    not g6798 ( n13331 , n31077 );
    or g6799 ( n5488 , n7664 , n29367 );
    or g6800 ( n34902 , n34054 , n5585 );
    or g6801 ( n22507 , n6658 , n36433 );
    nor g6802 ( n19432 , n19025 , n40726 );
    or g6803 ( n16087 , n12355 , n7253 );
    or g6804 ( n16698 , n20331 , n11984 );
    nor g6805 ( n19158 , n20134 , n27985 );
    or g6806 ( n2159 , n24772 , n19701 );
    or g6807 ( n10759 , n29891 , n16345 );
    or g6808 ( n29689 , n9957 , n18881 );
    and g6809 ( n27060 , n26195 , n20329 );
    not g6810 ( n433 , n42016 );
    or g6811 ( n1628 , n31452 , n40432 );
    xnor g6812 ( n29911 , n4546 , n32327 );
    or g6813 ( n20372 , n15254 , n31651 );
    not g6814 ( n31050 , n42355 );
    or g6815 ( n35513 , n8871 , n25704 );
    or g6816 ( n20158 , n34052 , n31368 );
    and g6817 ( n25102 , n21911 , n1530 );
    and g6818 ( n40428 , n40005 , n39084 );
    or g6819 ( n16409 , n25704 , n15318 );
    or g6820 ( n16457 , n30152 , n17404 );
    xnor g6821 ( n5975 , n35867 , n33482 );
    nor g6822 ( n38053 , n33926 , n6898 );
    nor g6823 ( n4264 , n7281 , n26336 );
    or g6824 ( n26110 , n726 , n22639 );
    or g6825 ( n29159 , n10625 , n42840 );
    not g6826 ( n38711 , n39832 );
    or g6827 ( n38561 , n42691 , n94 );
    or g6828 ( n23095 , n37505 , n16465 );
    not g6829 ( n3542 , n18832 );
    or g6830 ( n17807 , n38665 , n41923 );
    or g6831 ( n8305 , n26653 , n36410 );
    and g6832 ( n26776 , n28797 , n22006 );
    or g6833 ( n26385 , n42862 , n34858 );
    and g6834 ( n6016 , n21648 , n10712 );
    or g6835 ( n25031 , n24847 , n33526 );
    or g6836 ( n37998 , n13885 , n26772 );
    nor g6837 ( n5149 , n26818 , n12860 );
    and g6838 ( n13525 , n10713 , n32734 );
    or g6839 ( n29618 , n20141 , n20734 );
    or g6840 ( n31952 , n19156 , n22858 );
    or g6841 ( n1963 , n17506 , n34561 );
    or g6842 ( n10843 , n1609 , n18102 );
    or g6843 ( n10634 , n14489 , n9649 );
    or g6844 ( n40360 , n4842 , n35045 );
    not g6845 ( n15010 , n21306 );
    or g6846 ( n30747 , n41479 , n23877 );
    or g6847 ( n18899 , n20209 , n42478 );
    not g6848 ( n9668 , n1478 );
    or g6849 ( n24110 , n30170 , n25142 );
    nor g6850 ( n34468 , n14490 , n6563 );
    not g6851 ( n14696 , n24000 );
    nor g6852 ( n4963 , n41698 , n21114 );
    not g6853 ( n42780 , n42650 );
    or g6854 ( n13405 , n28153 , n17071 );
    nor g6855 ( n22778 , n2292 , n3402 );
    or g6856 ( n35388 , n39501 , n20696 );
    and g6857 ( n1192 , n23823 , n33983 );
    or g6858 ( n38895 , n36179 , n4660 );
    and g6859 ( n18716 , n13801 , n21055 );
    and g6860 ( n8602 , n37209 , n39982 );
    not g6861 ( n20185 , n8911 );
    xnor g6862 ( n16732 , n42064 , n12546 );
    xnor g6863 ( n22534 , n22899 , n4688 );
    not g6864 ( n35443 , n27570 );
    xnor g6865 ( n17200 , n31099 , n10222 );
    or g6866 ( n27400 , n35309 , n30097 );
    and g6867 ( n12395 , n16087 , n36129 );
    or g6868 ( n19738 , n37427 , n21942 );
    or g6869 ( n3440 , n5769 , n8239 );
    not g6870 ( n2535 , n24447 );
    or g6871 ( n18037 , n33419 , n16818 );
    not g6872 ( n29052 , n13140 );
    and g6873 ( n18188 , n10970 , n4351 );
    not g6874 ( n8276 , n6021 );
    and g6875 ( n1724 , n6995 , n41626 );
    or g6876 ( n30560 , n8025 , n11257 );
    or g6877 ( n25962 , n5257 , n28887 );
    and g6878 ( n575 , n16329 , n34455 );
    or g6879 ( n34724 , n14777 , n30842 );
    and g6880 ( n37637 , n40558 , n12682 );
    not g6881 ( n13657 , n15166 );
    or g6882 ( n27770 , n9349 , n9738 );
    and g6883 ( n15766 , n41489 , n34246 );
    nor g6884 ( n11718 , n708 , n29965 );
    or g6885 ( n37620 , n42460 , n12095 );
    or g6886 ( n15042 , n23274 , n12087 );
    or g6887 ( n3422 , n5619 , n16495 );
    or g6888 ( n32773 , n27841 , n11050 );
    not g6889 ( n16544 , n14068 );
    xnor g6890 ( n21012 , n20487 , n11192 );
    or g6891 ( n5697 , n24453 , n23547 );
    and g6892 ( n33239 , n17056 , n16346 );
    or g6893 ( n11359 , n15866 , n23943 );
    xnor g6894 ( n8810 , n42715 , n1273 );
    and g6895 ( n22910 , n15764 , n13274 );
    xnor g6896 ( n21264 , n33584 , n38144 );
    and g6897 ( n3562 , n16963 , n7108 );
    and g6898 ( n40151 , n24833 , n17095 );
    and g6899 ( n15294 , n14977 , n32864 );
    nor g6900 ( n42820 , n26803 , n30205 );
    xnor g6901 ( n14650 , n26907 , n30986 );
    or g6902 ( n37272 , n14471 , n31127 );
    or g6903 ( n3404 , n27310 , n41643 );
    xnor g6904 ( n28276 , n31099 , n575 );
    nor g6905 ( n17702 , n32916 , n14714 );
    or g6906 ( n17210 , n30039 , n34522 );
    or g6907 ( n6007 , n2719 , n32923 );
    xnor g6908 ( n669 , n28443 , n20821 );
    xnor g6909 ( n29922 , n35646 , n7324 );
    and g6910 ( n25790 , n33994 , n7940 );
    or g6911 ( n9976 , n26714 , n15632 );
    or g6912 ( n15083 , n16598 , n39256 );
    and g6913 ( n39191 , n15055 , n9239 );
    not g6914 ( n37942 , n25644 );
    xnor g6915 ( n3378 , n912 , n17120 );
    or g6916 ( n23346 , n5536 , n7244 );
    not g6917 ( n33901 , n26949 );
    or g6918 ( n27167 , n13367 , n38533 );
    not g6919 ( n4839 , n12308 );
    or g6920 ( n28915 , n25459 , n328 );
    not g6921 ( n31334 , n40119 );
    and g6922 ( n32820 , n17960 , n16486 );
    or g6923 ( n29301 , n37043 , n34091 );
    xnor g6924 ( n40238 , n8063 , n9117 );
    and g6925 ( n41553 , n24113 , n11428 );
    or g6926 ( n37613 , n19573 , n33740 );
    or g6927 ( n41412 , n7839 , n26171 );
    or g6928 ( n37409 , n15556 , n41927 );
    or g6929 ( n41806 , n2599 , n7349 );
    or g6930 ( n11851 , n13780 , n13894 );
    or g6931 ( n21714 , n18998 , n41513 );
    not g6932 ( n2572 , n41464 );
    or g6933 ( n8118 , n18080 , n1387 );
    or g6934 ( n11441 , n42368 , n17254 );
    or g6935 ( n15458 , n28143 , n12492 );
    or g6936 ( n40106 , n39330 , n38998 );
    not g6937 ( n4907 , n36010 );
    and g6938 ( n32722 , n17379 , n38361 );
    or g6939 ( n17421 , n21687 , n41354 );
    xnor g6940 ( n9050 , n5891 , n39576 );
    xnor g6941 ( n32176 , n3146 , n1251 );
    not g6942 ( n1013 , n22134 );
    nor g6943 ( n41776 , n36117 , n15167 );
    or g6944 ( n36728 , n19702 , n7695 );
    or g6945 ( n4179 , n2472 , n8113 );
    and g6946 ( n37679 , n26566 , n41778 );
    or g6947 ( n947 , n4843 , n12579 );
    and g6948 ( n29092 , n27024 , n24489 );
    or g6949 ( n27338 , n20165 , n25950 );
    or g6950 ( n29860 , n29254 , n12706 );
    or g6951 ( n120 , n8192 , n26670 );
    not g6952 ( n35217 , n40299 );
    and g6953 ( n3554 , n23215 , n4380 );
    not g6954 ( n13299 , n2085 );
    or g6955 ( n32853 , n9151 , n25546 );
    not g6956 ( n30555 , n40387 );
    not g6957 ( n8182 , n33889 );
    or g6958 ( n33765 , n935 , n41527 );
    or g6959 ( n12331 , n23844 , n40588 );
    not g6960 ( n33735 , n32766 );
    xnor g6961 ( n26091 , n40 , n1668 );
    xnor g6962 ( n19945 , n10256 , n18898 );
    nor g6963 ( n25529 , n29265 , n21445 );
    or g6964 ( n40143 , n29974 , n4488 );
    xnor g6965 ( n41375 , n3032 , n42548 );
    or g6966 ( n39397 , n9383 , n6512 );
    nor g6967 ( n4667 , n4091 , n8133 );
    and g6968 ( n7013 , n24122 , n24435 );
    and g6969 ( n14859 , n5195 , n23494 );
    or g6970 ( n37095 , n3473 , n30242 );
    xnor g6971 ( n3822 , n3277 , n24885 );
    or g6972 ( n35947 , n14604 , n4180 );
    or g6973 ( n652 , n18242 , n32750 );
    or g6974 ( n852 , n12511 , n3270 );
    nor g6975 ( n13535 , n13174 , n22249 );
    xnor g6976 ( n15601 , n3125 , n4041 );
    or g6977 ( n6877 , n26886 , n7114 );
    xnor g6978 ( n47 , n19300 , n41676 );
    and g6979 ( n21002 , n40834 , n27074 );
    or g6980 ( n26054 , n8696 , n2527 );
    nor g6981 ( n4107 , n39266 , n16315 );
    or g6982 ( n17043 , n33817 , n21960 );
    and g6983 ( n28971 , n31210 , n19827 );
    xnor g6984 ( n30485 , n7661 , n31463 );
    or g6985 ( n649 , n5602 , n15780 );
    not g6986 ( n31284 , n27447 );
    or g6987 ( n17882 , n24053 , n1648 );
    or g6988 ( n36785 , n35087 , n36507 );
    or g6989 ( n36679 , n388 , n34267 );
    or g6990 ( n39538 , n34634 , n10546 );
    and g6991 ( n13509 , n19626 , n38692 );
    and g6992 ( n42357 , n20563 , n5875 );
    not g6993 ( n27769 , n7825 );
    nor g6994 ( n17950 , n17039 , n42890 );
    and g6995 ( n40446 , n5834 , n16376 );
    nor g6996 ( n23437 , n24048 , n14228 );
    nor g6997 ( n12369 , n2856 , n2312 );
    or g6998 ( n35568 , n2181 , n5713 );
    and g6999 ( n28231 , n19386 , n5690 );
    or g7000 ( n3022 , n38556 , n16643 );
    and g7001 ( n3278 , n37719 , n11397 );
    and g7002 ( n35371 , n19799 , n8882 );
    or g7003 ( n15124 , n19253 , n25424 );
    and g7004 ( n33653 , n5371 , n8606 );
    and g7005 ( n25674 , n42339 , n5963 );
    or g7006 ( n3177 , n16736 , n16227 );
    or g7007 ( n32723 , n34141 , n7376 );
    nor g7008 ( n10532 , n18051 , n5042 );
    nor g7009 ( n11139 , n2257 , n1181 );
    and g7010 ( n16146 , n5998 , n29128 );
    or g7011 ( n23014 , n10688 , n20174 );
    and g7012 ( n37056 , n7908 , n4179 );
    or g7013 ( n27469 , n30101 , n35713 );
    xnor g7014 ( n28706 , n32591 , n35494 );
    not g7015 ( n16590 , n22361 );
    or g7016 ( n38923 , n32100 , n23177 );
    or g7017 ( n31022 , n37868 , n18091 );
    or g7018 ( n32385 , n33643 , n2345 );
    or g7019 ( n37125 , n22193 , n256 );
    or g7020 ( n25725 , n29989 , n21807 );
    or g7021 ( n22786 , n10009 , n12669 );
    nor g7022 ( n1882 , n38836 , n25583 );
    and g7023 ( n8040 , n4547 , n38000 );
    xnor g7024 ( n38156 , n784 , n38039 );
    or g7025 ( n35024 , n29135 , n19158 );
    xnor g7026 ( n36607 , n14758 , n3247 );
    or g7027 ( n30663 , n29479 , n36848 );
    and g7028 ( n27326 , n28342 , n6121 );
    xnor g7029 ( n945 , n16998 , n15948 );
    or g7030 ( n7491 , n30502 , n16771 );
    and g7031 ( n12698 , n23526 , n21009 );
    not g7032 ( n31775 , n33974 );
    xnor g7033 ( n19981 , n16998 , n24271 );
    nor g7034 ( n1314 , n2199 , n25401 );
    not g7035 ( n32100 , n1794 );
    or g7036 ( n41469 , n40277 , n14668 );
    xnor g7037 ( n36836 , n29712 , n7356 );
    and g7038 ( n30210 , n14832 , n5145 );
    or g7039 ( n12023 , n37010 , n10926 );
    not g7040 ( n38408 , n32660 );
    or g7041 ( n34667 , n36584 , n41038 );
    nor g7042 ( n37840 , n10135 , n18077 );
    and g7043 ( n40486 , n9871 , n38790 );
    xnor g7044 ( n36778 , n5144 , n25656 );
    or g7045 ( n14713 , n14139 , n4897 );
    nor g7046 ( n30019 , n20411 , n12284 );
    nor g7047 ( n36949 , n21891 , n13135 );
    not g7048 ( n14578 , n9385 );
    nor g7049 ( n13024 , n15437 , n38963 );
    or g7050 ( n33538 , n33216 , n36176 );
    not g7051 ( n5961 , n40604 );
    or g7052 ( n21058 , n25850 , n25847 );
    and g7053 ( n22815 , n32238 , n24137 );
    xnor g7054 ( n42739 , n36998 , n159 );
    or g7055 ( n11371 , n28989 , n3223 );
    or g7056 ( n25510 , n24953 , n11417 );
    xnor g7057 ( n20286 , n41636 , n6449 );
    nor g7058 ( n27458 , n24553 , n9339 );
    or g7059 ( n36043 , n28707 , n33261 );
    nor g7060 ( n8188 , n13389 , n187 );
    nor g7061 ( n9092 , n9953 , n7013 );
    or g7062 ( n11010 , n19089 , n37253 );
    or g7063 ( n17728 , n36844 , n35782 );
    or g7064 ( n15920 , n18095 , n31326 );
    or g7065 ( n23820 , n11798 , n29008 );
    and g7066 ( n25108 , n26313 , n11858 );
    or g7067 ( n21731 , n32109 , n11455 );
    not g7068 ( n23491 , n27555 );
    xnor g7069 ( n27368 , n4784 , n16136 );
    or g7070 ( n39271 , n38249 , n35617 );
    not g7071 ( n33720 , n659 );
    not g7072 ( n8017 , n30305 );
    or g7073 ( n40020 , n33407 , n22906 );
    not g7074 ( n36899 , n27764 );
    not g7075 ( n40389 , n22310 );
    nor g7076 ( n34232 , n7990 , n24462 );
    or g7077 ( n36375 , n9427 , n37893 );
    or g7078 ( n22620 , n732 , n35337 );
    nor g7079 ( n41130 , n5398 , n24254 );
    or g7080 ( n35172 , n27719 , n23935 );
    or g7081 ( n7806 , n3582 , n30744 );
    not g7082 ( n13696 , n40772 );
    or g7083 ( n34506 , n21037 , n34790 );
    or g7084 ( n654 , n4619 , n10413 );
    and g7085 ( n24006 , n37281 , n5809 );
    xnor g7086 ( n36615 , n9827 , n29320 );
    xnor g7087 ( n27102 , n15936 , n41812 );
    or g7088 ( n27382 , n12031 , n20420 );
    xnor g7089 ( n28680 , n28981 , n37133 );
    or g7090 ( n42103 , n29782 , n196 );
    or g7091 ( n36706 , n19753 , n17936 );
    xnor g7092 ( n31121 , n32379 , n4082 );
    or g7093 ( n5116 , n30013 , n23703 );
    or g7094 ( n11406 , n26094 , n37273 );
    or g7095 ( n23220 , n40619 , n4775 );
    not g7096 ( n19459 , n11525 );
    or g7097 ( n1777 , n328 , n17664 );
    xnor g7098 ( n15568 , n42567 , n18243 );
    xnor g7099 ( n36123 , n9775 , n41103 );
    and g7100 ( n8535 , n25237 , n8217 );
    and g7101 ( n23782 , n35555 , n28808 );
    not g7102 ( n39720 , n31569 );
    or g7103 ( n36209 , n17393 , n17396 );
    xnor g7104 ( n4118 , n23080 , n16092 );
    or g7105 ( n1118 , n29314 , n26437 );
    not g7106 ( n34785 , n13893 );
    xnor g7107 ( n15372 , n31099 , n22985 );
    or g7108 ( n34803 , n39149 , n36675 );
    and g7109 ( n35378 , n12971 , n31359 );
    nor g7110 ( n13226 , n34565 , n22186 );
    and g7111 ( n27447 , n33593 , n15559 );
    or g7112 ( n16758 , n441 , n177 );
    or g7113 ( n34130 , n6632 , n37149 );
    or g7114 ( n1125 , n21294 , n29144 );
    not g7115 ( n16216 , n40635 );
    and g7116 ( n33127 , n10954 , n32951 );
    nor g7117 ( n19649 , n18974 , n31767 );
    and g7118 ( n3690 , n4780 , n22893 );
    nor g7119 ( n32663 , n5168 , n746 );
    or g7120 ( n26412 , n20856 , n27504 );
    or g7121 ( n31536 , n32965 , n19643 );
    or g7122 ( n32162 , n7175 , n26536 );
    or g7123 ( n33913 , n9151 , n12975 );
    and g7124 ( n31948 , n16023 , n31396 );
    and g7125 ( n19152 , n24149 , n39319 );
    or g7126 ( n22895 , n1733 , n14308 );
    xnor g7127 ( n14169 , n7943 , n22250 );
    nor g7128 ( n19280 , n10276 , n19341 );
    or g7129 ( n1676 , n29968 , n17829 );
    and g7130 ( n10268 , n17376 , n9027 );
    not g7131 ( n18134 , n21515 );
    and g7132 ( n32411 , n38624 , n28176 );
    and g7133 ( n42321 , n7721 , n37398 );
    or g7134 ( n40156 , n9319 , n3940 );
    nor g7135 ( n31190 , n5270 , n6140 );
    and g7136 ( n33394 , n20688 , n36069 );
    or g7137 ( n28927 , n2184 , n10330 );
    not g7138 ( n34559 , n33915 );
    nor g7139 ( n17908 , n21592 , n42840 );
    xnor g7140 ( n5712 , n6508 , n30503 );
    xnor g7141 ( n26489 , n4244 , n34506 );
    and g7142 ( n39995 , n18246 , n42639 );
    or g7143 ( n41473 , n15936 , n30386 );
    not g7144 ( n4552 , n16566 );
    xnor g7145 ( n17904 , n2637 , n17940 );
    not g7146 ( n8087 , n14219 );
    nor g7147 ( n37150 , n14052 , n20207 );
    or g7148 ( n20432 , n28919 , n32095 );
    and g7149 ( n23523 , n1875 , n28802 );
    or g7150 ( n28923 , n34994 , n10690 );
    nor g7151 ( n35272 , n7769 , n29760 );
    or g7152 ( n32131 , n18088 , n4718 );
    not g7153 ( n37005 , n67 );
    or g7154 ( n41434 , n38475 , n34561 );
    nor g7155 ( n26286 , n8044 , n33091 );
    or g7156 ( n23516 , n38004 , n31557 );
    nor g7157 ( n25716 , n29535 , n34346 );
    or g7158 ( n5130 , n14407 , n29177 );
    or g7159 ( n18565 , n1701 , n11258 );
    and g7160 ( n4361 , n17098 , n10432 );
    and g7161 ( n31339 , n13208 , n23050 );
    or g7162 ( n25019 , n33673 , n33301 );
    nor g7163 ( n25009 , n6762 , n1733 );
    nor g7164 ( n19258 , n26643 , n12969 );
    or g7165 ( n35182 , n6075 , n37633 );
    not g7166 ( n30764 , n32667 );
    nor g7167 ( n25557 , n3769 , n28359 );
    not g7168 ( n24116 , n19571 );
    xnor g7169 ( n9582 , n6375 , n29471 );
    or g7170 ( n2925 , n34775 , n23646 );
    and g7171 ( n4321 , n40353 , n30229 );
    and g7172 ( n21947 , n35481 , n7527 );
    and g7173 ( n1367 , n9751 , n33381 );
    or g7174 ( n23825 , n25788 , n12220 );
    nor g7175 ( n6582 , n36828 , n18765 );
    or g7176 ( n9893 , n4880 , n10496 );
    xnor g7177 ( n28601 , n10078 , n36335 );
    or g7178 ( n3488 , n13558 , n28251 );
    or g7179 ( n38564 , n5881 , n28494 );
    or g7180 ( n37021 , n14811 , n38798 );
    or g7181 ( n3847 , n11685 , n12286 );
    and g7182 ( n2584 , n35436 , n15243 );
    nor g7183 ( n14992 , n23491 , n6672 );
    nor g7184 ( n12203 , n35748 , n2549 );
    xnor g7185 ( n1616 , n38371 , n2545 );
    and g7186 ( n35629 , n29166 , n28640 );
    and g7187 ( n23742 , n4003 , n33627 );
    or g7188 ( n40161 , n24026 , n3973 );
    or g7189 ( n8463 , n2856 , n29791 );
    or g7190 ( n39667 , n27951 , n39199 );
    not g7191 ( n19385 , n25370 );
    and g7192 ( n39505 , n5787 , n9193 );
    and g7193 ( n8500 , n10026 , n34043 );
    not g7194 ( n25302 , n13032 );
    and g7195 ( n15784 , n28910 , n24087 );
    xnor g7196 ( n21649 , n20487 , n24238 );
    and g7197 ( n27047 , n32490 , n35919 );
    nor g7198 ( n4998 , n32928 , n28992 );
    not g7199 ( n1174 , n26607 );
    or g7200 ( n2699 , n19473 , n23703 );
    and g7201 ( n21076 , n10036 , n40749 );
    not g7202 ( n12722 , n41153 );
    xnor g7203 ( n5442 , n29347 , n29772 );
    and g7204 ( n25647 , n4031 , n19681 );
    xnor g7205 ( n1088 , n455 , n8372 );
    xnor g7206 ( n9585 , n25849 , n34448 );
    or g7207 ( n11493 , n27414 , n32310 );
    or g7208 ( n41296 , n40598 , n21703 );
    or g7209 ( n39769 , n17952 , n2597 );
    and g7210 ( n36506 , n19176 , n18248 );
    or g7211 ( n21824 , n19727 , n34198 );
    not g7212 ( n23201 , n31433 );
    or g7213 ( n6049 , n15604 , n41975 );
    and g7214 ( n5357 , n8436 , n17217 );
    nor g7215 ( n41322 , n14652 , n39513 );
    nor g7216 ( n21829 , n30237 , n39786 );
    and g7217 ( n13383 , n33096 , n24753 );
    not g7218 ( n19958 , n33741 );
    or g7219 ( n18418 , n27106 , n24785 );
    xnor g7220 ( n9990 , n42064 , n38297 );
    or g7221 ( n11967 , n19969 , n33762 );
    and g7222 ( n19858 , n10112 , n37351 );
    and g7223 ( n21894 , n22027 , n13351 );
    and g7224 ( n8874 , n39613 , n31962 );
    or g7225 ( n31126 , n30360 , n1322 );
    and g7226 ( n4382 , n8638 , n26064 );
    not g7227 ( n10952 , n28816 );
    and g7228 ( n40955 , n10209 , n25065 );
    or g7229 ( n25260 , n21948 , n25225 );
    and g7230 ( n13718 , n38598 , n30762 );
    not g7231 ( n16088 , n23401 );
    or g7232 ( n33839 , n13838 , n10781 );
    not g7233 ( n18558 , n40173 );
    or g7234 ( n14323 , n9584 , n9962 );
    or g7235 ( n28942 , n31652 , n17104 );
    not g7236 ( n6573 , n16987 );
    or g7237 ( n27199 , n4492 , n3083 );
    not g7238 ( n7815 , n4202 );
    nor g7239 ( n11921 , n37005 , n27465 );
    xnor g7240 ( n35150 , n17561 , n16362 );
    or g7241 ( n1176 , n5341 , n16267 );
    or g7242 ( n40220 , n25072 , n32787 );
    or g7243 ( n23680 , n33815 , n41456 );
    or g7244 ( n7063 , n6632 , n24868 );
    or g7245 ( n12294 , n14732 , n3259 );
    nor g7246 ( n8954 , n24625 , n20375 );
    and g7247 ( n27264 , n31375 , n18772 );
    xnor g7248 ( n27754 , n35727 , n18542 );
    not g7249 ( n19099 , n18469 );
    or g7250 ( n25765 , n12981 , n14441 );
    nor g7251 ( n35735 , n12570 , n10361 );
    not g7252 ( n3420 , n7702 );
    nor g7253 ( n10042 , n993 , n10840 );
    not g7254 ( n13495 , n14219 );
    and g7255 ( n16553 , n37915 , n30686 );
    xnor g7256 ( n5767 , n32178 , n20654 );
    xnor g7257 ( n32023 , n25884 , n39342 );
    not g7258 ( n11759 , n2355 );
    and g7259 ( n18742 , n8910 , n8771 );
    nor g7260 ( n23788 , n14707 , n17297 );
    not g7261 ( n22074 , n22980 );
    nor g7262 ( n18823 , n33331 , n883 );
    and g7263 ( n2280 , n21638 , n18598 );
    or g7264 ( n15018 , n36553 , n24457 );
    nor g7265 ( n42055 , n34565 , n20018 );
    and g7266 ( n14524 , n10453 , n5566 );
    and g7267 ( n13568 , n26802 , n36664 );
    or g7268 ( n41656 , n3622 , n19540 );
    or g7269 ( n20793 , n16887 , n28994 );
    and g7270 ( n17506 , n38649 , n41470 );
    not g7271 ( n41738 , n9706 );
    and g7272 ( n11970 , n21099 , n10262 );
    and g7273 ( n27538 , n26796 , n24236 );
    or g7274 ( n35605 , n42269 , n32255 );
    not g7275 ( n26443 , n7502 );
    and g7276 ( n40705 , n51 , n18818 );
    or g7277 ( n34619 , n40389 , n10861 );
    and g7278 ( n7786 , n18408 , n6670 );
    nor g7279 ( n23297 , n36094 , n11641 );
    xnor g7280 ( n36332 , n28891 , n15769 );
    not g7281 ( n20469 , n32201 );
    xnor g7282 ( n24401 , n16885 , n36842 );
    nor g7283 ( n21839 , n37419 , n11576 );
    or g7284 ( n22362 , n8653 , n17888 );
    xnor g7285 ( n29674 , n27250 , n36573 );
    or g7286 ( n21518 , n41942 , n36909 );
    and g7287 ( n9382 , n40452 , n38055 );
    or g7288 ( n41508 , n4709 , n38403 );
    and g7289 ( n33241 , n24139 , n3250 );
    and g7290 ( n26000 , n32925 , n10805 );
    or g7291 ( n14 , n9574 , n11178 );
    not g7292 ( n31016 , n2709 );
    and g7293 ( n26258 , n41486 , n32254 );
    or g7294 ( n6040 , n1944 , n4270 );
    not g7295 ( n996 , n19168 );
    xnor g7296 ( n30651 , n34358 , n36082 );
    not g7297 ( n1911 , n27623 );
    or g7298 ( n23447 , n5419 , n35091 );
    not g7299 ( n20737 , n19119 );
    or g7300 ( n29079 , n42777 , n1202 );
    and g7301 ( n14047 , n41367 , n25473 );
    nor g7302 ( n3748 , n28053 , n25531 );
    or g7303 ( n22856 , n38011 , n31851 );
    xnor g7304 ( n5695 , n29563 , n17787 );
    not g7305 ( n36137 , n20714 );
    or g7306 ( n28670 , n37720 , n36481 );
    nor g7307 ( n20484 , n23941 , n14680 );
    or g7308 ( n38457 , n21300 , n22620 );
    or g7309 ( n32035 , n35386 , n12594 );
    and g7310 ( n22164 , n24520 , n42208 );
    or g7311 ( n29333 , n41216 , n9508 );
    or g7312 ( n20922 , n17586 , n9434 );
    and g7313 ( n32276 , n26691 , n29756 );
    xnor g7314 ( n14627 , n38749 , n20283 );
    not g7315 ( n35526 , n35936 );
    not g7316 ( n4790 , n31128 );
    and g7317 ( n1024 , n9156 , n20052 );
    xnor g7318 ( n28983 , n542 , n16007 );
    nor g7319 ( n20330 , n32226 , n11844 );
    or g7320 ( n14781 , n23204 , n36313 );
    or g7321 ( n18724 , n33134 , n1334 );
    not g7322 ( n4105 , n23381 );
    or g7323 ( n37003 , n10177 , n3863 );
    and g7324 ( n5653 , n13973 , n32122 );
    and g7325 ( n7490 , n2365 , n28121 );
    or g7326 ( n21911 , n25039 , n40705 );
    nor g7327 ( n29318 , n8406 , n18551 );
    and g7328 ( n15695 , n28605 , n32235 );
    or g7329 ( n38746 , n28154 , n40352 );
    not g7330 ( n16285 , n28269 );
    nor g7331 ( n14934 , n41480 , n9308 );
    not g7332 ( n13486 , n12418 );
    and g7333 ( n36851 , n18430 , n5376 );
    xnor g7334 ( n19219 , n8873 , n4701 );
    or g7335 ( n13557 , n972 , n12242 );
    or g7336 ( n21841 , n20138 , n41685 );
    and g7337 ( n28743 , n11436 , n24 );
    nor g7338 ( n22544 , n8494 , n9212 );
    or g7339 ( n35173 , n34881 , n21770 );
    and g7340 ( n40347 , n20902 , n24360 );
    or g7341 ( n12123 , n37250 , n25674 );
    or g7342 ( n7536 , n14471 , n23751 );
    xnor g7343 ( n25836 , n20239 , n33981 );
    xnor g7344 ( n15324 , n105 , n21375 );
    not g7345 ( n15116 , n40197 );
    or g7346 ( n39845 , n29305 , n34084 );
    or g7347 ( n4975 , n35301 , n18490 );
    not g7348 ( n21948 , n14121 );
    nor g7349 ( n1293 , n32603 , n19617 );
    and g7350 ( n16614 , n40404 , n34155 );
    nor g7351 ( n35218 , n2059 , n33519 );
    not g7352 ( n25325 , n17130 );
    or g7353 ( n1515 , n4007 , n3261 );
    and g7354 ( n30600 , n13304 , n10911 );
    and g7355 ( n40563 , n13378 , n14203 );
    or g7356 ( n32610 , n7410 , n19676 );
    and g7357 ( n18308 , n31394 , n36208 );
    or g7358 ( n6814 , n37512 , n5390 );
    or g7359 ( n41161 , n25547 , n30875 );
    and g7360 ( n8146 , n34370 , n33177 );
    or g7361 ( n31304 , n2457 , n30998 );
    and g7362 ( n39112 , n3471 , n36497 );
    or g7363 ( n18 , n37863 , n39389 );
    and g7364 ( n9176 , n41568 , n21271 );
    or g7365 ( n18359 , n5906 , n11412 );
    or g7366 ( n22908 , n34907 , n39837 );
    not g7367 ( n30434 , n9596 );
    or g7368 ( n36065 , n11261 , n32353 );
    nor g7369 ( n7792 , n23139 , n38570 );
    or g7370 ( n37574 , n36344 , n940 );
    or g7371 ( n332 , n37827 , n6279 );
    not g7372 ( n34373 , n38263 );
    or g7373 ( n15810 , n20446 , n38876 );
    or g7374 ( n21411 , n10090 , n8796 );
    not g7375 ( n34652 , n31294 );
    nor g7376 ( n42804 , n20323 , n34215 );
    or g7377 ( n33578 , n34565 , n24308 );
    not g7378 ( n14945 , n4886 );
    or g7379 ( n37421 , n13160 , n5472 );
    or g7380 ( n6332 , n10119 , n32446 );
    and g7381 ( n5083 , n33303 , n28106 );
    not g7382 ( n40886 , n42550 );
    or g7383 ( n7325 , n35377 , n27130 );
    nor g7384 ( n34893 , n4906 , n23418 );
    or g7385 ( n11307 , n36071 , n4865 );
    or g7386 ( n12889 , n36393 , n11190 );
    or g7387 ( n17029 , n38867 , n31497 );
    or g7388 ( n21567 , n28721 , n41487 );
    and g7389 ( n13629 , n20829 , n28536 );
    or g7390 ( n3111 , n13830 , n34217 );
    or g7391 ( n27309 , n38191 , n37972 );
    and g7392 ( n5828 , n12155 , n20104 );
    or g7393 ( n4440 , n17114 , n1409 );
    not g7394 ( n5105 , n30081 );
    nor g7395 ( n24467 , n8186 , n40308 );
    or g7396 ( n20046 , n31015 , n5049 );
    nor g7397 ( n35978 , n33981 , n42084 );
    xnor g7398 ( n40525 , n38679 , n35907 );
    or g7399 ( n18904 , n38547 , n3728 );
    or g7400 ( n25587 , n38211 , n31700 );
    not g7401 ( n33693 , n20641 );
    or g7402 ( n18288 , n18300 , n31271 );
    and g7403 ( n3308 , n33863 , n33247 );
    and g7404 ( n33563 , n16009 , n30303 );
    and g7405 ( n26943 , n13793 , n17799 );
    xnor g7406 ( n31916 , n34235 , n40226 );
    and g7407 ( n27452 , n23229 , n15724 );
    and g7408 ( n41386 , n31233 , n30650 );
    or g7409 ( n12589 , n42446 , n28155 );
    or g7410 ( n29283 , n31187 , n7616 );
    xnor g7411 ( n20459 , n7827 , n36117 );
    not g7412 ( n10165 , n32382 );
    nor g7413 ( n18406 , n14475 , n17321 );
    xnor g7414 ( n8456 , n5457 , n5678 );
    not g7415 ( n8676 , n38282 );
    or g7416 ( n13716 , n22038 , n14204 );
    and g7417 ( n18057 , n15228 , n1310 );
    xnor g7418 ( n18144 , n15886 , n22421 );
    not g7419 ( n14298 , n10587 );
    and g7420 ( n41460 , n5003 , n25569 );
    or g7421 ( n11020 , n30071 , n29162 );
    not g7422 ( n27594 , n7510 );
    xnor g7423 ( n4697 , n32297 , n6745 );
    and g7424 ( n13260 , n11806 , n13813 );
    nor g7425 ( n30290 , n39882 , n9463 );
    or g7426 ( n1227 , n7322 , n21509 );
    nor g7427 ( n13333 , n15123 , n33025 );
    and g7428 ( n33864 , n5103 , n13424 );
    and g7429 ( n23467 , n22477 , n42736 );
    or g7430 ( n38579 , n28080 , n42061 );
    nor g7431 ( n7149 , n27745 , n30232 );
    not g7432 ( n37883 , n7656 );
    or g7433 ( n18989 , n37587 , n15335 );
    or g7434 ( n5516 , n41752 , n37401 );
    and g7435 ( n13380 , n17672 , n36013 );
    or g7436 ( n744 , n4391 , n26046 );
    or g7437 ( n18768 , n24626 , n30008 );
    or g7438 ( n15697 , n19558 , n36848 );
    not g7439 ( n10213 , n24726 );
    xnor g7440 ( n12493 , n29571 , n1971 );
    and g7441 ( n41312 , n38139 , n18936 );
    or g7442 ( n23306 , n16736 , n38465 );
    or g7443 ( n22198 , n26144 , n15882 );
    nor g7444 ( n2025 , n10929 , n20666 );
    and g7445 ( n17061 , n29966 , n26732 );
    nor g7446 ( n23695 , n2214 , n3525 );
    or g7447 ( n2636 , n1122 , n904 );
    not g7448 ( n35073 , n42369 );
    or g7449 ( n13627 , n8177 , n14479 );
    xnor g7450 ( n37326 , n1255 , n779 );
    nor g7451 ( n16367 , n10417 , n38846 );
    or g7452 ( n28759 , n25033 , n42751 );
    or g7453 ( n18232 , n12867 , n4987 );
    or g7454 ( n7185 , n28698 , n24229 );
    xnor g7455 ( n4760 , n38029 , n14001 );
    or g7456 ( n14940 , n15285 , n37862 );
    or g7457 ( n36780 , n5681 , n6359 );
    or g7458 ( n36592 , n11431 , n10568 );
    nor g7459 ( n10789 , n8611 , n23590 );
    or g7460 ( n34104 , n33043 , n36575 );
    or g7461 ( n29188 , n30782 , n36509 );
    or g7462 ( n18254 , n26861 , n3589 );
    not g7463 ( n37523 , n37245 );
    or g7464 ( n7137 , n614 , n30482 );
    xnor g7465 ( n1169 , n28916 , n10920 );
    or g7466 ( n19046 , n33870 , n40610 );
    and g7467 ( n2576 , n1209 , n26525 );
    or g7468 ( n34089 , n22091 , n12606 );
    xnor g7469 ( n4353 , n37543 , n15466 );
    and g7470 ( n42052 , n32546 , n11402 );
    or g7471 ( n34630 , n5168 , n34289 );
    or g7472 ( n15622 , n39719 , n24183 );
    or g7473 ( n1869 , n34648 , n23280 );
    or g7474 ( n22509 , n13639 , n32752 );
    or g7475 ( n23355 , n5720 , n6019 );
    or g7476 ( n19820 , n33433 , n37220 );
    nor g7477 ( n14957 , n3067 , n40112 );
    and g7478 ( n14899 , n1397 , n860 );
    and g7479 ( n28141 , n21705 , n9179 );
    xnor g7480 ( n20278 , n40155 , n19286 );
    and g7481 ( n32104 , n33790 , n34944 );
    nor g7482 ( n42886 , n27593 , n22464 );
    nor g7483 ( n29524 , n7613 , n14856 );
    or g7484 ( n17123 , n28205 , n6819 );
    or g7485 ( n10923 , n15867 , n29583 );
    xnor g7486 ( n33790 , n34329 , n11648 );
    and g7487 ( n41766 , n11869 , n3610 );
    xnor g7488 ( n12799 , n32507 , n19353 );
    or g7489 ( n35148 , n6628 , n37219 );
    xnor g7490 ( n20647 , n105 , n17432 );
    or g7491 ( n26676 , n29924 , n6124 );
    and g7492 ( n7079 , n9361 , n6814 );
    and g7493 ( n570 , n19226 , n36688 );
    not g7494 ( n18589 , n19010 );
    or g7495 ( n10339 , n12019 , n3740 );
    not g7496 ( n38080 , n22212 );
    and g7497 ( n29649 , n40030 , n42799 );
    or g7498 ( n25153 , n12930 , n32478 );
    and g7499 ( n22373 , n42029 , n1052 );
    nor g7500 ( n25812 , n30864 , n22448 );
    not g7501 ( n23285 , n5819 );
    or g7502 ( n41418 , n12008 , n40032 );
    and g7503 ( n30620 , n23840 , n30827 );
    or g7504 ( n11094 , n10511 , n32002 );
    or g7505 ( n8826 , n39318 , n27738 );
    or g7506 ( n18613 , n33998 , n22278 );
    xnor g7507 ( n22742 , n17267 , n35124 );
    nor g7508 ( n31418 , n11380 , n41833 );
    or g7509 ( n5076 , n39489 , n17569 );
    xnor g7510 ( n3704 , n40 , n31315 );
    or g7511 ( n37795 , n20486 , n18321 );
    or g7512 ( n40858 , n8976 , n440 );
    or g7513 ( n2447 , n10610 , n3988 );
    and g7514 ( n9536 , n29819 , n9237 );
    nor g7515 ( n38558 , n1722 , n849 );
    xnor g7516 ( n14922 , n29646 , n23530 );
    not g7517 ( n34419 , n21503 );
    not g7518 ( n41358 , n3334 );
    nor g7519 ( n11678 , n13921 , n12575 );
    or g7520 ( n397 , n15282 , n16441 );
    and g7521 ( n32525 , n4878 , n35786 );
    or g7522 ( n33975 , n37783 , n42300 );
    or g7523 ( n17298 , n5964 , n37303 );
    and g7524 ( n37675 , n11499 , n10144 );
    or g7525 ( n27649 , n28337 , n27179 );
    nor g7526 ( n26553 , n4879 , n2153 );
    or g7527 ( n25385 , n16920 , n37689 );
    and g7528 ( n2380 , n3 , n31942 );
    or g7529 ( n30056 , n16744 , n22991 );
    or g7530 ( n24004 , n35450 , n9851 );
    xnor g7531 ( n30136 , n30833 , n6133 );
    or g7532 ( n33389 , n20978 , n13854 );
    and g7533 ( n23826 , n4857 , n5596 );
    or g7534 ( n42897 , n3773 , n5984 );
    not g7535 ( n16094 , n4468 );
    or g7536 ( n1343 , n7219 , n37804 );
    and g7537 ( n18534 , n32084 , n25609 );
    xnor g7538 ( n13032 , n39705 , n1380 );
    and g7539 ( n22859 , n25253 , n13660 );
    xnor g7540 ( n37216 , n8602 , n17193 );
    or g7541 ( n26222 , n27070 , n33929 );
    and g7542 ( n24012 , n38253 , n28287 );
    nor g7543 ( n16588 , n1683 , n16359 );
    and g7544 ( n8828 , n32648 , n5948 );
    and g7545 ( n33547 , n10187 , n27 );
    and g7546 ( n3066 , n7886 , n34443 );
    not g7547 ( n12279 , n12342 );
    or g7548 ( n38968 , n14677 , n19497 );
    or g7549 ( n28637 , n37099 , n14137 );
    or g7550 ( n23222 , n34554 , n32367 );
    not g7551 ( n39036 , n40168 );
    not g7552 ( n35732 , n8465 );
    and g7553 ( n20025 , n36053 , n18160 );
    and g7554 ( n35332 , n42279 , n25825 );
    and g7555 ( n17065 , n42426 , n11965 );
    not g7556 ( n14996 , n2769 );
    nor g7557 ( n33649 , n14148 , n6747 );
    nor g7558 ( n9860 , n3608 , n27391 );
    not g7559 ( n36114 , n20076 );
    xnor g7560 ( n10294 , n22054 , n38622 );
    and g7561 ( n2440 , n8609 , n23443 );
    or g7562 ( n31816 , n41356 , n25445 );
    or g7563 ( n19426 , n7178 , n12484 );
    or g7564 ( n1021 , n39991 , n16083 );
    not g7565 ( n23947 , n246 );
    nor g7566 ( n1769 , n10971 , n6069 );
    not g7567 ( n12156 , n24498 );
    xnor g7568 ( n32016 , n21973 , n38067 );
    xnor g7569 ( n8206 , n4651 , n16597 );
    nor g7570 ( n25829 , n8494 , n16354 );
    or g7571 ( n38858 , n6503 , n2762 );
    not g7572 ( n27879 , n3695 );
    xnor g7573 ( n26131 , n11109 , n13709 );
    or g7574 ( n4135 , n32731 , n8284 );
    nor g7575 ( n36037 , n22408 , n25138 );
    nor g7576 ( n42630 , n36636 , n22024 );
    xnor g7577 ( n20154 , n27246 , n19221 );
    and g7578 ( n4922 , n28300 , n31842 );
    or g7579 ( n15249 , n33951 , n22502 );
    nor g7580 ( n24261 , n19586 , n29248 );
    and g7581 ( n26078 , n25619 , n17085 );
    or g7582 ( n15378 , n22281 , n42311 );
    or g7583 ( n28738 , n22440 , n14126 );
    or g7584 ( n17365 , n5408 , n27146 );
    nor g7585 ( n16541 , n40698 , n17721 );
    nor g7586 ( n1619 , n25237 , n8217 );
    and g7587 ( n26494 , n15558 , n3509 );
    nor g7588 ( n9039 , n19262 , n25500 );
    xnor g7589 ( n23746 , n20487 , n6436 );
    or g7590 ( n41599 , n15424 , n24718 );
    nor g7591 ( n6199 , n22461 , n21626 );
    or g7592 ( n8606 , n11443 , n4625 );
    xnor g7593 ( n16113 , n18303 , n35202 );
    nor g7594 ( n36852 , n5897 , n127 );
    and g7595 ( n28164 , n31425 , n4152 );
    not g7596 ( n33397 , n35966 );
    xnor g7597 ( n30242 , n17436 , n26177 );
    not g7598 ( n39640 , n28362 );
    not g7599 ( n15917 , n8652 );
    or g7600 ( n15104 , n6664 , n8483 );
    not g7601 ( n36461 , n20873 );
    or g7602 ( n23175 , n12130 , n20985 );
    nor g7603 ( n18326 , n3817 , n21814 );
    not g7604 ( n42118 , n19952 );
    not g7605 ( n21019 , n19571 );
    or g7606 ( n7098 , n3459 , n26207 );
    or g7607 ( n8896 , n28887 , n1924 );
    not g7608 ( n36203 , n32637 );
    and g7609 ( n12215 , n36595 , n23668 );
    nor g7610 ( n3346 , n38879 , n4171 );
    not g7611 ( n18390 , n36665 );
    or g7612 ( n36060 , n17232 , n8132 );
    not g7613 ( n30561 , n22848 );
    not g7614 ( n33730 , n34042 );
    nor g7615 ( n33562 , n42760 , n42301 );
    or g7616 ( n4414 , n24050 , n16410 );
    xnor g7617 ( n14828 , n24505 , n12243 );
    and g7618 ( n15895 , n29535 , n34346 );
    xnor g7619 ( n10825 , n18874 , n40082 );
    and g7620 ( n17891 , n11841 , n16000 );
    or g7621 ( n32935 , n24736 , n27127 );
    or g7622 ( n21257 , n31343 , n27725 );
    not g7623 ( n11132 , n35983 );
    or g7624 ( n4685 , n3684 , n33297 );
    or g7625 ( n1606 , n28643 , n8213 );
    and g7626 ( n25614 , n38294 , n747 );
    nor g7627 ( n17008 , n31698 , n35007 );
    or g7628 ( n40715 , n19135 , n28038 );
    nor g7629 ( n38170 , n12328 , n25199 );
    xnor g7630 ( n35983 , n34226 , n1279 );
    xnor g7631 ( n19231 , n37309 , n29510 );
    and g7632 ( n21103 , n14151 , n24936 );
    or g7633 ( n23244 , n15185 , n16089 );
    or g7634 ( n9846 , n8180 , n20078 );
    or g7635 ( n25842 , n473 , n41772 );
    or g7636 ( n30385 , n6423 , n38297 );
    or g7637 ( n31576 , n23691 , n17383 );
    not g7638 ( n22824 , n40063 );
    or g7639 ( n39403 , n30123 , n33770 );
    or g7640 ( n26415 , n33135 , n3937 );
    xnor g7641 ( n28226 , n27421 , n24981 );
    and g7642 ( n34481 , n1542 , n33613 );
    or g7643 ( n29789 , n36117 , n15070 );
    or g7644 ( n20959 , n21524 , n10667 );
    or g7645 ( n27170 , n1817 , n20446 );
    or g7646 ( n27587 , n25407 , n26578 );
    xnor g7647 ( n33654 , n37175 , n1226 );
    nor g7648 ( n15734 , n18757 , n35857 );
    or g7649 ( n14203 , n10544 , n39328 );
    or g7650 ( n33564 , n29027 , n13852 );
    or g7651 ( n13988 , n37836 , n20923 );
    or g7652 ( n23219 , n33049 , n41829 );
    or g7653 ( n4769 , n32041 , n30702 );
    or g7654 ( n41272 , n41773 , n6241 );
    or g7655 ( n35556 , n2830 , n33464 );
    or g7656 ( n6768 , n8076 , n22704 );
    xnor g7657 ( n7239 , n9237 , n29819 );
    or g7658 ( n35436 , n18344 , n40323 );
    nor g7659 ( n29080 , n8540 , n2006 );
    not g7660 ( n27398 , n24498 );
    or g7661 ( n1366 , n19221 , n14899 );
    or g7662 ( n30649 , n5964 , n11639 );
    or g7663 ( n16378 , n42109 , n27127 );
    and g7664 ( n4654 , n37525 , n19650 );
    or g7665 ( n5736 , n38557 , n3854 );
    or g7666 ( n40291 , n23745 , n36373 );
    xnor g7667 ( n32146 , n26609 , n18712 );
    nor g7668 ( n7204 , n9001 , n41857 );
    or g7669 ( n28966 , n21032 , n22614 );
    or g7670 ( n9431 , n28887 , n24288 );
    or g7671 ( n7002 , n20328 , n15342 );
    or g7672 ( n27007 , n11976 , n6183 );
    not g7673 ( n25193 , n24372 );
    not g7674 ( n19159 , n13668 );
    or g7675 ( n1998 , n38463 , n36536 );
    and g7676 ( n16903 , n7344 , n20008 );
    and g7677 ( n26585 , n10838 , n42503 );
    not g7678 ( n7943 , n34922 );
    or g7679 ( n23208 , n40253 , n18492 );
    and g7680 ( n6679 , n6656 , n22338 );
    xnor g7681 ( n40559 , n10394 , n18108 );
    or g7682 ( n18245 , n1211 , n42706 );
    not g7683 ( n40695 , n20736 );
    and g7684 ( n2303 , n25503 , n41503 );
    or g7685 ( n31479 , n36163 , n7170 );
    nor g7686 ( n36967 , n1448 , n25329 );
    not g7687 ( n8662 , n10052 );
    xnor g7688 ( n28840 , n784 , n12629 );
    nor g7689 ( n42525 , n14707 , n12931 );
    nor g7690 ( n6388 , n21759 , n8508 );
    and g7691 ( n26841 , n29014 , n31667 );
    not g7692 ( n26512 , n41391 );
    not g7693 ( n19611 , n41427 );
    or g7694 ( n40348 , n23862 , n31475 );
    and g7695 ( n3235 , n36879 , n1103 );
    or g7696 ( n7917 , n13223 , n5124 );
    nor g7697 ( n1378 , n25588 , n16768 );
    or g7698 ( n35561 , n30899 , n13751 );
    or g7699 ( n23729 , n21639 , n1631 );
    or g7700 ( n15991 , n34114 , n1527 );
    xnor g7701 ( n29845 , n105 , n7682 );
    and g7702 ( n4270 , n13845 , n6298 );
    or g7703 ( n4315 , n36727 , n35284 );
    not g7704 ( n8930 , n37749 );
    or g7705 ( n40344 , n12072 , n11374 );
    or g7706 ( n28910 , n2818 , n39680 );
    xnor g7707 ( n762 , n21888 , n29738 );
    or g7708 ( n22135 , n32269 , n7289 );
    or g7709 ( n28008 , n28891 , n15769 );
    nor g7710 ( n13961 , n30862 , n25945 );
    not g7711 ( n25642 , n18915 );
    or g7712 ( n40021 , n38808 , n16575 );
    and g7713 ( n32235 , n160 , n31028 );
    not g7714 ( n25893 , n27463 );
    nor g7715 ( n38552 , n14188 , n8951 );
    or g7716 ( n22107 , n39266 , n22564 );
    or g7717 ( n33515 , n33556 , n7793 );
    xnor g7718 ( n12339 , n18530 , n31776 );
    or g7719 ( n37089 , n14471 , n26897 );
    or g7720 ( n15533 , n16350 , n42810 );
    not g7721 ( n18298 , n24526 );
    nor g7722 ( n34013 , n13474 , n673 );
    or g7723 ( n31042 , n33931 , n17978 );
    or g7724 ( n40750 , n7802 , n7159 );
    nor g7725 ( n23051 , n34565 , n38483 );
    or g7726 ( n36984 , n1039 , n24307 );
    and g7727 ( n33481 , n33631 , n2491 );
    xnor g7728 ( n14876 , n1622 , n23300 );
    not g7729 ( n22440 , n35966 );
    nor g7730 ( n19870 , n29053 , n33350 );
    or g7731 ( n24270 , n31542 , n22876 );
    or g7732 ( n40706 , n18534 , n33984 );
    or g7733 ( n2150 , n35732 , n13421 );
    and g7734 ( n35160 , n21980 , n3349 );
    and g7735 ( n17720 , n15414 , n9545 );
    or g7736 ( n37135 , n39922 , n19842 );
    and g7737 ( n11190 , n21529 , n35902 );
    or g7738 ( n18555 , n14941 , n38127 );
    not g7739 ( n5205 , n38802 );
    or g7740 ( n28019 , n22709 , n23085 );
    or g7741 ( n12102 , n26601 , n41923 );
    nor g7742 ( n7793 , n36074 , n12534 );
    and g7743 ( n944 , n25856 , n13943 );
    not g7744 ( n9035 , n36154 );
    or g7745 ( n12230 , n4899 , n33175 );
    not g7746 ( n11072 , n31015 );
    nor g7747 ( n42912 , n22967 , n10296 );
    not g7748 ( n20115 , n369 );
    or g7749 ( n20836 , n37805 , n6326 );
    xnor g7750 ( n42671 , n10352 , n11623 );
    or g7751 ( n24329 , n25136 , n31019 );
    not g7752 ( n18990 , n14870 );
    not g7753 ( n40512 , n25325 );
    and g7754 ( n17759 , n5301 , n41977 );
    or g7755 ( n26011 , n21894 , n27949 );
    or g7756 ( n20827 , n23694 , n42582 );
    xnor g7757 ( n25283 , n898 , n21782 );
    or g7758 ( n36635 , n5110 , n1127 );
    xnor g7759 ( n32234 , n24546 , n29488 );
    or g7760 ( n28131 , n15157 , n39619 );
    xnor g7761 ( n23439 , n41013 , n20004 );
    or g7762 ( n12940 , n24439 , n34665 );
    or g7763 ( n27283 , n23902 , n19446 );
    not g7764 ( n17492 , n42848 );
    not g7765 ( n42501 , n27395 );
    or g7766 ( n35666 , n28486 , n14819 );
    and g7767 ( n23670 , n31331 , n37568 );
    and g7768 ( n29627 , n5297 , n12720 );
    not g7769 ( n2348 , n6642 );
    or g7770 ( n31062 , n240 , n12343 );
    and g7771 ( n2085 , n31290 , n23568 );
    or g7772 ( n17986 , n17851 , n23290 );
    or g7773 ( n38171 , n4842 , n12683 );
    and g7774 ( n31012 , n4804 , n4126 );
    not g7775 ( n2005 , n8663 );
    nor g7776 ( n32514 , n4796 , n7768 );
    or g7777 ( n33075 , n18447 , n33464 );
    not g7778 ( n13753 , n26871 );
    and g7779 ( n2470 , n22497 , n3523 );
    or g7780 ( n42216 , n8626 , n42180 );
    and g7781 ( n268 , n14471 , n41727 );
    and g7782 ( n39851 , n20584 , n21455 );
    nor g7783 ( n41573 , n1457 , n22761 );
    xnor g7784 ( n25380 , n22103 , n34095 );
    nor g7785 ( n9562 , n1002 , n41653 );
    not g7786 ( n13506 , n34021 );
    or g7787 ( n35784 , n31077 , n2119 );
    and g7788 ( n28115 , n4971 , n11026 );
    nor g7789 ( n33802 , n38157 , n42052 );
    or g7790 ( n37048 , n11947 , n1021 );
    xnor g7791 ( n3065 , n27968 , n4323 );
    or g7792 ( n7736 , n20484 , n13525 );
    not g7793 ( n32912 , n24444 );
    or g7794 ( n32567 , n18480 , n10437 );
    or g7795 ( n32687 , n34873 , n33691 );
    nor g7796 ( n22755 , n36625 , n35907 );
    or g7797 ( n6225 , n24660 , n12939 );
    or g7798 ( n35299 , n39118 , n1024 );
    or g7799 ( n16175 , n5264 , n13938 );
    and g7800 ( n1173 , n37422 , n13035 );
    and g7801 ( n3408 , n12900 , n9570 );
    or g7802 ( n24630 , n3347 , n9804 );
    and g7803 ( n14898 , n4918 , n28137 );
    nor g7804 ( n34775 , n27762 , n26710 );
    and g7805 ( n6704 , n11436 , n35082 );
    or g7806 ( n4811 , n35564 , n30334 );
    and g7807 ( n10244 , n4057 , n36026 );
    not g7808 ( n9492 , n570 );
    or g7809 ( n36341 , n41571 , n6094 );
    not g7810 ( n33626 , n24531 );
    not g7811 ( n26235 , n40058 );
    or g7812 ( n9235 , n22538 , n929 );
    and g7813 ( n35489 , n22586 , n37463 );
    or g7814 ( n34255 , n36949 , n29545 );
    and g7815 ( n10108 , n9600 , n28951 );
    or g7816 ( n15171 , n28651 , n11374 );
    or g7817 ( n21764 , n18196 , n26087 );
    xnor g7818 ( n39442 , n9412 , n37699 );
    nor g7819 ( n37323 , n5356 , n20171 );
    or g7820 ( n5542 , n37730 , n16465 );
    and g7821 ( n30400 , n30497 , n14453 );
    not g7822 ( n22054 , n14870 );
    or g7823 ( n7808 , n32722 , n25249 );
    and g7824 ( n42814 , n36009 , n18830 );
    not g7825 ( n33755 , n341 );
    nor g7826 ( n2750 , n39266 , n36485 );
    xnor g7827 ( n22139 , n41947 , n32975 );
    and g7828 ( n40984 , n6580 , n24756 );
    nor g7829 ( n10468 , n29577 , n15331 );
    and g7830 ( n18213 , n16183 , n4058 );
    and g7831 ( n13930 , n41711 , n22717 );
    or g7832 ( n15755 , n32986 , n30586 );
    nor g7833 ( n28009 , n16885 , n28598 );
    and g7834 ( n17303 , n9154 , n10865 );
    xnor g7835 ( n10721 , n9460 , n19445 );
    and g7836 ( n36389 , n39086 , n34471 );
    or g7837 ( n4871 , n37520 , n25273 );
    nor g7838 ( n15965 , n7987 , n40437 );
    nor g7839 ( n25169 , n28593 , n38678 );
    or g7840 ( n11396 , n39367 , n36771 );
    not g7841 ( n7993 , n41223 );
    not g7842 ( n10822 , n34500 );
    nor g7843 ( n39047 , n34566 , n10529 );
    nor g7844 ( n27316 , n1278 , n27368 );
    and g7845 ( n13400 , n42573 , n34946 );
    not g7846 ( n965 , n31764 );
    or g7847 ( n3188 , n15523 , n12129 );
    and g7848 ( n35333 , n22331 , n13452 );
    nor g7849 ( n33088 , n13336 , n28607 );
    or g7850 ( n32461 , n9319 , n11787 );
    xnor g7851 ( n31432 , n15106 , n8494 );
    or g7852 ( n24842 , n14134 , n20570 );
    or g7853 ( n11019 , n17310 , n19402 );
    xnor g7854 ( n33505 , n35727 , n7854 );
    or g7855 ( n42716 , n12188 , n26338 );
    nor g7856 ( n38320 , n14990 , n18164 );
    or g7857 ( n9816 , n7498 , n29884 );
    or g7858 ( n1536 , n39991 , n385 );
    and g7859 ( n3120 , n12893 , n17534 );
    and g7860 ( n40483 , n5964 , n2176 );
    and g7861 ( n35111 , n40513 , n32613 );
    or g7862 ( n11263 , n4535 , n37182 );
    or g7863 ( n36329 , n1444 , n42095 );
    and g7864 ( n14695 , n10338 , n37178 );
    not g7865 ( n8735 , n21764 );
    xnor g7866 ( n5721 , n39051 , n3913 );
    nor g7867 ( n6120 , n14265 , n38427 );
    xnor g7868 ( n22537 , n29740 , n39171 );
    xnor g7869 ( n32813 , n10414 , n18964 );
    or g7870 ( n16781 , n40604 , n21117 );
    or g7871 ( n4528 , n8356 , n697 );
    not g7872 ( n42725 , n41427 );
    or g7873 ( n4269 , n425 , n17394 );
    or g7874 ( n20627 , n11976 , n19839 );
    or g7875 ( n9966 , n23774 , n30071 );
    or g7876 ( n2027 , n20296 , n31211 );
    or g7877 ( n15694 , n28551 , n20460 );
    or g7878 ( n42000 , n22419 , n18938 );
    or g7879 ( n16130 , n7356 , n17503 );
    not g7880 ( n17049 , n22777 );
    and g7881 ( n4290 , n37330 , n15381 );
    nor g7882 ( n23283 , n15388 , n19010 );
    and g7883 ( n34588 , n17093 , n29442 );
    not g7884 ( n38662 , n34880 );
    nor g7885 ( n23862 , n30641 , n8424 );
    and g7886 ( n14561 , n5749 , n10931 );
    or g7887 ( n37529 , n524 , n30453 );
    not g7888 ( n36667 , n26749 );
    or g7889 ( n23913 , n2599 , n4171 );
    or g7890 ( n10237 , n37144 , n4128 );
    not g7891 ( n26334 , n28655 );
    xnor g7892 ( n14652 , n13444 , n19404 );
    and g7893 ( n21014 , n35844 , n10899 );
    not g7894 ( n37120 , n27925 );
    or g7895 ( n26438 , n30872 , n40702 );
    or g7896 ( n26169 , n35879 , n6126 );
    and g7897 ( n310 , n40469 , n10319 );
    nor g7898 ( n2260 , n27767 , n21084 );
    not g7899 ( n7659 , n36256 );
    or g7900 ( n30469 , n14929 , n19887 );
    xnor g7901 ( n958 , n38497 , n41659 );
    and g7902 ( n36103 , n32031 , n10236 );
    nor g7903 ( n8983 , n2896 , n32698 );
    nor g7904 ( n21420 , n16870 , n22811 );
    not g7905 ( n17942 , n24945 );
    and g7906 ( n27424 , n36974 , n19290 );
    xnor g7907 ( n36120 , n28079 , n38879 );
    and g7908 ( n33752 , n1573 , n36123 );
    not g7909 ( n35268 , n4981 );
    nor g7910 ( n24262 , n17744 , n9609 );
    and g7911 ( n16441 , n32776 , n12229 );
    nor g7912 ( n42381 , n36486 , n17045 );
    or g7913 ( n6184 , n16161 , n4374 );
    or g7914 ( n5773 , n38999 , n16999 );
    not g7915 ( n16649 , n42803 );
    not g7916 ( n29396 , n39248 );
    xnor g7917 ( n33493 , n36998 , n3155 );
    xnor g7918 ( n36484 , n4334 , n37791 );
    or g7919 ( n26434 , n1584 , n33401 );
    or g7920 ( n42297 , n31636 , n2910 );
    or g7921 ( n7135 , n29219 , n36713 );
    and g7922 ( n15248 , n24207 , n5617 );
    and g7923 ( n1318 , n8191 , n7312 );
    and g7924 ( n37862 , n5000 , n39220 );
    xnor g7925 ( n19281 , n42572 , n36103 );
    not g7926 ( n4517 , n31075 );
    or g7927 ( n17501 , n2801 , n28642 );
    or g7928 ( n23991 , n35269 , n16181 );
    or g7929 ( n26673 , n33892 , n32244 );
    nor g7930 ( n30967 , n24129 , n4142 );
    or g7931 ( n30474 , n8494 , n15278 );
    or g7932 ( n37568 , n30984 , n8990 );
    or g7933 ( n38439 , n38066 , n42670 );
    or g7934 ( n40076 , n8195 , n17777 );
    nor g7935 ( n20587 , n13832 , n8180 );
    nor g7936 ( n25427 , n12593 , n2250 );
    or g7937 ( n30332 , n31410 , n18242 );
    and g7938 ( n35533 , n4032 , n8176 );
    or g7939 ( n5157 , n3082 , n3543 );
    not g7940 ( n11404 , n36792 );
    or g7941 ( n1936 , n39436 , n39378 );
    or g7942 ( n8869 , n9040 , n4486 );
    xnor g7943 ( n13407 , n9486 , n15821 );
    nor g7944 ( n40313 , n13793 , n17799 );
    not g7945 ( n37880 , n30047 );
    nor g7946 ( n18097 , n31187 , n42317 );
    or g7947 ( n8815 , n32277 , n36861 );
    nor g7948 ( n4624 , n9906 , n18699 );
    and g7949 ( n4701 , n34834 , n37174 );
    or g7950 ( n19043 , n37983 , n19405 );
    and g7951 ( n19226 , n33209 , n14968 );
    xnor g7952 ( n34706 , n35154 , n9049 );
    or g7953 ( n39728 , n28883 , n17422 );
    and g7954 ( n28722 , n32888 , n15458 );
    nor g7955 ( n21408 , n11451 , n22515 );
    not g7956 ( n24072 , n32071 );
    nor g7957 ( n35674 , n1555 , n23786 );
    and g7958 ( n31765 , n20171 , n26754 );
    or g7959 ( n4000 , n8373 , n16248 );
    or g7960 ( n30249 , n904 , n6080 );
    xnor g7961 ( n18659 , n39957 , n40009 );
    and g7962 ( n42532 , n35881 , n19595 );
    or g7963 ( n34700 , n7994 , n2599 );
    or g7964 ( n12134 , n42404 , n35541 );
    nor g7965 ( n19601 , n6564 , n12401 );
    nor g7966 ( n37855 , n38760 , n39272 );
    or g7967 ( n40031 , n16911 , n28447 );
    or g7968 ( n17755 , n29454 , n30352 );
    not g7969 ( n15236 , n16246 );
    and g7970 ( n42006 , n35075 , n31835 );
    or g7971 ( n7274 , n4598 , n14053 );
    or g7972 ( n28930 , n5650 , n35540 );
    nor g7973 ( n21013 , n28801 , n39298 );
    or g7974 ( n5762 , n42333 , n42245 );
    or g7975 ( n41199 , n34604 , n37129 );
    nor g7976 ( n35283 , n12156 , n39506 );
    or g7977 ( n35052 , n31261 , n27699 );
    or g7978 ( n1710 , n20100 , n32068 );
    or g7979 ( n26008 , n42314 , n5881 );
    or g7980 ( n40925 , n33348 , n21708 );
    or g7981 ( n5572 , n33719 , n35190 );
    not g7982 ( n38676 , n42821 );
    or g7983 ( n31416 , n27762 , n3424 );
    or g7984 ( n23580 , n35443 , n4124 );
    xnor g7985 ( n28007 , n40941 , n3594 );
    or g7986 ( n2083 , n8293 , n18293 );
    or g7987 ( n25046 , n20364 , n8262 );
    or g7988 ( n41816 , n14944 , n15082 );
    not g7989 ( n4529 , n15691 );
    or g7990 ( n4754 , n6636 , n34978 );
    or g7991 ( n42194 , n27924 , n36494 );
    or g7992 ( n26517 , n21711 , n39151 );
    xnor g7993 ( n41004 , n24093 , n3548 );
    not g7994 ( n7864 , n15396 );
    or g7995 ( n9070 , n5210 , n24626 );
    and g7996 ( n7201 , n27590 , n26151 );
    or g7997 ( n10663 , n19563 , n34955 );
    xnor g7998 ( n29348 , n19665 , n23977 );
    and g7999 ( n31440 , n6778 , n20873 );
    nor g8000 ( n37606 , n526 , n35476 );
    and g8001 ( n17657 , n16110 , n7007 );
    not g8002 ( n42810 , n28089 );
    or g8003 ( n39895 , n30298 , n34201 );
    or g8004 ( n3352 , n3815 , n9800 );
    and g8005 ( n15077 , n29124 , n15664 );
    not g8006 ( n35934 , n31953 );
    not g8007 ( n8473 , n32828 );
    or g8008 ( n7698 , n14821 , n3564 );
    and g8009 ( n26479 , n20794 , n8789 );
    xnor g8010 ( n19180 , n21381 , n18101 );
    and g8011 ( n16092 , n554 , n15909 );
    or g8012 ( n14244 , n37771 , n25427 );
    not g8013 ( n30752 , n12634 );
    or g8014 ( n33499 , n11916 , n18009 );
    and g8015 ( n33152 , n12709 , n5397 );
    xnor g8016 ( n18461 , n41013 , n22020 );
    or g8017 ( n12197 , n31950 , n28148 );
    or g8018 ( n10151 , n36117 , n36587 );
    and g8019 ( n3018 , n7154 , n2321 );
    xnor g8020 ( n6892 , n19495 , n16021 );
    not g8021 ( n37787 , n23667 );
    or g8022 ( n42590 , n20094 , n21500 );
    nor g8023 ( n38059 , n20299 , n25801 );
    nor g8024 ( n29233 , n5896 , n30101 );
    not g8025 ( n39741 , n29662 );
    xnor g8026 ( n21097 , n836 , n20666 );
    or g8027 ( n35817 , n34565 , n23542 );
    or g8028 ( n31040 , n20746 , n31497 );
    nor g8029 ( n41597 , n10273 , n7895 );
    nor g8030 ( n38420 , n14981 , n2945 );
    or g8031 ( n39240 , n24745 , n441 );
    not g8032 ( n3802 , n34142 );
    or g8033 ( n38090 , n7139 , n17240 );
    or g8034 ( n1085 , n23925 , n27857 );
    xnor g8035 ( n10356 , n37896 , n24229 );
    or g8036 ( n16662 , n35292 , n5934 );
    xnor g8037 ( n31821 , n27035 , n2140 );
    or g8038 ( n1194 , n5874 , n12021 );
    nor g8039 ( n37197 , n2232 , n38786 );
    or g8040 ( n7394 , n31298 , n16575 );
    or g8041 ( n3594 , n7971 , n30785 );
    or g8042 ( n15114 , n33297 , n39490 );
    and g8043 ( n37414 , n18372 , n9535 );
    and g8044 ( n17812 , n28631 , n20195 );
    or g8045 ( n36204 , n24626 , n29982 );
    or g8046 ( n41455 , n33205 , n21175 );
    or g8047 ( n8446 , n34732 , n211 );
    and g8048 ( n30867 , n11370 , n17357 );
    nor g8049 ( n23700 , n589 , n11346 );
    and g8050 ( n42396 , n25782 , n18056 );
    and g8051 ( n11979 , n41395 , n34025 );
    nor g8052 ( n87 , n40001 , n16258 );
    and g8053 ( n19475 , n39051 , n3913 );
    or g8054 ( n39801 , n31944 , n6390 );
    xnor g8055 ( n21537 , n11255 , n14471 );
    or g8056 ( n4199 , n27902 , n4346 );
    or g8057 ( n35655 , n1581 , n33727 );
    or g8058 ( n5069 , n23445 , n14998 );
    or g8059 ( n9624 , n4119 , n35231 );
    nor g8060 ( n41598 , n30623 , n12655 );
    not g8061 ( n35471 , n8182 );
    or g8062 ( n32302 , n18481 , n31156 );
    or g8063 ( n16128 , n7020 , n31831 );
    xnor g8064 ( n6227 , n17724 , n1160 );
    or g8065 ( n36285 , n5027 , n11456 );
    and g8066 ( n15879 , n6222 , n19501 );
    or g8067 ( n13543 , n2614 , n8162 );
    or g8068 ( n13673 , n4018 , n14691 );
    not g8069 ( n26991 , n15228 );
    or g8070 ( n35065 , n315 , n4669 );
    and g8071 ( n36163 , n16991 , n7405 );
    nor g8072 ( n35529 , n34686 , n6669 );
    and g8073 ( n456 , n5226 , n4935 );
    nor g8074 ( n14093 , n236 , n40037 );
    nor g8075 ( n8865 , n4257 , n27284 );
    or g8076 ( n6834 , n26531 , n27592 );
    xnor g8077 ( n14990 , n6625 , n34670 );
    or g8078 ( n31287 , n26587 , n41963 );
    xnor g8079 ( n22556 , n32132 , n2899 );
    and g8080 ( n9713 , n23979 , n41076 );
    and g8081 ( n8155 , n548 , n6305 );
    or g8082 ( n17699 , n32711 , n33254 );
    nor g8083 ( n10914 , n37115 , n1830 );
    and g8084 ( n12498 , n9568 , n1108 );
    and g8085 ( n2664 , n22117 , n28396 );
    or g8086 ( n13680 , n32319 , n19742 );
    not g8087 ( n16418 , n13714 );
    or g8088 ( n32073 , n13830 , n24602 );
    not g8089 ( n22091 , n28202 );
    not g8090 ( n40728 , n3265 );
    xnor g8091 ( n27100 , n20487 , n16047 );
    and g8092 ( n38570 , n33286 , n12043 );
    or g8093 ( n24079 , n25005 , n9360 );
    or g8094 ( n40565 , n18249 , n24751 );
    or g8095 ( n17572 , n15986 , n20446 );
    not g8096 ( n40544 , n25397 );
    xnor g8097 ( n18338 , n29740 , n30447 );
    or g8098 ( n12958 , n37502 , n10530 );
    and g8099 ( n19143 , n10492 , n2028 );
    or g8100 ( n15669 , n17494 , n10682 );
    or g8101 ( n21266 , n5564 , n7436 );
    and g8102 ( n40212 , n5230 , n16036 );
    and g8103 ( n19284 , n14050 , n14872 );
    not g8104 ( n16403 , n18186 );
    and g8105 ( n41226 , n20455 , n28462 );
    xnor g8106 ( n25436 , n16820 , n30840 );
    or g8107 ( n17207 , n40240 , n34436 );
    nor g8108 ( n19970 , n8909 , n39431 );
    and g8109 ( n33708 , n29887 , n38076 );
    and g8110 ( n20049 , n12708 , n30236 );
    or g8111 ( n430 , n26746 , n342 );
    or g8112 ( n23133 , n21111 , n12879 );
    and g8113 ( n691 , n9706 , n17096 );
    and g8114 ( n17754 , n26293 , n3496 );
    nor g8115 ( n39030 , n12349 , n17278 );
    or g8116 ( n16674 , n7874 , n41079 );
    not g8117 ( n17704 , n4526 );
    or g8118 ( n27437 , n13368 , n6467 );
    and g8119 ( n3236 , n34601 , n23887 );
    and g8120 ( n474 , n29728 , n13792 );
    not g8121 ( n36696 , n8463 );
    nor g8122 ( n16802 , n5964 , n38532 );
    and g8123 ( n27962 , n36989 , n15896 );
    xnor g8124 ( n30534 , n24546 , n19962 );
    or g8125 ( n32282 , n22997 , n28958 );
    and g8126 ( n20680 , n4299 , n8291 );
    nor g8127 ( n31766 , n31818 , n18290 );
    not g8128 ( n28968 , n1794 );
    and g8129 ( n5079 , n39371 , n20731 );
    and g8130 ( n10751 , n16275 , n7132 );
    nor g8131 ( n7037 , n1507 , n6413 );
    or g8132 ( n14435 , n5142 , n33775 );
    or g8133 ( n38037 , n12245 , n10916 );
    not g8134 ( n36973 , n24876 );
    nor g8135 ( n31711 , n37874 , n29814 );
    or g8136 ( n35122 , n37212 , n3709 );
    or g8137 ( n30751 , n7186 , n25115 );
    and g8138 ( n34041 , n17677 , n3497 );
    not g8139 ( n41976 , n5282 );
    or g8140 ( n40242 , n14707 , n17499 );
    and g8141 ( n4987 , n12204 , n16758 );
    and g8142 ( n41674 , n2229 , n14637 );
    nor g8143 ( n19449 , n24441 , n2649 );
    and g8144 ( n20436 , n19995 , n41743 );
    and g8145 ( n28531 , n40721 , n42459 );
    or g8146 ( n7579 , n36844 , n33127 );
    or g8147 ( n10112 , n1470 , n41720 );
    nor g8148 ( n9080 , n31857 , n24776 );
    or g8149 ( n6062 , n41835 , n34715 );
    nor g8150 ( n5027 , n40092 , n26572 );
    or g8151 ( n27674 , n16267 , n14664 );
    not g8152 ( n9809 , n22306 );
    not g8153 ( n9608 , n40631 );
    xnor g8154 ( n25949 , n37235 , n18081 );
    and g8155 ( n25318 , n12301 , n30692 );
    not g8156 ( n768 , n25892 );
    and g8157 ( n41461 , n37159 , n22547 );
    or g8158 ( n33934 , n30030 , n9162 );
    or g8159 ( n6215 , n33027 , n6388 );
    nor g8160 ( n17034 , n20323 , n14853 );
    nor g8161 ( n31347 , n16620 , n39940 );
    or g8162 ( n11934 , n30420 , n15388 );
    and g8163 ( n9400 , n13389 , n187 );
    nor g8164 ( n40888 , n17120 , n29520 );
    or g8165 ( n30898 , n40501 , n40485 );
    nor g8166 ( n29532 , n15272 , n38040 );
    and g8167 ( n17346 , n1856 , n15583 );
    or g8168 ( n34709 , n27815 , n24931 );
    xnor g8169 ( n21520 , n19385 , n4256 );
    and g8170 ( n31011 , n18610 , n11343 );
    nor g8171 ( n12788 , n19045 , n9547 );
    and g8172 ( n9970 , n2048 , n19785 );
    nor g8173 ( n32043 , n35660 , n15232 );
    and g8174 ( n9647 , n27031 , n21688 );
    not g8175 ( n15894 , n35230 );
    and g8176 ( n20311 , n30474 , n1831 );
    xnor g8177 ( n12809 , n27960 , n40961 );
    and g8178 ( n23141 , n15686 , n12602 );
    or g8179 ( n8450 , n24499 , n40157 );
    xnor g8180 ( n2139 , n36009 , n7833 );
    xnor g8181 ( n17508 , n4712 , n10821 );
    not g8182 ( n31966 , n41155 );
    or g8183 ( n26610 , n26217 , n15267 );
    not g8184 ( n12068 , n39309 );
    or g8185 ( n34613 , n37333 , n40529 );
    xnor g8186 ( n38474 , n25041 , n17022 );
    or g8187 ( n34454 , n33511 , n2968 );
    or g8188 ( n5875 , n36250 , n22119 );
    and g8189 ( n32027 , n6785 , n10944 );
    or g8190 ( n24101 , n10306 , n39254 );
    and g8191 ( n30488 , n3186 , n3189 );
    nor g8192 ( n7526 , n10989 , n447 );
    not g8193 ( n9318 , n13720 );
    not g8194 ( n9833 , n13124 );
    or g8195 ( n1544 , n6509 , n1283 );
    nor g8196 ( n19675 , n11431 , n414 );
    xnor g8197 ( n17875 , n5146 , n6113 );
    not g8198 ( n34786 , n271 );
    and g8199 ( n9942 , n17393 , n15977 );
    xnor g8200 ( n20678 , n24113 , n11428 );
    not g8201 ( n33655 , n4756 );
    nor g8202 ( n17280 , n15590 , n7293 );
    not g8203 ( n23304 , n20737 );
    or g8204 ( n11686 , n327 , n27986 );
    or g8205 ( n30478 , n167 , n22364 );
    or g8206 ( n9493 , n29027 , n12913 );
    nor g8207 ( n14529 , n33351 , n23564 );
    and g8208 ( n13464 , n41137 , n26530 );
    nor g8209 ( n42693 , n23736 , n17135 );
    or g8210 ( n29839 , n7087 , n16967 );
    and g8211 ( n11152 , n17612 , n4536 );
    or g8212 ( n20433 , n23399 , n12947 );
    nor g8213 ( n2830 , n39605 , n32917 );
    and g8214 ( n10423 , n3840 , n35598 );
    or g8215 ( n10461 , n26099 , n6726 );
    not g8216 ( n20714 , n23915 );
    nor g8217 ( n13500 , n17592 , n26355 );
    not g8218 ( n10646 , n5254 );
    and g8219 ( n38245 , n2162 , n26602 );
    nor g8220 ( n39999 , n35501 , n24866 );
    or g8221 ( n37527 , n28847 , n15556 );
    nor g8222 ( n26873 , n28010 , n17157 );
    and g8223 ( n12317 , n7264 , n8779 );
    or g8224 ( n14332 , n4193 , n16027 );
    xnor g8225 ( n18062 , n7943 , n30216 );
    xnor g8226 ( n31337 , n38242 , n18458 );
    or g8227 ( n3605 , n2199 , n14608 );
    or g8228 ( n19292 , n19061 , n32060 );
    or g8229 ( n34312 , n1738 , n4669 );
    or g8230 ( n13198 , n22371 , n26403 );
    or g8231 ( n38083 , n13794 , n31232 );
    or g8232 ( n1955 , n17504 , n34939 );
    or g8233 ( n24860 , n31072 , n19793 );
    or g8234 ( n33090 , n15384 , n34670 );
    or g8235 ( n38683 , n19726 , n3764 );
    xnor g8236 ( n25723 , n1841 , n38623 );
    and g8237 ( n24893 , n34020 , n22747 );
    and g8238 ( n6592 , n26436 , n8605 );
    and g8239 ( n40859 , n12237 , n35669 );
    or g8240 ( n34801 , n27468 , n2599 );
    or g8241 ( n14165 , n24955 , n22885 );
    or g8242 ( n33880 , n38387 , n36432 );
    nor g8243 ( n11765 , n30506 , n34438 );
    nor g8244 ( n6189 , n5896 , n14949 );
    not g8245 ( n9353 , n15978 );
    or g8246 ( n22402 , n42115 , n29598 );
    xnor g8247 ( n23118 , n33937 , n42341 );
    and g8248 ( n9937 , n36031 , n28340 );
    nor g8249 ( n25686 , n761 , n12695 );
    and g8250 ( n19778 , n25891 , n707 );
    and g8251 ( n7028 , n36814 , n14249 );
    or g8252 ( n40251 , n27730 , n42296 );
    nor g8253 ( n28442 , n10716 , n28430 );
    or g8254 ( n9317 , n7616 , n30964 );
    or g8255 ( n21358 , n38042 , n19261 );
    not g8256 ( n5993 , n33199 );
    not g8257 ( n3317 , n25592 );
    or g8258 ( n39882 , n8501 , n33454 );
    xnor g8259 ( n35522 , n32470 , n5059 );
    or g8260 ( n31993 , n8848 , n31939 );
    or g8261 ( n40938 , n24879 , n20474 );
    not g8262 ( n29034 , n5842 );
    not g8263 ( n3034 , n13105 );
    or g8264 ( n34836 , n6220 , n41007 );
    or g8265 ( n17140 , n38797 , n23926 );
    nor g8266 ( n36738 , n37444 , n28296 );
    or g8267 ( n39931 , n8299 , n11814 );
    nor g8268 ( n25506 , n35310 , n25179 );
    not g8269 ( n7987 , n32009 );
    xnor g8270 ( n12137 , n22726 , n26079 );
    nor g8271 ( n1791 , n42481 , n16661 );
    not g8272 ( n35198 , n30557 );
    or g8273 ( n38234 , n15087 , n25677 );
    and g8274 ( n25047 , n12795 , n16979 );
    and g8275 ( n41497 , n35891 , n34210 );
    not g8276 ( n1927 , n29675 );
    or g8277 ( n4601 , n29367 , n37713 );
    not g8278 ( n17478 , n19127 );
    xnor g8279 ( n7881 , n19700 , n33623 );
    and g8280 ( n31914 , n40076 , n2613 );
    or g8281 ( n1342 , n36934 , n439 );
    nor g8282 ( n1090 , n33647 , n26595 );
    or g8283 ( n25944 , n3931 , n17456 );
    and g8284 ( n6073 , n24686 , n33881 );
    nor g8285 ( n31854 , n28502 , n23698 );
    xnor g8286 ( n29866 , n11436 , n34896 );
    and g8287 ( n4666 , n22228 , n40162 );
    or g8288 ( n20947 , n2095 , n20677 );
    or g8289 ( n14411 , n11737 , n14489 );
    not g8290 ( n37545 , n39298 );
    xnor g8291 ( n38392 , n13858 , n23644 );
    and g8292 ( n30312 , n13395 , n14409 );
    xnor g8293 ( n28907 , n32154 , n20354 );
    and g8294 ( n1638 , n36106 , n3614 );
    and g8295 ( n27252 , n34180 , n16954 );
    and g8296 ( n16715 , n40922 , n35609 );
    or g8297 ( n35008 , n31760 , n35732 );
    nor g8298 ( n32028 , n21987 , n6479 );
    not g8299 ( n12367 , n36843 );
    not g8300 ( n32543 , n21685 );
    xnor g8301 ( n3191 , n4218 , n20191 );
    xnor g8302 ( n40414 , n6841 , n19214 );
    not g8303 ( n8434 , n6148 );
    not g8304 ( n27 , n36315 );
    or g8305 ( n22852 , n7257 , n23392 );
    xnor g8306 ( n40707 , n8928 , n38255 );
    or g8307 ( n38681 , n5262 , n40646 );
    not g8308 ( n3557 , n38925 );
    and g8309 ( n24452 , n1402 , n12622 );
    and g8310 ( n30939 , n18446 , n22185 );
    and g8311 ( n4999 , n619 , n24990 );
    or g8312 ( n12222 , n19128 , n34681 );
    or g8313 ( n39111 , n36234 , n35425 );
    not g8314 ( n18381 , n20062 );
    not g8315 ( n41380 , n4086 );
    and g8316 ( n21499 , n8766 , n35137 );
    or g8317 ( n4430 , n37520 , n38016 );
    xnor g8318 ( n14342 , n13350 , n11792 );
    or g8319 ( n1566 , n34830 , n19095 );
    or g8320 ( n4498 , n10821 , n28028 );
    or g8321 ( n26315 , n24053 , n24740 );
    and g8322 ( n6798 , n8320 , n42213 );
    or g8323 ( n18210 , n19308 , n38266 );
    and g8324 ( n15882 , n2059 , n33519 );
    nor g8325 ( n12479 , n24917 , n37538 );
    xnor g8326 ( n33131 , n14969 , n41985 );
    xnor g8327 ( n34603 , n27363 , n32277 );
    or g8328 ( n11214 , n17256 , n4499 );
    or g8329 ( n42506 , n41066 , n19399 );
    and g8330 ( n26976 , n21566 , n4981 );
    or g8331 ( n26106 , n10902 , n11339 );
    and g8332 ( n27295 , n13543 , n20506 );
    or g8333 ( n19669 , n5956 , n34164 );
    or g8334 ( n14838 , n37980 , n31657 );
    and g8335 ( n25693 , n2369 , n28284 );
    or g8336 ( n12099 , n18236 , n36322 );
    and g8337 ( n28525 , n40817 , n3612 );
    and g8338 ( n13854 , n8937 , n6931 );
    not g8339 ( n24152 , n33028 );
    or g8340 ( n34484 , n28683 , n42098 );
    nor g8341 ( n4648 , n34298 , n42070 );
    and g8342 ( n28078 , n31143 , n32434 );
    xnor g8343 ( n15224 , n5658 , n7356 );
    or g8344 ( n28219 , n26910 , n1264 );
    or g8345 ( n18518 , n40184 , n14002 );
    or g8346 ( n28820 , n32087 , n35631 );
    nor g8347 ( n40989 , n16598 , n19325 );
    and g8348 ( n25789 , n32205 , n16880 );
    xnor g8349 ( n26063 , n35874 , n34199 );
    and g8350 ( n20231 , n14842 , n33123 );
    or g8351 ( n16238 , n29071 , n28447 );
    nor g8352 ( n14009 , n2199 , n14963 );
    or g8353 ( n42690 , n34477 , n41767 );
    and g8354 ( n8088 , n6172 , n12624 );
    nor g8355 ( n4236 , n6540 , n9944 );
    and g8356 ( n36944 , n42771 , n24381 );
    and g8357 ( n30070 , n17593 , n28284 );
    and g8358 ( n26149 , n31931 , n8520 );
    and g8359 ( n36647 , n17138 , n13722 );
    or g8360 ( n21890 , n22127 , n17921 );
    or g8361 ( n3031 , n3522 , n17044 );
    xnor g8362 ( n39846 , n4341 , n2563 );
    or g8363 ( n35821 , n35989 , n32402 );
    and g8364 ( n36456 , n18037 , n148 );
    nor g8365 ( n15563 , n5413 , n32258 );
    or g8366 ( n9954 , n18577 , n8531 );
    and g8367 ( n42349 , n21930 , n40793 );
    or g8368 ( n26564 , n41961 , n37143 );
    and g8369 ( n7874 , n33510 , n21964 );
    or g8370 ( n37704 , n13040 , n42694 );
    or g8371 ( n4328 , n35364 , n42786 );
    or g8372 ( n31660 , n36226 , n11989 );
    not g8373 ( n14098 , n20290 );
    or g8374 ( n17289 , n16467 , n1247 );
    not g8375 ( n21513 , n16646 );
    and g8376 ( n35010 , n1943 , n13225 );
    xnor g8377 ( n18829 , n21332 , n17062 );
    or g8378 ( n7769 , n39594 , n39520 );
    not g8379 ( n35382 , n35221 );
    or g8380 ( n887 , n10967 , n28130 );
    nor g8381 ( n8590 , n31542 , n12791 );
    xnor g8382 ( n32661 , n17087 , n38529 );
    nor g8383 ( n39409 , n1601 , n33500 );
    nor g8384 ( n17735 , n21736 , n30087 );
    nor g8385 ( n36171 , n31777 , n41972 );
    and g8386 ( n19115 , n35920 , n7369 );
    and g8387 ( n22896 , n4364 , n29691 );
    or g8388 ( n8804 , n11065 , n42533 );
    nor g8389 ( n9701 , n33981 , n15958 );
    or g8390 ( n25479 , n26565 , n9087 );
    and g8391 ( n1823 , n41945 , n27029 );
    or g8392 ( n2262 , n24062 , n32172 );
    or g8393 ( n38046 , n12687 , n20087 );
    xnor g8394 ( n25480 , n8175 , n23179 );
    not g8395 ( n32132 , n36372 );
    or g8396 ( n39352 , n23528 , n23053 );
    not g8397 ( n3343 , n1417 );
    or g8398 ( n29506 , n38132 , n20580 );
    not g8399 ( n42652 , n30826 );
    xnor g8400 ( n36656 , n36998 , n24521 );
    not g8401 ( n35931 , n8402 );
    nor g8402 ( n41447 , n14038 , n40122 );
    or g8403 ( n35975 , n41736 , n18299 );
    nor g8404 ( n16487 , n39571 , n19303 );
    xnor g8405 ( n8779 , n26794 , n41327 );
    nor g8406 ( n14145 , n20904 , n17504 );
    xnor g8407 ( n22843 , n41013 , n21481 );
    and g8408 ( n8886 , n8135 , n28509 );
    or g8409 ( n29759 , n33040 , n30935 );
    nor g8410 ( n4369 , n22482 , n37419 );
    or g8411 ( n7761 , n14407 , n22046 );
    or g8412 ( n22588 , n1507 , n2821 );
    not g8413 ( n5099 , n21480 );
    and g8414 ( n29140 , n8231 , n22508 );
    nor g8415 ( n2980 , n4919 , n22070 );
    and g8416 ( n42522 , n37874 , n29814 );
    or g8417 ( n11204 , n40702 , n37855 );
    nor g8418 ( n21663 , n14471 , n30511 );
    not g8419 ( n13121 , n5561 );
    not g8420 ( n6774 , n28530 );
    or g8421 ( n40804 , n9444 , n24371 );
    not g8422 ( n28152 , n33466 );
    or g8423 ( n24412 , n14313 , n256 );
    nor g8424 ( n37172 , n30430 , n41619 );
    not g8425 ( n16387 , n14823 );
    not g8426 ( n21697 , n15708 );
    or g8427 ( n17450 , n6560 , n9459 );
    or g8428 ( n24134 , n26744 , n38211 );
    and g8429 ( n3670 , n40779 , n3180 );
    and g8430 ( n4436 , n34484 , n2343 );
    xnor g8431 ( n12694 , n36046 , n40607 );
    and g8432 ( n40661 , n34852 , n23159 );
    or g8433 ( n35935 , n27452 , n6852 );
    and g8434 ( n31459 , n35397 , n35976 );
    xnor g8435 ( n8277 , n15524 , n19123 );
    not g8436 ( n37136 , n31205 );
    or g8437 ( n858 , n38 , n14290 );
    not g8438 ( n41642 , n29232 );
    and g8439 ( n23747 , n23976 , n16960 );
    or g8440 ( n36846 , n26611 , n21536 );
    or g8441 ( n13959 , n35629 , n23130 );
    and g8442 ( n29106 , n40506 , n35947 );
    not g8443 ( n28289 , n31728 );
    and g8444 ( n5380 , n18033 , n2979 );
    or g8445 ( n24853 , n14707 , n41129 );
    and g8446 ( n29422 , n16974 , n32517 );
    and g8447 ( n31472 , n32916 , n14714 );
    xnor g8448 ( n35107 , n26406 , n42177 );
    or g8449 ( n30933 , n24160 , n27700 );
    not g8450 ( n12808 , n24510 );
    not g8451 ( n12954 , n42554 );
    xnor g8452 ( n21039 , n1316 , n11494 );
    or g8453 ( n20226 , n41116 , n15794 );
    nor g8454 ( n3409 , n33981 , n4766 );
    not g8455 ( n38044 , n29334 );
    nor g8456 ( n20813 , n15426 , n3167 );
    not g8457 ( n22879 , n31089 );
    not g8458 ( n40725 , n5186 );
    nor g8459 ( n15048 , n30084 , n10405 );
    or g8460 ( n18218 , n3359 , n14410 );
    xnor g8461 ( n10390 , n17038 , n18889 );
    and g8462 ( n19179 , n37908 , n31212 );
    and g8463 ( n18705 , n29130 , n22966 );
    xnor g8464 ( n8831 , n32896 , n41672 );
    and g8465 ( n33902 , n40739 , n4167 );
    or g8466 ( n8472 , n1152 , n3746 );
    xnor g8467 ( n10647 , n39566 , n9096 );
    nor g8468 ( n32675 , n18275 , n18292 );
    nor g8469 ( n15348 , n37988 , n32209 );
    xnor g8470 ( n34083 , n3146 , n8330 );
    and g8471 ( n33585 , n15454 , n33005 );
    and g8472 ( n41238 , n39750 , n19222 );
    and g8473 ( n731 , n15378 , n12174 );
    nor g8474 ( n35548 , n38356 , n20604 );
    xnor g8475 ( n7405 , n12146 , n24740 );
    and g8476 ( n10574 , n6763 , n31275 );
    or g8477 ( n507 , n17943 , n27020 );
    xnor g8478 ( n12995 , n6420 , n26182 );
    xnor g8479 ( n10801 , n42047 , n2942 );
    or g8480 ( n41925 , n28876 , n30041 );
    nor g8481 ( n17180 , n36638 , n32932 );
    not g8482 ( n34187 , n24013 );
    not g8483 ( n13604 , n28362 );
    or g8484 ( n42729 , n6087 , n24571 );
    and g8485 ( n24583 , n24591 , n24649 );
    and g8486 ( n40947 , n11853 , n2090 );
    or g8487 ( n26109 , n14434 , n5466 );
    nor g8488 ( n1718 , n19227 , n6997 );
    or g8489 ( n8575 , n4108 , n22487 );
    or g8490 ( n27428 , n30971 , n9393 );
    or g8491 ( n18957 , n13783 , n30614 );
    and g8492 ( n35081 , n4324 , n22795 );
    xnor g8493 ( n35908 , n17087 , n21050 );
    or g8494 ( n2004 , n20728 , n10241 );
    or g8495 ( n5580 , n12397 , n15918 );
    or g8496 ( n6593 , n5718 , n17491 );
    nor g8497 ( n5476 , n14658 , n22671 );
    not g8498 ( n21561 , n9116 );
    not g8499 ( n27658 , n40912 );
    nor g8500 ( n27008 , n25727 , n23406 );
    nor g8501 ( n217 , n18948 , n32979 );
    nor g8502 ( n42088 , n12316 , n32323 );
    or g8503 ( n1805 , n6258 , n34344 );
    xnor g8504 ( n41525 , n37303 , n5964 );
    or g8505 ( n2505 , n14883 , n42544 );
    and g8506 ( n882 , n8727 , n13988 );
    not g8507 ( n8210 , n19861 );
    nor g8508 ( n27432 , n41293 , n14232 );
    or g8509 ( n30279 , n40815 , n11786 );
    xnor g8510 ( n34236 , n42118 , n21923 );
    or g8511 ( n39177 , n25600 , n2912 );
    not g8512 ( n27741 , n33455 );
    or g8513 ( n20267 , n13963 , n42344 );
    not g8514 ( n11393 , n9253 );
    and g8515 ( n33767 , n31395 , n11160 );
    or g8516 ( n40846 , n32879 , n32514 );
    not g8517 ( n42399 , n16247 );
    not g8518 ( n8031 , n14468 );
    xnor g8519 ( n38701 , n1838 , n13294 );
    and g8520 ( n10455 , n20507 , n40356 );
    xnor g8521 ( n29441 , n2839 , n23786 );
    not g8522 ( n13160 , n19178 );
    and g8523 ( n41927 , n22813 , n2606 );
    not g8524 ( n18840 , n23681 );
    and g8525 ( n24528 , n24095 , n15654 );
    or g8526 ( n3578 , n36806 , n16734 );
    or g8527 ( n19125 , n6889 , n34957 );
    nor g8528 ( n36323 , n7648 , n36387 );
    or g8529 ( n21017 , n94 , n37510 );
    or g8530 ( n36544 , n36929 , n18102 );
    and g8531 ( n31692 , n2702 , n18231 );
    and g8532 ( n18645 , n34349 , n21182 );
    and g8533 ( n42177 , n41085 , n4440 );
    or g8534 ( n15892 , n23880 , n7884 );
    not g8535 ( n29833 , n597 );
    or g8536 ( n34540 , n34939 , n36741 );
    nor g8537 ( n5789 , n17087 , n33813 );
    not g8538 ( n42256 , n40653 );
    or g8539 ( n14174 , n13665 , n904 );
    or g8540 ( n18682 , n15384 , n16692 );
    or g8541 ( n40030 , n35012 , n14909 );
    and g8542 ( n37690 , n5392 , n31816 );
    or g8543 ( n19585 , n24656 , n19533 );
    or g8544 ( n31885 , n37229 , n20921 );
    or g8545 ( n9746 , n34997 , n39786 );
    not g8546 ( n11445 , n10239 );
    nor g8547 ( n16142 , n907 , n37509 );
    or g8548 ( n27672 , n29593 , n19548 );
    xnor g8549 ( n28156 , n10078 , n26710 );
    or g8550 ( n8478 , n38259 , n15508 );
    or g8551 ( n14916 , n37662 , n12898 );
    xnor g8552 ( n34679 , n40883 , n32492 );
    xnor g8553 ( n15058 , n28443 , n41712 );
    nor g8554 ( n18105 , n34565 , n10694 );
    or g8555 ( n35485 , n17826 , n20273 );
    xnor g8556 ( n22285 , n29740 , n19915 );
    or g8557 ( n41949 , n27037 , n8746 );
    and g8558 ( n22450 , n3013 , n40892 );
    or g8559 ( n4359 , n31795 , n13447 );
    or g8560 ( n30789 , n41393 , n32252 );
    nor g8561 ( n28672 , n26377 , n24885 );
    and g8562 ( n8468 , n26392 , n27404 );
    or g8563 ( n16516 , n16052 , n22891 );
    and g8564 ( n28165 , n13593 , n17414 );
    not g8565 ( n11482 , n701 );
    not g8566 ( n5212 , n20423 );
    or g8567 ( n32845 , n16342 , n10149 );
    not g8568 ( n40305 , n3841 );
    or g8569 ( n17769 , n15116 , n32502 );
    xnor g8570 ( n20956 , n25884 , n5434 );
    and g8571 ( n1246 , n5561 , n16468 );
    or g8572 ( n20764 , n38224 , n9414 );
    nor g8573 ( n33017 , n29120 , n839 );
    not g8574 ( n19545 , n29379 );
    or g8575 ( n32906 , n29646 , n34688 );
    or g8576 ( n20255 , n779 , n4301 );
    or g8577 ( n30664 , n27792 , n33945 );
    or g8578 ( n21073 , n25669 , n9177 );
    nor g8579 ( n37945 , n2445 , n6464 );
    or g8580 ( n29456 , n34037 , n24056 );
    and g8581 ( n21128 , n28179 , n27569 );
    xnor g8582 ( n18529 , n8873 , n26288 );
    not g8583 ( n16575 , n13430 );
    not g8584 ( n36776 , n22812 );
    and g8585 ( n9501 , n26290 , n28744 );
    nor g8586 ( n5935 , n13474 , n25790 );
    or g8587 ( n6736 , n41283 , n5202 );
    or g8588 ( n30722 , n16897 , n41689 );
    or g8589 ( n19550 , n1816 , n12217 );
    or g8590 ( n40737 , n25906 , n467 );
    or g8591 ( n6805 , n2372 , n33635 );
    or g8592 ( n35875 , n22744 , n35382 );
    and g8593 ( n37793 , n24553 , n9339 );
    or g8594 ( n20233 , n17138 , n42407 );
    and g8595 ( n14124 , n25884 , n9007 );
    or g8596 ( n6888 , n787 , n5 );
    xnor g8597 ( n9311 , n18272 , n16918 );
    or g8598 ( n37985 , n30811 , n25030 );
    nor g8599 ( n15868 , n7763 , n36540 );
    or g8600 ( n8382 , n20311 , n2611 );
    xnor g8601 ( n26157 , n38629 , n33228 );
    or g8602 ( n27268 , n5428 , n1659 );
    and g8603 ( n3501 , n29689 , n12201 );
    or g8604 ( n24478 , n12652 , n7218 );
    or g8605 ( n26153 , n15837 , n29299 );
    or g8606 ( n42808 , n38485 , n14980 );
    or g8607 ( n848 , n28714 , n27127 );
    and g8608 ( n11189 , n29584 , n26610 );
    not g8609 ( n41513 , n13485 );
    or g8610 ( n10134 , n10090 , n3301 );
    not g8611 ( n8573 , n39766 );
    or g8612 ( n10919 , n13279 , n27782 );
    or g8613 ( n39496 , n10939 , n9044 );
    xnor g8614 ( n34856 , n4501 , n10237 );
    and g8615 ( n12740 , n13038 , n39052 );
    or g8616 ( n35820 , n4798 , n27779 );
    or g8617 ( n872 , n42192 , n27887 );
    and g8618 ( n40898 , n36009 , n5572 );
    or g8619 ( n10703 , n1292 , n16881 );
    not g8620 ( n13181 , n9671 );
    and g8621 ( n20302 , n16446 , n16400 );
    nor g8622 ( n29018 , n37146 , n40853 );
    and g8623 ( n31601 , n22580 , n20346 );
    and g8624 ( n8778 , n557 , n9230 );
    nor g8625 ( n2526 , n34752 , n12519 );
    not g8626 ( n17035 , n32078 );
    or g8627 ( n40438 , n6604 , n20127 );
    and g8628 ( n16578 , n39401 , n10189 );
    not g8629 ( n14307 , n20509 );
    not g8630 ( n17249 , n23430 );
    not g8631 ( n38973 , n10245 );
    xnor g8632 ( n29293 , n31989 , n31459 );
    xnor g8633 ( n40523 , n23964 , n27673 );
    not g8634 ( n23478 , n35871 );
    and g8635 ( n17037 , n6347 , n38539 );
    not g8636 ( n22597 , n21876 );
    not g8637 ( n6917 , n6309 );
    xnor g8638 ( n19468 , n27786 , n7148 );
    and g8639 ( n5729 , n23440 , n8856 );
    or g8640 ( n11219 , n13586 , n34716 );
    not g8641 ( n28185 , n18134 );
    or g8642 ( n29416 , n12526 , n31045 );
    or g8643 ( n10713 , n16793 , n12423 );
    nor g8644 ( n4757 , n4430 , n36083 );
    or g8645 ( n41174 , n21078 , n38550 );
    or g8646 ( n5421 , n21096 , n13500 );
    or g8647 ( n676 , n15718 , n20633 );
    and g8648 ( n27640 , n23248 , n10463 );
    or g8649 ( n39319 , n6673 , n11202 );
    nor g8650 ( n35336 , n30689 , n26537 );
    or g8651 ( n23433 , n31033 , n16145 );
    xnor g8652 ( n28851 , n19514 , n30603 );
    or g8653 ( n18301 , n13495 , n28441 );
    not g8654 ( n28725 , n28968 );
    or g8655 ( n18729 , n25784 , n14695 );
    or g8656 ( n883 , n8218 , n15757 );
    xnor g8657 ( n18153 , n34352 , n29241 );
    or g8658 ( n38551 , n11516 , n35643 );
    and g8659 ( n41326 , n27552 , n6675 );
    xnor g8660 ( n28293 , n38827 , n16568 );
    not g8661 ( n35992 , n8578 );
    or g8662 ( n38440 , n34974 , n34626 );
    or g8663 ( n20605 , n40784 , n39328 );
    xnor g8664 ( n37832 , n35965 , n6900 );
    or g8665 ( n25871 , n21152 , n38414 );
    and g8666 ( n25589 , n17431 , n22594 );
    or g8667 ( n14107 , n7341 , n27612 );
    or g8668 ( n39362 , n27329 , n18701 );
    and g8669 ( n17509 , n24648 , n23985 );
    or g8670 ( n3070 , n6423 , n27480 );
    or g8671 ( n30706 , n8897 , n24875 );
    not g8672 ( n13947 , n12786 );
    or g8673 ( n15298 , n13448 , n25303 );
    xnor g8674 ( n14521 , n28464 , n24195 );
    nor g8675 ( n13626 , n37939 , n33278 );
    or g8676 ( n40869 , n27388 , n36733 );
    or g8677 ( n34251 , n37678 , n15640 );
    or g8678 ( n13554 , n24797 , n6929 );
    and g8679 ( n21782 , n9707 , n6339 );
    nor g8680 ( n41348 , n23311 , n19922 );
    nor g8681 ( n20546 , n38454 , n14056 );
    and g8682 ( n39459 , n21101 , n1923 );
    or g8683 ( n15899 , n11629 , n9068 );
    xnor g8684 ( n20272 , n40391 , n7482 );
    not g8685 ( n10239 , n11830 );
    not g8686 ( n3379 , n41533 );
    or g8687 ( n12353 , n30756 , n11084 );
    or g8688 ( n18113 , n14434 , n26288 );
    or g8689 ( n26264 , n14487 , n40193 );
    and g8690 ( n35918 , n6579 , n40150 );
    or g8691 ( n29497 , n42792 , n39556 );
    not g8692 ( n26846 , n16075 );
    not g8693 ( n14467 , n35238 );
    and g8694 ( n3119 , n13719 , n19745 );
    and g8695 ( n11794 , n9669 , n12917 );
    or g8696 ( n36212 , n37854 , n18534 );
    or g8697 ( n29683 , n18070 , n25803 );
    xnor g8698 ( n32710 , n25118 , n3525 );
    nor g8699 ( n2345 , n38474 , n18202 );
    or g8700 ( n8609 , n2373 , n15035 );
    not g8701 ( n35663 , n33132 );
    not g8702 ( n8713 , n38055 );
    or g8703 ( n21213 , n31011 , n30896 );
    and g8704 ( n41331 , n40553 , n3354 );
    xnor g8705 ( n38697 , n37765 , n33953 );
    or g8706 ( n41257 , n7400 , n29895 );
    nor g8707 ( n32740 , n23052 , n2585 );
    or g8708 ( n238 , n13866 , n33630 );
    or g8709 ( n15017 , n20728 , n9406 );
    or g8710 ( n40582 , n27969 , n17475 );
    and g8711 ( n4333 , n8620 , n7880 );
    or g8712 ( n10761 , n22647 , n13572 );
    or g8713 ( n17177 , n40926 , n37951 );
    and g8714 ( n10913 , n9033 , n30805 );
    xnor g8715 ( n11014 , n8873 , n7 );
    nor g8716 ( n16305 , n1158 , n27 );
    nor g8717 ( n11773 , n24356 , n41080 );
    nor g8718 ( n27201 , n26185 , n7251 );
    and g8719 ( n36217 , n32868 , n33493 );
    or g8720 ( n32941 , n22920 , n19151 );
    not g8721 ( n30287 , n40600 );
    not g8722 ( n39744 , n33593 );
    and g8723 ( n7398 , n29359 , n15494 );
    or g8724 ( n37655 , n4006 , n11404 );
    or g8725 ( n31020 , n7486 , n40695 );
    or g8726 ( n14451 , n11798 , n32038 );
    nor g8727 ( n16504 , n19079 , n12835 );
    or g8728 ( n21379 , n20623 , n17937 );
    xnor g8729 ( n32139 , n3052 , n2842 );
    not g8730 ( n38761 , n26056 );
    not g8731 ( n32913 , n31702 );
    or g8732 ( n2851 , n20611 , n23856 );
    xnor g8733 ( n9810 , n24093 , n40492 );
    or g8734 ( n39534 , n38494 , n5555 );
    xnor g8735 ( n15219 , n32297 , n4580 );
    and g8736 ( n282 , n5019 , n7271 );
    and g8737 ( n4241 , n42611 , n20188 );
    not g8738 ( n8617 , n11851 );
    not g8739 ( n19326 , n26846 );
    nor g8740 ( n6891 , n23723 , n17733 );
    or g8741 ( n24788 , n10054 , n12565 );
    not g8742 ( n22056 , n23664 );
    not g8743 ( n1341 , n14380 );
    or g8744 ( n42352 , n17670 , n42544 );
    or g8745 ( n41874 , n19469 , n8159 );
    or g8746 ( n34455 , n4717 , n12545 );
    or g8747 ( n19524 , n29930 , n24723 );
    xnor g8748 ( n31177 , n2659 , n41706 );
    xnor g8749 ( n18187 , n18146 , n37867 );
    or g8750 ( n2325 , n39821 , n425 );
    nor g8751 ( n27238 , n31675 , n4566 );
    and g8752 ( n21069 , n14918 , n7919 );
    nor g8753 ( n30027 , n1355 , n36671 );
    or g8754 ( n15535 , n36099 , n4411 );
    and g8755 ( n28308 , n10653 , n31412 );
    nor g8756 ( n32325 , n22725 , n42403 );
    or g8757 ( n37374 , n30566 , n37848 );
    or g8758 ( n27197 , n22354 , n2296 );
    or g8759 ( n23361 , n23462 , n26704 );
    and g8760 ( n38429 , n18988 , n758 );
    not g8761 ( n41633 , n36509 );
    or g8762 ( n17040 , n28883 , n180 );
    not g8763 ( n23158 , n34126 );
    and g8764 ( n4076 , n34439 , n34615 );
    xnor g8765 ( n7850 , n41607 , n26073 );
    not g8766 ( n13899 , n8232 );
    or g8767 ( n38889 , n27412 , n9195 );
    or g8768 ( n15929 , n37548 , n24077 );
    xnor g8769 ( n25342 , n17225 , n11093 );
    nor g8770 ( n18523 , n10675 , n5982 );
    xnor g8771 ( n20705 , n37539 , n33746 );
    nor g8772 ( n18585 , n41844 , n22689 );
    or g8773 ( n8181 , n20073 , n40541 );
    not g8774 ( n7076 , n1151 );
    and g8775 ( n34907 , n24476 , n24971 );
    not g8776 ( n12640 , n7658 );
    and g8777 ( n34415 , n12817 , n34068 );
    or g8778 ( n4042 , n32217 , n17398 );
    or g8779 ( n3272 , n20538 , n37204 );
    nor g8780 ( n40038 , n24745 , n28375 );
    not g8781 ( n18070 , n30845 );
    not g8782 ( n9827 , n10614 );
    or g8783 ( n37052 , n17845 , n19363 );
    or g8784 ( n4966 , n25335 , n26316 );
    nor g8785 ( n42108 , n4140 , n16311 );
    xnor g8786 ( n6473 , n20487 , n35948 );
    xnor g8787 ( n29781 , n11133 , n29965 );
    not g8788 ( n24674 , n6469 );
    not g8789 ( n41767 , n30014 );
    and g8790 ( n39997 , n16918 , n18272 );
    nor g8791 ( n12981 , n33430 , n33409 );
    or g8792 ( n17718 , n20030 , n3155 );
    xnor g8793 ( n6133 , n11051 , n17569 );
    or g8794 ( n10298 , n36807 , n37468 );
    xnor g8795 ( n16314 , n9927 , n31929 );
    not g8796 ( n28177 , n40496 );
    not g8797 ( n18238 , n10611 );
    and g8798 ( n40080 , n19295 , n15155 );
    or g8799 ( n16961 , n12130 , n2901 );
    not g8800 ( n14851 , n341 );
    and g8801 ( n42395 , n20347 , n4476 );
    xnor g8802 ( n6232 , n28573 , n29802 );
    or g8803 ( n1764 , n15218 , n2152 );
    or g8804 ( n24312 , n14481 , n10178 );
    not g8805 ( n24449 , n22745 );
    not g8806 ( n12153 , n30826 );
    or g8807 ( n27716 , n42800 , n35701 );
    or g8808 ( n38294 , n28149 , n23542 );
    or g8809 ( n37827 , n722 , n15573 );
    or g8810 ( n14559 , n28837 , n27458 );
    nor g8811 ( n7093 , n41941 , n28164 );
    nor g8812 ( n39495 , n31284 , n35279 );
    or g8813 ( n17920 , n18798 , n293 );
    or g8814 ( n31251 , n34997 , n10718 );
    not g8815 ( n24914 , n26706 );
    xnor g8816 ( n1818 , n31989 , n40241 );
    or g8817 ( n34137 , n25150 , n22126 );
    or g8818 ( n31483 , n870 , n33926 );
    or g8819 ( n17562 , n33356 , n36182 );
    or g8820 ( n36239 , n2265 , n15186 );
    nor g8821 ( n7651 , n38242 , n1300 );
    or g8822 ( n41274 , n20699 , n21569 );
    or g8823 ( n29353 , n35289 , n37161 );
    or g8824 ( n28144 , n40455 , n2202 );
    not g8825 ( n23880 , n205 );
    and g8826 ( n34616 , n39240 , n28833 );
    or g8827 ( n37162 , n42260 , n2565 );
    or g8828 ( n19754 , n37208 , n24042 );
    and g8829 ( n41305 , n35575 , n41696 );
    or g8830 ( n35516 , n36345 , n26463 );
    or g8831 ( n7734 , n6802 , n19479 );
    xnor g8832 ( n35245 , n17823 , n20660 );
    or g8833 ( n3830 , n33337 , n500 );
    and g8834 ( n35422 , n42292 , n41882 );
    or g8835 ( n22540 , n12166 , n29322 );
    not g8836 ( n13771 , n38478 );
    or g8837 ( n21565 , n31004 , n36962 );
    or g8838 ( n17203 , n41288 , n30841 );
    or g8839 ( n13456 , n25964 , n19370 );
    xnor g8840 ( n40578 , n8694 , n3192 );
    nor g8841 ( n30390 , n18488 , n19974 );
    and g8842 ( n7374 , n32896 , n41672 );
    nor g8843 ( n4195 , n18866 , n38999 );
    not g8844 ( n5888 , n35027 );
    or g8845 ( n40592 , n6929 , n3959 );
    not g8846 ( n36661 , n39764 );
    or g8847 ( n6223 , n11823 , n1703 );
    or g8848 ( n9505 , n2056 , n33859 );
    and g8849 ( n3884 , n22237 , n39610 );
    and g8850 ( n18480 , n20110 , n7709 );
    and g8851 ( n11904 , n40575 , n30724 );
    or g8852 ( n14447 , n12666 , n38036 );
    xnor g8853 ( n13418 , n10427 , n24902 );
    and g8854 ( n39814 , n28819 , n21841 );
    xnor g8855 ( n6104 , n40 , n23888 );
    not g8856 ( n21006 , n1931 );
    and g8857 ( n28913 , n1046 , n5483 );
    or g8858 ( n38199 , n40773 , n17547 );
    not g8859 ( n12947 , n5661 );
    and g8860 ( n36971 , n17020 , n26721 );
    nor g8861 ( n21100 , n20167 , n1226 );
    not g8862 ( n15185 , n22634 );
    or g8863 ( n20188 , n33410 , n39098 );
    xnor g8864 ( n19174 , n28648 , n14800 );
    or g8865 ( n10273 , n22221 , n40955 );
    or g8866 ( n31668 , n2735 , n25597 );
    or g8867 ( n24460 , n38223 , n31997 );
    and g8868 ( n28405 , n2962 , n381 );
    and g8869 ( n11034 , n25066 , n27739 );
    or g8870 ( n31342 , n16748 , n13866 );
    xnor g8871 ( n15390 , n15776 , n39243 );
    or g8872 ( n10712 , n29440 , n29659 );
    and g8873 ( n18728 , n10993 , n38154 );
    and g8874 ( n37730 , n7002 , n22080 );
    and g8875 ( n37526 , n2186 , n977 );
    and g8876 ( n18787 , n36998 , n8647 );
    nor g8877 ( n895 , n9793 , n32133 );
    or g8878 ( n11251 , n24585 , n31879 );
    or g8879 ( n38692 , n32185 , n12867 );
    or g8880 ( n36228 , n31897 , n5796 );
    or g8881 ( n22257 , n12136 , n8676 );
    or g8882 ( n37370 , n18274 , n28140 );
    or g8883 ( n30520 , n4292 , n32766 );
    and g8884 ( n29653 , n29 , n18769 );
    or g8885 ( n38811 , n28795 , n31083 );
    and g8886 ( n27785 , n17787 , n29563 );
    or g8887 ( n21795 , n37090 , n36848 );
    or g8888 ( n28964 , n6577 , n28117 );
    nor g8889 ( n23627 , n3817 , n32503 );
    or g8890 ( n18223 , n23627 , n14267 );
    not g8891 ( n40318 , n35536 );
    xnor g8892 ( n7409 , n42825 , n38671 );
    or g8893 ( n11343 , n17984 , n24340 );
    or g8894 ( n31610 , n11184 , n39932 );
    and g8895 ( n38797 , n2568 , n32280 );
    nor g8896 ( n18267 , n1719 , n34143 );
    xnor g8897 ( n32187 , n7922 , n38980 );
    and g8898 ( n8094 , n16644 , n35641 );
    xnor g8899 ( n12261 , n17377 , n35280 );
    or g8900 ( n10948 , n23509 , n12238 );
    or g8901 ( n5880 , n4140 , n1123 );
    or g8902 ( n15902 , n17214 , n41337 );
    and g8903 ( n2777 , n29875 , n22223 );
    and g8904 ( n13428 , n21491 , n13026 );
    nor g8905 ( n34155 , n32922 , n11455 );
    xnor g8906 ( n40664 , n10004 , n7594 );
    xnor g8907 ( n14361 , n32134 , n25227 );
    or g8908 ( n38186 , n11129 , n3543 );
    and g8909 ( n27162 , n3721 , n25405 );
    nor g8910 ( n722 , n14566 , n41991 );
    or g8911 ( n35893 , n2193 , n15088 );
    nor g8912 ( n1890 , n34731 , n22483 );
    or g8913 ( n40399 , n38157 , n1141 );
    not g8914 ( n21470 , n23145 );
    xnor g8915 ( n28101 , n27184 , n37706 );
    xnor g8916 ( n30539 , n36009 , n26984 );
    xnor g8917 ( n25797 , n105 , n35554 );
    nor g8918 ( n28540 , n22484 , n26667 );
    and g8919 ( n21926 , n26347 , n8497 );
    xnor g8920 ( n11203 , n7969 , n33093 );
    or g8921 ( n13167 , n7678 , n1412 );
    and g8922 ( n30031 , n38997 , n19046 );
    or g8923 ( n15786 , n12850 , n14749 );
    or g8924 ( n8677 , n18595 , n19484 );
    xnor g8925 ( n9535 , n7922 , n1583 );
    and g8926 ( n12696 , n11384 , n9053 );
    not g8927 ( n7172 , n9814 );
    xnor g8928 ( n25209 , n18972 , n13189 );
    or g8929 ( n18979 , n27932 , n16921 );
    nor g8930 ( n32962 , n33652 , n28421 );
    and g8931 ( n7663 , n5182 , n11358 );
    and g8932 ( n20866 , n29351 , n20550 );
    or g8933 ( n5705 , n30957 , n12051 );
    nor g8934 ( n29962 , n11923 , n25151 );
    xnor g8935 ( n40922 , n29476 , n29071 );
    or g8936 ( n23785 , n42191 , n4043 );
    not g8937 ( n9884 , n35199 );
    not g8938 ( n18435 , n33885 );
    and g8939 ( n38849 , n4210 , n18939 );
    and g8940 ( n35157 , n2890 , n18568 );
    nor g8941 ( n11790 , n41380 , n13924 );
    and g8942 ( n20068 , n10210 , n37986 );
    or g8943 ( n9249 , n4798 , n10563 );
    xnor g8944 ( n11609 , n36998 , n9574 );
    or g8945 ( n13417 , n20684 , n22071 );
    or g8946 ( n23338 , n5718 , n30920 );
    xnor g8947 ( n10319 , n9783 , n39939 );
    and g8948 ( n23171 , n10613 , n32984 );
    not g8949 ( n13050 , n21818 );
    xnor g8950 ( n38101 , n18880 , n33487 );
    not g8951 ( n29163 , n29948 );
    and g8952 ( n9012 , n17824 , n15810 );
    not g8953 ( n20608 , n11264 );
    xnor g8954 ( n28604 , n36622 , n42879 );
    or g8955 ( n35404 , n25101 , n23956 );
    or g8956 ( n26618 , n12790 , n22675 );
    and g8957 ( n28572 , n36375 , n41552 );
    or g8958 ( n15713 , n32087 , n37435 );
    xnor g8959 ( n13929 , n36073 , n2199 );
    and g8960 ( n39612 , n21493 , n8298 );
    or g8961 ( n13037 , n18186 , n25035 );
    and g8962 ( n10727 , n17076 , n17801 );
    or g8963 ( n14094 , n34017 , n13702 );
    xnor g8964 ( n1437 , n37709 , n12729 );
    xnor g8965 ( n23070 , n4511 , n8078 );
    and g8966 ( n2412 , n5487 , n36650 );
    not g8967 ( n33674 , n20691 );
    not g8968 ( n3751 , n11418 );
    and g8969 ( n6328 , n42326 , n40268 );
    and g8970 ( n18822 , n16218 , n27937 );
    not g8971 ( n39687 , n4929 );
    nor g8972 ( n3325 , n13006 , n21414 );
    and g8973 ( n12888 , n36980 , n17389 );
    or g8974 ( n41299 , n38640 , n17631 );
    not g8975 ( n22191 , n16820 );
    not g8976 ( n19347 , n22784 );
    nor g8977 ( n25039 , n10456 , n31869 );
    and g8978 ( n10326 , n622 , n6345 );
    not g8979 ( n6621 , n21246 );
    or g8980 ( n35389 , n21387 , n7355 );
    or g8981 ( n9875 , n38996 , n3083 );
    xnor g8982 ( n30950 , n21888 , n28765 );
    or g8983 ( n1873 , n25033 , n12371 );
    or g8984 ( n16019 , n5913 , n31561 );
    not g8985 ( n26268 , n3137 );
    and g8986 ( n3907 , n17156 , n35943 );
    or g8987 ( n18108 , n26582 , n17575 );
    or g8988 ( n19906 , n26431 , n23012 );
    nor g8989 ( n40302 , n28036 , n10025 );
    and g8990 ( n30072 , n2509 , n2139 );
    or g8991 ( n29204 , n463 , n32285 );
    xnor g8992 ( n14571 , n37484 , n10598 );
    and g8993 ( n21277 , n25231 , n20725 );
    nor g8994 ( n12658 , n23942 , n10087 );
    not g8995 ( n41614 , n30048 );
    or g8996 ( n34558 , n27980 , n25078 );
    or g8997 ( n25745 , n24903 , n23328 );
    or g8998 ( n22834 , n36367 , n22631 );
    or g8999 ( n3474 , n18282 , n41035 );
    nor g9000 ( n30536 , n1683 , n36335 );
    nor g9001 ( n20394 , n3864 , n40376 );
    or g9002 ( n1660 , n2372 , n5210 );
    and g9003 ( n23743 , n26883 , n10415 );
    or g9004 ( n7270 , n5072 , n10666 );
    and g9005 ( n15113 , n1400 , n1492 );
    or g9006 ( n10492 , n19509 , n41981 );
    nor g9007 ( n32645 , n5625 , n27576 );
    and g9008 ( n38799 , n37473 , n38425 );
    or g9009 ( n42456 , n24167 , n41336 );
    not g9010 ( n2990 , n24899 );
    or g9011 ( n36497 , n26932 , n15137 );
    or g9012 ( n26510 , n35294 , n30967 );
    and g9013 ( n37960 , n37148 , n11252 );
    or g9014 ( n33614 , n9417 , n7878 );
    xnor g9015 ( n16339 , n3934 , n5707 );
    or g9016 ( n37145 , n8222 , n3487 );
    or g9017 ( n13674 , n5525 , n5458 );
    or g9018 ( n4805 , n41356 , n25245 );
    or g9019 ( n17517 , n28551 , n15212 );
    xnor g9020 ( n33400 , n31989 , n31751 );
    or g9021 ( n34541 , n1205 , n7935 );
    xnor g9022 ( n32161 , n21605 , n10342 );
    not g9023 ( n36298 , n29648 );
    and g9024 ( n42821 , n29775 , n35936 );
    and g9025 ( n12807 , n9348 , n1498 );
    or g9026 ( n24247 , n5408 , n4575 );
    and g9027 ( n5173 , n42752 , n22082 );
    xnor g9028 ( n15288 , n29667 , n17985 );
    or g9029 ( n23595 , n33030 , n14837 );
    xnor g9030 ( n4791 , n30576 , n14760 );
    or g9031 ( n16274 , n30288 , n23878 );
    and g9032 ( n42511 , n12488 , n34915 );
    or g9033 ( n16240 , n8426 , n19360 );
    or g9034 ( n27222 , n17486 , n5022 );
    and g9035 ( n37552 , n1130 , n24270 );
    or g9036 ( n2038 , n15184 , n26205 );
    not g9037 ( n32455 , n3599 );
    or g9038 ( n3966 , n1107 , n42420 );
    and g9039 ( n24107 , n5064 , n20915 );
    and g9040 ( n18660 , n12066 , n36695 );
    or g9041 ( n14127 , n40186 , n1961 );
    not g9042 ( n821 , n21419 );
    nor g9043 ( n661 , n31987 , n28070 );
    xnor g9044 ( n39477 , n8255 , n15942 );
    xnor g9045 ( n37085 , n41515 , n29111 );
    not g9046 ( n21631 , n41618 );
    and g9047 ( n21176 , n29976 , n2474 );
    not g9048 ( n19361 , n33214 );
    and g9049 ( n23917 , n34154 , n13363 );
    and g9050 ( n27353 , n10443 , n33221 );
    or g9051 ( n35854 , n37038 , n8595 );
    nor g9052 ( n8970 , n24991 , n10191 );
    or g9053 ( n7748 , n27835 , n37622 );
    nor g9054 ( n26023 , n5674 , n33872 );
    or g9055 ( n15132 , n20120 , n4281 );
    not g9056 ( n3465 , n14280 );
    or g9057 ( n15767 , n42367 , n5315 );
    xnor g9058 ( n3894 , n14953 , n2178 );
    not g9059 ( n19512 , n12810 );
    xnor g9060 ( n23256 , n26700 , n38714 );
    or g9061 ( n35415 , n1507 , n1203 );
    or g9062 ( n18479 , n16602 , n34079 );
    and g9063 ( n38338 , n30765 , n42330 );
    nor g9064 ( n37411 , n14537 , n11729 );
    and g9065 ( n25194 , n20483 , n28084 );
    or g9066 ( n18595 , n19103 , n36962 );
    or g9067 ( n6785 , n40389 , n31902 );
    or g9068 ( n40373 , n9794 , n4569 );
    or g9069 ( n35022 , n20626 , n425 );
    xnor g9070 ( n11902 , n32297 , n3860 );
    or g9071 ( n38253 , n9809 , n9283 );
    not g9072 ( n17955 , n24700 );
    or g9073 ( n5191 , n15547 , n27663 );
    or g9074 ( n31189 , n28675 , n32406 );
    or g9075 ( n13451 , n9752 , n32114 );
    or g9076 ( n26702 , n10953 , n12015 );
    or g9077 ( n3800 , n34544 , n21064 );
    or g9078 ( n25183 , n30737 , n3708 );
    and g9079 ( n2649 , n19489 , n42271 );
    or g9080 ( n2229 , n27714 , n28351 );
    or g9081 ( n34837 , n16792 , n16224 );
    and g9082 ( n26869 , n31793 , n11422 );
    or g9083 ( n30388 , n40685 , n42856 );
    xnor g9084 ( n20113 , n35090 , n20982 );
    and g9085 ( n37016 , n11945 , n17206 );
    xnor g9086 ( n10808 , n4558 , n30690 );
    xnor g9087 ( n41335 , n26745 , n14720 );
    not g9088 ( n18902 , n12548 );
    not g9089 ( n30788 , n23650 );
    xnor g9090 ( n38100 , n7978 , n30221 );
    or g9091 ( n6511 , n40422 , n17229 );
    not g9092 ( n8649 , n40772 );
    and g9093 ( n11575 , n18803 , n12660 );
    and g9094 ( n37258 , n5032 , n25211 );
    xnor g9095 ( n26534 , n31099 , n3097 );
    or g9096 ( n33551 , n3446 , n10687 );
    or g9097 ( n1119 , n16505 , n20328 );
    or g9098 ( n14644 , n16663 , n30652 );
    or g9099 ( n9442 , n4669 , n3598 );
    nor g9100 ( n23422 , n6072 , n267 );
    and g9101 ( n37842 , n23166 , n40850 );
    not g9102 ( n2017 , n20403 );
    or g9103 ( n26141 , n20934 , n40245 );
    or g9104 ( n37104 , n20250 , n5892 );
    not g9105 ( n617 , n22958 );
    and g9106 ( n15526 , n11550 , n35547 );
    or g9107 ( n10711 , n20138 , n24572 );
    not g9108 ( n34281 , n29959 );
    not g9109 ( n40 , n17120 );
    nor g9110 ( n12169 , n25173 , n42518 );
    and g9111 ( n38781 , n31987 , n28070 );
    or g9112 ( n2329 , n39276 , n17692 );
    or g9113 ( n6610 , n1380 , n20503 );
    or g9114 ( n26883 , n17654 , n34503 );
    not g9115 ( n37760 , n27942 );
    nor g9116 ( n21636 , n38879 , n23621 );
    or g9117 ( n34530 , n28402 , n25038 );
    not g9118 ( n6379 , n40136 );
    or g9119 ( n6603 , n31584 , n22770 );
    or g9120 ( n12327 , n37191 , n4209 );
    and g9121 ( n41547 , n10919 , n4835 );
    or g9122 ( n32759 , n10673 , n15900 );
    or g9123 ( n13497 , n10996 , n42185 );
    or g9124 ( n12976 , n40384 , n35294 );
    and g9125 ( n14963 , n3865 , n5381 );
    and g9126 ( n24521 , n3376 , n989 );
    nor g9127 ( n13490 , n3139 , n20460 );
    and g9128 ( n35045 , n2351 , n30813 );
    and g9129 ( n1717 , n22255 , n32404 );
    not g9130 ( n4512 , n6205 );
    or g9131 ( n42040 , n10467 , n9145 );
    and g9132 ( n17985 , n4080 , n4051 );
    or g9133 ( n7345 , n6319 , n23551 );
    or g9134 ( n38144 , n23714 , n20712 );
    or g9135 ( n18369 , n2754 , n16902 );
    and g9136 ( n12620 , n29040 , n1998 );
    or g9137 ( n7211 , n28745 , n33950 );
    nor g9138 ( n959 , n16598 , n13852 );
    not g9139 ( n5915 , n36762 );
    and g9140 ( n33269 , n15495 , n34701 );
    and g9141 ( n36370 , n4334 , n22856 );
    or g9142 ( n22062 , n36671 , n38569 );
    and g9143 ( n28297 , n17966 , n26605 );
    xnor g9144 ( n18362 , n6052 , n27828 );
    xnor g9145 ( n11469 , n30264 , n12831 );
    and g9146 ( n37749 , n39435 , n28427 );
    xnor g9147 ( n28183 , n22263 , n2791 );
    and g9148 ( n34750 , n9094 , n4118 );
    and g9149 ( n31578 , n9968 , n17223 );
    and g9150 ( n40608 , n7642 , n32849 );
    xnor g9151 ( n38344 , n31099 , n26638 );
    and g9152 ( n38538 , n2485 , n5135 );
    nor g9153 ( n32855 , n32753 , n20905 );
    or g9154 ( n9053 , n10860 , n34085 );
    or g9155 ( n24673 , n40218 , n9040 );
    not g9156 ( n33332 , n29025 );
    or g9157 ( n26215 , n39195 , n22439 );
    and g9158 ( n28344 , n34379 , n34541 );
    or g9159 ( n36194 , n1148 , n16236 );
    and g9160 ( n9357 , n4186 , n7517 );
    xnor g9161 ( n2274 , n23686 , n18139 );
    or g9162 ( n36463 , n34642 , n18622 );
    or g9163 ( n21758 , n40710 , n20526 );
    nor g9164 ( n6392 , n27190 , n5514 );
    and g9165 ( n844 , n16788 , n40903 );
    not g9166 ( n39159 , n20592 );
    xnor g9167 ( n28026 , n33884 , n5440 );
    or g9168 ( n38365 , n39457 , n6316 );
    nor g9169 ( n19003 , n24115 , n1988 );
    or g9170 ( n4741 , n1387 , n27709 );
    or g9171 ( n14774 , n13385 , n41584 );
    or g9172 ( n32763 , n38996 , n10130 );
    or g9173 ( n21274 , n40283 , n18574 );
    xnor g9174 ( n630 , n25367 , n5896 );
    and g9175 ( n27270 , n9149 , n30026 );
    or g9176 ( n5112 , n41228 , n6628 );
    not g9177 ( n30308 , n33554 );
    or g9178 ( n13561 , n801 , n30436 );
    xnor g9179 ( n16279 , n18530 , n39196 );
    or g9180 ( n24690 , n38960 , n14776 );
    or g9181 ( n27665 , n3853 , n24307 );
    or g9182 ( n36361 , n41247 , n35159 );
    not g9183 ( n18946 , n22399 );
    not g9184 ( n5186 , n36696 );
    or g9185 ( n25358 , n39559 , n4363 );
    or g9186 ( n2942 , n29039 , n33724 );
    and g9187 ( n7824 , n23506 , n32761 );
    nor g9188 ( n20429 , n36009 , n5572 );
    nor g9189 ( n14016 , n8494 , n36130 );
    xnor g9190 ( n26243 , n31099 , n23420 );
    or g9191 ( n12571 , n40389 , n20424 );
    xnor g9192 ( n31092 , n10005 , n10529 );
    or g9193 ( n10280 , n20720 , n36608 );
    and g9194 ( n19828 , n32834 , n16289 );
    or g9195 ( n20962 , n8494 , n42510 );
    not g9196 ( n325 , n25406 );
    nor g9197 ( n42502 , n17932 , n4779 );
    and g9198 ( n35070 , n19597 , n30618 );
    and g9199 ( n27292 , n29866 , n38700 );
    or g9200 ( n8950 , n13486 , n18222 );
    xnor g9201 ( n35472 , n40886 , n33504 );
    and g9202 ( n4212 , n3731 , n22775 );
    or g9203 ( n29036 , n31111 , n37336 );
    or g9204 ( n26381 , n26961 , n16578 );
    or g9205 ( n38575 , n25588 , n42746 );
    xnor g9206 ( n4324 , n2182 , n42408 );
    and g9207 ( n364 , n9433 , n35444 );
    or g9208 ( n21629 , n21582 , n4463 );
    or g9209 ( n15583 , n26884 , n36613 );
    xnor g9210 ( n23945 , n32351 , n30064 );
    or g9211 ( n17462 , n15934 , n40238 );
    not g9212 ( n15696 , n10881 );
    or g9213 ( n7594 , n31264 , n39357 );
    and g9214 ( n40748 , n2572 , n35345 );
    and g9215 ( n13155 , n35968 , n28220 );
    and g9216 ( n19450 , n1285 , n25114 );
    or g9217 ( n20073 , n1006 , n20210 );
    not g9218 ( n40612 , n22953 );
    xnor g9219 ( n17698 , n6841 , n5983 );
    nor g9220 ( n38185 , n21745 , n16168 );
    or g9221 ( n10644 , n14140 , n30926 );
    or g9222 ( n8990 , n13737 , n1404 );
    or g9223 ( n27625 , n32100 , n38969 );
    xnor g9224 ( n19628 , n20548 , n39033 );
    not g9225 ( n28065 , n38662 );
    or g9226 ( n6341 , n7008 , n19387 );
    or g9227 ( n33627 , n32369 , n8599 );
    or g9228 ( n25328 , n7992 , n34102 );
    or g9229 ( n22629 , n19810 , n1707 );
    xnor g9230 ( n15290 , n9827 , n11507 );
    and g9231 ( n2113 , n29417 , n37934 );
    or g9232 ( n32002 , n25279 , n31534 );
    or g9233 ( n32560 , n10282 , n38319 );
    or g9234 ( n1909 , n10634 , n32239 );
    not g9235 ( n37547 , n17638 );
    nor g9236 ( n20580 , n20039 , n13807 );
    xnor g9237 ( n1129 , n24584 , n5143 );
    and g9238 ( n37579 , n29873 , n28299 );
    nor g9239 ( n26225 , n36426 , n25914 );
    or g9240 ( n34587 , n1189 , n40455 );
    and g9241 ( n21084 , n26645 , n8016 );
    or g9242 ( n19934 , n12197 , n990 );
    or g9243 ( n29878 , n33772 , n34209 );
    or g9244 ( n297 , n33981 , n35013 );
    xnor g9245 ( n26165 , n6625 , n41888 );
    or g9246 ( n6391 , n25904 , n11629 );
    not g9247 ( n15662 , n10757 );
    or g9248 ( n35108 , n22824 , n15930 );
    nor g9249 ( n12943 , n14813 , n21243 );
    nor g9250 ( n8768 , n3248 , n21910 );
    or g9251 ( n28569 , n2022 , n924 );
    not g9252 ( n25715 , n11430 );
    or g9253 ( n35062 , n41428 , n13158 );
    not g9254 ( n17855 , n26095 );
    or g9255 ( n24413 , n37274 , n13710 );
    or g9256 ( n5913 , n4205 , n1940 );
    xnor g9257 ( n23996 , n35035 , n41238 );
    and g9258 ( n8721 , n29079 , n23287 );
    and g9259 ( n4956 , n41118 , n25159 );
    and g9260 ( n36902 , n16048 , n6793 );
    or g9261 ( n41765 , n30206 , n15232 );
    or g9262 ( n18791 , n10386 , n21365 );
    nor g9263 ( n13653 , n41761 , n29982 );
    nor g9264 ( n202 , n10716 , n20413 );
    or g9265 ( n36921 , n28490 , n8765 );
    or g9266 ( n33406 , n20854 , n29010 );
    nor g9267 ( n36347 , n9839 , n21271 );
    and g9268 ( n26036 , n11764 , n13379 );
    or g9269 ( n38634 , n832 , n18102 );
    not g9270 ( n4245 , n2369 );
    xnor g9271 ( n28860 , n14946 , n6682 );
    xnor g9272 ( n7620 , n15467 , n6524 );
    or g9273 ( n23643 , n22254 , n41176 );
    xnor g9274 ( n41232 , n35154 , n29521 );
    or g9275 ( n34180 , n5889 , n4660 );
    not g9276 ( n21837 , n23096 );
    or g9277 ( n34878 , n20040 , n4833 );
    nor g9278 ( n26219 , n33652 , n1320 );
    and g9279 ( n33954 , n10369 , n14071 );
    or g9280 ( n13583 , n28119 , n7949 );
    or g9281 ( n30339 , n12768 , n30128 );
    or g9282 ( n5860 , n23694 , n7995 );
    xnor g9283 ( n10200 , n31991 , n32277 );
    and g9284 ( n11641 , n2331 , n15760 );
    and g9285 ( n38063 , n23845 , n40123 );
    or g9286 ( n30052 , n10476 , n5813 );
    not g9287 ( n9916 , n36541 );
    nor g9288 ( n24125 , n28502 , n40943 );
    or g9289 ( n3239 , n22582 , n39468 );
    and g9290 ( n34315 , n24296 , n29810 );
    or g9291 ( n11621 , n36277 , n29550 );
    not g9292 ( n4852 , n13613 );
    and g9293 ( n27425 , n41805 , n17086 );
    nor g9294 ( n23101 , n27917 , n30627 );
    and g9295 ( n34911 , n39444 , n24568 );
    or g9296 ( n38745 , n6909 , n39520 );
    not g9297 ( n41981 , n9964 );
    nor g9298 ( n41570 , n8494 , n18522 );
    or g9299 ( n9723 , n14291 , n13085 );
    xnor g9300 ( n37860 , n11633 , n12690 );
    and g9301 ( n41287 , n21664 , n31602 );
    nor g9302 ( n8738 , n40666 , n77 );
    or g9303 ( n14358 , n12286 , n22683 );
    or g9304 ( n9650 , n21703 , n37519 );
    or g9305 ( n39451 , n32326 , n25243 );
    and g9306 ( n18078 , n34901 , n40103 );
    not g9307 ( n5574 , n15148 );
    and g9308 ( n17488 , n3609 , n25344 );
    nor g9309 ( n14433 , n35568 , n11329 );
    or g9310 ( n22252 , n40703 , n30767 );
    or g9311 ( n36673 , n11322 , n31707 );
    and g9312 ( n40116 , n22238 , n15660 );
    nor g9313 ( n6075 , n38391 , n41127 );
    nor g9314 ( n23162 , n17836 , n35085 );
    nor g9315 ( n15303 , n42699 , n33569 );
    or g9316 ( n37151 , n18601 , n21277 );
    and g9317 ( n21870 , n18901 , n1877 );
    or g9318 ( n18277 , n8244 , n2451 );
    not g9319 ( n13681 , n14301 );
    and g9320 ( n7267 , n4528 , n36204 );
    or g9321 ( n32021 , n3080 , n3414 );
    nor g9322 ( n30953 , n14840 , n35960 );
    or g9323 ( n25365 , n16469 , n29809 );
    or g9324 ( n39758 , n27503 , n31832 );
    xnor g9325 ( n39198 , n2799 , n10130 );
    not g9326 ( n12874 , n23848 );
    not g9327 ( n23598 , n25700 );
    and g9328 ( n11950 , n20456 , n5446 );
    xnor g9329 ( n39796 , n29740 , n21488 );
    nor g9330 ( n33102 , n3437 , n20436 );
    not g9331 ( n31539 , n38828 );
    and g9332 ( n15430 , n1469 , n26665 );
    or g9333 ( n39706 , n25522 , n35531 );
    and g9334 ( n35930 , n37570 , n41952 );
    not g9335 ( n5763 , n35882 );
    xnor g9336 ( n11131 , n40 , n6874 );
    not g9337 ( n16817 , n3925 );
    not g9338 ( n41698 , n166 );
    xnor g9339 ( n36126 , n7904 , n35249 );
    and g9340 ( n12477 , n34899 , n35312 );
    and g9341 ( n41249 , n11706 , n39129 );
    xnor g9342 ( n41970 , n22263 , n42913 );
    and g9343 ( n7030 , n9140 , n29397 );
    and g9344 ( n1999 , n25081 , n39518 );
    or g9345 ( n13365 , n4809 , n10710 );
    nor g9346 ( n355 , n27745 , n19224 );
    not g9347 ( n1301 , n8232 );
    or g9348 ( n39736 , n40764 , n20842 );
    nor g9349 ( n32117 , n36684 , n28355 );
    and g9350 ( n31412 , n39161 , n7036 );
    not g9351 ( n22746 , n28770 );
    or g9352 ( n21572 , n19723 , n21064 );
    and g9353 ( n2039 , n23343 , n34176 );
    xnor g9354 ( n24135 , n12146 , n19359 );
    or g9355 ( n9069 , n24615 , n40340 );
    xnor g9356 ( n15102 , n784 , n17187 );
    and g9357 ( n13712 , n24707 , n7311 );
    and g9358 ( n16890 , n1541 , n11011 );
    or g9359 ( n26849 , n7063 , n14457 );
    xnor g9360 ( n13353 , n527 , n4593 );
    or g9361 ( n30574 , n29612 , n2936 );
    or g9362 ( n29439 , n10778 , n8048 );
    and g9363 ( n22020 , n26054 , n31893 );
    and g9364 ( n17176 , n11115 , n32677 );
    nor g9365 ( n7364 , n9480 , n26998 );
    or g9366 ( n35891 , n12782 , n10106 );
    xnor g9367 ( n23804 , n5144 , n315 );
    not g9368 ( n37029 , n18138 );
    not g9369 ( n20304 , n23635 );
    not g9370 ( n24917 , n18583 );
    and g9371 ( n27126 , n27588 , n39163 );
    xnor g9372 ( n10815 , n32218 , n37097 );
    or g9373 ( n27975 , n25346 , n2877 );
    and g9374 ( n32686 , n11636 , n39278 );
    or g9375 ( n5512 , n7864 , n39304 );
    or g9376 ( n32947 , n31806 , n25907 );
    or g9377 ( n41630 , n31717 , n3290 );
    not g9378 ( n26817 , n42273 );
    and g9379 ( n32038 , n1306 , n3585 );
    and g9380 ( n3280 , n34283 , n2163 );
    not g9381 ( n465 , n33639 );
    or g9382 ( n15652 , n13244 , n14053 );
    and g9383 ( n23924 , n31154 , n19999 );
    or g9384 ( n39360 , n13396 , n13215 );
    xnor g9385 ( n22572 , n26406 , n42691 );
    nor g9386 ( n34961 , n18866 , n5216 );
    or g9387 ( n1725 , n15200 , n34634 );
    and g9388 ( n16472 , n25256 , n10001 );
    and g9389 ( n25129 , n8392 , n2450 );
    and g9390 ( n33419 , n11730 , n18153 );
    nor g9391 ( n235 , n16063 , n18632 );
    and g9392 ( n42565 , n6540 , n9944 );
    nor g9393 ( n38933 , n5253 , n42043 );
    and g9394 ( n16631 , n36304 , n8919 );
    or g9395 ( n27868 , n644 , n35257 );
    or g9396 ( n8314 , n28080 , n26389 );
    not g9397 ( n21907 , n19178 );
    not g9398 ( n25727 , n10279 );
    or g9399 ( n41478 , n2419 , n4908 );
    or g9400 ( n34088 , n16163 , n15871 );
    xnor g9401 ( n10411 , n37074 , n3606 );
    and g9402 ( n40879 , n14742 , n20017 );
    nor g9403 ( n12641 , n33222 , n10430 );
    or g9404 ( n25549 , n20442 , n10570 );
    and g9405 ( n14853 , n42093 , n41613 );
    or g9406 ( n20053 , n14606 , n11619 );
    nor g9407 ( n31264 , n22057 , n20680 );
    or g9408 ( n7291 , n22039 , n33965 );
    xnor g9409 ( n2625 , n14953 , n24784 );
    nor g9410 ( n23221 , n32462 , n17484 );
    or g9411 ( n261 , n17120 , n17944 );
    xnor g9412 ( n2290 , n27767 , n28345 );
    or g9413 ( n26616 , n10430 , n28551 );
    not g9414 ( n37131 , n40141 );
    or g9415 ( n32925 , n12450 , n25818 );
    nor g9416 ( n29812 , n17120 , n22095 );
    nor g9417 ( n29490 , n25172 , n42704 );
    and g9418 ( n12538 , n27860 , n14916 );
    nor g9419 ( n28481 , n25639 , n18329 );
    not g9420 ( n34586 , n35611 );
    or g9421 ( n13827 , n22821 , n23496 );
    not g9422 ( n23266 , n3634 );
    or g9423 ( n23793 , n16586 , n31998 );
    xnor g9424 ( n35667 , n25258 , n36840 );
    and g9425 ( n25963 , n10175 , n9025 );
    nor g9426 ( n1509 , n17790 , n39006 );
    not g9427 ( n11426 , n2919 );
    not g9428 ( n33314 , n32824 );
    not g9429 ( n5140 , n8641 );
    nor g9430 ( n23552 , n1507 , n42476 );
    or g9431 ( n42233 , n8015 , n38096 );
    nor g9432 ( n14067 , n36579 , n40672 );
    or g9433 ( n27547 , n28065 , n24195 );
    nor g9434 ( n18342 , n24745 , n37380 );
    and g9435 ( n28935 , n7859 , n38839 );
    or g9436 ( n470 , n26971 , n5422 );
    or g9437 ( n1782 , n28292 , n42218 );
    nor g9438 ( n10633 , n35813 , n35981 );
    or g9439 ( n20488 , n30652 , n28448 );
    or g9440 ( n27321 , n19695 , n41977 );
    and g9441 ( n2538 , n14709 , n21908 );
    xnor g9442 ( n36547 , n10088 , n16637 );
    or g9443 ( n42050 , n32656 , n14902 );
    or g9444 ( n32314 , n8501 , n20501 );
    and g9445 ( n26876 , n3269 , n41866 );
    and g9446 ( n21539 , n39330 , n24506 );
    xnor g9447 ( n24075 , n35371 , n27440 );
    xnor g9448 ( n6367 , n20015 , n19707 );
    or g9449 ( n33078 , n22250 , n5910 );
    nor g9450 ( n13965 , n33981 , n8198 );
    not g9451 ( n37256 , n22344 );
    or g9452 ( n11358 , n21473 , n23250 );
    or g9453 ( n1373 , n4083 , n16891 );
    or g9454 ( n38202 , n31844 , n12037 );
    and g9455 ( n23790 , n21727 , n19492 );
    and g9456 ( n34638 , n14178 , n648 );
    or g9457 ( n21010 , n38157 , n30269 );
    nor g9458 ( n27969 , n19221 , n30067 );
    not g9459 ( n32795 , n19798 );
    and g9460 ( n39821 , n13986 , n29699 );
    or g9461 ( n23685 , n33134 , n20366 );
    nor g9462 ( n41501 , n14707 , n17037 );
    nor g9463 ( n14436 , n38328 , n31304 );
    or g9464 ( n6424 , n7150 , n41501 );
    or g9465 ( n16951 , n39635 , n30665 );
    nor g9466 ( n21641 , n16023 , n31396 );
    and g9467 ( n11539 , n37476 , n42313 );
    nor g9468 ( n10253 , n37149 , n16995 );
    or g9469 ( n26852 , n5044 , n425 );
    and g9470 ( n688 , n20487 , n26022 );
    and g9471 ( n8864 , n42647 , n5550 );
    xnor g9472 ( n1639 , n11531 , n21564 );
    nor g9473 ( n8183 , n5964 , n33468 );
    or g9474 ( n4044 , n11640 , n30223 );
    or g9475 ( n40083 , n31918 , n4631 );
    or g9476 ( n23571 , n17903 , n10073 );
    or g9477 ( n40027 , n33981 , n36568 );
    not g9478 ( n26620 , n27446 );
    and g9479 ( n27071 , n35652 , n8644 );
    xnor g9480 ( n40590 , n784 , n41783 );
    and g9481 ( n10398 , n25556 , n11207 );
    or g9482 ( n13933 , n31958 , n37824 );
    not g9483 ( n5938 , n11181 );
    nor g9484 ( n34779 , n24411 , n31765 );
    or g9485 ( n1010 , n12220 , n25813 );
    or g9486 ( n10729 , n34011 , n33755 );
    not g9487 ( n7566 , n24177 );
    and g9488 ( n33665 , n32590 , n40842 );
    not g9489 ( n20384 , n35569 );
    not g9490 ( n19293 , n25357 );
    xnor g9491 ( n36232 , n41013 , n39661 );
    nor g9492 ( n25500 , n12041 , n13445 );
    xnor g9493 ( n3739 , n31989 , n24801 );
    and g9494 ( n26809 , n22479 , n6977 );
    or g9495 ( n24214 , n10987 , n36669 );
    and g9496 ( n7275 , n15129 , n5740 );
    or g9497 ( n29263 , n15510 , n39804 );
    or g9498 ( n41673 , n14471 , n35273 );
    nor g9499 ( n33947 , n13697 , n9581 );
    or g9500 ( n4749 , n28424 , n11864 );
    xnor g9501 ( n8612 , n5457 , n33557 );
    or g9502 ( n11244 , n9888 , n969 );
    not g9503 ( n7210 , n3008 );
    and g9504 ( n38255 , n41506 , n42790 );
    or g9505 ( n1242 , n13456 , n12038 );
    and g9506 ( n2270 , n1458 , n35591 );
    nor g9507 ( n13441 , n5605 , n10733 );
    and g9508 ( n19325 , n12485 , n23543 );
    or g9509 ( n22267 , n3323 , n17453 );
    or g9510 ( n34431 , n25526 , n17164 );
    or g9511 ( n18276 , n3901 , n26845 );
    or g9512 ( n34501 , n39382 , n39293 );
    xnor g9513 ( n19034 , n6338 , n25947 );
    and g9514 ( n34406 , n11624 , n24290 );
    or g9515 ( n40369 , n8292 , n28641 );
    and g9516 ( n10250 , n26292 , n21086 );
    xnor g9517 ( n19558 , n5159 , n36191 );
    and g9518 ( n31343 , n18445 , n14942 );
    not g9519 ( n21466 , n3680 );
    nor g9520 ( n7351 , n34483 , n15547 );
    or g9521 ( n30918 , n8150 , n31271 );
    or g9522 ( n6304 , n3498 , n5813 );
    or g9523 ( n12732 , n33328 , n38384 );
    nor g9524 ( n27090 , n27762 , n41848 );
    not g9525 ( n30477 , n1818 );
    xnor g9526 ( n21490 , n18696 , n259 );
    xnor g9527 ( n12530 , n1309 , n14471 );
    not g9528 ( n6760 , n37873 );
    xnor g9529 ( n8655 , n21192 , n38424 );
    and g9530 ( n15738 , n11691 , n41579 );
    or g9531 ( n2937 , n34528 , n7616 );
    or g9532 ( n28285 , n40544 , n4191 );
    and g9533 ( n30483 , n15668 , n41291 );
    and g9534 ( n14120 , n18383 , n30705 );
    and g9535 ( n16929 , n6143 , n39797 );
    or g9536 ( n15182 , n15934 , n598 );
    and g9537 ( n28209 , n258 , n14147 );
    nor g9538 ( n11527 , n5896 , n23467 );
    or g9539 ( n28838 , n4140 , n31125 );
    or g9540 ( n9018 , n32711 , n932 );
    not g9541 ( n11503 , n13044 );
    not g9542 ( n27781 , n8081 );
    or g9543 ( n28242 , n24062 , n12592 );
    or g9544 ( n17018 , n17440 , n27951 );
    or g9545 ( n17308 , n7143 , n39732 );
    nor g9546 ( n14958 , n36112 , n35761 );
    or g9547 ( n21209 , n18051 , n8372 );
    not g9548 ( n39933 , n3716 );
    not g9549 ( n15561 , n17338 );
    and g9550 ( n25969 , n5088 , n3699 );
    or g9551 ( n39259 , n22631 , n5180 );
    xnor g9552 ( n32375 , n33885 , n19498 );
    and g9553 ( n1191 , n8741 , n28635 );
    or g9554 ( n7145 , n22130 , n8087 );
    or g9555 ( n8936 , n23297 , n28715 );
    xnor g9556 ( n16308 , n25917 , n26924 );
    or g9557 ( n3952 , n20787 , n17576 );
    or g9558 ( n11416 , n16104 , n20367 );
    or g9559 ( n14950 , n34939 , n21076 );
    or g9560 ( n8730 , n35633 , n38296 );
    not g9561 ( n14233 , n38125 );
    nor g9562 ( n2731 , n16493 , n30154 );
    and g9563 ( n770 , n10403 , n31521 );
    not g9564 ( n36979 , n33108 );
    or g9565 ( n37035 , n34515 , n27385 );
    or g9566 ( n18721 , n27297 , n12198 );
    not g9567 ( n38532 , n36124 );
    or g9568 ( n26180 , n31679 , n29930 );
    not g9569 ( n30931 , n32427 );
    and g9570 ( n26982 , n30545 , n21601 );
    not g9571 ( n34151 , n23541 );
    xnor g9572 ( n18158 , n27658 , n42418 );
    or g9573 ( n913 , n6560 , n4323 );
    and g9574 ( n12607 , n22028 , n5439 );
    and g9575 ( n16759 , n1297 , n6680 );
    or g9576 ( n22466 , n11891 , n35758 );
    xnor g9577 ( n2554 , n4024 , n7104 );
    and g9578 ( n21875 , n21138 , n28830 );
    or g9579 ( n30746 , n33120 , n37141 );
    or g9580 ( n15097 , n26646 , n27196 );
    or g9581 ( n16053 , n39635 , n20514 );
    xnor g9582 ( n12440 , n302 , n6118 );
    or g9583 ( n37973 , n5307 , n34569 );
    nor g9584 ( n42651 , n23363 , n16070 );
    nor g9585 ( n13725 , n31242 , n23136 );
    not g9586 ( n19298 , n30406 );
    not g9587 ( n37983 , n17632 );
    or g9588 ( n29040 , n25471 , n26657 );
    or g9589 ( n4285 , n22298 , n69 );
    or g9590 ( n36455 , n14558 , n29322 );
    or g9591 ( n24949 , n33297 , n4310 );
    xnor g9592 ( n24266 , n37335 , n40665 );
    or g9593 ( n40392 , n33330 , n6013 );
    nor g9594 ( n13209 , n3581 , n16682 );
    and g9595 ( n28729 , n28616 , n39377 );
    or g9596 ( n7419 , n35320 , n1318 );
    not g9597 ( n31242 , n22121 );
    or g9598 ( n26449 , n14471 , n8479 );
    not g9599 ( n341 , n28202 );
    nor g9600 ( n27916 , n33222 , n42408 );
    or g9601 ( n38978 , n5964 , n38222 );
    not g9602 ( n7414 , n33362 );
    nor g9603 ( n17296 , n11702 , n31254 );
    xnor g9604 ( n34382 , n11449 , n26330 );
    or g9605 ( n11420 , n10803 , n17691 );
    or g9606 ( n18752 , n22750 , n5443 );
    or g9607 ( n32190 , n35514 , n24932 );
    not g9608 ( n34014 , n14042 );
    and g9609 ( n13580 , n39565 , n3651 );
    and g9610 ( n24349 , n30807 , n7133 );
    or g9611 ( n20852 , n6632 , n38894 );
    and g9612 ( n32215 , n16849 , n12164 );
    or g9613 ( n32045 , n10088 , n22868 );
    not g9614 ( n3834 , n26558 );
    not g9615 ( n22574 , n39487 );
    or g9616 ( n14878 , n15775 , n31544 );
    or g9617 ( n18306 , n26851 , n281 );
    not g9618 ( n18233 , n41484 );
    xnor g9619 ( n23960 , n2488 , n12559 );
    xnor g9620 ( n25525 , n11426 , n2322 );
    not g9621 ( n36355 , n25414 );
    or g9622 ( n31852 , n16365 , n30247 );
    nor g9623 ( n16331 , n34565 , n8374 );
    xnor g9624 ( n39222 , n25673 , n5831 );
    nor g9625 ( n38233 , n27927 , n24274 );
    and g9626 ( n28273 , n17965 , n18259 );
    xnor g9627 ( n6506 , n13683 , n10191 );
    xnor g9628 ( n27905 , n34731 , n34359 );
    or g9629 ( n34990 , n952 , n41015 );
    nor g9630 ( n41721 , n794 , n15822 );
    not g9631 ( n11001 , n15816 );
    and g9632 ( n33817 , n19167 , n26774 );
    xnor g9633 ( n24335 , n21954 , n5033 );
    nor g9634 ( n34465 , n16802 , n24759 );
    xnor g9635 ( n10954 , n36667 , n15952 );
    and g9636 ( n21068 , n6049 , n6934 );
    and g9637 ( n41914 , n30792 , n41469 );
    xnor g9638 ( n18968 , n36632 , n12310 );
    not g9639 ( n30473 , n22571 );
    and g9640 ( n41833 , n28677 , n39767 );
    not g9641 ( n4331 , n37839 );
    or g9642 ( n2557 , n10456 , n9390 );
    and g9643 ( n8301 , n7518 , n15345 );
    not g9644 ( n2840 , n8927 );
    not g9645 ( n8274 , n11713 );
    or g9646 ( n2294 , n12867 , n29778 );
    xnor g9647 ( n18444 , n19665 , n31720 );
    nor g9648 ( n1723 , n9629 , n39419 );
    and g9649 ( n42743 , n2996 , n37923 );
    not g9650 ( n39449 , n26941 );
    and g9651 ( n39445 , n15841 , n16712 );
    not g9652 ( n11682 , n4907 );
    or g9653 ( n2938 , n4843 , n17385 );
    nor g9654 ( n35043 , n1507 , n33462 );
    and g9655 ( n2607 , n15070 , n14260 );
    nor g9656 ( n17224 , n12311 , n23539 );
    or g9657 ( n10970 , n37018 , n33137 );
    not g9658 ( n22456 , n14975 );
    and g9659 ( n12818 , n35448 , n30952 );
    xnor g9660 ( n20783 , n18530 , n35736 );
    or g9661 ( n38195 , n21978 , n30680 );
    and g9662 ( n5323 , n41733 , n38360 );
    or g9663 ( n35750 , n31644 , n5941 );
    nor g9664 ( n8853 , n5459 , n22205 );
    or g9665 ( n24741 , n13255 , n35382 );
    or g9666 ( n9956 , n34596 , n485 );
    and g9667 ( n5403 , n18982 , n42175 );
    nor g9668 ( n6296 , n38084 , n7547 );
    xnor g9669 ( n10412 , n21534 , n24286 );
    nor g9670 ( n26606 , n5896 , n8363 );
    and g9671 ( n13223 , n14127 , n3171 );
    and g9672 ( n3975 , n31778 , n17773 );
    not g9673 ( n22790 , n16801 );
    or g9674 ( n30426 , n36535 , n14955 );
    xnor g9675 ( n12728 , n31992 , n10788 );
    or g9676 ( n29468 , n4355 , n33577 );
    or g9677 ( n41948 , n5673 , n13529 );
    or g9678 ( n14865 , n20830 , n20184 );
    not g9679 ( n3487 , n2062 );
    or g9680 ( n8723 , n28837 , n24743 );
    or g9681 ( n33673 , n38373 , n21268 );
    xnor g9682 ( n6020 , n14739 , n42789 );
    not g9683 ( n23583 , n27817 );
    and g9684 ( n42180 , n20524 , n36698 );
    or g9685 ( n21099 , n18866 , n33486 );
    nor g9686 ( n23307 , n8494 , n930 );
    not g9687 ( n3137 , n280 );
    or g9688 ( n42208 , n16161 , n39515 );
    or g9689 ( n3156 , n21807 , n13067 );
    not g9690 ( n40792 , n27687 );
    not g9691 ( n11813 , n20334 );
    or g9692 ( n3011 , n13176 , n33878 );
    nor g9693 ( n39580 , n12264 , n28732 );
    or g9694 ( n20347 , n12105 , n37957 );
    or g9695 ( n24586 , n14707 , n20424 );
    or g9696 ( n6746 , n5348 , n24349 );
    not g9697 ( n11417 , n13759 );
    or g9698 ( n33021 , n25228 , n35713 );
    or g9699 ( n29672 , n27359 , n25528 );
    not g9700 ( n35058 , n37485 );
    and g9701 ( n3736 , n4930 , n28776 );
    or g9702 ( n7805 , n23703 , n5900 );
    or g9703 ( n33622 , n11272 , n971 );
    or g9704 ( n30709 , n22821 , n19404 );
    xnor g9705 ( n39263 , n11785 , n17574 );
    or g9706 ( n30907 , n26542 , n41927 );
    nor g9707 ( n4050 , n39174 , n11820 );
    and g9708 ( n25288 , n4643 , n39010 );
    or g9709 ( n28365 , n24621 , n36528 );
    or g9710 ( n39917 , n36549 , n24367 );
    and g9711 ( n20759 , n31549 , n23843 );
    not g9712 ( n17225 , n3759 );
    or g9713 ( n15826 , n7758 , n12480 );
    not g9714 ( n37771 , n13668 );
    not g9715 ( n41903 , n20870 );
    or g9716 ( n20257 , n36296 , n207 );
    nor g9717 ( n12374 , n36053 , n18160 );
    or g9718 ( n3161 , n26935 , n20406 );
    xnor g9719 ( n24579 , n16693 , n15718 );
    xnor g9720 ( n33519 , n21765 , n5770 );
    and g9721 ( n11601 , n2118 , n1131 );
    or g9722 ( n38286 , n31145 , n29396 );
    or g9723 ( n32531 , n7414 , n30155 );
    and g9724 ( n25011 , n37067 , n23460 );
    not g9725 ( n30832 , n40927 );
    xnor g9726 ( n27520 , n16320 , n19858 );
    xnor g9727 ( n17315 , n1216 , n11797 );
    xnor g9728 ( n26496 , n13444 , n41581 );
    and g9729 ( n29774 , n32696 , n2361 );
    not g9730 ( n38214 , n27052 );
    nor g9731 ( n27357 , n38058 , n26820 );
    xnor g9732 ( n23267 , n28648 , n41425 );
    and g9733 ( n5278 , n30773 , n37532 );
    xnor g9734 ( n2400 , n13046 , n8526 );
    and g9735 ( n41700 , n1398 , n10978 );
    or g9736 ( n23414 , n3748 , n31618 );
    or g9737 ( n41168 , n28904 , n30616 );
    xnor g9738 ( n24410 , n18874 , n2765 );
    and g9739 ( n40449 , n7089 , n66 );
    and g9740 ( n29020 , n37375 , n6137 );
    not g9741 ( n29305 , n39738 );
    or g9742 ( n13240 , n18335 , n29757 );
    and g9743 ( n19503 , n2494 , n20693 );
    and g9744 ( n12166 , n4945 , n24109 );
    nor g9745 ( n20941 , n3839 , n25274 );
    and g9746 ( n27508 , n25511 , n40548 );
    and g9747 ( n21218 , n5304 , n14435 );
    and g9748 ( n34319 , n29886 , n18136 );
    and g9749 ( n19698 , n4516 , n16059 );
    or g9750 ( n32682 , n40865 , n29608 );
    and g9751 ( n25583 , n22700 , n18780 );
    and g9752 ( n6966 , n32850 , n20377 );
    xnor g9753 ( n28537 , n15860 , n11890 );
    or g9754 ( n41096 , n12490 , n29218 );
    nor g9755 ( n33820 , n26763 , n34971 );
    or g9756 ( n7776 , n7475 , n14103 );
    not g9757 ( n1978 , n35923 );
    and g9758 ( n37849 , n39013 , n4534 );
    or g9759 ( n37877 , n23762 , n40612 );
    and g9760 ( n12465 , n15755 , n14936 );
    and g9761 ( n6180 , n19833 , n30500 );
    not g9762 ( n17100 , n9062 );
    and g9763 ( n41314 , n19550 , n23638 );
    or g9764 ( n30645 , n33981 , n35823 );
    nor g9765 ( n30213 , n26921 , n24319 );
    nor g9766 ( n14427 , n4470 , n15642 );
    xnor g9767 ( n17095 , n12146 , n24400 );
    or g9768 ( n577 , n3801 , n22671 );
    or g9769 ( n38709 , n27432 , n8171 );
    nor g9770 ( n22524 , n32953 , n8629 );
    or g9771 ( n18397 , n26915 , n16798 );
    not g9772 ( n19419 , n32560 );
    nor g9773 ( n32064 , n17744 , n38213 );
    or g9774 ( n5792 , n26076 , n41608 );
    xnor g9775 ( n11283 , n8994 , n38879 );
    and g9776 ( n40766 , n29471 , n6375 );
    not g9777 ( n32048 , n36309 );
    or g9778 ( n38030 , n34060 , n11369 );
    or g9779 ( n39855 , n32711 , n14982 );
    or g9780 ( n30377 , n30519 , n40989 );
    or g9781 ( n34018 , n18376 , n12055 );
    and g9782 ( n4952 , n34800 , n40095 );
    or g9783 ( n19663 , n33464 , n28514 );
    or g9784 ( n20057 , n10598 , n1290 );
    or g9785 ( n9224 , n32124 , n6197 );
    or g9786 ( n16639 , n34686 , n29888 );
    not g9787 ( n36255 , n19724 );
    or g9788 ( n16290 , n6559 , n10754 );
    xnor g9789 ( n29684 , n35553 , n4006 );
    nor g9790 ( n24923 , n26394 , n15421 );
    and g9791 ( n17139 , n36871 , n36146 );
    or g9792 ( n28107 , n38704 , n14141 );
    xnor g9793 ( n38989 , n18530 , n9 );
    nor g9794 ( n36199 , n21979 , n30364 );
    or g9795 ( n6921 , n7388 , n37806 );
    xnor g9796 ( n8842 , n31989 , n18485 );
    nor g9797 ( n21041 , n10822 , n4688 );
    nor g9798 ( n16082 , n36104 , n18893 );
    not g9799 ( n7056 , n21270 );
    or g9800 ( n23223 , n1613 , n32820 );
    nor g9801 ( n4658 , n15288 , n36732 );
    and g9802 ( n6453 , n20892 , n17708 );
    or g9803 ( n5272 , n3747 , n5682 );
    or g9804 ( n27944 , n23082 , n5852 );
    or g9805 ( n4471 , n21553 , n28291 );
    or g9806 ( n19454 , n15968 , n27884 );
    nor g9807 ( n10490 , n13041 , n28969 );
    not g9808 ( n32983 , n33631 );
    nor g9809 ( n20401 , n20817 , n37690 );
    xnor g9810 ( n10034 , n21888 , n32027 );
    and g9811 ( n19035 , n7943 , n37378 );
    or g9812 ( n2504 , n40794 , n8455 );
    and g9813 ( n14063 , n31639 , n10764 );
    not g9814 ( n20446 , n36025 );
    or g9815 ( n13666 , n25588 , n30152 );
    nor g9816 ( n11854 , n6145 , n25146 );
    and g9817 ( n33228 , n36589 , n41167 );
    or g9818 ( n4019 , n42352 , n26788 );
    xnor g9819 ( n21190 , n11595 , n35153 );
    not g9820 ( n26377 , n6260 );
    or g9821 ( n28355 , n34748 , n1409 );
    nor g9822 ( n40652 , n2441 , n42474 );
    and g9823 ( n4617 , n22311 , n25766 );
    xnor g9824 ( n13932 , n42064 , n23426 );
    not g9825 ( n28882 , n31010 );
    nor g9826 ( n18515 , n31208 , n35983 );
    or g9827 ( n23257 , n22872 , n39083 );
    or g9828 ( n29373 , n41684 , n4737 );
    xnor g9829 ( n39858 , n34731 , n9837 );
    and g9830 ( n34320 , n29416 , n709 );
    xnor g9831 ( n34884 , n13597 , n35636 );
    or g9832 ( n23333 , n26133 , n8940 );
    not g9833 ( n4375 , n33883 );
    xnor g9834 ( n40964 , n28979 , n14873 );
    and g9835 ( n41131 , n23613 , n1284 );
    or g9836 ( n39893 , n42405 , n8865 );
    and g9837 ( n13883 , n28519 , n13241 );
    or g9838 ( n32496 , n16717 , n19809 );
    or g9839 ( n21181 , n30188 , n27586 );
    or g9840 ( n13110 , n4045 , n20877 );
    xnor g9841 ( n1467 , n10612 , n12744 );
    or g9842 ( n28240 , n14471 , n1039 );
    nor g9843 ( n10248 , n24509 , n17890 );
    or g9844 ( n15363 , n14707 , n27161 );
    xnor g9845 ( n8110 , n31099 , n15688 );
    nor g9846 ( n6691 , n41195 , n19263 );
    not g9847 ( n22611 , n7268 );
    or g9848 ( n28703 , n28020 , n33637 );
    or g9849 ( n12447 , n6019 , n13331 );
    and g9850 ( n39201 , n693 , n18562 );
    xnor g9851 ( n473 , n20487 , n475 );
    and g9852 ( n19068 , n16697 , n19157 );
    or g9853 ( n11399 , n3525 , n7375 );
    and g9854 ( n748 , n15225 , n35393 );
    or g9855 ( n11002 , n1626 , n38509 );
    not g9856 ( n7628 , n40225 );
    or g9857 ( n35324 , n23553 , n28241 );
    or g9858 ( n13808 , n35963 , n13347 );
    or g9859 ( n13976 , n34060 , n14220 );
    xnor g9860 ( n4836 , n4972 , n37809 );
    not g9861 ( n33013 , n35062 );
    or g9862 ( n36850 , n1574 , n15573 );
    not g9863 ( n41805 , n26706 );
    xnor g9864 ( n28584 , n965 , n40577 );
    or g9865 ( n29014 , n7839 , n12559 );
    or g9866 ( n23978 , n16109 , n21782 );
    nor g9867 ( n14374 , n18424 , n33128 );
    xnor g9868 ( n10293 , n10558 , n15907 );
    or g9869 ( n419 , n9031 , n6181 );
    nor g9870 ( n35757 , n13749 , n10056 );
    xnor g9871 ( n35353 , n5144 , n1334 );
    not g9872 ( n4228 , n28530 );
    and g9873 ( n4716 , n13217 , n40435 );
    nor g9874 ( n17472 , n4556 , n18262 );
    nor g9875 ( n22467 , n37771 , n28222 );
    not g9876 ( n14819 , n25800 );
    and g9877 ( n33173 , n941 , n2724 );
    and g9878 ( n2007 , n39556 , n24406 );
    and g9879 ( n39 , n13195 , n3533 );
    and g9880 ( n1177 , n5112 , n23661 );
    or g9881 ( n39329 , n35289 , n27383 );
    xnor g9882 ( n33444 , n18530 , n23757 );
    or g9883 ( n24769 , n25053 , n20801 );
    nor g9884 ( n17783 , n15221 , n31234 );
    or g9885 ( n34442 , n35515 , n34184 );
    and g9886 ( n25623 , n27415 , n33244 );
    and g9887 ( n24704 , n28068 , n33934 );
    or g9888 ( n22621 , n31060 , n41333 );
    or g9889 ( n2331 , n15269 , n29212 );
    or g9890 ( n9220 , n825 , n35 );
    or g9891 ( n21346 , n37651 , n12598 );
    or g9892 ( n18776 , n35883 , n25144 );
    xnor g9893 ( n23883 , n11023 , n39663 );
    or g9894 ( n27255 , n7223 , n17129 );
    and g9895 ( n17190 , n32197 , n2504 );
    nor g9896 ( n32754 , n39028 , n18626 );
    or g9897 ( n35958 , n15271 , n34960 );
    nor g9898 ( n7413 , n41534 , n1993 );
    and g9899 ( n36023 , n11726 , n14043 );
    xnor g9900 ( n30874 , n24278 , n37703 );
    or g9901 ( n41918 , n17194 , n28500 );
    and g9902 ( n35662 , n33325 , n5858 );
    or g9903 ( n16203 , n41097 , n29930 );
    not g9904 ( n27473 , n31337 );
    and g9905 ( n2132 , n28435 , n580 );
    xnor g9906 ( n19418 , n34945 , n6105 );
    or g9907 ( n12443 , n28173 , n17703 );
    not g9908 ( n36275 , n31287 );
    or g9909 ( n14190 , n16890 , n38810 );
    or g9910 ( n22992 , n9376 , n1279 );
    not g9911 ( n40957 , n20841 );
    and g9912 ( n2979 , n21343 , n5888 );
    or g9913 ( n19021 , n14531 , n41950 );
    xnor g9914 ( n40836 , n4467 , n22671 );
    xnor g9915 ( n29685 , n1629 , n4761 );
    not g9916 ( n33679 , n29694 );
    nor g9917 ( n13222 , n16221 , n10452 );
    not g9918 ( n38263 , n21183 );
    not g9919 ( n28614 , n13111 );
    nor g9920 ( n16190 , n26952 , n29205 );
    nor g9921 ( n39164 , n349 , n13995 );
    and g9922 ( n31072 , n39961 , n31604 );
    xnor g9923 ( n18947 , n16884 , n35762 );
    not g9924 ( n25994 , n22980 );
    or g9925 ( n31798 , n3545 , n39064 );
    or g9926 ( n20967 , n16696 , n20925 );
    nor g9927 ( n377 , n38835 , n1829 );
    and g9928 ( n19170 , n22453 , n15805 );
    or g9929 ( n20989 , n1583 , n7321 );
    and g9930 ( n42816 , n32620 , n5689 );
    nor g9931 ( n42183 , n9777 , n20114 );
    or g9932 ( n13973 , n37629 , n34911 );
    xnor g9933 ( n5030 , n542 , n23779 );
    or g9934 ( n19128 , n19486 , n8494 );
    or g9935 ( n24040 , n31387 , n42220 );
    not g9936 ( n20792 , n19614 );
    not g9937 ( n36009 , n1507 );
    or g9938 ( n2423 , n36413 , n1215 );
    or g9939 ( n39421 , n19102 , n22606 );
    xnor g9940 ( n25231 , n28225 , n30895 );
    or g9941 ( n11127 , n32478 , n1099 );
    or g9942 ( n9183 , n23971 , n3024 );
    xnor g9943 ( n8047 , n30189 , n20865 );
    not g9944 ( n20030 , n29731 );
    nor g9945 ( n733 , n5182 , n11358 );
    not g9946 ( n5457 , n27148 );
    or g9947 ( n2610 , n27928 , n5261 );
    xnor g9948 ( n41764 , n2339 , n14223 );
    or g9949 ( n23664 , n22642 , n40997 );
    or g9950 ( n3708 , n28456 , n6512 );
    and g9951 ( n41361 , n2823 , n41701 );
    and g9952 ( n30665 , n31449 , n15234 );
    not g9953 ( n41288 , n35450 );
    or g9954 ( n26083 , n7637 , n19706 );
    nor g9955 ( n23803 , n34611 , n34840 );
    or g9956 ( n33012 , n3571 , n34769 );
    xnor g9957 ( n19071 , n40 , n21817 );
    and g9958 ( n252 , n23034 , n11122 );
    or g9959 ( n1446 , n15625 , n37385 );
    nor g9960 ( n22739 , n33981 , n29065 );
    xnor g9961 ( n17391 , n42064 , n216 );
    and g9962 ( n23726 , n26678 , n21083 );
    or g9963 ( n24646 , n1752 , n15519 );
    or g9964 ( n8756 , n42792 , n17720 );
    not g9965 ( n9637 , n5337 );
    xnor g9966 ( n27560 , n22128 , n37182 );
    or g9967 ( n23677 , n14741 , n782 );
    and g9968 ( n14001 , n4349 , n2201 );
    and g9969 ( n36494 , n31598 , n41627 );
    or g9970 ( n31441 , n22427 , n29862 );
    xnor g9971 ( n17098 , n23947 , n12783 );
    not g9972 ( n794 , n2630 );
    xnor g9973 ( n10812 , n7904 , n40473 );
    and g9974 ( n27776 , n22449 , n21043 );
    nor g9975 ( n2225 , n26627 , n7482 );
    or g9976 ( n11060 , n11444 , n15158 );
    or g9977 ( n12884 , n28629 , n27884 );
    not g9978 ( n27899 , n34339 );
    and g9979 ( n36091 , n1746 , n34351 );
    xnor g9980 ( n5240 , n36998 , n41827 );
    nor g9981 ( n25911 , n33981 , n40947 );
    nor g9982 ( n11753 , n38168 , n13601 );
    not g9983 ( n12314 , n4646 );
    nor g9984 ( n7250 , n31610 , n20047 );
    nor g9985 ( n8960 , n19000 , n16234 );
    or g9986 ( n32685 , n33297 , n17355 );
    and g9987 ( n41374 , n4334 , n4971 );
    xnor g9988 ( n32376 , n5891 , n35332 );
    not g9989 ( n42851 , n29369 );
    and g9990 ( n1439 , n30054 , n40683 );
    and g9991 ( n40137 , n13476 , n23410 );
    and g9992 ( n10255 , n38952 , n38065 );
    nor g9993 ( n11025 , n16620 , n21695 );
    and g9994 ( n24901 , n12216 , n40783 );
    or g9995 ( n19109 , n17120 , n3254 );
    and g9996 ( n37564 , n42241 , n19710 );
    or g9997 ( n27299 , n3373 , n2021 );
    and g9998 ( n14861 , n23333 , n35102 );
    not g9999 ( n24058 , n42608 );
    nor g10000 ( n38813 , n26398 , n39353 );
    or g10001 ( n25 , n17744 , n11 );
    or g10002 ( n2824 , n2280 , n17404 );
    or g10003 ( n40416 , n3223 , n1527 );
    and g10004 ( n27624 , n23850 , n4182 );
    or g10005 ( n41933 , n32712 , n28457 );
    and g10006 ( n1874 , n16003 , n35246 );
    xnor g10007 ( n25641 , n36046 , n17919 );
    or g10008 ( n1652 , n32739 , n16220 );
    not g10009 ( n24892 , n8949 );
    not g10010 ( n29964 , n3704 );
    nor g10011 ( n39318 , n12250 , n36248 );
    or g10012 ( n30726 , n18777 , n42706 );
    and g10013 ( n23995 , n41272 , n32171 );
    nor g10014 ( n19134 , n35793 , n5655 );
    and g10015 ( n30097 , n41244 , n1236 );
    or g10016 ( n13297 , n34546 , n13885 );
    or g10017 ( n42576 , n37933 , n24503 );
    and g10018 ( n7297 , n11436 , n34644 );
    or g10019 ( n41234 , n15563 , n33976 );
    nor g10020 ( n22605 , n23234 , n18476 );
    or g10021 ( n39009 , n28349 , n1403 );
    not g10022 ( n14153 , n11047 );
    or g10023 ( n31425 , n14250 , n35116 );
    xnor g10024 ( n1055 , n41013 , n41732 );
    nor g10025 ( n31454 , n31228 , n39675 );
    not g10026 ( n3154 , n24616 );
    not g10027 ( n24328 , n21308 );
    and g10028 ( n38657 , n16640 , n34989 );
    nor g10029 ( n12938 , n2763 , n9569 );
    or g10030 ( n42259 , n14061 , n6271 );
    or g10031 ( n12404 , n25932 , n18771 );
    or g10032 ( n2336 , n4670 , n14035 );
    nor g10033 ( n135 , n18433 , n6194 );
    or g10034 ( n2788 , n5913 , n42119 );
    or g10035 ( n29827 , n32093 , n33118 );
    or g10036 ( n15712 , n23139 , n42125 );
    not g10037 ( n16999 , n25910 );
    nor g10038 ( n31730 , n41906 , n21193 );
    or g10039 ( n18463 , n27186 , n41990 );
    not g10040 ( n22036 , n29809 );
    and g10041 ( n12616 , n13768 , n28270 );
    not g10042 ( n42264 , n522 );
    or g10043 ( n20534 , n26264 , n5588 );
    or g10044 ( n3099 , n11149 , n19753 );
    xnor g10045 ( n3013 , n40 , n19971 );
    or g10046 ( n15357 , n16197 , n2492 );
    or g10047 ( n9666 , n42792 , n33527 );
    and g10048 ( n24801 , n28142 , n42362 );
    nor g10049 ( n31662 , n33283 , n5672 );
    or g10050 ( n18092 , n41860 , n23262 );
    or g10051 ( n4597 , n20025 , n24534 );
    or g10052 ( n41486 , n22396 , n22968 );
    and g10053 ( n37419 , n21209 , n3460 );
    nor g10054 ( n10365 , n10427 , n32719 );
    or g10055 ( n1162 , n38216 , n41413 );
    and g10056 ( n27355 , n11999 , n11505 );
    nor g10057 ( n6948 , n41773 , n15062 );
    xnor g10058 ( n42360 , n24165 , n31591 );
    or g10059 ( n12324 , n10582 , n18070 );
    and g10060 ( n39791 , n14965 , n14031 );
    xnor g10061 ( n39763 , n34731 , n37891 );
    not g10062 ( n14056 , n28499 );
    xnor g10063 ( n14993 , n22263 , n18428 );
    or g10064 ( n194 , n41433 , n16929 );
    xnor g10065 ( n19033 , n22263 , n28633 );
    and g10066 ( n21024 , n4983 , n32505 );
    xnor g10067 ( n208 , n15051 , n38816 );
    and g10068 ( n3020 , n7228 , n36450 );
    or g10069 ( n3958 , n14707 , n14868 );
    not g10070 ( n2832 , n24956 );
    xnor g10071 ( n31947 , n30768 , n3230 );
    xnor g10072 ( n4437 , n22346 , n832 );
    nor g10073 ( n257 , n19907 , n16152 );
    and g10074 ( n28109 , n35451 , n21122 );
    and g10075 ( n20390 , n36206 , n18284 );
    or g10076 ( n3733 , n11722 , n6792 );
    or g10077 ( n5811 , n4502 , n1667 );
    not g10078 ( n17467 , n4587 );
    or g10079 ( n32360 , n30412 , n25784 );
    or g10080 ( n5519 , n1635 , n31238 );
    not g10081 ( n10716 , n6054 );
    nor g10082 ( n15264 , n11563 , n19199 );
    and g10083 ( n40987 , n3426 , n35873 );
    or g10084 ( n33063 , n32390 , n39883 );
    or g10085 ( n22916 , n9300 , n37186 );
    not g10086 ( n5447 , n8361 );
    xnor g10087 ( n37546 , n37176 , n11949 );
    or g10088 ( n37810 , n13551 , n16759 );
    not g10089 ( n16397 , n18142 );
    or g10090 ( n30023 , n12728 , n39992 );
    not g10091 ( n5324 , n17918 );
    or g10092 ( n1613 , n13821 , n439 );
    or g10093 ( n10684 , n24656 , n8454 );
    and g10094 ( n29173 , n11686 , n13494 );
    or g10095 ( n15100 , n34378 , n38981 );
    nor g10096 ( n33074 , n26904 , n31680 );
    and g10097 ( n41678 , n20669 , n8376 );
    or g10098 ( n41983 , n28066 , n684 );
    or g10099 ( n11751 , n34626 , n30326 );
    nor g10100 ( n35541 , n36667 , n34430 );
    or g10101 ( n17761 , n3557 , n36326 );
    nor g10102 ( n22468 , n35711 , n36518 );
    and g10103 ( n2077 , n7472 , n35244 );
    and g10104 ( n23254 , n38337 , n11400 );
    nor g10105 ( n24775 , n383 , n10521 );
    or g10106 ( n23458 , n18115 , n16260 );
    not g10107 ( n26493 , n12969 );
    xnor g10108 ( n12917 , n30022 , n5357 );
    and g10109 ( n11617 , n18681 , n33371 );
    not g10110 ( n28577 , n41841 );
    nor g10111 ( n33467 , n18914 , n12925 );
    nor g10112 ( n15364 , n8494 , n25614 );
    or g10113 ( n42350 , n25551 , n42831 );
    or g10114 ( n42756 , n26961 , n869 );
    or g10115 ( n23723 , n21082 , n18104 );
    not g10116 ( n36932 , n25207 );
    not g10117 ( n2659 , n12224 );
    nor g10118 ( n38645 , n20227 , n3031 );
    not g10119 ( n28263 , n15412 );
    not g10120 ( n31780 , n3101 );
    not g10121 ( n21965 , n19233 );
    xnor g10122 ( n12304 , n174 , n27910 );
    nor g10123 ( n31844 , n17823 , n10121 );
    xnor g10124 ( n32563 , n16717 , n4356 );
    nor g10125 ( n12612 , n5605 , n42225 );
    not g10126 ( n14658 , n8759 );
    or g10127 ( n63 , n9409 , n10899 );
    or g10128 ( n31316 , n19366 , n40495 );
    or g10129 ( n38871 , n28226 , n40271 );
    or g10130 ( n10838 , n28634 , n40984 );
    and g10131 ( n14491 , n36390 , n13169 );
    nor g10132 ( n19549 , n24064 , n22589 );
    or g10133 ( n29836 , n22171 , n3157 );
    xnor g10134 ( n34012 , n34731 , n12298 );
    or g10135 ( n34776 , n10090 , n1344 );
    or g10136 ( n28477 , n21847 , n22129 );
    not g10137 ( n20726 , n25123 );
    and g10138 ( n39822 , n30161 , n42162 );
    not g10139 ( n40015 , n38046 );
    and g10140 ( n29023 , n32647 , n13778 );
    not g10141 ( n18937 , n37770 );
    and g10142 ( n38216 , n12538 , n14012 );
    or g10143 ( n35702 , n37763 , n24897 );
    not g10144 ( n40764 , n13641 );
    not g10145 ( n14944 , n25288 );
    not g10146 ( n15280 , n41688 );
    or g10147 ( n33525 , n6636 , n9435 );
    or g10148 ( n16352 , n33054 , n26101 );
    or g10149 ( n406 , n24068 , n6299 );
    xnor g10150 ( n22922 , n18530 , n8891 );
    xnor g10151 ( n2957 , n18146 , n4654 );
    or g10152 ( n39767 , n22705 , n11504 );
    or g10153 ( n34464 , n29221 , n1054 );
    or g10154 ( n7326 , n29803 , n4489 );
    or g10155 ( n14429 , n39608 , n28831 );
    or g10156 ( n38366 , n3518 , n1735 );
    and g10157 ( n28013 , n3299 , n16946 );
    or g10158 ( n17546 , n10939 , n26588 );
    not g10159 ( n1457 , n9062 );
    or g10160 ( n16634 , n12112 , n14860 );
    and g10161 ( n10685 , n5160 , n15249 );
    not g10162 ( n13316 , n9389 );
    or g10163 ( n26566 , n17053 , n32604 );
    nor g10164 ( n1511 , n27658 , n3818 );
    not g10165 ( n7920 , n41200 );
    or g10166 ( n4458 , n9720 , n5545 );
    nor g10167 ( n19652 , n15102 , n5569 );
    and g10168 ( n8973 , n6877 , n17439 );
    xnor g10169 ( n19007 , n10601 , n24484 );
    or g10170 ( n18737 , n20772 , n34225 );
    not g10171 ( n6000 , n36110 );
    or g10172 ( n14994 , n14361 , n2193 );
    nor g10173 ( n39395 , n1338 , n40675 );
    nor g10174 ( n12035 , n40247 , n18505 );
    or g10175 ( n39914 , n40427 , n11757 );
    not g10176 ( n27026 , n32384 );
    nor g10177 ( n30313 , n4265 , n39071 );
    and g10178 ( n9015 , n4677 , n11017 );
    xnor g10179 ( n25620 , n11596 , n21069 );
    or g10180 ( n14576 , n37656 , n25959 );
    nor g10181 ( n3257 , n35861 , n3873 );
    or g10182 ( n10167 , n26122 , n4187 );
    and g10183 ( n5863 , n22880 , n34950 );
    nor g10184 ( n3174 , n9001 , n23459 );
    and g10185 ( n27176 , n23379 , n21792 );
    or g10186 ( n35574 , n32358 , n8676 );
    xnor g10187 ( n39254 , n34401 , n19447 );
    nor g10188 ( n16393 , n17057 , n27954 );
    or g10189 ( n23429 , n36108 , n14811 );
    not g10190 ( n19120 , n36010 );
    or g10191 ( n41154 , n8916 , n31185 );
    and g10192 ( n40325 , n12328 , n25199 );
    or g10193 ( n18709 , n36992 , n37264 );
    and g10194 ( n17559 , n16943 , n26720 );
    nor g10195 ( n30888 , n2183 , n18777 );
    and g10196 ( n12336 , n32717 , n29083 );
    or g10197 ( n13575 , n12011 , n4883 );
    not g10198 ( n29754 , n38874 );
    and g10199 ( n23138 , n31283 , n25338 );
    or g10200 ( n12064 , n5935 , n25710 );
    nor g10201 ( n34790 , n38157 , n38799 );
    and g10202 ( n7086 , n23514 , n8815 );
    and g10203 ( n601 , n15040 , n10858 );
    xnor g10204 ( n36263 , n898 , n38123 );
    nor g10205 ( n9384 , n40086 , n20194 );
    and g10206 ( n5782 , n11692 , n14254 );
    xnor g10207 ( n4201 , n22604 , n29434 );
    xnor g10208 ( n2471 , n42567 , n27934 );
    or g10209 ( n35618 , n12187 , n36240 );
    or g10210 ( n29691 , n40752 , n38119 );
    and g10211 ( n34502 , n40441 , n17782 );
    nor g10212 ( n42226 , n6617 , n39403 );
    and g10213 ( n8145 , n1562 , n39564 );
    or g10214 ( n27085 , n7851 , n35337 );
    or g10215 ( n5366 , n34292 , n25798 );
    xnor g10216 ( n22193 , n35107 , n20291 );
    nor g10217 ( n14722 , n7535 , n16841 );
    and g10218 ( n8410 , n39926 , n9082 );
    not g10219 ( n13769 , n38752 );
    not g10220 ( n40409 , n7739 );
    nor g10221 ( n21670 , n38879 , n18181 );
    and g10222 ( n30603 , n10016 , n37989 );
    or g10223 ( n41465 , n10486 , n15927 );
    nor g10224 ( n23829 , n1002 , n3862 );
    not g10225 ( n36625 , n11677 );
    xnor g10226 ( n21865 , n5746 , n6607 );
    not g10227 ( n39883 , n18510 );
    xnor g10228 ( n23069 , n24745 , n28297 );
    and g10229 ( n30368 , n11884 , n23212 );
    or g10230 ( n13319 , n26260 , n42123 );
    or g10231 ( n19583 , n30020 , n15509 );
    and g10232 ( n8294 , n27870 , n34912 );
    not g10233 ( n2565 , n28269 );
    xnor g10234 ( n24096 , n15051 , n6718 );
    and g10235 ( n29958 , n38925 , n9077 );
    or g10236 ( n24293 , n4669 , n24271 );
    and g10237 ( n36832 , n36999 , n8461 );
    not g10238 ( n41236 , n3280 );
    or g10239 ( n4814 , n28777 , n14416 );
    not g10240 ( n35501 , n42039 );
    and g10241 ( n4222 , n4194 , n5591 );
    not g10242 ( n4833 , n30286 );
    or g10243 ( n10368 , n26302 , n19355 );
    and g10244 ( n818 , n7277 , n10644 );
    nor g10245 ( n22853 , n41241 , n21920 );
    or g10246 ( n41235 , n3668 , n28772 );
    and g10247 ( n16982 , n12143 , n19767 );
    nor g10248 ( n21815 , n9240 , n11389 );
    or g10249 ( n34265 , n32605 , n21362 );
    and g10250 ( n4599 , n33514 , n4739 );
    or g10251 ( n7642 , n228 , n2104 );
    not g10252 ( n27393 , n11937 );
    not g10253 ( n29475 , n3140 );
    and g10254 ( n5128 , n18067 , n5758 );
    or g10255 ( n31813 , n22577 , n17930 );
    and g10256 ( n19909 , n9759 , n2873 );
    not g10257 ( n3960 , n40330 );
    or g10258 ( n25691 , n25721 , n26930 );
    or g10259 ( n30996 , n20990 , n36500 );
    and g10260 ( n24738 , n2824 , n19941 );
    or g10261 ( n12608 , n33523 , n6576 );
    and g10262 ( n39342 , n22196 , n33601 );
    or g10263 ( n30299 , n5896 , n22373 );
    and g10264 ( n12403 , n19428 , n9039 );
    xnor g10265 ( n12401 , n26579 , n39849 );
    or g10266 ( n7592 , n14892 , n3542 );
    or g10267 ( n28878 , n14696 , n8086 );
    nor g10268 ( n24232 , n42430 , n33163 );
    and g10269 ( n16170 , n38782 , n18744 );
    not g10270 ( n22490 , n7215 );
    xnor g10271 ( n19834 , n4334 , n12505 );
    or g10272 ( n582 , n28841 , n3034 );
    nor g10273 ( n29952 , n28252 , n29772 );
    or g10274 ( n28886 , n22957 , n21893 );
    not g10275 ( n32420 , n60 );
    xnor g10276 ( n9626 , n16693 , n41561 );
    and g10277 ( n15907 , n12556 , n11335 );
    xnor g10278 ( n31314 , n6861 , n33497 );
    or g10279 ( n20159 , n40787 , n23015 );
    or g10280 ( n20981 , n1724 , n30019 );
    or g10281 ( n29779 , n40773 , n2108 );
    or g10282 ( n13096 , n8083 , n37434 );
    not g10283 ( n11981 , n4628 );
    and g10284 ( n16684 , n30817 , n34724 );
    and g10285 ( n28869 , n33346 , n41510 );
    xnor g10286 ( n1029 , n25701 , n11968 );
    or g10287 ( n9026 , n1149 , n24783 );
    nor g10288 ( n36139 , n9882 , n20154 );
    or g10289 ( n21896 , n32515 , n37128 );
    xnor g10290 ( n13649 , n4538 , n3630 );
    xnor g10291 ( n19806 , n34236 , n38705 );
    or g10292 ( n8368 , n28634 , n15973 );
    not g10293 ( n32824 , n2562 );
    and g10294 ( n25223 , n41737 , n4487 );
    not g10295 ( n3014 , n3087 );
    or g10296 ( n38987 , n5896 , n25367 );
    and g10297 ( n9459 , n20255 , n37313 );
    or g10298 ( n24660 , n15729 , n2565 );
    nor g10299 ( n41009 , n32542 , n23655 );
    xnor g10300 ( n7077 , n329 , n13125 );
    or g10301 ( n21489 , n38995 , n14583 );
    or g10302 ( n4142 , n7370 , n5138 );
    or g10303 ( n21315 , n12754 , n31439 );
    or g10304 ( n16177 , n30030 , n38544 );
    nor g10305 ( n25956 , n24551 , n36627 );
    and g10306 ( n2315 , n6514 , n3063 );
    nor g10307 ( n37785 , n12381 , n889 );
    nor g10308 ( n11328 , n12837 , n27468 );
    and g10309 ( n41863 , n31409 , n23866 );
    or g10310 ( n32769 , n591 , n21855 );
    xnor g10311 ( n10386 , n9275 , n4564 );
    or g10312 ( n26124 , n31791 , n34817 );
    and g10313 ( n14299 , n32833 , n16432 );
    or g10314 ( n37310 , n15339 , n28309 );
    not g10315 ( n38035 , n26575 );
    nor g10316 ( n16609 , n11609 , n38970 );
    nor g10317 ( n7166 , n41140 , n16510 );
    not g10318 ( n15093 , n2730 );
    not g10319 ( n28339 , n41004 );
    or g10320 ( n36994 , n38034 , n33321 );
    and g10321 ( n13381 , n31853 , n41585 );
    not g10322 ( n18581 , n18216 );
    or g10323 ( n20137 , n15560 , n27840 );
    and g10324 ( n20431 , n28620 , n8632 );
    not g10325 ( n40075 , n710 );
    or g10326 ( n38482 , n818 , n3467 );
    or g10327 ( n18205 , n19523 , n10531 );
    xnor g10328 ( n41491 , n38749 , n12375 );
    or g10329 ( n35902 , n21513 , n28062 );
    or g10330 ( n28069 , n16891 , n39008 );
    or g10331 ( n15628 , n41621 , n9216 );
    nor g10332 ( n34661 , n16773 , n2596 );
    nor g10333 ( n23560 , n31592 , n11441 );
    or g10334 ( n42548 , n12987 , n22092 );
    nor g10335 ( n22932 , n12501 , n4687 );
    or g10336 ( n27328 , n21912 , n29458 );
    or g10337 ( n13533 , n37647 , n8160 );
    or g10338 ( n21409 , n31162 , n11822 );
    nor g10339 ( n15021 , n1971 , n23670 );
    and g10340 ( n39715 , n18303 , n35202 );
    or g10341 ( n16205 , n41215 , n15600 );
    and g10342 ( n20974 , n36642 , n38468 );
    or g10343 ( n13055 , n15116 , n908 );
    and g10344 ( n10130 , n31047 , n35532 );
    or g10345 ( n22225 , n36415 , n39230 );
    or g10346 ( n34466 , n16424 , n18427 );
    nor g10347 ( n22974 , n9318 , n33768 );
    and g10348 ( n8716 , n12065 , n21808 );
    or g10349 ( n19227 , n6044 , n22468 );
    or g10350 ( n35570 , n32743 , n38191 );
    not g10351 ( n33409 , n20001 );
    or g10352 ( n4664 , n9259 , n13341 );
    or g10353 ( n14918 , n26013 , n40239 );
    or g10354 ( n38322 , n8968 , n16941 );
    and g10355 ( n1412 , n25718 , n19948 );
    and g10356 ( n2454 , n15970 , n36987 );
    and g10357 ( n29912 , n25598 , n40213 );
    and g10358 ( n26321 , n37515 , n16769 );
    xnor g10359 ( n4653 , n28443 , n31081 );
    or g10360 ( n36510 , n24569 , n18726 );
    xnor g10361 ( n12282 , n11109 , n38036 );
    not g10362 ( n19407 , n26591 );
    xnor g10363 ( n7969 , n38886 , n23463 );
    nor g10364 ( n30975 , n5398 , n13613 );
    not g10365 ( n3675 , n25763 );
    or g10366 ( n13902 , n29792 , n19935 );
    and g10367 ( n35848 , n17334 , n15207 );
    or g10368 ( n20892 , n32425 , n8128 );
    nor g10369 ( n31996 , n4271 , n29607 );
    nor g10370 ( n12181 , n32572 , n17727 );
    and g10371 ( n2101 , n15614 , n2473 );
    nor g10372 ( n20954 , n4205 , n28907 );
    xnor g10373 ( n5416 , n4697 , n7748 );
    or g10374 ( n29553 , n9022 , n39398 );
    and g10375 ( n32729 , n33052 , n20462 );
    or g10376 ( n41978 , n7864 , n41528 );
    and g10377 ( n24659 , n35781 , n7692 );
    not g10378 ( n27585 , n40918 );
    and g10379 ( n1668 , n42216 , n427 );
    and g10380 ( n8574 , n36382 , n31564 );
    not g10381 ( n22783 , n3629 );
    not g10382 ( n32548 , n47 );
    nor g10383 ( n6422 , n12409 , n5684 );
    nor g10384 ( n19950 , n38879 , n29407 );
    or g10385 ( n11659 , n30381 , n12495 );
    or g10386 ( n37293 , n24282 , n30235 );
    or g10387 ( n22236 , n30947 , n35997 );
    nor g10388 ( n36602 , n8282 , n1140 );
    not g10389 ( n10095 , n14468 );
    and g10390 ( n27278 , n1085 , n11458 );
    and g10391 ( n22211 , n35599 , n28307 );
    or g10392 ( n37406 , n27712 , n8582 );
    nor g10393 ( n17713 , n38381 , n3344 );
    not g10394 ( n7508 , n5016 );
    or g10395 ( n21843 , n38537 , n13329 );
    or g10396 ( n18380 , n40679 , n23601 );
    and g10397 ( n1648 , n20859 , n24284 );
    or g10398 ( n13661 , n38284 , n10525 );
    not g10399 ( n9852 , n31170 );
    and g10400 ( n38733 , n9906 , n18699 );
    not g10401 ( n10946 , n19712 );
    xnor g10402 ( n11506 , n12876 , n38012 );
    or g10403 ( n7319 , n26896 , n31326 );
    nor g10404 ( n33528 , n5175 , n13394 );
    xnor g10405 ( n6123 , n29740 , n20494 );
    and g10406 ( n24240 , n1398 , n22559 );
    and g10407 ( n13412 , n10310 , n2650 );
    and g10408 ( n20934 , n36178 , n9826 );
    or g10409 ( n21354 , n16393 , n20027 );
    xnor g10410 ( n13350 , n2317 , n30493 );
    or g10411 ( n8706 , n7888 , n428 );
    and g10412 ( n32243 , n10799 , n23429 );
    nor g10413 ( n90 , n23507 , n35663 );
    xnor g10414 ( n11990 , n27968 , n31773 );
    xnor g10415 ( n9219 , n31973 , n27103 );
    or g10416 ( n33689 , n35621 , n42086 );
    or g10417 ( n27097 , n12289 , n28859 );
    nor g10418 ( n13185 , n37212 , n28416 );
    or g10419 ( n33230 , n20412 , n27897 );
    and g10420 ( n26019 , n15319 , n21355 );
    or g10421 ( n13218 , n11012 , n37053 );
    nor g10422 ( n26784 , n17744 , n21176 );
    and g10423 ( n1248 , n12906 , n22756 );
    or g10424 ( n34964 , n8552 , n28289 );
    or g10425 ( n36572 , n4140 , n20382 );
    xnor g10426 ( n8116 , n29646 , n9044 );
    not g10427 ( n31123 , n6212 );
    nor g10428 ( n16239 , n41545 , n39379 );
    nor g10429 ( n29449 , n11784 , n38547 );
    nor g10430 ( n28343 , n41446 , n2723 );
    nor g10431 ( n22912 , n30862 , n6027 );
    or g10432 ( n10415 , n6560 , n24363 );
    or g10433 ( n25163 , n15874 , n29762 );
    or g10434 ( n27198 , n19794 , n40637 );
    xnor g10435 ( n38770 , n21309 , n19294 );
    not g10436 ( n34731 , n33981 );
    and g10437 ( n31466 , n14767 , n39219 );
    not g10438 ( n30453 , n37592 );
    or g10439 ( n15914 , n30435 , n39274 );
    or g10440 ( n25294 , n9781 , n12871 );
    and g10441 ( n15922 , n33255 , n40167 );
    nor g10442 ( n4081 , n7015 , n8991 );
    nor g10443 ( n22348 , n3124 , n7611 );
    or g10444 ( n12297 , n9151 , n14200 );
    or g10445 ( n13134 , n22359 , n37084 );
    and g10446 ( n18139 , n13618 , n20540 );
    nor g10447 ( n15385 , n26247 , n13679 );
    or g10448 ( n22418 , n32668 , n25784 );
    and g10449 ( n33860 , n34213 , n17200 );
    nor g10450 ( n23319 , n17193 , n20373 );
    xnor g10451 ( n28864 , n16742 , n40855 );
    not g10452 ( n33918 , n18444 );
    and g10453 ( n29278 , n19994 , n14235 );
    xnor g10454 ( n11423 , n3462 , n9341 );
    nor g10455 ( n3312 , n25588 , n9047 );
    or g10456 ( n31283 , n17654 , n29990 );
    not g10457 ( n19811 , n25592 );
    xnor g10458 ( n6112 , n25673 , n25488 );
    and g10459 ( n40574 , n5956 , n34164 );
    xnor g10460 ( n35236 , n12769 , n1211 );
    not g10461 ( n42111 , n30037 );
    or g10462 ( n36311 , n29782 , n8198 );
    or g10463 ( n38369 , n5438 , n26216 );
    not g10464 ( n3140 , n40979 );
    and g10465 ( n22988 , n6382 , n3953 );
    not g10466 ( n28831 , n20260 );
    or g10467 ( n29726 , n19041 , n27501 );
    nor g10468 ( n4376 , n38157 , n21314 );
    or g10469 ( n21182 , n33710 , n17815 );
    xnor g10470 ( n36622 , n35727 , n38538 );
    xnor g10471 ( n19660 , n29296 , n37656 );
    xnor g10472 ( n7193 , n36938 , n414 );
    nor g10473 ( n38151 , n10806 , n7869 );
    or g10474 ( n35547 , n19396 , n37872 );
    nor g10475 ( n10232 , n955 , n18341 );
    and g10476 ( n39083 , n28915 , n22431 );
    nor g10477 ( n40363 , n18477 , n37489 );
    not g10478 ( n21106 , n40531 );
    nor g10479 ( n42057 , n34419 , n34004 );
    not g10480 ( n1416 , n15476 );
    xnor g10481 ( n25809 , n25884 , n11647 );
    or g10482 ( n1277 , n17804 , n22560 );
    or g10483 ( n17824 , n36474 , n34436 );
    nor g10484 ( n35795 , n33026 , n9908 );
    nor g10485 ( n30964 , n29896 , n34183 );
    xnor g10486 ( n2962 , n31099 , n34998 );
    xnor g10487 ( n27918 , n17868 , n31952 );
    or g10488 ( n6641 , n25382 , n25298 );
    nor g10489 ( n36669 , n40902 , n34537 );
    or g10490 ( n36960 , n33235 , n22767 );
    not g10491 ( n26969 , n3280 );
    and g10492 ( n12417 , n4819 , n20809 );
    or g10493 ( n604 , n34131 , n27573 );
    and g10494 ( n40265 , n11937 , n57 );
    and g10495 ( n39072 , n32394 , n23898 );
    xnor g10496 ( n1188 , n20908 , n22838 );
    or g10497 ( n16653 , n28482 , n29075 );
    and g10498 ( n39824 , n27133 , n27899 );
    nor g10499 ( n40321 , n29575 , n6831 );
    not g10500 ( n35911 , n31169 );
    not g10501 ( n11456 , n40387 );
    or g10502 ( n35919 , n20156 , n41914 );
    not g10503 ( n23745 , n26959 );
    and g10504 ( n6425 , n11902 , n20663 );
    not g10505 ( n20254 , n12012 );
    or g10506 ( n856 , n21111 , n21420 );
    or g10507 ( n16776 , n27936 , n42870 );
    nor g10508 ( n22977 , n28752 , n36035 );
    or g10509 ( n20298 , n16108 , n7565 );
    or g10510 ( n3371 , n26922 , n16455 );
    xnor g10511 ( n13882 , n16693 , n25575 );
    or g10512 ( n37884 , n31258 , n8142 );
    xnor g10513 ( n24034 , n21534 , n22721 );
    or g10514 ( n19572 , n16671 , n9693 );
    and g10515 ( n20290 , n32131 , n4077 );
    and g10516 ( n39253 , n28753 , n2228 );
    not g10517 ( n34810 , n20737 );
    or g10518 ( n40308 , n9032 , n19057 );
    and g10519 ( n29562 , n22461 , n21626 );
    or g10520 ( n37657 , n33027 , n9335 );
    not g10521 ( n13200 , n12644 );
    and g10522 ( n33294 , n7120 , n1623 );
    and g10523 ( n17149 , n1909 , n19579 );
    or g10524 ( n13018 , n34469 , n41684 );
    and g10525 ( n34676 , n36113 , n887 );
    or g10526 ( n31455 , n25033 , n11637 );
    or g10527 ( n26037 , n9388 , n15064 );
    not g10528 ( n403 , n9694 );
    xnor g10529 ( n5487 , n13677 , n24049 );
    xnor g10530 ( n8884 , n7489 , n7350 );
    not g10531 ( n38355 , n22533 );
    not g10532 ( n35379 , n38332 );
    or g10533 ( n20765 , n12675 , n40323 );
    not g10534 ( n6171 , n24624 );
    or g10535 ( n33583 , n34855 , n7242 );
    or g10536 ( n12983 , n29080 , n29322 );
    or g10537 ( n11514 , n39249 , n11314 );
    or g10538 ( n31212 , n24488 , n41415 );
    or g10539 ( n12407 , n9234 , n29020 );
    nor g10540 ( n39127 , n4879 , n40077 );
    not g10541 ( n23053 , n17455 );
    and g10542 ( n24832 , n4912 , n20254 );
    xnor g10543 ( n21229 , n38105 , n31807 );
    and g10544 ( n22143 , n30058 , n7722 );
    and g10545 ( n32407 , n29946 , n40257 );
    xnor g10546 ( n24590 , n29129 , n32136 );
    nor g10547 ( n19144 , n17193 , n36563 );
    and g10548 ( n42705 , n16816 , n718 );
    or g10549 ( n3249 , n42735 , n10898 );
    or g10550 ( n23147 , n13662 , n18211 );
    or g10551 ( n19317 , n19144 , n28491 );
    xnor g10552 ( n20555 , n784 , n5466 );
    or g10553 ( n6028 , n23555 , n15564 );
    xnor g10554 ( n38260 , n16746 , n13573 );
    xnor g10555 ( n33437 , n2003 , n40105 );
    xnor g10556 ( n34633 , n26548 , n31957 );
    nor g10557 ( n35746 , n36215 , n32065 );
    or g10558 ( n25783 , n22117 , n20138 );
    or g10559 ( n22264 , n17744 , n4124 );
    or g10560 ( n20125 , n32046 , n21819 );
    nor g10561 ( n18784 , n39017 , n32220 );
    xnor g10562 ( n7046 , n15489 , n37931 );
    or g10563 ( n7280 , n3034 , n7011 );
    xnor g10564 ( n41844 , n6625 , n27374 );
    or g10565 ( n42267 , n18277 , n12812 );
    nor g10566 ( n17214 , n9513 , n41807 );
    not g10567 ( n34704 , n7999 );
    or g10568 ( n10752 , n13503 , n37779 );
    and g10569 ( n25036 , n14169 , n20667 );
    xnor g10570 ( n22318 , n28872 , n30112 );
    or g10571 ( n3448 , n30263 , n37728 );
    not g10572 ( n24709 , n23205 );
    not g10573 ( n18472 , n42394 );
    or g10574 ( n18540 , n7335 , n34955 );
    or g10575 ( n10747 , n37533 , n27869 );
    not g10576 ( n40768 , n6797 );
    nor g10577 ( n14140 , n20167 , n3736 );
    not g10578 ( n1219 , n32558 );
    or g10579 ( n19184 , n10542 , n29402 );
    not g10580 ( n140 , n18969 );
    nor g10581 ( n35001 , n15241 , n4184 );
    or g10582 ( n11999 , n34485 , n23468 );
    or g10583 ( n16231 , n35018 , n10351 );
    and g10584 ( n16345 , n13644 , n29599 );
    or g10585 ( n23501 , n27683 , n23063 );
    nor g10586 ( n26896 , n30161 , n3805 );
    and g10587 ( n31357 , n10990 , n19429 );
    nor g10588 ( n29874 , n42832 , n32926 );
    or g10589 ( n27809 , n9696 , n34634 );
    and g10590 ( n33604 , n12748 , n29502 );
    nor g10591 ( n22677 , n40985 , n25191 );
    nor g10592 ( n18071 , n16842 , n17423 );
    and g10593 ( n33085 , n1260 , n3861 );
    and g10594 ( n25943 , n8296 , n5965 );
    and g10595 ( n37340 , n15431 , n37246 );
    and g10596 ( n22599 , n27995 , n8077 );
    and g10597 ( n22623 , n6417 , n3683 );
    xnor g10598 ( n13570 , n21534 , n2335 );
    or g10599 ( n27152 , n20375 , n13566 );
    nor g10600 ( n1974 , n20852 , n19245 );
    not g10601 ( n3361 , n8430 );
    nor g10602 ( n25003 , n6710 , n599 );
    nor g10603 ( n28222 , n3599 , n41769 );
    and g10604 ( n26930 , n21459 , n30298 );
    or g10605 ( n42268 , n32072 , n12724 );
    or g10606 ( n26743 , n41913 , n36926 );
    or g10607 ( n26547 , n4887 , n20633 );
    or g10608 ( n648 , n28774 , n13065 );
    or g10609 ( n3232 , n19122 , n6966 );
    not g10610 ( n30036 , n16139 );
    or g10611 ( n20640 , n15107 , n22715 );
    or g10612 ( n27155 , n8494 , n37558 );
    or g10613 ( n15673 , n18490 , n32698 );
    or g10614 ( n6274 , n13710 , n21100 );
    or g10615 ( n2098 , n11025 , n42349 );
    or g10616 ( n29453 , n29181 , n34388 );
    or g10617 ( n16668 , n14642 , n21442 );
    or g10618 ( n11841 , n14868 , n19497 );
    or g10619 ( n12247 , n29625 , n28570 );
    or g10620 ( n13987 , n12192 , n34793 );
    and g10621 ( n24007 , n774 , n27541 );
    or g10622 ( n5744 , n5310 , n40428 );
    and g10623 ( n42161 , n26884 , n36613 );
    or g10624 ( n31010 , n18123 , n12892 );
    not g10625 ( n16945 , n29258 );
    nor g10626 ( n3485 , n14471 , n2077 );
    or g10627 ( n41010 , n42634 , n9752 );
    not g10628 ( n33262 , n29713 );
    or g10629 ( n25044 , n16862 , n33439 );
    not g10630 ( n12570 , n10247 );
    not g10631 ( n42514 , n17682 );
    not g10632 ( n30164 , n25821 );
    or g10633 ( n4162 , n5850 , n15199 );
    or g10634 ( n1923 , n41819 , n15077 );
    xnor g10635 ( n41542 , n17038 , n3670 );
    nor g10636 ( n8218 , n4796 , n40492 );
    or g10637 ( n17465 , n34847 , n13468 );
    and g10638 ( n1398 , n40878 , n27050 );
    and g10639 ( n8407 , n31104 , n18044 );
    xnor g10640 ( n27243 , n32048 , n9075 );
    or g10641 ( n4061 , n35722 , n14646 );
    or g10642 ( n37482 , n754 , n11128 );
    or g10643 ( n30986 , n8340 , n33081 );
    or g10644 ( n20839 , n35495 , n23857 );
    xnor g10645 ( n4229 , n31675 , n4566 );
    xnor g10646 ( n29177 , n11528 , n18616 );
    or g10647 ( n8096 , n19260 , n28863 );
    xnor g10648 ( n39537 , n36548 , n5605 );
    nor g10649 ( n10156 , n9319 , n23694 );
    and g10650 ( n34477 , n21567 , n20534 );
    or g10651 ( n21696 , n33556 , n29555 );
    or g10652 ( n10776 , n17805 , n27331 );
    or g10653 ( n12287 , n3679 , n19860 );
    or g10654 ( n29517 , n17744 , n25364 );
    not g10655 ( n40927 , n2832 );
    xnor g10656 ( n37254 , n13261 , n31216 );
    or g10657 ( n39340 , n31828 , n37250 );
    nor g10658 ( n32607 , n42048 , n24204 );
    or g10659 ( n6955 , n29430 , n38149 );
    xnor g10660 ( n23273 , n23761 , n24530 );
    xnor g10661 ( n8225 , n542 , n13807 );
    and g10662 ( n27904 , n33506 , n3967 );
    and g10663 ( n27934 , n17572 , n30104 );
    and g10664 ( n19177 , n39738 , n31826 );
    or g10665 ( n31206 , n39059 , n10191 );
    not g10666 ( n38898 , n15441 );
    or g10667 ( n16579 , n37372 , n15811 );
    not g10668 ( n10871 , n35956 );
    or g10669 ( n645 , n28211 , n6906 );
    and g10670 ( n22176 , n36093 , n31587 );
    xnor g10671 ( n8186 , n42118 , n37675 );
    and g10672 ( n34023 , n27486 , n35228 );
    or g10673 ( n4834 , n1840 , n5851 );
    and g10674 ( n35276 , n24640 , n21556 );
    and g10675 ( n31403 , n23105 , n17671 );
    and g10676 ( n23396 , n18549 , n32725 );
    and g10677 ( n2893 , n35525 , n32440 );
    and g10678 ( n6876 , n647 , n13471 );
    nor g10679 ( n26586 , n42340 , n339 );
    or g10680 ( n24145 , n25273 , n34311 );
    or g10681 ( n3964 , n22079 , n7242 );
    and g10682 ( n391 , n28845 , n31896 );
    nor g10683 ( n34877 , n34565 , n10595 );
    or g10684 ( n10662 , n9808 , n9628 );
    not g10685 ( n40261 , n13989 );
    not g10686 ( n14589 , n41841 );
    or g10687 ( n41921 , n16123 , n19267 );
    or g10688 ( n39727 , n17082 , n41082 );
    xnor g10689 ( n41165 , n20920 , n32745 );
    xnor g10690 ( n32529 , n1224 , n38574 );
    or g10691 ( n38002 , n8924 , n26845 );
    or g10692 ( n37940 , n9543 , n31321 );
    not g10693 ( n25015 , n2021 );
    or g10694 ( n39595 , n19615 , n38022 );
    or g10695 ( n23018 , n24691 , n32007 );
    or g10696 ( n19399 , n25600 , n21962 );
    nor g10697 ( n30347 , n2803 , n14779 );
    xnor g10698 ( n7655 , n4304 , n33479 );
    not g10699 ( n15429 , n14954 );
    xnor g10700 ( n8165 , n37235 , n13255 );
    nor g10701 ( n21509 , n3096 , n31767 );
    or g10702 ( n16480 , n28458 , n31892 );
    nor g10703 ( n4373 , n762 , n27839 );
    or g10704 ( n8654 , n38305 , n5813 );
    or g10705 ( n24512 , n28625 , n41990 );
    or g10706 ( n38318 , n33114 , n31976 );
    not g10707 ( n28710 , n32938 );
    and g10708 ( n12794 , n37109 , n14640 );
    xnor g10709 ( n12174 , n23080 , n10632 );
    nor g10710 ( n28639 , n19221 , n13436 );
    not g10711 ( n13488 , n15353 );
    and g10712 ( n8172 , n41986 , n14045 );
    and g10713 ( n36107 , n2389 , n645 );
    not g10714 ( n14370 , n11525 );
    not g10715 ( n6710 , n1546 );
    not g10716 ( n39941 , n29784 );
    and g10717 ( n34491 , n17330 , n41042 );
    or g10718 ( n8168 , n28235 , n28143 );
    nor g10719 ( n16328 , n38430 , n27103 );
    and g10720 ( n4997 , n3023 , n14592 );
    xnor g10721 ( n6899 , n12806 , n7048 );
    nor g10722 ( n20719 , n39266 , n36233 );
    xnor g10723 ( n20509 , n15800 , n36407 );
    and g10724 ( n19350 , n7583 , n31314 );
    nor g10725 ( n32508 , n7264 , n8779 );
    nor g10726 ( n35845 , n23311 , n12802 );
    not g10727 ( n26575 , n6196 );
    not g10728 ( n8311 , n37753 );
    or g10729 ( n1328 , n8613 , n21752 );
    not g10730 ( n19842 , n37446 );
    or g10731 ( n32399 , n29958 , n26329 );
    not g10732 ( n15706 , n12984 );
    or g10733 ( n21554 , n18914 , n853 );
    or g10734 ( n19204 , n18333 , n23417 );
    or g10735 ( n13472 , n33750 , n30701 );
    or g10736 ( n10372 , n31725 , n41709 );
    or g10737 ( n22111 , n1644 , n18498 );
    and g10738 ( n23557 , n27674 , n28378 );
    nor g10739 ( n37092 , n17120 , n13014 );
    not g10740 ( n23017 , n37919 );
    and g10741 ( n32958 , n31698 , n35007 );
    or g10742 ( n37331 , n8035 , n35639 );
    or g10743 ( n39480 , n4798 , n34827 );
    nor g10744 ( n40294 , n22011 , n39228 );
    or g10745 ( n23460 , n15715 , n36810 );
    or g10746 ( n24827 , n3606 , n36687 );
    or g10747 ( n14751 , n9063 , n24594 );
    xnor g10748 ( n29806 , n12146 , n42020 );
    or g10749 ( n14480 , n4843 , n8355 );
    and g10750 ( n38867 , n25203 , n29572 );
    xnor g10751 ( n33024 , n42499 , n19967 );
    not g10752 ( n37262 , n10116 );
    or g10753 ( n5054 , n41819 , n25125 );
    and g10754 ( n12337 , n20664 , n19972 );
    nor g10755 ( n26314 , n29079 , n23287 );
    not g10756 ( n27786 , n9671 );
    or g10757 ( n9803 , n8280 , n7028 );
    and g10758 ( n6521 , n10988 , n28558 );
    and g10759 ( n20823 , n40356 , n16523 );
    or g10760 ( n42602 , n29782 , n35809 );
    and g10761 ( n37249 , n1800 , n21144 );
    and g10762 ( n34095 , n14757 , n17996 );
    or g10763 ( n18556 , n34409 , n39602 );
    not g10764 ( n15111 , n25370 );
    xnor g10765 ( n24951 , n542 , n3556 );
    not g10766 ( n13785 , n36776 );
    and g10767 ( n42099 , n38879 , n11479 );
    or g10768 ( n16278 , n13308 , n15689 );
    or g10769 ( n21310 , n6717 , n4316 );
    and g10770 ( n13186 , n21427 , n1605 );
    or g10771 ( n5164 , n30071 , n22945 );
    nor g10772 ( n31889 , n36510 , n14477 );
    or g10773 ( n23877 , n21342 , n10953 );
    nor g10774 ( n14600 , n42042 , n5075 );
    nor g10775 ( n14387 , n36135 , n30042 );
    not g10776 ( n27313 , n1411 );
    or g10777 ( n4894 , n31542 , n8601 );
    and g10778 ( n20133 , n784 , n16983 );
    or g10779 ( n8142 , n19969 , n16078 );
    or g10780 ( n29125 , n23261 , n32494 );
    and g10781 ( n22230 , n13902 , n21350 );
    and g10782 ( n38343 , n31402 , n8250 );
    or g10783 ( n19988 , n17848 , n28510 );
    or g10784 ( n16342 , n8035 , n38869 );
    and g10785 ( n30314 , n25832 , n10578 );
    and g10786 ( n39849 , n35254 , n31253 );
    nor g10787 ( n38755 , n39367 , n27551 );
    xnor g10788 ( n429 , n22082 , n42752 );
    or g10789 ( n31744 , n4018 , n38902 );
    and g10790 ( n23426 , n1983 , n37997 );
    or g10791 ( n24473 , n30629 , n20618 );
    not g10792 ( n14553 , n33438 );
    xnor g10793 ( n13420 , n15796 , n35631 );
    not g10794 ( n17888 , n861 );
    xnor g10795 ( n41769 , n30397 , n4815 );
    or g10796 ( n1241 , n14434 , n11797 );
    xnor g10797 ( n32926 , n24527 , n17924 );
    not g10798 ( n30614 , n21175 );
    xnor g10799 ( n18231 , n35727 , n41493 );
    and g10800 ( n40790 , n2293 , n19749 );
    or g10801 ( n29544 , n18475 , n15265 );
    nor g10802 ( n4479 , n20668 , n10221 );
    or g10803 ( n39833 , n40156 , n8401 );
    or g10804 ( n30803 , n28149 , n17620 );
    xnor g10805 ( n34310 , n28691 , n9076 );
    xnor g10806 ( n26402 , n26579 , n20407 );
    or g10807 ( n20930 , n13030 , n12179 );
    or g10808 ( n39835 , n16999 , n8864 );
    or g10809 ( n36805 , n31898 , n2044 );
    not g10810 ( n14969 , n2135 );
    and g10811 ( n13130 , n29999 , n35659 );
    and g10812 ( n2052 , n29005 , n42758 );
    or g10813 ( n33618 , n8539 , n35095 );
    nor g10814 ( n7131 , n3430 , n22262 );
    or g10815 ( n8131 , n36703 , n22127 );
    or g10816 ( n6520 , n6381 , n34792 );
    nor g10817 ( n6286 , n30543 , n38747 );
    and g10818 ( n33845 , n39124 , n3039 );
    nor g10819 ( n25850 , n34565 , n9823 );
    not g10820 ( n32838 , n22303 );
    not g10821 ( n38836 , n9977 );
    or g10822 ( n5686 , n2867 , n425 );
    and g10823 ( n38405 , n10059 , n11219 );
    or g10824 ( n8801 , n15116 , n42570 );
    and g10825 ( n19173 , n24978 , n9209 );
    and g10826 ( n12887 , n21401 , n25095 );
    or g10827 ( n26880 , n38441 , n4760 );
    and g10828 ( n41839 , n33364 , n17784 );
    nor g10829 ( n38201 , n5896 , n37817 );
    not g10830 ( n35505 , n23814 );
    not g10831 ( n8093 , n13251 );
    not g10832 ( n2031 , n21255 );
    or g10833 ( n6378 , n20486 , n42034 );
    not g10834 ( n11455 , n3680 );
    or g10835 ( n37534 , n24307 , n21203 );
    or g10836 ( n38330 , n28470 , n37371 );
    nor g10837 ( n20122 , n22473 , n4928 );
    or g10838 ( n12875 , n7572 , n42243 );
    or g10839 ( n19595 , n31130 , n34456 );
    xnor g10840 ( n812 , n12146 , n13337 );
    and g10841 ( n39923 , n37168 , n33827 );
    or g10842 ( n14284 , n20437 , n30710 );
    or g10843 ( n5326 , n18413 , n17983 );
    and g10844 ( n18387 , n20070 , n10548 );
    not g10845 ( n17522 , n8508 );
    not g10846 ( n27715 , n39955 );
    xnor g10847 ( n7074 , n3277 , n30241 );
    and g10848 ( n13958 , n41024 , n21039 );
    and g10849 ( n7953 , n36341 , n35676 );
    xnor g10850 ( n42843 , n13444 , n24349 );
    nor g10851 ( n26296 , n14642 , n9459 );
    xnor g10852 ( n11817 , n4877 , n12562 );
    nor g10853 ( n25157 , n30220 , n19477 );
    nor g10854 ( n37075 , n24699 , n27954 );
    not g10855 ( n12105 , n40861 );
    nor g10856 ( n14432 , n32023 , n1480 );
    xnor g10857 ( n20047 , n6625 , n29909 );
    not g10858 ( n20571 , n10835 );
    xnor g10859 ( n509 , n136 , n25390 );
    and g10860 ( n7719 , n28814 , n41135 );
    nor g10861 ( n9365 , n10271 , n38660 );
    or g10862 ( n19604 , n27598 , n1067 );
    nor g10863 ( n24595 , n39266 , n31679 );
    and g10864 ( n40345 , n14824 , n37085 );
    and g10865 ( n9663 , n25915 , n15449 );
    not g10866 ( n32728 , n34476 );
    and g10867 ( n13081 , n8634 , n29160 );
    xnor g10868 ( n37907 , n42064 , n18426 );
    and g10869 ( n30895 , n22581 , n10348 );
    and g10870 ( n42891 , n11481 , n23061 );
    and g10871 ( n41297 , n40224 , n42863 );
    or g10872 ( n2357 , n15791 , n17827 );
    and g10873 ( n4227 , n10270 , n31085 );
    or g10874 ( n4393 , n2007 , n33139 );
    or g10875 ( n39561 , n14287 , n9341 );
    or g10876 ( n4344 , n12235 , n699 );
    nor g10877 ( n26834 , n25602 , n6188 );
    nor g10878 ( n5200 , n35259 , n6406 );
    or g10879 ( n41138 , n29043 , n17752 );
    not g10880 ( n24437 , n13896 );
    or g10881 ( n26324 , n8970 , n15940 );
    and g10882 ( n871 , n28717 , n26209 );
    and g10883 ( n10851 , n10154 , n40776 );
    or g10884 ( n18047 , n22933 , n8535 );
    not g10885 ( n23778 , n11137 );
    or g10886 ( n3233 , n11885 , n3580 );
    nor g10887 ( n948 , n18424 , n5039 );
    or g10888 ( n8392 , n15770 , n27384 );
    or g10889 ( n13925 , n5663 , n11321 );
    or g10890 ( n30431 , n5670 , n21297 );
    not g10891 ( n17084 , n38444 );
    not g10892 ( n2727 , n36745 );
    and g10893 ( n35405 , n29823 , n4876 );
    or g10894 ( n17263 , n8847 , n41787 );
    or g10895 ( n35630 , n37903 , n21924 );
    or g10896 ( n41020 , n3387 , n23700 );
    not g10897 ( n10698 , n41956 );
    or g10898 ( n42541 , n26114 , n12260 );
    or g10899 ( n6922 , n30368 , n1017 );
    or g10900 ( n20445 , n32193 , n27552 );
    not g10901 ( n18476 , n29673 );
    and g10902 ( n12072 , n24211 , n21163 );
    or g10903 ( n15328 , n12397 , n477 );
    and g10904 ( n13852 , n28806 , n3658 );
    or g10905 ( n1071 , n4998 , n12153 );
    and g10906 ( n25960 , n37750 , n19895 );
    or g10907 ( n21369 , n2199 , n27091 );
    xnor g10908 ( n16301 , n4767 , n5964 );
    or g10909 ( n34581 , n22117 , n328 );
    and g10910 ( n37803 , n38318 , n31289 );
    or g10911 ( n29362 , n30458 , n4995 );
    and g10912 ( n37315 , n4967 , n31340 );
    or g10913 ( n13257 , n9400 , n41932 );
    or g10914 ( n16737 , n42588 , n13368 );
    or g10915 ( n37959 , n8433 , n30652 );
    not g10916 ( n2022 , n18637 );
    nor g10917 ( n21160 , n16387 , n38636 );
    or g10918 ( n22132 , n35933 , n14569 );
    xnor g10919 ( n2923 , n784 , n10476 );
    and g10920 ( n25694 , n15291 , n23791 );
    and g10921 ( n4696 , n30160 , n36043 );
    nor g10922 ( n26156 , n35009 , n20283 );
    and g10923 ( n21109 , n15156 , n40565 );
    or g10924 ( n34309 , n26108 , n25418 );
    nor g10925 ( n37560 , n18320 , n10505 );
    or g10926 ( n39547 , n3855 , n21942 );
    or g10927 ( n35964 , n12722 , n2739 );
    nor g10928 ( n36653 , n18866 , n24801 );
    xnor g10929 ( n16366 , n8529 , n42606 );
    or g10930 ( n5777 , n17033 , n1812 );
    and g10931 ( n3920 , n25927 , n31558 );
    or g10932 ( n11630 , n8419 , n10707 );
    not g10933 ( n41356 , n40197 );
    or g10934 ( n30823 , n35722 , n9735 );
    not g10935 ( n27987 , n4517 );
    or g10936 ( n27800 , n29646 , n23530 );
    nor g10937 ( n508 , n1254 , n1804 );
    or g10938 ( n18693 , n29767 , n19961 );
    not g10939 ( n9880 , n36154 );
    and g10940 ( n23005 , n494 , n33939 );
    not g10941 ( n11439 , n16982 );
    and g10942 ( n13335 , n26100 , n26866 );
    or g10943 ( n27498 , n41197 , n3414 );
    or g10944 ( n24561 , n31981 , n39267 );
    not g10945 ( n16527 , n7771 );
    or g10946 ( n12659 , n40174 , n16073 );
    xnor g10947 ( n20333 , n6625 , n17037 );
    and g10948 ( n21091 , n39020 , n1272 );
    or g10949 ( n27046 , n22821 , n32884 );
    and g10950 ( n19587 , n37999 , n25786 );
    not g10951 ( n32297 , n10598 );
    or g10952 ( n31484 , n15064 , n4408 );
    or g10953 ( n39643 , n15820 , n26111 );
    or g10954 ( n27849 , n20241 , n14776 );
    or g10955 ( n18669 , n11688 , n2802 );
    or g10956 ( n30904 , n42416 , n16476 );
    or g10957 ( n25974 , n1327 , n170 );
    or g10958 ( n13800 , n2701 , n12818 );
    xnor g10959 ( n4537 , n5891 , n6029 );
    not g10960 ( n14389 , n16535 );
    and g10961 ( n3006 , n7806 , n16111 );
    or g10962 ( n41329 , n2132 , n23921 );
    or g10963 ( n39530 , n41201 , n6472 );
    or g10964 ( n5731 , n34365 , n10455 );
    nor g10965 ( n19278 , n16598 , n21164 );
    and g10966 ( n36024 , n13491 , n42737 );
    xnor g10967 ( n30641 , n35727 , n12619 );
    xnor g10968 ( n8408 , n16722 , n21497 );
    or g10969 ( n33371 , n30971 , n16164 );
    or g10970 ( n12154 , n13048 , n7716 );
    or g10971 ( n37772 , n38249 , n8577 );
    or g10972 ( n1831 , n8907 , n19293 );
    xnor g10973 ( n9167 , n30549 , n27998 );
    or g10974 ( n14516 , n19186 , n37399 );
    and g10975 ( n3275 , n7688 , n6983 );
    or g10976 ( n18512 , n26874 , n17992 );
    or g10977 ( n3585 , n37910 , n421 );
    not g10978 ( n15137 , n38344 );
    nor g10979 ( n41824 , n31682 , n10686 );
    nor g10980 ( n40444 , n35301 , n24349 );
    not g10981 ( n39330 , n10848 );
    or g10982 ( n38442 , n3583 , n34432 );
    and g10983 ( n13165 , n10502 , n7698 );
    or g10984 ( n7420 , n14668 , n1928 );
    nor g10985 ( n26951 , n20456 , n5446 );
    or g10986 ( n8807 , n6170 , n8893 );
    not g10987 ( n3905 , n37170 );
    not g10988 ( n38191 , n4331 );
    or g10989 ( n17237 , n14125 , n15837 );
    or g10990 ( n31308 , n40446 , n29500 );
    or g10991 ( n19800 , n20138 , n33990 );
    and g10992 ( n22666 , n13257 , n36981 );
    nor g10993 ( n20180 , n38543 , n14376 );
    not g10994 ( n13731 , n22383 );
    and g10995 ( n19352 , n23994 , n29569 );
    or g10996 ( n2783 , n7821 , n38006 );
    nor g10997 ( n25201 , n40757 , n9863 );
    or g10998 ( n22238 , n32324 , n36641 );
    or g10999 ( n42101 , n39699 , n10534 );
    and g11000 ( n21152 , n15237 , n40219 );
    not g11001 ( n30877 , n3898 );
    xnor g11002 ( n14779 , n27734 , n7504 );
    or g11003 ( n35435 , n30113 , n32068 );
    xnor g11004 ( n19785 , n2659 , n15211 );
    and g11005 ( n41176 , n13749 , n10056 );
    or g11006 ( n3613 , n13250 , n39744 );
    or g11007 ( n24009 , n20138 , n5481 );
    nor g11008 ( n27231 , n10969 , n11963 );
    not g11009 ( n1214 , n33199 );
    and g11010 ( n20403 , n37745 , n32592 );
    or g11011 ( n26069 , n23397 , n27187 );
    xnor g11012 ( n36684 , n20557 , n17145 );
    and g11013 ( n1353 , n32560 , n10508 );
    and g11014 ( n25038 , n14318 , n1834 );
    or g11015 ( n29317 , n3389 , n39408 );
    and g11016 ( n16095 , n22360 , n22083 );
    not g11017 ( n24657 , n10210 );
    not g11018 ( n31857 , n17454 );
    and g11019 ( n41777 , n24804 , n41874 );
    not g11020 ( n16617 , n1542 );
    or g11021 ( n28771 , n6004 , n23315 );
    not g11022 ( n15617 , n10962 );
    or g11023 ( n35892 , n39187 , n33139 );
    nor g11024 ( n1968 , n37393 , n5221 );
    and g11025 ( n15346 , n30275 , n1405 );
    not g11026 ( n7197 , n4424 );
    or g11027 ( n28521 , n11599 , n15149 );
    or g11028 ( n20132 , n35684 , n20402 );
    or g11029 ( n20915 , n32957 , n18707 );
    or g11030 ( n17490 , n9501 , n36189 );
    nor g11031 ( n2883 , n30766 , n9450 );
    and g11032 ( n18441 , n34216 , n28450 );
    not g11033 ( n10863 , n13453 );
    nor g11034 ( n3962 , n7840 , n15610 );
    not g11035 ( n1611 , n36497 );
    not g11036 ( n3769 , n9691 );
    not g11037 ( n11938 , n29879 );
    not g11038 ( n4807 , n19430 );
    or g11039 ( n14296 , n21242 , n39924 );
    or g11040 ( n7876 , n18475 , n27933 );
    and g11041 ( n34607 , n41937 , n20864 );
    nor g11042 ( n26459 , n18131 , n3588 );
    or g11043 ( n26750 , n24698 , n9536 );
    or g11044 ( n23889 , n21805 , n9160 );
    not g11045 ( n26226 , n4382 );
    and g11046 ( n39000 , n38101 , n12865 );
    and g11047 ( n20276 , n35653 , n18050 );
    xnor g11048 ( n12109 , n27968 , n19960 );
    not g11049 ( n39108 , n1013 );
    and g11050 ( n24468 , n30456 , n901 );
    or g11051 ( n27911 , n18606 , n25451 );
    xnor g11052 ( n20964 , n17220 , n11433 );
    or g11053 ( n16642 , n27752 , n10234 );
    and g11054 ( n8610 , n21577 , n13183 );
    not g11055 ( n24122 , n20481 );
    or g11056 ( n18982 , n42220 , n206 );
    and g11057 ( n35544 , n5703 , n35955 );
    nor g11058 ( n239 , n37287 , n4073 );
    or g11059 ( n16405 , n15070 , n1651 );
    nor g11060 ( n21620 , n68 , n9756 );
    not g11061 ( n41119 , n7801 );
    or g11062 ( n36612 , n20802 , n12403 );
    and g11063 ( n4276 , n39458 , n14570 );
    or g11064 ( n24854 , n40044 , n22991 );
    nor g11065 ( n21085 , n1313 , n29331 );
    xnor g11066 ( n28767 , n42127 , n9485 );
    or g11067 ( n20620 , n20650 , n14569 );
    not g11068 ( n21856 , n17406 );
    and g11069 ( n15935 , n36982 , n23899 );
    and g11070 ( n24055 , n42113 , n42845 );
    or g11071 ( n42313 , n9797 , n38317 );
    or g11072 ( n22254 , n35757 , n9617 );
    and g11073 ( n6501 , n12723 , n42081 );
    not g11074 ( n5203 , n32001 );
    and g11075 ( n32102 , n40751 , n17605 );
    not g11076 ( n5082 , n9127 );
    or g11077 ( n22774 , n32245 , n18208 );
    not g11078 ( n28211 , n28016 );
    and g11079 ( n26590 , n1515 , n36592 );
    or g11080 ( n15477 , n12291 , n560 );
    or g11081 ( n16385 , n23034 , n11122 );
    and g11082 ( n28214 , n995 , n38062 );
    or g11083 ( n9558 , n20684 , n18851 );
    or g11084 ( n13900 , n13965 , n26713 );
    or g11085 ( n2873 , n24523 , n35016 );
    nor g11086 ( n38138 , n36117 , n30672 );
    or g11087 ( n36270 , n34256 , n28239 );
    and g11088 ( n25933 , n4430 , n36083 );
    and g11089 ( n6769 , n9872 , n6404 );
    nor g11090 ( n3985 , n40585 , n13205 );
    or g11091 ( n3523 , n41567 , n19788 );
    or g11092 ( n12160 , n22569 , n14992 );
    xnor g11093 ( n8132 , n14377 , n12492 );
    or g11094 ( n22165 , n40324 , n3570 );
    and g11095 ( n12991 , n17917 , n20467 );
    or g11096 ( n22673 , n6924 , n21807 );
    not g11097 ( n71 , n13111 );
    nor g11098 ( n5037 , n42583 , n35399 );
    nor g11099 ( n24421 , n1458 , n35591 );
    or g11100 ( n31396 , n8090 , n46 );
    and g11101 ( n33031 , n20487 , n33341 );
    or g11102 ( n17444 , n4145 , n23372 );
    xnor g11103 ( n41518 , n34875 , n4850 );
    and g11104 ( n11188 , n26124 , n13537 );
    and g11105 ( n34925 , n33568 , n2730 );
    or g11106 ( n37661 , n8289 , n36514 );
    or g11107 ( n12380 , n36850 , n35265 );
    or g11108 ( n16050 , n41705 , n9722 );
    not g11109 ( n20983 , n13386 );
    or g11110 ( n4985 , n11739 , n19074 );
    nor g11111 ( n27059 , n33981 , n32884 );
    and g11112 ( n19957 , n25257 , n23074 );
    not g11113 ( n34637 , n18046 );
    or g11114 ( n29578 , n35328 , n18100 );
    not g11115 ( n39519 , n32633 );
    nor g11116 ( n33237 , n17744 , n5647 );
    not g11117 ( n38784 , n10857 );
    nor g11118 ( n36167 , n14356 , n8211 );
    not g11119 ( n32475 , n10587 );
    not g11120 ( n1581 , n36811 );
    or g11121 ( n1915 , n3342 , n2626 );
    xnor g11122 ( n26509 , n2174 , n21218 );
    or g11123 ( n32202 , n10284 , n10586 );
    or g11124 ( n15539 , n25265 , n14064 );
    nor g11125 ( n26211 , n19522 , n21433 );
    xnor g11126 ( n9110 , n10427 , n18353 );
    and g11127 ( n36646 , n38739 , n15219 );
    xnor g11128 ( n1490 , n105 , n36946 );
    or g11129 ( n25492 , n35292 , n17795 );
    xnor g11130 ( n4360 , n14052 , n31165 );
    or g11131 ( n21456 , n4538 , n12814 );
    and g11132 ( n42845 , n5855 , n29213 );
    nor g11133 ( n24341 , n14168 , n34891 );
    nor g11134 ( n24470 , n31639 , n10764 );
    or g11135 ( n11484 , n3583 , n4606 );
    or g11136 ( n40817 , n3559 , n17542 );
    or g11137 ( n10006 , n10092 , n13673 );
    not g11138 ( n10612 , n18134 );
    not g11139 ( n34093 , n29086 );
    or g11140 ( n25955 , n41406 , n30231 );
    or g11141 ( n42190 , n650 , n33826 );
    or g11142 ( n5549 , n14281 , n12035 );
    not g11143 ( n38685 , n27895 );
    xnor g11144 ( n27708 , n8868 , n6816 );
    xnor g11145 ( n42542 , n105 , n41787 );
    or g11146 ( n17358 , n4969 , n41496 );
    not g11147 ( n37466 , n42560 );
    not g11148 ( n24972 , n28578 );
    or g11149 ( n32950 , n32217 , n37803 );
    xnor g11150 ( n35682 , n15343 , n38889 );
    or g11151 ( n14359 , n27445 , n1199 );
    and g11152 ( n31323 , n18867 , n29620 );
    and g11153 ( n27680 , n34336 , n30047 );
    and g11154 ( n40154 , n379 , n9124 );
    not g11155 ( n803 , n37961 );
    or g11156 ( n5667 , n35247 , n8998 );
    or g11157 ( n2324 , n851 , n8661 );
    or g11158 ( n640 , n972 , n33809 );
    or g11159 ( n21419 , n4904 , n2561 );
    not g11160 ( n1785 , n27274 );
    and g11161 ( n3084 , n41023 , n11354 );
    not g11162 ( n36853 , n21870 );
    or g11163 ( n24207 , n26915 , n24123 );
    nor g11164 ( n22567 , n32461 , n32706 );
    and g11165 ( n21195 , n41805 , n8969 );
    or g11166 ( n7619 , n11373 , n25742 );
    and g11167 ( n5526 , n31454 , n2779 );
    or g11168 ( n29397 , n17108 , n29685 );
    nor g11169 ( n33143 , n17226 , n11041 );
    or g11170 ( n20902 , n20292 , n8314 );
    and g11171 ( n29521 , n4733 , n31645 );
    or g11172 ( n14857 , n27130 , n13830 );
    not g11173 ( n19653 , n21974 );
    not g11174 ( n40275 , n25623 );
    and g11175 ( n987 , n17974 , n25075 );
    or g11176 ( n37926 , n23478 , n20201 );
    or g11177 ( n23185 , n2012 , n25061 );
    nor g11178 ( n17066 , n42272 , n12072 );
    or g11179 ( n2634 , n13416 , n31503 );
    or g11180 ( n9198 , n34091 , n24857 );
    and g11181 ( n1296 , n32059 , n41794 );
    and g11182 ( n7966 , n4034 , n4830 );
    not g11183 ( n13607 , n29150 );
    nor g11184 ( n26628 , n38640 , n31427 );
    nor g11185 ( n3305 , n14707 , n38740 );
    and g11186 ( n6125 , n5857 , n37301 );
    or g11187 ( n31739 , n2811 , n22355 );
    or g11188 ( n22431 , n12666 , n17975 );
    and g11189 ( n18583 , n29740 , n19674 );
    or g11190 ( n32493 , n22065 , n30373 );
    xnor g11191 ( n27751 , n784 , n17356 );
    and g11192 ( n14216 , n20671 , n25632 );
    not g11193 ( n41649 , n20513 );
    and g11194 ( n7795 , n12779 , n12673 );
    nor g11195 ( n14029 , n20945 , n26629 );
    and g11196 ( n9825 , n30292 , n21798 );
    not g11197 ( n29988 , n18041 );
    not g11198 ( n41583 , n4139 );
    or g11199 ( n16118 , n29054 , n16654 );
    nor g11200 ( n22935 , n41856 , n35511 );
    nor g11201 ( n34400 , n11799 , n2140 );
    or g11202 ( n36079 , n5742 , n41413 );
    not g11203 ( n6919 , n22483 );
    and g11204 ( n37622 , n20487 , n475 );
    or g11205 ( n15027 , n6944 , n9858 );
    not g11206 ( n6273 , n5097 );
    or g11207 ( n29850 , n30068 , n30912 );
    xnor g11208 ( n352 , n31539 , n20680 );
    and g11209 ( n12845 , n33536 , n18845 );
    and g11210 ( n31720 , n22890 , n14175 );
    and g11211 ( n14325 , n33376 , n27115 );
    and g11212 ( n11004 , n41531 , n6256 );
    and g11213 ( n10632 , n1195 , n3228 );
    nor g11214 ( n15951 , n20016 , n10732 );
    or g11215 ( n17265 , n19580 , n22203 );
    xnor g11216 ( n8832 , n25809 , n3221 );
    xnor g11217 ( n17121 , n38084 , n31120 );
    or g11218 ( n14482 , n17359 , n22430 );
    not g11219 ( n40881 , n39873 );
    and g11220 ( n33272 , n16165 , n12736 );
    nor g11221 ( n9577 , n28938 , n33505 );
    xnor g11222 ( n29037 , n24573 , n22111 );
    or g11223 ( n28437 , n33683 , n38924 );
    not g11224 ( n23591 , n22872 );
    nor g11225 ( n33472 , n33532 , n29674 );
    not g11226 ( n6145 , n10279 );
    nor g11227 ( n14691 , n12362 , n4851 );
    or g11228 ( n4604 , n27156 , n16610 );
    or g11229 ( n17987 , n38093 , n36844 );
    or g11230 ( n32030 , n14945 , n25309 );
    or g11231 ( n11101 , n25121 , n38196 );
    or g11232 ( n12507 , n3164 , n10215 );
    or g11233 ( n38108 , n13265 , n2654 );
    or g11234 ( n38071 , n35143 , n18494 );
    or g11235 ( n1041 , n26689 , n18173 );
    or g11236 ( n13252 , n1507 , n19017 );
    and g11237 ( n28453 , n23402 , n17818 );
    not g11238 ( n9417 , n17327 );
    and g11239 ( n18860 , n39994 , n39427 );
    nor g11240 ( n1550 , n29308 , n26232 );
    xnor g11241 ( n20560 , n34731 , n28721 );
    not g11242 ( n34951 , n12651 );
    and g11243 ( n37321 , n34476 , n8521 );
    and g11244 ( n30631 , n30516 , n20884 );
    not g11245 ( n42791 , n9974 );
    or g11246 ( n34526 , n10880 , n36619 );
    not g11247 ( n836 , n22454 );
    nor g11248 ( n19826 , n14471 , n4312 );
    not g11249 ( n25483 , n19196 );
    not g11250 ( n6290 , n14888 );
    or g11251 ( n7584 , n31051 , n9752 );
    or g11252 ( n39836 , n35170 , n31444 );
    xnor g11253 ( n31874 , n34951 , n24602 );
    or g11254 ( n11698 , n2183 , n38034 );
    or g11255 ( n20600 , n35633 , n29063 );
    or g11256 ( n19860 , n11976 , n8107 );
    or g11257 ( n32557 , n38508 , n23703 );
    not g11258 ( n29214 , n30845 );
    or g11259 ( n3823 , n4422 , n35695 );
    xnor g11260 ( n24120 , n5144 , n2713 );
    and g11261 ( n26448 , n27866 , n38049 );
    not g11262 ( n10397 , n3335 );
    or g11263 ( n32854 , n4335 , n39282 );
    nor g11264 ( n20634 , n20223 , n1101 );
    and g11265 ( n32125 , n40158 , n31744 );
    and g11266 ( n34338 , n24507 , n36906 );
    xnor g11267 ( n27623 , n30830 , n38639 );
    or g11268 ( n1672 , n21544 , n29914 );
    or g11269 ( n42172 , n37248 , n15784 );
    or g11270 ( n6256 , n7394 , n15410 );
    or g11271 ( n35819 , n7356 , n29712 );
    not g11272 ( n1011 , n3539 );
    or g11273 ( n3757 , n1183 , n24366 );
    or g11274 ( n25139 , n14139 , n39117 );
    not g11275 ( n22427 , n14233 );
    and g11276 ( n33558 , n38749 , n8821 );
    or g11277 ( n36480 , n10845 , n15409 );
    nor g11278 ( n28965 , n41665 , n32153 );
    or g11279 ( n14187 , n35930 , n24709 );
    and g11280 ( n20561 , n12299 , n2888 );
    or g11281 ( n2725 , n11327 , n12359 );
    or g11282 ( n8622 , n30144 , n14405 );
    or g11283 ( n37801 , n5362 , n19131 );
    and g11284 ( n19259 , n18109 , n26648 );
    nor g11285 ( n36477 , n42700 , n23470 );
    nor g11286 ( n24934 , n34565 , n40722 );
    and g11287 ( n19460 , n17227 , n9966 );
    or g11288 ( n4640 , n34728 , n10108 );
    and g11289 ( n12541 , n6967 , n20798 );
    or g11290 ( n2425 , n3472 , n5183 );
    or g11291 ( n24398 , n19576 , n42749 );
    not g11292 ( n34277 , n20889 );
    nor g11293 ( n20153 , n6929 , n31059 );
    or g11294 ( n23798 , n12618 , n18354 );
    nor g11295 ( n1408 , n15179 , n39512 );
    or g11296 ( n17316 , n16318 , n22885 );
    not g11297 ( n14501 , n9588 );
    and g11298 ( n40517 , n21012 , n1235 );
    nor g11299 ( n24098 , n12885 , n32114 );
    or g11300 ( n31635 , n33529 , n7289 );
    and g11301 ( n9670 , n41755 , n98 );
    and g11302 ( n12787 , n16230 , n37618 );
    and g11303 ( n145 , n4425 , n32735 );
    nor g11304 ( n17858 , n18866 , n29693 );
    not g11305 ( n21172 , n25756 );
    or g11306 ( n35904 , n37119 , n3563 );
    nor g11307 ( n4656 , n4004 , n23669 );
    or g11308 ( n8095 , n14634 , n39108 );
    not g11309 ( n8123 , n42332 );
    xnor g11310 ( n2278 , n33420 , n33315 );
    xnor g11311 ( n40227 , n8502 , n21047 );
    or g11312 ( n20444 , n1248 , n12153 );
    not g11313 ( n37890 , n34858 );
    or g11314 ( n9716 , n3629 , n15982 );
    xnor g11315 ( n19154 , n1762 , n34007 );
    or g11316 ( n42063 , n4608 , n24701 );
    nor g11317 ( n6504 , n35073 , n25302 );
    not g11318 ( n23282 , n12629 );
    or g11319 ( n42573 , n39962 , n4700 );
    nor g11320 ( n32097 , n15070 , n31101 );
    and g11321 ( n22359 , n20462 , n21753 );
    or g11322 ( n41647 , n9646 , n19890 );
    and g11323 ( n3785 , n28703 , n31239 );
    or g11324 ( n32330 , n25313 , n18705 );
    or g11325 ( n12029 , n42746 , n2701 );
    or g11326 ( n28681 , n24027 , n10837 );
    and g11327 ( n8267 , n18787 , n18583 );
    or g11328 ( n24112 , n35188 , n38293 );
    or g11329 ( n27391 , n3213 , n11907 );
    or g11330 ( n42141 , n28515 , n2913 );
    xnor g11331 ( n14229 , n11436 , n15935 );
    and g11332 ( n20694 , n16554 , n24655 );
    or g11333 ( n32617 , n16738 , n12352 );
    and g11334 ( n7463 , n38916 , n34770 );
    not g11335 ( n11879 , n19248 );
    and g11336 ( n35581 , n25388 , n26660 );
    and g11337 ( n20760 , n33335 , n18603 );
    or g11338 ( n29576 , n15445 , n108 );
    or g11339 ( n33404 , n37212 , n13664 );
    and g11340 ( n15500 , n8671 , n36465 );
    not g11341 ( n40531 , n12068 );
    xnor g11342 ( n9441 , n41218 , n22928 );
    not g11343 ( n1117 , n7740 );
    and g11344 ( n326 , n21692 , n21436 );
    or g11345 ( n9006 , n17435 , n24281 );
    not g11346 ( n35802 , n14619 );
    or g11347 ( n22813 , n16605 , n12122 );
    or g11348 ( n38310 , n7835 , n14708 );
    and g11349 ( n11732 , n33061 , n39362 );
    nor g11350 ( n40384 , n19039 , n28259 );
    and g11351 ( n5927 , n4027 , n19947 );
    or g11352 ( n15532 , n23977 , n16150 );
    or g11353 ( n15750 , n3351 , n34569 );
    or g11354 ( n31280 , n26777 , n24559 );
    not g11355 ( n8790 , n20761 );
    xnor g11356 ( n31819 , n31917 , n12541 );
    and g11357 ( n30216 , n39041 , n12142 );
    or g11358 ( n7038 , n14730 , n18200 );
    and g11359 ( n23757 , n28622 , n41693 );
    or g11360 ( n35326 , n10934 , n26090 );
    xnor g11361 ( n26182 , n25582 , n15545 );
    xnor g11362 ( n4962 , n9268 , n31377 );
    or g11363 ( n36039 , n42340 , n34981 );
    xnor g11364 ( n40555 , n16929 , n5605 );
    not g11365 ( n19486 , n14224 );
    and g11366 ( n37642 , n3842 , n1045 );
    not g11367 ( n25877 , n9401 );
    nor g11368 ( n25285 , n2753 , n38909 );
    not g11369 ( n19398 , n39450 );
    or g11370 ( n17778 , n23300 , n28065 );
    or g11371 ( n7318 , n36902 , n2802 );
    and g11372 ( n32839 , n29891 , n16345 );
    not g11373 ( n25649 , n40496 );
    nor g11374 ( n22396 , n40476 , n41799 );
    not g11375 ( n1078 , n3512 );
    and g11376 ( n35764 , n17993 , n29379 );
    or g11377 ( n37192 , n6279 , n23189 );
    or g11378 ( n28926 , n5795 , n10013 );
    not g11379 ( n33770 , n24046 );
    or g11380 ( n31740 , n31494 , n8104 );
    not g11381 ( n24179 , n29470 );
    not g11382 ( n21710 , n31780 );
    not g11383 ( n34793 , n26836 );
    or g11384 ( n39007 , n6911 , n26158 );
    xnor g11385 ( n18442 , n31895 , n33156 );
    and g11386 ( n18830 , n42064 , n25598 );
    or g11387 ( n40822 , n35291 , n31007 );
    xnor g11388 ( n27820 , n15324 , n37267 );
    or g11389 ( n13091 , n6658 , n11523 );
    or g11390 ( n21405 , n31299 , n23121 );
    not g11391 ( n17957 , n26722 );
    and g11392 ( n15448 , n39280 , n16763 );
    xnor g11393 ( n24067 , n42725 , n36169 );
    and g11394 ( n37208 , n39527 , n18290 );
    not g11395 ( n18812 , n36776 );
    not g11396 ( n2733 , n42451 );
    or g11397 ( n1922 , n38057 , n18393 );
    nor g11398 ( n15327 , n4516 , n16059 );
    not g11399 ( n12878 , n17610 );
    or g11400 ( n12363 , n34849 , n37250 );
    xnor g11401 ( n2266 , n39279 , n26019 );
    and g11402 ( n5647 , n628 , n37575 );
    and g11403 ( n27221 , n12009 , n25555 );
    or g11404 ( n36150 , n39802 , n20446 );
    not g11405 ( n6956 , n12370 );
    or g11406 ( n1195 , n17867 , n39924 );
    or g11407 ( n10186 , n18347 , n17370 );
    not g11408 ( n1054 , n21744 );
    not g11409 ( n11594 , n32175 );
    xnor g11410 ( n34936 , n6625 , n31961 );
    or g11411 ( n29267 , n14434 , n8516 );
    and g11412 ( n17239 , n2727 , n24091 );
    not g11413 ( n15039 , n37499 );
    or g11414 ( n12749 , n40995 , n15671 );
    or g11415 ( n14041 , n10200 , n31292 );
    nor g11416 ( n40204 , n6623 , n23186 );
    not g11417 ( n30851 , n2427 );
    nor g11418 ( n11125 , n22947 , n10791 );
    not g11419 ( n31156 , n28269 );
    or g11420 ( n32088 , n8711 , n2125 );
    or g11421 ( n29638 , n23556 , n37952 );
    xnor g11422 ( n31565 , n38749 , n36571 );
    or g11423 ( n7102 , n20921 , n10568 );
    nor g11424 ( n1233 , n6261 , n42259 );
    and g11425 ( n10523 , n32426 , n40508 );
    and g11426 ( n2881 , n27813 , n14156 );
    and g11427 ( n28785 , n23398 , n33421 );
    and g11428 ( n33066 , n36360 , n8580 );
    not g11429 ( n2419 , n30738 );
    or g11430 ( n38602 , n21372 , n28471 );
    or g11431 ( n29366 , n1104 , n5048 );
    not g11432 ( n15860 , n21480 );
    and g11433 ( n4803 , n29301 , n19228 );
    not g11434 ( n11526 , n22342 );
    nor g11435 ( n16827 , n13080 , n15188 );
    nor g11436 ( n11632 , n22521 , n5219 );
    xnor g11437 ( n1349 , n21230 , n19137 );
    or g11438 ( n6265 , n16938 , n31475 );
    and g11439 ( n11821 , n6746 , n38442 );
    or g11440 ( n25002 , n41583 , n29939 );
    not g11441 ( n20921 , n14900 );
    and g11442 ( n1048 , n5738 , n3404 );
    and g11443 ( n2635 , n19611 , n18368 );
    xnor g11444 ( n38246 , n13984 , n41163 );
    nor g11445 ( n7415 , n36486 , n25125 );
    not g11446 ( n20618 , n28496 );
    not g11447 ( n13175 , n27101 );
    and g11448 ( n24255 , n40468 , n35239 );
    and g11449 ( n31364 , n29530 , n24851 );
    xnor g11450 ( n11108 , n5320 , n41420 );
    and g11451 ( n30365 , n41900 , n14444 );
    or g11452 ( n28346 , n13830 , n36492 );
    and g11453 ( n41561 , n25925 , n2986 );
    or g11454 ( n42079 , n41943 , n16785 );
    and g11455 ( n5292 , n32374 , n25301 );
    not g11456 ( n31099 , n38879 );
    or g11457 ( n27597 , n35995 , n22334 );
    not g11458 ( n4535 , n32284 );
    and g11459 ( n15973 , n19148 , n13328 );
    or g11460 ( n35749 , n41526 , n20638 );
    or g11461 ( n7226 , n38019 , n40157 );
    or g11462 ( n22962 , n8447 , n34972 );
    not g11463 ( n40787 , n35221 );
    xnor g11464 ( n24584 , n36009 , n25116 );
    xnor g11465 ( n10417 , n12146 , n41691 );
    xnor g11466 ( n24241 , n36656 , n31980 );
    or g11467 ( n41621 , n14406 , n28837 );
    xnor g11468 ( n29861 , n38081 , n17862 );
    or g11469 ( n22921 , n20597 , n15302 );
    not g11470 ( n25730 , n36426 );
    or g11471 ( n36708 , n18905 , n20265 );
    or g11472 ( n6902 , n2786 , n20687 );
    xnor g11473 ( n28485 , n21937 , n11450 );
    nor g11474 ( n7044 , n27762 , n33129 );
    or g11475 ( n32505 , n420 , n1874 );
    and g11476 ( n9414 , n30396 , n5268 );
    and g11477 ( n34456 , n36135 , n30042 );
    not g11478 ( n26366 , n36298 );
    or g11479 ( n5309 , n24894 , n18101 );
    xnor g11480 ( n35720 , n15972 , n13625 );
    or g11481 ( n24880 , n41650 , n10960 );
    xnor g11482 ( n31017 , n27035 , n21221 );
    and g11483 ( n25888 , n1072 , n42082 );
    or g11484 ( n15059 , n10674 , n38639 );
    or g11485 ( n3609 , n7869 , n2022 );
    or g11486 ( n30289 , n1726 , n16189 );
    or g11487 ( n11491 , n42668 , n17570 );
    or g11488 ( n13870 , n5910 , n30386 );
    not g11489 ( n889 , n35179 );
    and g11490 ( n39902 , n33391 , n7778 );
    nor g11491 ( n26346 , n10542 , n12189 );
    or g11492 ( n35546 , n4108 , n28275 );
    or g11493 ( n24937 , n21855 , n16940 );
    not g11494 ( n32585 , n20793 );
    or g11495 ( n4117 , n4018 , n21828 );
    or g11496 ( n19051 , n33837 , n6289 );
    and g11497 ( n793 , n11982 , n7137 );
    or g11498 ( n38312 , n24626 , n18742 );
    and g11499 ( n36080 , n16274 , n4524 );
    not g11500 ( n24063 , n30322 );
    or g11501 ( n7950 , n4176 , n36651 );
    xnor g11502 ( n8089 , n39852 , n38001 );
    nor g11503 ( n19212 , n19522 , n12306 );
    xnor g11504 ( n25927 , n33884 , n8536 );
    and g11505 ( n24480 , n37221 , n38045 );
    not g11506 ( n13138 , n25570 );
    not g11507 ( n38022 , n4961 );
    xnor g11508 ( n32572 , n12057 , n9159 );
    not g11509 ( n20904 , n38263 );
    not g11510 ( n31087 , n23882 );
    or g11511 ( n10389 , n33926 , n30493 );
    not g11512 ( n29310 , n20544 );
    and g11513 ( n5444 , n6823 , n14456 );
    xnor g11514 ( n42140 , n14942 , n18445 );
    or g11515 ( n30157 , n15013 , n4301 );
    or g11516 ( n18457 , n32245 , n36931 );
    nor g11517 ( n36722 , n33098 , n3894 );
    not g11518 ( n10491 , n14888 );
    nor g11519 ( n23614 , n11460 , n25356 );
    or g11520 ( n29191 , n3034 , n40568 );
    or g11521 ( n38247 , n1995 , n9466 );
    nor g11522 ( n38231 , n13476 , n14966 );
    nor g11523 ( n34469 , n6640 , n21963 );
    xnor g11524 ( n42815 , n20467 , n17917 );
    and g11525 ( n26280 , n12857 , n10895 );
    or g11526 ( n17521 , n17750 , n10849 );
    nor g11527 ( n13547 , n8494 , n31664 );
    xnor g11528 ( n20008 , n35553 , n42225 );
    nor g11529 ( n25104 , n33981 , n14126 );
    not g11530 ( n25811 , n28584 );
    or g11531 ( n29959 , n35175 , n29708 );
    xnor g11532 ( n3179 , n21973 , n31911 );
    or g11533 ( n30962 , n33926 , n17065 );
    nor g11534 ( n1799 , n12004 , n35634 );
    or g11535 ( n28024 , n30488 , n32666 );
    xnor g11536 ( n35858 , n28983 , n12608 );
    or g11537 ( n30276 , n38022 , n7189 );
    nor g11538 ( n3320 , n5896 , n21481 );
    nor g11539 ( n32952 , n30166 , n33272 );
    or g11540 ( n16453 , n38492 , n34609 );
    not g11541 ( n18672 , n35971 );
    or g11542 ( n37967 , n36848 , n11044 );
    and g11543 ( n37978 , n19557 , n5050 );
    and g11544 ( n39168 , n38738 , n41593 );
    not g11545 ( n27738 , n10307 );
    or g11546 ( n5749 , n10898 , n2715 );
    not g11547 ( n18511 , n2406 );
    or g11548 ( n38386 , n8870 , n1861 );
    not g11549 ( n28867 , n19861 );
    or g11550 ( n38888 , n37722 , n31153 );
    not g11551 ( n36843 , n17489 );
    and g11552 ( n30451 , n27656 , n32805 );
    and g11553 ( n6053 , n16526 , n40528 );
    nor g11554 ( n6779 , n32506 , n35418 );
    and g11555 ( n10180 , n7387 , n17125 );
    and g11556 ( n853 , n23688 , n9148 );
    nor g11557 ( n22789 , n31989 , n20178 );
    not g11558 ( n12130 , n14712 );
    not g11559 ( n9667 , n28971 );
    nor g11560 ( n14283 , n19903 , n20103 );
    or g11561 ( n34313 , n23951 , n38150 );
    xnor g11562 ( n22382 , n10414 , n42185 );
    nor g11563 ( n26052 , n23861 , n24455 );
    and g11564 ( n24662 , n5836 , n41751 );
    or g11565 ( n13435 , n23487 , n15894 );
    not g11566 ( n13566 , n37446 );
    not g11567 ( n20978 , n25910 );
    xnor g11568 ( n40017 , n10774 , n32665 );
    or g11569 ( n17266 , n31810 , n11915 );
    or g11570 ( n30181 , n31451 , n26174 );
    not g11571 ( n37122 , n28833 );
    nor g11572 ( n36220 , n38640 , n33562 );
    or g11573 ( n23927 , n22314 , n27273 );
    or g11574 ( n8246 , n20269 , n644 );
    and g11575 ( n13752 , n35147 , n29119 );
    and g11576 ( n32435 , n105 , n8630 );
    and g11577 ( n5800 , n24116 , n8652 );
    not g11578 ( n26972 , n28404 );
    not g11579 ( n28870 , n34482 );
    xnor g11580 ( n14313 , n4857 , n5596 );
    not g11581 ( n34536 , n36688 );
    not g11582 ( n42694 , n263 );
    or g11583 ( n38455 , n28009 , n9935 );
    not g11584 ( n19728 , n4834 );
    or g11585 ( n48 , n13830 , n23589 );
    and g11586 ( n24816 , n16519 , n1784 );
    xnor g11587 ( n4927 , n36423 , n42171 );
    and g11588 ( n25360 , n5442 , n41465 );
    or g11589 ( n13208 , n20156 , n30610 );
    or g11590 ( n32737 , n40312 , n15064 );
    and g11591 ( n8927 , n42696 , n6034 );
    or g11592 ( n20339 , n6000 , n6342 );
    not g11593 ( n19645 , n34990 );
    not g11594 ( n9160 , n30555 );
    xnor g11595 ( n36690 , n38694 , n29342 );
    nor g11596 ( n39552 , n37797 , n25797 );
    or g11597 ( n31327 , n3014 , n29554 );
    and g11598 ( n31373 , n24587 , n25586 );
    or g11599 ( n27336 , n18785 , n20827 );
    or g11600 ( n23534 , n2420 , n40678 );
    or g11601 ( n9611 , n22619 , n30199 );
    xnor g11602 ( n36140 , n22753 , n30933 );
    not g11603 ( n39443 , n36060 );
    or g11604 ( n8393 , n35843 , n13282 );
    xnor g11605 ( n9573 , n21145 , n35962 );
    and g11606 ( n24723 , n27441 , n35996 );
    or g11607 ( n23737 , n34728 , n33728 );
    xnor g11608 ( n34848 , n5891 , n32494 );
    xnor g11609 ( n33251 , n16742 , n27444 );
    xnor g11610 ( n37218 , n25388 , n26660 );
    and g11611 ( n33171 , n34731 , n32435 );
    xnor g11612 ( n32463 , n1255 , n34074 );
    xnor g11613 ( n15110 , n9180 , n33293 );
    nor g11614 ( n2308 , n9880 , n27910 );
    or g11615 ( n26009 , n40318 , n20058 );
    or g11616 ( n29393 , n30230 , n31879 );
    not g11617 ( n37444 , n28076 );
    xnor g11618 ( n33827 , n36158 , n1971 );
    and g11619 ( n12120 , n31172 , n42325 );
    nor g11620 ( n9383 , n31124 , n35395 );
    or g11621 ( n32641 , n17256 , n28737 );
    not g11622 ( n22695 , n31975 );
    or g11623 ( n32648 , n42508 , n11294 );
    or g11624 ( n10501 , n29615 , n7220 );
    and g11625 ( n11769 , n36175 , n5425 );
    and g11626 ( n38074 , n26247 , n13679 );
    nor g11627 ( n30458 , n18866 , n18485 );
    not g11628 ( n21332 , n19407 );
    nor g11629 ( n8023 , n28749 , n21337 );
    or g11630 ( n36768 , n32728 , n27085 );
    nor g11631 ( n30780 , n34565 , n37510 );
    or g11632 ( n25972 , n17320 , n10890 );
    or g11633 ( n39341 , n7142 , n23764 );
    or g11634 ( n25045 , n19913 , n25935 );
    or g11635 ( n5644 , n29833 , n42766 );
    or g11636 ( n6689 , n32411 , n1788 );
    or g11637 ( n749 , n15149 , n8631 );
    xnor g11638 ( n19681 , n39279 , n9299 );
    or g11639 ( n20984 , n20634 , n21772 );
    xnor g11640 ( n28791 , n1956 , n14707 );
    nor g11641 ( n1345 , n26418 , n18537 );
    or g11642 ( n42438 , n29027 , n1251 );
    xnor g11643 ( n31616 , n40064 , n7403 );
    nor g11644 ( n6827 , n5964 , n6006 );
    or g11645 ( n25569 , n2012 , n4094 );
    nor g11646 ( n27375 , n24105 , n28089 );
    or g11647 ( n6540 , n26787 , n39647 );
    or g11648 ( n9288 , n30975 , n19535 );
    xnor g11649 ( n32865 , n27907 , n24363 );
    or g11650 ( n15664 , n21703 , n23313 );
    or g11651 ( n41828 , n34429 , n24635 );
    and g11652 ( n10901 , n12146 , n26579 );
    or g11653 ( n38178 , n5896 , n40232 );
    or g11654 ( n36581 , n36079 , n4401 );
    and g11655 ( n27947 , n2546 , n38848 );
    xnor g11656 ( n33193 , n20161 , n17912 );
    not g11657 ( n25443 , n905 );
    nor g11658 ( n30714 , n30563 , n9340 );
    xnor g11659 ( n11277 , n41013 , n31779 );
    xnor g11660 ( n10347 , n3146 , n13493 );
    xnor g11661 ( n150 , n2214 , n39299 );
    nor g11662 ( n21913 , n19174 , n3895 );
    or g11663 ( n42254 , n40295 , n23651 );
    xnor g11664 ( n212 , n29476 , n18121 );
    not g11665 ( n12630 , n3898 );
    or g11666 ( n4251 , n38157 , n12610 );
    not g11667 ( n38847 , n10465 );
    or g11668 ( n17331 , n35301 , n14695 );
    nor g11669 ( n18971 , n7870 , n38088 );
    and g11670 ( n25213 , n13977 , n16317 );
    and g11671 ( n11122 , n13240 , n32306 );
    or g11672 ( n3914 , n30496 , n13019 );
    nor g11673 ( n23320 , n13151 , n13815 );
    or g11674 ( n10572 , n15040 , n15722 );
    or g11675 ( n34435 , n7065 , n14074 );
    not g11676 ( n25526 , n8274 );
    or g11677 ( n12013 , n37680 , n5910 );
    and g11678 ( n35032 , n9921 , n17168 );
    or g11679 ( n24757 , n5881 , n26314 );
    or g11680 ( n36059 , n39367 , n31619 );
    xnor g11681 ( n9495 , n42917 , n4390 );
    or g11682 ( n7192 , n40289 , n34536 );
    xnor g11683 ( n19605 , n6565 , n21753 );
    xnor g11684 ( n4986 , n37969 , n6848 );
    or g11685 ( n42718 , n6458 , n29449 );
    or g11686 ( n3383 , n9697 , n6250 );
    and g11687 ( n19781 , n26509 , n39335 );
    xnor g11688 ( n22110 , n2722 , n29615 );
    nor g11689 ( n21325 , n27808 , n38919 );
    nor g11690 ( n31919 , n35352 , n10575 );
    not g11691 ( n3218 , n2494 );
    and g11692 ( n30547 , n10343 , n17607 );
    nor g11693 ( n31801 , n33190 , n36205 );
    nor g11694 ( n33849 , n15070 , n14245 );
    and g11695 ( n18075 , n21769 , n4614 );
    and g11696 ( n26887 , n17675 , n28975 );
    not g11697 ( n20531 , n4480 );
    and g11698 ( n7482 , n13870 , n26457 );
    nor g11699 ( n22882 , n8904 , n16178 );
    or g11700 ( n14241 , n11232 , n38618 );
    or g11701 ( n22576 , n16740 , n9004 );
    not g11702 ( n42446 , n11900 );
    and g11703 ( n6413 , n30758 , n20002 );
    not g11704 ( n23859 , n25624 );
    or g11705 ( n39880 , n29983 , n14917 );
    and g11706 ( n41625 , n5464 , n15945 );
    and g11707 ( n9569 , n34794 , n10188 );
    xnor g11708 ( n8058 , n40 , n5673 );
    not g11709 ( n42591 , n22864 );
    and g11710 ( n11645 , n16307 , n26322 );
    and g11711 ( n4206 , n3151 , n42861 );
    or g11712 ( n24274 , n39127 , n12199 );
    or g11713 ( n31960 , n22631 , n10599 );
    or g11714 ( n5388 , n34234 , n20814 );
    xnor g11715 ( n16015 , n31956 , n1648 );
    and g11716 ( n28691 , n42482 , n24959 );
    or g11717 ( n32022 , n4869 , n24006 );
    or g11718 ( n2528 , n24035 , n14108 );
    or g11719 ( n35458 , n30700 , n27241 );
    xnor g11720 ( n23165 , n38269 , n14664 );
    nor g11721 ( n5471 , n28174 , n2902 );
    and g11722 ( n9851 , n38741 , n3575 );
    or g11723 ( n6395 , n23489 , n225 );
    xnor g11724 ( n18067 , n16693 , n34828 );
    and g11725 ( n38931 , n42275 , n34369 );
    xnor g11726 ( n7254 , n3607 , n33246 );
    and g11727 ( n3517 , n34200 , n6205 );
    or g11728 ( n31289 , n33330 , n32332 );
    or g11729 ( n39431 , n28988 , n3649 );
    nor g11730 ( n36597 , n42056 , n42718 );
    xnor g11731 ( n33178 , n18061 , n33906 );
    and g11732 ( n4936 , n11850 , n28606 );
    xnor g11733 ( n12969 , n15842 , n18078 );
    not g11734 ( n20553 , n2832 );
    xnor g11735 ( n23716 , n19665 , n29076 );
    and g11736 ( n30970 , n17050 , n41973 );
    not g11737 ( n4129 , n1549 );
    xnor g11738 ( n36909 , n31127 , n14471 );
    nor g11739 ( n34016 , n11578 , n24111 );
    or g11740 ( n12624 , n30614 , n11312 );
    xnor g11741 ( n8729 , n34444 , n31914 );
    and g11742 ( n36038 , n17809 , n33076 );
    xnor g11743 ( n29085 , n34731 , n5663 );
    not g11744 ( n18749 , n691 );
    xnor g11745 ( n11676 , n4351 , n10970 );
    or g11746 ( n18493 , n29349 , n25392 );
    or g11747 ( n26762 , n35185 , n3689 );
    and g11748 ( n18394 , n40362 , n30991 );
    xnor g11749 ( n32910 , n42064 , n5863 );
    not g11750 ( n40160 , n10264 );
    xnor g11751 ( n28073 , n38749 , n41361 );
    nor g11752 ( n29690 , n8494 , n13244 );
    and g11753 ( n17360 , n36927 , n20121 );
    xnor g11754 ( n7626 , n12536 , n7261 );
    xnor g11755 ( n33544 , n6552 , n7570 );
    and g11756 ( n13066 , n40613 , n4628 );
    and g11757 ( n25179 , n38171 , n32314 );
    and g11758 ( n40319 , n11103 , n15834 );
    nor g11759 ( n30223 , n36911 , n18883 );
    not g11760 ( n15165 , n20927 );
    and g11761 ( n39296 , n17080 , n33062 );
    or g11762 ( n3121 , n38255 , n4301 );
    or g11763 ( n5815 , n2302 , n16603 );
    or g11764 ( n25908 , n22778 , n39911 );
    and g11765 ( n20215 , n42417 , n39725 );
    or g11766 ( n3509 , n14388 , n25361 );
    or g11767 ( n10543 , n41327 , n11134 );
    or g11768 ( n17348 , n4098 , n40245 );
    not g11769 ( n32602 , n10347 );
    or g11770 ( n35943 , n12808 , n388 );
    or g11771 ( n17261 , n866 , n177 );
    xnor g11772 ( n17571 , n28612 , n13514 );
    and g11773 ( n27119 , n28109 , n40555 );
    or g11774 ( n14102 , n6418 , n42425 );
    xnor g11775 ( n19245 , n35217 , n15547 );
    not g11776 ( n3982 , n23379 );
    nor g11777 ( n18294 , n34565 , n11036 );
    or g11778 ( n11802 , n21625 , n42667 );
    xnor g11779 ( n37240 , n10078 , n25928 );
    or g11780 ( n10203 , n18690 , n13745 );
    nor g11781 ( n17253 , n5203 , n40876 );
    or g11782 ( n28582 , n7045 , n8270 );
    not g11783 ( n18881 , n39212 );
    or g11784 ( n11172 , n12685 , n38662 );
    not g11785 ( n1838 , n37811 );
    or g11786 ( n9102 , n10561 , n14668 );
    and g11787 ( n32319 , n9013 , n4457 );
    not g11788 ( n30682 , n15998 );
    not g11789 ( n10639 , n2857 );
    not g11790 ( n25706 , n39310 );
    nor g11791 ( n8978 , n5826 , n35739 );
    not g11792 ( n27025 , n29253 );
    or g11793 ( n16344 , n18116 , n2761 );
    and g11794 ( n1578 , n26014 , n39192 );
    or g11795 ( n31209 , n23849 , n41870 );
    or g11796 ( n538 , n32341 , n12140 );
    xnor g11797 ( n4244 , n25619 , n37332 );
    or g11798 ( n33206 , n17382 , n5850 );
    and g11799 ( n3333 , n24347 , n22922 );
    or g11800 ( n1492 , n15055 , n9239 );
    nor g11801 ( n7885 , n35748 , n20069 );
    and g11802 ( n34577 , n36674 , n41091 );
    and g11803 ( n17514 , n22173 , n17343 );
    or g11804 ( n14460 , n3434 , n16891 );
    nor g11805 ( n19480 , n3502 , n31403 );
    and g11806 ( n6859 , n5306 , n6897 );
    and g11807 ( n724 , n42662 , n224 );
    or g11808 ( n35502 , n14069 , n22219 );
    nor g11809 ( n30239 , n22625 , n35662 );
    xnor g11810 ( n4609 , n12693 , n39667 );
    not g11811 ( n9090 , n42096 );
    and g11812 ( n23011 , n21236 , n23143 );
    or g11813 ( n29286 , n23509 , n11113 );
    not g11814 ( n27766 , n33927 );
    or g11815 ( n24433 , n26988 , n2599 );
    not g11816 ( n35743 , n14340 );
    not g11817 ( n12129 , n24221 );
    nor g11818 ( n11222 , n18732 , n38709 );
    nor g11819 ( n24267 , n40472 , n34287 );
    or g11820 ( n25930 , n42655 , n18035 );
    and g11821 ( n17473 , n13588 , n23677 );
    and g11822 ( n5628 , n22527 , n42795 );
    or g11823 ( n17093 , n10598 , n29368 );
    and g11824 ( n39639 , n9090 , n32906 );
    or g11825 ( n42354 , n28673 , n41997 );
    and g11826 ( n20889 , n14968 , n19202 );
    xnor g11827 ( n38667 , n34875 , n27936 );
    nor g11828 ( n11745 , n39778 , n4484 );
    and g11829 ( n32951 , n24891 , n22384 );
    or g11830 ( n9477 , n6231 , n12153 );
    xnor g11831 ( n536 , n27334 , n40527 );
    not g11832 ( n37763 , n26142 );
    xnor g11833 ( n42117 , n34562 , n41528 );
    or g11834 ( n13399 , n17485 , n18763 );
    not g11835 ( n23052 , n21931 );
    or g11836 ( n19741 , n25126 , n10974 );
    nor g11837 ( n33320 , n35074 , n34135 );
    or g11838 ( n31814 , n24062 , n3556 );
    not g11839 ( n30837 , n770 );
    not g11840 ( n29489 , n23766 );
    xnor g11841 ( n3805 , n12605 , n39974 );
    or g11842 ( n1545 , n23971 , n36072 );
    nor g11843 ( n38384 , n22822 , n39070 );
    or g11844 ( n21202 , n7668 , n28324 );
    and g11845 ( n14493 , n41450 , n4000 );
    xnor g11846 ( n23310 , n40939 , n2955 );
    xnor g11847 ( n21525 , n15972 , n9912 );
    or g11848 ( n18965 , n25600 , n22411 );
    and g11849 ( n35127 , n3239 , n28112 );
    and g11850 ( n24602 , n42589 , n26771 );
    nor g11851 ( n28210 , n8157 , n40023 );
    or g11852 ( n19745 , n27205 , n14275 );
    nor g11853 ( n29549 , n35965 , n8294 );
    or g11854 ( n29417 , n27624 , n32744 );
    or g11855 ( n19492 , n41667 , n10490 );
    not g11856 ( n3732 , n23099 );
    nor g11857 ( n15227 , n20067 , n11647 );
    or g11858 ( n22435 , n14379 , n21060 );
    or g11859 ( n7126 , n2197 , n9217 );
    xnor g11860 ( n3172 , n13769 , n22568 );
    not g11861 ( n14308 , n32056 );
    nor g11862 ( n19473 , n26612 , n7521 );
    and g11863 ( n8083 , n7871 , n12838 );
    and g11864 ( n29742 , n8446 , n37974 );
    and g11865 ( n8429 , n21003 , n13763 );
    xnor g11866 ( n7678 , n28113 , n25588 );
    not g11867 ( n27654 , n36863 );
    or g11868 ( n5249 , n40366 , n13637 );
    or g11869 ( n26457 , n29600 , n30561 );
    or g11870 ( n26683 , n37944 , n1620 );
    or g11871 ( n10775 , n38157 , n38257 );
    and g11872 ( n16440 , n31078 , n34867 );
    and g11873 ( n42114 , n19413 , n7231 );
    and g11874 ( n3886 , n3474 , n11029 );
    or g11875 ( n16477 , n17848 , n12759 );
    and g11876 ( n28780 , n35108 , n27215 );
    not g11877 ( n41623 , n13409 );
    or g11878 ( n5735 , n13701 , n33502 );
    or g11879 ( n18810 , n33655 , n16325 );
    and g11880 ( n8926 , n26521 , n16171 );
    not g11881 ( n7621 , n25607 );
    xnor g11882 ( n16 , n20245 , n555 );
    not g11883 ( n38155 , n25838 );
    or g11884 ( n1798 , n13492 , n7331 );
    nor g11885 ( n39493 , n18215 , n17621 );
    or g11886 ( n26006 , n35368 , n5850 );
    nor g11887 ( n9665 , n1507 , n18703 );
    xnor g11888 ( n33310 , n21133 , n30715 );
    not g11889 ( n4873 , n20714 );
    or g11890 ( n38361 , n42039 , n4642 );
    or g11891 ( n32523 , n10878 , n29884 );
    and g11892 ( n39429 , n28090 , n22332 );
    or g11893 ( n25898 , n33311 , n5252 );
    or g11894 ( n10218 , n3835 , n12477 );
    or g11895 ( n29995 , n37664 , n28113 );
    xnor g11896 ( n29567 , n38105 , n21650 );
    or g11897 ( n2568 , n12286 , n23463 );
    and g11898 ( n35838 , n26568 , n14221 );
    nor g11899 ( n31345 , n2194 , n2822 );
    nor g11900 ( n1949 , n13336 , n35859 );
    and g11901 ( n20205 , n21447 , n23135 );
    or g11902 ( n14604 , n24341 , n3543 );
    not g11903 ( n29857 , n26344 );
    or g11904 ( n19205 , n27678 , n10095 );
    and g11905 ( n12509 , n13611 , n30594 );
    or g11906 ( n2778 , n17204 , n22445 );
    and g11907 ( n35530 , n27 , n15554 );
    or g11908 ( n34092 , n18798 , n9207 );
    or g11909 ( n12854 , n26226 , n10113 );
    nor g11910 ( n20578 , n38563 , n117 );
    xnor g11911 ( n18925 , n4573 , n24654 );
    and g11912 ( n3155 , n16606 , n26328 );
    or g11913 ( n26042 , n11445 , n20175 );
    and g11914 ( n40561 , n26067 , n28810 );
    or g11915 ( n18923 , n11327 , n2426 );
    xnor g11916 ( n30724 , n5144 , n10385 );
    and g11917 ( n42580 , n30657 , n39756 );
    nor g11918 ( n40821 , n10480 , n25368 );
    xnor g11919 ( n6067 , n31848 , n15960 );
    nor g11920 ( n39959 , n18401 , n4066 );
    or g11921 ( n26798 , n404 , n13064 );
    and g11922 ( n18710 , n17533 , n11191 );
    nor g11923 ( n30294 , n27754 , n11503 );
    or g11924 ( n34870 , n41823 , n11814 );
    and g11925 ( n13317 , n7865 , n1787 );
    xnor g11926 ( n28296 , n27704 , n39294 );
    and g11927 ( n1058 , n11437 , n594 );
    and g11928 ( n22564 , n15845 , n16240 );
    not g11929 ( n27396 , n7673 );
    not g11930 ( n32217 , n12318 );
    nor g11931 ( n16284 , n10598 , n8418 );
    nor g11932 ( n29273 , n30281 , n3214 );
    and g11933 ( n3564 , n37504 , n36442 );
    or g11934 ( n28142 , n31950 , n35734 );
    xnor g11935 ( n18208 , n42847 , n4201 );
    xnor g11936 ( n24940 , n14596 , n28348 );
    or g11937 ( n31959 , n20819 , n3838 );
    or g11938 ( n33477 , n4274 , n27903 );
    and g11939 ( n32489 , n17945 , n18913 );
    nor g11940 ( n28754 , n16573 , n10028 );
    and g11941 ( n20570 , n17558 , n18565 );
    or g11942 ( n28280 , n23782 , n4056 );
    nor g11943 ( n36991 , n40067 , n1995 );
    or g11944 ( n2321 , n34854 , n13071 );
    and g11945 ( n4646 , n36345 , n35993 );
    and g11946 ( n23530 , n28000 , n10368 );
    or g11947 ( n25763 , n2533 , n8514 );
    or g11948 ( n36874 , n30002 , n17109 );
    not g11949 ( n31694 , n2093 );
    nor g11950 ( n9359 , n19221 , n34229 );
    nor g11951 ( n19736 , n25917 , n8908 );
    nor g11952 ( n40663 , n34103 , n17196 );
    and g11953 ( n38176 , n24477 , n22148 );
    not g11954 ( n12302 , n38004 );
    or g11955 ( n29870 , n40073 , n6794 );
    and g11956 ( n11786 , n23723 , n17733 );
    or g11957 ( n35056 , n36299 , n24560 );
    or g11958 ( n10933 , n32800 , n40602 );
    and g11959 ( n20381 , n37449 , n19717 );
    or g11960 ( n31305 , n29455 , n36550 );
    nor g11961 ( n30401 , n22317 , n31013 );
    or g11962 ( n36460 , n2368 , n42730 );
    and g11963 ( n24396 , n26565 , n27807 );
    and g11964 ( n11737 , n6773 , n32456 );
    or g11965 ( n38221 , n9191 , n7604 );
    or g11966 ( n10059 , n9748 , n18055 );
    not g11967 ( n6671 , n27764 );
    nor g11968 ( n23492 , n7572 , n12352 );
    nor g11969 ( n17160 , n20994 , n42303 );
    or g11970 ( n41068 , n12706 , n14680 );
    xnor g11971 ( n41407 , n34691 , n42173 );
    nor g11972 ( n26851 , n34816 , n457 );
    and g11973 ( n35331 , n29456 , n13638 );
    nor g11974 ( n33669 , n42064 , n29168 );
    not g11975 ( n11344 , n27141 );
    nor g11976 ( n29192 , n5073 , n19858 );
    or g11977 ( n29710 , n19333 , n42694 );
    not g11978 ( n18722 , n38514 );
    and g11979 ( n8542 , n19316 , n41372 );
    and g11980 ( n36865 , n34731 , n23270 );
    nor g11981 ( n14470 , n41859 , n28991 );
    nor g11982 ( n24387 , n23011 , n27954 );
    or g11983 ( n12792 , n1503 , n27127 );
    and g11984 ( n2791 , n32334 , n18693 );
    and g11985 ( n40697 , n32567 , n5107 );
    nor g11986 ( n37282 , n3776 , n26339 );
    or g11987 ( n13038 , n287 , n7034 );
    not g11988 ( n21551 , n36313 );
    xnor g11989 ( n33526 , n26627 , n13568 );
    xnor g11990 ( n25571 , n40391 , n25583 );
    and g11991 ( n22671 , n27381 , n6531 );
    or g11992 ( n23885 , n35101 , n40639 );
    and g11993 ( n42751 , n30535 , n30245 );
    and g11994 ( n31625 , n24032 , n16749 );
    not g11995 ( n29113 , n13720 );
    nor g11996 ( n30968 , n20074 , n1786 );
    or g11997 ( n26400 , n38864 , n13566 );
    not g11998 ( n40673 , n11297 );
    not g11999 ( n16267 , n26201 );
    xnor g12000 ( n14353 , n32672 , n27946 );
    xnor g12001 ( n20055 , n39178 , n36733 );
    or g12002 ( n3990 , n34686 , n17022 );
    not g12003 ( n28159 , n13445 );
    or g12004 ( n26738 , n17736 , n9702 );
    or g12005 ( n30104 , n41036 , n34436 );
    xnor g12006 ( n21733 , n22263 , n25669 );
    and g12007 ( n23043 , n30675 , n7440 );
    or g12008 ( n33016 , n39537 , n21849 );
    xnor g12009 ( n29319 , n9767 , n34565 );
    not g12010 ( n4642 , n24866 );
    not g12011 ( n39065 , n570 );
    or g12012 ( n33369 , n9031 , n22076 );
    or g12013 ( n5381 , n7649 , n4843 );
    not g12014 ( n37610 , n3119 );
    and g12015 ( n39984 , n37236 , n18374 );
    nor g12016 ( n37598 , n21199 , n24450 );
    nor g12017 ( n37404 , n15070 , n22021 );
    and g12018 ( n27551 , n21181 , n1476 );
    or g12019 ( n15819 , n3420 , n1740 );
    nor g12020 ( n6472 , n34651 , n23876 );
    or g12021 ( n24523 , n40294 , n28837 );
    not g12022 ( n5988 , n38372 );
    or g12023 ( n27386 , n4751 , n29147 );
    xnor g12024 ( n11403 , n10456 , n27330 );
    nor g12025 ( n10002 , n8656 , n4098 );
    or g12026 ( n30054 , n40265 , n272 );
    or g12027 ( n33890 , n41366 , n38814 );
    nor g12028 ( n2754 , n22010 , n27742 );
    not g12029 ( n26490 , n23048 );
    and g12030 ( n30601 , n36761 , n10452 );
    nor g12031 ( n36428 , n14231 , n5562 );
    not g12032 ( n19562 , n1582 );
    nor g12033 ( n40699 , n31791 , n41351 );
    not g12034 ( n17850 , n34886 );
    or g12035 ( n32266 , n21064 , n13622 );
    and g12036 ( n24365 , n31840 , n32838 );
    or g12037 ( n720 , n19858 , n33655 );
    nor g12038 ( n38443 , n7266 , n28317 );
    and g12039 ( n18086 , n28925 , n35698 );
    or g12040 ( n22190 , n25682 , n1658 );
    and g12041 ( n20893 , n42104 , n10621 );
    nor g12042 ( n30491 , n1507 , n34132 );
    or g12043 ( n15383 , n11049 , n26493 );
    or g12044 ( n17068 , n18431 , n10450 );
    xnor g12045 ( n11217 , n31607 , n25309 );
    xnor g12046 ( n6542 , n35876 , n40894 );
    xnor g12047 ( n20677 , n22698 , n33086 );
    and g12048 ( n29065 , n28227 , n38656 );
    not g12049 ( n6885 , n31694 );
    or g12050 ( n33613 , n32589 , n14913 );
    nor g12051 ( n40865 , n36117 , n924 );
    and g12052 ( n42096 , n27394 , n3243 );
    or g12053 ( n764 , n17744 , n37056 );
    xnor g12054 ( n15099 , n31539 , n29752 );
    or g12055 ( n36006 , n16599 , n9411 );
    and g12056 ( n6411 , n40208 , n10807 );
    or g12057 ( n8671 , n2382 , n30820 );
    or g12058 ( n2103 , n13848 , n29110 );
    nor g12059 ( n13369 , n35512 , n34786 );
    and g12060 ( n4307 , n24933 , n32306 );
    or g12061 ( n31701 , n37270 , n24643 );
    not g12062 ( n17722 , n28755 );
    and g12063 ( n27260 , n26410 , n3177 );
    and g12064 ( n2556 , n36354 , n19047 );
    or g12065 ( n7055 , n6180 , n29798 );
    not g12066 ( n24745 , n426 );
    not g12067 ( n32078 , n13144 );
    or g12068 ( n34111 , n14980 , n35443 );
    xnor g12069 ( n13897 , n37914 , n430 );
    and g12070 ( n33293 , n42012 , n17565 );
    or g12071 ( n25662 , n20741 , n36757 );
    or g12072 ( n27556 , n22478 , n15631 );
    or g12073 ( n40969 , n5225 , n16783 );
    and g12074 ( n22589 , n40622 , n28043 );
    or g12075 ( n16638 , n7288 , n32980 );
    and g12076 ( n18575 , n20785 , n21971 );
    or g12077 ( n25975 , n39258 , n7802 );
    or g12078 ( n9759 , n30653 , n41079 );
    or g12079 ( n17557 , n42158 , n40016 );
    or g12080 ( n10708 , n16718 , n25119 );
    nor g12081 ( n6717 , n532 , n4827 );
    or g12082 ( n6766 , n29593 , n9406 );
    and g12083 ( n22823 , n10083 , n39467 );
    or g12084 ( n7206 , n29013 , n11346 );
    xnor g12085 ( n10396 , n18606 , n34292 );
    and g12086 ( n23558 , n34312 , n29734 );
    or g12087 ( n42720 , n20288 , n26956 );
    and g12088 ( n24653 , n16180 , n34620 );
    not g12089 ( n32716 , n4517 );
    or g12090 ( n36698 , n35818 , n16216 );
    or g12091 ( n37619 , n13701 , n35539 );
    xnor g12092 ( n21244 , n10612 , n38909 );
    or g12093 ( n42663 , n24633 , n21926 );
    xnor g12094 ( n40183 , n35887 , n2432 );
    or g12095 ( n34394 , n32217 , n25546 );
    and g12096 ( n40732 , n37940 , n41785 );
    nor g12097 ( n14545 , n14786 , n34355 );
    or g12098 ( n27300 , n22371 , n25686 );
    not g12099 ( n5423 , n25046 );
    or g12100 ( n8174 , n17772 , n5978 );
    nor g12101 ( n31632 , n6565 , n37628 );
    or g12102 ( n1888 , n10244 , n37384 );
    or g12103 ( n41880 , n33738 , n24068 );
    or g12104 ( n31112 , n2848 , n32563 );
    nor g12105 ( n26559 , n3837 , n39184 );
    or g12106 ( n34438 , n8432 , n37768 );
    nor g12107 ( n17092 , n32495 , n35691 );
    or g12108 ( n8185 , n2977 , n33671 );
    nor g12109 ( n17262 , n36539 , n34720 );
    or g12110 ( n42503 , n31452 , n31136 );
    or g12111 ( n12798 , n862 , n1641 );
    or g12112 ( n26413 , n40748 , n11262 );
    and g12113 ( n5989 , n34629 , n29576 );
    xnor g12114 ( n8796 , n4123 , n35744 );
    and g12115 ( n41420 , n2033 , n5511 );
    xnor g12116 ( n11293 , n9155 , n29898 );
    or g12117 ( n5460 , n425 , n39634 );
    not g12118 ( n34933 , n17131 );
    and g12119 ( n34537 , n22019 , n42397 );
    not g12120 ( n27171 , n26581 );
    or g12121 ( n29758 , n33423 , n23056 );
    or g12122 ( n795 , n1693 , n9026 );
    not g12123 ( n33636 , n5289 );
    and g12124 ( n19235 , n12297 , n9786 );
    not g12125 ( n8888 , n16348 );
    nor g12126 ( n19838 , n37729 , n4734 );
    and g12127 ( n15371 , n15153 , n40394 );
    or g12128 ( n25855 , n1507 , n23968 );
    or g12129 ( n18852 , n23858 , n36235 );
    and g12130 ( n653 , n9101 , n29116 );
    nor g12131 ( n24173 , n130 , n11758 );
    nor g12132 ( n26986 , n13936 , n33009 );
    and g12133 ( n34037 , n12584 , n24811 );
    nor g12134 ( n2711 , n23067 , n9883 );
    or g12135 ( n23699 , n42870 , n25851 );
    nor g12136 ( n38009 , n35790 , n28495 );
    or g12137 ( n25541 , n23971 , n35232 );
    or g12138 ( n18396 , n333 , n1678 );
    or g12139 ( n30427 , n14471 , n35258 );
    not g12140 ( n29432 , n34677 );
    nor g12141 ( n38517 , n7777 , n24869 );
    not g12142 ( n37521 , n20929 );
    or g12143 ( n25196 , n5848 , n6262 );
    not g12144 ( n20322 , n20792 );
    xnor g12145 ( n3881 , n12156 , n16199 );
    and g12146 ( n15377 , n36598 , n33426 );
    or g12147 ( n4475 , n13775 , n25507 );
    not g12148 ( n35009 , n1572 );
    nor g12149 ( n32439 , n14188 , n36091 );
    or g12150 ( n8818 , n35273 , n18236 );
    and g12151 ( n5426 , n34859 , n41093 );
    not g12152 ( n40032 , n14968 );
    not g12153 ( n8004 , n37094 );
    or g12154 ( n27166 , n27037 , n35849 );
    nor g12155 ( n39197 , n5650 , n17442 );
    or g12156 ( n2275 , n13357 , n6543 );
    or g12157 ( n42120 , n17193 , n28633 );
    nor g12158 ( n31061 , n18550 , n1286 );
    or g12159 ( n12343 , n19009 , n20370 );
    or g12160 ( n21713 , n34685 , n19701 );
    and g12161 ( n5513 , n26324 , n29956 );
    not g12162 ( n9808 , n26593 );
    xnor g12163 ( n15056 , n11785 , n41927 );
    or g12164 ( n12941 , n2104 , n10559 );
    nor g12165 ( n13658 , n18275 , n36279 );
    nor g12166 ( n8244 , n21621 , n37522 );
    xnor g12167 ( n11442 , n35727 , n5518 );
    nor g12168 ( n13220 , n6179 , n39152 );
    or g12169 ( n33916 , n28534 , n26590 );
    or g12170 ( n17899 , n23085 , n26708 );
    not g12171 ( n25657 , n26114 );
    not g12172 ( n1884 , n12273 );
    or g12173 ( n14662 , n41207 , n13594 );
    or g12174 ( n21707 , n23598 , n20179 );
    and g12175 ( n18000 , n39114 , n25450 );
    or g12176 ( n13246 , n12582 , n8658 );
    or g12177 ( n17408 , n39312 , n4421 );
    nor g12178 ( n34995 , n28664 , n31204 );
    nor g12179 ( n2739 , n30761 , n15587 );
    and g12180 ( n17401 , n20840 , n34763 );
    xnor g12181 ( n5015 , n36009 , n2556 );
    xnor g12182 ( n24111 , n41358 , n12056 );
    and g12183 ( n18485 , n8452 , n23633 );
    nor g12184 ( n21760 , n25187 , n19114 );
    xnor g12185 ( n39045 , n4334 , n1141 );
    or g12186 ( n30634 , n26035 , n18450 );
    xnor g12187 ( n38328 , n11434 , n16509 );
    xnor g12188 ( n8187 , n11855 , n22714 );
    or g12189 ( n400 , n23489 , n25743 );
    or g12190 ( n21980 , n3583 , n23131 );
    and g12191 ( n9298 , n32443 , n4337 );
    nor g12192 ( n14812 , n6751 , n29934 );
    and g12193 ( n17031 , n32017 , n11158 );
    and g12194 ( n37641 , n11664 , n27078 );
    or g12195 ( n19023 , n37759 , n21372 );
    and g12196 ( n22721 , n7592 , n18163 );
    or g12197 ( n36086 , n28402 , n6119 );
    or g12198 ( n28151 , n40252 , n41923 );
    not g12199 ( n24991 , n5915 );
    and g12200 ( n17856 , n2676 , n17444 );
    and g12201 ( n4841 , n38316 , n29877 );
    or g12202 ( n18322 , n42633 , n21847 );
    xnor g12203 ( n36467 , n29376 , n28071 );
    or g12204 ( n10257 , n21831 , n15478 );
    xnor g12205 ( n38147 , n23561 , n39266 );
    and g12206 ( n29598 , n40260 , n2852 );
    or g12207 ( n26519 , n16121 , n4915 );
    and g12208 ( n4274 , n37132 , n14631 );
    or g12209 ( n33686 , n34631 , n28335 );
    or g12210 ( n11521 , n19372 , n3100 );
    and g12211 ( n7350 , n38699 , n18099 );
    xnor g12212 ( n10381 , n30764 , n21094 );
    not g12213 ( n31871 , n33425 );
    and g12214 ( n23856 , n3843 , n39143 );
    not g12215 ( n12835 , n32146 );
    or g12216 ( n32403 , n12212 , n34577 );
    or g12217 ( n27707 , n1653 , n39481 );
    or g12218 ( n26774 , n15579 , n9782 );
    xnor g12219 ( n34276 , n34783 , n7049 );
    and g12220 ( n3254 , n9898 , n24422 );
    or g12221 ( n7132 , n16366 , n42446 );
    and g12222 ( n10486 , n26517 , n8036 );
    nor g12223 ( n22593 , n37078 , n37126 );
    or g12224 ( n26143 , n15429 , n2272 );
    or g12225 ( n29745 , n24974 , n35174 );
    not g12226 ( n12777 , n25697 );
    xnor g12227 ( n11342 , n18736 , n10272 );
    nor g12228 ( n8870 , n14515 , n9338 );
    and g12229 ( n32295 , n23666 , n39291 );
    xnor g12230 ( n10799 , n13261 , n6734 );
    and g12231 ( n4156 , n19542 , n32664 );
    or g12232 ( n27997 , n40462 , n823 );
    or g12233 ( n34604 , n23519 , n17321 );
    nor g12234 ( n38345 , n465 , n32237 );
    or g12235 ( n10661 , n25648 , n33607 );
    and g12236 ( n8235 , n14246 , n28966 );
    xnor g12237 ( n30559 , n11436 , n26988 );
    not g12238 ( n21759 , n28576 );
    not g12239 ( n3437 , n33632 );
    or g12240 ( n21158 , n30235 , n16600 );
    xnor g12241 ( n14239 , n32470 , n14856 );
    or g12242 ( n18487 , n10900 , n1871 );
    nor g12243 ( n42457 , n16598 , n17021 );
    or g12244 ( n35244 , n31091 , n16115 );
    or g12245 ( n5598 , n33380 , n21240 );
    and g12246 ( n16281 , n19689 , n3159 );
    or g12247 ( n15164 , n36235 , n37096 );
    xnor g12248 ( n12090 , n8058 , n9605 );
    nor g12249 ( n17044 , n35892 , n39824 );
    not g12250 ( n30616 , n29777 );
    or g12251 ( n36732 , n41143 , n29385 );
    nor g12252 ( n26349 , n22086 , n38977 );
    or g12253 ( n17889 , n39733 , n34569 );
    or g12254 ( n3577 , n20407 , n21025 );
    and g12255 ( n5462 , n27565 , n35535 );
    and g12256 ( n24979 , n33618 , n13531 );
    nor g12257 ( n33877 , n22407 , n34396 );
    not g12258 ( n10460 , n30510 );
    xnor g12259 ( n25942 , n30264 , n2559 );
    nor g12260 ( n29790 , n2183 , n40036 );
    and g12261 ( n11901 , n23066 , n13541 );
    or g12262 ( n662 , n40567 , n33040 );
    nor g12263 ( n27471 , n21340 , n38033 );
    not g12264 ( n22631 , n25994 );
    nor g12265 ( n9129 , n35678 , n35010 );
    nor g12266 ( n11082 , n32701 , n21239 );
    xnor g12267 ( n36895 , n2501 , n35070 );
    or g12268 ( n21251 , n32430 , n19842 );
    not g12269 ( n28432 , n29674 );
    not g12270 ( n39573 , n23274 );
    nor g12271 ( n34094 , n24750 , n35636 );
    and g12272 ( n27352 , n2942 , n42047 );
    or g12273 ( n5107 , n18424 , n13130 );
    and g12274 ( n2646 , n17674 , n4978 );
    xnor g12275 ( n4002 , n22255 , n32404 );
    xnor g12276 ( n10123 , n21457 , n28086 );
    or g12277 ( n21074 , n18806 , n31361 );
    or g12278 ( n4009 , n17120 , n34885 );
    nor g12279 ( n40413 , n30161 , n42162 );
    nor g12280 ( n28035 , n28581 , n30246 );
    nor g12281 ( n28599 , n16598 , n159 );
    xnor g12282 ( n36314 , n37662 , n5889 );
    not g12283 ( n5823 , n20788 );
    not g12284 ( n33978 , n19614 );
    or g12285 ( n30689 , n42745 , n5760 );
    and g12286 ( n10669 , n9715 , n18422 );
    xnor g12287 ( n9027 , n29740 , n11637 );
    or g12288 ( n16107 , n37905 , n7260 );
    and g12289 ( n26424 , n27064 , n23458 );
    and g12290 ( n6711 , n7098 , n1483 );
    nor g12291 ( n34096 , n27728 , n2665 );
    nor g12292 ( n4682 , n35011 , n1590 );
    or g12293 ( n17966 , n27772 , n30378 );
    xnor g12294 ( n19403 , n10639 , n39922 );
    or g12295 ( n31276 , n3222 , n12003 );
    or g12296 ( n24502 , n15139 , n39730 );
    not g12297 ( n40954 , n3361 );
    and g12298 ( n16147 , n9310 , n13931 );
    nor g12299 ( n19411 , n12389 , n40422 );
    not g12300 ( n34446 , n2497 );
    not g12301 ( n35790 , n17567 );
    or g12302 ( n647 , n26964 , n30404 );
    nor g12303 ( n10736 , n3117 , n23298 );
    and g12304 ( n12846 , n38156 , n2869 );
    or g12305 ( n19165 , n18473 , n9802 );
    and g12306 ( n42701 , n38290 , n16353 );
    xnor g12307 ( n19268 , n37829 , n40287 );
    and g12308 ( n17359 , n35665 , n25412 );
    nor g12309 ( n19092 , n15068 , n28767 );
    or g12310 ( n26718 , n38879 , n323 );
    xnor g12311 ( n21677 , n30870 , n34125 );
    not g12312 ( n32446 , n13668 );
    or g12313 ( n6706 , n42429 , n15425 );
    or g12314 ( n22686 , n9601 , n24114 );
    or g12315 ( n17671 , n33624 , n6845 );
    nor g12316 ( n25419 , n3621 , n22163 );
    or g12317 ( n33571 , n7989 , n36027 );
    or g12318 ( n30366 , n27884 , n33232 );
    nor g12319 ( n19083 , n33595 , n30798 );
    or g12320 ( n32207 , n15565 , n24440 );
    and g12321 ( n35280 , n3099 , n10479 );
    and g12322 ( n32956 , n12775 , n21490 );
    or g12323 ( n33593 , n514 , n4621 );
    or g12324 ( n24678 , n26576 , n5385 );
    or g12325 ( n10566 , n19927 , n14053 );
    xnor g12326 ( n32204 , n33875 , n40518 );
    xnor g12327 ( n38648 , n34687 , n11603 );
    or g12328 ( n3614 , n12413 , n30428 );
    or g12329 ( n36188 , n15936 , n19259 );
    or g12330 ( n25946 , n38931 , n28447 );
    and g12331 ( n14607 , n7734 , n36907 );
    nor g12332 ( n10240 , n2445 , n23973 );
    or g12333 ( n18746 , n4391 , n1088 );
    xnor g12334 ( n27978 , n3193 , n10109 );
    not g12335 ( n28551 , n22312 );
    not g12336 ( n14202 , n8047 );
    or g12337 ( n8153 , n18618 , n27494 );
    not g12338 ( n24202 , n34887 );
    or g12339 ( n25837 , n13486 , n9258 );
    xnor g12340 ( n24915 , n19319 , n36469 );
    nor g12341 ( n33174 , n17193 , n15473 );
    or g12342 ( n40622 , n7989 , n14283 );
    and g12343 ( n519 , n27235 , n6981 );
    or g12344 ( n38535 , n7651 , n22889 );
    not g12345 ( n19744 , n41200 );
    or g12346 ( n5576 , n41546 , n25683 );
    or g12347 ( n5321 , n14800 , n6842 );
    and g12348 ( n13285 , n36994 , n29745 );
    or g12349 ( n24425 , n26116 , n8559 );
    and g12350 ( n31809 , n8639 , n21398 );
    or g12351 ( n18145 , n19899 , n8722 );
    not g12352 ( n16471 , n27822 );
    not g12353 ( n5245 , n32319 );
    or g12354 ( n9639 , n39954 , n24926 );
    or g12355 ( n28609 , n33294 , n42703 );
    nor g12356 ( n41665 , n19055 , n25314 );
    nor g12357 ( n5121 , n26964 , n13193 );
    or g12358 ( n35986 , n9544 , n36858 );
    or g12359 ( n6682 , n36399 , n4220 );
    nor g12360 ( n10935 , n7509 , n5537 );
    not g12361 ( n27767 , n38504 );
    xnor g12362 ( n23727 , n9951 , n22336 );
    and g12363 ( n38309 , n8612 , n11179 );
    and g12364 ( n41543 , n20981 , n24862 );
    or g12365 ( n33373 , n3653 , n6541 );
    and g12366 ( n31282 , n11606 , n9571 );
    or g12367 ( n36429 , n39927 , n41812 );
    or g12368 ( n3260 , n31263 , n14216 );
    or g12369 ( n36366 , n33737 , n12956 );
    or g12370 ( n8203 , n36253 , n36997 );
    or g12371 ( n82 , n36820 , n13912 );
    not g12372 ( n30235 , n15133 );
    nor g12373 ( n19336 , n19787 , n29330 );
    nor g12374 ( n2457 , n10929 , n5256 );
    and g12375 ( n27831 , n2540 , n2246 );
    not g12376 ( n34105 , n1615 );
    not g12377 ( n21249 , n1398 );
    and g12378 ( n27103 , n17690 , n35888 );
    or g12379 ( n20669 , n6657 , n32410 );
    and g12380 ( n6937 , n12585 , n38809 );
    or g12381 ( n14960 , n28647 , n32745 );
    and g12382 ( n37270 , n3487 , n5945 );
    not g12383 ( n13623 , n17373 );
    or g12384 ( n16621 , n4635 , n10946 );
    not g12385 ( n9480 , n27667 );
    nor g12386 ( n32032 , n14707 , n19802 );
    and g12387 ( n36790 , n38627 , n33360 );
    not g12388 ( n17406 , n16507 );
    nor g12389 ( n31905 , n34474 , n21400 );
    or g12390 ( n4710 , n18308 , n35566 );
    and g12391 ( n27273 , n30319 , n20555 );
    or g12392 ( n8348 , n20118 , n946 );
    or g12393 ( n23830 , n33484 , n41810 );
    xnor g12394 ( n34582 , n37309 , n24618 );
    nor g12395 ( n39448 , n14347 , n14372 );
    not g12396 ( n20412 , n41153 );
    or g12397 ( n20426 , n10172 , n14749 );
    nor g12398 ( n41429 , n24356 , n19888 );
    and g12399 ( n26113 , n37616 , n9037 );
    or g12400 ( n40377 , n38494 , n32483 );
    xnor g12401 ( n26659 , n4143 , n2500 );
    or g12402 ( n12292 , n38879 , n8994 );
    and g12403 ( n39003 , n24619 , n27418 );
    not g12404 ( n12806 , n38828 );
    or g12405 ( n8077 , n32662 , n40554 );
    or g12406 ( n40121 , n35243 , n25036 );
    or g12407 ( n31572 , n26617 , n23302 );
    xnor g12408 ( n29376 , n2799 , n1064 );
    or g12409 ( n19998 , n20567 , n2308 );
    or g12410 ( n875 , n15967 , n2850 );
    or g12411 ( n20844 , n32475 , n41287 );
    or g12412 ( n21790 , n21011 , n1061 );
    xnor g12413 ( n9751 , n136 , n37683 );
    and g12414 ( n552 , n24272 , n17403 );
    xnor g12415 ( n29865 , n15353 , n1495 );
    and g12416 ( n3569 , n12428 , n31752 );
    and g12417 ( n37030 , n41979 , n7184 );
    or g12418 ( n31922 , n9145 , n27640 );
    not g12419 ( n28252 , n11677 );
    not g12420 ( n32605 , n11900 );
    not g12421 ( n11049 , n26643 );
    nor g12422 ( n30265 , n7356 , n42288 );
    or g12423 ( n39574 , n16738 , n29407 );
    xnor g12424 ( n35506 , n18520 , n7635 );
    not g12425 ( n40299 , n18524 );
    and g12426 ( n20454 , n13252 , n3058 );
    or g12427 ( n37286 , n17860 , n4646 );
    not g12428 ( n32793 , n26941 );
    or g12429 ( n26818 , n34123 , n36084 );
    or g12430 ( n32928 , n29108 , n34308 );
    or g12431 ( n3505 , n5571 , n34491 );
    nor g12432 ( n35951 , n32128 , n24120 );
    or g12433 ( n21445 , n16715 , n38336 );
    and g12434 ( n31021 , n15427 , n21270 );
    or g12435 ( n8605 , n21983 , n31690 );
    not g12436 ( n10440 , n8290 );
    or g12437 ( n24444 , n3758 , n14556 );
    or g12438 ( n27342 , n23479 , n17139 );
    not g12439 ( n33843 , n18969 );
    xnor g12440 ( n10653 , n3837 , n28572 );
    and g12441 ( n30208 , n22627 , n22414 );
    nor g12442 ( n30499 , n22753 , n23450 );
    not g12443 ( n33051 , n1058 );
    or g12444 ( n2282 , n17077 , n20032 );
    and g12445 ( n7227 , n16065 , n11088 );
    xnor g12446 ( n36914 , n26345 , n23618 );
    and g12447 ( n16271 , n26507 , n3976 );
    not g12448 ( n37911 , n40008 );
    nor g12449 ( n29287 , n37639 , n4160 );
    nor g12450 ( n37713 , n15590 , n21393 );
    or g12451 ( n32659 , n11710 , n38411 );
    and g12452 ( n36205 , n16665 , n1271 );
    or g12453 ( n24280 , n8550 , n35483 );
    xnor g12454 ( n27906 , n4784 , n10028 );
    not g12455 ( n37397 , n30003 );
    or g12456 ( n17693 , n17108 , n7674 );
    nor g12457 ( n5011 , n40099 , n13196 );
    and g12458 ( n35689 , n15419 , n10033 );
    or g12459 ( n28397 , n6170 , n12555 );
    or g12460 ( n21680 , n2742 , n29155 );
    or g12461 ( n23195 , n24526 , n17373 );
    and g12462 ( n279 , n111 , n30526 );
    and g12463 ( n7307 , n4828 , n11221 );
    or g12464 ( n32636 , n9755 , n24828 );
    xnor g12465 ( n8008 , n41053 , n14259 );
    and g12466 ( n40566 , n35055 , n4932 );
    and g12467 ( n16920 , n26621 , n22488 );
    or g12468 ( n21739 , n33055 , n1539 );
    and g12469 ( n1933 , n4024 , n7104 );
    and g12470 ( n38845 , n30664 , n21093 );
    not g12471 ( n28632 , n3140 );
    or g12472 ( n7691 , n1273 , n21025 );
    or g12473 ( n25111 , n13007 , n29742 );
    not g12474 ( n31925 , n27182 );
    not g12475 ( n6319 , n19948 );
    xnor g12476 ( n38403 , n455 , n21060 );
    xnor g12477 ( n41901 , n31607 , n20683 );
    or g12478 ( n4198 , n19452 , n3409 );
    or g12479 ( n18193 , n30864 , n15484 );
    or g12480 ( n28682 , n3037 , n39675 );
    not g12481 ( n174 , n12634 );
    not g12482 ( n30413 , n15258 );
    xnor g12483 ( n29421 , n34690 , n9251 );
    and g12484 ( n24104 , n12593 , n2250 );
    not g12485 ( n21752 , n17205 );
    or g12486 ( n41495 , n40887 , n38438 );
    xnor g12487 ( n759 , n27574 , n20764 );
    or g12488 ( n14084 , n24286 , n26922 );
    and g12489 ( n39457 , n9404 , n3488 );
    or g12490 ( n8975 , n4447 , n18353 );
    or g12491 ( n1675 , n23572 , n12492 );
    or g12492 ( n12936 , n6346 , n14501 );
    or g12493 ( n706 , n27804 , n21015 );
    or g12494 ( n12667 , n16247 , n16633 );
    or g12495 ( n25028 , n35982 , n18234 );
    and g12496 ( n15832 , n36818 , n24532 );
    or g12497 ( n6269 , n17295 , n39144 );
    or g12498 ( n6927 , n39121 , n5629 );
    or g12499 ( n8845 , n23990 , n30064 );
    or g12500 ( n5515 , n35344 , n26063 );
    or g12501 ( n14173 , n15095 , n31616 );
    xnor g12502 ( n7894 , n37856 , n8494 );
    not g12503 ( n20085 , n18434 );
    or g12504 ( n18671 , n18236 , n33705 );
    not g12505 ( n16126 , n29310 );
    not g12506 ( n17874 , n28660 );
    nor g12507 ( n6712 , n17744 , n39972 );
    nor g12508 ( n36395 , n20026 , n42167 );
    xnor g12509 ( n40333 , n10590 , n24966 );
    nor g12510 ( n12245 , n28361 , n14188 );
    and g12511 ( n24539 , n32099 , n20973 );
    and g12512 ( n6371 , n539 , n42731 );
    not g12513 ( n6170 , n19832 );
    nor g12514 ( n20280 , n36070 , n6653 );
    not g12515 ( n25310 , n31162 );
    and g12516 ( n39922 , n35884 , n5499 );
    nor g12517 ( n16772 , n15178 , n20983 );
    xnor g12518 ( n36403 , n31291 , n10481 );
    or g12519 ( n10621 , n948 , n28950 );
    or g12520 ( n17458 , n28673 , n8322 );
    or g12521 ( n25931 , n16012 , n14287 );
    and g12522 ( n21770 , n58 , n17351 );
    and g12523 ( n27186 , n17316 , n42846 );
    nor g12524 ( n31939 , n21592 , n38622 );
    xnor g12525 ( n40833 , n6663 , n2369 );
    or g12526 ( n22907 , n5904 , n41549 );
    and g12527 ( n34228 , n666 , n8445 );
    or g12528 ( n27227 , n6953 , n16676 );
    nor g12529 ( n14820 , n13455 , n2633 );
    or g12530 ( n37189 , n15070 , n19359 );
    not g12531 ( n13759 , n28202 );
    or g12532 ( n25747 , n5798 , n14363 );
    xnor g12533 ( n40774 , n330 , n35933 );
    and g12534 ( n15986 , n312 , n29102 );
    not g12535 ( n34274 , n3085 );
    not g12536 ( n13332 , n41301 );
    not g12537 ( n11725 , n31172 );
    and g12538 ( n12531 , n18414 , n23169 );
    and g12539 ( n1767 , n1249 , n16185 );
    not g12540 ( n9488 , n29929 );
    nor g12541 ( n17254 , n11319 , n39922 );
    not g12542 ( n23895 , n14575 );
    or g12543 ( n30057 , n2440 , n34267 );
    or g12544 ( n34727 , n121 , n14770 );
    not g12545 ( n34052 , n34151 );
    or g12546 ( n1960 , n25672 , n40157 );
    or g12547 ( n3194 , n40790 , n38417 );
    nor g12548 ( n20299 , n41534 , n13473 );
    or g12549 ( n28940 , n13919 , n30570 );
    not g12550 ( n16404 , n13066 );
    not g12551 ( n9409 , n35844 );
    not g12552 ( n40770 , n9232 );
    and g12553 ( n333 , n9945 , n5214 );
    not g12554 ( n19844 , n34925 );
    or g12555 ( n4576 , n7657 , n27320 );
    or g12556 ( n12965 , n18105 , n23400 );
    or g12557 ( n17760 , n26693 , n33448 );
    or g12558 ( n39945 , n10505 , n17723 );
    not g12559 ( n36110 , n33362 );
    not g12560 ( n25961 , n39247 );
    xnor g12561 ( n26190 , n30549 , n41346 );
    or g12562 ( n22445 , n19969 , n10285 );
    xnor g12563 ( n2698 , n2127 , n3901 );
    xnor g12564 ( n29370 , n27710 , n14995 );
    nor g12565 ( n24820 , n3949 , n14609 );
    or g12566 ( n32665 , n20305 , n21822 );
    or g12567 ( n7941 , n42133 , n10374 );
    nor g12568 ( n18631 , n39406 , n30816 );
    not g12569 ( n34235 , n12984 );
    or g12570 ( n39172 , n1961 , n19750 );
    not g12571 ( n37702 , n18033 );
    and g12572 ( n38237 , n35235 , n16727 );
    and g12573 ( n18172 , n35119 , n30943 );
    or g12574 ( n522 , n1365 , n31748 );
    or g12575 ( n11910 , n30690 , n28239 );
    xnor g12576 ( n8457 , n2182 , n11487 );
    and g12577 ( n28157 , n6460 , n42172 );
    or g12578 ( n13910 , n2096 , n22525 );
    and g12579 ( n13642 , n37661 , n16878 );
    or g12580 ( n6475 , n12557 , n12832 );
    nor g12581 ( n20499 , n17120 , n8698 );
    not g12582 ( n31865 , n39426 );
    nor g12583 ( n34517 , n19020 , n39775 );
    and g12584 ( n5185 , n13203 , n3605 );
    or g12585 ( n25740 , n32961 , n4861 );
    or g12586 ( n23451 , n14272 , n3381 );
    xnor g12587 ( n35569 , n21929 , n38998 );
    nor g12588 ( n27642 , n4093 , n25400 );
    xnor g12589 ( n26522 , n42916 , n7054 );
    not g12590 ( n4180 , n9592 );
    or g12591 ( n14505 , n35338 , n23953 );
    or g12592 ( n21071 , n28021 , n1769 );
    nor g12593 ( n28789 , n27030 , n39678 );
    not g12594 ( n23342 , n5303 );
    xnor g12595 ( n30660 , n9304 , n20081 );
    xnor g12596 ( n3132 , n18850 , n830 );
    or g12597 ( n41850 , n21874 , n27034 );
    or g12598 ( n26304 , n10402 , n13282 );
    or g12599 ( n14257 , n12867 , n37332 );
    not g12600 ( n39021 , n29596 );
    or g12601 ( n4254 , n41403 , n11950 );
    or g12602 ( n4837 , n15044 , n2034 );
    not g12603 ( n4879 , n29474 );
    or g12604 ( n29747 , n19633 , n34772 );
    or g12605 ( n33979 , n35959 , n34019 );
    xnor g12606 ( n31719 , n18880 , n40478 );
    and g12607 ( n23657 , n11056 , n41334 );
    and g12608 ( n18578 , n5674 , n33872 );
    xnor g12609 ( n14356 , n5144 , n37954 );
    or g12610 ( n9385 , n33792 , n8699 );
    and g12611 ( n39949 , n15204 , n26395 );
    or g12612 ( n10567 , n20278 , n17654 );
    not g12613 ( n10454 , n41243 );
    not g12614 ( n9671 , n928 );
    or g12615 ( n4455 , n26488 , n35567 );
    or g12616 ( n15881 , n6006 , n38556 );
    nor g12617 ( n223 , n26345 , n33032 );
    or g12618 ( n40145 , n7096 , n17321 );
    and g12619 ( n1500 , n3395 , n6562 );
    xnor g12620 ( n11350 , n36009 , n3927 );
    xnor g12621 ( n11551 , n24388 , n13788 );
    nor g12622 ( n24196 , n9368 , n6266 );
    or g12623 ( n34395 , n18362 , n32605 );
    not g12624 ( n19667 , n42844 );
    or g12625 ( n34846 , n25047 , n11876 );
    and g12626 ( n657 , n19516 , n13227 );
    xnor g12627 ( n30433 , n19116 , n30757 );
    or g12628 ( n8342 , n3980 , n31871 );
    or g12629 ( n13704 , n23674 , n17576 );
    nor g12630 ( n27957 , n41728 , n39033 );
    not g12631 ( n39363 , n6653 );
    and g12632 ( n36891 , n275 , n7877 );
    or g12633 ( n9342 , n2701 , n41783 );
    or g12634 ( n7563 , n32350 , n42618 );
    or g12635 ( n33841 , n33569 , n21172 );
    and g12636 ( n10007 , n21346 , n40744 );
    and g12637 ( n4688 , n32301 , n32250 );
    or g12638 ( n42757 , n16910 , n19852 );
    not g12639 ( n4753 , n38194 );
    not g12640 ( n25552 , n2857 );
    nor g12641 ( n21928 , n17178 , n37717 );
    nor g12642 ( n25018 , n5964 , n30472 );
    or g12643 ( n29409 , n39337 , n893 );
    or g12644 ( n21391 , n2334 , n18393 );
    or g12645 ( n12827 , n36455 , n37654 );
    or g12646 ( n39062 , n23085 , n3616 );
    nor g12647 ( n27628 , n33981 , n1520 );
    and g12648 ( n27956 , n1713 , n3158 );
    or g12649 ( n40937 , n8657 , n2701 );
    xnor g12650 ( n22022 , n36998 , n21444 );
    nor g12651 ( n38962 , n18866 , n42180 );
    and g12652 ( n20328 , n27609 , n37483 );
    or g12653 ( n23769 , n40455 , n25659 );
    not g12654 ( n2182 , n29457 );
    or g12655 ( n22245 , n22493 , n13954 );
    nor g12656 ( n6173 , n29971 , n28909 );
    or g12657 ( n34900 , n3885 , n16216 );
    and g12658 ( n6094 , n42676 , n17459 );
    not g12659 ( n22355 , n39452 );
    xnor g12660 ( n34040 , n20920 , n38786 );
    or g12661 ( n19946 , n24496 , n36128 );
    or g12662 ( n35696 , n3767 , n12376 );
    and g12663 ( n4623 , n5146 , n6113 );
    xnor g12664 ( n25918 , n39532 , n2835 );
    not g12665 ( n7723 , n1681 );
    nor g12666 ( n36958 , n18866 , n19659 );
    or g12667 ( n29514 , n12152 , n42309 );
    and g12668 ( n28556 , n11668 , n11715 );
    or g12669 ( n38566 , n38193 , n41674 );
    nor g12670 ( n10497 , n25588 , n28329 );
    or g12671 ( n31658 , n15403 , n16199 );
    and g12672 ( n15473 , n36566 , n29876 );
    or g12673 ( n22804 , n6596 , n28837 );
    nor g12674 ( n5378 , n20991 , n13939 );
    not g12675 ( n7222 , n36015 );
    nor g12676 ( n1893 , n14707 , n40669 );
    not g12677 ( n10110 , n19029 );
    not g12678 ( n35238 , n39158 );
    xnor g12679 ( n35710 , n37085 , n14824 );
    and g12680 ( n36374 , n11070 , n30588 );
    or g12681 ( n37009 , n18689 , n262 );
    or g12682 ( n29413 , n18944 , n42152 );
    xnor g12683 ( n32225 , n37175 , n37566 );
    or g12684 ( n35855 , n40304 , n25303 );
    xnor g12685 ( n39864 , n28225 , n30717 );
    or g12686 ( n26144 , n18083 , n35218 );
    or g12687 ( n38003 , n18552 , n21869 );
    and g12688 ( n32770 , n15274 , n28265 );
    xnor g12689 ( n22941 , n105 , n25585 );
    not g12690 ( n26925 , n24504 );
    not g12691 ( n6943 , n34446 );
    xnor g12692 ( n3681 , n18756 , n14707 );
    and g12693 ( n20428 , n12800 , n26103 );
    not g12694 ( n3015 , n28775 );
    or g12695 ( n6357 , n3274 , n27457 );
    or g12696 ( n27935 , n28382 , n39528 );
    not g12697 ( n6548 , n26932 );
    and g12698 ( n9351 , n20489 , n17846 );
    xnor g12699 ( n39454 , n30318 , n8494 );
    and g12700 ( n32792 , n6477 , n24922 );
    not g12701 ( n33927 , n36696 );
    xnor g12702 ( n6052 , n8928 , n9338 );
    or g12703 ( n8719 , n4108 , n15925 );
    or g12704 ( n23327 , n40709 , n23626 );
    not g12705 ( n38573 , n5825 );
    or g12706 ( n19504 , n39196 , n27179 );
    not g12707 ( n18735 , n9321 );
    nor g12708 ( n39040 , n2223 , n42857 );
    not g12709 ( n6985 , n26637 );
    and g12710 ( n31522 , n41805 , n35089 );
    and g12711 ( n4124 , n18029 , n28728 );
    xnor g12712 ( n15257 , n37012 , n26543 );
    or g12713 ( n41171 , n2766 , n5978 );
    xnor g12714 ( n26082 , n5246 , n30600 );
    not g12715 ( n33617 , n9977 );
    or g12716 ( n9676 , n20837 , n25626 );
    or g12717 ( n13125 , n2639 , n38755 );
    or g12718 ( n21223 , n42152 , n23910 );
    xnor g12719 ( n12077 , n5099 , n20514 );
    or g12720 ( n10746 , n39061 , n8069 );
    or g12721 ( n9034 , n20453 , n37433 );
    and g12722 ( n5646 , n417 , n26748 );
    xnor g12723 ( n14942 , n2632 , n15440 );
    not g12724 ( n19364 , n13979 );
    not g12725 ( n4099 , n40655 );
    or g12726 ( n42800 , n31361 , n10785 );
    and g12727 ( n31216 , n11096 , n16778 );
    or g12728 ( n3054 , n17703 , n35878 );
    and g12729 ( n22133 , n8660 , n28172 );
    nor g12730 ( n22142 , n26187 , n39295 );
    not g12731 ( n29942 , n29094 );
    and g12732 ( n23302 , n4246 , n27402 );
    or g12733 ( n11256 , n16891 , n38673 );
    and g12734 ( n17069 , n21754 , n20170 );
    or g12735 ( n32121 , n13867 , n35829 );
    or g12736 ( n30335 , n34896 , n19762 );
    and g12737 ( n36468 , n17552 , n36847 );
    or g12738 ( n5028 , n13993 , n6916 );
    not g12739 ( n2608 , n570 );
    and g12740 ( n5974 , n11633 , n31431 );
    nor g12741 ( n756 , n1683 , n19349 );
    or g12742 ( n23970 , n7844 , n41347 );
    not g12743 ( n15858 , n30168 );
    xnor g12744 ( n8802 , n35322 , n41080 );
    or g12745 ( n33478 , n16564 , n35960 );
    and g12746 ( n28474 , n30649 , n29516 );
    or g12747 ( n31912 , n6558 , n23641 );
    or g12748 ( n29448 , n1042 , n4043 );
    or g12749 ( n38316 , n2199 , n35949 );
    nor g12750 ( n31696 , n6351 , n29668 );
    not g12751 ( n949 , n10631 );
    or g12752 ( n6325 , n18314 , n27983 );
    xnor g12753 ( n38936 , n784 , n8582 );
    or g12754 ( n34076 , n6046 , n32844 );
    or g12755 ( n35974 , n27172 , n19885 );
    or g12756 ( n2588 , n20293 , n31156 );
    or g12757 ( n28300 , n26265 , n5170 );
    nor g12758 ( n12459 , n12266 , n29701 );
    nor g12759 ( n10258 , n37237 , n20042 );
    or g12760 ( n37745 , n38256 , n32215 );
    or g12761 ( n12510 , n12721 , n30712 );
    not g12762 ( n14144 , n11087 );
    and g12763 ( n36861 , n17831 , n6096 );
    xnor g12764 ( n10865 , n24926 , n5964 );
    xnor g12765 ( n27158 , n5985 , n1561 );
    not g12766 ( n24599 , n28279 );
    and g12767 ( n18159 , n28692 , n7798 );
    or g12768 ( n36147 , n23880 , n35417 );
    and g12769 ( n16655 , n8931 , n42027 );
    and g12770 ( n7175 , n41325 , n35376 );
    or g12771 ( n32436 , n3627 , n11178 );
    or g12772 ( n12637 , n30647 , n12456 );
    or g12773 ( n5666 , n7379 , n8401 );
    and g12774 ( n31897 , n21058 , n37932 );
    and g12775 ( n37912 , n9017 , n3075 );
    xnor g12776 ( n12849 , n27808 , n27261 );
    not g12777 ( n17087 , n11677 );
    xnor g12778 ( n39887 , n31099 , n16529 );
    not g12779 ( n19189 , n30782 );
    or g12780 ( n29512 , n1136 , n23218 );
    xnor g12781 ( n8624 , n7268 , n25432 );
    or g12782 ( n19570 , n24173 , n11346 );
    and g12783 ( n398 , n11943 , n23663 );
    or g12784 ( n36565 , n24656 , n5624 );
    or g12785 ( n8709 , n9720 , n20653 );
    or g12786 ( n20736 , n26903 , n29709 );
    or g12787 ( n5267 , n9653 , n22610 );
    xnor g12788 ( n30489 , n11671 , n37049 );
    or g12789 ( n11401 , n17367 , n34939 );
    nor g12790 ( n34107 , n40053 , n38805 );
    and g12791 ( n26944 , n16063 , n18632 );
    xnor g12792 ( n9447 , n4651 , n3417 );
    not g12793 ( n19561 , n1384 );
    or g12794 ( n23987 , n13626 , n7679 );
    or g12795 ( n36382 , n17869 , n40931 );
    or g12796 ( n20672 , n30601 , n32518 );
    or g12797 ( n23376 , n1940 , n28139 );
    and g12798 ( n2258 , n26857 , n15497 );
    or g12799 ( n29822 , n28335 , n32819 );
    xnor g12800 ( n31375 , n1838 , n21977 );
    xnor g12801 ( n16221 , n36140 , n21376 );
    nor g12802 ( n12014 , n16069 , n40398 );
    or g12803 ( n7804 , n38704 , n36819 );
    or g12804 ( n2970 , n1072 , n42082 );
    xnor g12805 ( n36889 , n9688 , n11840 );
    and g12806 ( n10450 , n15711 , n35419 );
    not g12807 ( n20633 , n5254 );
    not g12808 ( n2387 , n37357 );
    or g12809 ( n16013 , n8387 , n30652 );
    and g12810 ( n24436 , n40658 , n12825 );
    xnor g12811 ( n35195 , n34875 , n22688 );
    and g12812 ( n12670 , n10444 , n42781 );
    not g12813 ( n14955 , n42652 );
    and g12814 ( n16712 , n34845 , n5917 );
    nor g12815 ( n19061 , n35301 , n35679 );
    or g12816 ( n29284 , n24015 , n5422 );
    not g12817 ( n25993 , n31583 );
    or g12818 ( n3104 , n10284 , n15009 );
    not g12819 ( n18192 , n10748 );
    or g12820 ( n18888 , n42896 , n22144 );
    or g12821 ( n15716 , n6606 , n10874 );
    not g12822 ( n30254 , n7505 );
    not g12823 ( n4702 , n11675 );
    and g12824 ( n8111 , n41369 , n24544 );
    xnor g12825 ( n4551 , n41395 , n34025 );
    not g12826 ( n19808 , n2368 );
    and g12827 ( n21204 , n27972 , n20577 );
    or g12828 ( n30849 , n37238 , n28239 );
    not g12829 ( n3023 , n13767 );
    and g12830 ( n29520 , n23185 , n19648 );
    and g12831 ( n315 , n1559 , n41948 );
    or g12832 ( n10348 , n15149 , n2026 );
    not g12833 ( n3937 , n19477 );
    or g12834 ( n27048 , n9248 , n9464 );
    or g12835 ( n11465 , n26122 , n32764 );
    or g12836 ( n18780 , n40443 , n8481 );
    and g12837 ( n35155 , n25373 , n41817 );
    nor g12838 ( n33205 , n28726 , n32990 );
    nor g12839 ( n29039 , n5964 , n39694 );
    and g12840 ( n14884 , n8018 , n41994 );
    not g12841 ( n12828 , n40300 );
    nor g12842 ( n2364 , n4275 , n34536 );
    or g12843 ( n13429 , n37646 , n14487 );
    and g12844 ( n42045 , n34837 , n30774 );
    or g12845 ( n4544 , n15500 , n22767 );
    and g12846 ( n19242 , n25196 , n12694 );
    and g12847 ( n21915 , n37624 , n12441 );
    or g12848 ( n2871 , n11925 , n2577 );
    or g12849 ( n19638 , n37806 , n30466 );
    not g12850 ( n29068 , n23835 );
    or g12851 ( n31230 , n37755 , n38279 );
    nor g12852 ( n42549 , n6549 , n23205 );
    not g12853 ( n5775 , n15944 );
    nor g12854 ( n16938 , n16817 , n37523 );
    or g12855 ( n38734 , n14626 , n11672 );
    or g12856 ( n12895 , n31924 , n36107 );
    or g12857 ( n15861 , n34584 , n23181 );
    or g12858 ( n35295 , n5833 , n31573 );
    not g12859 ( n902 , n16794 );
    and g12860 ( n37848 , n34892 , n8287 );
    or g12861 ( n176 , n4335 , n18779 );
    not g12862 ( n28161 , n10743 );
    xnor g12863 ( n18944 , n28631 , n20195 );
    or g12864 ( n22485 , n10332 , n16427 );
    or g12865 ( n10917 , n9072 , n14553 );
    and g12866 ( n15359 , n26770 , n23799 );
    or g12867 ( n23169 , n10928 , n40993 );
    not g12868 ( n15900 , n32019 );
    or g12869 ( n18152 , n12972 , n12867 );
    or g12870 ( n32674 , n32898 , n12754 );
    not g12871 ( n40642 , n5794 );
    and g12872 ( n29440 , n6313 , n21645 );
    or g12873 ( n18415 , n4946 , n34949 );
    or g12874 ( n41830 , n14945 , n14618 );
    nor g12875 ( n13819 , n26172 , n37182 );
    nor g12876 ( n11496 , n19957 , n16234 );
    or g12877 ( n464 , n32035 , n42765 );
    or g12878 ( n31867 , n7302 , n20112 );
    or g12879 ( n21171 , n34007 , n33655 );
    or g12880 ( n13928 , n40930 , n31321 );
    not g12881 ( n34433 , n41357 );
    or g12882 ( n8292 , n35526 , n37826 );
    and g12883 ( n33407 , n33368 , n9167 );
    and g12884 ( n9936 , n20779 , n17409 );
    or g12885 ( n32823 , n11980 , n12843 );
    or g12886 ( n22481 , n11038 , n37244 );
    or g12887 ( n42633 , n32449 , n36962 );
    or g12888 ( n31028 , n28109 , n40555 );
    and g12889 ( n5042 , n20059 , n36100 );
    not g12890 ( n28647 , n12318 );
    and g12891 ( n4522 , n2045 , n29975 );
    or g12892 ( n18448 , n21942 , n29619 );
    and g12893 ( n27234 , n14828 , n35186 );
    and g12894 ( n28316 , n32530 , n15819 );
    and g12895 ( n33179 , n14498 , n8315 );
    or g12896 ( n28332 , n2105 , n25951 );
    or g12897 ( n35183 , n28647 , n40665 );
    not g12898 ( n18285 , n22660 );
    or g12899 ( n16576 , n40350 , n35469 );
    nor g12900 ( n14671 , n41040 , n7087 );
    not g12901 ( n36922 , n20800 );
    not g12902 ( n29027 , n30611 );
    and g12903 ( n54 , n38399 , n32468 );
    nor g12904 ( n30444 , n14105 , n20760 );
    or g12905 ( n13103 , n22935 , n13747 );
    not g12906 ( n32892 , n29429 );
    or g12907 ( n128 , n41525 , n31094 );
    and g12908 ( n24864 , n33579 , n42329 );
    and g12909 ( n28721 , n19910 , n23276 );
    not g12910 ( n16316 , n5726 );
    or g12911 ( n40863 , n7623 , n35732 );
    and g12912 ( n28766 , n10076 , n24545 );
    and g12913 ( n34941 , n14798 , n15788 );
    and g12914 ( n42440 , n490 , n39899 );
    nor g12915 ( n16408 , n40777 , n28906 );
    or g12916 ( n25433 , n39277 , n16466 );
    nor g12917 ( n41996 , n9234 , n21218 );
    or g12918 ( n23483 , n21451 , n28428 );
    or g12919 ( n18253 , n3712 , n27109 );
    or g12920 ( n38210 , n36641 , n31403 );
    not g12921 ( n101 , n2093 );
    and g12922 ( n20850 , n4072 , n25533 );
    and g12923 ( n23077 , n9948 , n28759 );
    not g12924 ( n35780 , n28675 );
    or g12925 ( n13644 , n38494 , n22757 );
    not g12926 ( n6648 , n9895 );
    or g12927 ( n32989 , n32683 , n9530 );
    xnor g12928 ( n29692 , n12630 , n37290 );
    nor g12929 ( n8369 , n35723 , n3391 );
    or g12930 ( n37982 , n35633 , n27316 );
    or g12931 ( n11194 , n2517 , n37294 );
    xnor g12932 ( n17325 , n29441 , n35325 );
    nor g12933 ( n6806 , n35310 , n17218 );
    nor g12934 ( n24344 , n34686 , n15271 );
    not g12935 ( n7870 , n3539 );
    or g12936 ( n5758 , n29183 , n32467 );
    not g12937 ( n41211 , n36557 );
    or g12938 ( n32652 , n28335 , n35777 );
    and g12939 ( n994 , n13230 , n21305 );
    nor g12940 ( n10692 , n34920 , n39100 );
    xnor g12941 ( n37224 , n25574 , n1156 );
    or g12942 ( n616 , n11327 , n13563 );
    and g12943 ( n36240 , n7047 , n32333 );
    not g12944 ( n9859 , n11015 );
    or g12945 ( n21834 , n37707 , n35070 );
    and g12946 ( n29167 , n34261 , n25328 );
    or g12947 ( n19621 , n32348 , n28461 );
    or g12948 ( n5909 , n25588 , n14847 );
    and g12949 ( n24484 , n7735 , n13856 );
    or g12950 ( n12034 , n2492 , n34199 );
    and g12951 ( n15889 , n3836 , n2625 );
    not g12952 ( n25626 , n3280 );
    not g12953 ( n40674 , n20076 );
    xnor g12954 ( n37297 , n36009 , n8143 );
    not g12955 ( n4779 , n12772 );
    or g12956 ( n24315 , n29803 , n13655 );
    or g12957 ( n17271 , n22333 , n12925 );
    or g12958 ( n2166 , n26057 , n19643 );
    and g12959 ( n584 , n27707 , n34649 );
    and g12960 ( n17721 , n9618 , n39396 );
    or g12961 ( n5228 , n14503 , n21620 );
    or g12962 ( n22894 , n13476 , n21287 );
    not g12963 ( n2631 , n26056 );
    not g12964 ( n19635 , n4021 );
    or g12965 ( n29590 , n38269 , n16730 );
    and g12966 ( n18517 , n27726 , n22459 );
    or g12967 ( n34701 , n30414 , n36443 );
    not g12968 ( n33187 , n13179 );
    or g12969 ( n3903 , n27840 , n6975 );
    not g12970 ( n5891 , n21975 );
    nor g12971 ( n5126 , n37671 , n30355 );
    or g12972 ( n36135 , n25424 , n1750 );
    and g12973 ( n10299 , n6650 , n33857 );
    or g12974 ( n14033 , n40679 , n8624 );
    not g12975 ( n1762 , n29475 );
    xnor g12976 ( n19320 , n22842 , n21747 );
    xnor g12977 ( n3285 , n18689 , n22589 );
    xnor g12978 ( n14301 , n14969 , n2404 );
    or g12979 ( n33159 , n4729 , n5904 );
    nor g12980 ( n2144 , n34837 , n30774 );
    and g12981 ( n28515 , n8887 , n25189 );
    xnor g12982 ( n40593 , n42822 , n24533 );
    or g12983 ( n4453 , n19727 , n6427 );
    or g12984 ( n42339 , n17828 , n30402 );
    and g12985 ( n14228 , n19859 , n11621 );
    or g12986 ( n38649 , n23489 , n6494 );
    or g12987 ( n3463 , n11275 , n7534 );
    nor g12988 ( n32775 , n35173 , n40061 );
    nor g12989 ( n26379 , n28939 , n6321 );
    not g12990 ( n19933 , n38974 );
    or g12991 ( n41677 , n26088 , n29996 );
    and g12992 ( n28846 , n33058 , n9095 );
    and g12993 ( n31127 , n16723 , n5783 );
    or g12994 ( n21593 , n20850 , n24175 );
    xnor g12995 ( n35968 , n4972 , n28684 );
    or g12996 ( n2072 , n6240 , n7415 );
    or g12997 ( n86 , n12235 , n33260 );
    xnor g12998 ( n11752 , n4343 , n13034 );
    or g12999 ( n26480 , n18798 , n5025 );
    or g13000 ( n34699 , n18130 , n41058 );
    and g13001 ( n17078 , n1714 , n29274 );
    not g13002 ( n1995 , n29429 );
    or g13003 ( n42261 , n27681 , n33345 );
    and g13004 ( n28130 , n2195 , n42673 );
    and g13005 ( n13061 , n32690 , n2826 );
    not g13006 ( n42060 , n6442 );
    not g13007 ( n30354 , n42406 );
    not g13008 ( n22989 , n27614 );
    or g13009 ( n24721 , n22967 , n9901 );
    and g13010 ( n23989 , n464 , n15360 );
    or g13011 ( n30003 , n32201 , n26994 );
    or g13012 ( n1779 , n27417 , n37315 );
    or g13013 ( n31502 , n36005 , n9635 );
    and g13014 ( n22462 , n32928 , n28992 );
    or g13015 ( n27689 , n8164 , n35655 );
    and g13016 ( n29361 , n9902 , n9071 );
    not g13017 ( n9001 , n14004 );
    and g13018 ( n36587 , n32915 , n16242 );
    xnor g13019 ( n6989 , n1965 , n14803 );
    and g13020 ( n2503 , n687 , n20744 );
    and g13021 ( n34011 , n32872 , n31397 );
    nor g13022 ( n41074 , n16728 , n22955 );
    or g13023 ( n5563 , n42723 , n36988 );
    nor g13024 ( n7750 , n38350 , n29254 );
    xnor g13025 ( n8851 , n28541 , n10410 );
    or g13026 ( n36906 , n27603 , n6907 );
    nor g13027 ( n40827 , n7476 , n22585 );
    nor g13028 ( n14381 , n105 , n36124 );
    and g13029 ( n17623 , n7782 , n36008 );
    xnor g13030 ( n28445 , n31202 , n39349 );
    xnor g13031 ( n19307 , n21184 , n30243 );
    or g13032 ( n28352 , n38594 , n36848 );
    or g13033 ( n3763 , n14705 , n27632 );
    not g13034 ( n15573 , n17406 );
    or g13035 ( n37740 , n20824 , n24068 );
    or g13036 ( n40330 , n20691 , n28479 );
    xnor g13037 ( n8063 , n31989 , n15799 );
    nor g13038 ( n6169 , n34857 , n34078 );
    not g13039 ( n20172 , n5372 );
    or g13040 ( n22180 , n18523 , n4099 );
    not g13041 ( n2585 , n9447 );
    or g13042 ( n32736 , n24305 , n22885 );
    or g13043 ( n39748 , n14281 , n40559 );
    xnor g13044 ( n11535 , n29740 , n33869 );
    and g13045 ( n29345 , n15739 , n19384 );
    not g13046 ( n9412 , n26268 );
    or g13047 ( n8643 , n20070 , n30081 );
    or g13048 ( n31467 , n11317 , n32654 );
    or g13049 ( n31179 , n42327 , n30143 );
    xnor g13050 ( n11636 , n28083 , n38986 );
    or g13051 ( n110 , n28696 , n3974 );
    or g13052 ( n23247 , n25934 , n38887 );
    and g13053 ( n3556 , n18457 , n24481 );
    and g13054 ( n36266 , n898 , n41840 );
    xnor g13055 ( n25473 , n23823 , n2379 );
    or g13056 ( n12093 , n42722 , n29012 );
    or g13057 ( n15471 , n22883 , n24083 );
    or g13058 ( n28439 , n12348 , n702 );
    or g13059 ( n14419 , n8770 , n10664 );
    not g13060 ( n10760 , n24466 );
    or g13061 ( n34071 , n37171 , n15951 );
    or g13062 ( n5319 , n29621 , n32243 );
    or g13063 ( n28543 , n38710 , n2234 );
    nor g13064 ( n8863 , n25588 , n39505 );
    not g13065 ( n9003 , n9533 );
    or g13066 ( n36675 , n7776 , n2149 );
    or g13067 ( n24019 , n21048 , n31129 );
    or g13068 ( n4389 , n40223 , n27178 );
    or g13069 ( n32492 , n35921 , n34285 );
    not g13070 ( n766 , n21263 );
    or g13071 ( n30135 , n33419 , n8246 );
    or g13072 ( n12973 , n1776 , n40612 );
    or g13073 ( n42219 , n2407 , n31399 );
    or g13074 ( n42430 , n30483 , n11077 );
    not g13075 ( n22842 , n10943 );
    or g13076 ( n39244 , n40139 , n29058 );
    or g13077 ( n36709 , n34797 , n35330 );
    and g13078 ( n13059 , n38252 , n21511 );
    or g13079 ( n4588 , n26667 , n11178 );
    not g13080 ( n18247 , n1986 );
    xnor g13081 ( n34835 , n11534 , n22900 );
    xnor g13082 ( n6164 , n28225 , n17401 );
    and g13083 ( n7689 , n39854 , n14906 );
    or g13084 ( n13521 , n38249 , n6933 );
    or g13085 ( n29107 , n10515 , n28028 );
    not g13086 ( n34329 , n28347 );
    nor g13087 ( n39915 , n22825 , n28993 );
    nor g13088 ( n8467 , n35255 , n20497 );
    nor g13089 ( n20293 , n13052 , n33589 );
    xnor g13090 ( n6617 , n4334 , n34415 );
    and g13091 ( n7814 , n18531 , n22341 );
    not g13092 ( n1719 , n35423 );
    not g13093 ( n24493 , n39457 );
    nor g13094 ( n16309 , n5367 , n25464 );
    or g13095 ( n21273 , n24001 , n30652 );
    or g13096 ( n5474 , n17927 , n6494 );
    or g13097 ( n36055 , n34433 , n21390 );
    xnor g13098 ( n8125 , n20582 , n19012 );
    or g13099 ( n10358 , n38313 , n22272 );
    or g13100 ( n14255 , n1640 , n17827 );
    xnor g13101 ( n3380 , n1305 , n40535 );
    or g13102 ( n37424 , n30302 , n617 );
    and g13103 ( n39520 , n40653 , n28161 );
    or g13104 ( n6163 , n22911 , n25440 );
    not g13105 ( n41993 , n32982 );
    or g13106 ( n38900 , n4856 , n12198 );
    and g13107 ( n25656 , n37696 , n6356 );
    or g13108 ( n34847 , n36047 , n39929 );
    or g13109 ( n1706 , n12346 , n15685 );
    not g13110 ( n29973 , n34933 );
    or g13111 ( n42858 , n41910 , n40459 );
    xnor g13112 ( n13071 , n19459 , n26081 );
    or g13113 ( n33359 , n4063 , n41092 );
    or g13114 ( n26266 , n37817 , n29930 );
    or g13115 ( n38069 , n34337 , n8289 );
    or g13116 ( n3347 , n18366 , n26740 );
    nor g13117 ( n32799 , n22760 , n19213 );
    xnor g13118 ( n24106 , n2903 , n13824 );
    nor g13119 ( n31144 , n34292 , n34828 );
    and g13120 ( n35461 , n41913 , n31713 );
    nor g13121 ( n4100 , n30880 , n38332 );
    not g13122 ( n5929 , n601 );
    and g13123 ( n39862 , n6706 , n4211 );
    or g13124 ( n1898 , n2050 , n18841 );
    or g13125 ( n36004 , n12063 , n41410 );
    or g13126 ( n29066 , n37652 , n30477 );
    not g13127 ( n7567 , n28003 );
    and g13128 ( n21258 , n22848 , n41473 );
    xnor g13129 ( n8386 , n536 , n38236 );
    nor g13130 ( n5068 , n39266 , n9 );
    or g13131 ( n21057 , n5431 , n32521 );
    and g13132 ( n24857 , n29768 , n15684 );
    or g13133 ( n10342 , n42449 , n25886 );
    not g13134 ( n30226 , n6668 );
    or g13135 ( n14005 , n4121 , n41570 );
    or g13136 ( n24222 , n1006 , n1332 );
    or g13137 ( n19824 , n38039 , n39481 );
    nor g13138 ( n14804 , n7700 , n2673 );
    nor g13139 ( n38219 , n14707 , n12923 );
    not g13140 ( n1612 , n15268 );
    xnor g13141 ( n2102 , n10466 , n13570 );
    or g13142 ( n16493 , n6050 , n40605 );
    or g13143 ( n17463 , n37011 , n8729 );
    not g13144 ( n40092 , n2916 );
    not g13145 ( n39385 , n3007 );
    nor g13146 ( n24043 , n30377 , n15566 );
    and g13147 ( n26500 , n37052 , n35937 );
    and g13148 ( n11709 , n32225 , n1802 );
    or g13149 ( n26695 , n958 , n26927 );
    xnor g13150 ( n535 , n11436 , n11651 );
    and g13151 ( n14462 , n26859 , n8709 );
    xnor g13152 ( n3683 , n34731 , n25778 );
    nor g13153 ( n14286 , n39669 , n38807 );
    or g13154 ( n15546 , n33134 , n3116 );
    or g13155 ( n23612 , n7093 , n18337 );
    or g13156 ( n6731 , n34248 , n5813 );
    xnor g13157 ( n42742 , n12161 , n24841 );
    or g13158 ( n39601 , n2095 , n23781 );
    or g13159 ( n11332 , n6733 , n23703 );
    or g13160 ( n5139 , n10065 , n42152 );
    or g13161 ( n6958 , n28322 , n313 );
    not g13162 ( n13840 , n36115 );
    xnor g13163 ( n305 , n42060 , n36787 );
    xnor g13164 ( n32254 , n23080 , n11711 );
    and g13165 ( n24447 , n5474 , n38308 );
    or g13166 ( n22441 , n11640 , n22567 );
    or g13167 ( n35212 , n33408 , n9351 );
    not g13168 ( n25600 , n12742 );
    or g13169 ( n24903 , n2517 , n41262 );
    xor g13170 ( n14040 , n10813 , n18953 );
    not g13171 ( n9793 , n369 );
    not g13172 ( n9556 , n20267 );
    or g13173 ( n9403 , n896 , n6310 );
    not g13174 ( n24715 , n1667 );
    or g13175 ( n40383 , n13362 , n27385 );
    or g13176 ( n29070 , n13991 , n3636 );
    xnor g13177 ( n18802 , n34875 , n14877 );
    nor g13178 ( n6615 , n38879 , n6092 );
    and g13179 ( n18567 , n11094 , n32202 );
    or g13180 ( n40054 , n29388 , n41710 );
    or g13181 ( n15170 , n39059 , n25107 );
    and g13182 ( n41145 , n6661 , n35209 );
    or g13183 ( n4095 , n17336 , n36848 );
    or g13184 ( n40124 , n32068 , n22599 );
    and g13185 ( n6673 , n32050 , n42552 );
    nor g13186 ( n2703 , n14840 , n34804 );
    nor g13187 ( n30464 , n2631 , n19378 );
    and g13188 ( n39316 , n19937 , n6155 );
    or g13189 ( n23200 , n972 , n680 );
    and g13190 ( n23673 , n2889 , n33905 );
    or g13191 ( n17765 , n34626 , n35036 );
    xnor g13192 ( n340 , n1713 , n3158 );
    or g13193 ( n24296 , n39489 , n22909 );
    nor g13194 ( n5495 , n21930 , n40793 );
    or g13195 ( n26813 , n22440 , n14462 );
    or g13196 ( n42336 , n40462 , n13824 );
    or g13197 ( n18821 , n24693 , n1326 );
    or g13198 ( n13946 , n8453 , n28918 );
    nor g13199 ( n29046 , n34483 , n30423 );
    and g13200 ( n35843 , n30029 , n31885 );
    not g13201 ( n1681 , n8573 );
    and g13202 ( n4336 , n37021 , n28242 );
    and g13203 ( n1251 , n26547 , n8331 );
    or g13204 ( n12746 , n33245 , n14157 );
    not g13205 ( n7218 , n7032 );
    nor g13206 ( n3010 , n5310 , n18816 );
    or g13207 ( n22215 , n14076 , n25148 );
    or g13208 ( n38985 , n9110 , n39791 );
    and g13209 ( n17983 , n21729 , n12338 );
    or g13210 ( n2798 , n21319 , n22619 );
    not g13211 ( n32752 , n14233 );
    or g13212 ( n10470 , n13625 , n11178 );
    not g13213 ( n39804 , n17598 );
    not g13214 ( n30897 , n38618 );
    and g13215 ( n40775 , n11130 , n15103 );
    and g13216 ( n20112 , n23554 , n27285 );
    or g13217 ( n22511 , n31447 , n10018 );
    not g13218 ( n12159 , n29701 );
    or g13219 ( n26856 , n30598 , n14470 );
    or g13220 ( n8492 , n27081 , n3406 );
    xnor g13221 ( n34766 , n30218 , n23727 );
    or g13222 ( n6010 , n7643 , n1095 );
    or g13223 ( n32086 , n4490 , n23827 );
    or g13224 ( n3047 , n28892 , n41413 );
    and g13225 ( n3632 , n6238 , n39175 );
    not g13226 ( n17109 , n32637 );
    xnor g13227 ( n39351 , n8968 , n34036 );
    or g13228 ( n15614 , n10505 , n36141 );
    nor g13229 ( n5134 , n30956 , n21837 );
    xnor g13230 ( n26239 , n41695 , n9162 );
    or g13231 ( n35686 , n10488 , n25303 );
    xnor g13232 ( n28702 , n2501 , n15208 );
    and g13233 ( n41090 , n21982 , n25293 );
    and g13234 ( n42904 , n26118 , n26137 );
    or g13235 ( n21063 , n22371 , n235 );
    nor g13236 ( n19756 , n5634 , n41604 );
    not g13237 ( n4492 , n426 );
    not g13238 ( n9838 , n20312 );
    or g13239 ( n16612 , n24621 , n32136 );
    and g13240 ( n30717 , n5698 , n3273 );
    or g13241 ( n30324 , n16564 , n9212 );
    xnor g13242 ( n40042 , n9178 , n29472 );
    and g13243 ( n5101 , n19584 , n26563 );
    not g13244 ( n7266 , n2111 );
    not g13245 ( n8462 , n34710 );
    xnor g13246 ( n27534 , n27660 , n27558 );
    or g13247 ( n29206 , n19269 , n29319 );
    or g13248 ( n38722 , n22440 , n16768 );
    or g13249 ( n9099 , n18916 , n16129 );
    xnor g13250 ( n21816 , n35154 , n19509 );
    and g13251 ( n5839 , n2314 , n31887 );
    and g13252 ( n4468 , n13641 , n32021 );
    and g13253 ( n39420 , n39324 , n20061 );
    or g13254 ( n37937 , n5124 , n16354 );
    and g13255 ( n25398 , n5159 , n36191 );
    or g13256 ( n31063 , n4881 , n13076 );
    nor g13257 ( n33457 , n42000 , n32187 );
    and g13258 ( n36500 , n25639 , n18329 );
    xnor g13259 ( n16607 , n32984 , n10613 );
    or g13260 ( n33899 , n36077 , n26758 );
    nor g13261 ( n18612 , n38957 , n7537 );
    and g13262 ( n33450 , n42286 , n17150 );
    or g13263 ( n22609 , n32892 , n41602 );
    not g13264 ( n37725 , n37396 );
    and g13265 ( n22900 , n9527 , n1992 );
    and g13266 ( n22776 , n4429 , n1529 );
    xnor g13267 ( n16069 , n27334 , n29522 );
    or g13268 ( n25998 , n16967 , n12733 );
    or g13269 ( n5743 , n37513 , n9332 );
    not g13270 ( n41722 , n17749 );
    or g13271 ( n27004 , n3291 , n32256 );
    xnor g13272 ( n38398 , n9783 , n20003 );
    and g13273 ( n1064 , n3401 , n1695 );
    and g13274 ( n8805 , n1885 , n21405 );
    not g13275 ( n42274 , n31188 );
    or g13276 ( n30179 , n7970 , n2015 );
    or g13277 ( n21146 , n41534 , n9825 );
    nor g13278 ( n37117 , n36895 , n10952 );
    or g13279 ( n1259 , n2477 , n17060 );
    nor g13280 ( n37202 , n25891 , n707 );
    or g13281 ( n7411 , n28667 , n8761 );
    not g13282 ( n16627 , n17463 );
    or g13283 ( n20052 , n22761 , n38191 );
    not g13284 ( n18375 , n41883 );
    and g13285 ( n20260 , n30062 , n31822 );
    not g13286 ( n7802 , n5305 );
    xnor g13287 ( n4934 , n42042 , n11775 );
    not g13288 ( n30197 , n5676 );
    not g13289 ( n29702 , n42575 );
    xnor g13290 ( n9190 , n37922 , n8613 );
    xnor g13291 ( n25828 , n42064 , n39949 );
    xnor g13292 ( n34813 , n28443 , n37759 );
    and g13293 ( n34723 , n36963 , n25676 );
    or g13294 ( n5604 , n6759 , n13388 );
    xnor g13295 ( n31895 , n10256 , n3709 );
    and g13296 ( n27506 , n3428 , n3831 );
    nor g13297 ( n39928 , n17676 , n11308 );
    or g13298 ( n39664 , n15006 , n2082 );
    or g13299 ( n9011 , n23574 , n37331 );
    and g13300 ( n17638 , n11101 , n20661 );
    or g13301 ( n18049 , n41534 , n14700 );
    not g13302 ( n15439 , n4432 );
    nor g13303 ( n8032 , n38234 , n5907 );
    or g13304 ( n7588 , n19780 , n36266 );
    not g13305 ( n29312 , n32014 );
    or g13306 ( n25531 , n37429 , n14025 );
    not g13307 ( n7385 , n3336 );
    or g13308 ( n8376 , n6765 , n23895 );
    and g13309 ( n41103 , n30918 , n6407 );
    or g13310 ( n22725 , n8476 , n1050 );
    nor g13311 ( n30567 , n33981 , n5663 );
    nor g13312 ( n30399 , n10598 , n20033 );
    and g13313 ( n7790 , n22758 , n1117 );
    nor g13314 ( n11696 , n26425 , n11089 );
    xnor g13315 ( n23898 , n22842 , n12845 );
    nor g13316 ( n33541 , n24991 , n22502 );
    and g13317 ( n42243 , n26778 , n40020 );
    not g13318 ( n35234 , n25684 );
    and g13319 ( n19639 , n6465 , n17579 );
    or g13320 ( n11874 , n12762 , n7699 );
    nor g13321 ( n35864 , n32539 , n7040 );
    xnor g13322 ( n41419 , n41013 , n35809 );
    nor g13323 ( n42008 , n16827 , n41121 );
    and g13324 ( n32405 , n8974 , n4649 );
    and g13325 ( n3720 , n29362 , n32013 );
    and g13326 ( n41032 , n14564 , n29741 );
    or g13327 ( n10409 , n19113 , n3625 );
    nor g13328 ( n31531 , n38629 , n35539 );
    nor g13329 ( n579 , n7356 , n28425 );
    and g13330 ( n5298 , n33713 , n41984 );
    or g13331 ( n30925 , n37263 , n41909 );
    nor g13332 ( n23479 , n22387 , n20545 );
    or g13333 ( n24321 , n20156 , n33447 );
    nor g13334 ( n20790 , n22425 , n34702 );
    or g13335 ( n19564 , n10845 , n42733 );
    xnor g13336 ( n21114 , n3549 , n22266 );
    not g13337 ( n7257 , n38286 );
    nor g13338 ( n27163 , n27557 , n42315 );
    or g13339 ( n39653 , n34485 , n21164 );
    or g13340 ( n11624 , n20474 , n7220 );
    or g13341 ( n28665 , n6243 , n19720 );
    or g13342 ( n16458 , n24760 , n35426 );
    or g13343 ( n39648 , n7001 , n9646 );
    xnor g13344 ( n15512 , n30864 , n39282 );
    or g13345 ( n822 , n9524 , n42513 );
    or g13346 ( n15252 , n34787 , n40885 );
    or g13347 ( n11556 , n21372 , n16615 );
    xnor g13348 ( n37747 , n12146 , n19115 );
    or g13349 ( n23577 , n15934 , n21501 );
    and g13350 ( n19310 , n221 , n10723 );
    not g13351 ( n38423 , n14233 );
    and g13352 ( n23724 , n29611 , n1918 );
    nor g13353 ( n356 , n21256 , n15783 );
    or g13354 ( n20472 , n34565 , n20451 );
    and g13355 ( n15404 , n9465 , n40715 );
    and g13356 ( n7207 , n36336 , n7024 );
    or g13357 ( n13203 , n28760 , n9328 );
    not g13358 ( n38430 , n36119 );
    or g13359 ( n4010 , n14018 , n26767 );
    and g13360 ( n8924 , n2757 , n10287 );
    xnor g13361 ( n38974 , n10527 , n38143 );
    not g13362 ( n1850 , n38790 );
    nor g13363 ( n30238 , n17011 , n28188 );
    or g13364 ( n18856 , n29228 , n23895 );
    or g13365 ( n24911 , n1159 , n5539 );
    not g13366 ( n7702 , n1287 );
    not g13367 ( n40912 , n36762 );
    not g13368 ( n38104 , n11726 );
    or g13369 ( n36601 , n35407 , n8164 );
    and g13370 ( n14860 , n19814 , n3418 );
    not g13371 ( n16373 , n31577 );
    not g13372 ( n40022 , n18575 );
    or g13373 ( n25160 , n1961 , n14699 );
    nor g13374 ( n13655 , n41837 , n27474 );
    nor g13375 ( n34480 , n28812 , n2995 );
    xnor g13376 ( n37744 , n18466 , n39184 );
    nor g13377 ( n28261 , n42008 , n35141 );
    nor g13378 ( n14551 , n27289 , n39763 );
    or g13379 ( n3631 , n39445 , n33558 );
    or g13380 ( n20456 , n15070 , n32293 );
    and g13381 ( n21212 , n18604 , n37799 );
    or g13382 ( n31689 , n40515 , n9961 );
    not g13383 ( n19266 , n36847 );
    nor g13384 ( n31657 , n3491 , n1431 );
    xnor g13385 ( n39415 , n105 , n2244 );
    xnor g13386 ( n19172 , n11436 , n40722 );
    and g13387 ( n36810 , n3763 , n40414 );
    nor g13388 ( n38352 , n5896 , n225 );
    not g13389 ( n13098 , n2261 );
    or g13390 ( n5568 , n5310 , n5286 );
    or g13391 ( n18936 , n15006 , n27114 );
    nor g13392 ( n27648 , n3437 , n30687 );
    xnor g13393 ( n20905 , n5144 , n12582 );
    or g13394 ( n28052 , n17500 , n31634 );
    and g13395 ( n11199 , n42644 , n13167 );
    not g13396 ( n4921 , n28486 );
    or g13397 ( n30604 , n435 , n20401 );
    not g13398 ( n36181 , n33676 );
    or g13399 ( n20166 , n33504 , n7863 );
    and g13400 ( n196 , n3326 , n40923 );
    or g13401 ( n17305 , n34697 , n13356 );
    and g13402 ( n6889 , n23516 , n28930 );
    nor g13403 ( n28264 , n1617 , n39131 );
    and g13404 ( n4312 , n2374 , n39285 );
    or g13405 ( n16282 , n25262 , n21054 );
    not g13406 ( n35814 , n7574 );
    xnor g13407 ( n25445 , n39743 , n30486 );
    or g13408 ( n34487 , n22292 , n8805 );
    and g13409 ( n11816 , n40465 , n37679 );
    or g13410 ( n34124 , n10533 , n4625 );
    nor g13411 ( n6835 , n34565 , n17153 );
    or g13412 ( n5514 , n13435 , n25652 );
    xnor g13413 ( n27684 , n34352 , n24815 );
    xnor g13414 ( n27483 , n784 , n9887 );
    and g13415 ( n17845 , n4556 , n18262 );
    or g13416 ( n26486 , n30082 , n2976 );
    and g13417 ( n434 , n20487 , n20657 );
    and g13418 ( n38358 , n14989 , n31438 );
    or g13419 ( n24090 , n22061 , n7727 );
    or g13420 ( n31180 , n34588 , n35985 );
    not g13421 ( n40499 , n22660 );
    and g13422 ( n1449 , n33678 , n13953 );
    or g13423 ( n35681 , n11614 , n25300 );
    and g13424 ( n12251 , n8403 , n42332 );
    not g13425 ( n33537 , n5661 );
    nor g13426 ( n26456 , n34565 , n3477 );
    or g13427 ( n32574 , n22976 , n2675 );
    not g13428 ( n5910 , n9182 );
    and g13429 ( n8898 , n10135 , n18077 );
    and g13430 ( n23621 , n5737 , n8678 );
    or g13431 ( n39361 , n16666 , n4435 );
    and g13432 ( n27661 , n29341 , n4395 );
    not g13433 ( n3804 , n32020 );
    nor g13434 ( n19358 , n34292 , n37564 );
    and g13435 ( n11443 , n32904 , n33358 );
    not g13436 ( n13742 , n24940 );
    and g13437 ( n25945 , n37194 , n32947 );
    or g13438 ( n20878 , n36660 , n7485 );
    not g13439 ( n13847 , n5409 );
    nor g13440 ( n39614 , n1507 , n11857 );
    not g13441 ( n12805 , n28843 );
    xnor g13442 ( n2037 , n8837 , n37072 );
    nor g13443 ( n18215 , n42792 , n3654 );
    or g13444 ( n15747 , n30192 , n9912 );
    not g13445 ( n40246 , n20131 );
    or g13446 ( n20417 , n36391 , n41641 );
    or g13447 ( n39695 , n39330 , n17548 );
    not g13448 ( n11374 , n5993 );
    or g13449 ( n32249 , n27577 , n25213 );
    xnor g13450 ( n16370 , n3053 , n28885 );
    not g13451 ( n39742 , n30438 );
    or g13452 ( n16546 , n12157 , n31593 );
    not g13453 ( n30754 , n24510 );
    or g13454 ( n23347 , n6455 , n21020 );
    and g13455 ( n25637 , n2963 , n17133 );
    and g13456 ( n42620 , n36144 , n37443 );
    and g13457 ( n710 , n21799 , n12986 );
    or g13458 ( n11080 , n6628 , n8934 );
    or g13459 ( n31229 , n7511 , n13000 );
    or g13460 ( n25214 , n16211 , n4356 );
    or g13461 ( n36933 , n39460 , n18070 );
    nor g13462 ( n40097 , n30420 , n33898 );
    or g13463 ( n38129 , n10530 , n16502 );
    or g13464 ( n32593 , n26212 , n19491 );
    or g13465 ( n5876 , n9733 , n34938 );
    and g13466 ( n8234 , n31492 , n16295 );
    or g13467 ( n31029 , n14776 , n32141 );
    and g13468 ( n13370 , n35506 , n2833 );
    or g13469 ( n20334 , n31975 , n4151 );
    or g13470 ( n8272 , n3981 , n5666 );
    or g13471 ( n13189 , n22850 , n21950 );
    xnor g13472 ( n12476 , n16693 , n30412 );
    not g13473 ( n29948 , n2358 );
    not g13474 ( n19522 , n19629 );
    or g13475 ( n27290 , n12587 , n2680 );
    or g13476 ( n13410 , n20138 , n18442 );
    or g13477 ( n25560 , n17000 , n38293 );
    or g13478 ( n28635 , n6510 , n41335 );
    and g13479 ( n10879 , n38203 , n38440 );
    nor g13480 ( n23593 , n24161 , n18619 );
    nor g13481 ( n37682 , n18131 , n22275 );
    and g13482 ( n26699 , n27012 , n11704 );
    or g13483 ( n24333 , n29455 , n2440 );
    or g13484 ( n34958 , n10088 , n2777 );
    nor g13485 ( n25566 , n35301 , n12913 );
    and g13486 ( n42391 , n24914 , n28424 );
    and g13487 ( n24840 , n5686 , n26015 );
    and g13488 ( n29829 , n7731 , n11556 );
    and g13489 ( n42195 , n6631 , n3011 );
    and g13490 ( n28086 , n4133 , n22975 );
    not g13491 ( n7035 , n29089 );
    and g13492 ( n14877 , n41459 , n27143 );
    or g13493 ( n27885 , n40426 , n20261 );
    and g13494 ( n2755 , n12796 , n22412 );
    nor g13495 ( n27457 , n14364 , n34324 );
    or g13496 ( n41105 , n30662 , n19702 );
    or g13497 ( n34615 , n29969 , n23760 );
    and g13498 ( n10462 , n430 , n37914 );
    nor g13499 ( n23176 , n37907 , n31714 );
    or g13500 ( n5970 , n42223 , n26219 );
    xnor g13501 ( n17498 , n37276 , n40171 );
    or g13502 ( n2558 , n31480 , n30446 );
    xnor g13503 ( n21318 , n36009 , n32668 );
    not g13504 ( n17872 , n36309 );
    and g13505 ( n16311 , n30323 , n11741 );
    xnor g13506 ( n26544 , n39432 , n25107 );
    xnor g13507 ( n33091 , n36998 , n23140 );
    and g13508 ( n12683 , n12390 , n26381 );
    xnor g13509 ( n26220 , n21448 , n26780 );
    xnor g13510 ( n6194 , n27721 , n29770 );
    or g13511 ( n17328 , n33295 , n28436 );
    or g13512 ( n8554 , n11267 , n3134 );
    and g13513 ( n10626 , n18949 , n3584 );
    nor g13514 ( n20388 , n14696 , n35153 );
    or g13515 ( n7998 , n32711 , n12219 );
    and g13516 ( n1340 , n955 , n18341 );
    xnor g13517 ( n22607 , n36009 , n32549 );
    not g13518 ( n41360 , n2981 );
    or g13519 ( n33779 , n35294 , n22307 );
    or g13520 ( n24811 , n3807 , n38326 );
    nor g13521 ( n31005 , n18866 , n2464 );
    not g13522 ( n19186 , n29715 );
    and g13523 ( n3092 , n20070 , n3327 );
    or g13524 ( n26905 , n19196 , n22688 );
    or g13525 ( n909 , n16564 , n8169 );
    not g13526 ( n2900 , n29792 );
    and g13527 ( n18870 , n25339 , n35480 );
    and g13528 ( n16690 , n3345 , n29081 );
    xnor g13529 ( n28952 , n39921 , n27062 );
    and g13530 ( n31806 , n12460 , n12396 );
    or g13531 ( n12478 , n969 , n3346 );
    and g13532 ( n24755 , n13192 , n37382 );
    xnor g13533 ( n38131 , n25582 , n20521 );
    or g13534 ( n11223 , n28029 , n26277 );
    and g13535 ( n37123 , n9674 , n36750 );
    or g13536 ( n2928 , n21857 , n5348 );
    or g13537 ( n30901 , n21665 , n25907 );
    not g13538 ( n37808 , n23963 );
    nor g13539 ( n22898 , n33716 , n37554 );
    or g13540 ( n24337 , n3287 , n4965 );
    or g13541 ( n42571 , n14266 , n9684 );
    or g13542 ( n37507 , n1866 , n35737 );
    and g13543 ( n33900 , n1646 , n38083 );
    not g13544 ( n36657 , n16677 );
    and g13545 ( n26646 , n29781 , n21658 );
    or g13546 ( n28124 , n39341 , n6209 );
    or g13547 ( n31790 , n15565 , n5277 );
    or g13548 ( n26756 , n32711 , n26780 );
    not g13549 ( n37074 , n36939 );
    nor g13550 ( n15339 , n13046 , n25228 );
    not g13551 ( n40757 , n32814 );
    or g13552 ( n25491 , n2142 , n24607 );
    nor g13553 ( n4579 , n13481 , n35199 );
    xnor g13554 ( n35680 , n38371 , n1063 );
    nor g13555 ( n21272 , n35074 , n6990 );
    not g13556 ( n25407 , n8407 );
    or g13557 ( n38586 , n38022 , n3370 );
    or g13558 ( n7586 , n5605 , n30610 );
    not g13559 ( n1432 , n37507 );
    nor g13560 ( n26536 , n14105 , n12726 );
    or g13561 ( n11959 , n13565 , n16084 );
    or g13562 ( n19148 , n23337 , n22355 );
    or g13563 ( n26697 , n30896 , n25702 );
    and g13564 ( n28457 , n37729 , n4734 );
    not g13565 ( n34654 , n23915 );
    and g13566 ( n30971 , n29499 , n10055 );
    xnor g13567 ( n17163 , n784 , n35662 );
    and g13568 ( n35852 , n41745 , n17648 );
    not g13569 ( n41079 , n6032 );
    not g13570 ( n20628 , n32388 );
    not g13571 ( n33671 , n32679 );
    nor g13572 ( n20826 , n17744 , n22157 );
    and g13573 ( n29334 , n12680 , n21369 );
    and g13574 ( n13851 , n4113 , n27622 );
    or g13575 ( n37302 , n33349 , n25940 );
    and g13576 ( n41111 , n15115 , n21104 );
    not g13577 ( n6878 , n20358 );
    xnor g13578 ( n4055 , n29740 , n22131 );
    and g13579 ( n33267 , n31846 , n41142 );
    and g13580 ( n9547 , n6649 , n11518 );
    or g13581 ( n2305 , n31003 , n38437 );
    and g13582 ( n20545 , n38116 , n27587 );
    or g13583 ( n13344 , n38407 , n30793 );
    or g13584 ( n26526 , n38119 , n22052 );
    not g13585 ( n5362 , n2681 );
    or g13586 ( n15313 , n5126 , n22752 );
    or g13587 ( n40901 , n2249 , n34206 );
    and g13588 ( n29800 , n35585 , n3300 );
    nor g13589 ( n26416 , n13181 , n6711 );
    or g13590 ( n687 , n14377 , n10467 );
    and g13591 ( n13944 , n7010 , n4295 );
    not g13592 ( n37723 , n19624 );
    not g13593 ( n14556 , n11153 );
    nor g13594 ( n19789 , n31274 , n28146 );
    nor g13595 ( n5771 , n35790 , n29288 );
    nor g13596 ( n8669 , n25775 , n13223 );
    and g13597 ( n23655 , n25799 , n35658 );
    xnor g13598 ( n42092 , n4901 , n35301 );
    nor g13599 ( n28208 , n22588 , n12337 );
    or g13600 ( n10122 , n29027 , n12601 );
    and g13601 ( n33772 , n29589 , n41125 );
    or g13602 ( n39220 , n15098 , n38196 );
    not g13603 ( n36962 , n34880 );
    or g13604 ( n20960 , n11087 , n21245 );
    or g13605 ( n6103 , n4121 , n1849 );
    or g13606 ( n8566 , n39208 , n23716 );
    or g13607 ( n33360 , n29598 , n38996 );
    nor g13608 ( n2388 , n19186 , n13469 );
    not g13609 ( n22772 , n9563 );
    not g13610 ( n31096 , n36724 );
    or g13611 ( n42126 , n29058 , n8468 );
    or g13612 ( n37492 , n25810 , n23591 );
    or g13613 ( n16450 , n34997 , n16166 );
    nor g13614 ( n31446 , n9275 , n15248 );
    or g13615 ( n11097 , n20848 , n22797 );
    or g13616 ( n37318 , n18646 , n10275 );
    not g13617 ( n6330 , n15967 );
    and g13618 ( n17332 , n1926 , n16530 );
    not g13619 ( n3416 , n2814 );
    nor g13620 ( n651 , n15070 , n646 );
    and g13621 ( n19479 , n27011 , n39370 );
    or g13622 ( n19666 , n30460 , n30652 );
    or g13623 ( n21474 , n4954 , n34576 );
    or g13624 ( n25334 , n23434 , n31255 );
    or g13625 ( n5757 , n41526 , n2776 );
    or g13626 ( n16974 , n25903 , n16209 );
    or g13627 ( n40919 , n37277 , n328 );
    nor g13628 ( n23758 , n6303 , n27326 );
    or g13629 ( n42861 , n3257 , n30462 );
    and g13630 ( n31447 , n34097 , n4248 );
    nor g13631 ( n6301 , n14598 , n2257 );
    or g13632 ( n15431 , n18912 , n20498 );
    nor g13633 ( n41861 , n16540 , n20439 );
    or g13634 ( n1112 , n10653 , n31412 );
    nor g13635 ( n21618 , n3061 , n3624 );
    and g13636 ( n10619 , n34758 , n6887 );
    or g13637 ( n31470 , n8005 , n21825 );
    nor g13638 ( n16414 , n27811 , n36594 );
    or g13639 ( n4819 , n15688 , n33775 );
    and g13640 ( n28857 , n5144 , n10738 );
    and g13641 ( n9443 , n8532 , n28033 );
    and g13642 ( n11492 , n30761 , n15587 );
    or g13643 ( n30618 , n18645 , n3142 );
    or g13644 ( n5333 , n26849 , n36540 );
    or g13645 ( n41060 , n35375 , n6024 );
    and g13646 ( n20784 , n39266 , n29145 );
    or g13647 ( n10236 , n38947 , n11591 );
    not g13648 ( n21067 , n5786 );
    and g13649 ( n1183 , n27557 , n42315 );
    and g13650 ( n21267 , n23813 , n37644 );
    and g13651 ( n17474 , n32612 , n35774 );
    or g13652 ( n23684 , n23776 , n37580 );
    and g13653 ( n28562 , n23486 , n33757 );
    not g13654 ( n8253 , n802 );
    or g13655 ( n10505 , n23103 , n38888 );
    xnor g13656 ( n34426 , n41098 , n18808 );
    xnor g13657 ( n31080 , n784 , n11071 );
    nor g13658 ( n42015 , n35301 , n26301 );
    or g13659 ( n35006 , n35550 , n30435 );
    xnor g13660 ( n42270 , n24524 , n28730 );
    and g13661 ( n15106 , n14488 , n40641 );
    and g13662 ( n23463 , n19048 , n32166 );
    and g13663 ( n12914 , n36617 , n34149 );
    or g13664 ( n24074 , n35822 , n16249 );
    and g13665 ( n12219 , n41209 , n15915 );
    xnor g13666 ( n16708 , n40 , n22683 );
    not g13667 ( n22169 , n493 );
    not g13668 ( n6374 , n39090 );
    not g13669 ( n41650 , n10281 );
    and g13670 ( n4928 , n8843 , n27177 );
    or g13671 ( n1711 , n31263 , n7749 );
    xnor g13672 ( n28118 , n41715 , n16990 );
    not g13673 ( n30405 , n42915 );
    or g13674 ( n33009 , n22654 , n5589 );
    or g13675 ( n26469 , n17025 , n24063 );
    nor g13676 ( n19843 , n33053 , n2354 );
    xnor g13677 ( n38324 , n36998 , n28483 );
    or g13678 ( n22970 , n5140 , n21047 );
    or g13679 ( n31169 , n38494 , n8901 );
    nor g13680 ( n24513 , n41534 , n10832 );
    and g13681 ( n29134 , n24321 , n12116 );
    not g13682 ( n42127 , n26650 );
    and g13683 ( n29320 , n22494 , n40440 );
    or g13684 ( n9545 , n42420 , n11545 );
    or g13685 ( n13706 , n14112 , n23902 );
    not g13686 ( n9977 , n2562 );
    or g13687 ( n13871 , n23059 , n15801 );
    nor g13688 ( n24367 , n19580 , n10690 );
    and g13689 ( n1659 , n36347 , n9257 );
    not g13690 ( n6500 , n16551 );
    nor g13691 ( n25659 , n38469 , n42347 );
    and g13692 ( n31371 , n20931 , n39820 );
    or g13693 ( n36740 , n5964 , n13464 );
    or g13694 ( n29500 , n405 , n26600 );
    and g13695 ( n26975 , n22034 , n30778 );
    and g13696 ( n25762 , n13166 , n20216 );
    xnor g13697 ( n892 , n13735 , n28701 );
    nor g13698 ( n40587 , n39640 , n932 );
    not g13699 ( n17819 , n36056 );
    and g13700 ( n39506 , n30537 , n5488 );
    nor g13701 ( n8543 , n38542 , n9152 );
    and g13702 ( n31030 , n21749 , n30102 );
    nor g13703 ( n36363 , n17371 , n9138 );
    nor g13704 ( n650 , n32807 , n11482 );
    or g13705 ( n12043 , n7375 , n6937 );
    and g13706 ( n42160 , n11878 , n1660 );
    or g13707 ( n21083 , n10898 , n41774 );
    and g13708 ( n36459 , n289 , n17887 );
    or g13709 ( n32464 , n5808 , n35036 );
    not g13710 ( n33134 , n40720 );
    or g13711 ( n39785 , n19366 , n16529 );
    not g13712 ( n2569 , n17512 );
    or g13713 ( n36404 , n123 , n33017 );
    not g13714 ( n6019 , n24929 );
    not g13715 ( n1057 , n29081 );
    and g13716 ( n11829 , n247 , n35482 );
    and g13717 ( n10832 , n28790 , n34028 );
    xnor g13718 ( n28559 , n8597 , n13567 );
    and g13719 ( n24612 , n32496 , n14162 );
    or g13720 ( n4500 , n2095 , n38572 );
    or g13721 ( n18960 , n1009 , n16989 );
    not g13722 ( n17182 , n6065 );
    and g13723 ( n36618 , n2890 , n6151 );
    nor g13724 ( n24844 , n8790 , n23496 );
    or g13725 ( n10079 , n31265 , n40056 );
    and g13726 ( n2312 , n13911 , n28923 );
    xnor g13727 ( n32000 , n32794 , n40509 );
    or g13728 ( n39089 , n34527 , n26019 );
    or g13729 ( n36562 , n38201 , n8587 );
    nor g13730 ( n33754 , n25060 , n8297 );
    or g13731 ( n20973 , n17947 , n25490 );
    or g13732 ( n10171 , n6454 , n35702 );
    xnor g13733 ( n32209 , n33287 , n18866 );
    xnor g13734 ( n12463 , n35928 , n14471 );
    not g13735 ( n14735 , n14162 );
    not g13736 ( n41381 , n12453 );
    or g13737 ( n14938 , n13517 , n684 );
    and g13738 ( n19066 , n29202 , n41800 );
    or g13739 ( n28196 , n1335 , n7780 );
    or g13740 ( n19356 , n34545 , n15232 );
    nor g13741 ( n29484 , n39896 , n19313 );
    and g13742 ( n26879 , n1278 , n27368 );
    and g13743 ( n27130 , n26618 , n14073 );
    or g13744 ( n8366 , n23599 , n4357 );
    xnor g13745 ( n8673 , n40 , n42302 );
    or g13746 ( n1579 , n24365 , n20048 );
    and g13747 ( n19333 , n40196 , n11018 );
    not g13748 ( n19538 , n3194 );
    and g13749 ( n13514 , n14320 , n3529 );
    or g13750 ( n29804 , n8994 , n26845 );
    or g13751 ( n41273 , n31580 , n20543 );
    nor g13752 ( n32477 , n5724 , n26243 );
    or g13753 ( n285 , n21054 , n810 );
    nor g13754 ( n41262 , n21653 , n30291 );
    or g13755 ( n26278 , n40808 , n13229 );
    not g13756 ( n15972 , n36526 );
    xnor g13757 ( n32608 , n32000 , n3319 );
    nor g13758 ( n3071 , n36798 , n8673 );
    and g13759 ( n40577 , n2251 , n7804 );
    xnor g13760 ( n32570 , n21301 , n17509 );
    not g13761 ( n20237 , n6161 );
    or g13762 ( n34532 , n22974 , n36000 );
    or g13763 ( n993 , n24035 , n34094 );
    not g13764 ( n30295 , n13523 );
    and g13765 ( n32894 , n32047 , n39234 );
    nor g13766 ( n26087 , n8439 , n933 );
    not g13767 ( n38149 , n22415 );
    nor g13768 ( n17687 , n33981 , n576 );
    not g13769 ( n12639 , n19503 );
    and g13770 ( n30123 , n21534 , n27246 );
    or g13771 ( n24161 , n24246 , n21207 );
    or g13772 ( n6165 , n41150 , n29545 );
    nor g13773 ( n3809 , n6246 , n15730 );
    not g13774 ( n33915 , n41321 );
    or g13775 ( n26815 , n17393 , n13576 );
    or g13776 ( n26249 , n7953 , n31608 );
    or g13777 ( n28858 , n328 , n39344 );
    and g13778 ( n4039 , n17958 , n10091 );
    not g13779 ( n4308 , n30997 );
    not g13780 ( n11960 , n19582 );
    xnor g13781 ( n39792 , n27035 , n35127 );
    xnor g13782 ( n39613 , n22103 , n22297 );
    xnor g13783 ( n25057 , n22604 , n2354 );
    or g13784 ( n40005 , n38711 , n27856 );
    or g13785 ( n9140 , n36038 , n40554 );
    or g13786 ( n33284 , n20826 , n4283 );
    or g13787 ( n1000 , n41560 , n35791 );
    not g13788 ( n18673 , n3631 );
    nor g13789 ( n32029 , n32731 , n37984 );
    or g13790 ( n33789 , n26752 , n33553 );
    or g13791 ( n10193 , n37837 , n40419 );
    or g13792 ( n23704 , n5324 , n338 );
    or g13793 ( n3674 , n23788 , n30129 );
    or g13794 ( n5368 , n21428 , n20462 );
    and g13795 ( n322 , n34709 , n23157 );
    and g13796 ( n18206 , n16463 , n36190 );
    not g13797 ( n1002 , n14004 );
    nor g13798 ( n38250 , n14808 , n5375 );
    and g13799 ( n13552 , n22053 , n36386 );
    and g13800 ( n29082 , n16061 , n31951 );
    nor g13801 ( n19973 , n12158 , n11541 );
    and g13802 ( n8582 , n15018 , n21017 );
    nor g13803 ( n36755 , n20851 , n39553 );
    xnor g13804 ( n5354 , n34810 , n39775 );
    not g13805 ( n17454 , n9682 );
    not g13806 ( n17420 , n11574 );
    and g13807 ( n42404 , n8724 , n35176 );
    xnor g13808 ( n2723 , n16320 , n17166 );
    or g13809 ( n35555 , n31762 , n1012 );
    xnor g13810 ( n6828 , n40701 , n9657 );
    not g13811 ( n25187 , n19307 );
    not g13812 ( n2088 , n13663 );
    and g13813 ( n34199 , n37369 , n14486 );
    nor g13814 ( n21687 , n32262 , n2257 );
    or g13815 ( n24014 , n9602 , n35362 );
    and g13816 ( n28684 , n31308 , n29390 );
    or g13817 ( n2119 , n10908 , n28335 );
    or g13818 ( n39762 , n25685 , n27296 );
    not g13819 ( n41215 , n5661 );
    or g13820 ( n31296 , n2016 , n29388 );
    xnor g13821 ( n17537 , n26579 , n31466 );
    or g13822 ( n21623 , n13176 , n5774 );
    nor g13823 ( n37621 , n36654 , n28621 );
    xnor g13824 ( n1066 , n16822 , n29853 );
    and g13825 ( n20883 , n7540 , n27351 );
    not g13826 ( n3457 , n39487 );
    or g13827 ( n25418 , n8207 , n32892 );
    not g13828 ( n6221 , n21739 );
    xnor g13829 ( n24577 , n31989 , n14686 );
    or g13830 ( n9148 , n964 , n9819 );
    and g13831 ( n16529 , n11256 , n32758 );
    and g13832 ( n16538 , n33855 , n37104 );
    or g13833 ( n31598 , n19217 , n25560 );
    or g13834 ( n18620 , n2701 , n31530 );
    and g13835 ( n37372 , n5171 , n30781 );
    or g13836 ( n1753 , n10081 , n39098 );
    not g13837 ( n38954 , n13708 );
    nor g13838 ( n6083 , n32277 , n22696 );
    and g13839 ( n30043 , n6433 , n36133 );
    not g13840 ( n34223 , n18039 );
    or g13841 ( n5748 , n28880 , n31119 );
    or g13842 ( n19255 , n28389 , n2908 );
    xnor g13843 ( n17893 , n10024 , n28920 );
    or g13844 ( n24041 , n7485 , n5363 );
    or g13845 ( n19797 , n35452 , n34160 );
    and g13846 ( n42893 , n39189 , n19906 );
    or g13847 ( n20117 , n18935 , n16309 );
    and g13848 ( n38507 , n20095 , n23662 );
    and g13849 ( n29996 , n6860 , n10127 );
    not g13850 ( n5398 , n29094 );
    or g13851 ( n27160 , n16143 , n35332 );
    or g13852 ( n27970 , n35748 , n41420 );
    xnor g13853 ( n29150 , n30251 , n34565 );
    nor g13854 ( n31704 , n35301 , n39884 );
    or g13855 ( n21348 , n23082 , n10075 );
    xnor g13856 ( n13123 , n13041 , n6188 );
    nor g13857 ( n10768 , n14277 , n28952 );
    or g13858 ( n19222 , n37616 , n24068 );
    and g13859 ( n37674 , n11497 , n33015 );
    or g13860 ( n24417 , n33537 , n28532 );
    or g13861 ( n17235 , n18986 , n34436 );
    and g13862 ( n21020 , n26666 , n20132 );
    or g13863 ( n39283 , n5565 , n22409 );
    or g13864 ( n9622 , n39195 , n118 );
    or g13865 ( n22043 , n22091 , n39928 );
    xnor g13866 ( n17672 , n40886 , n20359 );
    or g13867 ( n27830 , n2232 , n33680 );
    not g13868 ( n12381 , n26492 );
    or g13869 ( n11704 , n21018 , n28031 );
    or g13870 ( n2359 , n17197 , n19329 );
    and g13871 ( n17053 , n25524 , n19257 );
    xnor g13872 ( n12661 , n24034 , n14097 );
    not g13873 ( n18675 , n8616 );
    or g13874 ( n19011 , n1917 , n23457 );
    or g13875 ( n9648 , n26276 , n38191 );
    not g13876 ( n17449 , n12483 );
    xnor g13877 ( n12325 , n18939 , n4210 );
    xnor g13878 ( n7277 , n3068 , n42751 );
    and g13879 ( n37506 , n10794 , n41196 );
    not g13880 ( n14740 , n7221 );
    and g13881 ( n14634 , n17305 , n38002 );
    and g13882 ( n6954 , n15836 , n10250 );
    and g13883 ( n33353 , n16696 , n20925 );
    nor g13884 ( n11907 , n1917 , n27337 );
    nor g13885 ( n40599 , n3769 , n37706 );
    and g13886 ( n2870 , n1920 , n35846 );
    and g13887 ( n5997 , n3647 , n20609 );
    and g13888 ( n29477 , n30823 , n41664 );
    or g13889 ( n42401 , n14201 , n15912 );
    not g13890 ( n17173 , n36110 );
    nor g13891 ( n40733 , n3769 , n11105 );
    or g13892 ( n26388 , n7840 , n4227 );
    or g13893 ( n41101 , n27851 , n11178 );
    or g13894 ( n6735 , n18424 , n18394 );
    xnor g13895 ( n8894 , n40 , n7921 );
    and g13896 ( n7710 , n13869 , n18191 );
    and g13897 ( n35470 , n30429 , n30464 );
    not g13898 ( n42042 , n31965 );
    or g13899 ( n29262 , n10885 , n1581 );
    not g13900 ( n41480 , n25738 );
    and g13901 ( n26305 , n13269 , n21785 );
    and g13902 ( n35362 , n34973 , n35326 );
    xnor g13903 ( n27426 , n42151 , n29386 );
    nor g13904 ( n14122 , n30295 , n21812 );
    or g13905 ( n2070 , n4949 , n39399 );
    not g13906 ( n20952 , n19014 );
    or g13907 ( n18467 , n3620 , n2589 );
    nor g13908 ( n9943 , n6349 , n14999 );
    not g13909 ( n13368 , n29117 );
    or g13910 ( n36743 , n25267 , n39250 );
    and g13911 ( n2322 , n32571 , n25083 );
    not g13912 ( n38860 , n21905 );
    not g13913 ( n23218 , n9786 );
    or g13914 ( n26218 , n14418 , n5520 );
    and g13915 ( n1329 , n16822 , n29853 );
    xnor g13916 ( n40532 , n20310 , n14677 );
    or g13917 ( n31800 , n17658 , n8035 );
    nor g13918 ( n13397 , n34816 , n11577 );
    or g13919 ( n8285 , n2231 , n10997 );
    or g13920 ( n29904 , n41601 , n13278 );
    not g13921 ( n12942 , n21643 );
    not g13922 ( n22807 , n19039 );
    xnor g13923 ( n19959 , n20548 , n41387 );
    and g13924 ( n34976 , n17507 , n32533 );
    or g13925 ( n4250 , n23253 , n34972 );
    not g13926 ( n26919 , n31067 );
    or g13927 ( n13227 , n42190 , n34774 );
    not g13928 ( n33691 , n16702 );
    and g13929 ( n38945 , n22407 , n34396 );
    or g13930 ( n23520 , n24656 , n11446 );
    or g13931 ( n20017 , n7227 , n35531 );
    or g13932 ( n7290 , n37131 , n28928 );
    xnor g13933 ( n4525 , n36973 , n28216 );
    xnor g13934 ( n27771 , n35367 , n39451 );
    and g13935 ( n11828 , n8085 , n39836 );
    and g13936 ( n39295 , n26674 , n1154 );
    or g13937 ( n31650 , n5964 , n26342 );
    and g13938 ( n36786 , n36412 , n26198 );
    or g13939 ( n5595 , n6666 , n28538 );
    and g13940 ( n31428 , n40083 , n22116 );
    nor g13941 ( n4473 , n12302 , n5055 );
    xnor g13942 ( n38652 , n36009 , n16095 );
    or g13943 ( n42564 , n3447 , n28348 );
    and g13944 ( n26245 , n13859 , n17483 );
    and g13945 ( n13093 , n15849 , n4235 );
    or g13946 ( n11428 , n38967 , n12127 );
    not g13947 ( n10011 , n36776 );
    xnor g13948 ( n34827 , n41500 , n14751 );
    not g13949 ( n39264 , n31741 );
    not g13950 ( n12656 , n25417 );
    not g13951 ( n25440 , n26969 );
    not g13952 ( n25704 , n8588 );
    and g13953 ( n24785 , n3857 , n7932 );
    and g13954 ( n3234 , n36730 , n33921 );
    xnor g13955 ( n44 , n40 , n9452 );
    and g13956 ( n19026 , n16907 , n4 );
    or g13957 ( n17245 , n2416 , n8637 );
    or g13958 ( n32116 , n29717 , n37621 );
    or g13959 ( n33896 , n9194 , n25264 );
    or g13960 ( n25633 , n1997 , n13464 );
    or g13961 ( n6285 , n17108 , n15160 );
    and g13962 ( n22372 , n16983 , n16682 );
    and g13963 ( n31303 , n36867 , n33087 );
    and g13964 ( n42240 , n31069 , n12012 );
    or g13965 ( n16865 , n15580 , n9771 );
    nor g13966 ( n30013 , n25871 , n17007 );
    xnor g13967 ( n30911 , n16106 , n40909 );
    nor g13968 ( n35835 , n32981 , n15326 );
    nor g13969 ( n17448 , n10676 , n15863 );
    xnor g13970 ( n40037 , n31956 , n21203 );
    not g13971 ( n7965 , n39789 );
    nor g13972 ( n42777 , n17744 , n25656 );
    and g13973 ( n19847 , n1308 , n26451 );
    or g13974 ( n10305 , n36094 , n39723 );
    or g13975 ( n24481 , n5324 , n34804 );
    and g13976 ( n6393 , n30624 , n20586 );
    nor g13977 ( n30937 , n23811 , n25921 );
    and g13978 ( n2464 , n27748 , n26779 );
    or g13979 ( n37991 , n40439 , n2951 );
    not g13980 ( n3139 , n30463 );
    or g13981 ( n41875 , n1617 , n8530 );
    or g13982 ( n15724 , n37494 , n1407 );
    not g13983 ( n37081 , n30074 );
    or g13984 ( n18312 , n1238 , n42642 );
    not g13985 ( n16705 , n690 );
    and g13986 ( n11755 , n28752 , n36035 );
    or g13987 ( n14103 , n991 , n29497 );
    xnor g13988 ( n36346 , n22054 , n22024 );
    or g13989 ( n24803 , n17162 , n1044 );
    and g13990 ( n12136 , n3473 , n30242 );
    not g13991 ( n40197 , n33978 );
    not g13992 ( n10427 , n32667 );
    xnor g13993 ( n38738 , n33917 , n26578 );
    or g13994 ( n30928 , n4085 , n4245 );
    not g13995 ( n597 , n13994 );
    or g13996 ( n37261 , n17754 , n15780 );
    or g13997 ( n8365 , n30192 , n14836 );
    or g13998 ( n31946 , n2185 , n12392 );
    not g13999 ( n24760 , n29816 );
    xnor g14000 ( n42626 , n13108 , n36816 );
    or g14001 ( n26645 , n39439 , n9159 );
    xnor g14002 ( n38732 , n142 , n17939 );
    xnor g14003 ( n17471 , n34562 , n8997 );
    not g14004 ( n27010 , n4178 );
    and g14005 ( n25940 , n29783 , n24456 );
    and g14006 ( n7243 , n26082 , n41851 );
    and g14007 ( n38117 , n30049 , n12719 );
    and g14008 ( n35260 , n36398 , n29237 );
    or g14009 ( n28265 , n22872 , n33930 );
    or g14010 ( n29507 , n7139 , n22375 );
    not g14011 ( n38504 , n27463 );
    nor g14012 ( n10584 , n2292 , n207 );
    or g14013 ( n24938 , n734 , n23174 );
    or g14014 ( n33886 , n10311 , n8380 );
    or g14015 ( n1508 , n10190 , n15299 );
    and g14016 ( n37628 , n7738 , n3449 );
    nor g14017 ( n6389 , n22519 , n4699 );
    not g14018 ( n42515 , n13140 );
    or g14019 ( n18940 , n2193 , n39572 );
    or g14020 ( n31882 , n32812 , n38913 );
    or g14021 ( n2047 , n18535 , n28947 );
    not g14022 ( n13367 , n9492 );
    not g14023 ( n11534 , n40753 );
    or g14024 ( n38390 , n24283 , n13057 );
    and g14025 ( n32208 , n29153 , n20927 );
    nor g14026 ( n35204 , n20173 , n18532 );
    nor g14027 ( n36027 , n19903 , n41789 );
    nor g14028 ( n20051 , n1359 , n40523 );
    or g14029 ( n26556 , n37804 , n41999 );
    and g14030 ( n41405 , n24512 , n10487 );
    or g14031 ( n27893 , n29900 , n37789 );
    not g14032 ( n8873 , n23170 );
    and g14033 ( n5570 , n25041 , n16546 );
    nor g14034 ( n41388 , n17188 , n21462 );
    or g14035 ( n8879 , n5351 , n4358 );
    not g14036 ( n27478 , n34654 );
    or g14037 ( n34683 , n15429 , n23993 );
    nor g14038 ( n41181 , n41766 , n20887 );
    or g14039 ( n39913 , n31618 , n2845 );
    or g14040 ( n14196 , n15946 , n11132 );
    and g14041 ( n1167 , n36017 , n20466 );
    or g14042 ( n33524 , n19511 , n18188 );
    and g14043 ( n11537 , n42170 , n8028 );
    or g14044 ( n39860 , n14407 , n7774 );
    xnor g14045 ( n36613 , n1224 , n23931 );
    or g14046 ( n2156 , n19471 , n13236 );
    and g14047 ( n21 , n37148 , n29727 );
    not g14048 ( n32829 , n24941 );
    nor g14049 ( n24780 , n36636 , n31011 );
    or g14050 ( n41366 , n16229 , n21268 );
    not g14051 ( n24186 , n4952 );
    and g14052 ( n38825 , n18223 , n36362 );
    or g14053 ( n37377 , n23491 , n23618 );
    and g14054 ( n40252 , n33300 , n40594 );
    or g14055 ( n32672 , n16331 , n41644 );
    or g14056 ( n13162 , n3801 , n24801 );
    and g14057 ( n30725 , n10256 , n20926 );
    and g14058 ( n697 , n36047 , n8733 );
    xnor g14059 ( n23784 , n17165 , n14707 );
    and g14060 ( n1067 , n29705 , n34299 );
    or g14061 ( n709 , n10460 , n31807 );
    or g14062 ( n5196 , n18727 , n34976 );
    or g14063 ( n8102 , n19811 , n1888 );
    xnor g14064 ( n39719 , n4604 , n29085 );
    and g14065 ( n13807 , n34801 , n30441 );
    or g14066 ( n9587 , n31258 , n38715 );
    or g14067 ( n10431 , n32605 , n36857 );
    xnor g14068 ( n15891 , n10527 , n6711 );
    or g14069 ( n20275 , n1178 , n21527 );
    not g14070 ( n951 , n30205 );
    xnor g14071 ( n21007 , n17909 , n14155 );
    not g14072 ( n23735 , n3671 );
    not g14073 ( n6658 , n6968 );
    nor g14074 ( n6707 , n10152 , n17120 );
    or g14075 ( n41989 , n6978 , n20196 );
    or g14076 ( n18122 , n19035 , n17092 );
    or g14077 ( n36282 , n34411 , n5651 );
    and g14078 ( n2899 , n5530 , n42500 );
    nor g14079 ( n3427 , n34358 , n6039 );
    or g14080 ( n2808 , n36296 , n18349 );
    xnor g14081 ( n18020 , n9401 , n13119 );
    or g14082 ( n39272 , n13239 , n35514 );
    or g14083 ( n39154 , n29513 , n29748 );
    or g14084 ( n17132 , n18426 , n34972 );
    or g14085 ( n27723 , n33926 , n30031 );
    or g14086 ( n4164 , n16382 , n2296 );
    not g14087 ( n31125 , n31840 );
    or g14088 ( n28606 , n4645 , n15039 );
    nor g14089 ( n25830 , n17120 , n31186 );
    not g14090 ( n2710 , n41578 );
    and g14091 ( n35304 , n40700 , n33800 );
    and g14092 ( n28594 , n13715 , n25731 );
    and g14093 ( n35370 , n32756 , n23025 );
    not g14094 ( n7020 , n13615 );
    not g14095 ( n12945 , n18201 );
    not g14096 ( n19116 , n27964 );
    and g14097 ( n20003 , n23095 , n22806 );
    or g14098 ( n12110 , n27503 , n26860 );
    nor g14099 ( n15927 , n38836 , n14829 );
    nor g14100 ( n37638 , n16728 , n32 );
    xnor g14101 ( n9502 , n19052 , n24611 );
    not g14102 ( n39732 , n21504 );
    or g14103 ( n35971 , n8136 , n10381 );
    nor g14104 ( n23692 , n15080 , n27954 );
    not g14105 ( n38068 , n34579 );
    and g14106 ( n7065 , n18669 , n32569 );
    nor g14107 ( n10260 , n34429 , n41373 );
    not g14108 ( n30403 , n17660 );
    or g14109 ( n12516 , n33288 , n17296 );
    or g14110 ( n32651 , n5884 , n30137 );
    and g14111 ( n16923 , n13829 , n30673 );
    or g14112 ( n3742 , n26970 , n18935 );
    nor g14113 ( n40994 , n9607 , n10821 );
    or g14114 ( n21329 , n34255 , n7956 );
    or g14115 ( n21237 , n36071 , n1704 );
    or g14116 ( n20815 , n26865 , n37415 );
    nor g14117 ( n26217 , n18866 , n18770 );
    and g14118 ( n4477 , n40156 , n35449 );
    or g14119 ( n27839 , n40293 , n16733 );
    nor g14120 ( n37471 , n12106 , n36148 );
    nor g14121 ( n13330 , n33850 , n42285 );
    or g14122 ( n40192 , n6385 , n2565 );
    and g14123 ( n12566 , n15821 , n9486 );
    xnor g14124 ( n30563 , n11596 , n34555 );
    or g14125 ( n35164 , n1110 , n13325 );
    or g14126 ( n23110 , n14898 , n24511 );
    not g14127 ( n23619 , n36132 );
    and g14128 ( n11947 , n29103 , n33400 );
    or g14129 ( n1751 , n202 , n29139 );
    or g14130 ( n27360 , n11417 , n5831 );
    not g14131 ( n11434 , n36309 );
    xnor g14132 ( n10360 , n24928 , n20316 );
    or g14133 ( n12548 , n40168 , n766 );
    or g14134 ( n6250 , n257 , n8035 );
    and g14135 ( n2089 , n18676 , n14580 );
    and g14136 ( n3765 , n38522 , n18497 );
    or g14137 ( n1262 , n5242 , n31943 );
    or g14138 ( n22590 , n40315 , n12196 );
    not g14139 ( n32408 , n39068 );
    or g14140 ( n9209 , n1453 , n11860 );
    and g14141 ( n36279 , n35408 , n18516 );
    nor g14142 ( n39847 , n15426 , n13524 );
    nor g14143 ( n7496 , n7356 , n7350 );
    or g14144 ( n35305 , n32963 , n38169 );
    nor g14145 ( n20219 , n29120 , n40784 );
    nor g14146 ( n4207 , n20871 , n17741 );
    not g14147 ( n9982 , n4358 );
    xnor g14148 ( n30107 , n36998 , n5541 );
    not g14149 ( n33870 , n32287 );
    xnor g14150 ( n36980 , n21534 , n25111 );
    and g14151 ( n41712 , n27168 , n32034 );
    and g14152 ( n19962 , n37286 , n12123 );
    or g14153 ( n14731 , n28942 , n6153 );
    or g14154 ( n2656 , n17862 , n22920 );
    not g14155 ( n27419 , n26749 );
    or g14156 ( n19297 , n28745 , n34197 );
    and g14157 ( n9621 , n15765 , n11689 );
    or g14158 ( n7396 , n7726 , n2565 );
    and g14159 ( n25702 , n38883 , n39232 );
    or g14160 ( n37432 , n25498 , n3868 );
    or g14161 ( n35077 , n1507 , n13194 );
    not g14162 ( n25625 , n1707 );
    or g14163 ( n1239 , n29980 , n1300 );
    nor g14164 ( n12508 , n7648 , n37116 );
    and g14165 ( n11546 , n26095 , n28194 );
    or g14166 ( n18918 , n4233 , n13495 );
    or g14167 ( n27939 , n33350 , n14944 );
    not g14168 ( n21480 , n40531 );
    xnor g14169 ( n32406 , n21309 , n14262 );
    xnor g14170 ( n13129 , n23478 , n23946 );
    not g14171 ( n10198 , n42235 );
    or g14172 ( n40546 , n25920 , n30795 );
    or g14173 ( n40810 , n5099 , n2643 );
    xnor g14174 ( n28563 , n13444 , n18827 );
    xnor g14175 ( n3640 , n2669 , n42628 );
    or g14176 ( n28697 , n17482 , n6057 );
    xnor g14177 ( n19346 , n23730 , n22113 );
    xnor g14178 ( n20789 , n10833 , n11978 );
    not g14179 ( n37863 , n37813 );
    nor g14180 ( n42305 , n1051 , n27834 );
    not g14181 ( n26253 , n15435 );
    or g14182 ( n638 , n19850 , n36161 );
    or g14183 ( n24302 , n8386 , n37733 );
    or g14184 ( n26687 , n28175 , n28666 );
    not g14185 ( n19868 , n19935 );
    or g14186 ( n24236 , n2608 , n6232 );
    and g14187 ( n26129 , n25942 , n27591 );
    and g14188 ( n32623 , n17676 , n11308 );
    or g14189 ( n27282 , n32415 , n33633 );
    not g14190 ( n30552 , n27754 );
    nor g14191 ( n16476 , n21347 , n5142 );
    and g14192 ( n9154 , n29357 , n27966 );
    or g14193 ( n36237 , n38505 , n26409 );
    and g14194 ( n27549 , n26877 , n7389 );
    xnor g14195 ( n23706 , n7943 , n39814 );
    and g14196 ( n5065 , n28681 , n10101 );
    and g14197 ( n33232 , n616 , n39990 );
    nor g14198 ( n6291 , n9240 , n13889 );
    not g14199 ( n17122 , n24398 );
    not g14200 ( n16389 , n24805 );
    and g14201 ( n17101 , n12501 , n4687 );
    and g14202 ( n1261 , n23617 , n4170 );
    xnor g14203 ( n2999 , n14643 , n5964 );
    nor g14204 ( n5900 , n42286 , n17150 );
    xnor g14205 ( n38882 , n19107 , n14505 );
    xnor g14206 ( n31 , n40902 , n33197 );
    nor g14207 ( n11322 , n18298 , n13623 );
    nor g14208 ( n29458 , n41715 , n7349 );
    or g14209 ( n4973 , n37503 , n4381 );
    and g14210 ( n16675 , n3880 , n2970 );
    not g14211 ( n16650 , n17347 );
    xnor g14212 ( n42475 , n41515 , n18777 );
    and g14213 ( n33725 , n725 , n18045 );
    or g14214 ( n25857 , n21310 , n37687 );
    and g14215 ( n1610 , n14951 , n18545 );
    or g14216 ( n4719 , n14787 , n33548 );
    not g14217 ( n42465 , n7820 );
    nor g14218 ( n24379 , n25508 , n31457 );
    and g14219 ( n42746 , n4254 , n9296 );
    and g14220 ( n8299 , n41109 , n38516 );
    nor g14221 ( n23235 , n35259 , n29017 );
    not g14222 ( n42383 , n23393 );
    or g14223 ( n42611 , n40754 , n27683 );
    xnor g14224 ( n41713 , n36998 , n36504 );
    or g14225 ( n22209 , n6503 , n33657 );
    or g14226 ( n4787 , n37093 , n13723 );
    or g14227 ( n21119 , n16439 , n23916 );
    or g14228 ( n19271 , n6247 , n3888 );
    and g14229 ( n20265 , n37326 , n3844 );
    and g14230 ( n20659 , n22357 , n41445 );
    and g14231 ( n35423 , n7676 , n18919 );
    or g14232 ( n1036 , n25600 , n29548 );
    nor g14233 ( n26031 , n7197 , n5852 );
    or g14234 ( n26472 , n16422 , n15996 );
    and g14235 ( n21650 , n42598 , n2627 );
    or g14236 ( n40873 , n2484 , n36570 );
    or g14237 ( n28342 , n25291 , n1220 );
    or g14238 ( n4279 , n363 , n26139 );
    not g14239 ( n2628 , n30797 );
    not g14240 ( n19803 , n16566 );
    nor g14241 ( n1062 , n40090 , n2280 );
    or g14242 ( n13550 , n5350 , n31221 );
    or g14243 ( n98 , n34337 , n1210 );
    not g14244 ( n11375 , n23567 );
    nor g14245 ( n25708 , n14707 , n26531 );
    not g14246 ( n28225 , n28150 );
    or g14247 ( n6407 , n16968 , n15808 );
    nor g14248 ( n4865 , n15176 , n820 );
    and g14249 ( n20354 , n5184 , n11807 );
    and g14250 ( n12925 , n38719 , n41821 );
    nor g14251 ( n4589 , n20357 , n21890 );
    or g14252 ( n37101 , n15096 , n5896 );
    or g14253 ( n31718 , n41871 , n34278 );
    or g14254 ( n15915 , n13398 , n21694 );
    or g14255 ( n5976 , n17034 , n6173 );
    nor g14256 ( n21821 , n39858 , n22536 );
    or g14257 ( n7007 , n17307 , n26714 );
    or g14258 ( n30813 , n31924 , n14601 );
    and g14259 ( n30493 , n35545 , n15898 );
    nor g14260 ( n14539 , n23502 , n34241 );
    or g14261 ( n30258 , n32221 , n9456 );
    not g14262 ( n20165 , n30634 );
    xnor g14263 ( n12405 , n5144 , n31809 );
    or g14264 ( n39683 , n42699 , n18779 );
    or g14265 ( n37993 , n19969 , n41061 );
    and g14266 ( n29548 , n28212 , n17474 );
    or g14267 ( n29699 , n19034 , n1416 );
    and g14268 ( n11294 , n37127 , n35484 );
    or g14269 ( n337 , n19737 , n21893 );
    or g14270 ( n33576 , n516 , n38676 );
    or g14271 ( n15361 , n36104 , n15960 );
    not g14272 ( n15272 , n33397 );
    nor g14273 ( n5637 , n26377 , n13629 );
    or g14274 ( n39114 , n18323 , n12740 );
    or g14275 ( n8 , n5605 , n20604 );
    and g14276 ( n17499 , n24889 , n24850 );
    and g14277 ( n7061 , n42287 , n6738 );
    or g14278 ( n15057 , n41974 , n1208 );
    or g14279 ( n2860 , n19084 , n3595 );
    xnor g14280 ( n9191 , n15488 , n25791 );
    not g14281 ( n37114 , n26297 );
    xnor g14282 ( n22383 , n5144 , n37056 );
    and g14283 ( n15098 , n38608 , n22801 );
    or g14284 ( n10715 , n34189 , n25986 );
    and g14285 ( n2924 , n42019 , n5118 );
    or g14286 ( n39514 , n10060 , n33475 );
    nor g14287 ( n24613 , n29579 , n4815 );
    nor g14288 ( n25204 , n15602 , n22713 );
    xnor g14289 ( n40105 , n22773 , n5852 );
    xnor g14290 ( n40150 , n7922 , n34011 );
    and g14291 ( n23092 , n8098 , n16851 );
    or g14292 ( n14162 , n23586 , n14676 );
    or g14293 ( n11616 , n3447 , n41071 );
    xnor g14294 ( n20208 , n29740 , n26391 );
    and g14295 ( n39904 , n5137 , n27097 );
    or g14296 ( n8336 , n42558 , n20687 );
    and g14297 ( n35258 , n8614 , n15229 );
    xnor g14298 ( n1104 , n19230 , n41960 );
    or g14299 ( n12861 , n19166 , n6590 );
    or g14300 ( n38265 , n40995 , n10998 );
    nor g14301 ( n34705 , n41558 , n28661 );
    or g14302 ( n22195 , n27670 , n36542 );
    not g14303 ( n33211 , n2068 );
    xnor g14304 ( n28110 , n42715 , n11539 );
    xnor g14305 ( n39344 , n28073 , n10573 );
    xnor g14306 ( n6298 , n11436 , n13000 );
    or g14307 ( n19961 , n21096 , n389 );
    or g14308 ( n37034 , n3218 , n11924 );
    and g14309 ( n41739 , n24472 , n8080 );
    not g14310 ( n26142 , n31043 );
    and g14311 ( n471 , n31872 , n29293 );
    or g14312 ( n10520 , n42361 , n8052 );
    xnor g14313 ( n34263 , n11436 , n11036 );
    nor g14314 ( n22969 , n24745 , n33873 );
    not g14315 ( n14394 , n35766 );
    and g14316 ( n4946 , n11064 , n40107 );
    nor g14317 ( n449 , n19221 , n13750 );
    xnor g14318 ( n19199 , n4341 , n6592 );
    and g14319 ( n17569 , n39641 , n511 );
    and g14320 ( n34828 , n41746 , n3577 );
    or g14321 ( n39488 , n8381 , n2710 );
    not g14322 ( n38197 , n12069 );
    not g14323 ( n1120 , n3393 );
    or g14324 ( n36113 , n17573 , n12486 );
    or g14325 ( n24534 , n22091 , n12374 );
    and g14326 ( n23259 , n19604 , n33916 );
    and g14327 ( n31166 , n28368 , n504 );
    xnor g14328 ( n15161 , n6969 , n12234 );
    or g14329 ( n5730 , n26253 , n40942 );
    xnor g14330 ( n20087 , n21665 , n8494 );
    or g14331 ( n10683 , n5951 , n20646 );
    not g14332 ( n5355 , n35470 );
    and g14333 ( n646 , n41059 , n4793 );
    or g14334 ( n36475 , n7020 , n6553 );
    xnor g14335 ( n11914 , n5370 , n28868 );
    and g14336 ( n28079 , n36935 , n8883 );
    and g14337 ( n38678 , n18194 , n10543 );
    or g14338 ( n34152 , n26627 , n15098 );
    nor g14339 ( n39986 , n179 , n2480 );
    not g14340 ( n10939 , n18247 );
    not g14341 ( n41306 , n32124 );
    and g14342 ( n13235 , n32418 , n16406 );
    and g14343 ( n37183 , n8251 , n11654 );
    nor g14344 ( n38956 , n172 , n8758 );
    xnor g14345 ( n33405 , n42064 , n18042 );
    not g14346 ( n27884 , n22160 );
    nor g14347 ( n29824 , n20557 , n13906 );
    or g14348 ( n30006 , n24503 , n18265 );
    nor g14349 ( n4243 , n3360 , n15745 );
    or g14350 ( n18869 , n15116 , n19432 );
    xnor g14351 ( n16921 , n40852 , n22914 );
    or g14352 ( n14391 , n13657 , n20514 );
    or g14353 ( n10474 , n42565 , n29846 );
    not g14354 ( n26974 , n34446 );
    and g14355 ( n21564 , n40803 , n3279 );
    nor g14356 ( n286 , n14687 , n16430 );
    or g14357 ( n4989 , n2153 , n6024 );
    not g14358 ( n38339 , n39989 );
    and g14359 ( n31165 , n16384 , n26267 );
    and g14360 ( n42529 , n37354 , n31695 );
    xnor g14361 ( n30945 , n24259 , n34292 );
    nor g14362 ( n23216 , n17120 , n22683 );
    and g14363 ( n9767 , n10201 , n38951 );
    or g14364 ( n40949 , n15287 , n19366 );
    or g14365 ( n19228 , n40750 , n37397 );
    or g14366 ( n34214 , n38733 , n571 );
    and g14367 ( n24722 , n17236 , n3841 );
    or g14368 ( n4616 , n1326 , n17145 );
    nor g14369 ( n12930 , n39705 , n6418 );
    or g14370 ( n7348 , n34696 , n31426 );
    nor g14371 ( n5802 , n27219 , n15782 );
    not g14372 ( n15989 , n36611 );
    and g14373 ( n13244 , n4544 , n16592 );
    or g14374 ( n41222 , n31114 , n36619 );
    or g14375 ( n9510 , n31605 , n12153 );
    or g14376 ( n9921 , n38374 , n35713 );
    nor g14377 ( n34873 , n26535 , n2536 );
    or g14378 ( n8546 , n37970 , n21019 );
    nor g14379 ( n31758 , n29757 , n16430 );
    nor g14380 ( n20013 , n12033 , n42599 );
    nor g14381 ( n7157 , n42676 , n17459 );
    or g14382 ( n28776 , n11394 , n8087 );
    and g14383 ( n32884 , n12052 , n37068 );
    or g14384 ( n9181 , n41598 , n20900 );
    nor g14385 ( n6596 , n14654 , n24337 );
    and g14386 ( n36976 , n20878 , n13307 );
    and g14387 ( n20171 , n34803 , n40243 );
    xnor g14388 ( n23663 , n34352 , n41592 );
    or g14389 ( n29212 , n15040 , n19863 );
    or g14390 ( n2090 , n8490 , n12853 );
    and g14391 ( n20041 , n12629 , n2257 );
    and g14392 ( n12926 , n33890 , n6605 );
    or g14393 ( n41687 , n24228 , n3020 );
    and g14394 ( n1518 , n37283 , n2248 );
    xnor g14395 ( n9316 , n37176 , n35260 );
    and g14396 ( n10737 , n2578 , n15376 );
    or g14397 ( n14372 , n8347 , n25818 );
    or g14398 ( n24314 , n25573 , n21618 );
    and g14399 ( n969 , n28132 , n30883 );
    not g14400 ( n24948 , n33441 );
    and g14401 ( n20184 , n8489 , n21274 );
    or g14402 ( n7104 , n29872 , n6270 );
    nor g14403 ( n41237 , n32868 , n33493 );
    xnor g14404 ( n2886 , n32297 , n8418 );
    or g14405 ( n24922 , n28733 , n39993 );
    or g14406 ( n8964 , n17352 , n21096 );
    nor g14407 ( n6633 , n1186 , n13347 );
    nor g14408 ( n30868 , n16866 , n7710 );
    and g14409 ( n12853 , n30059 , n4586 );
    or g14410 ( n40918 , n31001 , n23718 );
    or g14411 ( n28327 , n20233 , n13284 );
    not g14412 ( n25055 , n20537 );
    xnor g14413 ( n39743 , n21973 , n23607 );
    and g14414 ( n39256 , n6844 , n26532 );
    or g14415 ( n13229 , n28883 , n7202 );
    or g14416 ( n25080 , n29455 , n36107 );
    or g14417 ( n22113 , n163 , n23071 );
    xnor g14418 ( n38136 , n23938 , n15408 );
    not g14419 ( n37654 , n6821 );
    not g14420 ( n19391 , n39669 );
    or g14421 ( n13427 , n20092 , n35667 );
    not g14422 ( n29560 , n24622 );
    or g14423 ( n23662 , n24448 , n8780 );
    or g14424 ( n27415 , n17663 , n17902 );
    xnor g14425 ( n36241 , n7791 , n5971 );
    or g14426 ( n6090 , n30491 , n39557 );
    nor g14427 ( n26140 , n17120 , n3116 );
    nor g14428 ( n5281 , n4492 , n5025 );
    and g14429 ( n29122 , n975 , n8238 );
    or g14430 ( n23626 , n4839 , n10692 );
    and g14431 ( n38713 , n13087 , n29244 );
    or g14432 ( n11198 , n6482 , n31763 );
    and g14433 ( n7921 , n34508 , n42187 );
    and g14434 ( n23280 , n18380 , n41422 );
    and g14435 ( n32318 , n34737 , n11819 );
    nor g14436 ( n11369 , n33053 , n33241 );
    or g14437 ( n21079 , n5324 , n21820 );
    and g14438 ( n34908 , n6127 , n42717 );
    nor g14439 ( n12993 , n5302 , n11324 );
    nor g14440 ( n38192 , n32542 , n10402 );
    nor g14441 ( n6622 , n39630 , n9615 );
    xnor g14442 ( n5639 , n21765 , n6913 );
    or g14443 ( n10981 , n33296 , n40605 );
    not g14444 ( n3423 , n36049 );
    nor g14445 ( n36458 , n5649 , n37081 );
    or g14446 ( n5477 , n14407 , n6486 );
    and g14447 ( n42188 , n39566 , n9096 );
    xnor g14448 ( n38677 , n16720 , n19939 );
    not g14449 ( n5097 , n22097 );
    or g14450 ( n21809 , n2880 , n27953 );
    nor g14451 ( n31465 , n7059 , n25879 );
    and g14452 ( n20691 , n37834 , n21809 );
    xnor g14453 ( n7439 , n25299 , n6408 );
    or g14454 ( n15816 , n3322 , n13316 );
    or g14455 ( n7052 , n1463 , n7663 );
    and g14456 ( n15661 , n35991 , n42629 );
    or g14457 ( n18708 , n25924 , n31595 );
    or g14458 ( n11292 , n22293 , n34079 );
    xnor g14459 ( n25428 , n34945 , n16293 );
    and g14460 ( n37759 , n33147 , n12583 );
    or g14461 ( n36834 , n1110 , n11381 );
    and g14462 ( n35636 , n23160 , n31852 );
    xnor g14463 ( n17206 , n34352 , n13524 );
    not g14464 ( n26426 , n585 );
    or g14465 ( n42234 , n1013 , n9969 );
    and g14466 ( n6718 , n26813 , n21750 );
    or g14467 ( n23264 , n5978 , n8984 );
    or g14468 ( n2398 , n23973 , n25451 );
    or g14469 ( n27055 , n16564 , n42504 );
    or g14470 ( n42868 , n16897 , n14949 );
    or g14471 ( n33761 , n1783 , n19091 );
    nor g14472 ( n2197 , n9272 , n21547 );
    or g14473 ( n39081 , n18543 , n39539 );
    not g14474 ( n14647 , n16099 );
    or g14475 ( n19812 , n20932 , n2774 );
    and g14476 ( n24263 , n35316 , n8043 );
    or g14477 ( n13527 , n40465 , n37679 );
    or g14478 ( n29408 , n18564 , n24262 );
    nor g14479 ( n13920 , n11120 , n29986 );
    xnor g14480 ( n260 , n34226 , n14761 );
    nor g14481 ( n9969 , n20483 , n28084 );
    nor g14482 ( n17694 , n8494 , n26947 );
    or g14483 ( n25889 , n18557 , n41340 );
    not g14484 ( n31279 , n14362 );
    or g14485 ( n42560 , n33588 , n28678 );
    or g14486 ( n13047 , n10284 , n41252 );
    xnor g14487 ( n17459 , n2903 , n26594 );
    nor g14488 ( n18687 , n32793 , n4790 );
    not g14489 ( n19636 , n35132 );
    or g14490 ( n5385 , n8130 , n17109 );
    nor g14491 ( n29186 , n26011 , n42199 );
    xnor g14492 ( n33996 , n8857 , n35010 );
    and g14493 ( n29909 , n34879 , n14247 );
    or g14494 ( n226 , n14642 , n35787 );
    and g14495 ( n39460 , n15741 , n8760 );
    and g14496 ( n3261 , n13884 , n15072 );
    nor g14497 ( n37755 , n16598 , n21900 );
    and g14498 ( n15012 , n22902 , n1022 );
    and g14499 ( n37885 , n95 , n41697 );
    and g14500 ( n14262 , n20012 , n5853 );
    xnor g14501 ( n38901 , n71 , n38544 );
    and g14502 ( n30581 , n41933 , n23120 );
    xnor g14503 ( n1114 , n38607 , n42571 );
    and g14504 ( n9955 , n11063 , n489 );
    or g14505 ( n22214 , n27977 , n14553 );
    or g14506 ( n7546 , n24722 , n11291 );
    xnor g14507 ( n30361 , n11691 , n41579 );
    and g14508 ( n11084 , n21385 , n26804 );
    xnor g14509 ( n35279 , n784 , n21031 );
    or g14510 ( n1313 , n16714 , n34140 );
    and g14511 ( n7349 , n8272 , n2446 );
    or g14512 ( n8580 , n30243 , n33858 );
    or g14513 ( n22906 , n7446 , n25136 );
    xnor g14514 ( n27516 , n34731 , n29023 );
    and g14515 ( n6643 , n23534 , n20240 );
    and g14516 ( n33609 , n37133 , n28981 );
    or g14517 ( n26236 , n13314 , n946 );
    xnor g14518 ( n2073 , n37146 , n19563 );
    nor g14519 ( n22883 , n25875 , n1653 );
    and g14520 ( n34555 , n6163 , n5285 );
    xnor g14521 ( n148 , n15842 , n29140 );
    or g14522 ( n34142 , n10681 , n28316 );
    and g14523 ( n23637 , n26952 , n29205 );
    xnor g14524 ( n3684 , n25473 , n41367 );
    and g14525 ( n42631 , n14961 , n5510 );
    xnor g14526 ( n9278 , n27684 , n23754 );
    and g14527 ( n27251 , n20423 , n29586 );
    nor g14528 ( n41964 , n28673 , n12914 );
    nor g14529 ( n32317 , n688 , n30821 );
    not g14530 ( n2117 , n40974 );
    or g14531 ( n21984 , n38179 , n3170 );
    or g14532 ( n27659 , n28634 , n34423 );
    xnor g14533 ( n9742 , n28443 , n13325 );
    or g14534 ( n5566 , n6432 , n42653 );
    or g14535 ( n9960 , n19260 , n7148 );
    and g14536 ( n42811 , n9273 , n32045 );
    not g14537 ( n2841 , n32499 );
    and g14538 ( n1396 , n29189 , n4817 );
    and g14539 ( n20169 , n26535 , n2536 );
    or g14540 ( n41960 , n14128 , n4786 );
    and g14541 ( n30118 , n11401 , n33650 );
    nor g14542 ( n23818 , n3893 , n3587 );
    or g14543 ( n42689 , n39804 , n2891 );
    nor g14544 ( n248 , n9041 , n28478 );
    and g14545 ( n30782 , n15076 , n32817 );
    and g14546 ( n4895 , n32015 , n28552 );
    nor g14547 ( n28408 , n5896 , n19691 );
    or g14548 ( n25226 , n36797 , n37299 );
    or g14549 ( n23524 , n25094 , n19616 );
    or g14550 ( n33893 , n11327 , n40059 );
    or g14551 ( n30288 , n28056 , n16466 );
    xnor g14552 ( n25665 , n16197 , n5964 );
    and g14553 ( n39134 , n24731 , n41402 );
    or g14554 ( n16312 , n34787 , n8341 );
    not g14555 ( n37357 , n26871 );
    and g14556 ( n35801 , n1710 , n17251 );
    xnor g14557 ( n15903 , n21012 , n1235 );
    xnor g14558 ( n36965 , n19448 , n32795 );
    xnor g14559 ( n6776 , n842 , n34984 );
    nor g14560 ( n21806 , n42884 , n11555 );
    not g14561 ( n14749 , n8734 );
    and g14562 ( n38088 , n37609 , n10627 );
    and g14563 ( n17457 , n42484 , n11182 );
    nor g14564 ( n10895 , n6929 , n30963 );
    not g14565 ( n41773 , n33927 );
    and g14566 ( n42877 , n25706 , n22282 );
    or g14567 ( n16569 , n1507 , n5799 );
    or g14568 ( n2058 , n24626 , n26688 );
    and g14569 ( n41243 , n33636 , n36330 );
    or g14570 ( n17951 , n26670 , n12751 );
    or g14571 ( n21104 , n3794 , n15818 );
    or g14572 ( n36770 , n1665 , n25528 );
    xnor g14573 ( n25772 , n11436 , n37510 );
    or g14574 ( n3784 , n35913 , n24583 );
    or g14575 ( n11185 , n14048 , n20063 );
    or g14576 ( n24752 , n6578 , n36477 );
    not g14577 ( n34618 , n937 );
    and g14578 ( n8374 , n26222 , n36984 );
    and g14579 ( n18026 , n17387 , n9500 );
    and g14580 ( n27275 , n27720 , n41033 );
    not g14581 ( n10559 , n294 );
    not g14582 ( n635 , n10089 );
    and g14583 ( n19632 , n18960 , n30124 );
    and g14584 ( n9471 , n36541 , n7991 );
    and g14585 ( n5833 , n21227 , n41913 );
    and g14586 ( n12435 , n30211 , n266 );
    not g14587 ( n1598 , n32007 );
    not g14588 ( n12383 , n12742 );
    and g14589 ( n9867 , n14428 , n625 );
    not g14590 ( n28872 , n27086 );
    or g14591 ( n39854 , n3172 , n18863 );
    nor g14592 ( n2255 , n26172 , n28900 );
    and g14593 ( n10172 , n17886 , n2973 );
    or g14594 ( n8958 , n6807 , n31321 );
    xnor g14595 ( n34264 , n25143 , n37238 );
    and g14596 ( n14526 , n35796 , n31719 );
    and g14597 ( n14043 , n1174 , n36385 );
    or g14598 ( n78 , n34565 , n17222 );
    or g14599 ( n40250 , n38546 , n17883 );
    or g14600 ( n35909 , n40110 , n36690 );
    or g14601 ( n11536 , n12867 , n10410 );
    or g14602 ( n42593 , n38525 , n16985 );
    or g14603 ( n11839 , n16155 , n17344 );
    and g14604 ( n28487 , n20026 , n42167 );
    xnor g14605 ( n39529 , n23120 , n41933 );
    nor g14606 ( n34545 , n36950 , n11538 );
    and g14607 ( n17258 , n25056 , n20747 );
    or g14608 ( n9361 , n39256 , n20383 );
    not g14609 ( n27764 , n41117 );
    and g14610 ( n3758 , n24586 , n36049 );
    and g14611 ( n16047 , n20875 , n31041 );
    or g14612 ( n26543 , n18474 , n41304 );
    or g14613 ( n4634 , n15384 , n10222 );
    or g14614 ( n15352 , n15470 , n16613 );
    nor g14615 ( n463 , n37639 , n10141 );
    not g14616 ( n1877 , n40696 );
    or g14617 ( n21299 , n20412 , n41156 );
    or g14618 ( n24924 , n35269 , n11593 );
    xnor g14619 ( n39815 , n16411 , n22267 );
    nor g14620 ( n23568 , n26565 , n1176 );
    or g14621 ( n9797 , n3307 , n25528 );
    not g14622 ( n11705 , n19721 );
    nor g14623 ( n26112 , n2637 , n18139 );
    or g14624 ( n17330 , n20271 , n25335 );
    and g14625 ( n39761 , n39447 , n10238 );
    or g14626 ( n10809 , n37031 , n30884 );
    nor g14627 ( n29771 , n15136 , n26814 );
    nor g14628 ( n13457 , n11360 , n6123 );
    or g14629 ( n10040 , n34359 , n17404 );
    or g14630 ( n41794 , n39055 , n2034 );
    or g14631 ( n20829 , n40978 , n26546 );
    not g14632 ( n16695 , n2880 );
    or g14633 ( n24071 , n14996 , n33463 );
    or g14634 ( n24099 , n16910 , n1191 );
    not g14635 ( n11353 , n9682 );
    xnor g14636 ( n19453 , n25582 , n39550 );
    or g14637 ( n15334 , n1449 , n11054 );
    nor g14638 ( n6183 , n39114 , n25450 );
    and g14639 ( n4630 , n32413 , n14335 );
    not g14640 ( n37494 , n22954 );
    and g14641 ( n30024 , n19898 , n6787 );
    or g14642 ( n36268 , n36998 , n42877 );
    xnor g14643 ( n39221 , n12120 , n6980 );
    and g14644 ( n31170 , n10739 , n1030 );
    or g14645 ( n5937 , n19056 , n40823 );
    or g14646 ( n22117 , n14112 , n55 );
    and g14647 ( n33657 , n26397 , n27508 );
    or g14648 ( n28043 , n15030 , n20103 );
    not g14649 ( n11610 , n27406 );
    or g14650 ( n42838 , n4790 , n39126 );
    not g14651 ( n28612 , n35759 );
    and g14652 ( n25216 , n26534 , n4198 );
    or g14653 ( n36986 , n5386 , n12011 );
    not g14654 ( n24856 , n40772 );
    and g14655 ( n40760 , n27044 , n11193 );
    xnor g14656 ( n7346 , n4188 , n11975 );
    or g14657 ( n18283 , n26122 , n29635 );
    or g14658 ( n4110 , n40210 , n12288 );
    and g14659 ( n34688 , n31477 , n1001 );
    or g14660 ( n31761 , n18233 , n28023 );
    or g14661 ( n26583 , n17904 , n40479 );
    or g14662 ( n16583 , n39700 , n27330 );
    or g14663 ( n41192 , n30283 , n4535 );
    and g14664 ( n39093 , n22809 , n4406 );
    not g14665 ( n35634 , n42738 );
    xnor g14666 ( n35449 , n35217 , n33546 );
    nor g14667 ( n36373 , n23549 , n11912 );
    nor g14668 ( n28234 , n23311 , n32988 );
    and g14669 ( n3210 , n19760 , n33829 );
    and g14670 ( n18438 , n40172 , n11611 );
    and g14671 ( n28421 , n18704 , n41692 );
    nor g14672 ( n1270 , n11147 , n35577 );
    or g14673 ( n8308 , n16147 , n16434 );
    or g14674 ( n20670 , n5327 , n31710 );
    nor g14675 ( n33382 , n9287 , n11406 );
    or g14676 ( n31178 , n40253 , n30114 );
    and g14677 ( n32133 , n19165 , n27405 );
    xnor g14678 ( n198 , n1768 , n21243 );
    or g14679 ( n4420 , n23502 , n35260 );
    xnor g14680 ( n35215 , n26579 , n16684 );
    and g14681 ( n35297 , n8859 , n35685 );
    not g14682 ( n20854 , n31393 );
    not g14683 ( n17238 , n1037 );
    and g14684 ( n3689 , n26881 , n3730 );
    xnor g14685 ( n39598 , n42725 , n23009 );
    nor g14686 ( n8491 , n21309 , n11539 );
    or g14687 ( n17648 , n28533 , n13346 );
    and g14688 ( n33115 , n8054 , n12755 );
    or g14689 ( n27662 , n11248 , n6391 );
    or g14690 ( n22565 , n31997 , n15942 );
    not g14691 ( n32175 , n7958 );
    or g14692 ( n1249 , n12880 , n2479 );
    not g14693 ( n10985 , n40284 );
    and g14694 ( n6595 , n21053 , n4071 );
    and g14695 ( n16719 , n29716 , n4943 );
    or g14696 ( n934 , n38921 , n10433 );
    or g14697 ( n21226 , n28745 , n22805 );
    or g14698 ( n22327 , n24843 , n31688 );
    xnor g14699 ( n33941 , n26168 , n33977 );
    not g14700 ( n26313 , n40447 );
    or g14701 ( n21005 , n16782 , n27220 );
    or g14702 ( n38425 , n39397 , n3891 );
    not g14703 ( n16797 , n40078 );
    xnor g14704 ( n6342 , n29917 , n10671 );
    or g14705 ( n40268 , n32104 , n3678 );
    or g14706 ( n41403 , n26951 , n9617 );
    or g14707 ( n37773 , n38056 , n25451 );
    not g14708 ( n19612 , n31892 );
    or g14709 ( n37892 , n37123 , n8148 );
    not g14710 ( n39105 , n28792 );
    and g14711 ( n37767 , n39740 , n16310 );
    nor g14712 ( n15987 , n6901 , n41078 );
    or g14713 ( n35214 , n22844 , n5800 );
    and g14714 ( n21312 , n36131 , n31509 );
    not g14715 ( n5842 , n4208 );
    not g14716 ( n12524 , n28632 );
    or g14717 ( n11081 , n9279 , n37545 );
    not g14718 ( n28861 , n41864 );
    nor g14719 ( n7159 , n20469 , n27955 );
    xnor g14720 ( n25447 , n21291 , n15177 );
    nor g14721 ( n10908 , n9552 , n38575 );
    or g14722 ( n2163 , n26346 , n20287 );
    and g14723 ( n20211 , n18678 , n3185 );
    or g14724 ( n218 , n25456 , n180 );
    or g14725 ( n5486 , n18966 , n21852 );
    and g14726 ( n42813 , n30949 , n13377 );
    nor g14727 ( n13694 , n36117 , n37972 );
    and g14728 ( n6666 , n13508 , n18286 );
    xnor g14729 ( n3368 , n35563 , n1914 );
    and g14730 ( n31071 , n37004 , n31369 );
    nor g14731 ( n35037 , n22484 , n1414 );
    xnor g14732 ( n25400 , n35727 , n13147 );
    and g14733 ( n4530 , n16228 , n4692 );
    or g14734 ( n3165 , n9757 , n12198 );
    or g14735 ( n29926 , n15025 , n26167 );
    or g14736 ( n38099 , n33581 , n776 );
    and g14737 ( n1231 , n16619 , n9221 );
    nor g14738 ( n6598 , n8933 , n35126 );
    or g14739 ( n20344 , n16598 , n21583 );
    or g14740 ( n5491 , n11976 , n2948 );
    nor g14741 ( n42637 , n12779 , n12673 );
    and g14742 ( n38389 , n38587 , n5792 );
    nor g14743 ( n24839 , n37057 , n10457 );
    or g14744 ( n6121 , n40752 , n14806 );
    not g14745 ( n16332 , n6768 );
    not g14746 ( n3309 , n42624 );
    and g14747 ( n17862 , n17882 , n30267 );
    and g14748 ( n29890 , n14187 , n6439 );
    not g14749 ( n14941 , n9062 );
    and g14750 ( n30185 , n29582 , n24777 );
    and g14751 ( n2912 , n20538 , n37204 );
    and g14752 ( n38107 , n14148 , n6747 );
    or g14753 ( n4049 , n18169 , n6740 );
    or g14754 ( n22223 , n2917 , n36848 );
    or g14755 ( n25114 , n2710 , n30521 );
    and g14756 ( n34567 , n29894 , n33064 );
    or g14757 ( n37775 , n1395 , n34991 );
    or g14758 ( n13253 , n16817 , n37733 );
    nor g14759 ( n8571 , n34356 , n32016 );
    not g14760 ( n9432 , n34277 );
    or g14761 ( n8425 , n10197 , n28191 );
    or g14762 ( n1235 , n39186 , n7496 );
    or g14763 ( n4582 , n20092 , n9438 );
    xnor g14764 ( n11903 , n35876 , n26025 );
    and g14765 ( n27812 , n26212 , n19491 );
    not g14766 ( n346 , n10337 );
    not g14767 ( n13539 , n30479 );
    or g14768 ( n26878 , n8592 , n40587 );
    or g14769 ( n15417 , n20629 , n19540 );
    nor g14770 ( n41110 , n13029 , n1966 );
    not g14771 ( n28150 , n34363 );
    and g14772 ( n39596 , n12691 , n1482 );
    or g14773 ( n27246 , n9612 , n30450 );
    not g14774 ( n35512 , n30894 );
    nor g14775 ( n36945 , n2372 , n9518 );
    and g14776 ( n19971 , n5773 , n1652 );
    not g14777 ( n25170 , n1267 );
    not g14778 ( n42072 , n28563 );
    nor g14779 ( n25753 , n41065 , n15791 );
    and g14780 ( n11389 , n32765 , n24009 );
    or g14781 ( n14891 , n21273 , n16659 );
    or g14782 ( n3252 , n29545 , n36537 );
    and g14783 ( n21825 , n21922 , n10151 );
    or g14784 ( n6829 , n7375 , n39884 );
    and g14785 ( n12354 , n21716 , n23616 );
    nor g14786 ( n19917 , n6671 , n30199 );
    or g14787 ( n29424 , n32458 , n32353 );
    xnor g14788 ( n24209 , n11436 , n14634 );
    nor g14789 ( n15632 , n14471 , n364 );
    nor g14790 ( n3298 , n4430 , n35424 );
    or g14791 ( n8106 , n10559 , n37435 );
    and g14792 ( n3680 , n5781 , n16942 );
    or g14793 ( n26007 , n8068 , n18014 );
    xnor g14794 ( n34163 , n20629 , n14707 );
    or g14795 ( n1966 , n27523 , n6016 );
    nor g14796 ( n32974 , n16011 , n2378 );
    or g14797 ( n2887 , n33556 , n19 );
    or g14798 ( n25404 , n3320 , n31232 );
    or g14799 ( n40783 , n26262 , n7474 );
    nor g14800 ( n1904 , n40755 , n39246 );
    and g14801 ( n15152 , n7183 , n16062 );
    xnor g14802 ( n22443 , n37394 , n35826 );
    and g14803 ( n19214 , n35022 , n38641 );
    not g14804 ( n10839 , n28024 );
    or g14805 ( n14247 , n8078 , n8658 );
    or g14806 ( n22684 , n10822 , n40746 );
    and g14807 ( n15511 , n40051 , n9425 );
    nor g14808 ( n118 , n20708 , n33895 );
    and g14809 ( n33427 , n15747 , n41308 );
    or g14810 ( n5224 , n25169 , n20378 );
    not g14811 ( n39511 , n22780 );
    or g14812 ( n13522 , n8062 , n42385 );
    and g14813 ( n14728 , n35041 , n7481 );
    or g14814 ( n4916 , n4114 , n37819 );
    not g14815 ( n2679 , n21193 );
    and g14816 ( n35949 , n24492 , n33194 );
    or g14817 ( n13775 , n37647 , n26986 );
    and g14818 ( n22288 , n26979 , n1957 );
    nor g14819 ( n22743 , n27137 , n35127 );
    or g14820 ( n28902 , n1581 , n7097 );
    xnor g14821 ( n13611 , n23304 , n22249 );
    not g14822 ( n32726 , n17350 );
    or g14823 ( n41128 , n25078 , n18508 );
    not g14824 ( n28313 , n6260 );
    not g14825 ( n1464 , n39200 );
    not g14826 ( n31541 , n19861 );
    not g14827 ( n19084 , n40078 );
    or g14828 ( n32595 , n33706 , n36842 );
    or g14829 ( n25717 , n28069 , n19734 );
    nor g14830 ( n24743 , n28603 , n1912 );
    nor g14831 ( n24403 , n25060 , n2870 );
    or g14832 ( n5106 , n26147 , n38706 );
    or g14833 ( n15419 , n25721 , n2865 );
    or g14834 ( n11611 , n3546 , n10792 );
    or g14835 ( n40684 , n37379 , n7398 );
    or g14836 ( n8278 , n33774 , n19143 );
    nor g14837 ( n2256 , n32120 , n13233 );
    and g14838 ( n6960 , n23594 , n10335 );
    not g14839 ( n38293 , n13668 );
    not g14840 ( n12316 , n35463 );
    not g14841 ( n14215 , n3790 );
    not g14842 ( n23800 , n36800 );
    or g14843 ( n1657 , n39523 , n21006 );
    and g14844 ( n37672 , n41075 , n42791 );
    xnor g14845 ( n41177 , n20958 , n23141 );
    or g14846 ( n33362 , n11658 , n29024 );
    or g14847 ( n32921 , n18132 , n30140 );
    not g14848 ( n2296 , n5661 );
    or g14849 ( n3050 , n4343 , n13034 );
    or g14850 ( n15117 , n25724 , n42470 );
    not g14851 ( n32978 , n26261 );
    nor g14852 ( n16292 , n5111 , n18290 );
    not g14853 ( n6699 , n30083 );
    and g14854 ( n36328 , n16200 , n32428 );
    or g14855 ( n25925 , n8004 , n11815 );
    and g14856 ( n33032 , n41926 , n27255 );
    or g14857 ( n12944 , n12616 , n30896 );
    and g14858 ( n5551 , n31972 , n22393 );
    or g14859 ( n9850 , n27140 , n8141 );
    not g14860 ( n36526 , n4149 );
    or g14861 ( n8325 , n42115 , n30909 );
    and g14862 ( n21535 , n38488 , n38229 );
    not g14863 ( n16688 , n23186 );
    xnor g14864 ( n13960 , n32018 , n4140 );
    or g14865 ( n1984 , n34860 , n27151 );
    or g14866 ( n16943 , n20978 , n17434 );
    and g14867 ( n23949 , n41837 , n27474 );
    and g14868 ( n6249 , n15168 , n29517 );
    and g14869 ( n17466 , n21171 , n34309 );
    xnor g14870 ( n11716 , n4470 , n39761 );
    and g14871 ( n33542 , n31197 , n34426 );
    and g14872 ( n24471 , n23439 , n9728 );
    not g14873 ( n1788 , n28850 );
    xnor g14874 ( n12646 , n24527 , n24738 );
    not g14875 ( n201 , n30451 );
    xnor g14876 ( n34924 , n40491 , n1698 );
    or g14877 ( n115 , n6929 , n36227 );
    and g14878 ( n8893 , n3756 , n18340 );
    xnor g14879 ( n10577 , n7922 , n40071 );
    nor g14880 ( n61 , n39718 , n19094 );
    or g14881 ( n37818 , n32587 , n28028 );
    not g14882 ( n23132 , n13721 );
    or g14883 ( n10026 , n1971 , n29571 );
    xnor g14884 ( n16624 , n19752 , n17099 );
    not g14885 ( n18532 , n33920 );
    not g14886 ( n2444 , n1679 );
    and g14887 ( n41860 , n30641 , n8424 );
    xnor g14888 ( n7306 , n4334 , n22661 );
    and g14889 ( n16508 , n39359 , n41790 );
    not g14890 ( n7125 , n10819 );
    or g14891 ( n28266 , n25958 , n38637 );
    xnor g14892 ( n6650 , n34810 , n4594 );
    or g14893 ( n11587 , n33580 , n22455 );
    not g14894 ( n36676 , n22318 );
    xnor g14895 ( n41607 , n542 , n22502 );
    xnor g14896 ( n35698 , n40 , n24299 );
    and g14897 ( n5284 , n7356 , n40081 );
    xnor g14898 ( n28916 , n3455 , n30051 );
    and g14899 ( n13762 , n26030 , n24390 );
    or g14900 ( n25051 , n38633 , n10926 );
    xnor g14901 ( n18054 , n19116 , n35577 );
    or g14902 ( n17379 , n15070 , n11674 );
    or g14903 ( n14306 , n32639 , n21111 );
    or g14904 ( n27630 , n23572 , n34080 );
    not g14905 ( n35573 , n4065 );
    not g14906 ( n32273 , n16507 );
    not g14907 ( n15778 , n2101 );
    nor g14908 ( n18734 , n15070 , n10375 );
    not g14909 ( n20458 , n12860 );
    and g14910 ( n20721 , n7522 , n40343 );
    or g14911 ( n11385 , n4926 , n918 );
    and g14912 ( n37461 , n4974 , n16071 );
    and g14913 ( n7857 , n9368 , n6266 );
    or g14914 ( n35240 , n41908 , n29545 );
    xnor g14915 ( n31640 , n41013 , n22373 );
    not g14916 ( n22777 , n7125 );
    not g14917 ( n40427 , n22337 );
    nor g14918 ( n22016 , n16598 , n41827 );
    not g14919 ( n21748 , n16666 );
    or g14920 ( n10093 , n13830 , n8601 );
    nor g14921 ( n742 , n2631 , n3648 );
    not g14922 ( n42774 , n40996 );
    or g14923 ( n25432 , n25812 , n14683 );
    not g14924 ( n4448 , n30948 );
    or g14925 ( n39094 , n2567 , n7337 );
    or g14926 ( n25874 , n5009 , n10798 );
    or g14927 ( n38543 , n21325 , n29249 );
    or g14928 ( n3129 , n15070 , n20274 );
    or g14929 ( n16959 , n36155 , n5170 );
    xnor g14930 ( n27440 , n10601 , n1895 );
    or g14931 ( n13884 , n19658 , n40896 );
    and g14932 ( n41081 , n14196 , n22992 );
    not g14933 ( n24154 , n25976 );
    or g14934 ( n17651 , n13830 , n13012 );
    or g14935 ( n554 , n25202 , n35732 );
    xnor g14936 ( n12464 , n7425 , n8289 );
    xnor g14937 ( n2426 , n27399 , n2544 );
    not g14938 ( n27070 , n29617 );
    and g14939 ( n29974 , n31115 , n35088 );
    xnor g14940 ( n31014 , n2471 , n2173 );
    xnor g14941 ( n42863 , n36998 , n5218 );
    or g14942 ( n31962 , n41757 , n7867 );
    not g14943 ( n2263 , n34330 );
    not g14944 ( n27733 , n13753 );
    xnor g14945 ( n9694 , n5144 , n7814 );
    xnor g14946 ( n6093 , n1135 , n33509 );
    and g14947 ( n8090 , n32910 , n461 );
    or g14948 ( n12475 , n41328 , n2989 );
    or g14949 ( n30644 , n36235 , n38429 );
    or g14950 ( n12711 , n33143 , n14153 );
    or g14951 ( n22258 , n1191 , n31997 );
    xnor g14952 ( n15506 , n38749 , n19308 );
    xnor g14953 ( n6207 , n105 , n15977 );
    and g14954 ( n1309 , n22315 , n3411 );
    not g14955 ( n17250 , n20459 );
    or g14956 ( n34203 , n41961 , n35249 );
    or g14957 ( n25095 , n30666 , n20030 );
    or g14958 ( n15845 , n25798 , n30140 );
    and g14959 ( n11808 , n42156 , n26905 );
    or g14960 ( n21989 , n36584 , n21550 );
    not g14961 ( n22493 , n36230 );
    or g14962 ( n33848 , n37707 , n22983 );
    nor g14963 ( n6575 , n28120 , n31513 );
    not g14964 ( n25990 , n39926 );
    nor g14965 ( n6677 , n41325 , n35376 );
    nor g14966 ( n41233 , n15630 , n14015 );
    and g14967 ( n36563 , n38612 , n25387 );
    xnor g14968 ( n17841 , n8739 , n7356 );
    not g14969 ( n11883 , n4452 );
    or g14970 ( n31207 , n26612 , n15900 );
    nor g14971 ( n30253 , n9318 , n12243 );
    or g14972 ( n10772 , n20932 , n10679 );
    nor g14973 ( n1026 , n16489 , n23462 );
    or g14974 ( n2393 , n12718 , n40245 );
    xnor g14975 ( n39248 , n12769 , n22531 );
    xnor g14976 ( n21939 , n29255 , n18641 );
    or g14977 ( n25381 , n11793 , n8038 );
    and g14978 ( n17954 , n29632 , n36645 );
    and g14979 ( n28197 , n24514 , n38984 );
    or g14980 ( n15913 , n1797 , n17104 );
    not g14981 ( n20145 , n22187 );
    or g14982 ( n38015 , n31864 , n6320 );
    or g14983 ( n22770 , n38595 , n3571 );
    nor g14984 ( n32866 , n17120 , n5403 );
    not g14985 ( n35867 , n3619 );
    or g14986 ( n32849 , n33441 , n9302 );
    or g14987 ( n19434 , n15040 , n34764 );
    or g14988 ( n1469 , n17016 , n5986 );
    xnor g14989 ( n7587 , n37335 , n37399 );
    and g14990 ( n41841 , n40986 , n23376 );
    or g14991 ( n15517 , n34561 , n24807 );
    or g14992 ( n42584 , n35165 , n33826 );
    xnor g14993 ( n20160 , n28415 , n23280 );
    or g14994 ( n37485 , n20970 , n28147 );
    xnor g14995 ( n36454 , n19463 , n40116 );
    and g14996 ( n29772 , n22155 , n10917 );
    nor g14997 ( n41058 , n8210 , n16914 );
    nor g14998 ( n26325 , n14026 , n9260 );
    xnor g14999 ( n4151 , n40296 , n11254 );
    not g15000 ( n28711 , n34943 );
    or g15001 ( n4940 , n21610 , n35841 );
    xnor g15002 ( n3782 , n30732 , n8204 );
    or g15003 ( n23911 , n8092 , n11282 );
    nor g15004 ( n24900 , n23252 , n17635 );
    or g15005 ( n39994 , n7956 , n8590 );
    not g15006 ( n35175 , n3124 );
    nor g15007 ( n41353 , n42467 , n40740 );
    nor g15008 ( n29880 , n1110 , n17611 );
    and g15009 ( n4730 , n40889 , n8737 );
    and g15010 ( n35637 , n2966 , n14523 );
    or g15011 ( n4465 , n19997 , n1489 );
    or g15012 ( n33606 , n8087 , n16131 );
    and g15013 ( n37687 , n532 , n4827 );
    or g15014 ( n27749 , n2181 , n30955 );
    xnor g15015 ( n25501 , n3739 , n14369 );
    or g15016 ( n18690 , n40588 , n5322 );
    or g15017 ( n34780 , n25433 , n10064 );
    and g15018 ( n33020 , n9355 , n33516 );
    nor g15019 ( n38684 , n22100 , n12415 );
    or g15020 ( n4364 , n25291 , n41971 );
    or g15021 ( n41334 , n18212 , n41211 );
    and g15022 ( n25575 , n17793 , n12999 );
    not g15023 ( n31184 , n36025 );
    xnor g15024 ( n10602 , n23937 , n28387 );
    or g15025 ( n10126 , n37258 , n7044 );
    xnor g15026 ( n28479 , n38840 , n14471 );
    or g15027 ( n18603 , n18754 , n28947 );
    not g15028 ( n41200 , n23500 );
    not g15029 ( n1186 , n25207 );
    or g15030 ( n11644 , n42234 , n25194 );
    xnor g15031 ( n4683 , n31099 , n39570 );
    and g15032 ( n12265 , n42609 , n23648 );
    or g15033 ( n3019 , n38772 , n3728 );
    and g15034 ( n26640 , n34343 , n40510 );
    and g15035 ( n3567 , n42917 , n4390 );
    not g15036 ( n1092 , n42521 );
    and g15037 ( n5466 , n36593 , n13818 );
    or g15038 ( n31255 , n40490 , n15069 );
    xnor g15039 ( n36529 , n11168 , n38647 );
    or g15040 ( n11262 , n22003 , n12484 );
    or g15041 ( n37881 , n14622 , n37586 );
    nor g15042 ( n19622 , n13855 , n22192 );
    and g15043 ( n8447 , n7115 , n14227 );
    or g15044 ( n8603 , n12084 , n5124 );
    or g15045 ( n1532 , n7041 , n32256 );
    or g15046 ( n39787 , n33624 , n27017 );
    or g15047 ( n27215 , n39439 , n8526 );
    or g15048 ( n3253 , n9748 , n13294 );
    or g15049 ( n25586 , n15423 , n21564 );
    or g15050 ( n4902 , n21178 , n26816 );
    or g15051 ( n24524 , n8199 , n23424 );
    or g15052 ( n22334 , n14859 , n28887 );
    or g15053 ( n36908 , n21048 , n25937 );
    and g15054 ( n26931 , n30038 , n12074 );
    and g15055 ( n18428 , n5005 , n34662 );
    or g15056 ( n780 , n11548 , n1044 );
    not g15057 ( n1374 , n23442 );
    not g15058 ( n25297 , n13158 );
    or g15059 ( n27143 , n19523 , n32988 );
    nor g15060 ( n10818 , n27051 , n39045 );
    nor g15061 ( n1669 , n31677 , n32580 );
    not g15062 ( n30995 , n30119 );
    and g15063 ( n31307 , n31974 , n41911 );
    xnor g15064 ( n37738 , n9783 , n2870 );
    or g15065 ( n39211 , n13043 , n12730 );
    or g15066 ( n13117 , n13526 , n40032 );
    or g15067 ( n31448 , n38571 , n21092 );
    xnor g15068 ( n9237 , n2839 , n12366 );
    not g15069 ( n378 , n23170 );
    not g15070 ( n30572 , n1758 );
    nor g15071 ( n17337 , n31471 , n24538 );
    not g15072 ( n4842 , n39392 );
    not g15073 ( n30298 , n5816 );
    xnor g15074 ( n37536 , n39760 , n2924 );
    xnor g15075 ( n2539 , n10168 , n17120 );
    nor g15076 ( n13843 , n35301 , n20436 );
    or g15077 ( n18996 , n40852 , n12574 );
    nor g15078 ( n17067 , n15800 , n24738 );
    and g15079 ( n4502 , n32778 , n5765 );
    xnor g15080 ( n32609 , n18509 , n10876 );
    nor g15081 ( n5391 , n42063 , n15394 );
    and g15082 ( n775 , n3923 , n250 );
    or g15083 ( n7834 , n29880 , n35198 );
    and g15084 ( n7732 , n34568 , n24201 );
    and g15085 ( n36371 , n28940 , n13946 );
    or g15086 ( n5597 , n12484 , n33957 );
    not g15087 ( n22303 , n31336 );
    nor g15088 ( n4011 , n35727 , n29878 );
    and g15089 ( n33824 , n23107 , n14926 );
    or g15090 ( n11652 , n31390 , n38573 );
    and g15091 ( n23808 , n6829 , n20308 );
    xnor g15092 ( n40099 , n16693 , n2666 );
    or g15093 ( n29868 , n7552 , n18581 );
    or g15094 ( n3611 , n26354 , n3750 );
    xnor g15095 ( n30454 , n542 , n13733 );
    xnor g15096 ( n25690 , n18657 , n35671 );
    nor g15097 ( n27494 , n41715 , n14561 );
    nor g15098 ( n14973 , n9394 , n13402 );
    nor g15099 ( n42508 , n26974 , n8511 );
    xnor g15100 ( n21362 , n22237 , n39610 );
    and g15101 ( n21814 , n32497 , n24788 );
    xnor g15102 ( n37383 , n20920 , n2977 );
    xnor g15103 ( n2000 , n38893 , n2678 );
    xnor g15104 ( n9362 , n22842 , n13355 );
    xnor g15105 ( n11819 , n4558 , n10242 );
    nor g15106 ( n41679 , n38974 , n23389 );
    or g15107 ( n39929 , n10972 , n25742 );
    xnor g15108 ( n1505 , n5237 , n31311 );
    or g15109 ( n6433 , n40296 , n6693 );
    and g15110 ( n38981 , n4693 , n16828 );
    or g15111 ( n22434 , n27924 , n853 );
    or g15112 ( n3553 , n25600 , n10217 );
    or g15113 ( n41295 , n18784 , n30496 );
    or g15114 ( n20609 , n27823 , n803 );
    or g15115 ( n16037 , n23473 , n8714 );
    or g15116 ( n2420 , n34001 , n33826 );
    or g15117 ( n19341 , n16207 , n7314 );
    or g15118 ( n35444 , n26938 , n34502 );
    xnor g15119 ( n26621 , n34562 , n21722 );
    or g15120 ( n2973 , n42382 , n15468 );
    and g15121 ( n788 , n5312 , n40248 );
    or g15122 ( n7959 , n20633 , n2258 );
    or g15123 ( n29706 , n18916 , n20865 );
    nor g15124 ( n40924 , n39266 , n1969 );
    or g15125 ( n23160 , n1470 , n22210 );
    or g15126 ( n17639 , n16052 , n23265 );
    nor g15127 ( n28699 , n17193 , n27431 );
    or g15128 ( n20147 , n22371 , n7966 );
    xnor g15129 ( n33379 , n18192 , n31747 );
    and g15130 ( n34849 , n34175 , n649 );
    or g15131 ( n33452 , n23745 , n39241 );
    nor g15132 ( n28168 , n15988 , n19016 );
    and g15133 ( n12663 , n23612 , n37366 );
    xnor g15134 ( n25574 , n28377 , n15265 );
    not g15135 ( n30443 , n36920 );
    nor g15136 ( n38402 , n4527 , n198 );
    and g15137 ( n6419 , n32033 , n17408 );
    or g15138 ( n12387 , n5340 , n26107 );
    xnor g15139 ( n19644 , n2620 , n17228 );
    or g15140 ( n5579 , n21402 , n12632 );
    or g15141 ( n37888 , n18197 , n27028 );
    nor g15142 ( n5932 , n34565 , n26988 );
    or g15143 ( n3842 , n980 , n15564 );
    and g15144 ( n40479 , n23195 , n3578 );
    and g15145 ( n21919 , n28694 , n36058 );
    and g15146 ( n11908 , n34603 , n18057 );
    nor g15147 ( n34930 , n22538 , n19942 );
    nor g15148 ( n33077 , n1507 , n35023 );
    and g15149 ( n30143 , n33406 , n3869 );
    and g15150 ( n30404 , n35206 , n21323 );
    or g15151 ( n21785 , n32062 , n22462 );
    xnor g15152 ( n19726 , n26199 , n10977 );
    not g15153 ( n7282 , n18134 );
    xnor g15154 ( n33001 , n33241 , n3834 );
    not g15155 ( n35347 , n41969 );
    or g15156 ( n40049 , n40295 , n13022 );
    or g15157 ( n24616 , n25846 , n30788 );
    nor g15158 ( n12334 , n38879 , n575 );
    xnor g15159 ( n37955 , n34382 , n39156 );
    and g15160 ( n21510 , n29759 , n27778 );
    or g15161 ( n32948 , n39663 , n41993 );
    and g15162 ( n42614 , n1881 , n35519 );
    and g15163 ( n10290 , n34602 , n22390 );
    or g15164 ( n25220 , n9263 , n36619 );
    not g15165 ( n10867 , n7532 );
    or g15166 ( n31404 , n32206 , n1044 );
    or g15167 ( n33830 , n781 , n788 );
    or g15168 ( n28163 , n33382 , n33345 );
    not g15169 ( n9329 , n34274 );
    or g15170 ( n2033 , n17293 , n21410 );
    and g15171 ( n19643 , n27844 , n5247 );
    nor g15172 ( n27006 , n26509 , n39335 );
    or g15173 ( n10706 , n35984 , n37477 );
    nor g15174 ( n38500 , n36721 , n21271 );
    and g15175 ( n38165 , n1826 , n36149 );
    or g15176 ( n13262 , n13600 , n15462 );
    not g15177 ( n38531 , n26985 );
    or g15178 ( n27456 , n30825 , n24040 );
    or g15179 ( n24578 , n21483 , n40455 );
    nor g15180 ( n42123 , n39640 , n20532 );
    xnor g15181 ( n2402 , n6625 , n4650 );
    not g15182 ( n37376 , n38389 );
    xnor g15183 ( n30465 , n784 , n32183 );
    nor g15184 ( n21779 , n26848 , n37475 );
    or g15185 ( n5376 , n32266 , n18946 );
    or g15186 ( n36519 , n18224 , n40592 );
    or g15187 ( n42434 , n20825 , n17229 );
    xnor g15188 ( n42436 , n42064 , n2172 );
    or g15189 ( n2875 , n6677 , n31227 );
    or g15190 ( n12563 , n34597 , n5243 );
    and g15191 ( n30672 , n25439 , n6938 );
    or g15192 ( n30310 , n11673 , n41767 );
    or g15193 ( n8650 , n30238 , n17109 );
    or g15194 ( n21417 , n14489 , n15327 );
    or g15195 ( n20917 , n15101 , n16982 );
    and g15196 ( n41999 , n9204 , n19715 );
    not g15197 ( n24176 , n11316 );
    and g15198 ( n8550 , n3448 , n18556 );
    or g15199 ( n26720 , n19985 , n5614 );
    or g15200 ( n41965 , n17124 , n32445 );
    or g15201 ( n33764 , n34275 , n41891 );
    xnor g15202 ( n22461 , n22604 , n34743 );
    and g15203 ( n25802 , n32710 , n15862 );
    or g15204 ( n24989 , n36548 , n14569 );
    or g15205 ( n18598 , n37119 , n4701 );
    or g15206 ( n22999 , n4787 , n15659 );
    not g15207 ( n8483 , n41508 );
    not g15208 ( n31302 , n15623 );
    and g15209 ( n20369 , n28399 , n22045 );
    or g15210 ( n20144 , n12495 , n10603 );
    or g15211 ( n23271 , n5065 , n21026 );
    and g15212 ( n39958 , n30258 , n37486 );
    nor g15213 ( n33355 , n9597 , n40563 );
    not g15214 ( n38708 , n11731 );
    and g15215 ( n8902 , n7943 , n3166 );
    not g15216 ( n37088 , n17738 );
    nor g15217 ( n36062 , n8591 , n8814 );
    or g15218 ( n26940 , n11749 , n31918 );
    not g15219 ( n3781 , n17252 );
    and g15220 ( n230 , n24813 , n29400 );
    or g15221 ( n22305 , n23352 , n14578 );
    nor g15222 ( n11270 , n22100 , n5770 );
    and g15223 ( n2143 , n34441 , n373 );
    or g15224 ( n40174 , n23114 , n7616 );
    not g15225 ( n22872 , n2932 );
    and g15226 ( n27052 , n14241 , n2760 );
    xnor g15227 ( n15305 , n36454 , n20805 );
    or g15228 ( n18163 , n9920 , n11340 );
    or g15229 ( n34815 , n29473 , n13675 );
    or g15230 ( n26452 , n12397 , n30717 );
    and g15231 ( n29969 , n26004 , n20091 );
    or g15232 ( n445 , n18367 , n42828 );
    nor g15233 ( n16981 , n31256 , n41977 );
    or g15234 ( n34876 , n25970 , n7172 );
    xnor g15235 ( n34177 , n34325 , n24795 );
    nor g15236 ( n10731 , n34492 , n27657 );
    and g15237 ( n33976 , n3944 , n18295 );
    or g15238 ( n8521 , n17193 , n10108 );
    and g15239 ( n5262 , n28276 , n8041 );
    or g15240 ( n8835 , n19067 , n18964 );
    xnor g15241 ( n8633 , n7489 , n11478 );
    xnor g15242 ( n38626 , n3769 , n30800 );
    or g15243 ( n6880 , n6558 , n16315 );
    xnor g15244 ( n17368 , n4334 , n21378 );
    xnor g15245 ( n22047 , n30139 , n28848 );
    and g15246 ( n27363 , n667 , n8236 );
    xnor g15247 ( n19822 , n21726 , n18866 );
    or g15248 ( n27727 , n22602 , n2507 );
    nor g15249 ( n39963 , n21382 , n10474 );
    or g15250 ( n9613 , n12429 , n13758 );
    not g15251 ( n26021 , n34118 );
    or g15252 ( n27867 , n40389 , n21444 );
    xnor g15253 ( n33987 , n22827 , n11859 );
    nor g15254 ( n22624 , n2183 , n9801 );
    or g15255 ( n39029 , n38074 , n4456 );
    or g15256 ( n12428 , n32307 , n42025 );
    xnor g15257 ( n2461 , n12146 , n28571 );
    or g15258 ( n31915 , n40086 , n1716 );
    or g15259 ( n39157 , n20138 , n4661 );
    or g15260 ( n7449 , n30306 , n1578 );
    and g15261 ( n18429 , n30088 , n18122 );
    or g15262 ( n29157 , n7313 , n19472 );
    or g15263 ( n36791 , n19184 , n38175 );
    xnor g15264 ( n23668 , n37153 , n4699 );
    or g15265 ( n21775 , n36296 , n9840 );
    or g15266 ( n38470 , n19303 , n40178 );
    nor g15267 ( n20271 , n6303 , n27871 );
    nor g15268 ( n41548 , n24892 , n189 );
    nor g15269 ( n2212 , n35215 , n24285 );
    and g15270 ( n12388 , n31765 , n9026 );
    not g15271 ( n6786 , n7327 );
    and g15272 ( n35340 , n37464 , n22630 );
    nor g15273 ( n16613 , n33038 , n31970 );
    xnor g15274 ( n29479 , n38906 , n24988 );
    nor g15275 ( n1750 , n10833 , n22104 );
    or g15276 ( n24804 , n94 , n6570 );
    xnor g15277 ( n11697 , n36998 , n26573 );
    or g15278 ( n42085 , n7020 , n7812 );
    or g15279 ( n29907 , n14287 , n10069 );
    xnor g15280 ( n4163 , n2645 , n17901 );
    or g15281 ( n17041 , n17268 , n24665 );
    and g15282 ( n38737 , n42432 , n9870 );
    or g15283 ( n25224 , n10674 , n3192 );
    or g15284 ( n37943 , n11404 , n9128 );
    not g15285 ( n22002 , n33861 );
    or g15286 ( n35271 , n39991 , n31066 );
    or g15287 ( n24047 , n40967 , n11769 );
    not g15288 ( n14885 , n14920 );
    nor g15289 ( n14300 , n34292 , n19748 );
    nor g15290 ( n2740 , n14125 , n32811 );
    or g15291 ( n40847 , n20196 , n28143 );
    nor g15292 ( n17709 , n37639 , n5678 );
    and g15293 ( n15787 , n36614 , n39222 );
    or g15294 ( n976 , n2199 , n39848 );
    xnor g15295 ( n33938 , n5144 , n3563 );
    not g15296 ( n17843 , n23043 );
    or g15297 ( n25052 , n7746 , n28309 );
    or g15298 ( n33949 , n9265 , n16636 );
    or g15299 ( n20301 , n34988 , n15573 );
    or g15300 ( n1822 , n15758 , n6135 );
    or g15301 ( n29112 , n13247 , n26740 );
    or g15302 ( n33506 , n18597 , n12976 );
    or g15303 ( n12747 , n21024 , n34655 );
    or g15304 ( n8404 , n28617 , n37468 );
    nor g15305 ( n16027 , n33981 , n27546 );
    and g15306 ( n40516 , n5899 , n37341 );
    not g15307 ( n12411 , n19288 );
    not g15308 ( n37692 , n41655 );
    or g15309 ( n2195 , n7506 , n42661 );
    or g15310 ( n8334 , n24454 , n41443 );
    or g15311 ( n41073 , n4798 , n9278 );
    or g15312 ( n4831 , n8716 , n38196 );
    not g15313 ( n42782 , n25159 );
    not g15314 ( n24198 , n31561 );
    or g15315 ( n15286 , n31648 , n9129 );
    not g15316 ( n11023 , n18134 );
    or g15317 ( n18730 , n16753 , n29073 );
    nor g15318 ( n40840 , n36117 , n19915 );
    and g15319 ( n22614 , n36228 , n17443 );
    nor g15320 ( n2752 , n23980 , n201 );
    not g15321 ( n4208 , n4147 );
    or g15322 ( n12528 , n1550 , n16530 );
    xnor g15323 ( n6488 , n2921 , n35779 );
    xnor g15324 ( n42848 , n13444 , n14695 );
    xnor g15325 ( n19907 , n18678 , n36652 );
    or g15326 ( n18135 , n30068 , n7371 );
    or g15327 ( n32416 , n27080 , n39328 );
    and g15328 ( n24348 , n35800 , n37975 );
    and g15329 ( n52 , n27160 , n31281 );
    or g15330 ( n8820 , n25878 , n8640 );
    and g15331 ( n5016 , n21001 , n33830 );
    nor g15332 ( n41069 , n11057 , n8324 );
    or g15333 ( n39953 , n4140 , n6187 );
    not g15334 ( n8968 , n24510 );
    and g15335 ( n19123 , n28439 , n37971 );
    nor g15336 ( n27341 , n11489 , n8651 );
    not g15337 ( n16198 , n12533 );
    nor g15338 ( n36649 , n39559 , n21446 );
    or g15339 ( n1463 , n35633 , n733 );
    xnor g15340 ( n27354 , n34691 , n13797 );
    not g15341 ( n13612 , n31837 );
    or g15342 ( n8915 , n21116 , n30981 );
    and g15343 ( n27165 , n37858 , n19105 );
    or g15344 ( n3095 , n41928 , n40787 );
    or g15345 ( n4785 , n39621 , n38416 );
    xnor g15346 ( n14214 , n41811 , n34256 );
    not g15347 ( n22899 , n16253 );
    and g15348 ( n6126 , n28943 , n9780 );
    or g15349 ( n40806 , n11895 , n4727 );
    or g15350 ( n20559 , n16117 , n25269 );
    or g15351 ( n13201 , n34460 , n17349 );
    or g15352 ( n18069 , n19082 , n2710 );
    not g15353 ( n32068 , n41758 );
    not g15354 ( n40618 , n39 );
    or g15355 ( n11580 , n42798 , n7046 );
    not g15356 ( n28949 , n11264 );
    and g15357 ( n25401 , n16932 , n42189 );
    xnor g15358 ( n30040 , n40889 , n8737 );
    and g15359 ( n18950 , n18979 , n16543 );
    or g15360 ( n12869 , n3462 , n41152 );
    nor g15361 ( n26044 , n17436 , n23872 );
    not g15362 ( n10220 , n25653 );
    not g15363 ( n23971 , n23285 );
    not g15364 ( n20157 , n1794 );
    xnor g15365 ( n23209 , n33917 , n28262 );
    nor g15366 ( n17199 , n38879 , n22985 );
    nor g15367 ( n39688 , n7963 , n4166 );
    xnor g15368 ( n9944 , n302 , n4267 );
    and g15369 ( n35180 , n12989 , n36503 );
    and g15370 ( n30871 , n25874 , n17185 );
    not g15371 ( n10315 , n9405 );
    or g15372 ( n36783 , n29932 , n32161 );
    or g15373 ( n1136 , n12947 , n27435 );
    nor g15374 ( n20343 , n39266 , n21280 );
    not g15375 ( n39176 , n15004 );
    not g15376 ( n313 , n3084 );
    nor g15377 ( n3712 , n30490 , n33082 );
    or g15378 ( n3987 , n4256 , n2034 );
    or g15379 ( n31842 , n28080 , n3258 );
    and g15380 ( n33054 , n14760 , n30576 );
    not g15381 ( n38284 , n27519 );
    and g15382 ( n31637 , n36046 , n18291 );
    or g15383 ( n15066 , n16899 , n7931 );
    and g15384 ( n26423 , n2864 , n16889 );
    and g15385 ( n42494 , n760 , n27583 );
    or g15386 ( n36678 , n31123 , n8223 );
    or g15387 ( n31980 , n29447 , n35111 );
    or g15388 ( n18704 , n5618 , n36067 );
    or g15389 ( n31183 , n21915 , n37835 );
    or g15390 ( n12865 , n21698 , n22217 );
    or g15391 ( n15414 , n10037 , n28725 );
    or g15392 ( n5231 , n4559 , n12020 );
    nor g15393 ( n4464 , n22403 , n18356 );
    or g15394 ( n5967 , n33948 , n29176 );
    or g15395 ( n39016 , n8369 , n25178 );
    or g15396 ( n27772 , n16586 , n3787 );
    or g15397 ( n5395 , n18051 , n30587 );
    or g15398 ( n36531 , n38613 , n27385 );
    or g15399 ( n31331 , n41819 , n24606 );
    xnor g15400 ( n25815 , n31989 , n38999 );
    xnor g15401 ( n32106 , n3317 , n40571 );
    nor g15402 ( n21032 , n5964 , n9876 );
    or g15403 ( n24873 , n37569 , n36673 );
    or g15404 ( n30481 , n11921 , n27127 );
    xnor g15405 ( n12300 , n27907 , n41102 );
    nor g15406 ( n27773 , n35142 , n38155 );
    xnor g15407 ( n24382 , n29174 , n6535 );
    or g15408 ( n25887 , n37990 , n5444 );
    not g15409 ( n11538 , n36030 );
    xnor g15410 ( n1925 , n7943 , n1975 );
    xnor g15411 ( n36513 , n17872 , n2525 );
    or g15412 ( n41852 , n12902 , n40481 );
    or g15413 ( n5714 , n32100 , n14722 );
    or g15414 ( n18579 , n11478 , n22920 );
    not g15415 ( n26623 , n34051 );
    xnor g15416 ( n30608 , n3080 , n3414 );
    or g15417 ( n7925 , n36848 , n11763 );
    or g15418 ( n815 , n31997 , n11320 );
    or g15419 ( n454 , n31889 , n3571 );
    or g15420 ( n3491 , n41964 , n18026 );
    not g15421 ( n31135 , n22642 );
    xnor g15422 ( n21305 , n18530 , n1969 );
    and g15423 ( n18456 , n1864 , n4968 );
    and g15424 ( n37872 , n37601 , n11027 );
    xnor g15425 ( n25301 , n17377 , n41438 );
    and g15426 ( n41376 , n2071 , n14629 );
    and g15427 ( n23698 , n39855 , n33483 );
    and g15428 ( n30349 , n17219 , n24150 );
    nor g15429 ( n9189 , n14821 , n13580 );
    or g15430 ( n23900 , n12945 , n31008 );
    not g15431 ( n25701 , n16699 );
    or g15432 ( n13966 , n28076 , n42423 );
    or g15433 ( n34556 , n36499 , n22456 );
    nor g15434 ( n79 , n10950 , n14653 );
    and g15435 ( n11619 , n10847 , n39102 );
    not g15436 ( n1932 , n7343 );
    or g15437 ( n8564 , n38022 , n27512 );
    or g15438 ( n41365 , n1377 , n40278 );
    not g15439 ( n41562 , n38049 );
    or g15440 ( n36794 , n33926 , n38123 );
    or g15441 ( n21968 , n31888 , n42636 );
    or g15442 ( n3027 , n19348 , n16752 );
    or g15443 ( n21423 , n12397 , n34406 );
    nor g15444 ( n28173 , n40222 , n7580 );
    nor g15445 ( n29385 , n7613 , n41594 );
    and g15446 ( n823 , n25117 , n40442 );
    or g15447 ( n35792 , n20338 , n39152 );
    nor g15448 ( n13765 , n38879 , n42006 );
    nor g15449 ( n33781 , n2449 , n17916 );
    and g15450 ( n16990 , n19916 , n1671 );
    and g15451 ( n32095 , n6574 , n23996 );
    or g15452 ( n22202 , n31150 , n25504 );
    or g15453 ( n22229 , n28774 , n23009 );
    not g15454 ( n19742 , n25283 );
    or g15455 ( n3983 , n5679 , n37043 );
    nor g15456 ( n19777 , n91 , n4542 );
    xnor g15457 ( n22940 , n24159 , n23860 );
    or g15458 ( n38608 , n10685 , n7265 );
    or g15459 ( n33514 , n26978 , n29686 );
    xnor g15460 ( n2905 , n6147 , n19966 );
    or g15461 ( n29093 , n14796 , n11712 );
    or g15462 ( n21468 , n41493 , n10646 );
    or g15463 ( n21443 , n27796 , n35880 );
    nor g15464 ( n24736 , n4129 , n28318 );
    and g15465 ( n15271 , n41551 , n36794 );
    not g15466 ( n5977 , n33988 );
    or g15467 ( n11226 , n31666 , n29312 );
    nor g15468 ( n468 , n35887 , n27816 );
    or g15469 ( n42910 , n39266 , n23561 );
    and g15470 ( n41812 , n28305 , n10225 );
    or g15471 ( n41982 , n40973 , n33859 );
    and g15472 ( n431 , n5008 , n27826 );
    and g15473 ( n11977 , n15636 , n8416 );
    not g15474 ( n22470 , n16755 );
    and g15475 ( n4311 , n14473 , n18290 );
    and g15476 ( n18719 , n8885 , n41742 );
    or g15477 ( n24960 , n19486 , n39675 );
    or g15478 ( n1433 , n35534 , n41619 );
    and g15479 ( n8180 , n22066 , n13761 );
    or g15480 ( n27847 , n39991 , n38744 );
    and g15481 ( n4028 , n30789 , n37930 );
    or g15482 ( n19546 , n3567 , n25824 );
    not g15483 ( n8518 , n28734 );
    or g15484 ( n12775 , n33887 , n34672 );
    and g15485 ( n11868 , n3319 , n32000 );
    xnor g15486 ( n502 , n836 , n13629 );
    or g15487 ( n24837 , n2859 , n12640 );
    not g15488 ( n2062 , n7824 );
    or g15489 ( n32026 , n30820 , n34328 );
    and g15490 ( n34715 , n15194 , n3461 );
    nor g15491 ( n28985 , n34686 , n19000 );
    or g15492 ( n31377 , n25750 , n3780 );
    nor g15493 ( n34044 , n34565 , n39753 );
    xnor g15494 ( n25306 , n27250 , n24015 );
    or g15495 ( n31630 , n37014 , n26385 );
    not g15496 ( n31618 , n14233 );
    not g15497 ( n27388 , n4784 );
    xnor g15498 ( n14801 , n13415 , n35981 );
    or g15499 ( n33879 , n35802 , n15720 );
    or g15500 ( n23644 , n31468 , n14703 );
    and g15501 ( n14312 , n27614 , n21728 );
    or g15502 ( n31487 , n433 , n17160 );
    and g15503 ( n30587 , n33290 , n23306 );
    not g15504 ( n18530 , n39266 );
    or g15505 ( n1958 , n12676 , n12286 );
    or g15506 ( n23499 , n40855 , n36687 );
    not g15507 ( n30125 , n6714 );
    not g15508 ( n8569 , n27446 );
    not g15509 ( n26587 , n20820 );
    or g15510 ( n33992 , n40588 , n1059 );
    not g15511 ( n39405 , n5332 );
    or g15512 ( n9656 , n32104 , n39092 );
    or g15513 ( n30375 , n1504 , n4355 );
    or g15514 ( n25807 , n24378 , n1828 );
    or g15515 ( n25455 , n8056 , n5610 );
    or g15516 ( n18358 , n39811 , n27510 );
    nor g15517 ( n10701 , n40558 , n12682 );
    and g15518 ( n3694 , n11055 , n24089 );
    or g15519 ( n26796 , n41998 , n38088 );
    and g15520 ( n3323 , n23324 , n11355 );
    or g15521 ( n17191 , n10986 , n27921 );
    and g15522 ( n39063 , n357 , n39782 );
    or g15523 ( n32911 , n2631 , n37408 );
    and g15524 ( n13609 , n1741 , n3375 );
    and g15525 ( n40944 , n4837 , n22466 );
    and g15526 ( n17901 , n11954 , n24004 );
    or g15527 ( n33158 , n7356 , n8739 );
    not g15528 ( n31475 , n30287 );
    not g15529 ( n9031 , n7508 );
    nor g15530 ( n23682 , n4410 , n12178 );
    not g15531 ( n19244 , n31193 );
    and g15532 ( n11284 , n39322 , n28422 );
    or g15533 ( n4197 , n2711 , n2061 );
    or g15534 ( n21909 , n2593 , n28339 );
    or g15535 ( n13408 , n25331 , n35058 );
    nor g15536 ( n17575 , n42115 , n23013 );
    xnor g15537 ( n26117 , n38261 , n9521 );
    or g15538 ( n40891 , n36405 , n21696 );
    and g15539 ( n39171 , n7462 , n37927 );
    or g15540 ( n27989 , n25100 , n1289 );
    xnor g15541 ( n37831 , n39279 , n28969 );
    nor g15542 ( n21295 , n6939 , n40355 );
    not g15543 ( n33120 , n24397 );
    not g15544 ( n24018 , n36246 );
    and g15545 ( n22980 , n34667 , n11098 );
    or g15546 ( n22332 , n586 , n31582 );
    or g15547 ( n42918 , n36951 , n25964 );
    and g15548 ( n20616 , n28990 , n22510 );
    or g15549 ( n6117 , n23374 , n24206 );
    xnor g15550 ( n3214 , n4491 , n8088 );
    not g15551 ( n26576 , n2996 );
    or g15552 ( n16844 , n19374 , n8087 );
    and g15553 ( n5342 , n25525 , n8379 );
    and g15554 ( n19563 , n30181 , n42028 );
    not g15555 ( n20092 , n2529 );
    not g15556 ( n17205 , n140 );
    or g15557 ( n26929 , n4096 , n22333 );
    xnor g15558 ( n11211 , n34210 , n35891 );
    nor g15559 ( n30730 , n33070 , n31152 );
    xnor g15560 ( n2065 , n17661 , n38089 );
    or g15561 ( n13142 , n41752 , n31686 );
    or g15562 ( n20216 , n31215 , n6415 );
    or g15563 ( n21656 , n9832 , n12768 );
    and g15564 ( n39187 , n19700 , n1621 );
    xnor g15565 ( n10725 , n41947 , n15084 );
    or g15566 ( n38642 , n28545 , n2290 );
    or g15567 ( n23016 , n29797 , n40475 );
    or g15568 ( n37311 , n5029 , n8777 );
    and g15569 ( n7209 , n5108 , n2306 );
    or g15570 ( n24533 , n38085 , n27988 );
    not g15571 ( n6263 , n23960 );
    or g15572 ( n29109 , n5555 , n36979 );
    not g15573 ( n27020 , n4404 );
    or g15574 ( n5924 , n41819 , n42221 );
    not g15575 ( n11830 , n3137 );
    xnor g15576 ( n11649 , n20310 , n23872 );
    not g15577 ( n25826 , n29474 );
    or g15578 ( n13942 , n28122 , n12059 );
    or g15579 ( n21516 , n19769 , n30573 );
    nor g15580 ( n32010 , n9001 , n8011 );
    xnor g15581 ( n39167 , n14242 , n19460 );
    xnor g15582 ( n15883 , n6308 , n24999 );
    and g15583 ( n14383 , n28653 , n20462 );
    xnor g15584 ( n9895 , n16693 , n41448 );
    nor g15585 ( n2853 , n19808 , n25790 );
    not g15586 ( n39602 , n13201 );
    or g15587 ( n34055 , n2927 , n14967 );
    nor g15588 ( n28970 , n21729 , n12338 );
    not g15589 ( n15368 , n20698 );
    and g15590 ( n7050 , n26981 , n10596 );
    nor g15591 ( n19694 , n27653 , n20129 );
    not g15592 ( n17634 , n31259 );
    nor g15593 ( n10182 , n36228 , n17443 );
    and g15594 ( n40437 , n18766 , n24434 );
    not g15595 ( n23318 , n25094 );
    or g15596 ( n25555 , n42466 , n41213 );
    not g15597 ( n11349 , n5147 );
    nor g15598 ( n26785 , n13338 , n18271 );
    or g15599 ( n17091 , n1004 , n41413 );
    or g15600 ( n38995 , n40350 , n3421 );
    or g15601 ( n6979 , n28683 , n32163 );
    nor g15602 ( n27136 , n1507 , n9000 );
    and g15603 ( n4933 , n30098 , n28764 );
    and g15604 ( n32123 , n13928 , n31708 );
    or g15605 ( n27084 , n23472 , n15473 );
    not g15606 ( n15138 , n22917 );
    or g15607 ( n40830 , n35835 , n33464 );
    not g15608 ( n38154 , n39048 );
    and g15609 ( n36197 , n7677 , n37215 );
    not g15610 ( n17476 , n8663 );
    not g15611 ( n25907 , n29777 );
    not g15612 ( n16766 , n1206 );
    not g15613 ( n39015 , n8308 );
    not g15614 ( n18859 , n21675 );
    not g15615 ( n376 , n26076 );
    or g15616 ( n4674 , n5538 , n7117 );
    or g15617 ( n20586 , n28198 , n5120 );
    and g15618 ( n7862 , n3755 , n33726 );
    or g15619 ( n42081 , n37031 , n1837 );
    or g15620 ( n10800 , n10906 , n9040 );
    nor g15621 ( n20914 , n24200 , n6798 );
    or g15622 ( n31407 , n14314 , n7853 );
    nor g15623 ( n16985 , n24200 , n4486 );
    and g15624 ( n7429 , n37322 , n29769 );
    not g15625 ( n30022 , n24800 );
    or g15626 ( n24434 , n36052 , n17390 );
    and g15627 ( n25132 , n32643 , n22960 );
    not g15628 ( n36415 , n21394 );
    or g15629 ( n6317 , n2244 , n22767 );
    nor g15630 ( n7194 , n26186 , n14521 );
    or g15631 ( n3723 , n42076 , n24521 );
    xnor g15632 ( n19680 , n21877 , n40838 );
    or g15633 ( n2264 , n40459 , n25897 );
    nor g15634 ( n37266 , n1073 , n2017 );
    or g15635 ( n9904 , n18244 , n4682 );
    and g15636 ( n33243 , n20516 , n8237 );
    or g15637 ( n3844 , n35359 , n26424 );
    and g15638 ( n27269 , n35462 , n29749 );
    xnor g15639 ( n18839 , n31989 , n16508 );
    nor g15640 ( n34403 , n24368 , n37295 );
    or g15641 ( n15304 , n26490 , n6018 );
    not g15642 ( n20410 , n25516 );
    nor g15643 ( n31812 , n35709 , n2574 );
    xnor g15644 ( n32157 , n35961 , n27770 );
    or g15645 ( n2773 , n35915 , n37373 );
    not g15646 ( n40157 , n17406 );
    nor g15647 ( n21140 , n28501 , n9284 );
    or g15648 ( n35517 , n8721 , n15737 );
    or g15649 ( n42445 , n36456 , n33372 );
    and g15650 ( n22683 , n37861 , n4199 );
    not g15651 ( n21876 , n18429 );
    and g15652 ( n35016 , n22011 , n39228 );
    or g15653 ( n18692 , n25129 , n14749 );
    or g15654 ( n21576 , n35524 , n31417 );
    and g15655 ( n13340 , n16358 , n29765 );
    not g15656 ( n15646 , n22331 );
    and g15657 ( n40478 , n26940 , n30553 );
    or g15658 ( n22658 , n2172 , n29382 );
    and g15659 ( n8127 , n6603 , n11175 );
    or g15660 ( n14413 , n34565 , n40335 );
    or g15661 ( n23870 , n21703 , n10155 );
    and g15662 ( n38078 , n33967 , n3742 );
    and g15663 ( n14068 , n13460 , n31583 );
    nor g15664 ( n10869 , n3687 , n32564 );
    or g15665 ( n11777 , n3886 , n11074 );
    not g15666 ( n23904 , n8446 );
    nor g15667 ( n18299 , n24879 , n40287 );
    not g15668 ( n5390 , n28182 );
    not g15669 ( n35497 , n25794 );
    or g15670 ( n6068 , n18314 , n1950 );
    or g15671 ( n20745 , n19729 , n2768 );
    nor g15672 ( n20975 , n30743 , n17258 );
    or g15673 ( n31749 , n19397 , n34485 );
    not g15674 ( n27566 , n7546 );
    or g15675 ( n13053 , n41356 , n6093 );
    xnor g15676 ( n26733 , n42567 , n2881 );
    not g15677 ( n38921 , n12318 );
    or g15678 ( n14336 , n21218 , n16999 );
    nor g15679 ( n12016 , n38821 , n274 );
    or g15680 ( n37525 , n40378 , n1533 );
    not g15681 ( n39236 , n21005 );
    or g15682 ( n36349 , n29290 , n32752 );
    and g15683 ( n30696 , n29753 , n20502 );
    or g15684 ( n16176 , n41957 , n32946 );
    and g15685 ( n12086 , n18201 , n36916 );
    or g15686 ( n38194 , n12442 , n42654 );
    or g15687 ( n36730 , n6327 , n5771 );
    not g15688 ( n5881 , n2018 );
    xnor g15689 ( n4731 , n41098 , n40784 );
    or g15690 ( n17106 , n17061 , n38196 );
    or g15691 ( n7455 , n21893 , n22914 );
    and g15692 ( n3941 , n23679 , n16656 );
    nor g15693 ( n33760 , n186 , n19308 );
    or g15694 ( n33192 , n27552 , n31894 );
    or g15695 ( n31909 , n8862 , n28370 );
    not g15696 ( n2036 , n13661 );
    xnor g15697 ( n8084 , n7489 , n29259 );
    xnor g15698 ( n2989 , n2222 , n32493 );
    or g15699 ( n29617 , n15368 , n34711 );
    and g15700 ( n107 , n6457 , n40525 );
    nor g15701 ( n34759 , n3092 , n19661 );
    nor g15702 ( n30522 , n7004 , n18730 );
    or g15703 ( n4406 , n4798 , n16113 );
    or g15704 ( n30202 , n14308 , n21655 );
    and g15705 ( n22533 , n5352 , n26589 );
    or g15706 ( n25941 , n11904 , n17963 );
    xnor g15707 ( n22561 , n41764 , n8929 );
    not g15708 ( n38378 , n3619 );
    nor g15709 ( n17686 , n17744 , n18114 );
    xnor g15710 ( n41025 , n2722 , n34941 );
    and g15711 ( n18273 , n29275 , n30910 );
    xnor g15712 ( n26952 , n20557 , n22512 );
    and g15713 ( n36431 , n28560 , n3926 );
    or g15714 ( n36699 , n31761 , n3790 );
    xnor g15715 ( n24781 , n14037 , n8570 );
    not g15716 ( n21836 , n1643 );
    and g15717 ( n38483 , n40584 , n37036 );
    or g15718 ( n30551 , n28111 , n20757 );
    xnor g15719 ( n11304 , n6625 , n33910 );
    and g15720 ( n40146 , n27670 , n36542 );
    or g15721 ( n26368 , n28114 , n12532 );
    or g15722 ( n15534 , n41314 , n29382 );
    or g15723 ( n7669 , n38175 , n37857 );
    xnor g15724 ( n34768 , n15706 , n37380 );
    or g15725 ( n28794 , n29992 , n10177 );
    or g15726 ( n7099 , n7336 , n25282 );
    nor g15727 ( n41254 , n41303 , n33956 );
    xnor g15728 ( n19833 , n36009 , n23974 );
    or g15729 ( n5241 , n21691 , n41981 );
    not g15730 ( n25303 , n27010 );
    and g15731 ( n10521 , n11894 , n19722 );
    or g15732 ( n27460 , n8966 , n22971 );
    xnor g15733 ( n26569 , n28303 , n32066 );
    nor g15734 ( n21210 , n38879 , n34998 );
    nor g15735 ( n16182 , n25348 , n7647 );
    or g15736 ( n20464 , n949 , n41880 );
    nor g15737 ( n39523 , n16619 , n9221 );
    nor g15738 ( n19815 , n40159 , n41610 );
    or g15739 ( n38628 , n27579 , n16250 );
    and g15740 ( n9725 , n27362 , n914 );
    and g15741 ( n25537 , n20181 , n382 );
    and g15742 ( n13448 , n41575 , n23810 );
    or g15743 ( n6276 , n38001 , n29980 );
    or g15744 ( n39269 , n5574 , n42713 );
    not g15745 ( n42738 , n31336 );
    and g15746 ( n28950 , n28974 , n9346 );
    or g15747 ( n10001 , n32116 , n33332 );
    not g15748 ( n23599 , n18683 );
    not g15749 ( n5546 , n18370 );
    or g15750 ( n13983 , n3782 , n27683 );
    xnor g15751 ( n18061 , n22899 , n34287 );
    and g15752 ( n3946 , n6217 , n9120 );
    or g15753 ( n6640 , n35534 , n25069 );
    and g15754 ( n10351 , n29408 , n2944 );
    and g15755 ( n11487 , n10765 , n8767 );
    or g15756 ( n22632 , n23599 , n22235 );
    nor g15757 ( n10477 , n18320 , n32683 );
    or g15758 ( n14849 , n9157 , n22892 );
    xnor g15759 ( n7401 , n14298 , n34160 );
    and g15760 ( n24380 , n38386 , n8057 );
    or g15761 ( n25599 , n15565 , n13587 );
    or g15762 ( n4263 , n37150 , n40556 );
    nor g15763 ( n10907 , n38762 , n18831 );
    or g15764 ( n12623 , n40462 , n4336 );
    not g15765 ( n14684 , n13037 );
    or g15766 ( n38844 , n19041 , n36856 );
    not g15767 ( n39139 , n25853 );
    nor g15768 ( n4286 , n41157 , n15232 );
    or g15769 ( n25685 , n36071 , n2237 );
    and g15770 ( n4990 , n25684 , n42463 );
    or g15771 ( n22166 , n3643 , n39328 );
    or g15772 ( n6887 , n40284 , n9563 );
    or g15773 ( n35420 , n259 , n12669 );
    and g15774 ( n35401 , n8719 , n11385 );
    not g15775 ( n8971 , n28595 );
    nor g15776 ( n2567 , n32408 , n26876 );
    or g15777 ( n20123 , n34267 , n12541 );
    nor g15778 ( n16209 , n15070 , n28571 );
    or g15779 ( n25971 , n10694 , n10646 );
    nor g15780 ( n38124 , n9743 , n18825 );
    not g15781 ( n34483 , n17454 );
    not g15782 ( n36815 , n20157 );
    and g15783 ( n32222 , n26190 , n31959 );
    not g15784 ( n18951 , n19667 );
    not g15785 ( n34278 , n18317 );
    or g15786 ( n13768 , n32326 , n41279 );
    or g15787 ( n27031 , n32471 , n20938 );
    not g15788 ( n14748 , n28474 );
    or g15789 ( n24220 , n37722 , n31153 );
    nor g15790 ( n29695 , n34565 , n5532 );
    not g15791 ( n19793 , n39246 );
    not g15792 ( n21184 , n41301 );
    and g15793 ( n3646 , n42030 , n33019 );
    xnor g15794 ( n25542 , n33253 , n7144 );
    and g15795 ( n2221 , n34402 , n35889 );
    and g15796 ( n32991 , n39684 , n6626 );
    and g15797 ( n35344 , n28410 , n12483 );
    or g15798 ( n13180 , n28468 , n32576 );
    or g15799 ( n25997 , n19811 , n12541 );
    or g15800 ( n35366 , n31190 , n37779 );
    and g15801 ( n21931 , n19430 , n14543 );
    and g15802 ( n20924 , n23625 , n12132 );
    not g15803 ( n18317 , n15476 );
    xnor g15804 ( n31456 , n37074 , n18742 );
    or g15805 ( n31504 , n8621 , n3915 );
    xnor g15806 ( n6337 , n27091 , n2199 );
    or g15807 ( n17116 , n9932 , n18888 );
    not g15808 ( n11962 , n37489 );
    and g15809 ( n12303 , n35543 , n16535 );
    and g15810 ( n27803 , n33273 , n8316 );
    nor g15811 ( n9938 , n17399 , n678 );
    xnor g15812 ( n33742 , n621 , n19998 );
    and g15813 ( n21438 , n41659 , n38497 );
    and g15814 ( n15440 , n12510 , n22961 );
    not g15815 ( n26358 , n35025 );
    or g15816 ( n35066 , n2459 , n3781 );
    xnor g15817 ( n6982 , n38749 , n24340 );
    or g15818 ( n15162 , n35458 , n40566 );
    nor g15819 ( n12427 , n23045 , n24763 );
    or g15820 ( n4698 , n2407 , n42023 );
    nor g15821 ( n35349 , n14812 , n30522 );
    or g15822 ( n36409 , n28143 , n32224 );
    or g15823 ( n37958 , n14768 , n31948 );
    nor g15824 ( n36817 , n14614 , n38038 );
    and g15825 ( n35850 , n7067 , n36834 );
    and g15826 ( n38977 , n3505 , n42493 );
    not g15827 ( n28057 , n36521 );
    and g15828 ( n36457 , n1699 , n39793 );
    or g15829 ( n37080 , n734 , n33604 );
    or g15830 ( n22406 , n16598 , n21103 );
    or g15831 ( n37555 , n15006 , n36889 );
    or g15832 ( n20109 , n13642 , n23857 );
    and g15833 ( n25545 , n23090 , n10516 );
    or g15834 ( n7822 , n24396 , n32781 );
    and g15835 ( n19596 , n37920 , n33159 );
    and g15836 ( n38574 , n37087 , n24073 );
    or g15837 ( n7512 , n23855 , n23211 );
    and g15838 ( n3230 , n37102 , n18819 );
    nor g15839 ( n25154 , n2900 , n19868 );
    or g15840 ( n38094 , n18119 , n30930 );
    xnor g15841 ( n15038 , n37297 , n445 );
    or g15842 ( n25764 , n39266 , n3885 );
    nor g15843 ( n37111 , n35301 , n30867 );
    or g15844 ( n30532 , n2829 , n7393 );
    xnor g15845 ( n9360 , n6106 , n6537 );
    nor g15846 ( n21874 , n15070 , n19115 );
    nor g15847 ( n29609 , n22537 , n23097 );
    or g15848 ( n5236 , n2466 , n11500 );
    not g15849 ( n17890 , n12307 );
    or g15850 ( n29365 , n41998 , n13815 );
    not g15851 ( n7729 , n990 );
    or g15852 ( n12615 , n25733 , n36081 );
    and g15853 ( n11510 , n38643 , n23108 );
    or g15854 ( n2894 , n40485 , n9306 );
    or g15855 ( n21464 , n13194 , n31918 );
    or g15856 ( n39649 , n2199 , n30326 );
    or g15857 ( n24580 , n64 , n20084 );
    nor g15858 ( n28778 , n20039 , n41999 );
    or g15859 ( n19306 , n39420 , n13617 );
    and g15860 ( n22845 , n28899 , n26593 );
    or g15861 ( n34579 , n37249 , n12491 );
    or g15862 ( n5517 , n24245 , n32222 );
    not g15863 ( n35871 , n41623 );
    or g15864 ( n21521 , n40133 , n11026 );
    or g15865 ( n27218 , n5324 , n967 );
    nor g15866 ( n36663 , n22473 , n37947 );
    and g15867 ( n3009 , n31592 , n11441 );
    and g15868 ( n13401 , n35650 , n31512 );
    nor g15869 ( n36835 , n13181 , n30687 );
    or g15870 ( n41276 , n30490 , n18639 );
    xnor g15871 ( n4677 , n29740 , n36155 );
    xnor g15872 ( n4235 , n10834 , n26808 );
    or g15873 ( n17 , n27311 , n23946 );
    or g15874 ( n13856 , n9008 , n31966 );
    not g15875 ( n35615 , n3758 );
    xnor g15876 ( n3768 , n4235 , n15849 );
    or g15877 ( n22488 , n309 , n19734 );
    not g15878 ( n12959 , n15739 );
    or g15879 ( n10628 , n40785 , n25714 );
    nor g15880 ( n33323 , n28248 , n24003 );
    or g15881 ( n39798 , n28088 , n12426 );
    and g15882 ( n13700 , n669 , n27688 );
    or g15883 ( n20236 , n23859 , n25876 );
    and g15884 ( n30884 , n26701 , n36020 );
    not g15885 ( n7397 , n9778 );
    nor g15886 ( n24623 , n17193 , n7327 );
    not g15887 ( n26749 , n14042 );
    or g15888 ( n39657 , n29842 , n6024 );
    or g15889 ( n23157 , n18775 , n8550 );
    xnor g15890 ( n8204 , n35813 , n29542 );
    nor g15891 ( n34413 , n16598 , n32919 );
    or g15892 ( n28387 , n10597 , n11467 );
    nor g15893 ( n9919 , n4914 , n34453 );
    nor g15894 ( n40796 , n16649 , n3714 );
    or g15895 ( n390 , n32026 , n23366 );
    nor g15896 ( n626 , n1110 , n4946 );
    xnor g15897 ( n20353 , n12190 , n20594 );
    and g15898 ( n28372 , n23784 , n3933 );
    nor g15899 ( n40534 , n12370 , n3115 );
    or g15900 ( n18670 , n3337 , n19714 );
    or g15901 ( n26805 , n675 , n28723 );
    nor g15902 ( n38042 , n24200 , n35856 );
    not g15903 ( n1674 , n31391 );
    and g15904 ( n23884 , n475 , n22205 );
    or g15905 ( n3672 , n13885 , n17273 );
    xnor g15906 ( n5481 , n18600 , n6058 );
    or g15907 ( n38270 , n24400 , n2647 );
    xnor g15908 ( n27576 , n7489 , n31114 );
    and g15909 ( n40676 , n21984 , n29410 );
    not g15910 ( n32105 , n7824 );
    and g15911 ( n17356 , n2744 , n6857 );
    and g15912 ( n22957 , n23919 , n36556 );
    xnor g15913 ( n10564 , n7922 , n31254 );
    nor g15914 ( n17869 , n16598 , n39746 );
    and g15915 ( n21912 , n1521 , n37448 );
    nor g15916 ( n15957 , n25781 , n2448 );
    or g15917 ( n38498 , n19068 , n13687 );
    not g15918 ( n1683 , n13714 );
    or g15919 ( n19872 , n1772 , n313 );
    xnor g15920 ( n40513 , n36009 , n15255 );
    or g15921 ( n3204 , n3387 , n2341 );
    or g15922 ( n1521 , n22505 , n769 );
    and g15923 ( n39131 , n6185 , n42291 );
    or g15924 ( n17582 , n12115 , n17888 );
    nor g15925 ( n42660 , n29362 , n32013 );
    nor g15926 ( n17485 , n33222 , n30613 );
    nor g15927 ( n18535 , n18754 , n26742 );
    or g15928 ( n17775 , n23060 , n41661 );
    or g15929 ( n1771 , n10193 , n27221 );
    or g15930 ( n3195 , n14945 , n19919 );
    not g15931 ( n36213 , n16395 );
    and g15932 ( n4101 , n3199 , n33119 );
    nor g15933 ( n9243 , n35009 , n12375 );
    and g15934 ( n34100 , n10757 , n2004 );
    not g15935 ( n36151 , n4574 );
    nor g15936 ( n28122 , n15648 , n2871 );
    and g15937 ( n5440 , n973 , n21489 );
    not g15938 ( n18199 , n25679 );
    and g15939 ( n39355 , n26064 , n23409 );
    or g15940 ( n8814 , n27941 , n4947 );
    or g15941 ( n1929 , n41203 , n12823 );
    and g15942 ( n40036 , n41421 , n29935 );
    and g15943 ( n5216 , n8174 , n29785 );
    not g15944 ( n27834 , n3900 );
    nor g15945 ( n28456 , n42050 , n4438 );
    and g15946 ( n8780 , n7545 , n4009 );
    and g15947 ( n33883 , n33734 , n25457 );
    or g15948 ( n41663 , n16007 , n4669 );
    and g15949 ( n3372 , n6727 , n34613 );
    or g15950 ( n33936 , n12653 , n10253 );
    not g15951 ( n20932 , n33843 );
    or g15952 ( n7940 , n21475 , n3036 );
    nor g15953 ( n13393 , n4266 , n855 );
    or g15954 ( n40142 , n34762 , n12523 );
    or g15955 ( n21657 , n13801 , n20145 );
    or g15956 ( n23104 , n21025 , n35339 );
    not g15957 ( n23497 , n31699 );
    or g15958 ( n25769 , n33216 , n30625 );
    and g15959 ( n27643 , n19740 , n8312 );
    xnor g15960 ( n32321 , n25889 , n16539 );
    or g15961 ( n36530 , n37455 , n42682 );
    or g15962 ( n15251 , n19770 , n15230 );
    nor g15963 ( n42428 , n35361 , n34406 );
    and g15964 ( n6589 , n8692 , n13663 );
    or g15965 ( n33374 , n1993 , n34652 );
    and g15966 ( n14492 , n15489 , n37931 );
    or g15967 ( n6191 , n10822 , n25127 );
    or g15968 ( n5067 , n30141 , n12129 );
    and g15969 ( n31238 , n960 , n11690 );
    or g15970 ( n20976 , n35340 , n21045 );
    or g15971 ( n4067 , n8494 , n37856 );
    or g15972 ( n27647 , n23472 , n30613 );
    xnor g15973 ( n7892 , n42064 , n10861 );
    or g15974 ( n13849 , n3660 , n22287 );
    not g15975 ( n6278 , n38080 );
    or g15976 ( n25757 , n19631 , n22105 );
    and g15977 ( n5539 , n9841 , n42294 );
    nor g15978 ( n37199 , n12639 , n18675 );
    and g15979 ( n9514 , n31219 , n10695 );
    or g15980 ( n16056 , n31794 , n32487 );
    not g15981 ( n10834 , n12651 );
    and g15982 ( n6613 , n7308 , n24600 );
    or g15983 ( n9115 , n34565 , n4510 );
    nor g15984 ( n29215 , n36088 , n14305 );
    or g15985 ( n40381 , n21096 , n19931 );
    and g15986 ( n23584 , n29494 , n20579 );
    not g15987 ( n23990 , n32597 );
    xnor g15988 ( n19760 , n36009 , n21357 );
    xnor g15989 ( n10399 , n13151 , n31727 );
    xnor g15990 ( n37448 , n37083 , n7349 );
    or g15991 ( n37904 , n30882 , n40702 );
    not g15992 ( n560 , n27654 );
    xnor g15993 ( n4073 , n29323 , n6886 );
    or g15994 ( n8300 , n30 , n1712 );
    or g15995 ( n11228 , n20684 , n12047 );
    xnor g15996 ( n23231 , n11595 , n35739 );
    not g15997 ( n19353 , n7548 );
    nor g15998 ( n9771 , n26627 , n17975 );
    and g15999 ( n16836 , n7068 , n16118 );
    or g16000 ( n29230 , n34762 , n41233 );
    or g16001 ( n22392 , n38479 , n36616 );
    or g16002 ( n28328 , n30131 , n8491 );
    not g16003 ( n41426 , n10847 );
    or g16004 ( n17618 , n23082 , n22480 );
    or g16005 ( n39498 , n42461 , n8156 );
    or g16006 ( n19821 , n42678 , n6832 );
    xnor g16007 ( n3702 , n5413 , n39616 );
    or g16008 ( n41800 , n5256 , n40787 );
    or g16009 ( n35870 , n18961 , n6004 );
    xnor g16010 ( n155 , n17561 , n41226 );
    or g16011 ( n37845 , n13801 , n30435 );
    nor g16012 ( n12053 , n2199 , n39949 );
    not g16013 ( n19260 , n17880 );
    and g16014 ( n39166 , n128 , n17298 );
    not g16015 ( n22039 , n15773 );
    or g16016 ( n7060 , n6827 , n8101 );
    xnor g16017 ( n20946 , n26579 , n38008 );
    or g16018 ( n37338 , n4535 , n14856 );
    or g16019 ( n4953 , n6423 , n35180 );
    or g16020 ( n21340 , n22667 , n10331 );
    xnor g16021 ( n36509 , n40090 , n10603 );
    or g16022 ( n30409 , n41474 , n11183 );
    or g16023 ( n24525 , n24062 , n18482 );
    or g16024 ( n42586 , n6370 , n20330 );
    nor g16025 ( n28881 , n34565 , n33539 );
    not g16026 ( n19463 , n25247 );
    or g16027 ( n38375 , n37603 , n35024 );
    xnor g16028 ( n27101 , n26897 , n14471 );
    and g16029 ( n30080 , n10356 , n16908 );
    and g16030 ( n23450 , n15962 , n15798 );
    or g16031 ( n33442 , n11325 , n31333 );
    and g16032 ( n11163 , n5040 , n18539 );
    and g16033 ( n29060 , n2207 , n25739 );
    xnor g16034 ( n10922 , n20972 , n37425 );
    or g16035 ( n3395 , n30110 , n35304 );
    and g16036 ( n38615 , n33055 , n1539 );
    and g16037 ( n28583 , n20386 , n36402 );
    and g16038 ( n34371 , n2595 , n13614 );
    not g16039 ( n5984 , n10307 );
    xnor g16040 ( n26299 , n18558 , n9399 );
    and g16041 ( n9047 , n13315 , n26365 );
    or g16042 ( n38434 , n12670 , n26789 );
    and g16043 ( n26119 , n41764 , n8929 );
    or g16044 ( n39290 , n20823 , n5316 );
    or g16045 ( n13192 , n18345 , n28865 );
    not g16046 ( n30984 , n8208 );
    or g16047 ( n18769 , n18798 , n17341 );
    not g16048 ( n41275 , n10482 );
    xnor g16049 ( n23237 , n31048 , n40539 );
    nor g16050 ( n15123 , n38073 , n6280 );
    or g16051 ( n7462 , n33010 , n13176 );
    not g16052 ( n21064 , n31825 );
    and g16053 ( n36399 , n1330 , n36615 );
    or g16054 ( n37910 , n37148 , n24220 );
    or g16055 ( n28873 , n14549 , n4159 );
    not g16056 ( n27913 , n703 );
    not g16057 ( n20492 , n5563 );
    and g16058 ( n37836 , n34857 , n34078 );
    or g16059 ( n26506 , n23812 , n23349 );
    and g16060 ( n3770 , n30861 , n11650 );
    and g16061 ( n23634 , n33060 , n1055 );
    and g16062 ( n10724 , n39042 , n8979 );
    or g16063 ( n9420 , n35208 , n33576 );
    nor g16064 ( n9730 , n10251 , n16857 );
    not g16065 ( n33592 , n28316 );
    and g16066 ( n779 , n2336 , n2058 );
    nor g16067 ( n8024 , n38879 , n40504 );
    not g16068 ( n5419 , n34274 );
    and g16069 ( n21819 , n5957 , n20465 );
    xnor g16070 ( n35910 , n39143 , n3843 );
    and g16071 ( n6220 , n25092 , n14582 );
    nor g16072 ( n37990 , n23478 , n27803 );
    nor g16073 ( n11259 , n9200 , n9982 );
    xnor g16074 ( n33122 , n20946 , n16527 );
    or g16075 ( n41563 , n3586 , n17979 );
    or g16076 ( n40189 , n21795 , n21187 );
    xnor g16077 ( n34086 , n12734 , n10330 );
    or g16078 ( n32469 , n39332 , n19160 );
    or g16079 ( n30905 , n7114 , n28818 );
    and g16080 ( n16562 , n16774 , n34113 );
    or g16081 ( n32620 , n22279 , n11716 );
    or g16082 ( n35097 , n40253 , n34004 );
    or g16083 ( n30577 , n33585 , n12741 );
    nor g16084 ( n33834 , n5099 , n7483 );
    or g16085 ( n34919 , n6796 , n22067 );
    or g16086 ( n16188 , n17108 , n30938 );
    nor g16087 ( n2688 , n21751 , n41449 );
    and g16088 ( n15433 , n25588 , n17706 );
    not g16089 ( n38242 , n38991 );
    not g16090 ( n28553 , n21155 );
    and g16091 ( n24815 , n22328 , n11315 );
    or g16092 ( n27668 , n3566 , n34290 );
    or g16093 ( n29226 , n15329 , n25216 );
    or g16094 ( n23404 , n22440 , n41145 );
    or g16095 ( n30468 , n31845 , n23676 );
    or g16096 ( n40788 , n34997 , n25300 );
    xnor g16097 ( n7080 , n42127 , n27468 );
    or g16098 ( n22780 , n6956 , n12636 );
    or g16099 ( n18246 , n28911 , n27333 );
    or g16100 ( n38236 , n31836 , n39002 );
    or g16101 ( n35987 , n9097 , n33168 );
    or g16102 ( n31237 , n8399 , n26927 );
    xnor g16103 ( n23135 , n6621 , n34004 );
    and g16104 ( n5986 , n1076 , n618 );
    or g16105 ( n6339 , n40380 , n16999 );
    or g16106 ( n3039 , n3080 , n15253 );
    xnor g16107 ( n16127 , n7840 , n13665 );
    xnor g16108 ( n4442 , n42064 , n14608 );
    not g16109 ( n33416 , n2919 );
    or g16110 ( n35162 , n28424 , n2364 );
    not g16111 ( n38918 , n42842 );
    and g16112 ( n41723 , n38244 , n40644 );
    xnor g16113 ( n20994 , n30429 , n18976 );
    or g16114 ( n5207 , n14551 , n17104 );
    nor g16115 ( n13571 , n23510 , n40170 );
    and g16116 ( n8816 , n3129 , n19105 );
    or g16117 ( n30923 , n9126 , n4043 );
    or g16118 ( n13242 , n37055 , n28320 );
    or g16119 ( n37531 , n22807 , n39609 );
    not g16120 ( n37388 , n28761 );
    not g16121 ( n17011 , n27881 );
    or g16122 ( n21577 , n5121 , n18716 );
    nor g16123 ( n13064 , n33981 , n12298 );
    or g16124 ( n27029 , n34565 , n42144 );
    or g16125 ( n41899 , n38773 , n27272 );
    nor g16126 ( n32298 , n12176 , n22205 );
    or g16127 ( n22646 , n15934 , n33476 );
    nor g16128 ( n740 , n38494 , n9543 );
    not g16129 ( n29437 , n30675 );
    and g16130 ( n30626 , n2523 , n42166 );
    not g16131 ( n9482 , n25005 );
    and g16132 ( n7971 , n26700 , n38714 );
    and g16133 ( n30344 , n12026 , n39169 );
    and g16134 ( n3709 , n20079 , n36159 );
    not g16135 ( n22173 , n4709 );
    or g16136 ( n41175 , n35386 , n27976 );
    or g16137 ( n11569 , n5754 , n1223 );
    or g16138 ( n35796 , n28741 , n40386 );
    and g16139 ( n12668 , n3294 , n30342 );
    not g16140 ( n38996 , n4756 );
    or g16141 ( n38850 , n42893 , n24092 );
    or g16142 ( n25872 , n25721 , n8372 );
    or g16143 ( n20695 , n32539 , n3630 );
    xnor g16144 ( n16658 , n18382 , n25805 );
    or g16145 ( n21594 , n35768 , n30208 );
    or g16146 ( n37133 , n2315 , n5012 );
    xnor g16147 ( n12631 , n36529 , n25463 );
    or g16148 ( n30900 , n14048 , n40388 );
    or g16149 ( n29302 , n19092 , n20900 );
    or g16150 ( n40932 , n29268 , n21220 );
    or g16151 ( n32054 , n22492 , n770 );
    or g16152 ( n37393 , n1091 , n42424 );
    nor g16153 ( n35072 , n16598 , n9574 );
    or g16154 ( n39453 , n32971 , n24053 );
    xnor g16155 ( n12772 , n5203 , n32215 );
    xnor g16156 ( n33919 , n37163 , n17442 );
    and g16157 ( n14677 , n32005 , n31031 );
    and g16158 ( n31964 , n37543 , n15466 );
    not g16159 ( n37653 , n20131 );
    or g16160 ( n29007 , n22050 , n22872 );
    or g16161 ( n3923 , n29058 , n3736 );
    and g16162 ( n19802 , n39931 , n23207 );
    not g16163 ( n14461 , n11922 );
    or g16164 ( n19302 , n20674 , n7406 );
    nor g16165 ( n26693 , n30295 , n37072 );
    or g16166 ( n592 , n552 , n16216 );
    or g16167 ( n24338 , n14707 , n25121 );
    or g16168 ( n13636 , n6705 , n15616 );
    or g16169 ( n25786 , n20728 , n36101 );
    and g16170 ( n23807 , n11263 , n2023 );
    or g16171 ( n31039 , n24656 , n29355 );
    or g16172 ( n8849 , n16719 , n16298 );
    not g16173 ( n10498 , n42164 );
    not g16174 ( n33652 , n32814 );
    or g16175 ( n36097 , n30812 , n38196 );
    not g16176 ( n6072 , n36681 );
    or g16177 ( n35703 , n12768 , n16102 );
    xnor g16178 ( n5985 , n1110 , n38043 );
    not g16179 ( n7342 , n38504 );
    xnor g16180 ( n34296 , n29758 , n1437 );
    and g16181 ( n5113 , n25071 , n30300 );
    xnor g16182 ( n3486 , n11168 , n17258 );
    and g16183 ( n27327 , n28100 , n8921 );
    or g16184 ( n4031 , n19982 , n28197 );
    or g16185 ( n17369 , n37771 , n37909 );
    and g16186 ( n1160 , n11276 , n26153 );
    or g16187 ( n41077 , n4541 , n36380 );
    not g16188 ( n25155 , n3635 );
    xnor g16189 ( n32782 , n4864 , n17655 );
    and g16190 ( n9424 , n17497 , n2109 );
    xnor g16191 ( n9138 , n18859 , n11068 );
    or g16192 ( n28270 , n17984 , n4866 );
    xnor g16193 ( n10335 , n8439 , n6716 );
    or g16194 ( n7902 , n35386 , n6662 );
    not g16195 ( n32350 , n11787 );
    or g16196 ( n15838 , n10963 , n30531 );
    not g16197 ( n6549 , n35930 );
    or g16198 ( n6678 , n5795 , n16787 );
    and g16199 ( n22325 , n11542 , n33608 );
    and g16200 ( n35948 , n36846 , n29933 );
    not g16201 ( n13481 , n13237 );
    xnor g16202 ( n32862 , n25042 , n31806 );
    and g16203 ( n20031 , n15626 , n39514 );
    xnor g16204 ( n3879 , n35509 , n2592 );
    or g16205 ( n3202 , n11039 , n39807 );
    xnor g16206 ( n31929 , n41013 , n37817 );
    or g16207 ( n5630 , n11331 , n25785 );
    nor g16208 ( n39975 , n14471 , n24369 );
    and g16209 ( n11779 , n33442 , n33642 );
    xnor g16210 ( n30571 , n4491 , n22957 );
    or g16211 ( n37596 , n5770 , n33926 );
    or g16212 ( n13287 , n42418 , n29299 );
    not g16213 ( n26624 , n23569 );
    not g16214 ( n35587 , n3278 );
    or g16215 ( n41945 , n24121 , n32978 );
    xnor g16216 ( n6997 , n1965 , n41386 );
    or g16217 ( n16907 , n14112 , n38819 );
    or g16218 ( n36670 , n39439 , n2835 );
    not g16219 ( n3713 , n10614 );
    nor g16220 ( n6907 , n5896 , n41909 );
    or g16221 ( n26822 , n22333 , n35115 );
    or g16222 ( n10783 , n12278 , n406 );
    nor g16223 ( n2087 , n22572 , n38482 );
    not g16224 ( n6243 , n40985 );
    xnor g16225 ( n16651 , n25673 , n26546 );
    and g16226 ( n17611 , n28866 , n23404 );
    not g16227 ( n7572 , n15166 );
    not g16228 ( n33620 , n6699 );
    nor g16229 ( n33485 , n14471 , n20341 );
    not g16230 ( n13249 , n27784 );
    and g16231 ( n36219 , n35114 , n3121 );
    not g16232 ( n31918 , n29777 );
    or g16233 ( n21089 , n37902 , n39635 );
    and g16234 ( n16955 , n14869 , n18048 );
    not g16235 ( n41684 , n2320 );
    and g16236 ( n18634 , n39450 , n41886 );
    or g16237 ( n22360 , n26569 , n18393 );
    or g16238 ( n7241 , n16996 , n38102 );
    or g16239 ( n34716 , n40429 , n8035 );
    nor g16240 ( n6315 , n18209 , n26716 );
    or g16241 ( n483 , n11349 , n2964 );
    and g16242 ( n23081 , n13567 , n8597 );
    or g16243 ( n11352 , n13556 , n16174 );
    and g16244 ( n23602 , n5557 , n24543 );
    not g16245 ( n500 , n41147 );
    nor g16246 ( n9677 , n7203 , n4483 );
    not g16247 ( n12768 , n7069 );
    xnor g16248 ( n31293 , n26579 , n39505 );
    not g16249 ( n42258 , n5248 );
    xnor g16250 ( n15588 , n33324 , n39658 );
    or g16251 ( n33647 , n25777 , n26539 );
    or g16252 ( n42325 , n14370 , n41258 );
    or g16253 ( n40650 , n9951 , n16990 );
    or g16254 ( n4075 , n27175 , n3868 );
    and g16255 ( n35761 , n30960 , n35601 );
    not g16256 ( n15402 , n5792 );
    not g16257 ( n36938 , n4746 );
    and g16258 ( n29588 , n29901 , n4526 );
    not g16259 ( n31332 , n20448 );
    and g16260 ( n27578 , n25057 , n35434 );
    and g16261 ( n25005 , n28878 , n7382 );
    or g16262 ( n15839 , n27999 , n35852 );
    and g16263 ( n39378 , n41554 , n16854 );
    and g16264 ( n13419 , n41390 , n10896 );
    not g16265 ( n18021 , n38758 );
    nor g16266 ( n36837 , n37868 , n27645 );
    xnor g16267 ( n1845 , n42064 , n12560 );
    or g16268 ( n20028 , n3162 , n40415 );
    and g16269 ( n7893 , n19886 , n16453 );
    xnor g16270 ( n20448 , n25694 , n38879 );
    and g16271 ( n42017 , n14628 , n22214 );
    or g16272 ( n15592 , n16725 , n30846 );
    nor g16273 ( n9472 , n20368 , n10034 );
    and g16274 ( n2549 , n21932 , n26511 );
    not g16275 ( n17131 , n9774 );
    xnor g16276 ( n32516 , n24216 , n9867 );
    not g16277 ( n25210 , n29356 );
    and g16278 ( n40088 , n3019 , n21148 );
    and g16279 ( n14623 , n33138 , n1259 );
    xnor g16280 ( n25766 , n33570 , n16311 );
    not g16281 ( n8380 , n21714 );
    or g16282 ( n3208 , n39266 , n190 );
    not g16283 ( n35167 , n5406 );
    xnor g16284 ( n3147 , n23325 , n27823 );
    xnor g16285 ( n38364 , n14596 , n37015 );
    or g16286 ( n5946 , n197 , n42525 );
    or g16287 ( n42605 , n30051 , n36296 );
    or g16288 ( n17895 , n405 , n22469 );
    or g16289 ( n14698 , n29135 , n2102 );
    and g16290 ( n40896 , n25097 , n3397 );
    xnor g16291 ( n15411 , n16455 , n38157 );
    or g16292 ( n6606 , n30161 , n33030 );
    xnor g16293 ( n6061 , n34844 , n24765 );
    nor g16294 ( n31499 , n25588 , n22998 );
    or g16295 ( n21986 , n16172 , n24783 );
    or g16296 ( n307 , n8670 , n23559 );
    not g16297 ( n42550 , n35391 );
    or g16298 ( n26125 , n25280 , n16216 );
    and g16299 ( n24143 , n2094 , n13776 );
    nor g16300 ( n11143 , n32033 , n17408 );
    or g16301 ( n3995 , n4798 , n4590 );
    not g16302 ( n36807 , n10867 );
    or g16303 ( n13761 , n29027 , n33653 );
    or g16304 ( n1052 , n22447 , n24451 );
    and g16305 ( n22172 , n36961 , n33069 );
    or g16306 ( n3846 , n981 , n22246 );
    and g16307 ( n36977 , n10956 , n12461 );
    not g16308 ( n25173 , n8649 );
    and g16309 ( n3246 , n13806 , n14469 );
    or g16310 ( n37483 , n42631 , n17827 );
    not g16311 ( n24408 , n6551 );
    xnor g16312 ( n12386 , n8502 , n14378 );
    not g16313 ( n30801 , n14241 );
    or g16314 ( n23950 , n39489 , n39570 );
    nor g16315 ( n7601 , n7344 , n20008 );
    and g16316 ( n5036 , n23546 , n3774 );
    not g16317 ( n26922 , n6032 );
    and g16318 ( n19688 , n29967 , n28768 );
    not g16319 ( n41207 , n1793 );
    and g16320 ( n25361 , n42581 , n3832 );
    and g16321 ( n22090 , n30596 , n24158 );
    and g16322 ( n2684 , n33059 , n6447 );
    or g16323 ( n1022 , n36466 , n772 );
    not g16324 ( n30845 , n22134 );
    nor g16325 ( n20897 , n28884 , n4884 );
    not g16326 ( n8422 , n26836 );
    and g16327 ( n33410 , n37739 , n12357 );
    xnor g16328 ( n2994 , n9180 , n6144 );
    nor g16329 ( n22719 , n30593 , n40185 );
    and g16330 ( n2761 , n23119 , n1614 );
    nor g16331 ( n34407 , n32544 , n9956 );
    xnor g16332 ( n17958 , n22263 , n32089 );
    not g16333 ( n42609 , n2523 );
    or g16334 ( n515 , n17297 , n30896 );
    or g16335 ( n23464 , n20122 , n22017 );
    nor g16336 ( n35151 , n15330 , n30388 );
    nor g16337 ( n12879 , n34852 , n23159 );
    and g16338 ( n1100 , n36074 , n12534 );
    not g16339 ( n40698 , n32118 );
    nor g16340 ( n10955 , n39645 , n28625 );
    and g16341 ( n42492 , n6355 , n15286 );
    xnor g16342 ( n3929 , n784 , n36522 );
    or g16343 ( n24249 , n12215 , n6389 );
    nor g16344 ( n11767 , n16780 , n23342 );
    or g16345 ( n39989 , n15890 , n3271 );
    and g16346 ( n28836 , n21459 , n40673 );
    and g16347 ( n29097 , n3723 , n40273 );
    or g16348 ( n32767 , n28745 , n9556 );
    or g16349 ( n2796 , n39589 , n33230 );
    nor g16350 ( n42205 , n1209 , n26525 );
    or g16351 ( n31438 , n34250 , n28556 );
    or g16352 ( n40009 , n37445 , n1729 );
    or g16353 ( n36523 , n14707 , n41888 );
    or g16354 ( n32976 , n425 , n16832 );
    xnor g16355 ( n17089 , n784 , n34863 );
    or g16356 ( n20523 , n2315 , n10772 );
    xnor g16357 ( n33441 , n10822 , n2104 );
    or g16358 ( n10813 , n15792 , n10532 );
    or g16359 ( n10636 , n38704 , n26868 );
    or g16360 ( n37997 , n4101 , n12210 );
    and g16361 ( n35708 , n12895 , n40433 );
    or g16362 ( n12108 , n3230 , n13368 );
    and g16363 ( n11896 , n24861 , n36109 );
    and g16364 ( n28678 , n31989 , n21726 );
    or g16365 ( n34508 , n30694 , n11901 );
    and g16366 ( n19517 , n8480 , n27890 );
    not g16367 ( n30350 , n29453 );
    or g16368 ( n19704 , n39954 , n23955 );
    or g16369 ( n16334 , n34292 , n41448 );
    or g16370 ( n20455 , n39023 , n41532 );
    or g16371 ( n13221 , n17888 , n27002 );
    or g16372 ( n16596 , n36946 , n20141 );
    or g16373 ( n36085 , n29082 , n6358 );
    and g16374 ( n17943 , n4903 , n2158 );
    xnor g16375 ( n17007 , n378 , n23354 );
    or g16376 ( n33559 , n28537 , n16119 );
    not g16377 ( n28461 , n9652 );
    not g16378 ( n10211 , n11546 );
    xnor g16379 ( n7962 , n13609 , n32755 );
    or g16380 ( n20838 , n19536 , n37058 );
    or g16381 ( n9117 , n19278 , n12498 );
    and g16382 ( n42385 , n17590 , n15597 );
    and g16383 ( n20853 , n35762 , n16884 );
    nor g16384 ( n14412 , n785 , n21546 );
    or g16385 ( n14995 , n24638 , n33469 );
    or g16386 ( n32442 , n37666 , n29232 );
    nor g16387 ( n24897 , n4141 , n8783 );
    or g16388 ( n38370 , n15703 , n21266 );
    xnor g16389 ( n14479 , n14070 , n12002 );
    and g16390 ( n5504 , n41826 , n40002 );
    or g16391 ( n21638 , n42454 , n20599 );
    and g16392 ( n16687 , n2241 , n4415 );
    and g16393 ( n38492 , n5436 , n25998 );
    or g16394 ( n39004 , n27037 , n25981 );
    xnor g16395 ( n142 , n21654 , n12449 );
    nor g16396 ( n22363 , n29303 , n27998 );
    nor g16397 ( n26886 , n29858 , n38748 );
    and g16398 ( n39373 , n18904 , n37474 );
    and g16399 ( n8010 , n35817 , n37355 );
    nor g16400 ( n18263 , n22175 , n31211 );
    or g16401 ( n14310 , n36067 , n42776 );
    xnor g16402 ( n23008 , n36587 , n36117 );
    and g16403 ( n6009 , n39534 , n30556 );
    not g16404 ( n36641 , n8422 );
    or g16405 ( n23943 , n5718 , n33281 );
    and g16406 ( n29937 , n17821 , n16389 );
    or g16407 ( n27794 , n9539 , n35890 );
    or g16408 ( n24821 , n6686 , n11278 );
    not g16409 ( n42765 , n5815 );
    or g16410 ( n25439 , n19808 , n10385 );
    xnor g16411 ( n37284 , n36009 , n14238 );
    or g16412 ( n35325 , n6566 , n11906 );
    or g16413 ( n17846 , n5704 , n12000 );
    nor g16414 ( n12547 , n1003 , n8431 );
    and g16415 ( n2379 , n16477 , n14693 );
    not g16416 ( n10904 , n16168 );
    nor g16417 ( n13970 , n1868 , n19019 );
    and g16418 ( n17643 , n737 , n28739 );
    and g16419 ( n35528 , n40406 , n4054 );
    and g16420 ( n15960 , n36777 , n29722 );
    or g16421 ( n15702 , n33708 , n22699 );
    not g16422 ( n13430 , n41595 );
    nor g16423 ( n11065 , n3934 , n7065 );
    and g16424 ( n30414 , n13585 , n31182 );
    xnor g16425 ( n5159 , n1841 , n40668 );
    not g16426 ( n5219 , n37296 );
    or g16427 ( n18970 , n16286 , n21466 );
    and g16428 ( n33082 , n28063 , n2940 );
    not g16429 ( n10974 , n37794 );
    xnor g16430 ( n36090 , n33902 , n1507 );
    or g16431 ( n9948 , n12378 , n21721 );
    nor g16432 ( n41653 , n12962 , n15831 );
    nor g16433 ( n9642 , n38163 , n18588 );
    and g16434 ( n4016 , n2603 , n20937 );
    not g16435 ( n38629 , n32667 );
    and g16436 ( n22134 , n14968 , n20615 );
    xnor g16437 ( n25676 , n12146 , n3874 );
    not g16438 ( n41515 , n5842 );
    or g16439 ( n4898 , n15064 , n39170 );
    or g16440 ( n34895 , n17231 , n24778 );
    not g16441 ( n1178 , n6065 );
    or g16442 ( n2189 , n16267 , n34829 );
    xnor g16443 ( n9981 , n27874 , n19036 );
    not g16444 ( n32094 , n3425 );
    nor g16445 ( n13116 , n8494 , n41783 );
    or g16446 ( n15814 , n34292 , n30412 );
    and g16447 ( n3882 , n10961 , n14527 );
    or g16448 ( n14573 , n35980 , n5077 );
    or g16449 ( n32739 , n24068 , n296 );
    not g16450 ( n21559 , n27895 );
    not g16451 ( n36848 , n36521 );
    or g16452 ( n13647 , n2087 , n1404 );
    nor g16453 ( n3245 , n2171 , n12877 );
    or g16454 ( n10741 , n24062 , n33272 );
    or g16455 ( n10862 , n7785 , n26815 );
    not g16456 ( n5340 , n39784 );
    not g16457 ( n41270 , n6230 );
    xnor g16458 ( n10927 , n36379 , n38879 );
    not g16459 ( n20817 , n4873 );
    not g16460 ( n267 , n18872 );
    or g16461 ( n2976 , n26166 , n39408 );
    and g16462 ( n2865 , n41815 , n16407 );
    xnor g16463 ( n19394 , n33458 , n34622 );
    or g16464 ( n1060 , n8539 , n35697 );
    not g16465 ( n28135 , n17189 );
    or g16466 ( n3572 , n9752 , n18973 );
    or g16467 ( n13442 , n25383 , n21215 );
    and g16468 ( n3357 , n23755 , n25542 );
    not g16469 ( n17079 , n18359 );
    xnor g16470 ( n2766 , n18231 , n2702 );
    or g16471 ( n21392 , n5896 , n788 );
    or g16472 ( n14767 , n28060 , n2518 );
    or g16473 ( n42224 , n33377 , n35745 );
    or g16474 ( n4485 , n1756 , n36694 );
    xnor g16475 ( n19339 , n17395 , n41083 );
    or g16476 ( n10893 , n16006 , n3715 );
    not g16477 ( n6784 , n28416 );
    or g16478 ( n6963 , n36111 , n19106 );
    or g16479 ( n7383 , n22892 , n39552 );
    or g16480 ( n42043 , n5280 , n19225 );
    xnor g16481 ( n41029 , n32874 , n1527 );
    and g16482 ( n39310 , n7799 , n5260 );
    and g16483 ( n23792 , n30091 , n22320 );
    or g16484 ( n37588 , n19469 , n2524 );
    nor g16485 ( n39980 , n19221 , n28547 );
    and g16486 ( n11087 , n11625 , n36769 );
    nor g16487 ( n12020 , n33796 , n10130 );
    xnor g16488 ( n42909 , n36146 , n36871 );
    or g16489 ( n6624 , n2387 , n20071 );
    or g16490 ( n33292 , n5581 , n16045 );
    or g16491 ( n23625 , n40090 , n2432 );
    or g16492 ( n20977 , n1110 , n34523 );
    and g16493 ( n26102 , n38920 , n11408 );
    and g16494 ( n8698 , n17248 , n40031 );
    or g16495 ( n4984 , n41545 , n11775 );
    or g16496 ( n39717 , n23502 , n39817 );
    not g16497 ( n9145 , n39392 );
    not g16498 ( n1806 , n29808 );
    or g16499 ( n23398 , n24234 , n40966 );
    not g16500 ( n3292 , n33551 );
    or g16501 ( n24213 , n34824 , n153 );
    or g16502 ( n7312 , n24547 , n11071 );
    or g16503 ( n31826 , n26542 , n11661 );
    or g16504 ( n26382 , n37688 , n42165 );
    nor g16505 ( n32985 , n21208 , n2721 );
    or g16506 ( n29207 , n10788 , n27663 );
    nor g16507 ( n36269 , n14471 , n41567 );
    not g16508 ( n10064 , n10000 );
    xnor g16509 ( n2523 , n21957 , n21143 );
    xnor g16510 ( n32465 , n85 , n29838 );
    or g16511 ( n16277 , n13866 , n16472 );
    xnor g16512 ( n41228 , n6014 , n20285 );
    and g16513 ( n26573 , n4268 , n6955 );
    or g16514 ( n12894 , n5161 , n35845 );
    or g16515 ( n1582 , n38935 , n5409 );
    and g16516 ( n37155 , n1563 , n16525 );
    not g16517 ( n41037 , n35620 );
    or g16518 ( n7597 , n4732 , n30451 );
    and g16519 ( n7498 , n30509 , n7345 );
    and g16520 ( n2525 , n21519 , n20649 );
    and g16521 ( n7543 , n30645 , n36392 );
    or g16522 ( n40900 , n41103 , n29930 );
    and g16523 ( n17788 , n13231 , n15872 );
    and g16524 ( n26017 , n9695 , n37718 );
    or g16525 ( n38764 , n36458 , n21064 );
    not g16526 ( n23444 , n38355 );
    not g16527 ( n38356 , n40725 );
    or g16528 ( n31799 , n38238 , n11374 );
    and g16529 ( n12975 , n4889 , n14960 );
    or g16530 ( n31295 , n25142 , n4505 );
    or g16531 ( n41282 , n17609 , n32774 );
    or g16532 ( n7913 , n32345 , n4595 );
    not g16533 ( n4567 , n24453 );
    or g16534 ( n28504 , n38530 , n29299 );
    nor g16535 ( n21730 , n37376 , n36397 );
    and g16536 ( n15950 , n5640 , n16888 );
    not g16537 ( n24998 , n26650 );
    and g16538 ( n33582 , n24502 , n10618 );
    nor g16539 ( n27501 , n19330 , n23987 );
    or g16540 ( n22094 , n27827 , n19196 );
    xnor g16541 ( n42761 , n11449 , n1817 );
    nor g16542 ( n372 , n37546 , n31599 );
    or g16543 ( n25713 , n15404 , n36033 );
    xnor g16544 ( n28597 , n2419 , n40144 );
    or g16545 ( n42019 , n26122 , n10758 );
    or g16546 ( n22395 , n9645 , n6512 );
    or g16547 ( n30333 , n31936 , n15950 );
    xnor g16548 ( n19949 , n6625 , n19802 );
    and g16549 ( n10916 , n10325 , n109 );
    xnor g16550 ( n3641 , n15911 , n22259 );
    nor g16551 ( n35338 , n7567 , n40999 );
    xnor g16552 ( n32734 , n39432 , n14680 );
    or g16553 ( n26881 , n39365 , n31303 );
    and g16554 ( n22909 , n12985 , n32198 );
    and g16555 ( n42458 , n31159 , n35230 );
    not g16556 ( n28500 , n23353 );
    nor g16557 ( n13466 , n13046 , n37234 );
    nor g16558 ( n10137 , n30539 , n14938 );
    and g16559 ( n25750 , n34731 , n41039 );
    and g16560 ( n9054 , n30178 , n37470 );
    xnor g16561 ( n29956 , n2956 , n6492 );
    and g16562 ( n24566 , n23869 , n24748 );
    xnor g16563 ( n24627 , n15309 , n17811 );
    not g16564 ( n19807 , n27815 );
    and g16565 ( n32977 , n38190 , n22382 );
    xnor g16566 ( n7541 , n29272 , n15321 );
    or g16567 ( n22570 , n26147 , n25182 );
    xnor g16568 ( n8193 , n28377 , n40270 );
    nor g16569 ( n22905 , n13340 , n16430 );
    or g16570 ( n17003 , n2807 , n10491 );
    or g16571 ( n1483 , n18916 , n39812 );
    or g16572 ( n9842 , n17684 , n4209 );
    or g16573 ( n7240 , n28723 , n32308 );
    or g16574 ( n6642 , n21373 , n7418 );
    not g16575 ( n14596 , n10962 );
    and g16576 ( n36524 , n23346 , n9762 );
    and g16577 ( n26594 , n34457 , n22236 );
    and g16578 ( n14730 , n38133 , n11137 );
    or g16579 ( n41529 , n30214 , n26559 );
    xnor g16580 ( n4232 , n41218 , n24973 );
    or g16581 ( n3058 , n11454 , n5586 );
    not g16582 ( n39712 , n23584 );
    and g16583 ( n29181 , n9716 , n30480 );
    and g16584 ( n30004 , n5508 , n3681 );
    and g16585 ( n2545 , n16024 , n18655 );
    and g16586 ( n41632 , n17039 , n42890 );
    not g16587 ( n14072 , n7627 );
    and g16588 ( n26854 , n12250 , n36248 );
    xnor g16589 ( n19380 , n31947 , n30632 );
    and g16590 ( n25460 , n33761 , n24768 );
    or g16591 ( n9769 , n12070 , n40485 );
    and g16592 ( n3586 , n35173 , n40061 );
    or g16593 ( n23712 , n11106 , n28754 );
    xnor g16594 ( n7887 , n28443 , n1857 );
    or g16595 ( n2849 , n12508 , n24116 );
    and g16596 ( n41227 , n6736 , n30202 );
    and g16597 ( n27735 , n11206 , n36543 );
    nor g16598 ( n26130 , n4228 , n12616 );
    or g16599 ( n32058 , n6393 , n14074 );
    not g16600 ( n25875 , n21503 );
    nor g16601 ( n30382 , n15447 , n1807 );
    or g16602 ( n30949 , n27760 , n33971 );
    xnor g16603 ( n39170 , n33512 , n36404 );
    or g16604 ( n11296 , n8556 , n26888 );
    and g16605 ( n4594 , n30726 , n29317 );
    xnor g16606 ( n14130 , n9429 , n31559 );
    and g16607 ( n30305 , n17148 , n27314 );
    and g16608 ( n699 , n27525 , n14850 );
    nor g16609 ( n9504 , n11460 , n41706 );
    not g16610 ( n15064 , n26245 );
    nor g16611 ( n14360 , n1046 , n5483 );
    or g16612 ( n19979 , n28757 , n9364 );
    or g16613 ( n30286 , n37032 , n4825 );
    xnor g16614 ( n26397 , n39150 , n27947 );
    or g16615 ( n5830 , n5964 , n41556 );
    not g16616 ( n31795 , n31088 );
    and g16617 ( n39884 , n15855 , n34765 );
    xnor g16618 ( n512 , n8210 , n11435 );
    not g16619 ( n41904 , n3044 );
    not g16620 ( n211 , n25326 );
    not g16621 ( n36063 , n20206 );
    or g16622 ( n10288 , n33541 , n80 );
    xnor g16623 ( n3339 , n7489 , n24606 );
    xnor g16624 ( n11586 , n17281 , n8936 );
    not g16625 ( n31074 , n8560 );
    and g16626 ( n8033 , n11448 , n16647 );
    not g16627 ( n27245 , n16253 );
    and g16628 ( n18762 , n23622 , n12506 );
    not g16629 ( n41891 , n17467 );
    or g16630 ( n38426 , n4219 , n19803 );
    nor g16631 ( n27208 , n40792 , n17420 );
    not g16632 ( n38747 , n36457 );
    xnor g16633 ( n19692 , n22263 , n23079 );
    or g16634 ( n38397 , n8088 , n5910 );
    or g16635 ( n23112 , n5173 , n19870 );
    or g16636 ( n8824 , n39016 , n36284 );
    or g16637 ( n10120 , n16593 , n10497 );
    or g16638 ( n20711 , n39210 , n12552 );
    or g16639 ( n4886 , n39204 , n7169 );
    xnor g16640 ( n21180 , n37383 , n18656 );
    or g16641 ( n1077 , n37917 , n26407 );
    or g16642 ( n40910 , n38586 , n27585 );
    and g16643 ( n15338 , n26579 , n12026 );
    or g16644 ( n8919 , n41227 , n7863 );
    and g16645 ( n293 , n38366 , n17557 );
    and g16646 ( n38120 , n9714 , n13321 );
    and g16647 ( n9680 , n4616 , n2324 );
    nor g16648 ( n30203 , n17393 , n30544 );
    or g16649 ( n40704 , n26782 , n2570 );
    xnor g16650 ( n42315 , n18880 , n15897 );
    or g16651 ( n8377 , n23201 , n23726 );
    not g16652 ( n42154 , n40078 );
    or g16653 ( n11162 , n42433 , n39879 );
    xnor g16654 ( n42552 , n7922 , n3240 );
    xnor g16655 ( n10394 , n2205 , n35708 );
    or g16656 ( n12060 , n18882 , n17229 );
    or g16657 ( n18284 , n12497 , n32568 );
    nor g16658 ( n25182 , n9525 , n17415 );
    not g16659 ( n22515 , n33133 );
    and g16660 ( n41304 , n35212 , n32138 );
    not g16661 ( n34551 , n6447 );
    not g16662 ( n26336 , n19171 );
    and g16663 ( n22447 , n24809 , n19555 );
    or g16664 ( n38941 , n8698 , n2647 );
    or g16665 ( n9498 , n40972 , n40160 );
    or g16666 ( n33909 , n26784 , n37060 );
    or g16667 ( n11944 , n41564 , n42247 );
    not g16668 ( n15149 , n22306 );
    not g16669 ( n38251 , n1879 );
    and g16670 ( n339 , n31653 , n37573 );
    xnor g16671 ( n3241 , n42064 , n35801 );
    or g16672 ( n35647 , n22493 , n32628 );
    or g16673 ( n15501 , n13043 , n26191 );
    or g16674 ( n6857 , n27761 , n33225 );
    or g16675 ( n17027 , n21863 , n10306 );
    and g16676 ( n36040 , n13497 , n18237 );
    or g16677 ( n12471 , n33691 , n8245 );
    and g16678 ( n88 , n10589 , n13971 );
    and g16679 ( n18123 , n24914 , n16939 );
    not g16680 ( n31859 , n28207 );
    and g16681 ( n34159 , n12039 , n32382 );
    nor g16682 ( n11202 , n30764 , n3240 );
    and g16683 ( n24708 , n30667 , n27256 );
    and g16684 ( n39716 , n22780 , n5925 );
    and g16685 ( n10075 , n27872 , n42858 );
    xnor g16686 ( n13891 , n16693 , n24581 );
    and g16687 ( n2328 , n3486 , n6450 );
    and g16688 ( n11024 , n21868 , n13729 );
    and g16689 ( n28370 , n2029 , n19642 );
    xnor g16690 ( n27706 , n25041 , n15271 );
    xnor g16691 ( n9995 , n1435 , n40190 );
    or g16692 ( n36963 , n6685 , n7152 );
    nor g16693 ( n12018 , n23920 , n38097 );
    and g16694 ( n25131 , n30765 , n39959 );
    and g16695 ( n40317 , n19851 , n3219 );
    not g16696 ( n1180 , n23060 );
    or g16697 ( n3390 , n14848 , n25451 );
    nor g16698 ( n31288 , n2751 , n13975 );
    and g16699 ( n3162 , n6354 , n22397 );
    or g16700 ( n6532 , n11694 , n8664 );
    or g16701 ( n39014 , n61 , n21807 );
    xnor g16702 ( n36200 , n31471 , n28361 );
    or g16703 ( n19150 , n32087 , n9265 );
    or g16704 ( n9826 , n7375 , n161 );
    not g16705 ( n37195 , n11456 );
    or g16706 ( n14495 , n5324 , n6505 );
    and g16707 ( n21234 , n34239 , n41383 );
    xnor g16708 ( n9931 , n4427 , n859 );
    not g16709 ( n26240 , n18363 );
    nor g16710 ( n8647 , n1507 , n5720 );
    or g16711 ( n19249 , n12722 , n29763 );
    or g16712 ( n35683 , n10598 , n24190 );
    and g16713 ( n17944 , n14727 , n14020 );
    nor g16714 ( n19673 , n19602 , n24475 );
    xnor g16715 ( n16010 , n34687 , n8778 );
    or g16716 ( n12163 , n39822 , n10584 );
    and g16717 ( n4432 , n5744 , n9280 );
    xnor g16718 ( n33421 , n21534 , n13750 );
    and g16719 ( n28748 , n9117 , n8063 );
    xnor g16720 ( n20511 , n10676 , n26228 );
    or g16721 ( n39918 , n7256 , n1735 );
    nor g16722 ( n1087 , n28490 , n25989 );
    not g16723 ( n13659 , n42159 );
    and g16724 ( n14235 , n3688 , n15533 );
    or g16725 ( n16829 , n24125 , n10485 );
    or g16726 ( n7434 , n3960 , n12797 );
    or g16727 ( n29202 , n11332 , n30998 );
    or g16728 ( n42406 , n35313 , n35490 );
    or g16729 ( n24358 , n34249 , n11456 );
    or g16730 ( n31942 , n22619 , n5628 );
    xnor g16731 ( n10835 , n4936 , n14707 );
    or g16732 ( n38488 , n7635 , n41207 );
    not g16733 ( n12125 , n14045 );
    not g16734 ( n14315 , n26268 );
    or g16735 ( n28033 , n28143 , n15277 );
    and g16736 ( n38331 , n32678 , n9726 );
    not g16737 ( n6065 , n42707 );
    or g16738 ( n41311 , n14466 , n11233 );
    or g16739 ( n5461 , n40995 , n11254 );
    or g16740 ( n1137 , n31027 , n9177 );
    and g16741 ( n26635 , n32270 , n34040 );
    or g16742 ( n15804 , n35790 , n21094 );
    and g16743 ( n19082 , n8268 , n29420 );
    nor g16744 ( n15200 , n14972 , n34120 );
    not g16745 ( n17796 , n25362 );
    not g16746 ( n10279 , n9116 );
    or g16747 ( n21435 , n40383 , n2476 );
    nor g16748 ( n11364 , n28945 , n26985 );
    and g16749 ( n16635 , n19580 , n2813 );
    or g16750 ( n26331 , n13555 , n5585 );
    or g16751 ( n6386 , n228 , n11312 );
    xnor g16752 ( n6476 , n32470 , n12683 );
    or g16753 ( n15229 , n23744 , n15780 );
    or g16754 ( n7684 , n39395 , n28134 );
    or g16755 ( n39202 , n8626 , n31776 );
    xnor g16756 ( n2806 , n27900 , n22727 );
    xnor g16757 ( n40061 , n34731 , n40175 );
    and g16758 ( n32172 , n24870 , n42658 );
    or g16759 ( n18605 , n13545 , n20846 );
    not g16760 ( n19089 , n38462 );
    or g16761 ( n40762 , n23826 , n18089 );
    nor g16762 ( n19190 , n18866 , n10816 );
    not g16763 ( n9051 , n41117 );
    not g16764 ( n21201 , n36661 );
    or g16765 ( n17592 , n38773 , n19265 );
    xnor g16766 ( n24994 , n4218 , n41897 );
    nor g16767 ( n23119 , n4183 , n21019 );
    or g16768 ( n42318 , n12792 , n27302 );
    or g16769 ( n11738 , n38816 , n20978 );
    xnor g16770 ( n36901 , n10376 , n26750 );
    or g16771 ( n15649 , n29214 , n15440 );
    and g16772 ( n32457 , n38046 , n38400 );
    nor g16773 ( n21953 , n39962 , n2277 );
    and g16774 ( n15009 , n17520 , n34157 );
    not g16775 ( n42481 , n19281 );
    not g16776 ( n36214 , n21114 );
    xnor g16777 ( n28336 , n34822 , n9497 );
    nor g16778 ( n37917 , n4681 , n14229 );
    nor g16779 ( n31195 , n23883 , n38506 );
    or g16780 ( n541 , n33907 , n17393 );
    or g16781 ( n31743 , n25407 , n18068 );
    and g16782 ( n2901 , n31537 , n40054 );
    or g16783 ( n34871 , n36117 , n7453 );
    not g16784 ( n40541 , n23269 );
    and g16785 ( n8661 , n36684 , n28355 );
    or g16786 ( n33550 , n19731 , n4781 );
    not g16787 ( n15389 , n26999 );
    or g16788 ( n18630 , n38763 , n34184 );
    or g16789 ( n33280 , n30790 , n38856 );
    or g16790 ( n28640 , n15698 , n10053 );
    not g16791 ( n136 , n38661 );
    xnor g16792 ( n30297 , n2174 , n24993 );
    or g16793 ( n5535 , n41373 , n15317 );
    and g16794 ( n42755 , n41852 , n2325 );
    and g16795 ( n13325 , n18168 , n15322 );
    not g16796 ( n14503 , n32905 );
    xnor g16797 ( n38589 , n892 , n10126 );
    or g16798 ( n26411 , n1396 , n25664 );
    or g16799 ( n5871 , n8512 , n41414 );
    or g16800 ( n36867 , n11294 , n18955 );
    or g16801 ( n24381 , n40374 , n28971 );
    nor g16802 ( n9426 , n8204 , n30732 );
    not g16803 ( n14530 , n25308 );
    nor g16804 ( n22335 , n8494 , n8582 );
    or g16805 ( n1391 , n8718 , n2095 );
    xnor g16806 ( n1134 , n28489 , n18091 );
    or g16807 ( n34662 , n26659 , n3954 );
    xnor g16808 ( n34113 , n40 , n29520 );
    nor g16809 ( n27106 , n10845 , n13065 );
    not g16810 ( n39645 , n32667 );
    and g16811 ( n15552 , n5052 , n34771 );
    xnor g16812 ( n36146 , n12487 , n20545 );
    and g16813 ( n4806 , n37039 , n12453 );
    or g16814 ( n25431 , n37305 , n29382 );
    not g16815 ( n5089 , n19763 );
    and g16816 ( n9913 , n4500 , n9088 );
    not g16817 ( n21173 , n16483 );
    nor g16818 ( n13004 , n15711 , n35419 );
    and g16819 ( n22750 , n14356 , n8211 );
    and g16820 ( n41750 , n26136 , n27301 );
    or g16821 ( n229 , n15272 , n34692 );
    not g16822 ( n5438 , n7038 );
    and g16823 ( n18833 , n34791 , n37774 );
    and g16824 ( n14552 , n39909 , n17331 );
    and g16825 ( n30325 , n29889 , n13487 );
    xnor g16826 ( n12494 , n2844 , n35301 );
    and g16827 ( n27760 , n32363 , n21474 );
    or g16828 ( n32338 , n28143 , n1266 );
    xnor g16829 ( n30250 , n22474 , n4958 );
    and g16830 ( n14586 , n28656 , n40711 );
    xnor g16831 ( n18176 , n2317 , n12850 );
    xnor g16832 ( n36362 , n26972 , n40602 );
    not g16833 ( n6351 , n37038 );
    and g16834 ( n36313 , n28480 , n22077 );
    and g16835 ( n2864 , n24491 , n35681 );
    and g16836 ( n20225 , n36297 , n25571 );
    not g16837 ( n17405 , n31637 );
    xnor g16838 ( n27815 , n14467 , n8550 );
    or g16839 ( n42066 , n33457 , n28335 );
    nor g16840 ( n15366 , n16848 , n36195 );
    or g16841 ( n22096 , n1971 , n35948 );
    xnor g16842 ( n36003 , n5679 , n4922 );
    xnor g16843 ( n6201 , n7004 , n11836 );
    or g16844 ( n21326 , n26489 , n18244 );
    not g16845 ( n1489 , n7624 );
    or g16846 ( n834 , n35803 , n18165 );
    or g16847 ( n26284 , n6434 , n22723 );
    and g16848 ( n13051 , n37655 , n36519 );
    and g16849 ( n165 , n17577 , n27605 );
    not g16850 ( n35938 , n24800 );
    and g16851 ( n34504 , n9990 , n4037 );
    nor g16852 ( n12490 , n14471 , n813 );
    or g16853 ( n7960 , n11913 , n6281 );
    or g16854 ( n12625 , n10549 , n26097 );
    nor g16855 ( n38024 , n20115 , n41485 );
    or g16856 ( n20050 , n17493 , n9617 );
    and g16857 ( n13584 , n17748 , n32014 );
    and g16858 ( n21711 , n10288 , n4392 );
    or g16859 ( n17784 , n29672 , n6517 );
    or g16860 ( n6846 , n9887 , n33262 );
    not g16861 ( n29682 , n3705 );
    or g16862 ( n1307 , n12970 , n12051 );
    or g16863 ( n33574 , n14723 , n28572 );
    or g16864 ( n29257 , n31200 , n24231 );
    or g16865 ( n24013 , n11977 , n17380 );
    xnor g16866 ( n38911 , n27184 , n29134 );
    and g16867 ( n2519 , n20319 , n20056 );
    not g16868 ( n36102 , n18660 );
    or g16869 ( n21622 , n27340 , n16636 );
    xnor g16870 ( n28879 , n42064 , n39155 );
    and g16871 ( n16335 , n28353 , n34264 );
    or g16872 ( n38204 , n31070 , n8829 );
    or g16873 ( n33663 , n6825 , n20556 );
    or g16874 ( n9491 , n14407 , n18774 );
    or g16875 ( n26913 , n33330 , n31458 );
    and g16876 ( n36630 , n34871 , n28133 );
    and g16877 ( n2140 , n3878 , n4770 );
    or g16878 ( n28842 , n7381 , n18360 );
    xnor g16879 ( n36707 , n25515 , n8206 );
    and g16880 ( n395 , n16807 , n1562 );
    nor g16881 ( n7488 , n19818 , n19121 );
    or g16882 ( n26602 , n6636 , n15373 );
    xnor g16883 ( n2467 , n11436 , n27701 );
    not g16884 ( n25504 , n11151 );
    or g16885 ( n24702 , n14657 , n10953 );
    and g16886 ( n3242 , n35605 , n42744 );
    and g16887 ( n34087 , n16416 , n22638 );
    xnor g16888 ( n34432 , n39912 , n42843 );
    or g16889 ( n28189 , n21199 , n12096 );
    not g16890 ( n33683 , n13540 );
    or g16891 ( n1650 , n35732 , n11405 );
    or g16892 ( n6222 , n4530 , n23438 );
    or g16893 ( n14159 , n11614 , n18541 );
    not g16894 ( n21512 , n41203 );
    or g16895 ( n5303 , n27539 , n20270 );
    nor g16896 ( n35490 , n32698 , n42225 );
    nor g16897 ( n5166 , n34566 , n20232 );
    and g16898 ( n22115 , n5479 , n36801 );
    or g16899 ( n29565 , n264 , n7894 );
    or g16900 ( n17752 , n5850 , n20568 );
    and g16901 ( n1138 , n40250 , n27649 );
    xnor g16902 ( n8043 , n18530 , n31679 );
    or g16903 ( n19895 , n23848 , n34115 );
    nor g16904 ( n32575 , n13728 , n727 );
    not g16905 ( n38953 , n33749 );
    not g16906 ( n9952 , n35774 );
    not g16907 ( n36584 , n34283 );
    or g16908 ( n23929 , n19702 , n26159 );
    nor g16909 ( n14703 , n2763 , n41897 );
    xnor g16910 ( n14330 , n18880 , n23632 );
    or g16911 ( n9927 , n36410 , n41588 );
    or g16912 ( n8600 , n29717 , n7121 );
    and g16913 ( n13147 , n13268 , n22026 );
    xnor g16914 ( n3258 , n28414 , n35200 );
    xnor g16915 ( n17579 , n35727 , n38601 );
    xnor g16916 ( n26451 , n40 , n8698 );
    not g16917 ( n10480 , n29247 );
    and g16918 ( n39588 , n13949 , n4507 );
    and g16919 ( n26433 , n3005 , n31320 );
    nor g16920 ( n11245 , n21598 , n25046 );
    and g16921 ( n8460 , n17097 , n18148 );
    or g16922 ( n23901 , n20145 , n11936 );
    or g16923 ( n11973 , n25990 , n41175 );
    and g16924 ( n31106 , n19628 , n29870 );
    nor g16925 ( n12702 , n16573 , n3330 );
    or g16926 ( n27797 , n34433 , n19509 );
    or g16927 ( n32834 , n33048 , n9752 );
    or g16928 ( n11448 , n29696 , n25705 );
    or g16929 ( n35402 , n1848 , n25637 );
    or g16930 ( n15159 , n19416 , n30715 );
    and g16931 ( n6182 , n14740 , n35853 );
    and g16932 ( n9785 , n38189 , n18527 );
    or g16933 ( n42662 , n27349 , n10306 );
    or g16934 ( n156 , n34485 , n15799 );
    or g16935 ( n22081 , n25959 , n18731 );
    or g16936 ( n40980 , n9314 , n4145 );
    not g16937 ( n36444 , n6442 );
    or g16938 ( n10336 , n31850 , n14262 );
    not g16939 ( n2802 , n37446 );
    or g16940 ( n14648 , n15894 , n34726 );
    and g16941 ( n11782 , n41673 , n23537 );
    xnor g16942 ( n21302 , n26972 , n36795 );
    and g16943 ( n27582 , n2797 , n3451 );
    not g16944 ( n29137 , n30680 );
    and g16945 ( n13492 , n32583 , n5922 );
    xnor g16946 ( n17646 , n14629 , n2071 );
    or g16947 ( n35137 , n32006 , n18206 );
    nor g16948 ( n12138 , n26609 , n27661 );
    or g16949 ( n10374 , n23374 , n6817 );
    xnor g16950 ( n4358 , n4659 , n26353 );
    not g16951 ( n7989 , n5250 );
    or g16952 ( n30770 , n38996 , n28918 );
    or g16953 ( n7897 , n28180 , n12153 );
    and g16954 ( n26607 , n12468 , n7332 );
    or g16955 ( n13754 , n7267 , n41007 );
    or g16956 ( n9158 , n17050 , n41973 );
    xnor g16957 ( n23363 , n11133 , n11362 );
    nor g16958 ( n28962 , n30338 , n33491 );
    not g16959 ( n19065 , n27966 );
    nor g16960 ( n27417 , n34292 , n19397 );
    nor g16961 ( n40185 , n31000 , n29950 );
    nor g16962 ( n3541 , n11506 , n28095 );
    and g16963 ( n18648 , n2266 , n16934 );
    nor g16964 ( n16207 , n15070 , n14142 );
    or g16965 ( n5753 , n22275 , n31497 );
    or g16966 ( n33661 , n24901 , n5813 );
    and g16967 ( n29127 , n32908 , n20447 );
    and g16968 ( n23711 , n36260 , n6489 );
    nor g16969 ( n24316 , n15285 , n12219 );
    or g16970 ( n32065 , n25873 , n21602 );
    xnor g16971 ( n18363 , n6769 , n15070 );
    or g16972 ( n21432 , n1662 , n3049 );
    xnor g16973 ( n31259 , n24998 , n16615 );
    or g16974 ( n6113 , n12993 , n42494 );
    xnor g16975 ( n18509 , n37953 , n19733 );
    xnor g16976 ( n40735 , n28917 , n37435 );
    not g16977 ( n21975 , n15004 );
    not g16978 ( n644 , n41321 );
    or g16979 ( n27732 , n40773 , n39409 );
    or g16980 ( n30529 , n24097 , n14508 );
    not g16981 ( n32980 , n16264 );
    xnor g16982 ( n4438 , n35553 , n25280 );
    not g16983 ( n6303 , n24856 );
    and g16984 ( n31168 , n21961 , n4931 );
    or g16985 ( n36476 , n15040 , n6459 );
    nor g16986 ( n22102 , n28617 , n38795 );
    or g16987 ( n6611 , n24745 , n24699 );
    and g16988 ( n21531 , n15367 , n38804 );
    xnor g16989 ( n11809 , n40993 , n10928 );
    nor g16990 ( n8265 , n32408 , n17509 );
    or g16991 ( n24889 , n11798 , n11381 );
    not g16992 ( n42516 , n33936 );
    nor g16993 ( n15365 , n39150 , n12690 );
    and g16994 ( n25126 , n28409 , n4025 );
    not g16995 ( n33484 , n15833 );
    or g16996 ( n40834 , n6247 , n1245 );
    and g16997 ( n1685 , n39658 , n33324 );
    not g16998 ( n33681 , n41311 );
    or g16999 ( n36508 , n7616 , n34661 );
    xnor g17000 ( n30492 , n31989 , n10816 );
    xnor g17001 ( n26199 , n31989 , n293 );
    nor g17002 ( n3623 , n15325 , n15208 );
    and g17003 ( n39955 , n28578 , n34710 );
    or g17004 ( n41771 , n6026 , n42880 );
    xnor g17005 ( n7926 , n898 , n13340 );
    xnor g17006 ( n32828 , n5013 , n25485 );
    nor g17007 ( n16324 , n1029 , n25122 );
    or g17008 ( n13406 , n37114 , n37748 );
    or g17009 ( n40615 , n19296 , n26811 );
    xnor g17010 ( n3948 , n23823 , n1928 );
    not g17011 ( n36948 , n13884 );
    nor g17012 ( n13346 , n34565 , n29564 );
    or g17013 ( n8962 , n10870 , n29545 );
    and g17014 ( n31845 , n14026 , n9260 );
    and g17015 ( n7150 , n20333 , n10377 );
    or g17016 ( n33521 , n3583 , n34218 );
    or g17017 ( n22012 , n2710 , n38554 );
    or g17018 ( n4817 , n32547 , n35413 );
    or g17019 ( n5709 , n25391 , n30852 );
    or g17020 ( n42187 , n6595 , n35866 );
    and g17021 ( n6886 , n32538 , n22132 );
    or g17022 ( n41320 , n8421 , n33943 );
    or g17023 ( n24733 , n2199 , n18927 );
    not g17024 ( n24826 , n8814 );
    or g17025 ( n41782 , n41351 , n34195 );
    not g17026 ( n32986 , n12278 );
    not g17027 ( n14252 , n20889 );
    and g17028 ( n14557 , n3388 , n24353 );
    not g17029 ( n27960 , n30877 );
    nor g17030 ( n17493 , n37130 , n12254 );
    nor g17031 ( n1647 , n31155 , n22169 );
    or g17032 ( n38179 , n4464 , n40323 );
    not g17033 ( n30110 , n1419 );
    not g17034 ( n1152 , n32337 );
    nor g17035 ( n20772 , n10594 , n23999 );
    xnor g17036 ( n26848 , n453 , n19963 );
    not g17037 ( n19126 , n7630 );
    or g17038 ( n3515 , n29027 , n31680 );
    or g17039 ( n33084 , n42076 , n19659 );
    or g17040 ( n3475 , n6560 , n16594 );
    xnor g17041 ( n40332 , n20204 , n20175 );
    or g17042 ( n27068 , n23261 , n15746 );
    not g17043 ( n4923 , n2377 );
    or g17044 ( n16788 , n9538 , n6713 );
    or g17045 ( n20470 , n10984 , n38691 );
    nor g17046 ( n13516 , n17120 , n21817 );
    or g17047 ( n10139 , n9264 , n37751 );
    or g17048 ( n13202 , n22173 , n5564 );
    or g17049 ( n2347 , n30887 , n17928 );
    not g17050 ( n26354 , n29389 );
    nor g17051 ( n18930 , n1507 , n27851 );
    or g17052 ( n18422 , n8948 , n39831 );
    xnor g17053 ( n40621 , n2182 , n30613 );
    and g17054 ( n38758 , n14632 , n24596 );
    or g17055 ( n28724 , n41705 , n24815 );
    nor g17056 ( n2619 , n10806 , n1774 );
    not g17057 ( n27967 , n8330 );
    xnor g17058 ( n9629 , n105 , n41460 );
    xnor g17059 ( n8003 , n26733 , n41522 );
    not g17060 ( n2971 , n33313 );
    not g17061 ( n18083 , n20156 );
    nor g17062 ( n26167 , n36806 , n30603 );
    or g17063 ( n23909 , n22069 , n27485 );
    and g17064 ( n4293 , n19077 , n16950 );
    not g17065 ( n14656 , n28755 );
    or g17066 ( n19136 , n10619 , n18987 );
    or g17067 ( n14371 , n37707 , n37663 );
    or g17068 ( n594 , n32212 , n40571 );
    or g17069 ( n41217 , n25526 , n36233 );
    and g17070 ( n7838 , n3430 , n22262 );
    or g17071 ( n15398 , n17054 , n4715 );
    and g17072 ( n4541 , n6564 , n12401 );
    nor g17073 ( n14483 , n38485 , n16012 );
    nor g17074 ( n27848 , n11497 , n33015 );
    and g17075 ( n41848 , n8544 , n39889 );
    xnor g17076 ( n585 , n4173 , n30158 );
    xnor g17077 ( n10133 , n10005 , n40437 );
    not g17078 ( n42792 , n31067 );
    or g17079 ( n12660 , n25588 , n7203 );
    or g17080 ( n6383 , n33179 , n41990 );
    and g17081 ( n14064 , n5803 , n31010 );
    or g17082 ( n8524 , n42546 , n29147 );
    and g17083 ( n39812 , n24873 , n11302 );
    or g17084 ( n21589 , n37821 , n31856 );
    and g17085 ( n30891 , n11833 , n12326 );
    not g17086 ( n18520 , n19014 );
    xnor g17087 ( n707 , n18146 , n8127 );
    or g17088 ( n24813 , n726 , n42538 );
    nor g17089 ( n12347 , n40662 , n42290 );
    or g17090 ( n7110 , n10956 , n12461 );
    or g17091 ( n27922 , n15594 , n40326 );
    or g17092 ( n39380 , n27804 , n1268 );
    xnor g17093 ( n22503 , n6625 , n11048 );
    or g17094 ( n15548 , n8220 , n9089 );
    and g17095 ( n31076 , n27370 , n26827 );
    nor g17096 ( n30407 , n13899 , n7267 );
    or g17097 ( n40403 , n9539 , n10839 );
    nor g17098 ( n4672 , n912 , n39368 );
    and g17099 ( n241 , n4325 , n31209 );
    nor g17100 ( n8283 , n7723 , n17362 );
    or g17101 ( n5846 , n21931 , n9447 );
    nor g17102 ( n11472 , n20345 , n1648 );
    or g17103 ( n36302 , n6153 , n37995 );
    and g17104 ( n37721 , n31655 , n1363 );
    and g17105 ( n33692 , n35644 , n10706 );
    not g17106 ( n21613 , n31685 );
    or g17107 ( n1678 , n8242 , n32194 );
    or g17108 ( n17637 , n12112 , n19115 );
    nor g17109 ( n36742 , n16554 , n24655 );
    nor g17110 ( n36116 , n39281 , n13770 );
    nor g17111 ( n12049 , n18233 , n15054 );
    or g17112 ( n25544 , n22603 , n29616 );
    not g17113 ( n2597 , n13979 );
    or g17114 ( n13908 , n1838 , n2726 );
    or g17115 ( n37624 , n10833 , n8716 );
    or g17116 ( n35638 , n6578 , n23003 );
    and g17117 ( n18536 , n36015 , n42682 );
    and g17118 ( n40126 , n16667 , n21432 );
    or g17119 ( n7103 , n31052 , n36767 );
    not g17120 ( n1006 , n41669 );
    or g17121 ( n33784 , n35445 , n33860 );
    or g17122 ( n19539 , n11620 , n4301 );
    or g17123 ( n12213 , n42530 , n22943 );
    nor g17124 ( n10886 , n32648 , n5948 );
    xnor g17125 ( n11541 , n2862 , n5035 );
    and g17126 ( n32640 , n36287 , n40687 );
    and g17127 ( n33453 , n38923 , n9236 );
    or g17128 ( n40314 , n7604 , n106 );
    or g17129 ( n17802 , n9031 , n10349 );
    nor g17130 ( n23019 , n42465 , n2607 );
    nor g17131 ( n12377 , n19181 , n20735 );
    nor g17132 ( n39404 , n11903 , n39710 );
    not g17133 ( n41132 , n27043 );
    and g17134 ( n30825 , n4927 , n35485 );
    and g17135 ( n41448 , n12029 , n35784 );
    and g17136 ( n4694 , n18906 , n18152 );
    and g17137 ( n18618 , n16969 , n6942 );
    or g17138 ( n17999 , n9400 , n42184 );
    xnor g17139 ( n3840 , n5246 , n699 );
    not g17140 ( n38146 , n7678 );
    xnor g17141 ( n36905 , n1196 , n243 );
    and g17142 ( n12555 , n32401 , n29198 );
    or g17143 ( n11221 , n27072 , n40485 );
    or g17144 ( n32961 , n11415 , n29856 );
    and g17145 ( n6772 , n30746 , n37814 );
    and g17146 ( n31953 , n22846 , n15944 );
    or g17147 ( n23997 , n23565 , n10623 );
    not g17148 ( n20360 , n15441 );
    nor g17149 ( n10738 , n17120 , n29789 );
    nor g17150 ( n5665 , n751 , n41227 );
    xnor g17151 ( n16554 , n16693 , n32185 );
    xnor g17152 ( n27994 , n4334 , n38465 );
    or g17153 ( n40230 , n2270 , n21615 );
    or g17154 ( n38614 , n34664 , n9420 );
    not g17155 ( n32213 , n32443 );
    xnor g17156 ( n21263 , n30832 , n25567 );
    and g17157 ( n28568 , n25584 , n4455 );
    nor g17158 ( n32255 , n4416 , n31216 );
    or g17159 ( n24567 , n33834 , n2576 );
    or g17160 ( n24768 , n37119 , n6848 );
    xnor g17161 ( n31811 , n19605 , n12767 );
    or g17162 ( n2365 , n3054 , n3675 );
    or g17163 ( n27813 , n14378 , n24626 );
    nor g17164 ( n11165 , n5896 , n31779 );
    or g17165 ( n15665 , n33241 , n23489 );
    or g17166 ( n28462 , n42324 , n37465 );
    or g17167 ( n19024 , n34838 , n31132 );
    or g17168 ( n16273 , n42596 , n12383 );
    xnor g17169 ( n33170 , n13415 , n35853 );
    and g17170 ( n29021 , n39235 , n42044 );
    not g17171 ( n13423 , n32567 );
    and g17172 ( n428 , n9546 , n18985 );
    xnor g17173 ( n35409 , n24645 , n23885 );
    or g17174 ( n16760 , n7017 , n34440 );
    not g17175 ( n14712 , n34880 );
    not g17176 ( n12532 , n9626 );
    and g17177 ( n17641 , n1971 , n18816 );
    and g17178 ( n37776 , n15605 , n42872 );
    xnor g17179 ( n2743 , n30862 , n40186 );
    or g17180 ( n36008 , n12830 , n21926 );
    or g17181 ( n27217 , n21179 , n19266 );
    or g17182 ( n30151 , n15150 , n27305 );
    or g17183 ( n39376 , n2131 , n42479 );
    and g17184 ( n41883 , n35154 , n41726 );
    and g17185 ( n41772 , n20014 , n35137 );
    not g17186 ( n35477 , n32573 );
    xnor g17187 ( n6421 , n31989 , n19371 );
    or g17188 ( n40820 , n23598 , n7263 );
    or g17189 ( n30509 , n28634 , n28330 );
    or g17190 ( n21185 , n36898 , n19701 );
    and g17191 ( n42448 , n16662 , n21591 );
    nor g17192 ( n10763 , n14707 , n13212 );
    not g17193 ( n32480 , n22389 );
    nor g17194 ( n2460 , n14471 , n38601 );
    xnor g17195 ( n21165 , n31370 , n19221 );
    or g17196 ( n36482 , n29021 , n39213 );
    and g17197 ( n7810 , n24654 , n4573 );
    or g17198 ( n21701 , n24547 , n1948 );
    and g17199 ( n17304 , n2960 , n15032 );
    not g17200 ( n33859 , n41759 );
    nor g17201 ( n20819 , n9336 , n9813 );
    xnor g17202 ( n22782 , n12806 , n32991 );
    or g17203 ( n42147 , n38266 , n14561 );
    nor g17204 ( n19982 , n22915 , n620 );
    or g17205 ( n36567 , n32977 , n26027 );
    not g17206 ( n21116 , n4030 );
    or g17207 ( n27996 , n42887 , n31227 );
    or g17208 ( n38198 , n29455 , n36717 );
    not g17209 ( n34818 , n31726 );
    nor g17210 ( n18180 , n39740 , n16310 );
    or g17211 ( n3741 , n25561 , n39627 );
    or g17212 ( n14834 , n14396 , n16970 );
    and g17213 ( n5210 , n26726 , n41832 );
    not g17214 ( n25602 , n34500 );
    or g17215 ( n13595 , n25836 , n39166 );
    and g17216 ( n14587 , n40377 , n27216 );
    not g17217 ( n8641 , n24610 );
    or g17218 ( n24809 , n5960 , n22739 );
    and g17219 ( n33597 , n14774 , n25946 );
    xnor g17220 ( n27877 , n6066 , n15576 );
    and g17221 ( n1279 , n24041 , n21506 );
    and g17222 ( n4402 , n15288 , n36732 );
    xnor g17223 ( n18537 , n8928 , n2434 );
    or g17224 ( n19295 , n28080 , n7997 );
    and g17225 ( n13573 , n29629 , n8965 );
    nor g17226 ( n7837 , n5605 , n4694 );
    xnor g17227 ( n6048 , n2327 , n35839 );
    or g17228 ( n36586 , n27840 , n17306 );
    or g17229 ( n17227 , n2946 , n5760 );
    or g17230 ( n25679 , n37059 , n32876 );
    or g17231 ( n24597 , n38464 , n37647 );
    and g17232 ( n14687 , n22208 , n13180 );
    and g17233 ( n34843 , n9686 , n10237 );
    or g17234 ( n10128 , n23698 , n30071 );
    xnor g17235 ( n12577 , n35967 , n23798 );
    or g17236 ( n13962 , n37967 , n21875 );
    nor g17237 ( n13360 , n19990 , n34884 );
    not g17238 ( n33794 , n25105 );
    xnor g17239 ( n11103 , n35727 , n24864 );
    and g17240 ( n14245 , n16356 , n16265 );
    not g17241 ( n23184 , n19614 );
    or g17242 ( n6259 , n14945 , n34300 );
    or g17243 ( n34402 , n1816 , n41873 );
    and g17244 ( n35539 , n29704 , n12689 );
    nor g17245 ( n11918 , n9793 , n34300 );
    or g17246 ( n26551 , n12722 , n41322 );
    nor g17247 ( n17042 , n14471 , n29012 );
    xnor g17248 ( n23060 , n456 , n33981 );
    not g17249 ( n13105 , n21643 );
    and g17250 ( n25234 , n10256 , n4568 );
    and g17251 ( n12778 , n28724 , n41073 );
    xnor g17252 ( n20822 , n30628 , n11843 );
    nor g17253 ( n20 , n2966 , n14523 );
    not g17254 ( n26279 , n32814 );
    not g17255 ( n40059 , n31506 );
    or g17256 ( n8406 , n4506 , n21829 );
    or g17257 ( n35075 , n35823 , n26961 );
    not g17258 ( n6111 , n42301 );
    xnor g17259 ( n4695 , n18736 , n3402 );
    not g17260 ( n21866 , n35793 );
    and g17261 ( n28128 , n32030 , n2764 );
    and g17262 ( n30326 , n21508 , n18448 );
    xnor g17263 ( n8507 , n11217 , n6357 );
    nor g17264 ( n30345 , n7297 , n10864 );
    or g17265 ( n24366 , n27163 , n25626 );
    and g17266 ( n20936 , n23245 , n20635 );
    or g17267 ( n22204 , n16409 , n8319 );
    not g17268 ( n34578 , n30178 );
    and g17269 ( n30737 , n42050 , n4438 );
    not g17270 ( n23136 , n23722 );
    xnor g17271 ( n24323 , n4949 , n39399 );
    and g17272 ( n8156 , n10379 , n25378 );
    not g17273 ( n41756 , n23896 );
    xnor g17274 ( n4087 , n8135 , n28509 );
    nor g17275 ( n32344 , n20952 , n33930 );
    or g17276 ( n22975 , n35083 , n39937 );
    xnor g17277 ( n36924 , n1249 , n16185 );
    or g17278 ( n9540 , n36719 , n31361 );
    xnor g17279 ( n3391 , n18530 , n3498 );
    not g17280 ( n8663 , n38992 );
    not g17281 ( n10674 , n41955 );
    xnor g17282 ( n19032 , n42060 , n13861 );
    and g17283 ( n8798 , n237 , n12884 );
    not g17284 ( n5041 , n8504 );
    or g17285 ( n13518 , n38463 , n30241 );
    and g17286 ( n466 , n9121 , n38158 );
    xnor g17287 ( n15711 , n6969 , n41714 );
    xnor g17288 ( n17902 , n19300 , n31458 );
    nor g17289 ( n157 , n8494 , n32183 );
    and g17290 ( n1380 , n42506 , n3284 );
    or g17291 ( n36694 , n16367 , n5984 );
    and g17292 ( n37180 , n36462 , n23412 );
    xnor g17293 ( n38607 , n9460 , n41871 );
    or g17294 ( n21627 , n35301 , n4901 );
    xnor g17295 ( n25412 , n27371 , n33864 );
    xnor g17296 ( n40680 , n5041 , n10037 );
    not g17297 ( n30985 , n18385 );
    or g17298 ( n4777 , n3636 , n30547 );
    or g17299 ( n22066 , n15529 , n2383 );
    and g17300 ( n17126 , n34970 , n41931 );
    not g17301 ( n25426 , n28051 );
    or g17302 ( n8858 , n25451 , n40527 );
    nor g17303 ( n29847 , n38927 , n29208 );
    and g17304 ( n5587 , n30209 , n7515 );
    and g17305 ( n29311 , n8906 , n22923 );
    or g17306 ( n20771 , n9636 , n12153 );
    or g17307 ( n23812 , n33513 , n17109 );
    or g17308 ( n32428 , n35779 , n2647 );
    nor g17309 ( n30137 , n14298 , n39304 );
    or g17310 ( n39466 , n27169 , n30821 );
    not g17311 ( n14502 , n33130 );
    and g17312 ( n2939 , n7140 , n5580 );
    and g17313 ( n34392 , n483 , n5238 );
    or g17314 ( n15091 , n33655 , n35540 );
    nor g17315 ( n3744 , n20015 , n832 );
    or g17316 ( n5429 , n36727 , n10204 );
    or g17317 ( n32257 , n11522 , n471 );
    or g17318 ( n15128 , n31109 , n38416 );
    or g17319 ( n37889 , n27960 , n7714 );
    not g17320 ( n34383 , n9353 );
    or g17321 ( n32742 , n41777 , n1788 );
    or g17322 ( n4378 , n13412 , n29833 );
    nor g17323 ( n42703 , n9020 , n11695 );
    nor g17324 ( n42449 , n17193 , n11597 );
    nor g17325 ( n27359 , n40950 , n32847 );
    not g17326 ( n22379 , n5097 );
    and g17327 ( n27330 , n24320 , n31173 );
    nor g17328 ( n19884 , n8694 , n3643 );
    or g17329 ( n11687 , n41535 , n2658 );
    xnor g17330 ( n23730 , n23944 , n29864 );
    and g17331 ( n1039 , n18357 , n8154 );
    or g17332 ( n6528 , n25575 , n21025 );
    or g17333 ( n18562 , n550 , n22868 );
    or g17334 ( n6783 , n24024 , n38196 );
    or g17335 ( n12697 , n14070 , n28904 );
    not g17336 ( n11085 , n3198 );
    xnor g17337 ( n34658 , n18812 , n4631 );
    nor g17338 ( n20010 , n29882 , n3285 );
    and g17339 ( n34885 , n26218 , n23230 );
    nor g17340 ( n6218 , n11136 , n13809 );
    or g17341 ( n35146 , n7478 , n9809 );
    or g17342 ( n31270 , n37312 , n7359 );
    and g17343 ( n42185 , n37985 , n19321 );
    nor g17344 ( n30772 , n24809 , n19555 );
    not g17345 ( n17272 , n19629 );
    not g17346 ( n13646 , n8849 );
    nor g17347 ( n40729 , n19905 , n19690 );
    not g17348 ( n23686 , n2857 );
    or g17349 ( n1529 , n27363 , n26922 );
    nor g17350 ( n30814 , n27229 , n2487 );
    or g17351 ( n35493 , n40358 , n9488 );
    or g17352 ( n29467 , n23634 , n39463 );
    not g17353 ( n13473 , n18894 );
    or g17354 ( n2693 , n11639 , n27540 );
    nor g17355 ( n19056 , n21907 , n22050 );
    not g17356 ( n1223 , n26817 );
    xnor g17357 ( n1046 , n21973 , n27372 );
    or g17358 ( n34230 , n25033 , n7465 );
    or g17359 ( n14488 , n42144 , n41993 );
    nor g17360 ( n30293 , n27026 , n12886 );
    or g17361 ( n19897 , n10247 , n11108 );
    and g17362 ( n24614 , n19528 , n23471 );
    or g17363 ( n21974 , n2099 , n31071 );
    or g17364 ( n1784 , n16416 , n22638 );
    or g17365 ( n10030 , n13370 , n21268 );
    or g17366 ( n18586 , n41433 , n42763 );
    or g17367 ( n29652 , n11346 , n1632 );
    not g17368 ( n36012 , n7984 );
    not g17369 ( n24180 , n5522 );
    and g17370 ( n39661 , n40537 , n35222 );
    and g17371 ( n9263 , n15913 , n2200 );
    or g17372 ( n37946 , n27681 , n3571 );
    or g17373 ( n31130 , n35267 , n14387 );
    not g17374 ( n26597 , n4836 );
    and g17375 ( n30735 , n36529 , n25463 );
    or g17376 ( n2081 , n32111 , n13367 );
    and g17377 ( n23986 , n26775 , n21449 );
    nor g17378 ( n23332 , n36607 , n39834 );
    and g17379 ( n27914 , n32669 , n22368 );
    xnor g17380 ( n10056 , n4467 , n24662 );
    and g17381 ( n16801 , n27893 , n18478 );
    and g17382 ( n4825 , n36048 , n40106 );
    and g17383 ( n9848 , n6518 , n2712 );
    or g17384 ( n42407 , n2628 , n15894 );
    or g17385 ( n28064 , n4672 , n498 );
    or g17386 ( n41362 , n11347 , n13190 );
    xnor g17387 ( n33231 , n25985 , n36195 );
    not g17388 ( n35578 , n37601 );
    not g17389 ( n32252 , n4476 );
    nor g17390 ( n11693 , n4651 , n18868 );
    or g17391 ( n18739 , n7771 , n16402 );
    nor g17392 ( n42461 , n22175 , n36328 );
    and g17393 ( n1558 , n4480 , n17555 );
    and g17394 ( n40913 , n8332 , n25604 );
    nor g17395 ( n31417 , n9084 , n13635 );
    not g17396 ( n801 , n6489 );
    or g17397 ( n39183 , n9998 , n35465 );
    or g17398 ( n17805 , n23092 , n21268 );
    or g17399 ( n4191 , n33210 , n23374 );
    or g17400 ( n1421 , n20138 , n23000 );
    or g17401 ( n15344 , n24831 , n15460 );
    or g17402 ( n1045 , n2041 , n5057 );
    not g17403 ( n32800 , n7824 );
    or g17404 ( n7047 , n17469 , n17865 );
    and g17405 ( n3814 , n29740 , n31453 );
    or g17406 ( n9193 , n13544 , n22365 );
    and g17407 ( n9802 , n39762 , n39894 );
    or g17408 ( n28104 , n15525 , n6435 );
    or g17409 ( n6738 , n34921 , n41765 );
    not g17410 ( n35087 , n1234 );
    or g17411 ( n21465 , n39195 , n31317 );
    or g17412 ( n10757 , n26350 , n22194 );
    and g17413 ( n23334 , n29584 , n20998 );
    or g17414 ( n23752 , n22201 , n39079 );
    xnor g17415 ( n23606 , n19700 , n6845 );
    nor g17416 ( n968 , n29859 , n10007 );
    xnor g17417 ( n23504 , n40 , n19004 );
    xnor g17418 ( n35956 , n20237 , n23435 );
    and g17419 ( n3981 , n14349 , n32450 );
    nor g17420 ( n28166 , n26394 , n32100 );
    nor g17421 ( n36032 , n11985 , n30433 );
    and g17422 ( n36491 , n9929 , n23685 );
    or g17423 ( n11547 , n36318 , n11829 );
    xnor g17424 ( n38725 , n38261 , n8309 );
    not g17425 ( n1735 , n31364 );
    or g17426 ( n2552 , n41122 , n42701 );
    not g17427 ( n27187 , n15383 );
    xnor g17428 ( n14814 , n35311 , n27473 );
    and g17429 ( n14161 , n14739 , n42789 );
    not g17430 ( n36272 , n2846 );
    and g17431 ( n12058 , n6300 , n17705 );
    or g17432 ( n34888 , n20446 , n20497 );
    or g17433 ( n23454 , n20451 , n34796 );
    and g17434 ( n41317 , n41325 , n39693 );
    or g17435 ( n15075 , n32635 , n42544 );
    or g17436 ( n10062 , n7048 , n24114 );
    nor g17437 ( n8149 , n38879 , n23420 );
    not g17438 ( n13144 , n39364 );
    xnor g17439 ( n31841 , n9478 , n20247 );
    or g17440 ( n29307 , n37637 , n39012 );
    or g17441 ( n30352 , n31999 , n41702 );
    nor g17442 ( n6162 , n1260 , n3861 );
    nor g17443 ( n38937 , n13174 , n1928 );
    or g17444 ( n38549 , n8730 , n16964 );
    not g17445 ( n22378 , n34654 );
    nor g17446 ( n22791 , n18866 , n293 );
    nor g17447 ( n15802 , n5964 , n29228 );
    or g17448 ( n12731 , n11941 , n35829 );
    or g17449 ( n21774 , n16805 , n12153 );
    or g17450 ( n30816 , n17700 , n42891 );
    and g17451 ( n20100 , n28040 , n39785 );
    or g17452 ( n829 , n10286 , n18016 );
    nor g17453 ( n5051 , n37953 , n1951 );
    nor g17454 ( n28803 , n15454 , n33005 );
    or g17455 ( n20961 , n27126 , n30983 );
    not g17456 ( n27570 , n4296 );
    or g17457 ( n3532 , n15593 , n24371 );
    nor g17458 ( n26205 , n18866 , n10691 );
    not g17459 ( n27420 , n1515 );
    or g17460 ( n36462 , n9799 , n14749 );
    or g17461 ( n16289 , n17108 , n28293 );
    or g17462 ( n23892 , n16564 , n11683 );
    xnor g17463 ( n9326 , n37403 , n2286 );
    nor g17464 ( n3001 , n35301 , n38783 );
    not g17465 ( n39878 , n33648 );
    or g17466 ( n3126 , n23786 , n29930 );
    or g17467 ( n3273 , n7412 , n27189 );
    xnor g17468 ( n30128 , n25584 , n4455 );
    not g17469 ( n9564 , n20960 );
    not g17470 ( n41253 , n36114 );
    nor g17471 ( n29033 , n14707 , n5455 );
    not g17472 ( n13476 , n15435 );
    and g17473 ( n7914 , n4413 , n800 );
    xnor g17474 ( n15309 , n4334 , n19927 );
    or g17475 ( n28105 , n17040 , n27817 );
    nor g17476 ( n14292 , n31723 , n13678 );
    or g17477 ( n17960 , n23548 , n29136 );
    and g17478 ( n23268 , n35986 , n37187 );
    and g17479 ( n24391 , n22304 , n40320 );
    or g17480 ( n2128 , n15295 , n21912 );
    nor g17481 ( n19247 , n15515 , n19959 );
    or g17482 ( n33424 , n16717 , n8803 );
    xnor g17483 ( n10767 , n27250 , n3643 );
    and g17484 ( n10568 , n27318 , n1982 );
    or g17485 ( n39425 , n33104 , n10704 );
    not g17486 ( n4484 , n14346 );
    xnor g17487 ( n4188 , n30022 , n34215 );
    not g17488 ( n18625 , n19861 );
    and g17489 ( n6385 , n2230 , n30523 );
    or g17490 ( n38719 , n6723 , n14668 );
    nor g17491 ( n10539 , n966 , n29836 );
    and g17492 ( n15707 , n9741 , n8257 );
    or g17493 ( n28819 , n17849 , n23880 );
    and g17494 ( n27988 , n3929 , n29718 );
    and g17495 ( n2061 , n2384 , n40822 );
    not g17496 ( n26475 , n33130 );
    nor g17497 ( n16031 , n4896 , n19379 );
    not g17498 ( n22948 , n16567 );
    and g17499 ( n40418 , n23191 , n25278 );
    not g17500 ( n15844 , n12728 );
    not g17501 ( n7476 , n19892 );
    or g17502 ( n4641 , n26258 , n25615 );
    or g17503 ( n5510 , n20138 , n18925 );
    xnor g17504 ( n1196 , n5144 , n21176 );
    or g17505 ( n35414 , n31437 , n36962 );
    or g17506 ( n25119 , n34411 , n35177 );
    not g17507 ( n25817 , n31138 );
    or g17508 ( n1308 , n1383 , n22645 );
    or g17509 ( n40743 , n13104 , n35538 );
    and g17510 ( n14326 , n32137 , n27981 );
    xnor g17511 ( n20872 , n21610 , n9569 );
    xnor g17512 ( n29852 , n42444 , n40045 );
    and g17513 ( n30232 , n5753 , n27304 );
    xnor g17514 ( n3435 , n330 , n134 );
    or g17515 ( n10000 , n30911 , n3907 );
    or g17516 ( n33357 , n6363 , n22413 );
    or g17517 ( n30108 , n9343 , n30455 );
    not g17518 ( n30684 , n1986 );
    xnor g17519 ( n29461 , n6625 , n3910 );
    not g17520 ( n8700 , n42244 );
    or g17521 ( n34963 , n38500 , n4772 );
    and g17522 ( n7043 , n13613 , n16777 );
    or g17523 ( n1243 , n15310 , n33537 );
    and g17524 ( n26546 , n42293 , n34314 );
    nor g17525 ( n23935 , n27705 , n35245 );
    or g17526 ( n33948 , n41913 , n15674 );
    xnor g17527 ( n19230 , n11534 , n1190 );
    or g17528 ( n33520 , n10925 , n6842 );
    or g17529 ( n5778 , n14481 , n36312 );
    and g17530 ( n40722 , n25156 , n5632 );
    or g17531 ( n20551 , n28725 , n18271 );
    nor g17532 ( n24001 , n39167 , n13755 );
    and g17533 ( n36430 , n20487 , n40917 );
    xnor g17534 ( n3889 , n13444 , n38783 );
    or g17535 ( n160 , n5605 , n16929 );
    and g17536 ( n19129 , n39914 , n32950 );
    and g17537 ( n38317 , n28787 , n12277 );
    xnor g17538 ( n20723 , n17272 , n41107 );
    not g17539 ( n7489 , n7356 );
    and g17540 ( n18073 , n41192 , n33688 );
    nor g17541 ( n15432 , n32297 , n27759 );
    not g17542 ( n38467 , n530 );
    and g17543 ( n8739 , n20765 , n33374 );
    and g17544 ( n26224 , n22758 , n41202 );
    or g17545 ( n24576 , n38921 , n14449 );
    or g17546 ( n26850 , n28134 , n7280 );
    or g17547 ( n36178 , n7429 , n12393 );
    and g17548 ( n32662 , n25680 , n24130 );
    and g17549 ( n11857 , n16743 , n21107 );
    nor g17550 ( n34640 , n36486 , n20321 );
    or g17551 ( n16425 , n38064 , n38109 );
    xnor g17552 ( n22397 , n42725 , n36040 );
    and g17553 ( n30570 , n29188 , n3858 );
    or g17554 ( n8607 , n27914 , n30630 );
    or g17555 ( n28181 , n13730 , n24108 );
    and g17556 ( n10410 , n31093 , n37735 );
    or g17557 ( n41648 , n11374 , n37353 );
    or g17558 ( n12309 , n4842 , n13861 );
    nor g17559 ( n41966 , n28974 , n9346 );
    and g17560 ( n4738 , n13858 , n23644 );
    and g17561 ( n8306 , n21200 , n5606 );
    not g17562 ( n35026 , n9818 );
    or g17563 ( n29200 , n22405 , n12392 );
    or g17564 ( n20873 , n9835 , n30467 );
    nor g17565 ( n18691 , n37643 , n39794 );
    not g17566 ( n23326 , n19735 );
    not g17567 ( n33464 , n26641 );
    xnor g17568 ( n32216 , n5487 , n36650 );
    xnor g17569 ( n11570 , n36998 , n15974 );
    or g17570 ( n11402 , n35320 , n27691 );
    nor g17571 ( n4726 , n16953 , n4986 );
    or g17572 ( n14208 , n8220 , n24260 );
    or g17573 ( n14339 , n22619 , n3648 );
    or g17574 ( n38490 , n10353 , n32588 );
    or g17575 ( n16503 , n11492 , n35964 );
    or g17576 ( n15518 , n5964 , n39237 );
    or g17577 ( n10219 , n8039 , n29856 );
    or g17578 ( n27966 , n8912 , n39454 );
    nor g17579 ( n21132 , n26443 , n8099 );
    xnor g17580 ( n41395 , n21654 , n6037 );
    nor g17581 ( n15912 , n21286 , n12371 );
    or g17582 ( n40681 , n41738 , n34144 );
    not g17583 ( n18260 , n27561 );
    and g17584 ( n8175 , n23997 , n35863 );
    or g17585 ( n16226 , n2353 , n20498 );
    and g17586 ( n7879 , n40130 , n38032 );
    and g17587 ( n20834 , n24102 , n32010 );
    xnor g17588 ( n149 , n25912 , n32629 );
    or g17589 ( n13113 , n6370 , n12988 );
    and g17590 ( n23094 , n16924 , n9213 );
    nor g17591 ( n22471 , n7300 , n39348 );
    or g17592 ( n32034 , n2430 , n27727 );
    not g17593 ( n38376 , n40508 );
    or g17594 ( n18819 , n20030 , n33008 );
    nor g17595 ( n11791 , n27524 , n35629 );
    not g17596 ( n41430 , n40979 );
    or g17597 ( n41188 , n31674 , n18305 );
    not g17598 ( n7355 , n18588 );
    not g17599 ( n41053 , n36309 );
    xnor g17600 ( n2650 , n26446 , n29082 );
    not g17601 ( n10044 , n27265 );
    xnor g17602 ( n12902 , n24118 , n13405 );
    xnor g17603 ( n15630 , n36009 , n35023 );
    or g17604 ( n34777 , n5294 , n34916 );
    xnor g17605 ( n39485 , n5144 , n5647 );
    or g17606 ( n5393 , n10244 , n34648 );
    and g17607 ( n18305 , n27850 , n11330 );
    or g17608 ( n20671 , n20229 , n8442 );
    or g17609 ( n42574 , n40228 , n6893 );
    nor g17610 ( n35190 , n36491 , n27954 );
    not g17611 ( n42251 , n24135 );
    not g17612 ( n41218 , n24610 );
    or g17613 ( n37259 , n40104 , n22892 );
    or g17614 ( n30805 , n35071 , n33679 );
    or g17615 ( n6047 , n5492 , n17915 );
    nor g17616 ( n23709 , n19813 , n13100 );
    and g17617 ( n26277 , n35666 , n29350 );
    or g17618 ( n5632 , n14851 , n38601 );
    or g17619 ( n40628 , n23656 , n33464 );
    or g17620 ( n36756 , n26172 , n30812 );
    or g17621 ( n5000 , n42320 , n15902 );
    and g17622 ( n1816 , n7059 , n25879 );
    not g17623 ( n6969 , n19485 );
    and g17624 ( n11495 , n32436 , n39654 );
    or g17625 ( n39185 , n11321 , n3975 );
    or g17626 ( n6108 , n23584 , n36922 );
    and g17627 ( n487 , n42048 , n24204 );
    xnor g17628 ( n30828 , n14364 , n1740 );
    or g17629 ( n8860 , n20921 , n6154 );
    and g17630 ( n25677 , n30420 , n33898 );
    nor g17631 ( n22271 , n1507 , n21357 );
    or g17632 ( n17813 , n14492 , n24375 );
    or g17633 ( n12632 , n14959 , n12059 );
    xnor g17634 ( n19996 , n10825 , n27083 );
    and g17635 ( n24340 , n32655 , n31814 );
    or g17636 ( n4838 , n30843 , n19159 );
    or g17637 ( n2409 , n2586 , n16966 );
    or g17638 ( n6217 , n25535 , n25481 );
    xnor g17639 ( n12675 , n19718 , n34077 );
    not g17640 ( n12308 , n24531 );
    and g17641 ( n19329 , n28170 , n34156 );
    nor g17642 ( n950 , n23995 , n11576 );
    or g17643 ( n31533 , n4446 , n3636 );
    not g17644 ( n20477 , n38094 );
    not g17645 ( n25577 , n37355 );
    not g17646 ( n26915 , n5947 );
    xnor g17647 ( n191 , n29889 , n13487 );
    or g17648 ( n16517 , n36374 , n17024 );
    nor g17649 ( n9745 , n36667 , n30653 );
    or g17650 ( n4182 , n4670 , n28849 );
    or g17651 ( n23537 , n12781 , n17457 );
    nor g17652 ( n38336 , n4659 , n29071 );
    or g17653 ( n6986 , n11316 , n29638 );
    or g17654 ( n8614 , n39976 , n38912 );
    xnor g17655 ( n30956 , n15972 , n25129 );
    xnor g17656 ( n30074 , n6978 , n8284 );
    or g17657 ( n29993 , n1971 , n1870 );
    or g17658 ( n31451 , n24883 , n29833 );
    xnor g17659 ( n17821 , n31099 , n25021 );
    or g17660 ( n41778 , n20811 , n10965 );
    and g17661 ( n42218 , n21599 , n9723 );
    and g17662 ( n25109 , n39631 , n27749 );
    and g17663 ( n17464 , n20562 , n10328 );
    or g17664 ( n32757 , n42699 , n29082 );
    not g17665 ( n12048 , n6069 );
    or g17666 ( n1258 , n8683 , n4627 );
    not g17667 ( n42097 , n4886 );
    nor g17668 ( n34250 , n5896 , n14491 );
    xnor g17669 ( n36546 , n25061 , n18866 );
    or g17670 ( n23864 , n12129 , n28559 );
    xnor g17671 ( n31226 , n37899 , n9680 );
    nor g17672 ( n29161 , n14746 , n15216 );
    and g17673 ( n32303 , n25595 , n5399 );
    not g17674 ( n4644 , n3706 );
    or g17675 ( n11966 , n6838 , n425 );
    or g17676 ( n16091 , n42007 , n15430 );
    or g17677 ( n16245 , n2583 , n24403 );
    xnor g17678 ( n22073 , n30271 , n41401 );
    or g17679 ( n4347 , n12700 , n2278 );
    not g17680 ( n14281 , n9432 );
    or g17681 ( n36068 , n38556 , n14963 );
    xnor g17682 ( n10457 , n37176 , n39817 );
    and g17683 ( n6744 , n26540 , n7457 );
    not g17684 ( n4298 , n116 );
    and g17685 ( n10936 , n18451 , n14243 );
    xnor g17686 ( n38372 , n21217 , n36117 );
    and g17687 ( n27836 , n37420 , n29795 );
    and g17688 ( n22578 , n12064 , n1552 );
    not g17689 ( n30281 , n21258 );
    and g17690 ( n34804 , n23903 , n41949 );
    or g17691 ( n32229 , n3813 , n14222 );
    or g17692 ( n11876 , n4900 , n31958 );
    or g17693 ( n28728 , n6792 , n32883 );
    and g17694 ( n12650 , n20836 , n15873 );
    or g17695 ( n8782 , n36117 , n39171 );
    and g17696 ( n23974 , n14253 , n34619 );
    not g17697 ( n32369 , n11889 );
    or g17698 ( n28382 , n11180 , n38423 );
    xnor g17699 ( n28507 , n4324 , n22795 );
    xnor g17700 ( n9732 , n40707 , n31280 );
    or g17701 ( n26705 , n36249 , n39898 );
    not g17702 ( n40109 , n32476 );
    not g17703 ( n10971 , n35998 );
    or g17704 ( n34879 , n16030 , n5984 );
    nor g17705 ( n38307 , n72 , n2503 );
    nor g17706 ( n30591 , n14471 , n7854 );
    not g17707 ( n1324 , n4851 );
    or g17708 ( n28027 , n22371 , n10935 );
    not g17709 ( n4949 , n14394 );
    not g17710 ( n7927 , n3509 );
    or g17711 ( n12204 , n32944 , n37122 );
    and g17712 ( n39400 , n15995 , n5609 );
    and g17713 ( n6327 , n42142 , n12089 );
    not g17714 ( n27087 , n22338 );
    not g17715 ( n28541 , n12514 );
    or g17716 ( n24167 , n10731 , n25528 );
    or g17717 ( n40442 , n30420 , n21096 );
    or g17718 ( n35243 , n2517 , n19073 );
    or g17719 ( n6364 , n18002 , n42065 );
    not g17720 ( n27463 , n7109 );
    or g17721 ( n15449 , n23125 , n32642 );
    nor g17722 ( n19409 , n21347 , n39460 );
    or g17723 ( n7828 , n7265 , n37234 );
    not g17724 ( n38693 , n18594 );
    or g17725 ( n30219 , n21002 , n22885 );
    nor g17726 ( n33549 , n25913 , n36145 );
    and g17727 ( n13172 , n38225 , n8666 );
    xnor g17728 ( n20387 , n35653 , n33052 );
    and g17729 ( n11433 , n33478 , n38842 );
    not g17730 ( n17415 , n7393 );
    xnor g17731 ( n11232 , n9796 , n12766 );
    or g17732 ( n16540 , n10571 , n15341 );
    or g17733 ( n29142 , n21794 , n11069 );
    xnor g17734 ( n33958 , n31973 , n17747 );
    and g17735 ( n27211 , n40949 , n18254 );
    or g17736 ( n27692 , n12926 , n16636 );
    or g17737 ( n31249 , n38421 , n26147 );
    or g17738 ( n24158 , n31480 , n10306 );
    or g17739 ( n18389 , n30741 , n21064 );
    or g17740 ( n36011 , n9553 , n4293 );
    or g17741 ( n37121 , n11773 , n16925 );
    xnor g17742 ( n27946 , n784 , n26502 );
    nor g17743 ( n35474 , n7278 , n3804 );
    not g17744 ( n4854 , n499 );
    xnor g17745 ( n32452 , n3053 , n18492 );
    nor g17746 ( n30759 , n37801 , n21504 );
    or g17747 ( n37312 , n12779 , n3573 );
    or g17748 ( n31461 , n24682 , n8888 );
    nor g17749 ( n36564 , n227 , n24577 );
    or g17750 ( n3328 , n17509 , n12210 );
    and g17751 ( n24501 , n10882 , n31921 );
    xnor g17752 ( n18551 , n2799 , n13145 );
    not g17753 ( n7169 , n2914 );
    or g17754 ( n20110 , n31261 , n26604 );
    or g17755 ( n39308 , n30829 , n23385 );
    not g17756 ( n27683 , n31122 );
    and g17757 ( n24416 , n28334 , n15716 );
    and g17758 ( n27444 , n36122 , n3628 );
    xnor g17759 ( n9065 , n37210 , n12926 );
    xnor g17760 ( n9638 , n2005 , n9128 );
    and g17761 ( n39042 , n27704 , n29041 );
    or g17762 ( n40258 , n4173 , n34475 );
    or g17763 ( n3073 , n40455 , n32754 );
    or g17764 ( n32530 , n39686 , n30828 );
    or g17765 ( n3082 , n34887 , n8485 );
    not g17766 ( n1073 , n6340 );
    and g17767 ( n12290 , n11150 , n23070 );
    nor g17768 ( n37225 , n34831 , n36263 );
    and g17769 ( n31680 , n31240 , n42498 );
    not g17770 ( n25118 , n26268 );
    or g17771 ( n15633 , n7807 , n13318 );
    or g17772 ( n18129 , n19771 , n25078 );
    xnor g17773 ( n36042 , n965 , n14317 );
    or g17774 ( n11882 , n14068 , n1086 );
    not g17775 ( n5522 , n28150 );
    or g17776 ( n31262 , n22626 , n34511 );
    or g17777 ( n2700 , n17119 , n39758 );
    or g17778 ( n27759 , n23884 , n29707 );
    xnor g17779 ( n13791 , n38081 , n12616 );
    or g17780 ( n3300 , n10953 , n5712 );
    nor g17781 ( n24575 , n18866 , n14000 );
    xnor g17782 ( n5221 , n5891 , n10940 );
    and g17783 ( n4177 , n18108 , n10394 );
    or g17784 ( n40968 , n5373 , n26729 );
    or g17785 ( n8458 , n19020 , n10846 );
    or g17786 ( n24427 , n11349 , n10897 );
    or g17787 ( n15698 , n35296 , n2597 );
    not g17788 ( n1153 , n20761 );
    or g17789 ( n24235 , n41439 , n3476 );
    not g17790 ( n42433 , n12901 );
    not g17791 ( n17587 , n21016 );
    and g17792 ( n9455 , n42346 , n40050 );
    or g17793 ( n4840 , n35578 , n8233 );
    nor g17794 ( n13058 , n16598 , n33473 );
    xnor g17795 ( n39978 , n6625 , n10488 );
    xnor g17796 ( n42244 , n20487 , n6252 );
    or g17797 ( n973 , n21372 , n11205 );
    not g17798 ( n9932 , n31638 );
    or g17799 ( n20309 , n41326 , n18536 );
    and g17800 ( n31892 , n34411 , n8495 );
    not g17801 ( n28284 , n22303 );
    xnor g17802 ( n41402 , n37235 , n8042 );
    nor g17803 ( n35567 , n30742 , n7742 );
    and g17804 ( n28216 , n14176 , n42865 );
    xnor g17805 ( n2382 , n15081 , n31536 );
    or g17806 ( n24916 , n39551 , n23340 );
    nor g17807 ( n38111 , n32534 , n24537 );
    not g17808 ( n12419 , n33646 );
    or g17809 ( n34125 , n40616 , n19283 );
    xnor g17810 ( n3331 , n1855 , n26208 );
    and g17811 ( n2404 , n20491 , n31740 );
    and g17812 ( n1670 , n13966 , n7974 );
    nor g17813 ( n13426 , n38324 , n33165 );
    and g17814 ( n9461 , n17751 , n39866 );
    or g17815 ( n41137 , n15106 , n13830 );
    or g17816 ( n38988 , n5273 , n3031 );
    and g17817 ( n26177 , n16374 , n42680 );
    not g17818 ( n14948 , n15677 );
    or g17819 ( n38045 , n14434 , n4688 );
    xnor g17820 ( n3930 , n29423 , n7216 );
    or g17821 ( n9260 , n18183 , n12179 );
    not g17822 ( n3447 , n15166 );
    nor g17823 ( n41907 , n8494 , n41126 );
    and g17824 ( n17747 , n11123 , n36933 );
    nor g17825 ( n13291 , n27762 , n6723 );
    and g17826 ( n34208 , n6166 , n32071 );
    not g17827 ( n2194 , n15191 );
    or g17828 ( n38012 , n25496 , n26801 );
    and g17829 ( n8479 , n33136 , n29321 );
    or g17830 ( n28145 , n33068 , n19746 );
    or g17831 ( n3839 , n8353 , n14923 );
    or g17832 ( n32462 , n40345 , n28229 );
    and g17833 ( n42733 , n17889 , n38680 );
    xnor g17834 ( n15373 , n11982 , n7137 );
    not g17835 ( n5312 , n743 );
    or g17836 ( n15300 , n20660 , n23895 );
    and g17837 ( n8536 , n29366 , n11831 );
    xnor g17838 ( n24045 , n37829 , n30010 );
    nor g17839 ( n22413 , n38621 , n13421 );
    and g17840 ( n10691 , n41365 , n18309 );
    nor g17841 ( n26198 , n2375 , n15728 );
    and g17842 ( n15238 , n9131 , n18586 );
    or g17843 ( n39780 , n3801 , n6464 );
    or g17844 ( n41185 , n15105 , n33867 );
    xnor g17845 ( n40658 , n36009 , n38405 );
    or g17846 ( n23419 , n19450 , n10491 );
    or g17847 ( n27609 , n38438 , n25707 );
    not g17848 ( n8453 , n37811 );
    or g17849 ( n6320 , n40350 , n777 );
    and g17850 ( n14756 , n38873 , n25796 );
    xnor g17851 ( n17319 , n11596 , n38570 );
    not g17852 ( n734 , n13373 );
    and g17853 ( n28207 , n3289 , n21714 );
    or g17854 ( n3721 , n20345 , n33746 );
    or g17855 ( n9704 , n41266 , n7477 );
    nor g17856 ( n13619 , n16505 , n18808 );
    and g17857 ( n41485 , n22539 , n25512 );
    or g17858 ( n30049 , n32748 , n32800 );
    not g17859 ( n14013 , n41951 );
    xnor g17860 ( n23507 , n30429 , n42733 );
    or g17861 ( n25112 , n18822 , n10045 );
    and g17862 ( n37566 , n1771 , n33739 );
    not g17863 ( n37952 , n12805 );
    nor g17864 ( n11031 , n25817 , n2939 );
    or g17865 ( n10660 , n32215 , n4660 );
    and g17866 ( n37656 , n37314 , n26837 );
    or g17867 ( n41886 , n15096 , n38640 );
    nor g17868 ( n1422 , n15620 , n41703 );
    and g17869 ( n29349 , n24802 , n35415 );
    or g17870 ( n2443 , n29864 , n29968 );
    nor g17871 ( n22651 , n1110 , n42073 );
    not g17872 ( n29892 , n4517 );
    xnor g17873 ( n18895 , n23869 , n24748 );
    not g17874 ( n28120 , n11353 );
    and g17875 ( n22814 , n37511 , n32882 );
    and g17876 ( n40515 , n23327 , n37251 );
    not g17877 ( n32938 , n6196 );
    and g17878 ( n38576 , n33701 , n5394 );
    not g17879 ( n19002 , n29711 );
    or g17880 ( n22125 , n17988 , n42265 );
    or g17881 ( n24219 , n40295 , n29015 );
    or g17882 ( n40095 , n14471 , n24979 );
    nor g17883 ( n6101 , n40210 , n30600 );
    or g17884 ( n27652 , n9813 , n25343 );
    xnor g17885 ( n8399 , n2998 , n22226 );
    and g17886 ( n22543 , n16571 , n17366 );
    not g17887 ( n29143 , n17247 );
    not g17888 ( n1009 , n35225 );
    or g17889 ( n18773 , n32542 , n31771 );
    or g17890 ( n21001 , n25742 , n25032 );
    not g17891 ( n32683 , n32105 );
    and g17892 ( n4256 , n6235 , n9166 );
    or g17893 ( n15944 , n40300 , n25616 );
    not g17894 ( n37478 , n20416 );
    nor g17895 ( n6258 , n22086 , n27934 );
    not g17896 ( n11051 , n15693 );
    and g17897 ( n40186 , n37766 , n24888 );
    or g17898 ( n33346 , n35348 , n27089 );
    nor g17899 ( n24877 , n4591 , n210 );
    xnor g17900 ( n22059 , n11436 , n37724 );
    and g17901 ( n42691 , n39673 , n31715 );
    or g17902 ( n19175 , n16848 , n28006 );
    not g17903 ( n31510 , n17738 );
    not g17904 ( n16618 , n20075 );
    or g17905 ( n39820 , n42045 , n26747 );
    not g17906 ( n9252 , n28921 );
    or g17907 ( n28626 , n5175 , n19009 );
    nor g17908 ( n18484 , n29481 , n6692 );
    or g17909 ( n24983 , n35320 , n37791 );
    or g17910 ( n23770 , n39730 , n14032 );
    xnor g17911 ( n36202 , n31989 , n24007 );
    or g17912 ( n41151 , n28796 , n37825 );
    or g17913 ( n12578 , n3806 , n1947 );
    or g17914 ( n22460 , n35193 , n22524 );
    not g17915 ( n16942 , n26595 );
    or g17916 ( n36289 , n32800 , n19986 );
    not g17917 ( n34389 , n20333 );
    not g17918 ( n22296 , n10962 );
    nor g17919 ( n42334 , n2686 , n28284 );
    and g17920 ( n33486 , n33067 , n4805 );
    xnor g17921 ( n20062 , n19385 , n9406 );
    or g17922 ( n2446 , n17229 , n31603 );
    or g17923 ( n6931 , n37566 , n41079 );
    nor g17924 ( n1889 , n23618 , n16430 );
    not g17925 ( n9743 , n9462 );
    not g17926 ( n402 , n26591 );
    and g17927 ( n22868 , n12595 , n37608 );
    or g17928 ( n12273 , n21336 , n495 );
    nor g17929 ( n40616 , n41534 , n35131 );
    or g17930 ( n37227 , n7404 , n1026 );
    not g17931 ( n22103 , n19485 );
    or g17932 ( n31253 , n36524 , n31091 );
    not g17933 ( n42505 , n34159 );
    and g17934 ( n26973 , n11933 , n39381 );
    xnor g17935 ( n7399 , n20548 , n11230 );
    xnor g17936 ( n6406 , n14105 , n27326 );
    or g17937 ( n5950 , n16939 , n16981 );
    not g17938 ( n35691 , n36024 );
    or g17939 ( n15831 , n8913 , n15705 );
    and g17940 ( n42173 , n28306 , n17734 );
    or g17941 ( n20808 , n13631 , n35795 );
    or g17942 ( n18941 , n17386 , n25355 );
    and g17943 ( n30412 , n37786 , n886 );
    not g17944 ( n24231 , n12451 );
    not g17945 ( n38314 , n27308 );
    nor g17946 ( n6284 , n16143 , n38255 );
    or g17947 ( n1157 , n38168 , n24755 );
    nor g17948 ( n9645 , n13913 , n25219 );
    nor g17949 ( n12256 , n7356 , n25304 );
    nor g17950 ( n4515 , n36932 , n41387 );
    not g17951 ( n38335 , n25692 );
    not g17952 ( n27599 , n23557 );
    nor g17953 ( n12399 , n1186 , n11230 );
    or g17954 ( n16144 , n23462 , n32699 );
    and g17955 ( n10473 , n5898 , n14171 );
    and g17956 ( n6480 , n6843 , n7733 );
    xnor g17957 ( n19108 , n25619 , n17559 );
    xnor g17958 ( n37729 , n38749 , n29585 );
    xnor g17959 ( n26200 , n34562 , n23174 );
    xnor g17960 ( n14037 , n18880 , n15294 );
    and g17961 ( n16882 , n2687 , n42446 );
    nor g17962 ( n1268 , n5959 , n37675 );
    and g17963 ( n17847 , n2674 , n32784 );
    and g17964 ( n28420 , n16305 , n16898 );
    and g17965 ( n42144 , n11212 , n8326 );
    or g17966 ( n5273 , n21249 , n24817 );
    and g17967 ( n30859 , n33928 , n9188 );
    and g17968 ( n34589 , n32461 , n10003 );
    or g17969 ( n39313 , n6703 , n42722 );
    or g17970 ( n7248 , n39757 , n35990 );
    not g17971 ( n10592 , n37478 );
    not g17972 ( n25978 , n34076 );
    or g17973 ( n12934 , n12657 , n29673 );
    nor g17974 ( n36293 , n4140 , n18929 );
    not g17975 ( n4542 , n10792 );
    and g17976 ( n38441 , n19932 , n25224 );
    or g17977 ( n26135 , n35866 , n28750 );
    and g17978 ( n20846 , n28374 , n411 );
    nor g17979 ( n1032 , n17319 , n36609 );
    or g17980 ( n3880 , n25588 , n5660 );
    or g17981 ( n16777 , n38614 , n39888 );
    or g17982 ( n23551 , n31452 , n19336 );
    xnor g17983 ( n30769 , n24588 , n36535 );
    or g17984 ( n28460 , n30320 , n25168 );
    nor g17985 ( n20756 , n2840 , n7760 );
    not g17986 ( n39642 , n5097 );
    or g17987 ( n1945 , n30806 , n32543 );
    nor g17988 ( n804 , n8494 , n9887 );
    or g17989 ( n25026 , n6632 , n36747 );
    not g17990 ( n33328 , n17130 );
    and g17991 ( n14787 , n17689 , n1132 );
    or g17992 ( n29516 , n665 , n31953 );
    not g17993 ( n24148 , n34459 );
    xnor g17994 ( n7963 , n22799 , n32770 );
    nor g17995 ( n40221 , n17193 , n23103 );
    or g17996 ( n9340 , n27730 , n17066 );
    or g17997 ( n24166 , n33743 , n42551 );
    not g17998 ( n1326 , n25756 );
    and g17999 ( n12177 , n32591 , n35494 );
    or g18000 ( n4703 , n18165 , n15026 );
    or g18001 ( n21137 , n40363 , n40350 );
    not g18002 ( n9988 , n35922 );
    and g18003 ( n16915 , n30873 , n41077 );
    not g18004 ( n39200 , n25025 );
    not g18005 ( n25853 , n3366 );
    and g18006 ( n29700 , n17645 , n31020 );
    and g18007 ( n28363 , n38304 , n15650 );
    or g18008 ( n3495 , n33480 , n18174 );
    nor g18009 ( n30872 , n18854 , n35542 );
    or g18010 ( n20641 , n41111 , n32186 );
    nor g18011 ( n22687 , n11847 , n40944 );
    xnor g18012 ( n38419 , n105 , n28731 );
    or g18013 ( n25093 , n67 , n14563 );
    not g18014 ( n25957 , n9205 );
    or g18015 ( n14605 , n14793 , n143 );
    not g18016 ( n6583 , n3730 );
    xnor g18017 ( n25442 , n13798 , n38291 );
    or g18018 ( n21344 , n36585 , n34228 );
    nor g18019 ( n17730 , n25041 , n8495 );
    or g18020 ( n2828 , n38822 , n39354 );
    xnor g18021 ( n41370 , n11852 , n20596 );
    not g18022 ( n2358 , n13409 );
    and g18023 ( n22761 , n11333 , n2220 );
    or g18024 ( n14147 , n6480 , n13547 );
    nor g18025 ( n35069 , n33620 , n39039 );
    not g18026 ( n34562 , n17275 );
    or g18027 ( n9422 , n13102 , n42603 );
    nor g18028 ( n12858 , n1531 , n40682 );
    nor g18029 ( n33970 , n39598 , n16710 );
    and g18030 ( n20359 , n21917 , n16050 );
    and g18031 ( n18104 , n42468 , n32528 );
    and g18032 ( n37565 , n32454 , n27013 );
    not g18033 ( n15095 , n8066 );
    and g18034 ( n3910 , n9578 , n2187 );
    or g18035 ( n5507 , n28021 , n15005 );
    nor g18036 ( n9395 , n3906 , n8277 );
    not g18037 ( n11633 , n2093 );
    and g18038 ( n38166 , n7489 , n31134 );
    or g18039 ( n34380 , n21673 , n31997 );
    or g18040 ( n37963 , n8401 , n31711 );
    or g18041 ( n13025 , n25964 , n11395 );
    and g18042 ( n7256 , n32196 , n4485 );
    not g18043 ( n42423 , n28296 );
    or g18044 ( n8829 , n10086 , n1995 );
    nor g18045 ( n37788 , n29782 , n17362 );
    xnor g18046 ( n1365 , n22484 , n22288 );
    nor g18047 ( n3915 , n5964 , n17844 );
    or g18048 ( n33271 , n1974 , n5110 );
    nor g18049 ( n40033 , n29882 , n37823 );
    xnor g18050 ( n41628 , n10157 , n27307 );
    not g18051 ( n4574 , n19521 );
    or g18052 ( n3779 , n23921 , n17530 );
    not g18053 ( n263 , n31267 );
    and g18054 ( n9205 , n23483 , n41935 );
    or g18055 ( n38707 , n40909 , n34267 );
    and g18056 ( n20305 , n18064 , n16651 );
    or g18057 ( n2792 , n20613 , n41413 );
    or g18058 ( n4818 , n38117 , n34184 );
    xnor g18059 ( n3979 , n40 , n15795 );
    or g18060 ( n17653 , n34796 , n19421 );
    or g18061 ( n42163 , n42786 , n34107 );
    not g18062 ( n14962 , n32526 );
    and g18063 ( n39911 , n41446 , n4695 );
    and g18064 ( n12063 , n16767 , n16646 );
    and g18065 ( n42655 , n33148 , n11289 );
    and g18066 ( n715 , n1093 , n35433 );
    not g18067 ( n34224 , n5145 );
    and g18068 ( n19308 , n956 , n11372 );
    not g18069 ( n42740 , n31440 );
    or g18070 ( n27074 , n29930 , n41509 );
    and g18071 ( n38601 , n7766 , n40858 );
    or g18072 ( n26072 , n31728 , n33029 );
    and g18073 ( n32771 , n31500 , n16068 );
    nor g18074 ( n4148 , n26579 , n16567 );
    not g18075 ( n39066 , n717 );
    not g18076 ( n31489 , n22712 );
    not g18077 ( n1615 , n40772 );
    nor g18078 ( n16349 , n3036 , n30932 );
    or g18079 ( n19542 , n7492 , n33812 );
    xnor g18080 ( n19876 , n36046 , n11641 );
    not g18081 ( n41082 , n10412 );
    and g18082 ( n34754 , n13510 , n28751 );
    or g18083 ( n35704 , n33581 , n22064 );
    nor g18084 ( n40805 , n7197 , n5434 );
    not g18085 ( n33385 , n28251 );
    not g18086 ( n10084 , n20737 );
    or g18087 ( n14773 , n3892 , n28241 );
    or g18088 ( n31709 , n16780 , n9928 );
    or g18089 ( n30449 , n15486 , n34858 );
    or g18090 ( n27209 , n37242 , n7838 );
    or g18091 ( n32300 , n42076 , n29770 );
    or g18092 ( n39770 , n34391 , n9934 );
    and g18093 ( n6507 , n14981 , n2945 );
    or g18094 ( n6804 , n33538 , n23421 );
    not g18095 ( n16244 , n19631 );
    nor g18096 ( n7573 , n16431 , n40680 );
    or g18097 ( n20512 , n12448 , n18427 );
    or g18098 ( n39867 , n29817 , n11484 );
    or g18099 ( n1684 , n40472 , n17940 );
    xnor g18100 ( n8059 , n35887 , n5210 );
    and g18101 ( n12535 , n39351 , n25158 );
    or g18102 ( n41585 , n2608 , n21264 );
    and g18103 ( n36796 , n42193 , n30528 );
    or g18104 ( n41884 , n31635 , n23959 );
    not g18105 ( n12706 , n8081 );
    xnor g18106 ( n31633 , n31989 , n42180 );
    not g18107 ( n10898 , n17598 );
    xnor g18108 ( n8871 , n36970 , n22679 );
    and g18109 ( n10595 , n7514 , n9109 );
    xnor g18110 ( n33584 , n36423 , n37628 );
    not g18111 ( n34361 , n15995 );
    or g18112 ( n2534 , n4088 , n10337 );
    not g18113 ( n2095 , n39487 );
    and g18114 ( n28483 , n37529 , n4053 );
    or g18115 ( n40558 , n25509 , n16501 );
    and g18116 ( n13654 , n17744 , n31296 );
    not g18117 ( n10859 , n9002 );
    or g18118 ( n625 , n39257 , n23793 );
    and g18119 ( n28731 , n34526 , n11296 );
    or g18120 ( n1512 , n23859 , n15588 );
    not g18121 ( n10845 , n12630 );
    and g18122 ( n36600 , n14753 , n34736 );
    not g18123 ( n6858 , n33959 );
    or g18124 ( n5062 , n35528 , n26757 );
    or g18125 ( n789 , n36272 , n42543 );
    and g18126 ( n36381 , n6444 , n33979 );
    or g18127 ( n26333 , n3275 , n8333 );
    xnor g18128 ( n680 , n37644 , n23813 );
    nor g18129 ( n39251 , n31378 , n38374 );
    nor g18130 ( n16997 , n22484 , n31907 );
    and g18131 ( n5280 , n5642 , n35602 );
    and g18132 ( n38407 , n23697 , n2541 );
    and g18133 ( n25221 , n37597 , n35623 );
    or g18134 ( n35059 , n31900 , n10290 );
    not g18135 ( n4018 , n16079 );
    or g18136 ( n29494 , n42547 , n20574 );
    not g18137 ( n26861 , n25645 );
    nor g18138 ( n5094 , n7421 , n26780 );
    not g18139 ( n13182 , n13103 );
    nor g18140 ( n9734 , n34415 , n28407 );
    or g18141 ( n3967 , n13701 , n21103 );
    and g18142 ( n33746 , n15532 , n5968 );
    or g18143 ( n3638 , n28869 , n1326 );
    or g18144 ( n34457 , n3247 , n40178 );
    xnor g18145 ( n11846 , n105 , n33468 );
    or g18146 ( n37325 , n12144 , n27274 );
    nor g18147 ( n12101 , n8300 , n38936 );
    nor g18148 ( n26166 , n9864 , n33308 );
    or g18149 ( n16629 , n14944 , n37984 );
    and g18150 ( n12232 , n17790 , n39006 );
    or g18151 ( n7264 , n35914 , n2152 );
    and g18152 ( n33451 , n38762 , n18831 );
    and g18153 ( n38132 , n8225 , n6594 );
    or g18154 ( n3388 , n39972 , n34559 );
    or g18155 ( n15308 , n23591 , n7365 );
    and g18156 ( n27546 , n4845 , n5878 );
    or g18157 ( n41012 , n11404 , n24238 );
    nor g18158 ( n1207 , n5964 , n40339 );
    and g18159 ( n35510 , n21190 , n16056 );
    not g18160 ( n36393 , n41758 );
    nor g18161 ( n26372 , n1782 , n4859 );
    not g18162 ( n23857 , n29131 );
    and g18163 ( n3135 , n22227 , n28781 );
    not g18164 ( n29646 , n18247 );
    or g18165 ( n13439 , n14423 , n32867 );
    and g18166 ( n36717 , n41432 , n16291 );
    not g18167 ( n25178 , n24466 );
    not g18168 ( n3583 , n37540 );
    not g18169 ( n25630 , n12332 );
    or g18170 ( n9324 , n34793 , n20558 );
    nor g18171 ( n13534 , n12430 , n36877 );
    not g18172 ( n17946 , n34302 );
    or g18173 ( n26014 , n36546 , n32633 );
    and g18174 ( n16893 , n10883 , n26920 );
    and g18175 ( n36155 , n6847 , n5014 );
    or g18176 ( n9831 , n22925 , n33464 );
    or g18177 ( n22878 , n36755 , n19182 );
    or g18178 ( n11505 , n13816 , n6195 );
    nor g18179 ( n30527 , n11201 , n24214 );
    not g18180 ( n22109 , n25893 );
    nor g18181 ( n26518 , n7987 , n31443 );
    nor g18182 ( n40819 , n22918 , n18479 );
    nor g18183 ( n38241 , n2199 , n38297 );
    or g18184 ( n14768 , n21641 , n27612 );
    xnor g18185 ( n33548 , n34444 , n6013 );
    nor g18186 ( n4017 , n2191 , n3979 );
    xnor g18187 ( n27881 , n14658 , n37751 );
    nor g18188 ( n23440 , n39923 , n9120 );
    and g18189 ( n25970 , n7318 , n9407 );
    and g18190 ( n12729 , n27290 , n19901 );
    nor g18191 ( n40946 , n17647 , n19682 );
    and g18192 ( n12687 , n9115 , n10442 );
    or g18193 ( n14702 , n13143 , n17249 );
    or g18194 ( n20300 , n23509 , n16846 );
    xnor g18195 ( n23837 , n21534 , n31307 );
    nor g18196 ( n29101 , n2199 , n22945 );
    and g18197 ( n26386 , n26923 , n35788 );
    or g18198 ( n35836 , n12243 , n12669 );
    or g18199 ( n27348 , n23563 , n38008 );
    not g18200 ( n36218 , n30020 );
    not g18201 ( n34626 , n41578 );
    or g18202 ( n34077 , n33802 , n37925 );
    or g18203 ( n11437 , n32106 , n29167 );
    and g18204 ( n32285 , n19286 , n40155 );
    or g18205 ( n26990 , n37665 , n14621 );
    and g18206 ( n29241 , n41481 , n12604 );
    or g18207 ( n3565 , n4594 , n26409 );
    nor g18208 ( n2438 , n13690 , n23567 );
    or g18209 ( n21799 , n38035 , n37015 );
    and g18210 ( n18031 , n36756 , n35389 );
    and g18211 ( n24650 , n25574 , n1156 );
    and g18212 ( n42569 , n31260 , n17089 );
    not g18213 ( n35604 , n36853 );
    nor g18214 ( n23073 , n28333 , n33923 );
    nor g18215 ( n20269 , n11730 , n18153 );
    nor g18216 ( n1205 , n3769 , n41163 );
    or g18217 ( n35121 , n29963 , n22222 );
    nor g18218 ( n16984 , n299 , n39886 );
    and g18219 ( n38066 , n36918 , n27559 );
    or g18220 ( n32267 , n18165 , n37956 );
    or g18221 ( n27514 , n25811 , n31175 );
    nor g18222 ( n10018 , n1507 , n12354 );
    not g18223 ( n29796 , n12514 );
    nor g18224 ( n19791 , n19835 , n35693 );
    or g18225 ( n23142 , n37588 , n10604 );
    not g18226 ( n13161 , n19387 );
    nor g18227 ( n29927 , n35522 , n33224 );
    or g18228 ( n28454 , n42801 , n6294 );
    or g18229 ( n35 , n36235 , n10042 );
    or g18230 ( n26831 , n9023 , n37793 );
    or g18231 ( n6830 , n19653 , n26223 );
    or g18232 ( n41846 , n14471 , n37894 );
    nor g18233 ( n10345 , n18512 , n25861 );
    nor g18234 ( n37727 , n16379 , n24116 );
    not g18235 ( n9177 , n22980 );
    xnor g18236 ( n21193 , n37175 , n2777 );
    and g18237 ( n31267 , n35230 , n42266 );
    not g18238 ( n39635 , n294 );
    and g18239 ( n33491 , n17546 , n3027 );
    nor g18240 ( n14997 , n10799 , n23429 );
    xnor g18241 ( n22121 , n7621 , n6119 );
    xnor g18242 ( n11848 , n29796 , n15014 );
    or g18243 ( n33123 , n12735 , n23456 );
    nor g18244 ( n6124 , n14471 , n15719 );
    and g18245 ( n668 , n41463 , n37593 );
    or g18246 ( n27083 , n28672 , n34117 );
    and g18247 ( n24808 , n1236 , n24676 );
    or g18248 ( n24370 , n28745 , n24684 );
    and g18249 ( n6881 , n23830 , n17106 );
    or g18250 ( n16307 , n21747 , n35382 );
    or g18251 ( n25332 , n31550 , n4328 );
    xnor g18252 ( n39572 , n24428 , n36808 );
    and g18253 ( n36789 , n20432 , n13283 );
    or g18254 ( n6623 , n22345 , n3520 );
    not g18255 ( n12437 , n22628 );
    or g18256 ( n24930 , n41387 , n39098 );
    or g18257 ( n36695 , n6602 , n32108 );
    xnor g18258 ( n24997 , n36973 , n7354 );
    and g18259 ( n27950 , n18110 , n23415 );
    or g18260 ( n32903 , n8914 , n27057 );
    and g18261 ( n8630 , n31099 , n41013 );
    not g18262 ( n39320 , n25323 );
    and g18263 ( n28076 , n32387 , n7334 );
    xnor g18264 ( n222 , n40771 , n22995 );
    xnor g18265 ( n11893 , n41013 , n16643 );
    xnor g18266 ( n36324 , n36365 , n3415 );
    and g18267 ( n5044 , n38843 , n5139 );
    nor g18268 ( n18838 , n24976 , n18359 );
    or g18269 ( n36229 , n23302 , n23017 );
    or g18270 ( n32145 , n12722 , n17311 );
    nor g18271 ( n833 , n31674 , n29542 );
    or g18272 ( n15427 , n27598 , n31727 );
    and g18273 ( n9308 , n9806 , n24946 );
    or g18274 ( n20689 , n17687 , n27459 );
    and g18275 ( n23286 , n2467 , n41096 );
    and g18276 ( n25281 , n10411 , n24672 );
    or g18277 ( n13915 , n28987 , n8442 );
    nor g18278 ( n4868 , n5064 , n20915 );
    or g18279 ( n10049 , n6866 , n17104 );
    or g18280 ( n12196 , n7020 , n9889 );
    nor g18281 ( n33825 , n33981 , n3091 );
    or g18282 ( n30946 , n34301 , n2221 );
    or g18283 ( n5698 , n40494 , n23386 );
    not g18284 ( n31957 , n39470 );
    nor g18285 ( n20507 , n15766 , n29739 );
    xnor g18286 ( n8002 , n14425 , n8456 );
    nor g18287 ( n22851 , n18212 , n21951 );
    or g18288 ( n17580 , n24243 , n36103 );
    nor g18289 ( n12426 , n3656 , n14983 );
    nor g18290 ( n32785 , n37257 , n28257 );
    nor g18291 ( n29766 , n19613 , n25671 );
    and g18292 ( n13467 , n25163 , n9119 );
    not g18293 ( n24108 , n29047 );
    or g18294 ( n23919 , n3580 , n8449 );
    xnor g18295 ( n20538 , n4659 , n27383 );
    or g18296 ( n29910 , n24070 , n21285 );
    or g18297 ( n12326 , n5896 , n20974 );
    not g18298 ( n41013 , n5896 );
    or g18299 ( n28546 , n7127 , n17754 );
    xnor g18300 ( n23486 , n9460 , n9461 );
    nor g18301 ( n18010 , n5400 , n18054 );
    and g18302 ( n19004 , n34347 , n5078 );
    nor g18303 ( n2774 , n27394 , n3243 );
    nor g18304 ( n34331 , n28872 , n37641 );
    or g18305 ( n27641 , n16967 , n10751 );
    not g18306 ( n9792 , n26903 );
    or g18307 ( n14270 , n1538 , n14072 );
    nor g18308 ( n29250 , n2183 , n9680 );
    xnor g18309 ( n19382 , n37953 , n4088 );
    and g18310 ( n19240 , n23658 , n3458 );
    or g18311 ( n18217 , n14074 , n15012 );
    or g18312 ( n41664 , n37312 , n37454 );
    or g18313 ( n26960 , n42748 , n35551 );
    nor g18314 ( n21112 , n9511 , n6437 );
    or g18315 ( n14415 , n1058 , n3335 );
    and g18316 ( n41928 , n23278 , n37937 );
    not g18317 ( n1863 , n1903 );
    or g18318 ( n19415 , n24692 , n24675 );
    or g18319 ( n2024 , n29288 , n10045 );
    nor g18320 ( n27532 , n34565 , n40984 );
    and g18321 ( n13414 , n6539 , n2978 );
    and g18322 ( n34170 , n30512 , n36959 );
    not g18323 ( n35083 , n26692 );
    or g18324 ( n14256 , n21023 , n36851 );
    or g18325 ( n24773 , n620 , n6290 );
    and g18326 ( n27908 , n24486 , n29022 );
    or g18327 ( n16794 , n38973 , n9344 );
    not g18328 ( n32410 , n7069 );
    and g18329 ( n12122 , n34321 , n15929 );
    or g18330 ( n34518 , n18873 , n9994 );
    or g18331 ( n25580 , n39636 , n24482 );
    and g18332 ( n19691 , n8305 , n19524 );
    nor g18333 ( n7896 , n28710 , n35417 );
    and g18334 ( n10544 , n11701 , n37676 );
    or g18335 ( n8720 , n16967 , n22517 );
    and g18336 ( n38123 , n38377 , n1228 );
    and g18337 ( n15547 , n38099 , n28626 );
    and g18338 ( n22007 , n22093 , n27118 );
    not g18339 ( n35377 , n40301 );
    or g18340 ( n9393 , n19969 , n9658 );
    and g18341 ( n38776 , n28879 , n10038 );
    or g18342 ( n25868 , n5814 , n41455 );
    nor g18343 ( n10528 , n25860 , n21403 );
    not g18344 ( n19508 , n42915 );
    or g18345 ( n21927 , n1070 , n2022 );
    nor g18346 ( n27753 , n34292 , n15718 );
    and g18347 ( n3873 , n36881 , n42485 );
    nor g18348 ( n8000 , n14707 , n24022 );
    xnor g18349 ( n690 , n6625 , n20424 );
    xnor g18350 ( n4351 , n41013 , n24807 );
    and g18351 ( n1866 , n8091 , n15773 );
    or g18352 ( n30439 , n30030 , n22896 );
    xnor g18353 ( n23316 , n7282 , n14114 );
    or g18354 ( n29756 , n10229 , n31996 );
    or g18355 ( n42847 , n25316 , n30418 );
    nor g18356 ( n9475 , n32910 , n461 );
    and g18357 ( n19294 , n32934 , n32466 );
    or g18358 ( n19671 , n9923 , n34057 );
    or g18359 ( n8201 , n38548 , n8073 );
    or g18360 ( n21861 , n14851 , n1520 );
    and g18361 ( n684 , n22918 , n18479 );
    and g18362 ( n15208 , n27790 , n31065 );
    nor g18363 ( n36157 , n4388 , n3670 );
    nor g18364 ( n25621 , n26523 , n24783 );
    not g18365 ( n36731 , n39287 );
    or g18366 ( n23276 , n39237 , n39536 );
    not g18367 ( n23920 , n40456 );
    or g18368 ( n9950 , n41453 , n22635 );
    and g18369 ( n9876 , n15652 , n1008 );
    and g18370 ( n33557 , n672 , n3866 );
    or g18371 ( n7909 , n8539 , n28995 );
    or g18372 ( n20483 , n38218 , n29340 );
    xnor g18373 ( n6437 , n28415 , n12627 );
    or g18374 ( n2491 , n4872 , n15084 );
    xnor g18375 ( n24140 , n28852 , n26220 );
    nor g18376 ( n27980 , n28110 , n39530 );
    and g18377 ( n13040 , n14256 , n35642 );
    and g18378 ( n42221 , n1388 , n13802 );
    not g18379 ( n40852 , n23948 );
    or g18380 ( n42417 , n23292 , n12435 );
    or g18381 ( n21580 , n7201 , n15582 );
    or g18382 ( n29967 , n29243 , n863 );
    or g18383 ( n18302 , n7882 , n25110 );
    and g18384 ( n21054 , n39410 , n27048 );
    or g18385 ( n32501 , n21201 , n23035 );
    nor g18386 ( n36631 , n15736 , n29132 );
    and g18387 ( n25309 , n14747 , n23084 );
    or g18388 ( n13802 , n36880 , n24841 );
    not g18389 ( n1940 , n29912 );
    or g18390 ( n22185 , n35923 , n20448 );
    and g18391 ( n32136 , n36626 , n20528 );
    not g18392 ( n28443 , n31780 );
    and g18393 ( n7468 , n28601 , n5976 );
    not g18394 ( n19366 , n21643 );
    xnor g18395 ( n23049 , n38914 , n20976 );
    or g18396 ( n4977 , n6033 , n38437 );
    nor g18397 ( n25954 , n22086 , n28417 );
    and g18398 ( n12278 , n34717 , n35776 );
    xnor g18399 ( n29435 , n119 , n6723 );
    or g18400 ( n6185 , n5952 , n9456 );
    and g18401 ( n516 , n5041 , n27505 );
    and g18402 ( n38897 , n14593 , n19520 );
    not g18403 ( n21282 , n14965 );
    not g18404 ( n7027 , n23002 );
    or g18405 ( n26993 , n40801 , n19159 );
    not g18406 ( n2734 , n37364 );
    or g18407 ( n10866 , n18107 , n36235 );
    xnor g18408 ( n10709 , n34628 , n20431 );
    not g18409 ( n15289 , n40006 );
    and g18410 ( n19798 , n42197 , n38451 );
    and g18411 ( n12716 , n21739 , n13878 );
    or g18412 ( n37499 , n41586 , n8249 );
    or g18413 ( n31202 , n38588 , n22624 );
    xnor g18414 ( n9098 , n36009 , n11218 );
    or g18415 ( n13462 , n5324 , n5357 );
    and g18416 ( n32633 , n10884 , n10393 );
    or g18417 ( n39740 , n13411 , n23559 );
    xnor g18418 ( n1605 , n15281 , n1173 );
    not g18419 ( n11585 , n33198 );
    or g18420 ( n1827 , n39422 , n4552 );
    not g18421 ( n41345 , n3201 );
    or g18422 ( n29591 , n14200 , n1735 );
    and g18423 ( n9213 , n878 , n4902 );
    nor g18424 ( n31597 , n13181 , n18731 );
    or g18425 ( n459 , n24574 , n15352 );
    or g18426 ( n29466 , n29058 , n5518 );
    and g18427 ( n34007 , n15669 , n8106 );
    not g18428 ( n16700 , n3100 );
    or g18429 ( n4605 , n28125 , n25366 );
    or g18430 ( n26734 , n19672 , n26961 );
    or g18431 ( n35460 , n22270 , n5183 );
    or g18432 ( n16374 , n39817 , n14379 );
    not g18433 ( n30796 , n29036 );
    nor g18434 ( n33349 , n40757 , n41284 );
    not g18435 ( n21259 , n854 );
    not g18436 ( n23292 , n37451 );
    not g18437 ( n42513 , n38444 );
    or g18438 ( n7704 , n41891 , n7830 );
    nor g18439 ( n25295 , n18833 , n35634 );
    or g18440 ( n28655 , n33466 , n17512 );
    and g18441 ( n18976 , n10186 , n31870 );
    or g18442 ( n6649 , n37663 , n4843 );
    xnor g18443 ( n32379 , n26972 , n5044 );
    or g18444 ( n4082 , n16299 , n38585 );
    nor g18445 ( n24927 , n39456 , n39679 );
    not g18446 ( n18775 , n23689 );
    and g18447 ( n8117 , n38675 , n12899 );
    xnor g18448 ( n25660 , n2488 , n40515 );
    not g18449 ( n7616 , n40246 );
    not g18450 ( n16791 , n29926 );
    or g18451 ( n12561 , n41363 , n4355 );
    and g18452 ( n7830 , n11042 , n19078 );
    or g18453 ( n10826 , n34373 , n30312 );
    or g18454 ( n25484 , n35879 , n33666 );
    and g18455 ( n159 , n23029 , n30922 );
    or g18456 ( n21959 , n4447 , n24902 );
    and g18457 ( n21632 , n40841 , n6022 );
    or g18458 ( n5787 , n13337 , n27179 );
    not g18459 ( n41603 , n29560 );
    xnor g18460 ( n2717 , n35727 , n41567 );
    not g18461 ( n21807 , n39487 );
    and g18462 ( n9135 , n37124 , n24249 );
    and g18463 ( n27709 , n29267 , n9972 );
    not g18464 ( n41302 , n4292 );
    or g18465 ( n35580 , n29571 , n32786 );
    and g18466 ( n24123 , n13288 , n24430 );
    not g18467 ( n32384 , n9682 );
    or g18468 ( n39012 , n10701 , n14503 );
    and g18469 ( n2215 , n36294 , n30342 );
    not g18470 ( n42870 , n17205 );
    or g18471 ( n39322 , n36115 , n11059 );
    and g18472 ( n37944 , n10590 , n24966 );
    or g18473 ( n3986 , n30771 , n24483 );
    or g18474 ( n3294 , n17182 , n24227 );
    or g18475 ( n37474 , n36236 , n6458 );
    or g18476 ( n33327 , n38129 , n40367 );
    nor g18477 ( n30268 , n3502 , n1389 );
    not g18478 ( n14027 , n37544 );
    not g18479 ( n6950 , n14415 );
    not g18480 ( n3265 , n34922 );
    and g18481 ( n21571 , n5395 , n23255 );
    or g18482 ( n6499 , n9660 , n7579 );
    and g18483 ( n20321 , n41292 , n29925 );
    or g18484 ( n12453 , n11440 , n26068 );
    not g18485 ( n16333 , n26561 );
    xnor g18486 ( n2611 , n15277 , n5964 );
    nor g18487 ( n30063 , n1002 , n36139 );
    nor g18488 ( n25920 , n1507 , n13582 );
    xnor g18489 ( n7510 , n6625 , n17499 );
    or g18490 ( n5752 , n38249 , n41027 );
    nor g18491 ( n36098 , n28502 , n29547 );
    or g18492 ( n36495 , n2517 , n11719 );
    and g18493 ( n13371 , n34699 , n16547 );
    or g18494 ( n38885 , n23453 , n21172 );
    and g18495 ( n4506 , n17525 , n29931 );
    or g18496 ( n9681 , n13677 , n7856 );
    and g18497 ( n23635 , n15629 , n24886 );
    not g18498 ( n8783 , n29774 );
    or g18499 ( n23679 , n41021 , n7745 );
    or g18500 ( n34181 , n26935 , n22919 );
    nor g18501 ( n1525 , n38852 , n29595 );
    or g18502 ( n30500 , n29817 , n41645 );
    nor g18503 ( n12614 , n4869 , n38305 );
    nor g18504 ( n27743 , n9113 , n5199 );
    or g18505 ( n25081 , n12509 , n13535 );
    or g18506 ( n8749 , n31850 , n27823 );
    or g18507 ( n6463 , n30578 , n37594 );
    and g18508 ( n7845 , n11728 , n33640 );
    nor g18509 ( n41003 , n34292 , n4499 );
    or g18510 ( n22800 , n5995 , n10332 );
    or g18511 ( n12893 , n35320 , n41163 );
    or g18512 ( n9029 , n6290 , n9299 );
    not g18513 ( n4587 , n8066 );
    or g18514 ( n19711 , n4267 , n12011 );
    xnor g18515 ( n34574 , n30227 , n36805 );
    nor g18516 ( n32992 , n42049 , n41541 );
    nor g18517 ( n35878 , n40799 , n38274 );
    or g18518 ( n8016 , n19049 , n16241 );
    or g18519 ( n24833 , n40840 , n13329 );
    and g18520 ( n18330 , n20247 , n9478 );
    xnor g18521 ( n29635 , n5442 , n41465 );
    or g18522 ( n12080 , n35301 , n882 );
    nor g18523 ( n50 , n15961 , n11992 );
    not g18524 ( n19735 , n15978 );
    or g18525 ( n21793 , n23078 , n30234 );
    or g18526 ( n38189 , n28699 , n8318 );
    and g18527 ( n35959 , n3384 , n16895 );
    xnor g18528 ( n16895 , n16693 , n8151 );
    or g18529 ( n18803 , n14146 , n14115 );
    not g18530 ( n21610 , n7221 );
    or g18531 ( n28224 , n34042 , n20896 );
    not g18532 ( n10614 , n19119 );
    and g18533 ( n4901 , n5576 , n41217 );
    nor g18534 ( n6819 , n3581 , n15681 );
    not g18535 ( n24003 , n31629 );
    or g18536 ( n26303 , n39832 , n5568 );
    or g18537 ( n10968 , n17938 , n30914 );
    xnor g18538 ( n9355 , n26579 , n42280 );
    not g18539 ( n22825 , n26712 );
    or g18540 ( n32556 , n5911 , n37195 );
    and g18541 ( n16964 , n19328 , n16708 );
    not g18542 ( n17870 , n30949 );
    not g18543 ( n17510 , n35764 );
    or g18544 ( n38717 , n30498 , n15127 );
    or g18545 ( n6620 , n23739 , n27340 );
    or g18546 ( n6567 , n34626 , n40857 );
    or g18547 ( n11099 , n5978 , n1811 );
    nor g18548 ( n42536 , n31792 , n3190 );
    nor g18549 ( n23805 , n40752 , n25845 );
    or g18550 ( n8811 , n8206 , n25515 );
    nor g18551 ( n38646 , n5896 , n12417 );
    or g18552 ( n39877 , n33908 , n750 );
    not g18553 ( n28662 , n8093 );
    nor g18554 ( n8757 , n42003 , n19273 );
    nor g18555 ( n5052 , n39037 , n39675 );
    or g18556 ( n8838 , n2710 , n11 );
    and g18557 ( n10844 , n42116 , n4583 );
    or g18558 ( n27413 , n17744 , n29118 );
    and g18559 ( n38102 , n23441 , n42545 );
    or g18560 ( n4390 , n10650 , n35584 );
    not g18561 ( n15314 , n3369 );
    or g18562 ( n3393 , n6369 , n27787 );
    and g18563 ( n26914 , n31555 , n36699 );
    or g18564 ( n33729 , n8945 , n16999 );
    or g18565 ( n20542 , n32852 , n14380 );
    or g18566 ( n22990 , n31737 , n22892 );
    or g18567 ( n5260 , n35949 , n18070 );
    not g18568 ( n10496 , n11887 );
    or g18569 ( n5432 , n9176 , n32208 );
    and g18570 ( n41092 , n1325 , n41700 );
    and g18571 ( n41332 , n12918 , n1764 );
    or g18572 ( n38769 , n9778 , n21661 );
    or g18573 ( n26208 , n29528 , n1633 );
    not g18574 ( n21271 , n36315 );
    or g18575 ( n27266 , n15095 , n11676 );
    nor g18576 ( n10325 , n24010 , n3344 );
    or g18577 ( n28132 , n34127 , n38657 );
    xnor g18578 ( n20698 , n35727 , n1039 );
    and g18579 ( n18492 , n23091 , n4319 );
    or g18580 ( n33065 , n39118 , n40303 );
    or g18581 ( n9596 , n22220 , n12953 );
    or g18582 ( n14329 , n30948 , n19763 );
    and g18583 ( n24929 , n9232 , n16845 );
    nor g18584 ( n30703 , n22442 , n22321 );
    xnor g18585 ( n27590 , n20204 , n29840 );
    and g18586 ( n35880 , n22771 , n18932 );
    not g18587 ( n1879 , n12332 );
    xnor g18588 ( n5726 , n22263 , n26197 );
    or g18589 ( n23149 , n16836 , n32695 );
    and g18590 ( n15094 , n34760 , n40626 );
    or g18591 ( n27366 , n37671 , n16047 );
    or g18592 ( n19137 , n10493 , n34244 );
    not g18593 ( n18314 , n11713 );
    xnor g18594 ( n28147 , n9376 , n13862 );
    and g18595 ( n5431 , n24354 , n6114 );
    or g18596 ( n1084 , n5341 , n36306 );
    or g18597 ( n8379 , n22351 , n16093 );
    or g18598 ( n27858 , n27840 , n15793 );
    and g18599 ( n6773 , n26466 , n38114 );
    nor g18600 ( n9747 , n376 , n13352 );
    or g18601 ( n15036 , n40451 , n29915 );
    xnor g18602 ( n24443 , n21457 , n4368 );
    or g18603 ( n34722 , n39195 , n14997 );
    or g18604 ( n33747 , n33649 , n12220 );
    or g18605 ( n12188 , n33297 , n38103 );
    or g18606 ( n25305 , n23044 , n440 );
    or g18607 ( n15723 , n1735 , n36716 );
    not g18608 ( n31622 , n41742 );
    or g18609 ( n16254 , n5258 , n17407 );
    and g18610 ( n30200 , n28976 , n40382 );
    nor g18611 ( n21604 , n34992 , n22106 );
    nor g18612 ( n38473 , n37322 , n29769 );
    or g18613 ( n18855 , n40617 , n2601 );
    nor g18614 ( n13846 , n21520 , n40976 );
    or g18615 ( n32897 , n8108 , n12626 );
    and g18616 ( n40943 , n22655 , n22591 );
    not g18617 ( n24454 , n3000 );
    or g18618 ( n14880 , n11464 , n30056 );
    or g18619 ( n37658 , n28745 , n30311 );
    and g18620 ( n13043 , n10969 , n11963 );
    not g18621 ( n14149 , n9502 );
    xnor g18622 ( n5334 , n784 , n16354 );
    xnor g18623 ( n17977 , n13400 , n3909 );
    nor g18624 ( n10107 , n27844 , n5247 );
    nor g18625 ( n34806 , n5896 , n26982 );
    or g18626 ( n21353 , n28475 , n23576 );
    or g18627 ( n42459 , n10845 , n24530 );
    xnor g18628 ( n39052 , n16693 , n29240 );
    or g18629 ( n37486 , n3868 , n33089 );
    and g18630 ( n24010 , n36200 , n24501 );
    not g18631 ( n35509 , n25607 );
    or g18632 ( n35434 , n4144 , n40733 );
    and g18633 ( n10940 , n24094 , n39109 );
    and g18634 ( n3933 , n40502 , n23048 );
    and g18635 ( n23406 , n33833 , n32976 );
    and g18636 ( n20151 , n11633 , n8902 );
    xnor g18637 ( n16057 , n13236 , n4814 );
    nor g18638 ( n35120 , n40128 , n21203 );
    not g18639 ( n26064 , n20797 );
    or g18640 ( n18430 , n15780 , n6643 );
    or g18641 ( n28824 , n25726 , n19317 );
    or g18642 ( n25534 , n3640 , n19701 );
    or g18643 ( n20319 , n31810 , n13226 );
    not g18644 ( n4926 , n2814 );
    nor g18645 ( n23983 , n14077 , n13995 );
    xnor g18646 ( n9283 , n28808 , n35555 );
    nor g18647 ( n28555 , n39456 , n32830 );
    and g18648 ( n36473 , n20647 , n38930 );
    and g18649 ( n31027 , n22451 , n38141 );
    not g18650 ( n41913 , n13668 );
    not g18651 ( n34498 , n32545 );
    or g18652 ( n28194 , n16910 , n33440 );
    or g18653 ( n21335 , n30616 , n24119 );
    not g18654 ( n28411 , n41430 );
    and g18655 ( n30432 , n9097 , n33168 );
    nor g18656 ( n3936 , n19054 , n1281 );
    or g18657 ( n4460 , n1440 , n25528 );
    xnor g18658 ( n23403 , n378 , n18882 );
    and g18659 ( n13179 , n37949 , n11948 );
    xnor g18660 ( n24913 , n27245 , n10269 );
    and g18661 ( n8451 , n23329 , n39548 );
    and g18662 ( n1083 , n34564 , n27620 );
    or g18663 ( n35334 , n17581 , n13700 );
    nor g18664 ( n11282 , n22820 , n20729 );
    not g18665 ( n37671 , n3465 );
    or g18666 ( n22326 , n19376 , n9508 );
    or g18667 ( n12185 , n1010 , n16335 );
    or g18668 ( n26323 , n20443 , n15215 );
    or g18669 ( n6771 , n9329 , n35333 );
    and g18670 ( n18901 , n10901 , n34038 );
    or g18671 ( n15764 , n12119 , n30735 );
    and g18672 ( n16718 , n18454 , n41775 );
    nor g18673 ( n29621 , n14941 , n6734 );
    xnor g18674 ( n25394 , n9959 , n34372 );
    nor g18675 ( n33283 , n10517 , n13276 );
    and g18676 ( n41342 , n26676 , n24668 );
    or g18677 ( n37265 , n23993 , n1970 );
    or g18678 ( n27486 , n38463 , n2545 );
    or g18679 ( n18077 , n6635 , n19549 );
    nor g18680 ( n13892 , n28682 , n9647 );
    xnor g18681 ( n9287 , n10005 , n39521 );
    and g18682 ( n35923 , n28770 , n41146 );
    or g18683 ( n13816 , n19969 , n15516 );
    or g18684 ( n18539 , n21047 , n36514 );
    xnor g18685 ( n30673 , n4334 , n42023 );
    not g18686 ( n29735 , n39469 );
    not g18687 ( n437 , n41733 );
    or g18688 ( n26727 , n486 , n34569 );
    not g18689 ( n25148 , n11944 );
    or g18690 ( n37754 , n11247 , n13868 );
    or g18691 ( n40826 , n17313 , n17927 );
    or g18692 ( n12364 , n30802 , n38463 );
    or g18693 ( n42398 , n7384 , n14577 );
    not g18694 ( n10005 , n31626 );
    not g18695 ( n6196 , n12068 );
    and g18696 ( n11648 , n33003 , n40436 );
    xnor g18697 ( n18956 , n21321 , n6498 );
    and g18698 ( n14968 , n8267 , n24929 );
    nor g18699 ( n38 , n16598 , n15974 );
    nor g18700 ( n30085 , n2254 , n24424 );
    or g18701 ( n13323 , n4532 , n39120 );
    not g18702 ( n8495 , n34311 );
    xnor g18703 ( n17842 , n21525 , n38285 );
    or g18704 ( n29895 , n29122 , n37763 );
    or g18705 ( n8166 , n33624 , n27551 );
    and g18706 ( n37603 , n20134 , n27985 );
    or g18707 ( n16873 , n38512 , n41943 );
    or g18708 ( n1592 , n4308 , n17638 );
    not g18709 ( n14508 , n2238 );
    nor g18710 ( n20712 , n36667 , n15963 );
    or g18711 ( n29279 , n20503 , n18091 );
    or g18712 ( n2782 , n251 , n41780 );
    or g18713 ( n41039 , n41739 , n9942 );
    or g18714 ( n5093 , n30067 , n21703 );
    not g18715 ( n18453 , n30808 );
    and g18716 ( n40824 , n26612 , n7521 );
    or g18717 ( n28133 , n29306 , n32398 );
    xnor g18718 ( n36474 , n17056 , n16346 );
    and g18719 ( n28566 , n17 , n409 );
    and g18720 ( n42171 , n5512 , n6193 );
    and g18721 ( n37652 , n25613 , n30048 );
    xnor g18722 ( n29917 , n8837 , n40170 );
    or g18723 ( n33087 , n8511 , n41649 );
    or g18724 ( n27365 , n40588 , n24043 );
    not g18725 ( n10456 , n41969 );
    not g18726 ( n5183 , n28403 );
    or g18727 ( n9025 , n2924 , n34184 );
    not g18728 ( n1095 , n18419 );
    or g18729 ( n21398 , n38743 , n35382 );
    or g18730 ( n7124 , n9370 , n11205 );
    or g18731 ( n27697 , n9868 , n7474 );
    not g18732 ( n5170 , n25794 );
    or g18733 ( n36543 , n29382 , n15167 );
    nor g18734 ( n31515 , n31917 , n29000 );
    nor g18735 ( n17529 , n15070 , n41691 );
    or g18736 ( n8736 , n30068 , n42660 );
    and g18737 ( n24849 , n16540 , n20439 );
    nor g18738 ( n22210 , n33856 , n30247 );
    xnor g18739 ( n25292 , n11436 , n10694 );
    and g18740 ( n11424 , n11243 , n20217 );
    xnor g18741 ( n807 , n8837 , n36219 );
    or g18742 ( n24683 , n18371 , n14910 );
    or g18743 ( n28049 , n28048 , n14385 );
    or g18744 ( n34334 , n34139 , n30496 );
    nor g18745 ( n27577 , n1507 , n19015 );
    not g18746 ( n21096 , n15778 );
    or g18747 ( n27369 , n21752 , n488 );
    or g18748 ( n774 , n20525 , n40931 );
    xnor g18749 ( n25181 , n31989 , n14000 );
    and g18750 ( n29234 , n25844 , n29820 );
    or g18751 ( n16568 , n17176 , n20755 );
    not g18752 ( n18165 , n12805 );
    or g18753 ( n26711 , n40010 , n4629 );
    and g18754 ( n9554 , n34389 , n33707 );
    not g18755 ( n19070 , n37158 );
    or g18756 ( n32400 , n22440 , n26897 );
    not g18757 ( n8928 , n4746 );
    not g18758 ( n17090 , n7807 );
    or g18759 ( n22067 , n11410 , n1591 );
    xnor g18760 ( n9832 , n20783 , n32075 );
    nor g18761 ( n6733 , n3429 , n23156 );
    and g18762 ( n10872 , n16589 , n10814 );
    not g18763 ( n9733 , n25365 );
    or g18764 ( n511 , n8442 , n5343 );
    or g18765 ( n38515 , n13820 , n35010 );
    and g18766 ( n42507 , n39829 , n3141 );
    or g18767 ( n28378 , n23165 , n1679 );
    xnor g18768 ( n6514 , n41013 , n23 );
    or g18769 ( n35481 , n21752 , n6035 );
    or g18770 ( n29095 , n37137 , n22991 );
    and g18771 ( n5287 , n15796 , n9659 );
    not g18772 ( n40872 , n26775 );
    and g18773 ( n41787 , n37198 , n2490 );
    or g18774 ( n18346 , n35633 , n39865 );
    xnor g18775 ( n29792 , n22482 , n5602 );
    nor g18776 ( n31252 , n14993 , n12321 );
    nor g18777 ( n19953 , n25826 , n10073 );
    or g18778 ( n32419 , n42440 , n42428 );
    or g18779 ( n15466 , n34733 , n21852 );
    and g18780 ( n30204 , n21826 , n4814 );
    not g18781 ( n18883 , n41729 );
    or g18782 ( n29042 , n1979 , n21016 );
    nor g18783 ( n23653 , n31917 , n8613 );
    or g18784 ( n38458 , n34565 , n2838 );
    or g18785 ( n5641 , n39367 , n18081 );
    not g18786 ( n18689 , n42204 );
    not g18787 ( n3780 , n29805 );
    and g18788 ( n21028 , n3438 , n12160 );
    or g18789 ( n2314 , n31120 , n2710 );
    or g18790 ( n835 , n1735 , n3356 );
    and g18791 ( n28630 , n2085 , n11675 );
    nor g18792 ( n25634 , n6663 , n18710 );
    or g18793 ( n39926 , n27484 , n14170 );
    not g18794 ( n32180 , n33362 );
    xnor g18795 ( n21462 , n31048 , n4227 );
    and g18796 ( n37173 , n24999 , n6308 );
    and g18797 ( n29344 , n16992 , n592 );
    not g18798 ( n16079 , n4574 );
    nor g18799 ( n21702 , n21066 , n30200 );
    not g18800 ( n7251 , n38197 );
    or g18801 ( n22472 , n32898 , n12754 );
    or g18802 ( n33829 , n10930 , n29957 );
    and g18803 ( n42773 , n13123 , n15479 );
    and g18804 ( n15158 , n38495 , n42360 );
    and g18805 ( n20874 , n35768 , n30208 );
    nor g18806 ( n6046 , n15850 , n39880 );
    and g18807 ( n18181 , n35050 , n26781 );
    and g18808 ( n18269 , n16652 , n36150 );
    nor g18809 ( n41002 , n42003 , n19214 );
    xnor g18810 ( n18793 , n25620 , n25887 );
    nor g18811 ( n20888 , n7644 , n25015 );
    not g18812 ( n24717 , n6026 );
    or g18813 ( n8196 , n18956 , n14281 );
    or g18814 ( n20667 , n29406 , n23007 );
    or g18815 ( n5290 , n17383 , n11260 );
    or g18816 ( n35194 , n17120 , n19082 );
    and g18817 ( n10141 , n3532 , n19539 );
    not g18818 ( n15508 , n23631 );
    nor g18819 ( n7151 , n35615 , n11153 );
    xnor g18820 ( n28340 , n30264 , n29156 );
    xnor g18821 ( n11899 , n20793 , n20982 );
    and g18822 ( n4969 , n39998 , n26441 );
    not g18823 ( n12235 , n35103 );
    or g18824 ( n3737 , n36163 , n25749 );
    or g18825 ( n15582 , n26793 , n14281 );
    and g18826 ( n1217 , n28585 , n37157 );
    not g18827 ( n1355 , n14124 );
    or g18828 ( n10637 , n19469 , n6599 );
    or g18829 ( n10793 , n11824 , n29426 );
    nor g18830 ( n16876 , n36667 , n30008 );
    or g18831 ( n8295 , n16738 , n38963 );
    and g18832 ( n33304 , n36643 , n11669 );
    or g18833 ( n3103 , n2755 , n9031 );
    and g18834 ( n15607 , n913 , n37754 );
    and g18835 ( n14686 , n17718 , n19678 );
    and g18836 ( n18080 , n27369 , n28697 );
    and g18837 ( n10784 , n1698 , n40491 );
    not g18838 ( n31769 , n19925 );
    and g18839 ( n5819 , n12854 , n39592 );
    xnor g18840 ( n2218 , n29044 , n20676 );
    or g18841 ( n34674 , n29419 , n22797 );
    or g18842 ( n38526 , n29671 , n41047 );
    or g18843 ( n35644 , n5896 , n35140 );
    or g18844 ( n26643 , n18875 , n32527 );
    or g18845 ( n13127 , n18775 , n28535 );
    and g18846 ( n28431 , n41805 , n15721 );
    and g18847 ( n10620 , n37870 , n3950 );
    xnor g18848 ( n6894 , n35727 , n17398 );
    not g18849 ( n26995 , n40051 );
    or g18850 ( n31990 , n23717 , n9958 );
    or g18851 ( n30596 , n35087 , n37447 );
    or g18852 ( n7191 , n4130 , n24967 );
    nor g18853 ( n30640 , n22979 , n10041 );
    not g18854 ( n37309 , n12651 );
    and g18855 ( n3544 , n6408 , n17393 );
    not g18856 ( n1931 , n4708 );
    or g18857 ( n38620 , n25775 , n38897 );
    or g18858 ( n10291 , n30317 , n24078 );
    and g18859 ( n19885 , n27083 , n10825 );
    xnor g18860 ( n26630 , n33979 , n6444 );
    xnor g18861 ( n1458 , n42567 , n1265 );
    xnor g18862 ( n17336 , n29845 , n9363 );
    or g18863 ( n12899 , n41859 , n1380 );
    nor g18864 ( n18498 , n2214 , n5033 );
    or g18865 ( n276 , n6811 , n5717 );
    nor g18866 ( n13954 , n26058 , n37733 );
    not g18867 ( n41941 , n38752 );
    not g18868 ( n27051 , n30001 );
    xnor g18869 ( n1003 , n5144 , n22157 );
    or g18870 ( n11740 , n1460 , n10689 );
    xnor g18871 ( n42823 , n5464 , n15945 );
    or g18872 ( n12396 , n11172 , n16930 );
    or g18873 ( n14864 , n12738 , n34110 );
    and g18874 ( n30082 , n9864 , n33308 );
    xnor g18875 ( n32218 , n784 , n18486 );
    or g18876 ( n5949 , n22042 , n22584 );
    xnor g18877 ( n29185 , n11220 , n5025 );
    or g18878 ( n27876 , n16088 , n2352 );
    xnor g18879 ( n23465 , n24527 , n20118 );
    not g18880 ( n12021 , n40091 );
    and g18881 ( n12968 , n16639 , n19612 );
    or g18882 ( n22539 , n21894 , n22138 );
    or g18883 ( n12031 , n11745 , n17576 );
    and g18884 ( n2742 , n3864 , n40376 );
    xnor g18885 ( n39925 , n31099 , n28434 );
    not g18886 ( n35772 , n4961 );
    or g18887 ( n9849 , n26584 , n21284 );
    and g18888 ( n7293 , n35704 , n32559 );
    or g18889 ( n42688 , n6775 , n19142 );
    and g18890 ( n20242 , n23865 , n5453 );
    or g18891 ( n15295 , n22828 , n33859 );
    not g18892 ( n3581 , n17441 );
    or g18893 ( n24870 , n3764 , n32216 );
    not g18894 ( n28083 , n35455 );
    or g18895 ( n27356 , n38915 , n11825 );
    or g18896 ( n8690 , n32245 , n13148 );
    xnor g18897 ( n12434 , n26299 , n23684 );
    nor g18898 ( n37362 , n42792 , n15918 );
    and g18899 ( n12812 , n21621 , n37522 );
    or g18900 ( n36860 , n29980 , n24840 );
    xnor g18901 ( n9820 , n40549 , n2984 );
    or g18902 ( n41725 , n22973 , n9836 );
    xnor g18903 ( n41688 , n31099 , n25833 );
    or g18904 ( n39113 , n38708 , n13654 );
    or g18905 ( n17048 , n29782 , n26301 );
    not g18906 ( n3000 , n12942 );
    or g18907 ( n16235 , n42361 , n35558 );
    and g18908 ( n19106 , n30309 , n5425 );
    xnor g18909 ( n10641 , n42064 , n9749 );
    or g18910 ( n19978 , n18866 , n14686 );
    or g18911 ( n27860 , n25024 , n14181 );
    and g18912 ( n6013 , n14541 , n2895 );
    or g18913 ( n32801 , n41397 , n27127 );
    or g18914 ( n23305 , n10646 , n5434 );
    xnor g18915 ( n34109 , n25611 , n36538 );
    xnor g18916 ( n21568 , n35727 , n15922 );
    or g18917 ( n13109 , n775 , n20288 );
    and g18918 ( n40509 , n33208 , n42319 );
    or g18919 ( n9714 , n22990 , n36757 );
    xnor g18920 ( n23045 , n36998 , n39746 );
    not g18921 ( n15232 , n14233 );
    not g18922 ( n21133 , n40753 );
    or g18923 ( n19903 , n32277 , n32486 );
    nor g18924 ( n22314 , n8494 , n5466 );
    xnor g18925 ( n27977 , n10721 , n38003 );
    or g18926 ( n40572 , n10202 , n23753 );
    and g18927 ( n41783 , n7006 , n2271 );
    or g18928 ( n9897 , n36880 , n36518 );
    nor g18929 ( n15090 , n41741 , n25326 );
    or g18930 ( n27387 , n15709 , n1393 );
    and g18931 ( n28330 , n42764 , n31739 );
    or g18932 ( n16918 , n17954 , n15768 );
    or g18933 ( n14324 , n12059 , n27775 );
    and g18934 ( n12601 , n1445 , n11958 );
    or g18935 ( n4527 , n16330 , n35094 );
    or g18936 ( n15177 , n12866 , n40202 );
    and g18937 ( n12575 , n42358 , n41055 );
    not g18938 ( n11239 , n22073 );
    or g18939 ( n8642 , n27746 , n17172 );
    or g18940 ( n3131 , n28779 , n23272 );
    or g18941 ( n35645 , n17553 , n24665 );
    and g18942 ( n11660 , n963 , n470 );
    and g18943 ( n33702 , n18901 , n347 );
    or g18944 ( n29873 , n31367 , n31856 );
    or g18945 ( n39444 , n24344 , n24652 );
    or g18946 ( n29371 , n7572 , n26869 );
    or g18947 ( n21042 , n28634 , n40660 );
    or g18948 ( n26241 , n34565 , n18908 );
    or g18949 ( n31735 , n38009 , n844 );
    not g18950 ( n25845 , n32694 );
    nor g18951 ( n20263 , n36765 , n16430 );
    and g18952 ( n15529 , n38234 , n5907 );
    or g18953 ( n12126 , n36928 , n15095 );
    and g18954 ( n14051 , n21859 , n2295 );
    or g18955 ( n14580 , n11706 , n39129 );
    or g18956 ( n30667 , n36374 , n39728 );
    xnor g18957 ( n18008 , n23964 , n12096 );
    xnor g18958 ( n7023 , n35867 , n7031 );
    not g18959 ( n3916 , n17935 );
    or g18960 ( n8139 , n26739 , n6496 );
    xnor g18961 ( n35029 , n21735 , n5890 );
    xnor g18962 ( n10617 , n30166 , n35295 );
    or g18963 ( n15970 , n5790 , n946 );
    or g18964 ( n38007 , n18484 , n38175 );
    not g18965 ( n34167 , n15001 );
    and g18966 ( n41080 , n20475 , n5255 );
    and g18967 ( n7901 , n22615 , n12493 );
    and g18968 ( n5983 , n12126 , n22386 );
    or g18969 ( n33763 , n37796 , n42786 );
    and g18970 ( n11734 , n22308 , n36482 );
    and g18971 ( n17373 , n27810 , n27470 );
    nor g18972 ( n31495 , n27610 , n24116 );
    or g18973 ( n21148 , n22124 , n25102 );
    or g18974 ( n4178 , n14697 , n12457 );
    and g18975 ( n3436 , n39212 , n8890 );
    nor g18976 ( n9045 , n21184 , n29998 );
    nor g18977 ( n10836 , n3735 , n17849 );
    xnor g18978 ( n23381 , n5650 , n41877 );
    and g18979 ( n8459 , n11251 , n15390 );
    xnor g18980 ( n36918 , n13296 , n11808 );
    or g18981 ( n21808 , n2095 , n28445 );
    and g18982 ( n207 , n6378 , n34581 );
    and g18983 ( n24271 , n14970 , n26619 );
    xnor g18984 ( n14640 , n7282 , n23042 );
    or g18985 ( n19321 , n9357 , n36393 );
    not g18986 ( n7220 , n8676 );
    not g18987 ( n28593 , n19014 );
    or g18988 ( n3394 , n26915 , n30186 );
    nor g18989 ( n40216 , n1940 , n21583 );
    or g18990 ( n32197 , n2492 , n24905 );
    not g18991 ( n5959 , n37478 );
    not g18992 ( n24956 , n9174 );
    xnor g18993 ( n300 , n10226 , n25453 );
    or g18994 ( n27159 , n28129 , n2399 );
    and g18995 ( n34792 , n31383 , n38128 );
    or g18996 ( n30807 , n21372 , n31697 );
    nor g18997 ( n39671 , n16598 , n1139 );
    and g18998 ( n1460 , n7090 , n23631 );
    and g18999 ( n9159 , n13905 , n35912 );
    or g19000 ( n22272 , n5355 , n23164 );
    or g19001 ( n22678 , n10967 , n23974 );
    and g19002 ( n2330 , n16645 , n8562 );
    or g19003 ( n24541 , n39536 , n1063 );
    or g19004 ( n27829 , n18279 , n15282 );
    or g19005 ( n28048 , n32980 , n18871 );
    nor g19006 ( n13821 , n17960 , n16486 );
    or g19007 ( n19272 , n23472 , n22884 );
    and g19008 ( n32397 , n6908 , n4010 );
    xnor g19009 ( n20134 , n31099 , n8111 );
    xnor g19010 ( n22706 , n17558 , n18565 );
    xnor g19011 ( n35737 , n3062 , n33981 );
    nor g19012 ( n13634 , n14707 , n16115 );
    or g19013 ( n3102 , n41442 , n8401 );
    and g19014 ( n36787 , n13053 , n26306 );
    or g19015 ( n39600 , n18293 , n12320 );
    and g19016 ( n19964 , n3540 , n23465 );
    or g19017 ( n20828 , n24170 , n27292 );
    and g19018 ( n25238 , n2340 , n33610 );
    and g19019 ( n6874 , n4203 , n7784 );
    not g19020 ( n9030 , n33220 );
    not g19021 ( n15468 , n38145 );
    and g19022 ( n36335 , n13983 , n19467 );
    not g19023 ( n3311 , n1214 );
    or g19024 ( n15961 , n9187 , n25911 );
    or g19025 ( n8215 , n13746 , n30651 );
    or g19026 ( n19088 , n3120 , n23926 );
    and g19027 ( n40936 , n1666 , n22633 );
    or g19028 ( n20435 , n37832 , n27113 );
    or g19029 ( n8227 , n429 , n42446 );
    xnor g19030 ( n35293 , n14740 , n1502 );
    xnor g19031 ( n35671 , n119 , n14586 );
    xnor g19032 ( n4859 , n14932 , n35544 );
    or g19033 ( n30745 , n32565 , n30750 );
    not g19034 ( n25033 , n15396 );
    not g19035 ( n7903 , n30151 );
    or g19036 ( n40470 , n27701 , n4717 );
    and g19037 ( n9128 , n16905 , n6383 );
    nor g19038 ( n1453 , n27398 , n8798 );
    not g19039 ( n30623 , n16339 );
    not g19040 ( n12634 , n30851 );
    or g19041 ( n40963 , n17823 , n7569 );
    and g19042 ( n14504 , n5975 , n1655 );
    and g19043 ( n41191 , n36665 , n32240 );
    and g19044 ( n16318 , n8367 , n3126 );
    and g19045 ( n36652 , n12027 , n1014 );
    or g19046 ( n18329 , n26113 , n11780 );
    and g19047 ( n866 , n36311 , n37307 );
    or g19048 ( n35123 , n42335 , n7544 );
    xnor g19049 ( n42615 , n7193 , n29195 );
    nor g19050 ( n22422 , n37597 , n35623 );
    and g19051 ( n33685 , n9987 , n18158 );
    and g19052 ( n30112 , n27829 , n22225 );
    or g19053 ( n15228 , n40759 , n9373 );
    and g19054 ( n20899 , n14911 , n13439 );
    or g19055 ( n42878 , n17436 , n10788 );
    nor g19056 ( n32886 , n10427 , n35115 );
    and g19057 ( n37576 , n4926 , n19243 );
    xnor g19058 ( n12455 , n2674 , n32784 );
    xnor g19059 ( n16302 , n32297 , n8178 );
    nor g19060 ( n26238 , n10640 , n3948 );
    xnor g19061 ( n5788 , n784 , n41126 );
    or g19062 ( n38839 , n14368 , n23895 );
    and g19063 ( n23457 , n19934 , n22686 );
    or g19064 ( n38790 , n6483 , n41729 );
    not g19065 ( n7015 , n36378 );
    xnor g19066 ( n40958 , n31928 , n13815 );
    or g19067 ( n39135 , n34960 , n31339 );
    or g19068 ( n16420 , n39174 , n12045 );
    or g19069 ( n3950 , n18462 , n18638 );
    not g19070 ( n13795 , n7451 );
    or g19071 ( n10514 , n20141 , n28547 );
    xnor g19072 ( n36164 , n26475 , n9543 );
    and g19073 ( n8688 , n33584 , n38144 );
    or g19074 ( n21922 , n23008 , n2514 );
    or g19075 ( n11922 , n2532 , n13903 );
    not g19076 ( n28760 , n4442 );
    not g19077 ( n40322 , n8622 );
    not g19078 ( n31208 , n15946 );
    nor g19079 ( n19991 , n17170 , n32293 );
    or g19080 ( n17363 , n20545 , n27663 );
    or g19081 ( n21818 , n8560 , n4905 );
    or g19082 ( n3203 , n30527 , n25626 );
    or g19083 ( n39920 , n39804 , n21647 );
    nor g19084 ( n41635 , n13344 , n35236 );
    xnor g19085 ( n18732 , n17159 , n21777 );
    not g19086 ( n41413 , n12578 );
    or g19087 ( n33480 , n16586 , n30408 );
    xnor g19088 ( n41140 , n3455 , n9087 );
    or g19089 ( n23647 , n8585 , n37657 );
    or g19090 ( n11243 , n6546 , n21807 );
    or g19091 ( n6352 , n20231 , n16465 );
    xnor g19092 ( n25498 , n13932 , n21027 );
    nor g19093 ( n1091 , n30685 , n5764 );
    and g19094 ( n35896 , n14263 , n3428 );
    not g19095 ( n35722 , n12421 );
    or g19096 ( n25469 , n5750 , n18332 );
    xnor g19097 ( n37792 , n34562 , n3978 );
    or g19098 ( n34521 , n32151 , n3728 );
    or g19099 ( n3711 , n189 , n8658 );
    or g19100 ( n21619 , n20535 , n34723 );
    or g19101 ( n6780 , n24588 , n13862 );
    and g19102 ( n25121 , n9333 , n23874 );
    and g19103 ( n41415 , n31161 , n15865 );
    not g19104 ( n41437 , n21136 );
    or g19105 ( n32083 , n26675 , n36087 );
    or g19106 ( n3087 , n230 , n28686 );
    not g19107 ( n18524 , n22558 );
    and g19108 ( n22532 , n892 , n10126 );
    not g19109 ( n31742 , n30977 );
    nor g19110 ( n28928 , n5169 , n1844 );
    and g19111 ( n15869 , n26556 , n23864 );
    or g19112 ( n772 , n850 , n28341 );
    or g19113 ( n15785 , n17744 , n24119 );
    xnor g19114 ( n28498 , n23964 , n7749 );
    xnor g19115 ( n8558 , n20044 , n12312 );
    or g19116 ( n41804 , n4416 , n24602 );
    and g19117 ( n28030 , n8457 , n36629 );
    or g19118 ( n29647 , n23513 , n36324 );
    xnor g19119 ( n42917 , n34951 , n6859 );
    or g19120 ( n9693 , n26002 , n4839 );
    or g19121 ( n14311 , n19783 , n38687 );
    or g19122 ( n21945 , n26468 , n41201 );
    nor g19123 ( n34410 , n7063 , n11154 );
    or g19124 ( n40644 , n31166 , n21697 );
    and g19125 ( n15709 , n16 , n40618 );
    or g19126 ( n32418 , n15154 , n2672 );
    not g19127 ( n35441 , n13817 );
    or g19128 ( n33195 , n24581 , n2022 );
    and g19129 ( n29407 , n24720 , n10894 );
    nor g19130 ( n22411 , n6812 , n19499 );
    nor g19131 ( n29236 , n17744 , n23224 );
    or g19132 ( n17776 , n14325 , n8572 );
    and g19133 ( n10205 , n6405 , n35792 );
    nor g19134 ( n19993 , n10083 , n39467 );
    and g19135 ( n6750 , n37938 , n2994 );
    and g19136 ( n23455 , n30105 , n15797 );
    and g19137 ( n34221 , n25608 , n32463 );
    not g19138 ( n5349 , n331 );
    or g19139 ( n41660 , n34889 , n16891 );
    not g19140 ( n15934 , n13886 );
    or g19141 ( n38367 , n24164 , n3618 );
    or g19142 ( n13890 , n29097 , n25451 );
    nor g19143 ( n41355 , n10011 , n41712 );
    not g19144 ( n22126 , n39403 );
    or g19145 ( n29006 , n18184 , n16770 );
    and g19146 ( n36453 , n39451 , n35367 );
    xnor g19147 ( n27433 , n21598 , n5113 );
    or g19148 ( n33840 , n14689 , n33033 );
    or g19149 ( n30916 , n3636 , n9749 );
    or g19150 ( n2147 , n26060 , n24107 );
    or g19151 ( n8280 , n41215 , n25661 );
    or g19152 ( n39795 , n17984 , n40241 );
    and g19153 ( n40082 , n18245 , n7788 );
    xnor g19154 ( n30588 , n29667 , n26433 );
    and g19155 ( n22952 , n4984 , n26034 );
    or g19156 ( n35942 , n42076 , n9277 );
    not g19157 ( n29677 , n16077 );
    or g19158 ( n21327 , n23803 , n22991 );
    and g19159 ( n37678 , n10580 , n21105 );
    or g19160 ( n36814 , n4428 , n20430 );
    and g19161 ( n11558 , n23099 , n6676 );
    and g19162 ( n16730 , n31327 , n16634 );
    or g19163 ( n16040 , n17683 , n27226 );
    or g19164 ( n27872 , n29909 , n38191 );
    or g19165 ( n31453 , n29498 , n8983 );
    or g19166 ( n36350 , n20911 , n20025 );
    xnor g19167 ( n32591 , n31973 , n32580 );
    not g19168 ( n22247 , n29064 );
    or g19169 ( n16270 , n20633 , n26391 );
    or g19170 ( n11772 , n7646 , n37716 );
    and g19171 ( n17907 , n7694 , n29060 );
    xnor g19172 ( n35705 , n1664 , n15253 );
    xnor g19173 ( n32357 , n21571 , n7356 );
    or g19174 ( n36304 , n18970 , n15848 );
    and g19175 ( n32474 , n16064 , n31638 );
    or g19176 ( n3717 , n2637 , n41099 );
    or g19177 ( n30087 , n40443 , n9243 );
    and g19178 ( n27302 , n37 , n33550 );
    and g19179 ( n5039 , n15029 , n10923 );
    xnor g19180 ( n17179 , n20237 , n32885 );
    nor g19181 ( n37062 , n7585 , n3702 );
    and g19182 ( n26667 , n14678 , n30617 );
    nor g19183 ( n24818 , n38629 , n40195 );
    or g19184 ( n33150 , n12686 , n27863 );
    not g19185 ( n25919 , n9718 );
    and g19186 ( n6029 , n2067 , n15328 );
    and g19187 ( n39039 , n19101 , n37892 );
    nor g19188 ( n14309 , n33652 , n5831 );
    or g19189 ( n213 , n30263 , n25963 );
    not g19190 ( n31089 , n19248 );
    xnor g19191 ( n12087 , n41941 , n22115 );
    or g19192 ( n41242 , n34292 , n203 );
    or g19193 ( n40506 , n814 , n10698 );
    or g19194 ( n30029 , n10183 , n168 );
    xnor g19195 ( n20386 , n30397 , n35515 );
    xnor g19196 ( n14012 , n38957 , n15392 );
    xnor g19197 ( n26307 , n11109 , n40944 );
    nor g19198 ( n11892 , n31378 , n36186 );
    xnor g19199 ( n39756 , n19282 , n8642 );
    or g19200 ( n26128 , n31761 , n26595 );
    xnor g19201 ( n12843 , n17872 , n8652 );
    not g19202 ( n18242 , n16395 );
    not g19203 ( n7506 , n20080 );
    or g19204 ( n20595 , n16863 , n38582 );
    and g19205 ( n26228 , n17651 , n16616 );
    or g19206 ( n10830 , n41752 , n10254 );
    or g19207 ( n42275 , n32256 , n13170 );
    and g19208 ( n10604 , n26636 , n9175 );
    or g19209 ( n14463 , n14075 , n35418 );
    or g19210 ( n18259 , n17883 , n16962 );
    not g19211 ( n13687 , n27570 );
    and g19212 ( n29141 , n41960 , n19230 );
    or g19213 ( n14789 , n37404 , n2836 );
    or g19214 ( n38578 , n13033 , n16891 );
    not g19215 ( n24248 , n34487 );
    not g19216 ( n2497 , n9691 );
    or g19217 ( n23030 , n21349 , n29835 );
    and g19218 ( n10525 , n27638 , n23592 );
    xnor g19219 ( n9991 , n6345 , n622 );
    nor g19220 ( n13033 , n29827 , n38131 );
    or g19221 ( n41974 , n25353 , n25626 );
    nor g19222 ( n18601 , n14696 , n30895 );
    or g19223 ( n23434 , n25456 , n41612 );
    or g19224 ( n19264 , n2660 , n4316 );
    or g19225 ( n18017 , n1996 , n32378 );
    or g19226 ( n6460 , n1153 , n22350 );
    or g19227 ( n17771 , n35829 , n20776 );
    or g19228 ( n37673 , n12912 , n41437 );
    and g19229 ( n5861 , n30454 , n11680 );
    nor g19230 ( n3582 , n20728 , n26265 );
    or g19231 ( n12817 , n12661 , n20699 );
    nor g19232 ( n7513 , n16454 , n23832 );
    or g19233 ( n25524 , n30685 , n27819 );
    xnor g19234 ( n15081 , n35727 , n35192 );
    or g19235 ( n12066 , n29455 , n41386 );
    or g19236 ( n3484 , n10796 , n6000 );
    nor g19237 ( n5556 , n18866 , n33287 );
    or g19238 ( n26100 , n31142 , n15280 );
    or g19239 ( n22829 , n24719 , n26338 );
    or g19240 ( n168 , n41288 , n34087 );
    or g19241 ( n26642 , n13375 , n25303 );
    or g19242 ( n31683 , n21752 , n11949 );
    nor g19243 ( n17786 , n35428 , n6795 );
    or g19244 ( n25454 , n35014 , n38691 );
    and g19245 ( n34665 , n29096 , n9257 );
    and g19246 ( n26081 , n1102 , n24081 );
    or g19247 ( n17143 , n21036 , n23566 );
    and g19248 ( n36306 , n20434 , n31798 );
    not g19249 ( n23303 , n11144 );
    and g19250 ( n23300 , n10128 , n20656 );
    and g19251 ( n40556 , n13801 , n10327 );
    nor g19252 ( n28301 , n22243 , n38986 );
    nor g19253 ( n36359 , n30345 , n42754 );
    or g19254 ( n23443 , n42733 , n1970 );
    or g19255 ( n21529 , n2143 , n30358 );
    or g19256 ( n42136 , n39967 , n29930 );
    not g19257 ( n36348 , n37999 );
    nor g19258 ( n4213 , n10937 , n42106 );
    and g19259 ( n1320 , n38221 , n36183 );
    nor g19260 ( n4083 , n7825 , n36274 );
    nor g19261 ( n5327 , n28946 , n33111 );
    or g19262 ( n8840 , n24142 , n35633 );
    or g19263 ( n22433 , n2054 , n8998 );
    or g19264 ( n29566 , n9113 , n39282 );
    or g19265 ( n18680 , n19350 , n16513 );
    or g19266 ( n215 , n8625 , n22316 );
    or g19267 ( n30701 , n37282 , n7242 );
    not g19268 ( n19243 , n7418 );
    not g19269 ( n17161 , n25432 );
    and g19270 ( n2965 , n19025 , n40726 );
    nor g19271 ( n18701 , n27026 , n26956 );
    nor g19272 ( n13146 , n20804 , n39802 );
    and g19273 ( n4802 , n1843 , n37889 );
    xnor g19274 ( n32780 , n1467 , n31276 );
    or g19275 ( n38534 , n5721 , n14489 );
    or g19276 ( n42879 , n13077 , n35715 );
    nor g19277 ( n23809 , n17744 , n2713 );
    or g19278 ( n31682 , n38241 , n34504 );
    and g19279 ( n31113 , n11575 , n7883 );
    and g19280 ( n38257 , n5727 , n32736 );
    or g19281 ( n35311 , n27488 , n36479 );
    xnor g19282 ( n25523 , n23237 , n10461 );
    or g19283 ( n33498 , n18310 , n1270 );
    xnor g19284 ( n27491 , n35727 , n37894 );
    not g19285 ( n32860 , n39680 );
    not g19286 ( n2284 , n26036 );
    xnor g19287 ( n39386 , n15111 , n8844 );
    xnor g19288 ( n28058 , n18365 , n17246 );
    or g19289 ( n32756 , n35350 , n22578 );
    or g19290 ( n23191 , n22088 , n28499 );
    not g19291 ( n27721 , n20761 );
    not g19292 ( n26792 , n21115 );
    and g19293 ( n1857 , n39111 , n41168 );
    not g19294 ( n299 , n12168 );
    or g19295 ( n30252 , n28415 , n8329 );
    and g19296 ( n2335 , n27217 , n7866 );
    and g19297 ( n10680 , n33373 , n6352 );
    not g19298 ( n19700 , n36526 );
    xnor g19299 ( n10526 , n2339 , n12171 );
    or g19300 ( n33799 , n40824 , n26408 );
    or g19301 ( n40519 , n26961 , n31619 );
    nor g19302 ( n10780 , n325 , n26061 );
    and g19303 ( n22478 , n32720 , n24863 );
    and g19304 ( n16497 , n1604 , n25454 );
    and g19305 ( n17595 , n29441 , n35325 );
    and g19306 ( n30992 , n34856 , n27481 );
    or g19307 ( n20178 , n24348 , n17461 );
    and g19308 ( n33487 , n19567 , n14528 );
    and g19309 ( n31006 , n24908 , n6534 );
    and g19310 ( n33124 , n27703 , n19132 );
    or g19311 ( n19537 , n783 , n34398 );
    not g19312 ( n38541 , n18031 );
    nor g19313 ( n19679 , n24991 , n42411 );
    or g19314 ( n33888 , n9464 , n11141 );
    or g19315 ( n38385 , n22336 , n16150 );
    or g19316 ( n17707 , n21170 , n24276 );
    and g19317 ( n31164 , n105 , n4074 );
    nor g19318 ( n17536 , n13489 , n7082 );
    not g19319 ( n27792 , n2423 );
    or g19320 ( n12997 , n5644 , n19443 );
    and g19321 ( n11285 , n18470 , n27861 );
    and g19322 ( n40043 , n5994 , n37818 );
    xnor g19323 ( n40781 , n27396 , n31012 );
    or g19324 ( n31590 , n22010 , n1631 );
    and g19325 ( n31049 , n1753 , n5636 );
    not g19326 ( n32479 , n29568 );
    or g19327 ( n5400 , n21 , n42886 );
    or g19328 ( n25744 , n3591 , n1083 );
    not g19329 ( n655 , n7074 );
    not g19330 ( n19928 , n499 );
    or g19331 ( n29807 , n24588 , n34393 );
    or g19332 ( n18747 , n16780 , n34686 );
    and g19333 ( n35999 , n18076 , n20770 );
    or g19334 ( n496 , n41998 , n10632 );
    not g19335 ( n656 , n15554 );
    not g19336 ( n21023 , n8734 );
    not g19337 ( n9272 , n26613 );
    and g19338 ( n22571 , n16693 , n15338 );
    not g19339 ( n30263 , n36298 );
    or g19340 ( n22357 , n23031 , n21239 );
    or g19341 ( n8331 , n15095 , n40042 );
    not g19342 ( n34290 , n42805 );
    xnor g19343 ( n1143 , n10414 , n7065 );
    and g19344 ( n12492 , n29042 , n93 );
    and g19345 ( n23468 , n13836 , n9603 );
    or g19346 ( n8727 , n28725 , n23423 );
    or g19347 ( n16151 , n34594 , n29380 );
    and g19348 ( n43 , n3961 , n38503 );
    or g19349 ( n2620 , n41090 , n24316 );
    xnor g19350 ( n42061 , n1813 , n32164 );
    nor g19351 ( n18938 , n39757 , n2538 );
    not g19352 ( n36872 , n3663 );
    and g19353 ( n8014 , n40149 , n3422 );
    or g19354 ( n14171 , n14490 , n17317 );
    or g19355 ( n2787 , n33655 , n6798 );
    nor g19356 ( n3661 , n10434 , n25966 );
    xnor g19357 ( n14629 , n34235 , n16472 );
    or g19358 ( n27397 , n34090 , n5707 );
    or g19359 ( n2859 , n19083 , n31671 );
    or g19360 ( n5925 , n35347 , n17934 );
    xnor g19361 ( n16889 , n1917 , n13285 );
    nor g19362 ( n23763 , n8971 , n4594 );
    and g19363 ( n30317 , n14133 , n8839 );
    or g19364 ( n31312 , n14471 , n18456 );
    or g19365 ( n17584 , n12434 , n35167 );
    not g19366 ( n8847 , n40720 );
    or g19367 ( n26501 , n30163 , n3881 );
    and g19368 ( n23517 , n13127 , n24646 );
    and g19369 ( n19133 , n30157 , n20585 );
    or g19370 ( n31035 , n28021 , n3298 );
    and g19371 ( n34906 , n35760 , n397 );
    and g19372 ( n40371 , n33396 , n37833 );
    not g19373 ( n23421 , n24730 );
    not g19374 ( n22197 , n13527 );
    or g19375 ( n27379 , n38142 , n19232 );
    xnor g19376 ( n20820 , n15972 , n10998 );
    and g19377 ( n24223 , n25261 , n14554 );
    xnor g19378 ( n42604 , n15426 , n34917 );
    and g19379 ( n36726 , n15145 , n39369 );
    xnor g19380 ( n15488 , n40176 , n20532 );
    or g19381 ( n8119 , n12645 , n29061 );
    not g19382 ( n37437 , n1903 );
    or g19383 ( n31628 , n16831 , n2675 );
    nor g19384 ( n11054 , n15860 , n15013 );
    or g19385 ( n21955 , n31838 , n41215 );
    or g19386 ( n28103 , n10137 , n38423 );
    or g19387 ( n26656 , n29058 , n22618 );
    or g19388 ( n15835 , n9408 , n18310 );
    or g19389 ( n20279 , n35732 , n16319 );
    not g19390 ( n6796 , n2431 );
    or g19391 ( n33306 , n23509 , n26361 );
    or g19392 ( n40435 , n2743 , n33196 );
    nor g19393 ( n9248 , n30166 , n11362 );
    or g19394 ( n20438 , n42870 , n22131 );
    or g19395 ( n31651 , n25483 , n26942 );
    or g19396 ( n13355 , n39662 , n36168 );
    and g19397 ( n14192 , n40280 , n19949 );
    or g19398 ( n20979 , n34036 , n21023 );
    or g19399 ( n9082 , n33794 , n21650 );
    nor g19400 ( n9354 , n18866 , n24007 );
    or g19401 ( n35063 , n27881 , n11592 );
    or g19402 ( n5837 , n6980 , n12120 );
    and g19403 ( n30511 , n14933 , n22583 );
    or g19404 ( n20080 , n21969 , n3236 );
    and g19405 ( n1484 , n12310 , n36632 );
    or g19406 ( n33722 , n26269 , n13960 );
    not g19407 ( n3939 , n6755 );
    and g19408 ( n28430 , n21434 , n12623 );
    nor g19409 ( n16602 , n5896 , n39661 );
    and g19410 ( n24563 , n38949 , n8488 );
    and g19411 ( n35288 , n34757 , n20344 );
    or g19412 ( n2249 , n29497 , n39149 );
    or g19413 ( n9366 , n4535 , n19251 );
    or g19414 ( n23633 , n23140 , n13368 );
    or g19415 ( n38106 , n3436 , n31643 );
    or g19416 ( n33507 , n6584 , n42839 );
    nor g19417 ( n37363 , n2468 , n35517 );
    or g19418 ( n4503 , n9222 , n34148 );
    xnor g19419 ( n752 , n31053 , n18013 );
    or g19420 ( n17710 , n22437 , n1168 );
    or g19421 ( n26145 , n13528 , n41981 );
    xnor g19422 ( n27349 , n33944 , n30215 );
    and g19423 ( n23400 , n25292 , n20918 );
    or g19424 ( n26514 , n21596 , n4099 );
    nor g19425 ( n8636 , n19004 , n32698 );
    or g19426 ( n7423 , n16443 , n21856 );
    or g19427 ( n39284 , n16738 , n31759 );
    and g19428 ( n38756 , n28018 , n24117 );
    or g19429 ( n34084 , n37266 , n1006 );
    not g19430 ( n22484 , n27086 );
    and g19431 ( n7335 , n10507 , n29972 );
    xnor g19432 ( n23001 , n25849 , n4747 );
    or g19433 ( n16774 , n8574 , n13438 );
    xnor g19434 ( n35291 , n23067 , n19580 );
    and g19435 ( n16148 , n30317 , n24078 );
    not g19436 ( n6565 , n32009 );
    xnor g19437 ( n6553 , n32138 , n35212 );
    or g19438 ( n34416 , n17817 , n40566 );
    or g19439 ( n27805 , n32242 , n3661 );
    nor g19440 ( n39463 , n5896 , n41732 );
    nor g19441 ( n35040 , n26446 , n20350 );
    xnor g19442 ( n33716 , n1316 , n35467 );
    or g19443 ( n4041 , n29314 , n29492 );
    or g19444 ( n33338 , n3571 , n7194 );
    not g19445 ( n21351 , n13178 );
    or g19446 ( n41445 , n35499 , n13885 );
    or g19447 ( n40228 , n1176 , n29002 );
    and g19448 ( n14959 , n38648 , n12868 );
    or g19449 ( n10259 , n9508 , n28128 );
    or g19450 ( n3869 , n4335 , n24255 );
    and g19451 ( n14738 , n22792 , n41700 );
    nor g19452 ( n33191 , n27439 , n23337 );
    or g19453 ( n11715 , n8173 , n8149 );
    or g19454 ( n29586 , n31674 , n21977 );
    or g19455 ( n11197 , n37707 , n38756 );
    or g19456 ( n11939 , n8453 , n30658 );
    or g19457 ( n18011 , n10530 , n17840 );
    xnor g19458 ( n37082 , n11633 , n35960 );
    not g19459 ( n26545 , n41956 );
    not g19460 ( n34205 , n29937 );
    or g19461 ( n31260 , n36466 , n25581 );
    or g19462 ( n29245 , n40457 , n4929 );
    nor g19463 ( n27719 , n15261 , n20660 );
    or g19464 ( n8243 , n31954 , n22201 );
    and g19465 ( n17389 , n18038 , n12940 );
    or g19466 ( n39476 , n5083 , n29652 );
    or g19467 ( n12142 , n19996 , n12220 );
    or g19468 ( n25344 , n29932 , n30514 );
    nor g19469 ( n911 , n12599 , n29929 );
    nor g19470 ( n7446 , n33368 , n9167 );
    nor g19471 ( n11471 , n8857 , n19765 );
    and g19472 ( n18316 , n4761 , n1629 );
    or g19473 ( n15994 , n4266 , n39056 );
    or g19474 ( n32322 , n4282 , n18528 );
    and g19475 ( n10177 , n9528 , n35810 );
    or g19476 ( n7829 , n32954 , n41215 );
    not g19477 ( n7701 , n3911 );
    and g19478 ( n3503 , n5694 , n36207 );
    or g19479 ( n23384 , n7954 , n4139 );
    or g19480 ( n40311 , n32775 , n17249 );
    and g19481 ( n6270 , n39077 , n31080 );
    or g19482 ( n28413 , n23480 , n28883 );
    and g19483 ( n8136 , n4035 , n27443 );
    or g19484 ( n36596 , n38068 , n14879 );
    not g19485 ( n38829 , n38263 );
    or g19486 ( n32031 , n22266 , n37250 );
    or g19487 ( n1682 , n15282 , n16192 );
    or g19488 ( n16442 , n33752 , n23640 );
    xnor g19489 ( n31969 , n9412 , n9725 );
    not g19490 ( n29038 , n26069 );
    xnor g19491 ( n35041 , n28185 , n7979 );
    nor g19492 ( n2265 , n42591 , n19878 );
    and g19493 ( n25909 , n40120 , n4603 );
    not g19494 ( n426 , n7946 );
    or g19495 ( n7743 , n38175 , n30172 );
    not g19496 ( n22831 , n14653 );
    or g19497 ( n1131 , n7165 , n36095 );
    or g19498 ( n38537 , n42708 , n2675 );
    or g19499 ( n34022 , n38528 , n10320 );
    not g19500 ( n11596 , n31764 );
    or g19501 ( n31320 , n16611 , n35830 );
    or g19502 ( n40545 , n22333 , n23435 );
    nor g19503 ( n6438 , n14707 , n40948 );
    or g19504 ( n3076 , n24621 , n27392 );
    nor g19505 ( n40011 , n33891 , n34427 );
    nor g19506 ( n39968 , n6188 , n35497 );
    or g19507 ( n132 , n25969 , n37787 );
    or g19508 ( n17351 , n23307 , n32259 );
    or g19509 ( n9262 , n27020 , n33129 );
    xnor g19510 ( n31647 , n42686 , n14752 );
    and g19511 ( n9923 , n8622 , n16420 );
    or g19512 ( n19593 , n23591 , n18814 );
    or g19513 ( n14904 , n16530 , n40574 );
    or g19514 ( n41316 , n41356 , n2065 );
    and g19515 ( n27851 , n31413 , n27659 );
    not g19516 ( n22740 , n22754 );
    xnor g19517 ( n11646 , n5013 , n1185 );
    and g19518 ( n27340 , n18952 , n32429 );
    nor g19519 ( n20099 , n11072 , n631 );
    xnor g19520 ( n33298 , n40774 , n2098 );
    and g19521 ( n30687 , n1810 , n29072 );
    or g19522 ( n35433 , n6203 , n20450 );
    or g19523 ( n4890 , n6572 , n1795 );
    or g19524 ( n31205 , n27769 , n11832 );
    and g19525 ( n13329 , n12327 , n22285 );
    and g19526 ( n10247 , n41805 , n6658 );
    and g19527 ( n29231 , n31206 , n7247 );
    or g19528 ( n22591 , n4843 , n36771 );
    and g19529 ( n38160 , n30901 , n15226 );
    or g19530 ( n16112 , n5203 , n26177 );
    or g19531 ( n2595 , n33289 , n6524 );
    or g19532 ( n41083 , n33677 , n11779 );
    and g19533 ( n40736 , n36679 , n22190 );
    or g19534 ( n35159 , n31707 , n22818 );
    and g19535 ( n520 , n7658 , n29529 );
    not g19536 ( n36809 , n37839 );
    or g19537 ( n38612 , n42447 , n1809 );
    and g19538 ( n27034 , n37747 , n35765 );
    and g19539 ( n10073 , n21416 , n11803 );
    or g19540 ( n14156 , n35287 , n30138 );
    xnor g19541 ( n21885 , n28600 , n35205 );
    nor g19542 ( n9584 , n32589 , n41314 );
    or g19543 ( n475 , n19218 , n23241 );
    and g19544 ( n21239 , n3741 , n32702 );
    not g19545 ( n15108 , n14054 );
    or g19546 ( n27069 , n240 , n22424 );
    not g19547 ( n26256 , n19406 );
    or g19548 ( n12216 , n12560 , n25303 );
    or g19549 ( n31899 , n40212 , n13039 );
    not g19550 ( n13760 , n31064 );
    nor g19551 ( n7113 , n2086 , n40895 );
    or g19552 ( n24710 , n16598 , n23897 );
    or g19553 ( n11544 , n28344 , n23577 );
    or g19554 ( n7908 , n29027 , n4563 );
    not g19555 ( n27644 , n31352 );
    or g19556 ( n36830 , n14723 , n13003 );
    not g19557 ( n36330 , n39809 );
    not g19558 ( n29057 , n1572 );
    and g19559 ( n27827 , n24242 , n25513 );
    and g19560 ( n18566 , n33801 , n17208 );
    or g19561 ( n36440 , n3487 , n1098 );
    or g19562 ( n12277 , n26640 , n31515 );
    or g19563 ( n14541 , n27317 , n13771 );
    or g19564 ( n21749 , n26927 , n7077 );
    or g19565 ( n1253 , n10182 , n21856 );
    and g19566 ( n24503 , n21340 , n38033 );
    or g19567 ( n16139 , n13058 , n36019 );
    and g19568 ( n116 , n5269 , n8342 );
    and g19569 ( n2416 , n26418 , n18537 );
    or g19570 ( n24556 , n2069 , n11520 );
    or g19571 ( n22226 , n23796 , n15943 );
    or g19572 ( n22099 , n40306 , n33321 );
    or g19573 ( n9979 , n1175 , n42544 );
    and g19574 ( n33154 , n31802 , n3065 );
    and g19575 ( n5153 , n3666 , n307 );
    or g19576 ( n36152 , n19562 , n31624 );
    or g19577 ( n42805 , n18950 , n10904 );
    or g19578 ( n10481 , n22910 , n24852 );
    and g19579 ( n27455 , n5270 , n6140 );
    not g19580 ( n17712 , n3026 );
    nor g19581 ( n7075 , n36667 , n24893 );
    not g19582 ( n6160 , n33526 );
    or g19583 ( n26160 , n31110 , n6635 );
    or g19584 ( n8474 , n6987 , n2565 );
    or g19585 ( n34668 , n14289 , n21579 );
    and g19586 ( n30690 , n39054 , n34914 );
    or g19587 ( n15073 , n9446 , n5294 );
    or g19588 ( n34543 , n1507 , n33902 );
    or g19589 ( n21541 , n2815 , n21471 );
    nor g19590 ( n8592 , n22827 , n11859 );
    not g19591 ( n19498 , n32709 );
    or g19592 ( n28888 , n28144 , n20273 );
    or g19593 ( n39879 , n7933 , n11410 );
    nor g19594 ( n35564 , n11445 , n9049 );
    nor g19595 ( n42464 , n26347 , n8497 );
    xnor g19596 ( n9306 , n5404 , n37649 );
    not g19597 ( n41811 , n29163 );
    and g19598 ( n32185 , n18128 , n8472 );
    or g19599 ( n32555 , n26281 , n2647 );
    or g19600 ( n10362 , n31741 , n36056 );
    or g19601 ( n786 , n41176 , n26639 );
    nor g19602 ( n42596 , n6894 , n32142 );
    xnor g19603 ( n18913 , n13444 , n21906 );
    xnor g19604 ( n25562 , n20502 , n29753 );
    or g19605 ( n38520 , n15571 , n15272 );
    and g19606 ( n16733 , n17854 , n28380 );
    nor g19607 ( n19533 , n18995 , n9520 );
    and g19608 ( n42504 , n7464 , n22931 );
    and g19609 ( n28937 , n1873 , n3407 );
    and g19610 ( n19375 , n13055 , n3260 );
    not g19611 ( n23968 , n22060 );
    or g19612 ( n40224 , n30860 , n42025 );
    or g19613 ( n40379 , n40329 , n22282 );
    or g19614 ( n40063 , n6148 , n2400 );
    nor g19615 ( n38193 , n4140 , n34284 );
    and g19616 ( n30064 , n25819 , n1512 );
    or g19617 ( n32071 , n29436 , n14351 );
    or g19618 ( n8027 , n15003 , n13603 );
    or g19619 ( n1807 , n29451 , n15276 );
    not g19620 ( n34358 , n28595 );
    and g19621 ( n36540 , n16334 , n35946 );
    or g19622 ( n42608 , n17121 , n25223 );
    xnor g19623 ( n1772 , n10577 , n20903 );
    or g19624 ( n27807 , n14379 , n21046 );
    or g19625 ( n23134 , n14644 , n15184 );
    xnor g19626 ( n8604 , n30271 , n20201 );
    not g19627 ( n17586 , n995 );
    nor g19628 ( n10484 , n6774 , n11487 );
    and g19629 ( n2399 , n3074 , n1302 );
    or g19630 ( n37941 , n20098 , n36052 );
    or g19631 ( n31449 , n28647 , n27303 );
    or g19632 ( n31755 , n30866 , n8898 );
    or g19633 ( n13015 , n38157 , n16455 );
    xnor g19634 ( n13128 , n27751 , n12965 );
    or g19635 ( n2219 , n2726 , n23489 );
    and g19636 ( n2297 , n9686 , n41172 );
    not g19637 ( n5581 , n21704 );
    or g19638 ( n10453 , n1499 , n29969 );
    or g19639 ( n8443 , n35732 , n5313 );
    xnor g19640 ( n6850 , n8951 , n41534 );
    not g19641 ( n40176 , n35307 );
    or g19642 ( n14002 , n28667 , n10355 );
    xnor g19643 ( n16168 , n36423 , n1191 );
    not g19644 ( n8502 , n26919 );
    or g19645 ( n39587 , n13392 , n10699 );
    or g19646 ( n39494 , n31452 , n11199 );
    or g19647 ( n3005 , n28774 , n37506 );
    and g19648 ( n7956 , n21891 , n13135 );
    or g19649 ( n14693 , n33582 , n6024 );
    or g19650 ( n41459 , n12856 , n20197 );
    and g19651 ( n25158 , n6782 , n11447 );
    and g19652 ( n28505 , n7571 , n10322 );
    xnor g19653 ( n3626 , n13046 , n28561 );
    and g19654 ( n27952 , n32651 , n17333 );
    xnor g19655 ( n24679 , n31564 , n36382 );
    not g19656 ( n22319 , n24984 );
    or g19657 ( n28853 , n28551 , n27367 );
    or g19658 ( n37480 , n20541 , n19545 );
    and g19659 ( n9430 , n38043 , n18290 );
    not g19660 ( n2183 , n1568 );
    nor g19661 ( n10194 , n32291 , n41084 );
    and g19662 ( n37724 , n1537 , n26564 );
    and g19663 ( n40004 , n11022 , n18483 );
    and g19664 ( n6014 , n15151 , n37189 );
    nor g19665 ( n13948 , n6049 , n6934 );
    or g19666 ( n11634 , n30153 , n34673 );
    xnor g19667 ( n39129 , n15285 , n36446 );
    or g19668 ( n16210 , n25840 , n5570 );
    not g19669 ( n10256 , n36372 );
    and g19670 ( n18543 , n37905 , n7260 );
    or g19671 ( n23064 , n3636 , n39775 );
    or g19672 ( n42818 , n8126 , n903 );
    and g19673 ( n18964 , n23825 , n3565 );
    or g19674 ( n9458 , n29980 , n8324 );
    nor g19675 ( n5620 , n25414 , n8163 );
    not g19676 ( n6525 , n24027 );
    and g19677 ( n17318 , n18098 , n21170 );
    or g19678 ( n15910 , n27625 , n8123 );
    nor g19679 ( n31298 , n12874 , n13881 );
    not g19680 ( n23760 , n19582 );
    not g19681 ( n25249 , n11557 );
    xnor g19682 ( n23287 , n29740 , n1948 );
    and g19683 ( n36158 , n3685 , n5730 );
    xnor g19684 ( n7688 , n22054 , n41252 );
    or g19685 ( n19200 , n8442 , n42620 );
    and g19686 ( n33447 , n18467 , n25550 );
    or g19687 ( n35285 , n24605 , n18495 );
    nor g19688 ( n39252 , n34483 , n22896 );
    or g19689 ( n35315 , n39438 , n41404 );
    or g19690 ( n40356 , n41489 , n34246 );
    or g19691 ( n7258 , n3764 , n16917 );
    or g19692 ( n827 , n40178 , n9709 );
    and g19693 ( n27329 , n29882 , n37823 );
    and g19694 ( n27261 , n39751 , n5470 );
    nor g19695 ( n17024 , n17906 , n26433 );
    or g19696 ( n19551 , n33655 , n26079 );
    nor g19697 ( n15981 , n5896 , n35809 );
    or g19698 ( n31478 , n9114 , n2311 );
    and g19699 ( n2682 , n11675 , n23106 );
    or g19700 ( n37781 , n11339 , n34267 );
    and g19701 ( n34158 , n11836 , n20462 );
    or g19702 ( n26259 , n8790 , n19828 );
    xnor g19703 ( n36968 , n21534 , n18822 );
    or g19704 ( n24073 , n15610 , n7265 );
    or g19705 ( n14951 , n38149 , n36197 );
    xnor g19706 ( n26077 , n4503 , n25058 );
    or g19707 ( n26308 , n3571 , n41169 );
    not g19708 ( n13474 , n21178 );
    and g19709 ( n4700 , n13403 , n32330 );
    nor g19710 ( n42046 , n23535 , n38281 );
    xnor g19711 ( n25895 , n29323 , n4892 );
    xnor g19712 ( n899 , n15617 , n724 );
    xnor g19713 ( n20845 , n13444 , n35679 );
    not g19714 ( n23941 , n33639 );
    or g19715 ( n37593 , n9880 , n38530 );
    or g19716 ( n34420 , n19663 , n25389 );
    nor g19717 ( n35566 , n17120 , n33705 );
    nor g19718 ( n41549 , n10245 , n37020 );
    and g19719 ( n40948 , n3819 , n26480 );
    or g19720 ( n6015 , n5299 , n6332 );
    xnor g19721 ( n24390 , n37899 , n19349 );
    and g19722 ( n12847 , n2894 , n1557 );
    or g19723 ( n18794 , n22242 , n22209 );
    and g19724 ( n40482 , n12124 , n15714 );
    xnor g19725 ( n7431 , n32632 , n19064 );
    or g19726 ( n40610 , n11021 , n38423 );
    and g19727 ( n29012 , n19239 , n20627 );
    or g19728 ( n2500 , n6125 , n17649 );
    or g19729 ( n41666 , n16343 , n37733 );
    nor g19730 ( n37144 , n33436 , n328 );
    xnor g19731 ( n28257 , n34352 , n19375 );
    or g19732 ( n29064 , n36681 , n18872 );
    or g19733 ( n36609 , n30863 , n6788 );
    or g19734 ( n5511 , n6606 , n14837 );
    or g19735 ( n13911 , n17393 , n8558 );
    or g19736 ( n34553 , n39042 , n8979 );
    not g19737 ( n3138 , n4794 );
    nor g19738 ( n15600 , n28601 , n5976 );
    xnor g19739 ( n33050 , n11534 , n33963 );
    or g19740 ( n1238 , n41943 , n31803 );
    or g19741 ( n13069 , n2756 , n14806 );
    not g19742 ( n11814 , n36942 );
    or g19743 ( n33015 , n31750 , n32489 );
    nor g19744 ( n11548 , n17965 , n18259 );
    nor g19745 ( n32126 , n30855 , n8982 );
    nor g19746 ( n32863 , n19221 , n18822 );
    xnor g19747 ( n10297 , n34875 , n35401 );
    nor g19748 ( n12674 , n24442 , n27105 );
    or g19749 ( n23143 , n12112 , n36379 );
    and g19750 ( n20950 , n15937 , n16814 );
    or g19751 ( n4172 , n41152 , n33321 );
    and g19752 ( n29915 , n27328 , n559 );
    or g19753 ( n38859 , n35184 , n25281 );
    nor g19754 ( n6559 , n14530 , n13752 );
    not g19755 ( n18800 , n40153 );
    nor g19756 ( n33957 , n10519 , n15141 );
    xnor g19757 ( n221 , n1863 , n27945 );
    not g19758 ( n34858 , n3084 );
    not g19759 ( n3373 , n7644 );
    and g19760 ( n37683 , n32417 , n9231 );
    not g19761 ( n2763 , n26613 );
    not g19762 ( n16505 , n27555 );
    nor g19763 ( n18576 , n4673 , n22793 );
    or g19764 ( n24373 , n9544 , n23390 );
    not g19765 ( n18544 , n6982 );
    xnor g19766 ( n23137 , n31017 , n7736 );
    not g19767 ( n38617 , n26791 );
    nor g19768 ( n29380 , n36730 , n33921 );
    not g19769 ( n25007 , n27740 );
    xnor g19770 ( n18356 , n41013 , n14766 );
    or g19771 ( n19146 , n25793 , n16576 );
    not g19772 ( n5564 , n31128 );
    or g19773 ( n5137 , n28116 , n17404 );
    not g19774 ( n7425 , n30083 );
    not g19775 ( n20995 , n24896 );
    and g19776 ( n38690 , n38745 , n34876 );
    not g19777 ( n3776 , n28597 );
    or g19778 ( n16233 , n12867 , n29065 );
    xnor g19779 ( n36645 , n6841 , n36401 );
    nor g19780 ( n22603 , n27598 , n33479 );
    or g19781 ( n28844 , n23296 , n22584 );
    not g19782 ( n24210 , n32485 );
    or g19783 ( n32968 , n38157 , n37791 );
    or g19784 ( n25008 , n23739 , n6013 );
    or g19785 ( n7861 , n18003 , n37633 );
    not g19786 ( n11835 , n26729 );
    nor g19787 ( n18552 , n21592 , n31482 );
    or g19788 ( n13588 , n12937 , n500 );
    or g19789 ( n10323 , n1997 , n36407 );
    nor g19790 ( n42745 , n20728 , n23774 );
    and g19791 ( n8432 , n31884 , n22829 );
    not g19792 ( n12418 , n41841 );
    not g19793 ( n6281 , n30372 );
    not g19794 ( n30083 , n9691 );
    and g19795 ( n4883 , n10777 , n5664 );
    nor g19796 ( n8398 , n1507 , n2556 );
    xnor g19797 ( n11852 , n12146 , n33304 );
    or g19798 ( n22298 , n21175 , n26093 );
    and g19799 ( n7916 , n27970 , n19897 );
    and g19800 ( n28987 , n24711 , n18415 );
    or g19801 ( n33096 , n19580 , n14687 );
    or g19802 ( n24205 , n25865 , n4305 );
    nor g19803 ( n24714 , n30634 , n12253 );
    not g19804 ( n5814 , n14221 );
    not g19805 ( n7690 , n22377 );
    nor g19806 ( n8070 , n33211 , n19401 );
    not g19807 ( n1702 , n28843 );
    or g19808 ( n7464 , n3801 , n17356 );
    or g19809 ( n35390 , n39260 , n10637 );
    or g19810 ( n24516 , n12017 , n39699 );
    or g19811 ( n906 , n29524 , n19840 );
    and g19812 ( n13347 , n25248 , n2938 );
    not g19813 ( n24301 , n2428 );
    or g19814 ( n6193 , n5884 , n6253 );
    and g19815 ( n39946 , n21484 , n7191 );
    not g19816 ( n21162 , n42290 );
    or g19817 ( n30198 , n14287 , n26193 );
    not g19818 ( n9372 , n23229 );
    not g19819 ( n4972 , n8182 );
    and g19820 ( n10350 , n24773 , n16014 );
    xnor g19821 ( n26075 , n42244 , n446 );
    or g19822 ( n27855 , n14490 , n29403 );
    and g19823 ( n14455 , n34307 , n13484 );
    or g19824 ( n27044 , n28745 , n19342 );
    or g19825 ( n29103 , n15542 , n28061 );
    and g19826 ( n10804 , n28 , n42483 );
    and g19827 ( n7758 , n33284 , n20208 );
    xnor g19828 ( n26840 , n8036 , n26517 );
    or g19829 ( n10671 , n21603 , n38115 );
    and g19830 ( n14811 , n22317 , n31013 );
    or g19831 ( n34443 , n10954 , n32951 );
    and g19832 ( n28375 , n15395 , n3724 );
    not g19833 ( n27308 , n30438 );
    or g19834 ( n39087 , n26089 , n5623 );
    and g19835 ( n24024 , n1438 , n20947 );
    and g19836 ( n33288 , n29235 , n10564 );
    or g19837 ( n16417 , n36203 , n11035 );
    and g19838 ( n10053 , n6175 , n39116 );
    not g19839 ( n12424 , n16069 );
    nor g19840 ( n14182 , n37367 , n18133 );
    or g19841 ( n374 , n37881 , n36590 );
    or g19842 ( n23832 , n36430 , n42830 );
    xnor g19843 ( n16894 , n27371 , n34557 );
    and g19844 ( n34308 , n27681 , n12537 );
    or g19845 ( n18999 , n34793 , n39615 );
    or g19846 ( n10920 , n15738 , n11778 );
    nor g19847 ( n4431 , n15285 , n8505 );
    or g19848 ( n24407 , n39930 , n13330 );
    nor g19849 ( n41514 , n2199 , n39155 );
    nor g19850 ( n28158 , n5964 , n22640 );
    or g19851 ( n1362 , n4639 , n29299 );
    not g19852 ( n9419 , n9571 );
    and g19853 ( n16455 , n33339 , n13682 );
    not g19854 ( n3303 , n42356 );
    not g19855 ( n8487 , n31955 );
    not g19856 ( n24729 , n35411 );
    or g19857 ( n31941 , n41162 , n25486 );
    xnor g19858 ( n13728 , n11168 , n36929 );
    and g19859 ( n27823 , n4453 , n30659 );
    or g19860 ( n42283 , n38648 , n12868 );
    or g19861 ( n2453 , n36496 , n35109 );
    not g19862 ( n1533 , n36048 );
    and g19863 ( n24378 , n27630 , n19136 );
    and g19864 ( n6197 , n35536 , n4251 );
    nor g19865 ( n37493 , n17964 , n1821 );
    or g19866 ( n27057 , n28667 , n19145 );
    and g19867 ( n13810 , n36763 , n34181 );
    or g19868 ( n5021 , n28215 , n41590 );
    not g19869 ( n37922 , n27148 );
    or g19870 ( n9131 , n38704 , n38943 );
    or g19871 ( n24453 , n11231 , n24240 );
    nor g19872 ( n29485 , n5356 , n10132 );
    and g19873 ( n41359 , n19428 , n27791 );
    not g19874 ( n9376 , n28595 );
    nor g19875 ( n36294 , n35700 , n27 );
    xnor g19876 ( n24772 , n29438 , n7126 );
    or g19877 ( n39377 , n27311 , n456 );
    or g19878 ( n4493 , n32212 , n14259 );
    and g19879 ( n34863 , n40049 , n25635 );
    xnor g19880 ( n18527 , n21534 , n24305 );
    or g19881 ( n3152 , n697 , n13653 );
    or g19882 ( n114 , n20338 , n12096 );
    nor g19883 ( n9195 , n7639 , n30043 );
    nor g19884 ( n14095 , n37707 , n30547 );
    or g19885 ( n4480 , n3113 , n7385 );
    not g19886 ( n36189 , n8045 );
    or g19887 ( n30476 , n42177 , n37120 );
    or g19888 ( n18099 , n17256 , n17559 );
    and g19889 ( n35933 , n19302 , n12833 );
    or g19890 ( n10322 , n5280 , n24881 );
    or g19891 ( n33650 , n38890 , n9487 );
    or g19892 ( n33862 , n22907 , n902 );
    xnor g19893 ( n36216 , n30521 , n16598 );
    or g19894 ( n9295 , n18324 , n26765 );
    and g19895 ( n1956 , n42695 , n7138 );
    nor g19896 ( n37974 , n19262 , n15090 );
    or g19897 ( n2764 , n14048 , n8507 );
    not g19898 ( n11489 , n2848 );
    or g19899 ( n8982 , n42778 , n14617 );
    not g19900 ( n34162 , n21983 );
    and g19901 ( n29817 , n5936 , n30787 );
    or g19902 ( n39961 , n8494 , n2600 );
    and g19903 ( n23717 , n33791 , n5697 );
    not g19904 ( n7548 , n26242 );
    nor g19905 ( n14128 , n1011 , n31166 );
    or g19906 ( n21492 , n33316 , n18236 );
    and g19907 ( n35187 , n6186 , n32854 );
    nor g19908 ( n29637 , n20039 , n27355 );
    xnor g19909 ( n5872 , n26996 , n36851 );
    or g19910 ( n31181 , n43 , n22646 );
    xnor g19911 ( n29132 , n34735 , n15077 );
    not g19912 ( n35840 , n21809 );
    or g19913 ( n39691 , n37954 , n20030 );
    and g19914 ( n3133 , n28477 , n34263 );
    or g19915 ( n22781 , n18648 , n14087 );
    or g19916 ( n16180 , n17062 , n39439 );
    and g19917 ( n19922 , n6581 , n32098 );
    or g19918 ( n8189 , n1417 , n6263 );
    or g19919 ( n27442 , n17393 , n31137 );
    or g19920 ( n393 , n36824 , n29932 );
    and g19921 ( n16192 , n23113 , n19506 );
    or g19922 ( n9427 , n1791 , n17576 );
    or g19923 ( n22796 , n11857 , n29058 );
    and g19924 ( n41584 , n23407 , n41149 );
    nor g19925 ( n19882 , n5957 , n20465 );
    nor g19926 ( n33233 , n39571 , n23540 );
    xnor g19927 ( n38744 , n14005 , n25212 );
    not g19928 ( n24498 , n12332 );
    and g19929 ( n3738 , n37069 , n33250 );
    or g19930 ( n2641 , n23420 , n36880 );
    nor g19931 ( n8352 , n13785 , n40660 );
    and g19932 ( n18795 , n25588 , n42746 );
    not g19933 ( n27045 , n4864 );
    or g19934 ( n5885 , n37056 , n7321 );
    or g19935 ( n6312 , n16826 , n19237 );
    or g19936 ( n15213 , n34466 , n24712 );
    xnor g19937 ( n34472 , n31677 , n4156 );
    or g19938 ( n40046 , n7813 , n2479 );
    and g19939 ( n16970 , n37257 , n28257 );
    or g19940 ( n1808 , n13880 , n33216 );
    not g19941 ( n19017 , n24354 );
    or g19942 ( n38212 , n13433 , n12528 );
    not g19943 ( n15384 , n25642 );
    and g19944 ( n7395 , n31815 , n11953 );
    xnor g19945 ( n15769 , n14515 , n20659 );
    not g19946 ( n38350 , n36137 );
    not g19947 ( n25793 , n11689 );
    or g19948 ( n35225 , n17596 , n10611 );
    nor g19949 ( n26735 , n37237 , n5482 );
    or g19950 ( n18304 , n31699 , n22441 );
    and g19951 ( n26843 , n1937 , n33919 );
    and g19952 ( n17000 , n37599 , n9085 );
    nor g19953 ( n6629 , n17583 , n12650 );
    or g19954 ( n12074 , n32705 , n34510 );
    and g19955 ( n20650 , n12368 , n16278 );
    xnor g19956 ( n3616 , n30721 , n12591 );
    and g19957 ( n37477 , n26718 , n13817 );
    nor g19958 ( n18432 , n27722 , n9722 );
    and g19959 ( n5899 , n31103 , n16794 );
    or g19960 ( n13763 , n9591 , n31875 );
    or g19961 ( n7484 , n11230 , n13529 );
    nor g19962 ( n3263 , n19001 , n24126 );
    not g19963 ( n28830 , n29843 );
    not g19964 ( n29980 , n21881 );
    or g19965 ( n6166 , n21373 , n36179 );
    or g19966 ( n17054 , n21560 , n37733 );
    and g19967 ( n21553 , n19418 , n16282 );
    or g19968 ( n1796 , n14645 , n22091 );
    or g19969 ( n15002 , n1075 , n11424 );
    or g19970 ( n27511 , n41446 , n781 );
    nor g19971 ( n16394 , n34565 , n21091 );
    or g19972 ( n27979 , n18471 , n35834 );
    nor g19973 ( n34073 , n13717 , n20082 );
    xnor g19974 ( n13505 , n35113 , n36910 );
    not g19975 ( n26716 , n28428 );
    or g19976 ( n35343 , n12808 , n6900 );
    or g19977 ( n5038 , n34730 , n22892 );
    or g19978 ( n26614 , n2662 , n34517 );
    xnor g19979 ( n32896 , n14594 , n5091 );
    not g19980 ( n4538 , n1419 );
    or g19981 ( n4133 , n21893 , n41107 );
    and g19982 ( n7354 , n40596 , n17885 );
    and g19983 ( n6254 , n3576 , n38593 );
    not g19984 ( n35267 , n23239 );
    and g19985 ( n7961 , n1016 , n32501 );
    xnor g19986 ( n24445 , n35711 , n32332 );
    and g19987 ( n30241 , n24304 , n5668 );
    or g19988 ( n39375 , n244 , n12887 );
    not g19989 ( n13215 , n4782 );
    not g19990 ( n39699 , n22863 );
    or g19991 ( n33573 , n24025 , n24535 );
    xnor g19992 ( n12586 , n20876 , n35334 );
    or g19993 ( n27736 , n10598 , n29970 );
    or g19994 ( n24435 , n37388 , n11705 );
    and g19995 ( n23821 , n10973 , n38811 );
    or g19996 ( n16689 , n13573 , n41007 );
    not g19997 ( n36014 , n29684 );
    and g19998 ( n16757 , n6203 , n20450 );
    or g19999 ( n37719 , n2868 , n466 );
    and g20000 ( n26051 , n22467 , n30989 );
    xnor g20001 ( n25237 , n25299 , n23015 );
    or g20002 ( n18203 , n122 , n34098 );
    xnor g20003 ( n22506 , n18990 , n38061 );
    or g20004 ( n17644 , n12198 , n42304 );
    nor g20005 ( n10673 , n4693 , n16828 );
    xnor g20006 ( n7895 , n3455 , n12352 );
    and g20007 ( n12432 , n10813 , n32838 );
    nor g20008 ( n17840 , n4322 , n22400 );
    or g20009 ( n21723 , n12920 , n40455 );
    or g20010 ( n4613 , n39951 , n38578 );
    and g20011 ( n8476 , n40190 , n1435 );
    and g20012 ( n31101 , n11138 , n20868 );
    and g20013 ( n31315 , n16503 , n34524 );
    or g20014 ( n6531 , n27761 , n13010 );
    or g20015 ( n233 , n1688 , n10691 );
    or g20016 ( n24819 , n16780 , n4871 );
    not g20017 ( n23057 , n26823 );
    not g20018 ( n38762 , n42391 );
    xnor g20019 ( n1776 , n24913 , n10228 );
    or g20020 ( n33645 , n15709 , n39595 );
    or g20021 ( n6409 , n19641 , n4706 );
    or g20022 ( n14132 , n5964 , n27211 );
    not g20023 ( n24617 , n40697 );
    xnor g20024 ( n41704 , n40176 , n39379 );
    or g20025 ( n34591 , n25619 , n12553 );
    or g20026 ( n4577 , n9437 , n16712 );
    or g20027 ( n36308 , n11558 , n32341 );
    nor g20028 ( n21879 , n19522 , n2977 );
    xnor g20029 ( n26018 , n31607 , n39460 );
    and g20030 ( n28816 , n23814 , n28189 );
    not g20031 ( n33926 , n29731 );
    nor g20032 ( n13080 , n17872 , n16344 );
    or g20033 ( n37971 , n27311 , n14547 );
    or g20034 ( n23813 , n27120 , n1999 );
    and g20035 ( n936 , n37918 , n33603 );
    or g20036 ( n35130 , n14884 , n29904 );
    not g20037 ( n5077 , n24886 );
    xnor g20038 ( n28089 , n21534 , n29531 );
    or g20039 ( n25844 , n32077 , n27632 );
    nor g20040 ( n2245 , n16817 , n38860 );
    or g20041 ( n25068 , n13332 , n19672 );
    or g20042 ( n22196 , n17984 , n13645 );
    xnor g20043 ( n34112 , n32132 , n40999 );
    and g20044 ( n4752 , n23037 , n21853 );
    nor g20045 ( n13413 , n27758 , n3247 );
    or g20046 ( n20718 , n26681 , n37462 );
    or g20047 ( n35778 , n7148 , n15780 );
    nor g20048 ( n37992 , n16885 , n19375 );
    xnor g20049 ( n41900 , n18990 , n36431 );
    or g20050 ( n14133 , n5896 , n20366 );
    nor g20051 ( n34571 , n17436 , n18984 );
    or g20052 ( n13309 , n35466 , n36751 );
    nor g20053 ( n38224 , n17193 , n7752 );
    nor g20054 ( n19488 , n41390 , n10896 );
    or g20055 ( n28446 , n33842 , n32318 );
    xnor g20056 ( n476 , n25884 , n13552 );
    or g20057 ( n8303 , n17193 , n9920 );
    xnor g20058 ( n40985 , n24265 , n18779 );
    and g20059 ( n29169 , n4433 , n24257 );
    and g20060 ( n18081 , n25931 , n30751 );
    xnor g20061 ( n7324 , n2464 , n18866 );
    not g20062 ( n28294 , n10409 );
    nor g20063 ( n7821 , n28152 , n2569 );
    or g20064 ( n24469 , n26025 , n41532 );
    nor g20065 ( n17010 , n17958 , n10091 );
    xnor g20066 ( n4906 , n12146 , n41639 );
    and g20067 ( n32311 , n30427 , n33249 );
    or g20068 ( n34301 , n36071 , n21059 );
    xnor g20069 ( n7764 , n42472 , n39979 );
    not g20070 ( n10132 , n40560 );
    or g20071 ( n32490 , n7142 , n21885 );
    or g20072 ( n2638 , n27311 , n16955 );
    xnor g20073 ( n29879 , n16952 , n6881 );
    and g20074 ( n22266 , n33006 , n20123 );
    or g20075 ( n32448 , n27619 , n17841 );
    or g20076 ( n236 , n21690 , n25933 );
    or g20077 ( n8233 , n1357 , n21268 );
    or g20078 ( n26004 , n20684 , n14402 );
    or g20079 ( n35300 , n4307 , n31758 );
    not g20080 ( n20610 , n5026 );
    nor g20081 ( n3441 , n2199 , n34423 );
    or g20082 ( n19428 , n7296 , n28159 );
    nor g20083 ( n42074 , n40067 , n41288 );
    and g20084 ( n15639 , n24871 , n10795 );
    not g20085 ( n31728 , n32596 );
    or g20086 ( n36436 , n22504 , n42351 );
    xnor g20087 ( n32955 , n16693 , n29343 );
    nor g20088 ( n4540 , n7585 , n13154 );
    or g20089 ( n24272 , n30519 , n115 );
    xnor g20090 ( n29203 , n13444 , n5129 );
    or g20091 ( n16225 , n26909 , n256 );
    xnor g20092 ( n7538 , n36009 , n34132 );
    xnor g20093 ( n9389 , n40391 , n3627 );
    not g20094 ( n25696 , n29442 );
    nor g20095 ( n18450 , n26345 , n30493 );
    or g20096 ( n16796 , n387 , n37911 );
    or g20097 ( n2157 , n15721 , n19603 );
    not g20098 ( n12877 , n34576 );
    or g20099 ( n37033 , n37494 , n3901 );
    and g20100 ( n40100 , n1680 , n38018 );
    or g20101 ( n20732 , n29192 , n41682 );
    or g20102 ( n25165 , n23634 , n15182 );
    xnor g20103 ( n16382 , n10641 , n41173 );
    or g20104 ( n40263 , n1554 , n14901 );
    or g20105 ( n24799 , n11283 , n31388 );
    not g20106 ( n13232 , n21753 );
    or g20107 ( n38287 , n32605 , n35603 );
    or g20108 ( n38656 , n37752 , n13687 );
    and g20109 ( n24965 , n39736 , n27498 );
    and g20110 ( n21164 , n7055 , n22678 );
    or g20111 ( n21999 , n10047 , n17083 );
    or g20112 ( n10932 , n40446 , n6291 );
    or g20113 ( n38491 , n23563 , n27275 );
    not g20114 ( n25910 , n26641 );
    or g20115 ( n33470 , n16412 , n32995 );
    not g20116 ( n4782 , n37653 );
    or g20117 ( n42035 , n22120 , n19240 );
    and g20118 ( n18718 , n3652 , n21685 );
    nor g20119 ( n1575 , n33876 , n9381 );
    and g20120 ( n8164 , n4821 , n15290 );
    or g20121 ( n23951 , n24459 , n21856 );
    nor g20122 ( n31731 , n39266 , n27507 );
    or g20123 ( n4025 , n23772 , n37756 );
    and g20124 ( n36560 , n7126 , n29438 );
    xnor g20125 ( n29760 , n542 , n19081 );
    and g20126 ( n10997 , n13849 , n12750 );
    not g20127 ( n30429 , n7221 );
    not g20128 ( n7907 , n31448 );
    or g20129 ( n34659 , n10979 , n7206 );
    or g20130 ( n9781 , n145 , n2565 );
    or g20131 ( n31715 , n13553 , n8243 );
    and g20132 ( n40961 , n3211 , n27846 );
    nor g20133 ( n29918 , n34483 , n18101 );
    or g20134 ( n42012 , n1455 , n35064 );
    or g20135 ( n34649 , n30201 , n40419 );
    or g20136 ( n35881 , n14345 , n29382 );
    and g20137 ( n16483 , n12502 , n40373 );
    not g20138 ( n2458 , n14170 );
    or g20139 ( n2712 , n37671 , n4338 );
    xnor g20140 ( n8026 , n5058 , n7298 );
    or g20141 ( n18094 , n26502 , n4843 );
    and g20142 ( n11603 , n26850 , n517 );
    not g20143 ( n37582 , n25308 );
    not g20144 ( n28021 , n14589 );
    nor g20145 ( n6713 , n6957 , n35843 );
    xnor g20146 ( n24127 , n23504 , n22680 );
    or g20147 ( n5171 , n29675 , n27052 );
    or g20148 ( n20840 , n30822 , n2039 );
    and g20149 ( n3274 , n9683 , n36356 );
    and g20150 ( n17883 , n12311 , n23539 );
    or g20151 ( n14176 , n33985 , n37804 );
    xnor g20152 ( n37932 , n784 , n10880 );
    not g20153 ( n30969 , n34279 );
    not g20154 ( n20572 , n21562 );
    or g20155 ( n15930 , n34138 , n35772 );
    nor g20156 ( n25341 , n14707 , n1820 );
    or g20157 ( n15453 , n37425 , n1326 );
    not g20158 ( n29651 , n10837 );
    not g20159 ( n2145 , n29606 );
    not g20160 ( n16751 , n9978 );
    or g20161 ( n31231 , n34778 , n17830 );
    or g20162 ( n39232 , n16587 , n38499 );
    nor g20163 ( n32168 , n27026 , n34552 );
    or g20164 ( n28192 , n23671 , n37921 );
    or g20165 ( n30628 , n8763 , n34270 );
    or g20166 ( n2670 , n16161 , n17390 );
    and g20167 ( n24037 , n35582 , n12373 );
    or g20168 ( n35658 , n21391 , n30214 );
    or g20169 ( n14401 , n724 , n32180 );
    and g20170 ( n3192 , n6129 , n31178 );
    and g20171 ( n7244 , n31882 , n728 );
    xnor g20172 ( n42916 , n12769 , n7710 );
    not g20173 ( n22821 , n13300 );
    or g20174 ( n36261 , n3580 , n18219 );
    or g20175 ( n41078 , n5189 , n33828 );
    or g20176 ( n37822 , n331 , n34624 );
    or g20177 ( n33855 , n28359 , n19084 );
    and g20178 ( n18003 , n12716 , n1639 );
    nor g20179 ( n39345 , n17906 , n41102 );
    xnor g20180 ( n27123 , n1429 , n34397 );
    or g20181 ( n36582 , n5324 , n8151 );
    not g20182 ( n23868 , n21710 );
    or g20183 ( n28172 , n37637 , n4155 );
    or g20184 ( n19253 , n20180 , n8401 );
    and g20185 ( n23435 , n29095 , n29151 );
    or g20186 ( n23890 , n34429 , n7815 );
    not g20187 ( n35879 , n39392 );
    and g20188 ( n39306 , n19912 , n39307 );
    nor g20189 ( n8039 , n25554 , n30707 );
    xnor g20190 ( n29265 , n28185 , n7275 );
    or g20191 ( n31623 , n10440 , n1725 );
    or g20192 ( n21461 , n13997 , n2602 );
    not g20193 ( n33838 , n16582 );
    not g20194 ( n9350 , n4829 );
    nor g20195 ( n2353 , n20847 , n12855 );
    not g20196 ( n19433 , n27671 );
    or g20197 ( n23061 , n32972 , n12028 );
    not g20198 ( n42115 , n8569 );
    not g20199 ( n25060 , n32009 );
    nor g20200 ( n40597 , n37223 , n29717 );
    or g20201 ( n5371 , n41620 , n19753 );
    not g20202 ( n17627 , n20648 );
    not g20203 ( n8787 , n24023 );
    or g20204 ( n22276 , n29655 , n27738 );
    or g20205 ( n13471 , n22294 , n33496 );
    or g20206 ( n27565 , n7356 , n5658 );
    xnor g20207 ( n7477 , n22263 , n8541 );
    and g20208 ( n12550 , n21431 , n36220 );
    nor g20209 ( n17240 , n25409 , n17549 );
    or g20210 ( n15274 , n6510 , n3918 );
    or g20211 ( n25699 , n3590 , n12153 );
    nor g20212 ( n5845 , n11542 , n33608 );
    xnor g20213 ( n27613 , n25619 , n20734 );
    and g20214 ( n15963 , n21967 , n8013 );
    or g20215 ( n33282 , n26934 , n15780 );
    or g20216 ( n1600 , n32715 , n6316 );
    and g20217 ( n4452 , n38929 , n8749 );
    nor g20218 ( n41890 , n39456 , n12084 );
    or g20219 ( n29032 , n18042 , n3801 );
    or g20220 ( n33399 , n34223 , n13425 );
    or g20221 ( n19920 , n5959 , n34179 );
    or g20222 ( n28358 , n19830 , n14884 );
    nor g20223 ( n38720 , n33981 , n4751 );
    and g20224 ( n14099 , n42196 , n36554 );
    and g20225 ( n27711 , n34018 , n40084 );
    or g20226 ( n27219 , n13565 , n7772 );
    or g20227 ( n8360 , n12194 , n31361 );
    or g20228 ( n3710 , n5087 , n18162 );
    and g20229 ( n10385 , n34934 , n6873 );
    and g20230 ( n23965 , n5336 , n19831 );
    and g20231 ( n23714 , n10109 , n3193 );
    and g20232 ( n40335 , n15023 , n41797 );
    and g20233 ( n8169 , n23264 , n30589 );
    or g20234 ( n13715 , n25579 , n7172 );
    xnor g20235 ( n14637 , n33570 , n34284 );
    or g20236 ( n15686 , n28164 , n13215 );
    and g20237 ( n7992 , n3512 , n37416 );
    or g20238 ( n14839 , n38021 , n12495 );
    or g20239 ( n31951 , n27699 , n15780 );
    not g20240 ( n3068 , n3759 );
    nor g20241 ( n11113 , n25081 , n39518 );
    nor g20242 ( n27482 , n41834 , n34348 );
    xnor g20243 ( n11694 , n36365 , n36902 );
    and g20244 ( n37317 , n20745 , n21681 );
    or g20245 ( n42231 , n41526 , n33336 );
    xnor g20246 ( n4614 , n21654 , n13549 );
    and g20247 ( n14000 , n23642 , n27867 );
    xnor g20248 ( n15008 , n25426 , n42221 );
    and g20249 ( n17247 , n19451 , n17233 );
    or g20250 ( n5470 , n19779 , n27082 );
    or g20251 ( n24555 , n16736 , n29259 );
    xnor g20252 ( n13563 , n5648 , n7530 );
    nor g20253 ( n30683 , n20571 , n40022 );
    or g20254 ( n6983 , n18465 , n3775 );
    or g20255 ( n21718 , n5119 , n38339 );
    not g20256 ( n18700 , n28621 );
    or g20257 ( n24087 , n2127 , n25963 );
    xnor g20258 ( n42444 , n13444 , n9632 );
    xnor g20259 ( n2665 , n29034 , n16359 );
    not g20260 ( n14188 , n38197 );
    or g20261 ( n20038 , n17397 , n12347 );
    or g20262 ( n33793 , n26989 , n36457 );
    or g20263 ( n11290 , n29980 , n7547 );
    not g20264 ( n12007 , n26650 );
    nor g20265 ( n1288 , n25643 , n12209 );
    nor g20266 ( n22290 , n898 , n5303 );
    nor g20267 ( n34168 , n23745 , n16148 );
    or g20268 ( n3386 , n26237 , n36844 );
    not g20269 ( n23767 , n39322 );
    not g20270 ( n15608 , n1096 );
    or g20271 ( n8343 , n40703 , n17126 );
    or g20272 ( n36826 , n6012 , n14776 );
    or g20273 ( n10246 , n1110 , n7473 );
    xnor g20274 ( n9397 , n12339 , n28272 );
    or g20275 ( n32945 , n12431 , n18566 );
    or g20276 ( n21360 , n6024 , n7144 );
    not g20277 ( n3906 , n18718 );
    nor g20278 ( n39312 , n1178 , n8155 );
    or g20279 ( n30630 , n28667 , n39430 );
    not g20280 ( n41695 , n6054 );
    and g20281 ( n11367 , n26233 , n26106 );
    nor g20282 ( n34642 , n26949 , n9833 );
    and g20283 ( n609 , n17147 , n20023 );
    and g20284 ( n9917 , n39873 , n27155 );
    and g20285 ( n7851 , n4217 , n33041 );
    not g20286 ( n34920 , n36793 );
    xnor g20287 ( n24954 , n20487 , n25522 );
    and g20288 ( n30183 , n1229 , n30016 );
    and g20289 ( n1370 , n33944 , n30215 );
    nor g20290 ( n36685 , n35371 , n27440 );
    xnor g20291 ( n15598 , n784 , n18522 );
    and g20292 ( n39621 , n2579 , n33659 );
    not g20293 ( n1287 , n18807 );
    not g20294 ( n5348 , n20072 );
    nor g20295 ( n23056 , n2971 , n3256 );
    and g20296 ( n18763 , n40621 , n32631 );
    and g20297 ( n32167 , n13518 , n26983 );
    and g20298 ( n4880 , n25827 , n11796 );
    xnor g20299 ( n13139 , n105 , n34169 );
    nor g20300 ( n3350 , n4225 , n5469 );
    or g20301 ( n38804 , n37119 , n39936 );
    or g20302 ( n15203 , n29037 , n5718 );
    and g20303 ( n33738 , n30945 , n16675 );
    and g20304 ( n37365 , n33023 , n16906 );
    or g20305 ( n7153 , n18235 , n6772 );
    not g20306 ( n1080 , n10739 );
    and g20307 ( n36130 , n829 , n42434 );
    or g20308 ( n5554 , n26681 , n11996 );
    xnor g20309 ( n6355 , n37210 , n41089 );
    nor g20310 ( n39478 , n33745 , n1640 );
    or g20311 ( n37726 , n36080 , n21023 );
    or g20312 ( n28744 , n37643 , n20231 );
    and g20313 ( n11106 , n27971 , n27906 );
    not g20314 ( n39149 , n35781 );
    not g20315 ( n37070 , n2878 );
    or g20316 ( n9542 , n7079 , n41487 );
    and g20317 ( n36573 , n2887 , n42524 );
    nor g20318 ( n21000 , n41677 , n41814 );
    xnor g20319 ( n21495 , n30752 , n24704 );
    nor g20320 ( n22716 , n708 , n34074 );
    not g20321 ( n2430 , n13008 );
    or g20322 ( n13788 , n16363 , n37659 );
    xnor g20323 ( n16434 , n1290 , n10598 );
    xnor g20324 ( n5167 , n17674 , n4978 );
    xnor g20325 ( n34690 , n7628 , n26876 );
    nor g20326 ( n30172 , n26307 , n18615 );
    and g20327 ( n7708 , n42267 , n40047 );
    and g20328 ( n1740 , n29868 , n35778 );
    or g20329 ( n4487 , n23550 , n22669 );
    and g20330 ( n25818 , n8271 , n42281 );
    and g20331 ( n24049 , n29591 , n29512 );
    not g20332 ( n2018 , n14008 );
    xnor g20333 ( n9760 , n26362 , n36708 );
    or g20334 ( n11098 , n19538 , n30621 );
    xnor g20335 ( n17150 , n36998 , n34534 );
    nor g20336 ( n10915 , n32042 , n24618 );
    or g20337 ( n26511 , n14314 , n18673 );
    or g20338 ( n31508 , n15934 , n162 );
    and g20339 ( n21387 , n353 , n39087 );
    or g20340 ( n37820 , n5896 , n17788 );
    not g20341 ( n6625 , n14707 );
    or g20342 ( n35625 , n41958 , n42544 );
    or g20343 ( n14111 , n42774 , n15181 );
    or g20344 ( n763 , n39930 , n32080 );
    or g20345 ( n25261 , n35632 , n6293 );
    nor g20346 ( n14754 , n30110 , n38078 );
    or g20347 ( n408 , n3162 , n33456 );
    not g20348 ( n19416 , n39065 );
    and g20349 ( n30487 , n27061 , n32403 );
    xnor g20350 ( n35112 , n14740 , n23396 );
    xnor g20351 ( n31995 , n1110 , n24699 );
    or g20352 ( n12065 , n35231 , n2410 );
    xnor g20353 ( n10013 , n24476 , n24971 );
    not g20354 ( n28092 , n13507 );
    not g20355 ( n25456 , n4382 );
    or g20356 ( n11517 , n4660 , n11661 );
    not g20357 ( n4632 , n2570 );
    and g20358 ( n14366 , n39338 , n25601 );
    and g20359 ( n38354 , n27723 , n22087 );
    or g20360 ( n1302 , n4262 , n21109 );
    not g20361 ( n16303 , n25091 );
    and g20362 ( n21375 , n12567 , n41268 );
    not g20363 ( n28362 , n28150 );
    or g20364 ( n40776 , n404 , n38050 );
    not g20365 ( n15163 , n9013 );
    and g20366 ( n38465 , n34022 , n238 );
    xnor g20367 ( n21008 , n12146 , n22021 );
    or g20368 ( n24046 , n22340 , n28283 );
    xnor g20369 ( n39656 , n9234 , n37680 );
    not g20370 ( n39314 , n34048 );
    and g20371 ( n15460 , n1582 , n8835 );
    or g20372 ( n20374 , n23079 , n35713 );
    nor g20373 ( n26096 , n31884 , n22829 );
    or g20374 ( n35400 , n7181 , n27648 );
    not g20375 ( n16996 , n27188 );
    or g20376 ( n10097 , n40588 , n21660 );
    nor g20377 ( n19625 , n37146 , n20035 );
    not g20378 ( n41046 , n30824 );
    and g20379 ( n31214 , n19468 , n40065 );
    or g20380 ( n17863 , n14060 , n12909 );
    and g20381 ( n17800 , n2931 , n6862 );
    not g20382 ( n9113 , n37357 );
    or g20383 ( n4058 , n303 , n39302 );
    or g20384 ( n11058 , n4717 , n4758 );
    not g20385 ( n12038 , n22775 );
    or g20386 ( n3374 , n32095 , n28107 );
    or g20387 ( n18688 , n27263 , n36955 );
    or g20388 ( n39175 , n22693 , n13566 );
    not g20389 ( n33581 , n7305 );
    or g20390 ( n10091 , n20622 , n40444 );
    not g20391 ( n6883 , n28255 );
    not g20392 ( n29851 , n757 );
    or g20393 ( n3998 , n39652 , n27037 );
    not g20394 ( n2919 , n26749 );
    and g20395 ( n7376 , n25539 , n33242 );
    or g20396 ( n20997 , n1265 , n31924 );
    not g20397 ( n1965 , n34030 );
    or g20398 ( n5276 , n20250 , n2547 );
    or g20399 ( n21645 , n35016 , n9745 );
    nor g20400 ( n26987 , n39639 , n21507 );
    or g20401 ( n14639 , n3824 , n18635 );
    or g20402 ( n11007 , n11775 , n42694 );
    and g20403 ( n24212 , n21568 , n22261 );
    xnor g20404 ( n8906 , n33884 , n3120 );
    and g20405 ( n29434 , n35152 , n15838 );
    xnor g20406 ( n16608 , n40928 , n38071 );
    and g20407 ( n33977 , n213 , n34335 );
    or g20408 ( n19447 , n18155 , n27618 );
    or g20409 ( n27301 , n4076 , n34626 );
    or g20410 ( n1770 , n17176 , n36125 );
    xnor g20411 ( n20933 , n18530 , n22701 );
    and g20412 ( n888 , n32299 , n11195 );
    or g20413 ( n23436 , n11340 , n37913 );
    or g20414 ( n24455 , n8313 , n1340 );
    or g20415 ( n4924 , n33464 , n36782 );
    and g20416 ( n18114 , n23652 , n40417 );
    xnor g20417 ( n9215 , n784 , n15287 );
    or g20418 ( n36424 , n26286 , n5904 );
    or g20419 ( n40584 , n7690 , n3103 );
    not g20420 ( n7384 , n21909 );
    or g20421 ( n14534 , n40785 , n33778 );
    nor g20422 ( n23041 , n33204 , n10953 );
    and g20423 ( n38999 , n25843 , n34746 );
    and g20424 ( n4171 , n27198 , n31151 );
    xnor g20425 ( n2950 , n542 , n23973 );
    not g20426 ( n21111 , n7508 );
    not g20427 ( n3313 , n40701 );
    not g20428 ( n38691 , n31122 );
    not g20429 ( n1495 , n36021 );
    and g20430 ( n16863 , n29602 , n298 );
    or g20431 ( n5711 , n3669 , n11084 );
    not g20432 ( n25985 , n23681 );
    and g20433 ( n34738 , n41647 , n21793 );
    and g20434 ( n19919 , n16629 , n34265 );
    and g20435 ( n11871 , n35716 , n22940 );
    or g20436 ( n20643 , n37562 , n31949 );
    and g20437 ( n15198 , n6989 , n12668 );
    nor g20438 ( n40521 , n40210 , n3120 );
    and g20439 ( n40400 , n8820 , n1939 );
    not g20440 ( n5 , n19154 );
    nor g20441 ( n1591 , n37692 , n17627 );
    and g20442 ( n3862 , n34461 , n23243 );
    nor g20443 ( n10934 , n13332 , n34095 );
    and g20444 ( n1123 , n24989 , n29391 );
    xnor g20445 ( n24620 , n39286 , n2199 );
    or g20446 ( n31257 , n13709 , n17903 );
    and g20447 ( n13530 , n21704 , n7204 );
    and g20448 ( n21708 , n38341 , n3956 );
    and g20449 ( n37043 , n41656 , n4247 );
    not g20450 ( n4625 , n5254 );
    and g20451 ( n14290 , n33329 , n11570 );
    or g20452 ( n23652 , n14107 , n20148 );
    or g20453 ( n24761 , n17488 , n34972 );
    or g20454 ( n34898 , n23295 , n12758 );
    not g20455 ( n22160 , n26245 );
    and g20456 ( n28565 , n11449 , n6171 );
    or g20457 ( n29622 , n15423 , n40477 );
    nor g20458 ( n1317 , n12208 , n35627 );
    and g20459 ( n28908 , n31276 , n1467 );
    not g20460 ( n38020 , n20228 );
    or g20461 ( n33386 , n37438 , n35043 );
    and g20462 ( n10337 , n9123 , n37440 );
    and g20463 ( n2582 , n33771 , n21657 );
    nor g20464 ( n10029 , n17049 , n32167 );
    and g20465 ( n36972 , n86 , n2159 );
    or g20466 ( n26666 , n38269 , n40400 );
    or g20467 ( n21616 , n20666 , n23261 );
    and g20468 ( n14259 , n31243 , n7939 );
    and g20469 ( n29343 , n39584 , n16457 );
    not g20470 ( n17321 , n13979 );
    not g20471 ( n32539 , n36132 );
    xnor g20472 ( n11502 , n25619 , n5741 );
    or g20473 ( n20449 , n28335 , n1299 );
    or g20474 ( n16861 , n21646 , n10898 );
    and g20475 ( n35960 , n1625 , n21124 );
    xnor g20476 ( n3074 , n11109 , n20399 );
    or g20477 ( n31163 , n33819 , n714 );
    or g20478 ( n39396 , n11569 , n32091 );
    and g20479 ( n19064 , n16776 , n17622 );
    or g20480 ( n27810 , n39150 , n23335 );
    xnor g20481 ( n11166 , n29098 , n40272 );
    not g20482 ( n22973 , n11351 );
    or g20483 ( n11898 , n841 , n21807 );
    not g20484 ( n3225 , n27750 );
    nor g20485 ( n16433 , n25404 , n17628 );
    nor g20486 ( n12113 , n4173 , n18421 );
    or g20487 ( n13801 , n37520 , n34136 );
    or g20488 ( n31131 , n1995 , n29484 );
    nor g20489 ( n35479 , n10592 , n40478 );
    and g20490 ( n15571 , n41547 , n3551 );
    not g20491 ( n295 , n34931 );
    not g20492 ( n14053 , n25594 );
    or g20493 ( n23442 , n12588 , n35747 );
    and g20494 ( n22349 , n39689 , n12494 );
    not g20495 ( n40255 , n41769 );
    xnor g20496 ( n6836 , n11886 , n42836 );
    and g20497 ( n30583 , n34617 , n13891 );
    xnor g20498 ( n713 , n34906 , n8494 );
    or g20499 ( n32817 , n3225 , n4990 );
    or g20500 ( n39163 , n14483 , n25115 );
    or g20501 ( n33057 , n8539 , n39830 );
    not g20502 ( n32887 , n30611 );
    nor g20503 ( n35129 , n33732 , n2953 );
    or g20504 ( n12439 , n27812 , n32980 );
    or g20505 ( n31393 , n23538 , n5974 );
    or g20506 ( n27373 , n13160 , n14677 );
    nor g20507 ( n7928 , n41941 , n10685 );
    or g20508 ( n36691 , n3402 , n7737 );
    or g20509 ( n30723 , n8967 , n553 );
    xnor g20510 ( n13685 , n35316 , n8043 );
    nor g20511 ( n5651 , n20432 , n13283 );
    or g20512 ( n31537 , n13387 , n34131 );
    xnor g20513 ( n7557 , n40762 , n25074 );
    not g20514 ( n38886 , n38898 );
    nor g20515 ( n4176 , n11451 , n34694 );
    or g20516 ( n5699 , n25821 , n42274 );
    and g20517 ( n287 , n31479 , n20987 );
    nor g20518 ( n39206 , n3181 , n39485 );
    not g20519 ( n81 , n32778 );
    xnor g20520 ( n7760 , n18859 , n37803 );
    and g20521 ( n21444 , n41899 , n8667 );
    xnor g20522 ( n13796 , n22263 , n15473 );
    or g20523 ( n17878 , n5639 , n11361 );
    nor g20524 ( n40520 , n9336 , n13480 );
    nor g20525 ( n42664 , n37079 , n38118 );
    xnor g20526 ( n9959 , n34875 , n17221 );
    or g20527 ( n31936 , n313 , n30304 );
    or g20528 ( n41470 , n20822 , n31950 );
    or g20529 ( n23370 , n25078 , n40068 );
    or g20530 ( n15586 , n7356 , n13172 );
    or g20531 ( n11550 , n38035 , n28920 );
    or g20532 ( n717 , n19683 , n2591 );
    or g20533 ( n29410 , n14766 , n31271 );
    and g20534 ( n35823 , n12365 , n31705 );
    nor g20535 ( n27799 , n33981 , n18471 );
    and g20536 ( n20232 , n27174 , n13987 );
    and g20537 ( n29703 , n15826 , n21935 );
    nor g20538 ( n23116 , n14969 , n33487 );
    and g20539 ( n38510 , n15828 , n40791 );
    and g20540 ( n19140 , n41834 , n34348 );
    and g20541 ( n19852 , n603 , n9620 );
    not g20542 ( n19780 , n40096 );
    and g20543 ( n13912 , n35720 , n16642 );
    xnor g20544 ( n10696 , n3013 , n40892 );
    nor g20545 ( n17555 , n16649 , n13757 );
    nor g20546 ( n521 , n33190 , n10719 );
    xnor g20547 ( n16033 , n2183 , n29598 );
    xnor g20548 ( n18382 , n26579 , n7498 );
    nor g20549 ( n19393 , n9607 , n25161 );
    and g20550 ( n27110 , n38422 , n3875 );
    xnor g20551 ( n2714 , n41718 , n35100 );
    and g20552 ( n24497 , n19377 , n23630 );
    and g20553 ( n20402 , n16041 , n17666 );
    or g20554 ( n31754 , n19005 , n27179 );
    not g20555 ( n27484 , n29567 );
    and g20556 ( n14126 , n42834 , n16737 );
    xnor g20557 ( n40967 , n36009 , n22060 );
    or g20558 ( n7303 , n32749 , n14553 );
    or g20559 ( n41265 , n42896 , n18097 );
    or g20560 ( n27256 , n28551 , n26433 );
    or g20561 ( n9602 , n1905 , n17321 );
    or g20562 ( n32931 , n8494 , n1113 );
    not g20563 ( n783 , n27415 );
    or g20564 ( n25683 , n6929 , n30937 );
    or g20565 ( n30229 , n19152 , n40526 );
    not g20566 ( n1989 , n34976 );
    xnor g20567 ( n39575 , n7180 , n18836 );
    or g20568 ( n24730 , n27425 , n16537 );
    and g20569 ( n189 , n35942 , n13589 );
    or g20570 ( n5689 , n1499 , n39761 );
    or g20571 ( n24069 , n13049 , n21850 );
    xnor g20572 ( n10739 , n28464 , n38505 );
    and g20573 ( n1004 , n8862 , n28370 );
    or g20574 ( n32864 , n2213 , n36198 );
    or g20575 ( n33668 , n20145 , n29519 );
    or g20576 ( n36764 , n35061 , n39050 );
    or g20577 ( n39110 , n220 , n42522 );
    xnor g20578 ( n41729 , n38554 , n1507 );
    not g20579 ( n26691 , n27419 );
    nor g20580 ( n29846 , n13604 , n4267 );
    or g20581 ( n19743 , n24386 , n30584 );
    or g20582 ( n39102 , n14070 , n19750 );
    or g20583 ( n23227 , n1071 , n22462 );
    and g20584 ( n17062 , n13458 , n13451 );
    or g20585 ( n24661 , n33572 , n32100 );
    or g20586 ( n33003 , n41767 , n30232 );
    or g20587 ( n27236 , n9319 , n6834 );
    xnor g20588 ( n20558 , n3486 , n6450 );
    and g20589 ( n19182 , n38413 , n33183 );
    or g20590 ( n18717 , n8891 , n35531 );
    or g20591 ( n41775 , n29104 , n24727 );
    or g20592 ( n4115 , n14622 , n39688 );
    or g20593 ( n19853 , n2332 , n35695 );
    or g20594 ( n4210 , n39850 , n6267 );
    xnor g20595 ( n22046 , n35259 , n29017 );
    and g20596 ( n5131 , n17929 , n34851 );
    or g20597 ( n42621 , n3726 , n30763 );
    or g20598 ( n18985 , n33981 , n28221 );
    xnor g20599 ( n29928 , n30429 , n9277 );
    xnor g20600 ( n36819 , n18297 , n18416 );
    xnor g20601 ( n14654 , n34562 , n4486 );
    and g20602 ( n9782 , n26176 , n40050 );
    not g20603 ( n1493 , n588 );
    or g20604 ( n534 , n19054 , n33977 );
    xnor g20605 ( n26772 , n15891 , n39907 );
    and g20606 ( n28223 , n33814 , n8706 );
    not g20607 ( n5768 , n34330 );
    or g20608 ( n42640 , n11461 , n22598 );
    or g20609 ( n37814 , n33330 , n37047 );
    or g20610 ( n11250 , n25596 , n1057 );
    xnor g20611 ( n39027 , n16732 , n29467 );
    and g20612 ( n41885 , n25527 , n8215 );
    xnor g20613 ( n8872 , n11595 , n33494 );
    xnor g20614 ( n31054 , n5891 , n14711 );
    and g20615 ( n5908 , n24002 , n16681 );
    or g20616 ( n7602 , n21706 , n26363 );
    not g20617 ( n2722 , n28530 );
    xnor g20618 ( n30194 , n36704 , n21748 );
    xnor g20619 ( n298 , n39178 , n15085 );
    not g20620 ( n15356 , n21975 );
    xnor g20621 ( n13579 , n2338 , n2277 );
    or g20622 ( n15424 , n8184 , n33345 );
    not g20623 ( n18491 , n26373 );
    not g20624 ( n42710 , n32520 );
    or g20625 ( n22376 , n33464 , n7367 );
    nor g20626 ( n8512 , n34292 , n11208 );
    or g20627 ( n40288 , n28461 , n35801 );
    or g20628 ( n9105 , n41977 , n21085 );
    nor g20629 ( n11498 , n18550 , n10350 );
    or g20630 ( n32908 , n25837 , n14743 );
    or g20631 ( n19091 , n6578 , n4726 );
    xnor g20632 ( n23099 , n33314 , n41314 );
    or g20633 ( n26152 , n37230 , n20799 );
    xnor g20634 ( n27621 , n25020 , n17417 );
    and g20635 ( n15952 , n16053 , n17897 );
    or g20636 ( n2653 , n36272 , n39221 );
    or g20637 ( n39889 , n41356 , n36700 );
    or g20638 ( n21694 , n7242 , n24230 );
    or g20639 ( n13996 , n30569 , n19493 );
    and g20640 ( n16354 , n39488 , n20758 );
    and g20641 ( n13861 , n20997 , n40230 );
    and g20642 ( n23750 , n30314 , n7422 );
    xnor g20643 ( n8508 , n5144 , n24162 );
    or g20644 ( n8628 , n23249 , n5578 );
    and g20645 ( n17452 , n3489 , n7724 );
    or g20646 ( n40324 , n35372 , n41684 );
    nor g20647 ( n13390 , n22607 , n1607 );
    and g20648 ( n13115 , n24385 , n126 );
    not g20649 ( n42124 , n37095 );
    not g20650 ( n7069 , n24447 );
    xnor g20651 ( n39117 , n36876 , n28719 );
    xnor g20652 ( n34279 , n7943 , n8344 );
    or g20653 ( n25457 , n8098 , n16851 );
    or g20654 ( n10459 , n29803 , n16321 );
    or g20655 ( n1402 , n40785 , n8832 );
    or g20656 ( n24514 , n8561 , n26459 );
    not g20657 ( n26210 , n3759 );
    or g20658 ( n8018 , n8967 , n31141 );
    or g20659 ( n11073 , n25817 , n32348 );
    and g20660 ( n22499 , n2166 , n3810 );
    and g20661 ( n30704 , n34538 , n31821 );
    xnor g20662 ( n39209 , n35217 , n21910 );
    or g20663 ( n41383 , n465 , n10790 );
    or g20664 ( n20221 , n34361 , n30331 );
    or g20665 ( n40410 , n14749 , n40736 );
    nor g20666 ( n27752 , n38350 , n22004 );
    xnor g20667 ( n15745 , n38679 , n8505 );
    nor g20668 ( n9314 , n16598 , n28483 );
    xnor g20669 ( n20329 , n25985 , n232 );
    or g20670 ( n9548 , n37980 , n5802 );
    and g20671 ( n23274 , n30560 , n24465 );
    not g20672 ( n6362 , n27550 );
    not g20673 ( n33532 , n17566 );
    or g20674 ( n31792 , n18951 , n25026 );
    or g20675 ( n21724 , n25650 , n33450 );
    or g20676 ( n37201 , n42202 , n31503 );
    and g20677 ( n16421 , n31299 , n23121 );
    and g20678 ( n27618 , n9959 , n34372 );
    xnor g20679 ( n36364 , n1219 , n36771 );
    or g20680 ( n20064 , n23694 , n18402 );
    or g20681 ( n3224 , n37029 , n3816 );
    or g20682 ( n14050 , n14048 , n3641 );
    nor g20683 ( n8913 , n30166 , n23254 );
    or g20684 ( n11086 , n31850 , n20098 );
    or g20685 ( n37825 , n15681 , n38611 );
    not g20686 ( n16141 , n1925 );
    nor g20687 ( n20427 , n35678 , n11749 );
    nor g20688 ( n14705 , n28710 , n23102 );
    or g20689 ( n13844 , n2582 , n29058 );
    or g20690 ( n18168 , n14431 , n4849 );
    nor g20691 ( n19637 , n40210 , n8536 );
    and g20692 ( n37706 , n32107 , n10382 );
    xnor g20693 ( n32291 , n31048 , n10433 );
    xnor g20694 ( n32709 , n35422 , n2199 );
    or g20695 ( n31712 , n27646 , n28950 );
    and g20696 ( n15216 , n3169 , n36728 );
    and g20697 ( n37817 , n26141 , n34747 );
    and g20698 ( n11906 , n16411 , n22267 );
    or g20699 ( n34814 , n19829 , n4926 );
    not g20700 ( n21380 , n791 );
    or g20701 ( n31397 , n13907 , n22419 );
    xnor g20702 ( n16917 , n13136 , n37714 );
    not g20703 ( n19952 , n18792 );
    and g20704 ( n19171 , n25362 , n21467 );
    nor g20705 ( n30130 , n36117 , n18788 );
    or g20706 ( n31987 , n9199 , n13141 );
    or g20707 ( n31555 , n6430 , n18945 );
    xnor g20708 ( n19689 , n19463 , n4630 );
    and g20709 ( n37360 , n27204 , n35855 );
    or g20710 ( n19640 , n21907 , n35090 );
    xnor g20711 ( n13245 , n15972 , n13664 );
    or g20712 ( n8640 , n9066 , n18165 );
    and g20713 ( n24251 , n41582 , n35600 );
    or g20714 ( n32680 , n1968 , n41328 );
    nor g20715 ( n28642 , n1301 , n26931 );
    not g20716 ( n16152 , n15460 );
    not g20717 ( n19629 , n9116 );
    and g20718 ( n35138 , n19008 , n15761 );
    and g20719 ( n13569 , n39845 , n11517 );
    or g20720 ( n40177 , n20412 , n15695 );
    nor g20721 ( n1155 , n4852 , n35208 );
    and g20722 ( n6195 , n39774 , n38275 );
    or g20723 ( n29732 , n14481 , n12963 );
    or g20724 ( n7730 , n37669 , n8401 );
    and g20725 ( n33010 , n21079 , n35825 );
    or g20726 ( n33961 , n24775 , n37678 );
    xnor g20727 ( n12358 , n965 , n17975 );
    or g20728 ( n38728 , n30696 , n24823 );
    or g20729 ( n19160 , n42450 , n6359 );
    or g20730 ( n9095 , n42174 , n19675 );
    or g20731 ( n36066 , n40786 , n13628 );
    or g20732 ( n39071 , n19449 , n11825 );
    and g20733 ( n6372 , n40161 , n3304 );
    or g20734 ( n9055 , n14546 , n40259 );
    or g20735 ( n11733 , n11546 , n32312 );
    xnor g20736 ( n35132 , n22014 , n12630 );
    or g20737 ( n3081 , n14110 , n31393 );
    or g20738 ( n27461 , n38622 , n22355 );
    or g20739 ( n13494 , n42513 , n14686 );
    and g20740 ( n24737 , n31179 , n38177 );
    nor g20741 ( n14883 , n8229 , n13831 );
    xnor g20742 ( n20907 , n24339 , n20753 );
    or g20743 ( n23956 , n972 , n29984 );
    nor g20744 ( n5154 , n17583 , n12562 );
    nor g20745 ( n17286 , n27387 , n35939 );
    xnor g20746 ( n33133 , n27081 , n22559 );
    and g20747 ( n18908 , n3734 , n23129 );
    not g20748 ( n27543 , n9501 );
    and g20749 ( n39033 , n10312 , n15036 );
    or g20750 ( n30542 , n3943 , n34195 );
    or g20751 ( n10552 , n41210 , n11868 );
    and g20752 ( n8092 , n22921 , n6614 );
    xnor g20753 ( n21858 , n9775 , n30086 );
    or g20754 ( n25085 , n36502 , n487 );
    or g20755 ( n18623 , n20152 , n42479 );
    or g20756 ( n22763 , n39851 , n4015 );
    and g20757 ( n27699 , n6312 , n32268 );
    or g20758 ( n8120 , n13282 , n26755 );
    xnor g20759 ( n19763 , n9113 , n1608 );
    and g20760 ( n6027 , n7803 , n33573 );
    or g20761 ( n6777 , n3420 , n16657 );
    and g20762 ( n14982 , n10761 , n15503 );
    and g20763 ( n38268 , n6369 , n27787 );
    or g20764 ( n23999 , n36891 , n14427 );
    not g20765 ( n24159 , n29457 );
    or g20766 ( n17447 , n10875 , n12129 );
    or g20767 ( n34610 , n35387 , n36599 );
    nor g20768 ( n37460 , n15403 , n24905 );
    or g20769 ( n33391 , n20583 , n34821 );
    or g20770 ( n33723 , n34513 , n42856 );
    not g20771 ( n7443 , n3265 );
    or g20772 ( n9589 , n29302 , n1280 );
    and g20773 ( n41609 , n39907 , n15891 );
    or g20774 ( n19893 , n6945 , n13397 );
    and g20775 ( n7714 , n20144 , n2690 );
    or g20776 ( n4371 , n38750 , n14487 );
    not g20777 ( n14569 , n39581 );
    not g20778 ( n244 , n38444 );
    not g20779 ( n42830 , n25698 );
    or g20780 ( n18079 , n37263 , n22528 );
    nor g20781 ( n42041 , n19262 , n6425 );
    and g20782 ( n22480 , n23062 , n19889 );
    xnor g20783 ( n21609 , n35477 , n15216 );
    or g20784 ( n3460 , n28912 , n11102 );
    or g20785 ( n14710 , n1735 , n22762 );
    not g20786 ( n708 , n4424 );
    or g20787 ( n13855 , n26173 , n35742 );
    nor g20788 ( n19792 , n27065 , n31839 );
    not g20789 ( n529 , n9828 );
    or g20790 ( n10765 , n33128 , n27712 );
    and g20791 ( n18119 , n24914 , n33581 );
    or g20792 ( n3110 , n16780 , n21782 );
    not g20793 ( n2492 , n30555 );
    nor g20794 ( n20601 , n14707 , n29403 );
    nor g20795 ( n27156 , n5964 , n3975 );
    xnor g20796 ( n22904 , n3277 , n34171 );
    or g20797 ( n13779 , n39266 , n31697 );
    nor g20798 ( n25776 , n27024 , n24489 );
    nor g20799 ( n8766 , n13013 , n13995 );
    and g20800 ( n42409 , n27814 , n13372 );
    or g20801 ( n7416 , n35963 , n9547 );
    or g20802 ( n9618 , n25651 , n19788 );
    and g20803 ( n32787 , n11139 , n37668 );
    and g20804 ( n31875 , n6789 , n38785 );
    or g20805 ( n20625 , n17108 , n20954 );
    and g20806 ( n15250 , n26411 , n5708 );
    and g20807 ( n28097 , n6089 , n12109 );
    and g20808 ( n22487 , n29207 , n36635 );
    or g20809 ( n8079 , n19755 , n40016 );
    or g20810 ( n19817 , n7209 , n10559 );
    or g20811 ( n36020 , n40232 , n38149 );
    nor g20812 ( n21608 , n26612 , n39209 );
    xnor g20813 ( n22011 , n17198 , n30653 );
    or g20814 ( n33968 , n34559 , n24497 );
    or g20815 ( n7677 , n35592 , n26065 );
    nor g20816 ( n528 , n33774 , n23463 );
    nor g20817 ( n15846 , n17744 , n42616 );
    or g20818 ( n13818 , n17657 , n27020 );
    nor g20819 ( n13622 , n28896 , n26825 );
    or g20820 ( n11804 , n14785 , n39741 );
    nor g20821 ( n16427 , n30327 , n26012 );
    and g20822 ( n3049 , n21736 , n30087 );
    nor g20823 ( n4036 , n14471 , n30767 );
    or g20824 ( n42332 , n19194 , n9917 );
    or g20825 ( n27078 , n15983 , n41891 );
    and g20826 ( n40730 , n31796 , n40836 );
    or g20827 ( n22848 , n40180 , n35379 );
    or g20828 ( n18816 , n32195 , n41038 );
    or g20829 ( n8461 , n7009 , n35531 );
    or g20830 ( n36360 , n8417 , n22343 );
    or g20831 ( n21313 , n22091 , n22457 );
    not g20832 ( n32540 , n31481 );
    or g20833 ( n21575 , n23881 , n2599 );
    and g20834 ( n27580 , n38683 , n17920 );
    and g20835 ( n3062 , n26378 , n15357 );
    and g20836 ( n2063 , n14572 , n7808 );
    nor g20837 ( n28501 , n26360 , n6627 );
    or g20838 ( n34451 , n26122 , n38077 );
    or g20839 ( n8397 , n23085 , n34109 );
    and g20840 ( n5741 , n15635 , n38172 );
    not g20841 ( n41517 , n16469 );
    not g20842 ( n3314 , n27635 );
    not g20843 ( n40169 , n4127 );
    and g20844 ( n34743 , n7632 , n20922 );
    not g20845 ( n39581 , n32273 );
    nor g20846 ( n14697 , n38676 , n21113 );
    not g20847 ( n13078 , n11626 );
    or g20848 ( n92 , n10485 , n17822 );
    or g20849 ( n8001 , n40295 , n24140 );
    and g20850 ( n40598 , n31023 , n14003 );
    or g20851 ( n22724 , n2967 , n42544 );
    or g20852 ( n12311 , n1199 , n12256 );
    or g20853 ( n31429 , n994 , n40924 );
    xnor g20854 ( n9268 , n31099 , n18315 );
    and g20855 ( n12980 , n26921 , n29756 );
    nor g20856 ( n38085 , n8494 , n36522 );
    not g20857 ( n16462 , n38635 );
    or g20858 ( n28677 , n42473 , n13150 );
    or g20859 ( n17697 , n28117 , n19841 );
    xnor g20860 ( n37336 , n16532 , n16928 );
    xnor g20861 ( n10195 , n31290 , n24450 );
    or g20862 ( n30831 , n11820 , n35382 );
    and g20863 ( n6900 , n22099 , n21191 );
    xnor g20864 ( n4610 , n36998 , n36862 );
    not g20865 ( n18137 , n15377 );
    not g20866 ( n16899 , n14280 );
    or g20867 ( n224 , n33922 , n36979 );
    not g20868 ( n17956 , n11045 );
    and g20869 ( n20942 , n23023 , n14624 );
    or g20870 ( n2744 , n26244 , n1387 );
    not g20871 ( n25914 , n29217 );
    nor g20872 ( n36660 , n13236 , n40270 );
    or g20873 ( n19147 , n38684 , n38853 );
    or g20874 ( n29280 , n31541 , n4492 );
    and g20875 ( n19734 , n41781 , n8513 );
    xnor g20876 ( n6975 , n32248 , n1258 );
    or g20877 ( n25098 , n26289 , n34140 );
    and g20878 ( n15555 , n20160 , n3364 );
    and g20879 ( n8750 , n21328 , n7703 );
    or g20880 ( n11419 , n37567 , n3916 );
    or g20881 ( n33594 , n9395 , n29322 );
    xnor g20882 ( n16454 , n32297 , n37010 );
    nor g20883 ( n41210 , n33935 , n40509 );
    and g20884 ( n25838 , n24733 , n7599 );
    xnor g20885 ( n30774 , n28614 , n17190 );
    and g20886 ( n6037 , n5360 , n13092 );
    not g20887 ( n11723 , n32572 );
    nor g20888 ( n11260 , n30582 , n102 );
    or g20889 ( n39950 , n37687 , n14090 );
    xnor g20890 ( n24253 , n38679 , n18842 );
    xnor g20891 ( n8493 , n8381 , n34565 );
    nor g20892 ( n30445 , n3826 , n5354 );
    not g20893 ( n41752 , n36488 );
    nor g20894 ( n8138 , n17120 , n27582 );
    not g20895 ( n39223 , n38228 );
    not g20896 ( n31326 , n15589 );
    nor g20897 ( n38632 , n15281 , n27112 );
    not g20898 ( n34992 , n17121 );
    xnor g20899 ( n11398 , n5891 , n37161 );
    or g20900 ( n40257 , n16736 , n19596 );
    or g20901 ( n15046 , n4970 , n18572 );
    nor g20902 ( n10990 , n37042 , n27 );
    nor g20903 ( n31636 , n41071 , n7251 );
    or g20904 ( n13359 , n13529 , n41820 );
    and g20905 ( n19057 , n4225 , n5469 );
    or g20906 ( n28934 , n33124 , n24068 );
    or g20907 ( n33276 , n8085 , n31444 );
    or g20908 ( n27402 , n19857 , n7604 );
    or g20909 ( n38741 , n29200 , n25520 );
    not g20910 ( n37770 , n36488 );
    xnor g20911 ( n12248 , n2205 , n34636 );
    or g20912 ( n6018 , n19655 , n5722 );
    not g20913 ( n4708 , n16552 );
    and g20914 ( n11012 , n26614 , n35925 );
    nor g20915 ( n28514 , n29226 , n19874 );
    and g20916 ( n12638 , n17737 , n16823 );
    or g20917 ( n14497 , n25246 , n3912 );
    not g20918 ( n39705 , n33313 );
    not g20919 ( n2692 , n9304 );
    nor g20920 ( n21802 , n15070 , n33113 );
    or g20921 ( n10578 , n29053 , n42418 );
    or g20922 ( n30688 , n19098 , n32958 );
    or g20923 ( n37930 , n37957 , n12896 );
    or g20924 ( n17402 , n30795 , n20162 );
    not g20925 ( n4548 , n32008 );
    nor g20926 ( n32335 , n5490 , n28844 );
    nor g20927 ( n14087 , n29057 , n26019 );
    and g20928 ( n34473 , n33952 , n34753 );
    and g20929 ( n9256 , n34833 , n20695 );
    not g20930 ( n24389 , n9886 );
    and g20931 ( n4680 , n25177 , n12997 );
    nor g20932 ( n16947 , n35255 , n9461 );
    or g20933 ( n19937 , n10306 , n16729 );
    nor g20934 ( n26471 , n19076 , n4710 );
    and g20935 ( n35907 , n21251 , n36276 );
    not g20936 ( n4154 , n27764 );
    and g20937 ( n1206 , n2651 , n3617 );
    or g20938 ( n9898 , n36585 , n26491 );
    and g20939 ( n12726 , n9481 , n36603 );
    and g20940 ( n10861 , n42868 , n4279 );
    or g20941 ( n16975 , n24885 , n34949 );
    not g20942 ( n35701 , n34104 );
    xnor g20943 ( n29519 , n36829 , n19187 );
    and g20944 ( n9727 , n24803 , n16238 );
    and g20945 ( n11675 , n40638 , n34930 );
    and g20946 ( n166 , n9818 , n24446 );
    or g20947 ( n26059 , n27612 , n39963 );
    or g20948 ( n33823 , n2225 , n26968 );
    xnor g20949 ( n36499 , n13045 , n41658 );
    not g20950 ( n30681 , n7198 );
    nor g20951 ( n7954 , n5041 , n24605 );
    nor g20952 ( n22281 , n2645 , n21923 );
    or g20953 ( n28298 , n33464 , n32959 );
    and g20954 ( n35841 , n41245 , n34436 );
    nor g20955 ( n13322 , n29170 , n30159 );
    or g20956 ( n24066 , n37643 , n11603 );
    nor g20957 ( n32789 , n38879 , n6807 );
    or g20958 ( n17507 , n31286 , n40515 );
    not g20959 ( n1216 , n31089 );
    or g20960 ( n40203 , n17256 , n33032 );
    or g20961 ( n29645 , n11908 , n41147 );
    or g20962 ( n34903 , n36600 , n13213 );
    not g20963 ( n13392 , n25804 );
    or g20964 ( n39500 , n39075 , n26783 );
    or g20965 ( n17731 , n38829 , n32488 );
    nor g20966 ( n5286 , n7489 , n22855 );
    not g20967 ( n9133 , n28632 );
    xnor g20968 ( n18681 , n36444 , n11685 );
    not g20969 ( n2253 , n21303 );
    or g20970 ( n37987 , n244 , n203 );
    nor g20971 ( n36943 , n14370 , n1063 );
    or g20972 ( n25870 , n38977 , n18236 );
    or g20973 ( n38476 , n3073 , n35227 );
    and g20974 ( n13601 , n11486 , n15491 );
    nor g20975 ( n22465 , n26394 , n28488 );
    or g20976 ( n22960 , n6694 , n29101 );
    or g20977 ( n38353 , n8881 , n33330 );
    or g20978 ( n18451 , n7789 , n16082 );
    or g20979 ( n31817 , n16920 , n39270 );
    xnor g20980 ( n37731 , n7904 , n18837 );
    and g20981 ( n14672 , n18680 , n15347 );
    or g20982 ( n35354 , n36687 , n24704 );
    nor g20983 ( n36936 , n18235 , n33709 );
    xnor g20984 ( n21607 , n26131 , n5709 );
    xnor g20985 ( n8241 , n32475 , n41287 );
    xnor g20986 ( n36956 , n42612 , n4175 );
    and g20987 ( n6464 , n35654 , n26300 );
    or g20988 ( n20690 , n34793 , n39885 );
    not g20989 ( n33238 , n21414 );
    or g20990 ( n21255 , n30210 , n20547 );
    nor g20991 ( n19623 , n5679 , n41681 );
    or g20992 ( n18372 , n27147 , n13081 );
    or g20993 ( n35117 , n38266 , n25689 );
    not g20994 ( n18320 , n3209 );
    or g20995 ( n25816 , n23894 , n42568 );
    and g20996 ( n35090 , n26616 , n11080 );
    or g20997 ( n28890 , n34626 , n18541 );
    not g20998 ( n34411 , n19326 );
    or g20999 ( n22430 , n8691 , n433 );
    not g21000 ( n21811 , n39791 );
    nor g21001 ( n175 , n17120 , n27865 );
    or g21002 ( n27963 , n36962 , n10886 );
    or g21003 ( n1843 , n12299 , n2888 );
    nor g21004 ( n40464 , n39571 , n8893 );
    and g21005 ( n32430 , n42578 , n5930 );
    nor g21006 ( n11032 , n13534 , n20276 );
    and g21007 ( n13631 , n23488 , n549 );
    and g21008 ( n16134 , n9254 , n30663 );
    or g21009 ( n39593 , n37647 , n24470 );
    not g21010 ( n12605 , n42204 );
    or g21011 ( n16560 , n15731 , n35530 );
    or g21012 ( n24681 , n34609 , n40036 );
    and g21013 ( n18777 , n37574 , n1835 );
    or g21014 ( n37152 , n41288 , n29546 );
    and g21015 ( n24326 , n14534 , n4634 );
    or g21016 ( n1553 , n42705 , n35319 );
    or g21017 ( n42641 , n6568 , n1416 );
    not g21018 ( n10184 , n10451 );
    and g21019 ( n38297 , n27266 , n15517 );
    not g21020 ( n17564 , n30467 );
    xnor g21021 ( n23120 , n22888 , n32114 );
    and g21022 ( n24015 , n12283 , n11465 );
    or g21023 ( n32067 , n41848 , n19842 );
    nor g21024 ( n17142 , n2183 , n34605 );
    or g21025 ( n27930 , n37973 , n165 );
    and g21026 ( n41780 , n33367 , n10495 );
    xnor g21027 ( n35318 , n41947 , n30802 );
    or g21028 ( n5919 , n13814 , n5813 );
    xnor g21029 ( n18056 , n35361 , n40494 );
    or g21030 ( n32412 , n34640 , n7340 );
    or g21031 ( n24188 , n11496 , n42157 );
    and g21032 ( n16597 , n39160 , n15637 );
    nor g21033 ( n2392 , n7068 , n16118 );
    nor g21034 ( n27573 , n7840 , n41710 );
    or g21035 ( n5865 , n70 , n32410 );
    and g21036 ( n34390 , n37201 , n23294 );
    not g21037 ( n14217 , n42338 );
    xnor g21038 ( n9570 , n41811 , n1286 );
    nor g21039 ( n19795 , n17893 , n33375 );
    or g21040 ( n27748 , n1788 , n15974 );
    not g21041 ( n33935 , n25630 );
    or g21042 ( n15230 , n6286 , n36203 );
    not g21043 ( n5401 , n42547 );
    or g21044 ( n9559 , n4018 , n33629 );
    or g21045 ( n25263 , n4579 , n15573 );
    and g21046 ( n11984 , n12271 , n20097 );
    or g21047 ( n37631 , n12791 , n19842 );
    nor g21048 ( n837 , n19020 , n2379 );
    and g21049 ( n7148 , n26283 , n5241 );
    and g21050 ( n37736 , n33682 , n19236 );
    or g21051 ( n12503 , n39839 , n12045 );
    or g21052 ( n37949 , n12954 , n37648 );
    nor g21053 ( n36913 , n23911 , n34086 );
    or g21054 ( n18045 , n18954 , n13493 );
    not g21055 ( n23377 , n30769 );
    or g21056 ( n30910 , n16562 , n18958 );
    not g21057 ( n16783 , n25757 );
    nor g21058 ( n5463 , n27158 , n18290 );
    nor g21059 ( n29862 , n2074 , n26596 );
    and g21060 ( n27920 , n1359 , n40523 );
    or g21061 ( n41183 , n11655 , n8693 );
    xnor g21062 ( n32392 , n35258 , n14471 );
    not g21063 ( n42801 , n5780 );
    not g21064 ( n23915 , n23150 );
    or g21065 ( n12117 , n23540 , n28028 );
    not g21066 ( n24265 , n27964 );
    and g21067 ( n15925 , n17363 , n25462 );
    and g21068 ( n12288 , n37024 , n5739 );
    nor g21069 ( n16481 , n5998 , n29128 );
    or g21070 ( n16953 , n36837 , n819 );
    nor g21071 ( n2889 , n17302 , n35634 );
    not g21072 ( n2624 , n14779 );
    or g21073 ( n14845 , n18358 , n9918 );
    xnor g21074 ( n13342 , n836 , n20763 );
    or g21075 ( n39912 , n5068 , n15242 );
    or g21076 ( n22754 , n25960 , n37595 );
    nor g21077 ( n11116 , n37582 , n7227 );
    nor g21078 ( n13007 , n22089 , n20373 );
    not g21079 ( n23708 , n20711 );
    or g21080 ( n3281 , n4567 , n2922 );
    or g21081 ( n14943 , n22606 , n8221 );
    or g21082 ( n2869 , n23206 , n26456 );
    and g21083 ( n31829 , n25258 , n36840 );
    nor g21084 ( n17030 , n8453 , n23522 );
    nor g21085 ( n35649 , n21634 , n41443 );
    and g21086 ( n22365 , n812 , n24561 );
    not g21087 ( n11887 , n42842 );
    xnor g21088 ( n31188 , n42060 , n10205 );
    not g21089 ( n10693 , n31119 );
    or g21090 ( n32538 , n33298 , n42544 );
    or g21091 ( n38610 , n20399 , n34652 );
    or g21092 ( n25311 , n8235 , n22901 );
    nor g21093 ( n24052 , n19189 , n41633 );
    not g21094 ( n40136 , n9604 );
    or g21095 ( n19080 , n4311 , n29536 );
    and g21096 ( n2356 , n9449 , n22878 );
    xnor g21097 ( n15836 , n14847 , n25588 );
    and g21098 ( n16046 , n27681 , n4437 );
    or g21099 ( n6190 , n22355 , n20936 );
    or g21100 ( n36648 , n31924 , n2432 );
    or g21101 ( n11333 , n10980 , n38691 );
    not g21102 ( n39150 , n21561 );
    not g21103 ( n16402 , n20946 );
    and g21104 ( n41107 , n12259 , n37492 );
    or g21105 ( n21921 , n41003 , n16915 );
    not g21106 ( n17808 , n28378 );
    or g21107 ( n23863 , n17193 , n13930 );
    not g21108 ( n14481 , n5582 );
    not g21109 ( n10806 , n21178 );
    or g21110 ( n21294 , n3516 , n31475 );
    or g21111 ( n41435 , n14471 , n670 );
    and g21112 ( n8329 , n24077 , n7950 );
    or g21113 ( n24676 , n32277 , n23710 );
    or g21114 ( n11564 , n26953 , n42513 );
    nor g21115 ( n5999 , n7489 , n23725 );
    and g21116 ( n25515 , n21425 , n37359 );
    or g21117 ( n25760 , n8216 , n41993 );
    or g21118 ( n3860 , n3215 , n653 );
    and g21119 ( n2877 , n24584 , n5143 );
    or g21120 ( n926 , n29231 , n17827 );
    or g21121 ( n17202 , n3553 , n13200 );
    or g21122 ( n14907 , n35874 , n19097 );
    or g21123 ( n4690 , n30169 , n5910 );
    or g21124 ( n9999 , n9338 , n2972 );
    or g21125 ( n18309 , n23897 , n13566 );
    or g21126 ( n32443 , n16690 , n6781 );
    not g21127 ( n6543 , n18338 );
    and g21128 ( n17434 , n23597 , n14084 );
    not g21129 ( n36435 , n41225 );
    xnor g21130 ( n3942 , n34562 , n17317 );
    nor g21131 ( n518 , n34618 , n38630 );
    or g21132 ( n24671 , n17548 , n28143 );
    nor g21133 ( n32954 , n31941 , n28463 );
    xnor g21134 ( n35439 , n26579 , n28329 );
    xnor g21135 ( n18261 , n20421 , n35056 );
    or g21136 ( n31380 , n2643 , n30614 );
    or g21137 ( n23072 , n14737 , n41573 );
    or g21138 ( n7334 , n31 , n25437 );
    or g21139 ( n34734 , n1838 , n13294 );
    and g21140 ( n34984 , n947 , n15422 );
    or g21141 ( n27581 , n26498 , n35834 );
    and g21142 ( n35467 , n33758 , n39497 );
    xnor g21143 ( n39418 , n40 , n29344 );
    not g21144 ( n26558 , n18090 );
    or g21145 ( n41537 , n2199 , n35422 );
    and g21146 ( n14685 , n9294 , n37668 );
    not g21147 ( n38766 , n40731 );
    or g21148 ( n21233 , n18953 , n40347 );
    nor g21149 ( n18214 , n38796 , n10294 );
    xnor g21150 ( n6868 , n18466 , n29829 );
    xnor g21151 ( n13307 , n13735 , n22145 );
    or g21152 ( n7763 , n39266 , n40826 );
    or g21153 ( n20251 , n22179 , n328 );
    xnor g21154 ( n2987 , n40601 , n28233 );
    not g21155 ( n20720 , n11666 );
    and g21156 ( n23214 , n42698 , n20595 );
    nor g21157 ( n27294 , n3835 , n34119 );
    and g21158 ( n4066 , n14236 , n37950 );
    and g21159 ( n38639 , n4769 , n42107 );
    xnor g21160 ( n4851 , n9180 , n36861 );
    or g21161 ( n6239 , n2588 , n10555 );
    and g21162 ( n17940 , n13287 , n27282 );
    not g21163 ( n4281 , n15110 );
    not g21164 ( n39141 , n31112 );
    and g21165 ( n19261 , n30389 , n14864 );
    or g21166 ( n27224 , n9264 , n11774 );
    and g21167 ( n19615 , n4676 , n39 );
    not g21168 ( n12497 , n30459 );
    and g21169 ( n23496 , n5021 , n12239 );
    or g21170 ( n38158 , n3951 , n5879 );
    or g21171 ( n18331 , n31568 , n28922 );
    nor g21172 ( n7847 , n26609 , n12839 );
    not g21173 ( n20766 , n37041 );
    not g21174 ( n18924 , n4212 );
    or g21175 ( n22749 , n30360 , n25967 );
    not g21176 ( n11319 , n35871 );
    and g21177 ( n5328 , n29961 , n7245 );
    not g21178 ( n12112 , n3465 );
    and g21179 ( n32494 , n18923 , n38315 );
    nor g21180 ( n34855 , n42110 , n30874 );
    not g21181 ( n39328 , n35103 );
    not g21182 ( n10677 , n39947 );
    and g21183 ( n13512 , n4514 , n23020 );
    not g21184 ( n31433 , n14925 );
    or g21185 ( n20482 , n25136 , n37199 );
    or g21186 ( n18460 , n1980 , n29165 );
    or g21187 ( n4808 , n42770 , n20145 );
    or g21188 ( n17326 , n12103 , n17353 );
    xnor g21189 ( n2482 , n24165 , n28417 );
    xnor g21190 ( n7008 , n4345 , n36550 );
    xnor g21191 ( n41620 , n28836 , n9118 );
    or g21192 ( n24906 , n18301 , n30648 );
    nor g21193 ( n10829 , n7566 , n42121 );
    and g21194 ( n19215 , n4427 , n859 );
    xnor g21195 ( n36886 , n27907 , n33008 );
    xnor g21196 ( n40432 , n27694 , n33784 );
    or g21197 ( n38949 , n38196 , n9087 );
    not g21198 ( n23710 , n6144 );
    xnor g21199 ( n38481 , n1656 , n5265 );
    xnor g21200 ( n26477 , n22879 , n2643 );
    nor g21201 ( n8062 , n16573 , n30470 );
    xnor g21202 ( n16023 , n36009 , n6400 );
    nor g21203 ( n1905 , n34973 , n35326 );
    xnor g21204 ( n41643 , n6110 , n14471 );
    not g21205 ( n16773 , n24722 );
    xnor g21206 ( n41636 , n9142 , n32856 );
    or g21207 ( n31891 , n7168 , n30334 );
    or g21208 ( n31583 , n39656 , n39716 );
    xnor g21209 ( n14305 , n18146 , n25579 );
    nor g21210 ( n7816 , n38989 , n12472 );
    or g21211 ( n41889 , n13830 , n35990 );
    or g21212 ( n37355 , n17967 , n16801 );
    or g21213 ( n6396 , n37557 , n39924 );
    not g21214 ( n35754 , n5799 );
    not g21215 ( n24750 , n11353 );
    and g21216 ( n23125 , n38920 , n16461 );
    and g21217 ( n20636 , n31112 , n25214 );
    and g21218 ( n753 , n19118 , n36317 );
    not g21219 ( n41615 , n35689 );
    and g21220 ( n30977 , n6191 , n21482 );
    and g21221 ( n1988 , n39414 , n38248 );
    and g21222 ( n22889 , n16419 , n13133 );
    nor g21223 ( n1680 , n15198 , n41619 );
    not g21224 ( n36620 , n42824 );
    not g21225 ( n4022 , n8351 );
    or g21226 ( n36866 , n22091 , n9467 );
    xnor g21227 ( n36969 , n13597 , n19333 );
    and g21228 ( n9042 , n41179 , n41576 );
    and g21229 ( n16756 , n7124 , n42024 );
    and g21230 ( n39647 , n7200 , n40040 );
    or g21231 ( n27731 , n9508 , n35459 );
    nor g21232 ( n20183 , n4896 , n39201 );
    and g21233 ( n15498 , n33525 , n21348 );
    xnor g21234 ( n6398 , n24409 , n25823 );
    or g21235 ( n15217 , n32866 , n32063 );
    or g21236 ( n19516 , n8086 , n803 );
    nor g21237 ( n13739 , n6929 , n21013 );
    and g21238 ( n22844 , n17713 , n32823 );
    or g21239 ( n6452 , n34858 , n33820 );
    xnor g21240 ( n24980 , n28225 , n3356 );
    and g21241 ( n36897 , n14907 , n33839 );
    or g21242 ( n1565 , n1917 , n25485 );
    or g21243 ( n2233 , n8538 , n3543 );
    and g21244 ( n8011 , n11188 , n16137 );
    nor g21245 ( n2170 , n30006 , n22047 );
    and g21246 ( n13545 , n5904 , n33983 );
    and g21247 ( n4621 , n41846 , n41976 );
    or g21248 ( n28590 , n32575 , n36962 );
    xnor g21249 ( n12135 , n105 , n3694 );
    not g21250 ( n39675 , n22444 );
    not g21251 ( n32618 , n4652 );
    or g21252 ( n11666 , n35882 , n6770 );
    or g21253 ( n6450 , n14179 , n12203 );
    and g21254 ( n15937 , n22697 , n28282 );
    and g21255 ( n17486 , n37396 , n29566 );
    or g21256 ( n42098 , n23509 , n34410 );
    or g21257 ( n10749 , n11453 , n29774 );
    or g21258 ( n10894 , n6636 , n4002 );
    or g21259 ( n32568 , n28468 , n12018 );
    or g21260 ( n35507 , n21572 , n36221 );
    not g21261 ( n18436 , n42141 );
    or g21262 ( n4733 , n27438 , n10953 );
    nor g21263 ( n22664 , n20698 , n18761 );
    and g21264 ( n30842 , n4906 , n23418 );
    or g21265 ( n27038 , n6011 , n41461 );
    and g21266 ( n36226 , n2183 , n27167 );
    nor g21267 ( n16654 , n15070 , n16591 );
    xnor g21268 ( n28123 , n25448 , n19221 );
    or g21269 ( n8548 , n33318 , n6753 );
    nor g21270 ( n12103 , n16598 , n26675 );
    or g21271 ( n37351 , n16365 , n7786 );
    xnor g21272 ( n24863 , n30513 , n431 );
    xnor g21273 ( n22162 , n4302 , n27121 );
    or g21274 ( n8846 , n40825 , n19041 );
    and g21275 ( n37025 , n15579 , n9782 );
    or g21276 ( n14887 , n30235 , n21677 );
    or g21277 ( n7018 , n33468 , n5258 );
    nor g21278 ( n27568 , n26964 , n2511 );
    xnor g21279 ( n30127 , n14932 , n12778 );
    and g21280 ( n33788 , n11161 , n10759 );
    and g21281 ( n11639 , n7523 , n11463 );
    or g21282 ( n9394 , n29848 , n15299 );
    not g21283 ( n330 , n10943 );
    or g21284 ( n22301 , n34565 , n11651 );
    and g21285 ( n18055 , n35675 , n15128 );
    xnor g21286 ( n25559 , n24745 , n4321 );
    or g21287 ( n12333 , n5910 , n796 );
    nor g21288 ( n42214 , n15156 , n40565 );
    or g21289 ( n24540 , n34244 , n4602 );
    or g21290 ( n5862 , n14696 , n29106 );
    and g21291 ( n12355 , n19835 , n35693 );
    not g21292 ( n38484 , n19006 );
    xnor g21293 ( n16979 , n5144 , n18114 );
    or g21294 ( n1130 , n31373 , n9661 );
    or g21295 ( n31402 , n38347 , n42289 );
    or g21296 ( n18036 , n2599 , n34534 );
    or g21297 ( n18459 , n13909 , n27241 );
    not g21298 ( n37045 , n4943 );
    not g21299 ( n31157 , n28269 );
    or g21300 ( n40526 , n39779 , n38293 );
    and g21301 ( n27526 , n25860 , n21403 );
    not g21302 ( n12348 , n30942 );
    not g21303 ( n30397 , n24800 );
    and g21304 ( n10080 , n15464 , n21010 );
    nor g21305 ( n28954 , n34292 , n2666 );
    not g21306 ( n38122 , n17025 );
    not g21307 ( n37116 , n26046 );
    and g21308 ( n35068 , n34519 , n19834 );
    nor g21309 ( n33378 , n37148 , n11252 );
    xnor g21310 ( n3608 , n7922 , n21390 );
    and g21311 ( n25180 , n23598 , n18605 );
    or g21312 ( n15969 , n28407 , n23467 );
    or g21313 ( n20009 , n17460 , n12210 );
    or g21314 ( n37087 , n39014 , n629 );
    or g21315 ( n38700 , n35360 , n19826 );
    not g21316 ( n28051 , n426 );
    and g21317 ( n21994 , n38249 , n26274 );
    not g21318 ( n6114 , n22444 );
    or g21319 ( n24376 , n41049 , n38006 );
    not g21320 ( n2 , n11284 );
    not g21321 ( n12011 , n23168 );
    or g21322 ( n3743 , n2648 , n12153 );
    or g21323 ( n37611 , n41526 , n16020 );
    or g21324 ( n17552 , n17193 , n2791 );
    or g21325 ( n18111 , n34762 , n16548 );
    or g21326 ( n41310 , n16598 , n8346 );
    or g21327 ( n30731 , n5643 , n38167 );
    not g21328 ( n33545 , n18800 );
    or g21329 ( n22887 , n35464 , n16332 );
    and g21330 ( n32244 , n4450 , n17775 );
    or g21331 ( n19942 , n186 , n41699 );
    or g21332 ( n26038 , n183 , n7616 );
    or g21333 ( n17650 , n18486 , n33671 );
    or g21334 ( n14818 , n24178 , n10032 );
    not g21335 ( n17833 , n41867 );
    and g21336 ( n11038 , n38071 , n40928 );
    and g21337 ( n22291 , n7529 , n26467 );
    or g21338 ( n22809 , n2333 , n41705 );
    and g21339 ( n25116 , n40583 , n37432 );
    and g21340 ( n8239 , n21456 , n29954 );
    xnor g21341 ( n13842 , n30768 , n36812 );
    and g21342 ( n12467 , n28857 , n22571 );
    or g21343 ( n24872 , n19789 , n17104 );
    or g21344 ( n12462 , n24855 , n17528 );
    or g21345 ( n35385 , n32100 , n4955 );
    and g21346 ( n22696 , n30351 , n16868 );
    or g21347 ( n22053 , n13429 , n22956 );
    or g21348 ( n30122 , n30473 , n19958 );
    or g21349 ( n26086 , n22230 , n28473 );
    or g21350 ( n39291 , n21479 , n39177 );
    or g21351 ( n12069 , n41019 , n39355 );
    and g21352 ( n11036 , n13312 , n2359 );
    not g21353 ( n1368 , n30517 );
    and g21354 ( n15992 , n12875 , n34162 );
    nor g21355 ( n17528 , n5168 , n25390 );
    or g21356 ( n4804 , n24077 , n25063 );
    xnor g21357 ( n21952 , n1965 , n8150 );
    and g21358 ( n15112 , n18499 , n29883 );
    or g21359 ( n34564 , n37173 , n21844 );
    nor g21360 ( n38519 , n29255 , n18641 );
    not g21361 ( n5818 , n20151 );
    or g21362 ( n4771 , n2051 , n10629 );
    or g21363 ( n19642 , n19490 , n29890 );
    or g21364 ( n22846 , n8494 , n3855 );
    or g21365 ( n42463 , n34704 , n10069 );
    or g21366 ( n36292 , n38704 , n19601 );
    or g21367 ( n7636 , n14615 , n3170 );
    nor g21368 ( n25487 , n1555 , n704 );
    nor g21369 ( n6033 , n11431 , n6082 );
    nor g21370 ( n31535 , n5871 , n16279 );
    or g21371 ( n39161 , n34273 , n29893 );
    or g21372 ( n25253 , n2959 , n24389 );
    not g21373 ( n13615 , n32284 );
    nor g21374 ( n38865 , n38908 , n2240 );
    or g21375 ( n40269 , n35337 , n38170 );
    and g21376 ( n31760 , n13754 , n4377 );
    and g21377 ( n14459 , n28085 , n7190 );
    not g21378 ( n15016 , n14385 );
    or g21379 ( n32359 , n13892 , n8960 );
    and g21380 ( n1527 , n42443 , n40181 );
    and g21381 ( n32999 , n14274 , n30794 );
    or g21382 ( n2373 , n90 , n3543 );
    xnor g21383 ( n13872 , n40992 , n33690 );
    or g21384 ( n39726 , n3570 , n37147 );
    or g21385 ( n15641 , n25940 , n12073 );
    and g21386 ( n4699 , n26819 , n11399 );
    xnor g21387 ( n30568 , n22263 , n36563 );
    and g21388 ( n15893 , n8450 , n4215 );
    xnor g21389 ( n31643 , n670 , n14471 );
    or g21390 ( n25339 , n31261 , n31720 );
    or g21391 ( n6022 , n27721 , n20431 );
    and g21392 ( n9699 , n20542 , n23387 );
    not g21393 ( n2006 , n11257 );
    not g21394 ( n11134 , n29799 );
    nor g21395 ( n41986 , n405 , n42773 );
    or g21396 ( n30836 , n21465 , n790 );
    nor g21397 ( n11444 , n12105 , n31591 );
    or g21398 ( n13660 , n26116 , n17829 );
    or g21399 ( n26151 , n12859 , n4177 );
    or g21400 ( n39567 , n1296 , n25440 );
    and g21401 ( n34772 , n25913 , n36145 );
    and g21402 ( n6904 , n20419 , n16779 );
    and g21403 ( n16615 , n11127 , n14102 );
    or g21404 ( n8892 , n29264 , n41034 );
    or g21405 ( n2246 , n37809 , n7737 );
    and g21406 ( n40560 , n39543 , n25670 );
    or g21407 ( n1775 , n9035 , n17901 );
    xnor g21408 ( n7777 , n10024 , n20460 );
    not g21409 ( n4823 , n5810 );
    or g21410 ( n29986 , n10918 , n37323 );
    or g21411 ( n41881 , n28402 , n34523 );
    not g21412 ( n3425 , n34014 );
    and g21413 ( n42588 , n31483 , n8600 );
    or g21414 ( n17217 , n40894 , n1735 );
    nor g21415 ( n8029 , n22073 , n33628 );
    not g21416 ( n8747 , n37222 );
    nor g21417 ( n1332 , n21705 , n9179 );
    not g21418 ( n18533 , n10291 );
    and g21419 ( n22955 , n23076 , n12897 );
    not g21420 ( n39927 , n38752 );
    not g21421 ( n32859 , n32115 );
    and g21422 ( n12579 , n27665 , n39582 );
    or g21423 ( n20864 , n30490 , n41062 );
    and g21424 ( n23779 , n37614 , n38834 );
    and g21425 ( n10035 , n35694 , n38180 );
    xnor g21426 ( n5769 , n32624 , n39527 );
    or g21427 ( n1880 , n34634 , n28783 );
    xnor g21428 ( n34210 , n20487 , n23670 );
    or g21429 ( n31684 , n16216 , n34829 );
    or g21430 ( n30954 , n8968 , n17385 );
    or g21431 ( n7606 , n24454 , n25367 );
    or g21432 ( n33508 , n17744 , n15774 );
    or g21433 ( n25530 , n23462 , n34942 );
    or g21434 ( n10158 , n25694 , n13282 );
    or g21435 ( n4516 , n26175 , n19964 );
    and g21436 ( n117 , n10216 , n31344 );
    or g21437 ( n17682 , n22178 , n36882 );
    and g21438 ( n42770 , n24336 , n37672 );
    and g21439 ( n40243 , n13613 , n16777 );
    and g21440 ( n41351 , n35824 , n27428 );
    xnor g21441 ( n4505 , n19591 , n3674 );
    not g21442 ( n4633 , n21440 );
    nor g21443 ( n27175 , n20117 , n37254 );
    nor g21444 ( n17599 , n34519 , n19834 );
    or g21445 ( n40659 , n8220 , n42616 );
    xnor g21446 ( n4060 , n33620 , n17593 );
    not g21447 ( n36792 , n11713 );
    xnor g21448 ( n10157 , n41811 , n10544 );
    nor g21449 ( n11184 , n41662 , n13991 );
    and g21450 ( n22704 , n13608 , n7546 );
    or g21451 ( n17114 , n36869 , n31580 );
    or g21452 ( n4821 , n16588 , n20199 );
    or g21453 ( n6820 , n1269 , n2679 );
    and g21454 ( n36501 , n4120 , n15214 );
    not g21455 ( n18088 , n19382 );
    not g21456 ( n37429 , n21999 );
    or g21457 ( n4925 , n17175 , n20515 );
    nor g21458 ( n35453 , n20573 , n24829 );
    not g21459 ( n26178 , n20511 );
    not g21460 ( n9043 , n31753 );
    and g21461 ( n40339 , n19824 , n37352 );
    not g21462 ( n21150 , n25405 );
    or g21463 ( n19276 , n40271 , n39180 );
    or g21464 ( n38768 , n40703 , n10665 );
    and g21465 ( n20953 , n5517 , n28217 );
    nor g21466 ( n33141 , n38084 , n38833 );
    and g21467 ( n22512 , n39101 , n9572 );
    or g21468 ( n2046 , n28953 , n29930 );
    and g21469 ( n12179 , n16018 , n31877 );
    and g21470 ( n41871 , n6146 , n8259 );
    and g21471 ( n29744 , n26186 , n14521 );
    not g21472 ( n11248 , n34709 );
    not g21473 ( n25948 , n36547 );
    or g21474 ( n28586 , n15134 , n16194 );
    or g21475 ( n1477 , n3635 , n10871 );
    or g21476 ( n37278 , n26741 , n41414 );
    not g21477 ( n40296 , n21293 );
    or g21478 ( n5822 , n13428 , n177 );
    not g21479 ( n34202 , n1568 );
    not g21480 ( n32142 , n41015 );
    and g21481 ( n9718 , n9293 , n21934 );
    or g21482 ( n35912 , n28643 , n1188 );
    nor g21483 ( n41178 , n10598 , n41509 );
    or g21484 ( n26890 , n34331 , n14431 );
    or g21485 ( n14527 , n37330 , n15381 );
    or g21486 ( n30707 , n34491 , n5840 );
    and g21487 ( n2951 , n17953 , n11851 );
    and g21488 ( n38238 , n22522 , n33520 );
    xnor g21489 ( n18066 , n35154 , n35539 );
    or g21490 ( n11842 , n40656 , n7375 );
    and g21491 ( n1891 , n21524 , n10667 );
    or g21492 ( n9592 , n29650 , n23357 );
    or g21493 ( n31887 , n24058 , n38095 );
    and g21494 ( n9720 , n26483 , n22269 );
    not g21495 ( n29276 , n42097 );
    xnor g21496 ( n36876 , n38105 , n17425 );
    or g21497 ( n9173 , n27232 , n22123 );
    and g21498 ( n2302 , n39683 , n28665 );
    not g21499 ( n9881 , n25151 );
    or g21500 ( n32697 , n2212 , n40419 );
    or g21501 ( n37184 , n7765 , n41207 );
    and g21502 ( n29031 , n921 , n19338 );
    xnor g21503 ( n23841 , n27422 , n3266 );
    nor g21504 ( n39533 , n38157 , n17164 );
    or g21505 ( n15964 , n10150 , n5584 );
    and g21506 ( n21668 , n38490 , n7536 );
    nor g21507 ( n32964 , n22719 , n15432 );
    xnor g21508 ( n14402 , n10432 , n17098 );
    nor g21509 ( n35731 , n30059 , n4586 );
    nor g21510 ( n7832 , n19221 , n7061 );
    or g21511 ( n38271 , n15045 , n39096 );
    or g21512 ( n42762 , n15934 , n17183 );
    and g21513 ( n12677 , n42597 , n20833 );
    and g21514 ( n38753 , n11579 , n10500 );
    or g21515 ( n37358 , n177 , n12627 );
    or g21516 ( n16771 , n20699 , n37428 );
    or g21517 ( n42031 , n4972 , n15789 );
    and g21518 ( n11435 , n5435 , n40411 );
    or g21519 ( n16859 , n32350 , n42566 );
    or g21520 ( n40264 , n19260 , n8390 );
    or g21521 ( n42150 , n10491 , n15642 );
    and g21522 ( n8711 , n31341 , n1237 );
    or g21523 ( n37301 , n31144 , n5128 );
    or g21524 ( n24887 , n25175 , n33859 );
    nor g21525 ( n21219 , n7568 , n39248 );
    not g21526 ( n21929 , n30405 );
    or g21527 ( n35430 , n41913 , n19134 );
    nor g21528 ( n19568 , n19262 , n31335 );
    not g21529 ( n24216 , n37811 );
    and g21530 ( n16004 , n12883 , n27 );
    and g21531 ( n41823 , n42215 , n21202 );
    or g21532 ( n461 , n16451 , n20089 );
    or g21533 ( n5807 , n4789 , n17685 );
    xnor g21534 ( n17764 , n9900 , n38897 );
    or g21535 ( n15829 , n30129 , n31324 );
    not g21536 ( n14166 , n32156 );
    nor g21537 ( n7640 , n38295 , n25232 );
    xnor g21538 ( n42132 , n42875 , n5605 );
    not g21539 ( n31850 , n42331 );
    nor g21540 ( n16451 , n5896 , n4101 );
    not g21541 ( n10575 , n18987 );
    or g21542 ( n9737 , n25588 , n23995 );
    xnor g21543 ( n42113 , n10088 , n22868 );
    or g21544 ( n15834 , n23917 , n25341 );
    or g21545 ( n3171 , n29885 , n19100 );
    and g21546 ( n11980 , n1614 , n25476 );
    or g21547 ( n7846 , n41767 , n38401 );
    or g21548 ( n7967 , n16804 , n27833 );
    not g21549 ( n18792 , n2427 );
    or g21550 ( n36664 , n22234 , n35901 );
    not g21551 ( n41995 , n24846 );
    or g21552 ( n11991 , n32217 , n22531 );
    or g21553 ( n7599 , n2111 , n2418 );
    and g21554 ( n41523 , n5024 , n10649 );
    or g21555 ( n29664 , n23462 , n20950 );
    not g21556 ( n29129 , n31352 );
    nor g21557 ( n5754 , n1731 , n11717 );
    or g21558 ( n13542 , n13769 , n39812 );
    or g21559 ( n2231 , n11827 , n25078 );
    or g21560 ( n11102 , n38640 , n36323 );
    or g21561 ( n32342 , n39301 , n32683 );
    and g21562 ( n9225 , n28800 , n17211 );
    nor g21563 ( n37981 , n20167 , n40855 );
    and g21564 ( n29067 , n36884 , n35670 );
    or g21565 ( n9662 , n4694 , n24592 );
    xnor g21566 ( n22320 , n36993 , n19957 );
    xnor g21567 ( n32120 , n34731 , n21283 );
    or g21568 ( n28602 , n19580 , n12968 );
    or g21569 ( n5084 , n25730 , n29217 );
    or g21570 ( n20481 , n9137 , n9663 );
    and g21571 ( n14766 , n38681 , n39073 );
    nor g21572 ( n13517 , n2199 , n24194 );
    or g21573 ( n22731 , n39346 , n42479 );
    and g21574 ( n26561 , n6361 , n34501 );
    or g21575 ( n9818 , n36640 , n18468 );
    or g21576 ( n13567 , n26843 , n39197 );
    xnor g21577 ( n31319 , n9084 , n4752 );
    not g21578 ( n12264 , n24687 );
    not g21579 ( n38249 , n36811 );
    or g21580 ( n23182 , n9554 , n25528 );
    or g21581 ( n5798 , n22278 , n452 );
    nor g21582 ( n40639 , n5896 , n38845 );
    not g21583 ( n42467 , n42813 );
    or g21584 ( n5297 , n32879 , n7531 );
    xnor g21585 ( n23811 , n18530 , n36233 );
    not g21586 ( n31153 , n42821 );
    or g21587 ( n7527 , n34762 , n17859 );
    or g21588 ( n30257 , n11925 , n7428 );
    xnor g21589 ( n29826 , n14217 , n2991 );
    and g21590 ( n35787 , n32523 , n26977 );
    and g21591 ( n10191 , n40327 , n32601 );
    or g21592 ( n14780 , n7113 , n32100 );
    and g21593 ( n32488 , n24473 , n6902 );
    not g21594 ( n27092 , n20777 );
    or g21595 ( n26095 , n35998 , n12048 );
    or g21596 ( n31360 , n41682 , n28190 );
    or g21597 ( n18580 , n27781 , n36971 );
    or g21598 ( n30878 , n30115 , n19041 );
    or g21599 ( n14701 , n32295 , n20503 );
    not g21600 ( n8126 , n23871 );
    nor g21601 ( n41193 , n22753 , n6492 );
    or g21602 ( n37497 , n16146 , n8695 );
    or g21603 ( n23575 , n22157 , n3801 );
    or g21604 ( n22536 , n38487 , n23027 );
    or g21605 ( n21471 , n29339 , n39408 );
    not g21606 ( n27503 , n15778 );
    or g21607 ( n15360 , n27092 , n31218 );
    or g21608 ( n24076 , n15384 , n7719 );
    nor g21609 ( n29688 , n32277 , n14976 );
    not g21610 ( n31825 , n4999 );
    and g21611 ( n6119 , n3996 , n11238 );
    or g21612 ( n6003 , n27264 , n38006 );
    and g21613 ( n32919 , n36960 , n29482 );
    nor g21614 ( n19363 , n30262 , n36128 );
    xnor g21615 ( n10897 , n8057 , n38386 );
    or g21616 ( n10762 , n36796 , n6842 );
    or g21617 ( n37900 , n34705 , n16466 );
    and g21618 ( n17291 , n4759 , n22252 );
    not g21619 ( n14808 , n1954 );
    or g21620 ( n36626 , n32264 , n28413 );
    or g21621 ( n1506 , n1335 , n35072 );
    not g21622 ( n23385 , n8554 );
    not g21623 ( n16369 , n25342 );
    or g21624 ( n4047 , n20818 , n21742 );
    or g21625 ( n13531 , n23201 , n8772 );
    not g21626 ( n37022 , n5974 );
    or g21627 ( n36629 , n3803 , n28913 );
    or g21628 ( n37681 , n11585 , n34075 );
    or g21629 ( n31577 , n6152 , n11533 );
    nor g21630 ( n24142 , n28800 , n17211 );
    or g21631 ( n39229 , n18953 , n2312 );
    xnor g21632 ( n25351 , n19373 , n37810 );
    nor g21633 ( n5500 , n30740 , n11000 );
    and g21634 ( n40823 , n19305 , n4985 );
    or g21635 ( n31056 , n33321 , n670 );
    and g21636 ( n28920 , n8519 , n2663 );
    xnor g21637 ( n29568 , n14315 , n8716 );
    or g21638 ( n39353 , n24441 , n9288 );
    not g21639 ( n14287 , n169 );
    or g21640 ( n27521 , n25968 , n29216 );
    and g21641 ( n12170 , n23831 , n35775 );
    nor g21642 ( n4422 , n36735 , n30180 );
    and g21643 ( n24955 , n12703 , n30923 );
    and g21644 ( n7223 , n30343 , n38092 );
    and g21645 ( n36077 , n29004 , n32899 );
    or g21646 ( n9330 , n39876 , n36153 );
    or g21647 ( n8579 , n42134 , n1044 );
    or g21648 ( n1728 , n39195 , n4069 );
    or g21649 ( n14382 , n36029 , n723 );
    xnor g21650 ( n29784 , n31460 , n35403 );
    xnor g21651 ( n17553 , n7249 , n2952 );
    or g21652 ( n39548 , n35511 , n34960 );
    or g21653 ( n1093 , n3139 , n29607 );
    or g21654 ( n41246 , n22876 , n26545 );
    not g21655 ( n17195 , n38282 );
    not g21656 ( n24605 , n29580 );
    not g21657 ( n12448 , n7692 );
    and g21658 ( n31613 , n16156 , n13245 );
    xnor g21659 ( n27438 , n21858 , n41965 );
    and g21660 ( n18882 , n29867 , n9198 );
    and g21661 ( n15462 , n8279 , n28670 );
    and g21662 ( n1969 , n2097 , n21198 );
    not g21663 ( n33212 , n11354 );
    not g21664 ( n40678 , n10502 );
    and g21665 ( n988 , n28944 , n15939 );
    or g21666 ( n39447 , n13549 , n28065 );
    or g21667 ( n35282 , n21375 , n18070 );
    nor g21668 ( n22535 , n33981 , n37891 );
    and g21669 ( n31751 , n17171 , n14328 );
    and g21670 ( n34258 , n30595 , n7911 );
    and g21671 ( n24318 , n17904 , n40479 );
    xnor g21672 ( n22637 , n31928 , n6798 );
    and g21673 ( n33440 , n16975 , n21454 );
    xnor g21674 ( n21712 , n13183 , n21577 );
    xnor g21675 ( n11781 , n14096 , n27548 );
    and g21676 ( n33387 , n24008 , n5473 );
    nor g21677 ( n37346 , n35301 , n12341 );
    not g21678 ( n8240 , n33807 );
    and g21679 ( n2277 , n35647 , n3377 );
    or g21680 ( n38393 , n17388 , n14057 );
    or g21681 ( n1526 , n42367 , n16765 );
    and g21682 ( n22037 , n27219 , n15782 );
    and g21683 ( n5874 , n19611 , n11509 );
    nor g21684 ( n26170 , n38879 , n28434 );
    or g21685 ( n37490 , n31081 , n19104 );
    and g21686 ( n933 , n14463 , n11455 );
    and g21687 ( n36521 , n29912 , n24198 );
    xnor g21688 ( n559 , n16746 , n21814 );
    nor g21689 ( n36437 , n15070 , n35815 );
    nor g21690 ( n28978 , n37017 , n34407 );
    and g21691 ( n704 , n41296 , n33552 );
    not g21692 ( n16949 , n38734 );
    and g21693 ( n35263 , n30163 , n3881 );
    not g21694 ( n19164 , n13714 );
    or g21695 ( n31549 , n14817 , n21903 );
    and g21696 ( n10570 , n25295 , n11833 );
    or g21697 ( n27177 , n38463 , n2617 );
    and g21698 ( n3406 , n14261 , n25147 );
    xnor g21699 ( n6546 , n33863 , n33247 );
    nor g21700 ( n25640 , n16598 , n5541 );
    xnor g21701 ( n13402 , n26579 , n5551 );
    not g21702 ( n35748 , n1615 );
    not g21703 ( n22979 , n41572 );
    not g21704 ( n17915 , n7217 );
    nor g21705 ( n28549 , n17744 , n37954 );
    and g21706 ( n8341 , n6597 , n34610 );
    nor g21707 ( n2759 , n33654 , n23852 );
    or g21708 ( n26290 , n42159 , n20566 );
    xnor g21709 ( n37630 , n2016 , n17120 );
    and g21710 ( n20729 , n35565 , n41967 );
    or g21711 ( n26560 , n28862 , n23148 );
    not g21712 ( n33570 , n4140 );
    or g21713 ( n40645 , n20498 , n23560 );
    xnor g21714 ( n7097 , n7399 , n8957 );
    or g21715 ( n26497 , n33262 , n2198 );
    and g21716 ( n26971 , n10167 , n22256 );
    and g21717 ( n29338 , n6783 , n31079 );
    or g21718 ( n11323 , n42875 , n5813 );
    nor g21719 ( n27949 , n9113 , n40154 );
    and g21720 ( n34575 , n7777 , n24869 );
    or g21721 ( n31705 , n1702 , n37303 );
    xnor g21722 ( n28905 , n136 , n746 );
    or g21723 ( n10228 , n32797 , n14063 );
    and g21724 ( n37567 , n3847 , n9379 );
    or g21725 ( n41967 , n34917 , n14308 );
    xnor g21726 ( n8728 , n26996 , n41458 );
    xnor g21727 ( n2630 , n13921 , n6872 );
    and g21728 ( n6563 , n12313 , n1963 );
    and g21729 ( n36975 , n2482 , n2930 );
    or g21730 ( n29195 , n25753 , n13633 );
    and g21731 ( n12832 , n30928 , n13242 );
    nor g21732 ( n33694 , n41323 , n40008 );
    or g21733 ( n28247 , n17072 , n3571 );
    or g21734 ( n36703 , n36873 , n30435 );
    and g21735 ( n28651 , n13011 , n34058 );
    and g21736 ( n2835 , n10424 , n33459 );
    or g21737 ( n3753 , n35963 , n40943 );
    nor g21738 ( n6739 , n29098 , n6898 );
    and g21739 ( n34882 , n2264 , n8428 );
    xnor g21740 ( n10991 , n37635 , n13319 );
    xnor g21741 ( n30126 , n28330 , n15070 );
    xnor g21742 ( n38188 , n10834 , n6505 );
    or g21743 ( n2933 , n4044 , n1850 );
    or g21744 ( n27495 , n39266 , n22670 );
    and g21745 ( n40853 , n41929 , n7424 );
    or g21746 ( n39729 , n18002 , n17803 );
    and g21747 ( n3900 , n32593 , n11197 );
    xnor g21748 ( n2281 , n34691 , n1733 );
    or g21749 ( n22826 , n2112 , n21023 );
    xnor g21750 ( n343 , n35102 , n23333 );
    or g21751 ( n19223 , n23005 , n36641 );
    or g21752 ( n40654 , n27761 , n34015 );
    not g21753 ( n4334 , n38157 );
    and g21754 ( n17911 , n20668 , n10221 );
    or g21755 ( n5611 , n26646 , n11718 );
    and g21756 ( n42418 , n15091 , n25396 );
    and g21757 ( n41023 , n26624 , n21377 );
    or g21758 ( n33956 , n38165 , n37778 );
    or g21759 ( n6972 , n40785 , n8527 );
    not g21760 ( n2032 , n22521 );
    not g21761 ( n13886 , n17107 );
    not g21762 ( n20174 , n33545 );
    xnor g21763 ( n35124 , n18471 , n33981 );
    or g21764 ( n15779 , n27862 , n33893 );
    or g21765 ( n23545 , n31789 , n37633 );
    or g21766 ( n34622 , n23216 , n16964 );
    not g21767 ( n6923 , n41919 );
    or g21768 ( n39707 , n7139 , n2035 );
    or g21769 ( n1844 , n28549 , n22750 );
    nor g21770 ( n4128 , n5701 , n17347 );
    or g21771 ( n4748 , n27049 , n36213 );
    or g21772 ( n10277 , n1930 , n34362 );
    not g21773 ( n34782 , n15397 );
    or g21774 ( n16968 , n40323 , n42519 );
    or g21775 ( n41627 , n31436 , n34960 );
    not g21776 ( n10419 , n39166 );
    or g21777 ( n21868 , n9544 , n418 );
    or g21778 ( n15821 , n37878 , n15808 );
    or g21779 ( n16656 , n5910 , n14114 );
    nor g21780 ( n2784 , n35301 , n2454 );
    or g21781 ( n24990 , n4308 , n13453 );
    and g21782 ( n9164 , n37516 , n29201 );
    nor g21783 ( n37308 , n39700 , n20683 );
    or g21784 ( n18843 , n30268 , n31076 );
    nor g21785 ( n35368 , n37052 , n35937 );
    or g21786 ( n2996 , n40608 , n8335 );
    and g21787 ( n34539 , n24205 , n7211 );
    or g21788 ( n2173 , n21004 , n817 );
    nor g21789 ( n12499 , n38157 , n12505 );
    nor g21790 ( n37850 , n13840 , n4508 );
    not g21791 ( n25643 , n35908 );
    xnor g21792 ( n11201 , n30513 , n40088 );
    xnor g21793 ( n42375 , n138 , n17324 );
    not g21794 ( n16117 , n20917 );
    nor g21795 ( n11600 , n7475 , n31165 );
    not g21796 ( n16276 , n26583 );
    or g21797 ( n26745 , n28385 , n34525 );
    and g21798 ( n28986 , n10416 , n39816 );
    nor g21799 ( n34059 , n32423 , n33402 );
    and g21800 ( n26287 , n28618 , n17601 );
    and g21801 ( n23671 , n41267 , n27408 );
    and g21802 ( n1185 , n35612 , n32837 );
    or g21803 ( n16815 , n4554 , n22282 );
    or g21804 ( n22903 , n32113 , n19782 );
    and g21805 ( n13339 , n12294 , n3288 );
    xnor g21806 ( n20652 , n22139 , n7501 );
    not g21807 ( n26230 , n19474 );
    or g21808 ( n1897 , n1457 , n10161 );
    or g21809 ( n15856 , n26252 , n39479 );
    and g21810 ( n39286 , n15969 , n22894 );
    xnor g21811 ( n26892 , n31989 , n35518 );
    xnor g21812 ( n22093 , n7425 , n33776 );
    not g21813 ( n31556 , n39512 );
    nor g21814 ( n27249 , n5615 , n20593 );
    or g21815 ( n2344 , n27840 , n5533 );
    or g21816 ( n19992 , n9701 , n38754 );
    nor g21817 ( n18120 , n18812 , n28780 );
    nor g21818 ( n27172 , n30189 , n40082 );
    or g21819 ( n26736 , n25529 , n17321 );
    or g21820 ( n8861 , n6139 , n16285 );
    or g21821 ( n21842 , n15485 , n6958 );
    not g21822 ( n2368 , n16623 );
    nor g21823 ( n9879 , n32277 , n25789 );
    and g21824 ( n12366 , n28072 , n3244 );
    xnor g21825 ( n2756 , n34037 , n24056 );
    or g21826 ( n34216 , n14490 , n35280 );
    or g21827 ( n3451 , n14894 , n34195 );
    or g21828 ( n26396 , n22849 , n19964 );
    xnor g21829 ( n18227 , n30022 , n42511 );
    or g21830 ( n25079 , n39822 , n37142 );
    nor g21831 ( n15999 , n30108 , n38246 );
    and g21832 ( n19975 , n18513 , n32554 );
    and g21833 ( n34160 , n146 , n32184 );
    and g21834 ( n36870 , n10252 , n6114 );
    or g21835 ( n23728 , n4479 , n10530 );
    and g21836 ( n28727 , n10735 , n11348 );
    not g21837 ( n2517 , n18862 );
    or g21838 ( n12195 , n2512 , n41987 );
    or g21839 ( n30160 , n4085 , n22957 );
    or g21840 ( n10393 , n16598 , n30521 );
    xnor g21841 ( n26844 , n40337 , n40035 );
    not g21842 ( n4335 , n20777 );
    and g21843 ( n27468 , n30915 , n11019 );
    and g21844 ( n11743 , n35185 , n3689 );
    or g21845 ( n6824 , n18517 , n4535 );
    or g21846 ( n10516 , n28932 , n41 );
    or g21847 ( n3866 , n40732 , n2647 );
    not g21848 ( n21634 , n24498 );
    nor g21849 ( n5992 , n25048 , n26181 );
    or g21850 ( n14965 , n30769 , n39446 );
    and g21851 ( n31979 , n15921 , n20493 );
    xnor g21852 ( n10047 , n542 , n5301 );
    and g21853 ( n10531 , n12512 , n24728 );
    nor g21854 ( n31963 , n3944 , n7164 );
    or g21855 ( n35220 , n5863 , n22379 );
    nor g21856 ( n8207 , n32598 , n19154 );
    and g21857 ( n1609 , n4289 , n38780 );
    or g21858 ( n21130 , n41699 , n40577 );
    or g21859 ( n36159 , n11834 , n27884 );
    or g21860 ( n9254 , n38940 , n33671 );
    xnor g21861 ( n11115 , n21781 , n3834 );
    not g21862 ( n14004 , n29271 );
    xnor g21863 ( n17414 , n25552 , n10350 );
    or g21864 ( n6318 , n7435 , n14955 );
    and g21865 ( n16136 , n18745 , n22322 );
    xnor g21866 ( n18624 , n20204 , n10121 );
    not g21867 ( n33352 , n33392 );
    and g21868 ( n29840 , n6932 , n35099 );
    or g21869 ( n6137 , n39828 , n36328 );
    or g21870 ( n1014 , n14681 , n22282 );
    or g21871 ( n17127 , n39507 , n19890 );
    xnor g21872 ( n13732 , n40836 , n31796 );
    or g21873 ( n37054 , n27762 , n32224 );
    and g21874 ( n33972 , n38390 , n6868 );
    not g21875 ( n29739 , n32657 );
    not g21876 ( n42238 , n20924 );
    xnor g21877 ( n35699 , n31099 , n39621 );
    not g21878 ( n14676 , n37423 );
    nor g21879 ( n3957 , n8638 , n10224 );
    xnor g21880 ( n11668 , n41013 , n14491 );
    nor g21881 ( n40426 , n7356 , n14985 );
    or g21882 ( n3761 , n1115 , n4839 );
    not g21883 ( n40297 , n20360 );
    xnor g21884 ( n16701 , n6625 , n2330 );
    not g21885 ( n4843 , n9652 );
    or g21886 ( n5571 , n11771 , n3410 );
    or g21887 ( n4602 , n10027 , n5795 );
    or g21888 ( n2775 , n17221 , n36979 );
    and g21889 ( n21117 , n31813 , n23030 );
    or g21890 ( n33376 , n32848 , n36786 );
    and g21891 ( n8657 , n20009 , n35696 );
    not g21892 ( n42722 , n3003 );
    and g21893 ( n8697 , n36436 , n26864 );
    or g21894 ( n42049 , n2210 , n33465 );
    and g21895 ( n11655 , n15136 , n26814 );
    not g21896 ( n369 , n6196 );
    nor g21897 ( n18931 , n19418 , n16282 );
    not g21898 ( n2080 , n2818 );
    not g21899 ( n27344 , n8542 );
    or g21900 ( n25739 , n31376 , n39470 );
    nor g21901 ( n30763 , n41695 , n4887 );
    and g21902 ( n8710 , n12033 , n42599 );
    or g21903 ( n36388 , n42521 , n9614 );
    or g21904 ( n19239 , n29058 , n12931 );
    not g21905 ( n18597 , n37531 );
    or g21906 ( n38730 , n4531 , n2785 );
    or g21907 ( n1182 , n2407 , n2178 );
    xnor g21908 ( n41452 , n41358 , n9863 );
    or g21909 ( n301 , n36325 , n31156 );
    or g21910 ( n32916 , n15096 , n30892 );
    xnor g21911 ( n21105 , n34875 , n10521 );
    or g21912 ( n37453 , n5966 , n39905 );
    or g21913 ( n3667 , n16109 , n9424 );
    and g21914 ( n2148 , n18910 , n41374 );
    or g21915 ( n41144 , n17035 , n38017 );
    and g21916 ( n19892 , n21530 , n34449 );
    or g21917 ( n41256 , n5872 , n36342 );
    or g21918 ( n23851 , n14707 , n20629 );
    nor g21919 ( n16438 , n14316 , n28734 );
    and g21920 ( n41893 , n28101 , n36350 );
    and g21921 ( n22568 , n5723 , n40891 );
    and g21922 ( n7359 , n39352 , n18764 );
    or g21923 ( n19995 , n2820 , n36921 );
    xnor g21924 ( n21653 , n14649 , n796 );
    and g21925 ( n40277 , n28619 , n23338 );
    xnor g21926 ( n16266 , n1255 , n30871 );
    xnor g21927 ( n37931 , n34731 , n17078 );
    not g21928 ( n33633 , n25832 );
    xnor g21929 ( n20991 , n31989 , n33486 );
    or g21930 ( n6324 , n12633 , n19866 );
    nor g21931 ( n33475 , n25777 , n13514 );
    nor g21932 ( n40956 , n6547 , n3632 );
    and g21933 ( n35473 , n27888 , n36545 );
    xnor g21934 ( n3096 , n42356 , n3048 );
    or g21935 ( n1331 , n15163 , n40177 );
    not g21936 ( n16395 , n15396 );
    and g21937 ( n34074 , n33153 , n27004 );
    or g21938 ( n39666 , n2180 , n20446 );
    or g21939 ( n35744 , n30810 , n36288 );
    or g21940 ( n38540 , n33635 , n32744 );
    or g21941 ( n16834 , n20446 , n11577 );
    and g21942 ( n13991 , n4588 , n22653 );
    or g21943 ( n17588 , n5140 , n10561 );
    xnor g21944 ( n18084 , n38413 , n33183 );
    and g21945 ( n30635 , n39598 , n16710 );
    not g21946 ( n29740 , n36117 );
    or g21947 ( n25284 , n21678 , n12761 );
    not g21948 ( n9040 , n6032 );
    and g21949 ( n10699 , n38645 , n13839 );
    or g21950 ( n1842 , n3573 , n37454 );
    or g21951 ( n36616 , n23374 , n35437 );
    or g21952 ( n33067 , n31263 , n26573 );
    or g21953 ( n10387 , n6399 , n34170 );
    xnor g21954 ( n35607 , n8638 , n40347 );
    xnor g21955 ( n2250 , n33570 , n31339 );
    not g21956 ( n21159 , n37756 );
    or g21957 ( n17437 , n23405 , n20498 );
    not g21958 ( n26680 , n39139 );
    not g21959 ( n27537 , n20959 );
    xnor g21960 ( n36627 , n32297 , n1138 );
    or g21961 ( n42004 , n20296 , n32691 );
    or g21962 ( n15855 , n15242 , n20614 );
    and g21963 ( n17232 , n39695 , n18688 );
    xnor g21964 ( n12402 , n8724 , n35176 );
    not g21965 ( n19041 , n13105 );
    or g21966 ( n4835 , n7613 , n2525 );
    and g21967 ( n27616 , n28669 , n3107 );
    and g21968 ( n21671 , n10259 , n14717 );
    and g21969 ( n20565 , n15284 , n14889 );
    and g21970 ( n714 , n28490 , n39300 );
    and g21971 ( n22876 , n36860 , n30333 );
    and g21972 ( n41938 , n36088 , n14305 );
    and g21973 ( n10022 , n26990 , n29383 );
    or g21974 ( n37422 , n5317 , n23591 );
    not g21975 ( n14975 , n27063 );
    and g21976 ( n1651 , n11560 , n22951 );
    or g21977 ( n5269 , n41534 , n33604 );
    xnor g21978 ( n25796 , n42064 , n13277 );
    and g21979 ( n31266 , n8833 , n9516 );
    and g21980 ( n21820 , n19606 , n28302 );
    not g21981 ( n2862 , n38898 );
    and g21982 ( n4394 , n32682 , n29806 );
    or g21983 ( n15086 , n8220 , n36425 );
    or g21984 ( n42601 , n25627 , n32564 );
    or g21985 ( n31823 , n36892 , n36962 );
    not g21986 ( n21941 , n11879 );
    not g21987 ( n29897 , n11602 );
    not g21988 ( n42715 , n32573 );
    not g21989 ( n27835 , n25842 );
    not g21990 ( n39382 , n33960 );
    and g21991 ( n11381 , n33390 , n28181 );
    or g21992 ( n23609 , n29693 , n18236 );
    or g21993 ( n21167 , n42173 , n18473 );
    not g21994 ( n9165 , n8805 );
    not g21995 ( n37498 , n30520 );
    and g21996 ( n40456 , n8756 , n22916 );
    and g21997 ( n20201 , n26127 , n42090 );
    or g21998 ( n30217 , n19406 , n5821 );
    nor g21999 ( n37347 , n33981 , n25778 );
    nor g22000 ( n19073 , n14169 , n20667 );
    or g22001 ( n10038 , n8020 , n35057 );
    not g22002 ( n7580 , n28436 );
    or g22003 ( n4652 , n38075 , n35581 );
    nor g22004 ( n29540 , n1092 , n35145 );
    xnor g22005 ( n26864 , n35322 , n19888 );
    or g22006 ( n32966 , n20633 , n34215 );
    and g22007 ( n28235 , n3143 , n28266 );
    or g22008 ( n25622 , n31563 , n39408 );
    not g22009 ( n34744 , n38907 );
    or g22010 ( n11875 , n36403 , n40679 );
    or g22011 ( n8085 , n39556 , n25646 );
    xnor g22012 ( n40825 , n33517 , n1213 );
    nor g22013 ( n18089 , n35301 , n17500 );
    xnor g22014 ( n34493 , n9149 , n30026 );
    and g22015 ( n38140 , n33370 , n16312 );
    xnor g22016 ( n9179 , n2338 , n41833 );
    not g22017 ( n17220 , n7035 );
    xnor g22018 ( n42575 , n13194 , n1507 );
    or g22019 ( n23525 , n5239 , n34943 );
    and g22020 ( n33648 , n18594 , n4618 );
    nor g22021 ( n30843 , n25333 , n39323 );
    not g22022 ( n30280 , n14606 );
    nor g22023 ( n25771 , n34377 , n41018 );
    or g22024 ( n32571 , n28745 , n1424 );
    or g22025 ( n42709 , n8687 , n35719 );
    or g22026 ( n18900 , n6316 , n19962 );
    and g22027 ( n42530 , n6856 , n29724 );
    xnor g22028 ( n42151 , n26579 , n9047 );
    or g22029 ( n24211 , n696 , n13348 );
    not g22030 ( n17576 , n13430 );
    and g22031 ( n21143 , n23448 , n22001 );
    and g22032 ( n10785 , n33043 , n36575 );
    xnor g22033 ( n40653 , n12057 , n25970 );
    and g22034 ( n20734 , n4698 , n19686 );
    not g22035 ( n3530 , n34553 );
    nor g22036 ( n31932 , n13832 , n4336 );
    or g22037 ( n39032 , n6074 , n1044 );
    and g22038 ( n209 , n25822 , n537 );
    or g22039 ( n14725 , n20789 , n32857 );
    or g22040 ( n2014 , n20984 , n8469 );
    or g22041 ( n29324 , n9329 , n16324 );
    nor g22042 ( n18945 , n33647 , n3790 );
    and g22043 ( n30750 , n17177 , n39978 );
    xnor g22044 ( n36974 , n18490 , n35301 );
    and g22045 ( n6944 , n11998 , n12940 );
    or g22046 ( n26060 , n39195 , n4868 );
    or g22047 ( n28941 , n31354 , n468 );
    nor g22048 ( n32997 , n5964 , n22909 );
    nor g22049 ( n10499 , n30176 , n31866 );
    xnor g22050 ( n40813 , n6625 , n5455 );
    or g22051 ( n37279 , n15388 , n2817 );
    not g22052 ( n13630 , n428 );
    not g22053 ( n22070 , n8586 );
    nor g22054 ( n10679 , n6514 , n3063 );
    and g22055 ( n41100 , n38522 , n29532 );
    and g22056 ( n13837 , n32721 , n14323 );
    or g22057 ( n18266 , n8955 , n38395 );
    and g22058 ( n7789 , n5746 , n6607 );
    xnor g22059 ( n10758 , n14841 , n14352 );
    not g22060 ( n28239 , n32679 );
    nor g22061 ( n30748 , n41995 , n942 );
    or g22062 ( n1848 , n19883 , n25626 );
    or g22063 ( n31423 , n4156 , n9160 );
    or g22064 ( n40603 , n15418 , n3042 );
    or g22065 ( n11638 , n19414 , n13211 );
    or g22066 ( n4988 , n12867 , n18703 );
    or g22067 ( n31196 , n31693 , n7303 );
    not g22068 ( n27184 , n38661 );
    or g22069 ( n24397 , n39426 , n1319 );
    not g22070 ( n6572 , n12441 );
    not g22071 ( n8104 , n39124 );
    nor g22072 ( n12062 , n36112 , n36571 );
    or g22073 ( n9454 , n6754 , n30328 );
    xnor g22074 ( n21880 , n3549 , n33597 );
    and g22075 ( n16845 , n4382 , n39955 );
    nor g22076 ( n13498 , n15273 , n11893 );
    and g22077 ( n29288 , n25167 , n5054 );
    xnor g22078 ( n1814 , n16717 , n41071 );
    and g22079 ( n33497 , n484 , n36957 );
    and g22080 ( n20071 , n19677 , n32381 );
    and g22081 ( n25885 , n35493 , n35226 );
    and g22082 ( n6716 , n20326 , n31586 );
    nor g22083 ( n21662 , n1847 , n16318 );
    or g22084 ( n25667 , n576 , n34561 );
    and g22085 ( n4715 , n2411 , n9496 );
    or g22086 ( n27843 , n21469 , n30440 );
    and g22087 ( n41581 , n15562 , n6202 );
    or g22088 ( n17969 , n9456 , n21143 );
    and g22089 ( n36417 , n21450 , n39472 );
    or g22090 ( n20639 , n40289 , n11285 );
    and g22091 ( n2311 , n35628 , n40096 );
    xnor g22092 ( n2235 , n6760 , n14442 );
    not g22093 ( n6790 , n2562 );
    nor g22094 ( n30392 , n27142 , n39316 );
    xnor g22095 ( n41179 , n784 , n36130 );
    or g22096 ( n36666 , n32557 , n8679 );
    or g22097 ( n25977 , n39112 , n14930 );
    or g22098 ( n36714 , n20446 , n20035 );
    or g22099 ( n21637 , n11951 , n32767 );
    nor g22100 ( n1946 , n34071 , n5015 );
    nor g22101 ( n26442 , n33981 , n28721 );
    or g22102 ( n33687 , n18000 , n2750 );
    or g22103 ( n38047 , n39376 , n20225 );
    not g22104 ( n27258 , n32473 );
    or g22105 ( n27873 , n40485 , n10643 );
    and g22106 ( n26816 , n6510 , n10237 );
    or g22107 ( n23666 , n26935 , n27383 );
    nor g22108 ( n34520 , n18997 , n3046 );
    nor g22109 ( n5133 , n22452 , n29534 );
    nor g22110 ( n25808 , n35705 , n20496 );
    or g22111 ( n11591 , n4963 , n14441 );
    and g22112 ( n42568 , n6357 , n11217 );
    or g22113 ( n7344 , n17111 , n9879 );
    and g22114 ( n28690 , n31311 , n5237 );
    and g22115 ( n42122 , n17289 , n20986 );
    or g22116 ( n34883 , n42473 , n23682 );
    and g22117 ( n12176 , n1814 , n25429 );
    and g22118 ( n40114 , n3348 , n21030 );
    not g22119 ( n25849 , n26268 );
    and g22120 ( n38436 , n8119 , n6061 );
    nor g22121 ( n1665 , n1085 , n11458 );
    not g22122 ( n2223 , n15166 );
    not g22123 ( n23739 , n21561 );
    or g22124 ( n36406 , n26439 , n3932 );
    and g22125 ( n23466 , n21261 , n26603 );
    or g22126 ( n11373 , n18375 , n23569 );
    and g22127 ( n12457 , n18106 , n41709 );
    and g22128 ( n2837 , n14619 , n20472 );
    or g22129 ( n25240 , n14746 , n24708 );
    xnor g22130 ( n13283 , n21598 , n22884 );
    or g22131 ( n42276 , n11374 , n21098 );
    nor g22132 ( n31037 , n33796 , n41332 );
    or g22133 ( n12929 , n23880 , n21812 );
    xnor g22134 ( n32456 , n42732 , n38157 );
    nor g22135 ( n7560 , n9951 , n40760 );
    and g22136 ( n17302 , n12175 , n8061 );
    or g22137 ( n36859 , n5408 , n39317 );
    and g22138 ( n14054 , n9590 , n4596 );
    xnor g22139 ( n29893 , n1555 , n25937 );
    xnor g22140 ( n26709 , n36998 , n19325 );
    or g22141 ( n36558 , n33259 , n33859 );
    xnor g22142 ( n41410 , n7127 , n18973 );
    xnor g22143 ( n26361 , n18433 , n6194 );
    nor g22144 ( n29294 , n14052 , n23965 );
    or g22145 ( n18903 , n27913 , n29324 );
    not g22146 ( n34566 , n22777 );
    not g22147 ( n13151 , n31965 );
    or g22148 ( n17345 , n34594 , n1946 );
    and g22149 ( n30081 , n41172 , n31326 );
    and g22150 ( n26824 , n39535 , n23393 );
    xnor g22151 ( n28570 , n41480 , n26755 );
    and g22152 ( n8067 , n14751 , n41500 );
    and g22153 ( n16591 , n11099 , n16270 );
    not g22154 ( n34393 , n14473 );
    and g22155 ( n14110 , n23966 , n40869 );
    not g22156 ( n41943 , n5305 );
    or g22157 ( n13351 , n19215 , n25084 );
    nor g22158 ( n23044 , n476 , n33717 );
    or g22159 ( n2134 , n37264 , n42613 );
    and g22160 ( n34244 , n32422 , n16175 );
    and g22161 ( n39709 , n42606 , n8529 );
    nor g22162 ( n15239 , n39757 , n28701 );
    or g22163 ( n28963 , n2170 , n41684 );
    and g22164 ( n35833 , n13910 , n12518 );
    or g22165 ( n22657 , n21538 , n21172 );
    nor g22166 ( n567 , n34704 , n22297 );
    or g22167 ( n2934 , n35690 , n9599 );
    and g22168 ( n29292 , n12928 , n29537 );
    or g22169 ( n39381 , n10044 , n16756 );
    and g22170 ( n22203 , n24789 , n13376 );
    and g22171 ( n31100 , n42847 , n4201 );
    not g22172 ( n41831 , n18525 );
    not g22173 ( n37685 , n14962 );
    or g22174 ( n33059 , n14471 , n11727 );
    xnor g22175 ( n15793 , n21190 , n16056 );
    not g22176 ( n15166 , n40531 );
    and g22177 ( n15837 , n24859 , n1654 );
    or g22178 ( n22034 , n209 , n38820 );
    or g22179 ( n5382 , n34397 , n1429 );
    not g22180 ( n15476 , n32596 );
    or g22181 ( n41369 , n13248 , n21137 );
    or g22182 ( n16218 , n20116 , n556 );
    or g22183 ( n1541 , n35301 , n18827 );
    or g22184 ( n39909 , n8523 , n17492 );
    and g22185 ( n19349 , n2219 , n25848 );
    xnor g22186 ( n33852 , n19548 , n10239 );
    and g22187 ( n20514 , n13978 , n1146 );
    or g22188 ( n31390 , n20932 , n2245 );
    not g22189 ( n10697 , n12465 );
    or g22190 ( n17541 , n6893 , n30192 );
    or g22191 ( n19557 , n14434 , n5278 );
    not g22192 ( n5310 , n16845 );
    or g22193 ( n22030 , n32832 , n19242 );
    not g22194 ( n41956 , n26655 );
    nor g22195 ( n367 , n16418 , n39055 );
    or g22196 ( n29815 , n19815 , n11026 );
    and g22197 ( n42384 , n21718 , n26085 );
    nor g22198 ( n9926 , n29053 , n42855 );
    not g22199 ( n39930 , n31091 );
    or g22200 ( n7481 , n18023 , n23959 );
    and g22201 ( n29384 , n7399 , n8957 );
    nor g22202 ( n24787 , n4388 , n10751 );
    and g22203 ( n32975 , n39787 , n27600 );
    xnor g22204 ( n3494 , n5013 , n33983 );
    nor g22205 ( n33372 , n36823 , n29140 );
    or g22206 ( n8310 , n16925 , n38126 );
    and g22207 ( n37902 , n23853 , n40606 );
    and g22208 ( n36198 , n36118 , n40809 );
    and g22209 ( n31557 , n20088 , n5811 );
    nor g22210 ( n1692 , n41545 , n24784 );
    xnor g22211 ( n23357 , n34052 , n814 );
    not g22212 ( n31256 , n17441 );
    xnor g22213 ( n22412 , n29700 , n14471 );
    xnor g22214 ( n30766 , n1316 , n13730 );
    or g22215 ( n32778 , n25795 , n3066 );
    or g22216 ( n35201 , n27251 , n4287 );
    not g22217 ( n27296 , n4487 );
    xnor g22218 ( n34576 , n9597 , n29755 );
    and g22219 ( n41336 , n34492 , n27657 );
    xnor g22220 ( n39090 , n11383 , n15789 );
    nor g22221 ( n16330 , n17100 , n20942 );
    or g22222 ( n10101 , n34565 , n7118 );
    and g22223 ( n41289 , n33384 , n17746 );
    or g22224 ( n21642 , n15033 , n17104 );
    nor g22225 ( n30461 , n12148 , n12737 );
    or g22226 ( n9469 , n42263 , n10996 );
    not g22227 ( n35834 , n15708 );
    nor g22228 ( n13362 , n18487 , n30559 );
    or g22229 ( n3615 , n23509 , n18926 );
    and g22230 ( n34287 , n20576 , n41663 );
    and g22231 ( n32061 , n42210 , n38018 );
    xnor g22232 ( n42403 , n31099 , n10851 );
    or g22233 ( n1501 , n25882 , n35078 );
    or g22234 ( n3206 , n21199 , n22531 );
    xnor g22235 ( n23475 , n10411 , n24672 );
    and g22236 ( n28221 , n15881 , n3470 );
    or g22237 ( n20849 , n27960 , n38574 );
    not g22238 ( n15007 , n18919 );
    not g22239 ( n3035 , n27901 );
    and g22240 ( n1758 , n14006 , n17682 );
    or g22241 ( n39668 , n29382 , n3588 );
    not g22242 ( n11291 , n2596 );
    not g22243 ( n7130 , n16782 );
    xnor g22244 ( n29253 , n25619 , n42299 );
    not g22245 ( n41098 , n19607 );
    not g22246 ( n40421 , n32592 );
    or g22247 ( n41045 , n41861 , n21006 );
    or g22248 ( n7779 , n31319 , n31282 );
    or g22249 ( n33644 , n4842 , n38483 );
    and g22250 ( n39848 , n7606 , n35940 );
    nor g22251 ( n21036 , n5896 , n22020 );
    and g22252 ( n28796 , n12864 , n8263 );
    nor g22253 ( n26832 , n13650 , n11241 );
    nor g22254 ( n5402 , n4561 , n584 );
    or g22255 ( n24995 , n29276 , n40988 );
    or g22256 ( n11958 , n15095 , n2079 );
    nor g22257 ( n3676 , n36117 , n12435 );
    or g22258 ( n30124 , n38196 , n29788 );
    and g22259 ( n23548 , n5490 , n28844 );
    nor g22260 ( n7823 , n5964 , n19989 );
    and g22261 ( n819 , n37006 , n40835 );
    and g22262 ( n21357 , n11751 , n24880 );
    or g22263 ( n22747 , n38695 , n856 );
    or g22264 ( n23654 , n9789 , n16222 );
    or g22265 ( n41209 , n33683 , n6588 );
    or g22266 ( n30093 , n16658 , n38691 );
    and g22267 ( n10113 , n28105 , n5939 );
    or g22268 ( n34 , n35908 , n16655 );
    and g22269 ( n7213 , n15574 , n31207 );
    or g22270 ( n30327 , n7452 , n41862 );
    not g22271 ( n17851 , n38016 );
    or g22272 ( n40385 , n1110 , n8309 );
    nor g22273 ( n29427 , n40898 , n7634 );
    or g22274 ( n26814 , n38849 , n7149 );
    xnor g22275 ( n14234 , n40012 , n7240 );
    or g22276 ( n32837 , n24713 , n25580 );
    and g22277 ( n33728 , n7238 , n42322 );
    and g22278 ( n17164 , n35211 , n19466 );
    nor g22279 ( n13334 , n38269 , n17985 );
    or g22280 ( n15562 , n38704 , n15683 );
    xnor g22281 ( n4330 , n12057 , n5631 );
    or g22282 ( n31060 , n40612 , n36247 );
    nor g22283 ( n1742 , n38922 , n19064 );
    and g22284 ( n25376 , n40500 , n14294 );
    nor g22285 ( n5493 , n8494 , n27878 );
    or g22286 ( n12810 , n11414 , n8117 );
    not g22287 ( n12456 , n25994 );
    or g22288 ( n3928 , n13413 , n35997 );
    and g22289 ( n35928 , n16022 , n12097 );
    and g22290 ( n25021 , n30121 , n5547 );
    not g22291 ( n31067 , n24610 );
    or g22292 ( n24137 , n27961 , n42479 );
    xnor g22293 ( n18211 , n39705 , n34985 );
    xnor g22294 ( n15587 , n31989 , n19664 );
    not g22295 ( n9911 , n23075 );
    and g22296 ( n27319 , n16977 , n29721 );
    and g22297 ( n42269 , n20117 , n37254 );
    nor g22298 ( n30593 , n1971 , n20706 );
    and g22299 ( n22491 , n6833 , n10195 );
    or g22300 ( n12797 , n26196 , n1589 );
    not g22301 ( n3277 , n27419 );
    xnor g22302 ( n9083 , n16998 , n24955 );
    or g22303 ( n25218 , n35216 , n28505 );
    xnor g22304 ( n19456 , n25744 , n18720 );
    or g22305 ( n13425 , n28080 , n5772 );
    nor g22306 ( n37018 , n38879 , n25762 );
    and g22307 ( n25846 , n9686 , n23038 );
    or g22308 ( n17886 , n24910 , n15780 );
    xnor g22309 ( n15815 , n30103 , n18517 );
    not g22310 ( n21558 , n23326 );
    or g22311 ( n19757 , n16936 , n19587 );
    and g22312 ( n11949 , n39600 , n32653 );
    or g22313 ( n33953 , n36534 , n5094 );
    or g22314 ( n24117 , n41641 , n13764 );
    or g22315 ( n36744 , n42646 , n36966 );
    xnor g22316 ( n9463 , n30139 , n33666 );
    nor g22317 ( n18060 , n37792 , n30961 );
    or g22318 ( n41502 , n17695 , n5261 );
    xnor g22319 ( n11561 , n6688 , n6898 );
    and g22320 ( n1840 , n37054 , n21974 );
    not g22321 ( n6914 , n40499 );
    nor g22322 ( n36720 , n10580 , n21105 );
    or g22323 ( n15503 , n25382 , n4255 );
    not g22324 ( n20331 , n34151 );
    or g22325 ( n41481 , n21265 , n36619 );
    or g22326 ( n2422 , n19206 , n36334 );
    and g22327 ( n40077 , n17604 , n22347 );
    and g22328 ( n8441 , n31384 , n23180 );
    and g22329 ( n20767 , n19454 , n14357 );
    and g22330 ( n12291 , n22279 , n11716 );
    and g22331 ( n37517 , n27975 , n2462 );
    not g22332 ( n5229 , n38195 );
    or g22333 ( n29960 , n20415 , n15006 );
    and g22334 ( n38127 , n28716 , n16296 );
    and g22335 ( n38276 , n25019 , n37184 );
    or g22336 ( n18878 , n37418 , n34793 );
    and g22337 ( n9269 , n41658 , n13045 );
    or g22338 ( n5152 , n30685 , n29522 );
    or g22339 ( n28620 , n41180 , n3829 );
    and g22340 ( n25651 , n23362 , n9973 );
    or g22341 ( n4313 , n10523 , n12159 );
    nor g22342 ( n17630 , n27245 , n12436 );
    or g22343 ( n32171 , n18051 , n646 );
    and g22344 ( n10511 , n6952 , n40402 );
    not g22345 ( n27250 , n25370 );
    or g22346 ( n19078 , n3431 , n16949 );
    or g22347 ( n2133 , n30847 , n19930 );
    not g22348 ( n30435 , n15439 );
    or g22349 ( n8221 , n8539 , n9410 );
    or g22350 ( n20588 , n13495 , n34807 );
    and g22351 ( n16501 , n35381 , n8822 );
    nor g22352 ( n600 , n26875 , n35021 );
    not g22353 ( n15589 , n23595 );
    nor g22354 ( n15606 , n16517 , n13842 );
    and g22355 ( n33995 , n32442 , n42619 );
    or g22356 ( n35985 , n31153 , n18571 );
    and g22357 ( n5243 , n32305 , n41407 );
    or g22358 ( n25186 , n25401 , n40787 );
    or g22359 ( n12833 , n18292 , n27179 );
    and g22360 ( n41071 , n9173 , n25638 );
    not g22361 ( n35633 , n13886 );
    or g22362 ( n16044 , n13795 , n34904 );
    not g22363 ( n27430 , n19125 );
    or g22364 ( n36781 , n34292 , n24259 );
    or g22365 ( n10408 , n25494 , n19965 );
    not g22366 ( n21981 , n6412 );
    not g22367 ( n40132 , n33277 );
    nor g22368 ( n24823 , n5964 , n14848 );
    xnor g22369 ( n18604 , n6053 , n18866 );
    or g22370 ( n37989 , n17903 , n34023 );
    or g22371 ( n30675 , n18884 , n23800 );
    or g22372 ( n26893 , n20199 , n40365 );
    xnor g22373 ( n40510 , n27900 , n29000 );
    or g22374 ( n39147 , n562 , n42614 );
    or g22375 ( n12 , n14471 , n11255 );
    and g22376 ( n24203 , n38908 , n2240 );
    not g22377 ( n14485 , n27452 );
    xnor g22378 ( n5018 , n38957 , n24910 );
    or g22379 ( n29196 , n21067 , n28195 );
    nor g22380 ( n16032 , n14876 , n20284 );
    or g22381 ( n15971 , n28527 , n256 );
    or g22382 ( n34660 , n34741 , n17942 );
    and g22383 ( n36640 , n38620 , n17825 );
    and g22384 ( n22752 , n29006 , n8875 );
    nor g22385 ( n30171 , n2372 , n259 );
    nor g22386 ( n29989 , n19689 , n3159 );
    or g22387 ( n35872 , n37699 , n31728 );
    not g22388 ( n27115 , n42738 );
    xnor g22389 ( n18286 , n25299 , n27859 );
    and g22390 ( n39294 , n38775 , n22826 );
    and g22391 ( n1990 , n16719 , n16298 );
    xnor g22392 ( n27022 , n4731 , n23086 );
    not g22393 ( n16628 , n9830 );
    and g22394 ( n38437 , n29698 , n20702 );
    or g22395 ( n21614 , n30036 , n36063 );
    and g22396 ( n20848 , n7295 , n10811 );
    or g22397 ( n33991 , n150 , n31571 );
    and g22398 ( n41425 , n29029 , n17027 );
    nor g22399 ( n21045 , n9370 , n2380 );
    or g22400 ( n26150 , n34555 , n11798 );
    or g22401 ( n41324 , n25304 , n31321 );
    or g22402 ( n42737 , n7943 , n5824 );
    nor g22403 ( n8981 , n996 , n21173 );
    or g22404 ( n6233 , n23087 , n31671 );
    or g22405 ( n39086 , n30228 , n32566 );
    nor g22406 ( n3798 , n4548 , n9252 );
    not g22407 ( n29616 , n7890 );
    or g22408 ( n2510 , n14886 , n30435 );
    or g22409 ( n24345 , n24915 , n31475 );
    or g22410 ( n26778 , n9748 , n27998 );
    nor g22411 ( n42783 , n3662 , n20938 );
    xnor g22412 ( n3773 , n36165 , n5104 );
    and g22413 ( n5688 , n8786 , n15511 );
    and g22414 ( n7215 , n20355 , n32365 );
    nor g22415 ( n10999 , n17823 , n36322 );
    or g22416 ( n9546 , n36196 , n28474 );
    not g22417 ( n10307 , n40600 );
    or g22418 ( n42376 , n38268 , n8676 );
    or g22419 ( n151 , n25600 , n19973 );
    xnor g22420 ( n39900 , n35727 , n15719 );
    not g22421 ( n23236 , n38364 );
    and g22422 ( n21906 , n37884 , n2872 );
    or g22423 ( n12774 , n27315 , n2310 );
    and g22424 ( n16761 , n5263 , n5240 );
    and g22425 ( n35998 , n24721 , n32148 );
    or g22426 ( n4348 , n21205 , n19084 );
    or g22427 ( n18005 , n39881 , n38211 );
    not g22428 ( n17288 , n11301 );
    and g22429 ( n30169 , n28886 , n39255 );
    and g22430 ( n583 , n12387 , n3253 );
    or g22431 ( n37554 , n28213 , n25590 );
    nor g22432 ( n5681 , n32394 , n23898 );
    not g22433 ( n24359 , n19608 );
    and g22434 ( n7026 , n2684 , n25324 );
    or g22435 ( n14178 , n19249 , n24785 );
    not g22436 ( n16150 , n37919 );
    and g22437 ( n13157 , n13537 , n34639 );
    or g22438 ( n39044 , n9036 , n22545 );
    or g22439 ( n21961 , n5283 , n42648 );
    or g22440 ( n39685 , n34160 , n6316 );
    and g22441 ( n17022 , n41264 , n23978 );
    or g22442 ( n10802 , n21096 , n26427 );
    and g22443 ( n26265 , n16739 , n26519 );
    or g22444 ( n6055 , n24528 , n34609 );
    or g22445 ( n22399 , n27680 , n21154 );
    xnor g22446 ( n28591 , n105 , n13396 );
    xnor g22447 ( n27030 , n40 , n4563 );
    not g22448 ( n14226 , n25607 );
    or g22449 ( n32868 , n6209 , n9665 );
    and g22450 ( n17729 , n7461 , n3733 );
    or g22451 ( n19506 , n16556 , n41993 );
    or g22452 ( n35591 , n40661 , n2395 );
    not g22453 ( n13606 , n18786 );
    or g22454 ( n38337 , n23173 , n11888 );
    or g22455 ( n39145 , n11653 , n26273 );
    not g22456 ( n10024 , n36939 );
    or g22457 ( n25892 , n40216 , n30850 );
    not g22458 ( n40462 , n22310 );
    or g22459 ( n19314 , n5910 , n17934 );
    and g22460 ( n29531 , n40573 , n16193 );
    and g22461 ( n2677 , n12705 , n12891 );
    xnor g22462 ( n39214 , n22799 , n375 );
    nor g22463 ( n39603 , n35301 , n36096 );
    nor g22464 ( n3828 , n42903 , n9026 );
    not g22465 ( n17111 , n26608 );
    and g22466 ( n39932 , n29375 , n18781 );
    xnor g22467 ( n34721 , n11436 , n29564 );
    and g22468 ( n3588 , n21322 , n23484 );
    nor g22469 ( n3353 , n19219 , n4471 );
    or g22470 ( n15454 , n677 , n4016 );
    nor g22471 ( n18265 , n37146 , n37232 );
    or g22472 ( n12263 , n14471 , n38840 );
    nor g22473 ( n37084 , n31811 , n31767 );
    nor g22474 ( n35141 , n19052 , n35214 );
    or g22475 ( n40013 , n19177 , n8717 );
    not g22476 ( n36408 , n9161 );
    and g22477 ( n12923 , n3852 , n41881 );
    xnor g22478 ( n13650 , n38867 , n39243 );
    not g22479 ( n6130 , n6870 );
    or g22480 ( n21431 , n36868 , n6111 );
    nor g22481 ( n36193 , n5896 , n31109 );
    or g22482 ( n27075 , n28290 , n22478 );
    or g22483 ( n29679 , n41961 , n20816 );
    and g22484 ( n23102 , n21713 , n21485 );
    not g22485 ( n40467 , n31916 );
    or g22486 ( n10983 , n28314 , n14295 );
    or g22487 ( n14496 , n11892 , n17026 );
    nor g22488 ( n31913 , n2435 , n36001 );
    xnor g22489 ( n29821 , n16693 , n25798 );
    or g22490 ( n28108 , n9485 , n30616 );
    and g22491 ( n410 , n3887 , n23501 );
    or g22492 ( n17300 , n16598 , n26573 );
    not g22493 ( n24289 , n37666 );
    and g22494 ( n15795 , n9542 , n37962 );
    or g22495 ( n30698 , n24194 , n35216 );
    not g22496 ( n2179 , n19322 );
    or g22497 ( n7107 , n22137 , n15164 );
    or g22498 ( n3755 , n17120 , n42302 );
    or g22499 ( n11249 , n22564 , n6842 );
    or g22500 ( n14357 , n15064 , n19465 );
    and g22501 ( n11128 , n26341 , n35527 );
    xnor g22502 ( n8859 , n36096 , n35301 );
    nor g22503 ( n7947 , n40752 , n9855 );
    or g22504 ( n16496 , n29661 , n3410 );
    and g22505 ( n20644 , n33342 , n12134 );
    not g22506 ( n2084 , n26501 );
    nor g22507 ( n32842 , n9030 , n30908 );
    xnor g22508 ( n5369 , n1297 , n6680 );
    not g22509 ( n42338 , n11830 );
    or g22510 ( n35451 , n32277 , n42763 );
    not g22511 ( n24442 , n30684 );
    nor g22512 ( n344 , n14707 , n38940 );
    or g22513 ( n34899 , n14599 , n26911 );
    nor g22514 ( n31387 , n4927 , n35485 );
    or g22515 ( n5503 , n10967 , n813 );
    or g22516 ( n26644 , n38494 , n39023 );
    or g22517 ( n28622 , n29343 , n37263 );
    nor g22518 ( n33874 , n10910 , n28183 );
    and g22519 ( n42372 , n26725 , n39484 );
    and g22520 ( n30163 , n27982 , n7448 );
    or g22521 ( n11011 , n42072 , n26230 );
    or g22522 ( n7062 , n22183 , n35405 );
    xnor g22523 ( n6261 , n21559 , n27355 );
    not g22524 ( n3813 , n7300 );
    or g22525 ( n3988 , n11935 , n30652 );
    or g22526 ( n15052 , n41839 , n6842 );
    or g22527 ( n17524 , n12351 , n36166 );
    and g22528 ( n18469 , n37436 , n37581 );
    not g22529 ( n8510 , n42881 );
    and g22530 ( n22014 , n18135 , n19139 );
    xnor g22531 ( n41611 , n4680 , n34565 );
    or g22532 ( n31984 , n1702 , n20239 );
    not g22533 ( n5728 , n37961 );
    nor g22534 ( n765 , n966 , n23409 );
    and g22535 ( n30328 , n27322 , n7366 );
    or g22536 ( n40929 , n13706 , n35626 );
    and g22537 ( n2795 , n37249 , n12491 );
    not g22538 ( n33130 , n19248 );
    or g22539 ( n34027 , n15349 , n33859 );
    and g22540 ( n25390 , n6996 , n10947 );
    not g22541 ( n8745 , n32403 );
    or g22542 ( n32914 , n28634 , n32183 );
    or g22543 ( n22656 , n34605 , n12669 );
    or g22544 ( n19111 , n2677 , n27039 );
    or g22545 ( n7249 , n42490 , n13477 );
    or g22546 ( n38351 , n4371 , n28392 );
    or g22547 ( n19042 , n20602 , n28379 );
    or g22548 ( n580 , n1765 , n16008 );
    not g22549 ( n33675 , n9726 );
    and g22550 ( n37503 , n7262 , n15502 );
    or g22551 ( n13159 , n4696 , n10214 );
    not g22552 ( n40557 , n41479 );
    or g22553 ( n8760 , n30443 , n5705 );
    and g22554 ( n40218 , n15298 , n33146 );
    or g22555 ( n28062 , n981 , n18063 );
    and g22556 ( n18014 , n12440 , n19147 );
    or g22557 ( n14896 , n7776 , n1149 );
    or g22558 ( n28250 , n3954 , n28931 );
    and g22559 ( n3256 , n27003 , n17933 );
    or g22560 ( n10640 , n17780 , n13291 );
    xnor g22561 ( n35523 , n1623 , n7120 );
    and g22562 ( n14278 , n35508 , n23482 );
    or g22563 ( n19569 , n39494 , n24674 );
    or g22564 ( n36045 , n4478 , n34561 );
    nor g22565 ( n37646 , n39599 , n24069 );
    or g22566 ( n3211 , n38240 , n10859 );
    not g22567 ( n11957 , n11010 );
    not g22568 ( n18548 , n21482 );
    xnor g22569 ( n18876 , n40 , n31552 );
    and g22570 ( n1141 , n14565 , n9850 );
    or g22571 ( n41167 , n10846 , n1387 );
    nor g22572 ( n36108 , n41293 , n12592 );
    not g22573 ( n39541 , n25618 );
    and g22574 ( n42674 , n3166 , n30027 );
    nor g22575 ( n2577 , n5959 , n11190 );
    or g22576 ( n15416 , n2972 , n27538 );
    not g22577 ( n37893 , n4571 );
    xnor g22578 ( n26421 , n24410 , n36624 );
    or g22579 ( n36310 , n22429 , n29562 );
    and g22580 ( n16388 , n21169 , n23024 );
    or g22581 ( n273 , n18392 , n32396 );
    and g22582 ( n23835 , n14896 , n7043 );
    or g22583 ( n2100 , n33594 , n9911 );
    not g22584 ( n4316 , n9078 );
    or g22585 ( n27042 , n11034 , n17383 );
    or g22586 ( n12603 , n37952 , n25737 );
    xnor g22587 ( n32378 , n20331 , n24440 );
    not g22588 ( n40285 , n38737 );
    and g22589 ( n33132 , n29154 , n39496 );
    nor g22590 ( n35558 , n37747 , n35765 );
    or g22591 ( n26589 , n37405 , n1194 );
    not g22592 ( n35456 , n2422 );
    or g22593 ( n20217 , n42462 , n5422 );
    or g22594 ( n36026 , n39541 , n19744 );
    or g22595 ( n288 , n11747 , n41191 );
    xnor g22596 ( n8708 , n10588 , n40737 );
    nor g22597 ( n18694 , n945 , n42401 );
    or g22598 ( n15122 , n4650 , n27712 );
    nor g22599 ( n42747 , n12775 , n21490 );
    or g22600 ( n24981 , n9269 , n3890 );
    or g22601 ( n36611 , n30977 , n4029 );
    or g22602 ( n19722 , n25012 , n26214 );
    nor g22603 ( n14987 , n19431 , n21597 );
    xnor g22604 ( n20593 , n22263 , n39731 );
    nor g22605 ( n31198 , n7200 , n40040 );
    or g22606 ( n37019 , n9197 , n16401 );
    or g22607 ( n1475 , n14365 , n12731 );
    or g22608 ( n27381 , n12171 , n4669 );
    or g22609 ( n21735 , n40807 , n1410 );
    or g22610 ( n29078 , n29579 , n41714 );
    not g22611 ( n42471 , n26920 );
    and g22612 ( n38653 , n20852 , n21368 );
    xnor g22613 ( n7479 , n25766 , n22311 );
    not g22614 ( n32586 , n34593 );
    not g22615 ( n23325 , n39082 );
    or g22616 ( n15919 , n42361 , n25087 );
    not g22617 ( n28993 , n14895 );
    or g22618 ( n30353 , n25699 , n5848 );
    and g22619 ( n37168 , n23866 , n32746 );
    or g22620 ( n5530 , n5558 , n24500 );
    nor g22621 ( n25430 , n8510 , n6421 );
    and g22622 ( n6693 , n13738 , n26257 );
    or g22623 ( n22923 , n17477 , n1367 );
    or g22624 ( n13544 , n14248 , n5261 );
    or g22625 ( n12679 , n14481 , n13320 );
    nor g22626 ( n14927 , n1494 , n10174 );
    or g22627 ( n22280 , n14245 , n35713 );
    not g22628 ( n31944 , n1230 );
    nor g22629 ( n38585 , n29973 , n17394 );
    and g22630 ( n4403 , n10545 , n15052 );
    not g22631 ( n21667 , n30217 );
    xnor g22632 ( n67 , n30818 , n3622 );
    or g22633 ( n31200 , n24350 , n41413 );
    not g22634 ( n11728 , n29730 );
    and g22635 ( n36534 , n28852 , n26220 );
    or g22636 ( n8668 , n28934 , n7210 );
    xnor g22637 ( n4065 , n25060 , n12677 );
    and g22638 ( n29585 , n13596 , n28151 );
    xnor g22639 ( n8733 , n30103 , n29982 );
    and g22640 ( n34942 , n12881 , n28236 );
    not g22641 ( n1977 , n18807 );
    and g22642 ( n5631 , n16875 , n17864 );
    and g22643 ( n41252 , n10421 , n12973 );
    not g22644 ( n13074 , n9182 );
    nor g22645 ( n8037 , n17120 , n19971 );
    or g22646 ( n35946 , n12606 , n6648 );
    or g22647 ( n6936 , n17193 , n23079 );
    not g22648 ( n14900 , n11085 );
    or g22649 ( n39107 , n41502 , n33033 );
    xnor g22650 ( n1487 , n6625 , n40669 );
    or g22651 ( n24742 , n42108 , n4617 );
    nor g22652 ( n20430 , n30295 , n3356 );
    or g22653 ( n26835 , n13380 , n8964 );
    or g22654 ( n2741 , n34565 , n9767 );
    not g22655 ( n34561 , n9588 );
    or g22656 ( n6749 , n26927 , n11236 );
    not g22657 ( n14506 , n36154 );
    nor g22658 ( n9787 , n24705 , n22136 );
    xnor g22659 ( n30943 , n31099 , n18181 );
    xnor g22660 ( n32804 , n21826 , n5343 );
    or g22661 ( n33757 , n30914 , n33625 );
    and g22662 ( n4964 , n38868 , n31712 );
    nor g22663 ( n16045 , n8494 , n35662 );
    not g22664 ( n12780 , n29345 );
    xnor g22665 ( n19857 , n21365 , n10386 );
    nor g22666 ( n42346 , n3344 , n26066 );
    nor g22667 ( n20210 , n7076 , n19192 );
    xnor g22668 ( n29978 , n28201 , n23464 );
    xnor g22669 ( n14554 , n36009 , n4403 );
    not g22670 ( n5407 , n28354 );
    or g22671 ( n34620 , n23028 , n6275 );
    or g22672 ( n17323 , n3034 , n17498 );
    and g22673 ( n16748 , n8743 , n18922 );
    or g22674 ( n1957 , n29857 , n31254 );
    or g22675 ( n26725 , n17120 , n2016 );
    not g22676 ( n30188 , n18887 );
    nor g22677 ( n20686 , n2134 , n21412 );
    nor g22678 ( n17322 , n14440 , n41230 );
    or g22679 ( n6491 , n28576 , n17522 );
    xnor g22680 ( n30854 , n32590 , n40842 );
    or g22681 ( n23979 , n34391 , n42823 );
    or g22682 ( n10424 , n5895 , n28457 );
    not g22683 ( n12172 , n34646 );
    or g22684 ( n28742 , n15429 , n10626 );
    or g22685 ( n28077 , n7141 , n33238 );
    and g22686 ( n11314 , n11010 , n13652 );
    xnor g22687 ( n5064 , n19385 , n12839 );
    or g22688 ( n37327 , n22776 , n20296 );
    nor g22689 ( n13028 , n35472 , n24669 );
    not g22690 ( n31175 , n28977 );
    or g22691 ( n2109 , n33262 , n22024 );
    or g22692 ( n8686 , n24379 , n42544 );
    xnor g22693 ( n12033 , n7943 , n3587 );
    or g22694 ( n25307 , n15911 , n22259 );
    or g22695 ( n8258 , n32344 , n25719 );
    or g22696 ( n253 , n13513 , n21772 );
    or g22697 ( n21052 , n3765 , n33131 );
    and g22698 ( n7144 , n37604 , n24589 );
    or g22699 ( n16399 , n900 , n33132 );
    and g22700 ( n28932 , n10812 , n29401 );
    and g22701 ( n39940 , n6766 , n35252 );
    and g22702 ( n42874 , n28467 , n14136 );
    and g22703 ( n17959 , n27041 , n23408 );
    or g22704 ( n1744 , n1724 , n2622 );
    xnor g22705 ( n3972 , n8416 , n15636 );
    or g22706 ( n40800 , n31471 , n5911 );
    or g22707 ( n31330 , n23724 , n42378 );
    nor g22708 ( n11864 , n4275 , n11285 );
    or g22709 ( n37966 , n30854 , n328 );
    and g22710 ( n14204 , n41242 , n33280 );
    and g22711 ( n40412 , n38725 , n13804 );
    xnor g22712 ( n38702 , n25822 , n537 );
    or g22713 ( n40522 , n1971 , n38354 );
    not g22714 ( n30606 , n32447 );
    not g22715 ( n41870 , n18829 );
    or g22716 ( n31324 , n3583 , n18631 );
    nor g22717 ( n8105 , n11986 , n20855 );
    or g22718 ( n11015 , n12809 , n21632 );
    xnor g22719 ( n3045 , n26279 , n11805 );
    xnor g22720 ( n1709 , n20160 , n3364 );
    not g22721 ( n24307 , n41758 );
    or g22722 ( n9736 , n34182 , n31100 );
    or g22723 ( n30580 , n10284 , n25470 );
    or g22724 ( n10076 , n7441 , n31192 );
    nor g22725 ( n7645 , n4896 , n11093 );
    and g22726 ( n41594 , n16337 , n27451 );
    or g22727 ( n21236 , n26995 , n28019 );
    or g22728 ( n1193 , n32051 , n7265 );
    or g22729 ( n6941 , n6327 , n24702 );
    and g22730 ( n30129 , n39406 , n30816 );
    nor g22731 ( n9687 , n21649 , n20665 );
    or g22732 ( n24495 , n10496 , n37471 );
    xnor g22733 ( n6059 , n40 , n21098 );
    and g22734 ( n30302 , n36998 , n33376 );
    not g22735 ( n22722 , n33852 );
    and g22736 ( n5313 , n13153 , n1343 );
    and g22737 ( n14608 , n15876 , n9517 );
    and g22738 ( n4368 , n21800 , n12102 );
    not g22739 ( n17935 , n15439 );
    not g22740 ( n41153 , n26846 );
    xnor g22741 ( n14246 , n34731 , n20650 );
    or g22742 ( n20540 , n26838 , n35713 );
    not g22743 ( n29473 , n1132 );
    or g22744 ( n41446 , n35534 , n23871 );
    xnor g22745 ( n17433 , n36452 , n40058 );
    not g22746 ( n29347 , n19407 );
    not g22747 ( n29987 , n14206 );
    nor g22748 ( n34596 , n5926 , n32407 );
    xnor g22749 ( n27423 , n21457 , n42411 );
    or g22750 ( n8834 , n23196 , n7942 );
    and g22751 ( n10215 , n40917 , n41977 );
    xnor g22752 ( n6443 , n28319 , n34605 );
    xnor g22753 ( n29592 , n13444 , n16550 );
    and g22754 ( n15461 , n35568 , n11329 );
    and g22755 ( n13603 , n24735 , n25441 );
    xnor g22756 ( n5955 , n12605 , n31513 );
    nor g22757 ( n25951 , n39449 , n40157 );
    xnor g22758 ( n20858 , n27734 , n6078 );
    nor g22759 ( n2696 , n34376 , n6737 );
    and g22760 ( n6719 , n10519 , n15141 );
    and g22761 ( n2496 , n25050 , n22481 );
    xnor g22762 ( n17854 , n7943 , n35489 );
    not g22763 ( n4282 , n20949 );
    not g22764 ( n41206 , n24221 );
    or g22765 ( n32664 , n27311 , n40714 );
    or g22766 ( n13734 , n5391 , n17104 );
    or g22767 ( n34149 , n15095 , n38732 );
    or g22768 ( n25512 , n21697 , n40154 );
    or g22769 ( n30106 , n18236 , n35577 );
    and g22770 ( n30168 , n18555 , n30459 );
    and g22771 ( n25174 , n21188 , n40822 );
    and g22772 ( n21044 , n41704 , n2590 );
    or g22773 ( n9274 , n4087 , n37806 );
    or g22774 ( n11159 , n42712 , n19009 );
    or g22775 ( n36710 , n10625 , n20616 );
    and g22776 ( n21933 , n20400 , n4577 );
    and g22777 ( n42253 , n36090 , n25434 );
    or g22778 ( n42724 , n36815 , n1279 );
    not g22779 ( n26056 , n8573 );
    and g22780 ( n19676 , n7543 , n25612 );
    nor g22781 ( n21011 , n38879 , n15688 );
    or g22782 ( n24735 , n25241 , n15402 );
    not g22783 ( n526 , n8897 );
    not g22784 ( n5685 , n10282 );
    xnor g22785 ( n17708 , n35727 , n24260 );
    or g22786 ( n2110 , n4099 , n41384 );
    not g22787 ( n16052 , n9005 );
    or g22788 ( n19914 , n30894 , n271 );
    or g22789 ( n5127 , n1839 , n6583 );
    and g22790 ( n29254 , n9324 , n6659 );
    or g22791 ( n1839 , n17907 , n20900 );
    xnor g22792 ( n42884 , n105 , n42504 );
    not g22793 ( n9597 , n32824 );
    nor g22794 ( n8068 , n42042 , n6118 );
    not g22795 ( n4401 , n41952 );
    and g22796 ( n24508 , n264 , n7894 );
    or g22797 ( n11171 , n1774 , n20288 );
    nor g22798 ( n25535 , n14614 , n24611 );
    and g22799 ( n6703 , n1627 , n26656 );
    or g22800 ( n34193 , n26764 , n905 );
    or g22801 ( n34970 , n9748 , n2777 );
    xnor g22802 ( n31721 , n36273 , n37190 );
    or g22803 ( n25162 , n4689 , n30670 );
    and g22804 ( n11838 , n13290 , n21358 );
    not g22805 ( n35216 , n40635 );
    not g22806 ( n40259 , n22953 );
    not g22807 ( n6260 , n35766 );
    nor g22808 ( n32815 , n38261 , n18482 );
    or g22809 ( n26622 , n38494 , n35473 );
    and g22810 ( n35685 , n13716 , n13090 );
    not g22811 ( n42627 , n28718 );
    xnor g22812 ( n6951 , n40 , n13744 );
    xnor g22813 ( n21051 , n36046 , n23253 );
    or g22814 ( n15079 , n41635 , n4552 );
    nor g22815 ( n4742 , n40617 , n4815 );
    xnor g22816 ( n8449 , n718 , n16816 );
    and g22817 ( n28863 , n18210 , n28102 );
    nor g22818 ( n34345 , n5896 , n12937 );
    or g22819 ( n3114 , n15003 , n8375 );
    not g22820 ( n21745 , n18950 );
    or g22821 ( n103 , n32752 , n21112 );
    or g22822 ( n21549 , n21021 , n36893 );
    and g22823 ( n41809 , n2772 , n25128 );
    or g22824 ( n36715 , n34828 , n34796 );
    and g22825 ( n15596 , n11870 , n40968 );
    or g22826 ( n23178 , n11337 , n15095 );
    and g22827 ( n28213 , n26848 , n37475 );
    or g22828 ( n13943 , n39118 , n24450 );
    or g22829 ( n6085 , n40455 , n20751 );
    not g22830 ( n23541 , n15004 );
    or g22831 ( n1363 , n9264 , n2563 );
    or g22832 ( n37933 , n27471 , n39408 );
    and g22833 ( n21388 , n7761 , n30439 );
    not g22834 ( n39018 , n3793 );
    xnor g22835 ( n23022 , n10705 , n6506 );
    nor g22836 ( n10560 , n31674 , n5357 );
    or g22837 ( n42241 , n27426 , n439 );
    not g22838 ( n34927 , n18907 );
    or g22839 ( n12032 , n22158 , n6284 );
    or g22840 ( n26668 , n2492 , n10976 );
    and g22841 ( n15618 , n32931 , n7122 );
    and g22842 ( n1633 , n28288 , n29945 );
    or g22843 ( n16512 , n24637 , n24254 );
    xnor g22844 ( n28800 , n31107 , n6937 );
    not g22845 ( n977 , n5584 );
    and g22846 ( n40882 , n34926 , n14011 );
    nor g22847 ( n9358 , n33981 , n161 );
    or g22848 ( n36763 , n39247 , n29541 );
    nor g22849 ( n20741 , n19221 , n31307 );
    or g22850 ( n34047 , n1735 , n31911 );
    or g22851 ( n32486 , n37520 , n38676 );
    or g22852 ( n11041 , n36280 , n10351 );
    or g22853 ( n37420 , n6943 , n40074 );
    or g22854 ( n16652 , n5695 , n35745 );
    not g22855 ( n20039 , n40912 );
    and g22856 ( n20366 , n20624 , n13538 );
    and g22857 ( n14317 , n7757 , n25758 );
    or g22858 ( n22055 , n23082 , n18893 );
    not g22859 ( n27371 , n4109 );
    not g22860 ( n35074 , n10072 );
    nor g22861 ( n37147 , n15800 , n27269 );
    or g22862 ( n22522 , n27487 , n37339 );
    or g22863 ( n5047 , n40978 , n3727 );
    and g22864 ( n6188 , n24519 , n20318 );
    xnor g22865 ( n23907 , n28288 , n29945 );
    or g22866 ( n3112 , n6370 , n12568 );
    or g22867 ( n16542 , n26504 , n6960 );
    and g22868 ( n27938 , n2099 , n31071 );
    and g22869 ( n27337 , n28967 , n9391 );
    and g22870 ( n40016 , n37830 , n22286 );
    or g22871 ( n19837 , n38029 , n42307 );
    and g22872 ( n8589 , n31989 , n20178 );
    and g22873 ( n28351 , n35553 , n39300 );
    or g22874 ( n42483 , n20921 , n16928 );
    and g22875 ( n3229 , n20945 , n26629 );
    or g22876 ( n3789 , n9021 , n25395 );
    or g22877 ( n40411 , n7396 , n21380 );
    and g22878 ( n16163 , n33697 , n13791 );
    xnor g22879 ( n29644 , n7628 , n32324 );
    nor g22880 ( n19902 , n29052 , n40342 );
    or g22881 ( n26937 , n5290 , n22740 );
    and g22882 ( n19232 , n1365 , n31748 );
    or g22883 ( n17860 , n14441 , n3469 );
    xnor g22884 ( n29383 , n10639 , n32024 );
    nor g22885 ( n25130 , n40915 , n10693 );
    or g22886 ( n34647 , n34411 , n35910 );
    not g22887 ( n11151 , n41595 );
    or g22888 ( n23645 , n31029 , n13085 );
    or g22889 ( n13853 , n39025 , n31120 );
    and g22890 ( n16901 , n35553 , n37019 );
    or g22891 ( n956 , n25959 , n21084 );
    and g22892 ( n25821 , n1936 , n11073 );
    nor g22893 ( n19237 , n28782 , n25863 );
    and g22894 ( n11231 , n35896 , n21408 );
    or g22895 ( n9690 , n23694 , n32969 );
    or g22896 ( n12717 , n9809 , n28508 );
    not g22897 ( n22557 , n34193 );
    or g22898 ( n14803 , n5323 , n34161 );
    xnor g22899 ( n34989 , n34731 , n23881 );
    nor g22900 ( n17626 , n8494 , n40431 );
    and g22901 ( n32320 , n20523 , n39586 );
    and g22902 ( n10976 , n24671 , n12067 );
    and g22903 ( n27923 , n12952 , n38448 );
    or g22904 ( n11193 , n13367 , n41706 );
    or g22905 ( n38671 , n23815 , n30868 );
    nor g22906 ( n29947 , n36667 , n19133 );
    nor g22907 ( n9335 , n5914 , n32361 );
    xnor g22908 ( n18720 , n40391 , n18710 );
    not g22909 ( n15620 , n19206 );
    nor g22910 ( n32445 , n15437 , n2020 );
    xnor g22911 ( n6843 , n784 , n31664 );
    nor g22912 ( n30356 , n24266 , n1989 );
    not g22913 ( n3898 , n4012 );
    and g22914 ( n5761 , n3032 , n42548 );
    and g22915 ( n18404 , n39390 , n11956 );
    or g22916 ( n7119 , n41433 , n35728 );
    not g22917 ( n37017 , n42803 );
    xnor g22918 ( n40249 , n898 , n41840 );
    nor g22919 ( n26942 , n35752 , n9694 );
    and g22920 ( n20399 , n5427 , n34327 );
    nor g22921 ( n10285 , n41281 , n36126 );
    and g22922 ( n8501 , n32331 , n6476 );
    or g22923 ( n19910 , n6858 , n16900 );
    or g22924 ( n19256 , n34719 , n5415 );
    and g22925 ( n38213 , n22260 , n18069 );
    xnor g22926 ( n306 , n4877 , n38748 );
    and g22927 ( n6174 , n42640 , n15058 );
    or g22928 ( n4137 , n36872 , n1823 );
    or g22929 ( n4134 , n31199 , n15292 );
    not g22930 ( n42478 , n1830 );
    or g22931 ( n41951 , n24957 , n33302 );
    and g22932 ( n14289 , n42000 , n32187 );
    nor g22933 ( n20802 , n14614 , n4797 );
    or g22934 ( n9756 , n16494 , n42793 );
    and g22935 ( n8545 , n34657 , n8553 );
    not g22936 ( n21373 , n7564 );
    and g22937 ( n39659 , n9878 , n7600 );
    or g22938 ( n1053 , n644 , n9416 );
    or g22939 ( n41044 , n7123 , n37880 );
    not g22940 ( n5048 , n9177 );
    not g22941 ( n6702 , n35607 );
    xnor g22942 ( n14841 , n42898 , n42017 );
    or g22943 ( n15536 , n41995 , n27831 );
    or g22944 ( n32497 , n37867 , n6290 );
    or g22945 ( n5878 , n39828 , n28731 );
    xnor g22946 ( n7268 , n15617 , n16008 );
    or g22947 ( n10773 , n3580 , n30361 );
    or g22948 ( n39278 , n12863 , n9857 );
    or g22949 ( n1964 , n36619 , n38281 );
    nor g22950 ( n8704 , n28489 , n42171 );
    and g22951 ( n14913 , n11162 , n11905 );
    or g22952 ( n32883 , n18314 , n28366 );
    xnor g22953 ( n2111 , n18927 , n2199 );
    and g22954 ( n15968 , n6824 , n22590 );
    or g22955 ( n8351 , n16033 , n36371 );
    or g22956 ( n11552 , n18093 , n37106 );
    nor g22957 ( n36570 , n6742 , n17919 );
    or g22958 ( n22630 , n2285 , n41740 );
    or g22959 ( n21376 , n15955 , n41240 );
    nor g22960 ( n32340 , n24745 , n10586 );
    not g22961 ( n2609 , n29377 );
    or g22962 ( n15679 , n6453 , n28127 );
    or g22963 ( n36642 , n4962 , n13697 );
    or g22964 ( n14935 , n11862 , n37779 );
    nor g22965 ( n34134 , n28593 , n31759 );
    or g22966 ( n32395 , n5818 , n14508 );
    and g22967 ( n8438 , n28871 , n42041 );
    nor g22968 ( n25314 , n24904 , n13322 );
    nor g22969 ( n9636 , n16251 , n14748 );
    and g22970 ( n31656 , n7503 , n28941 );
    or g22971 ( n21582 , n5396 , n38691 );
    or g22972 ( n17307 , n14503 , n28998 );
    not g22973 ( n22991 , n14233 );
    and g22974 ( n4441 , n12094 , n32074 );
    or g22975 ( n27622 , n38939 , n5864 );
    and g22976 ( n24226 , n22903 , n20803 );
    or g22977 ( n38292 , n27388 , n22266 );
    not g22978 ( n20453 , n5171 );
    or g22979 ( n10860 , n34059 , n40157 );
    xnor g22980 ( n13838 , n18496 , n19097 );
    or g22981 ( n25054 , n24879 , n29100 );
    not g22982 ( n40023 , n31540 );
    or g22983 ( n27436 , n20942 , n41819 );
    not g22984 ( n40350 , n12745 );
    and g22985 ( n9390 , n3161 , n41282 );
    and g22986 ( n42517 , n14613 , n2126 );
    or g22987 ( n29151 , n26386 , n35216 );
    or g22988 ( n38000 , n33976 , n33188 );
    nor g22989 ( n30844 , n2199 , n12104 );
    not g22990 ( n33640 , n29968 );
    or g22991 ( n36654 , n37028 , n32886 );
    and g22992 ( n24609 , n5743 , n6228 );
    and g22993 ( n7537 , n16034 , n41320 );
    not g22994 ( n9301 , n30775 );
    or g22995 ( n23372 , n17393 , n13426 );
    and g22996 ( n42649 , n11280 , n40964 );
    or g22997 ( n7576 , n19630 , n14699 );
    or g22998 ( n13364 , n23374 , n7500 );
    or g22999 ( n41409 , n41239 , n3743 );
    not g23000 ( n38983 , n38166 );
    or g23001 ( n1264 , n35526 , n17730 );
    or g23002 ( n42594 , n1291 , n27037 );
    xnor g23003 ( n14537 , n42064 , n32320 );
    and g23004 ( n9823 , n14731 , n132 );
    nor g23005 ( n12150 , n6978 , n41962 );
    or g23006 ( n2300 , n36446 , n34955 );
    not g23007 ( n5897 , n16158 );
    not g23008 ( n2921 , n402 );
    not g23009 ( n26579 , n25588 );
    and g23010 ( n41922 , n5236 , n41177 );
    xnor g23011 ( n37012 , n3277 , n9541 );
    or g23012 ( n17887 , n26795 , n35483 );
    xnor g23013 ( n14376 , n7922 , n22104 );
    not g23014 ( n16582 , n27463 );
    and g23015 ( n15287 , n3672 , n33644 );
    and g23016 ( n16657 , n18886 , n6920 );
    not g23017 ( n3030 , n39045 );
    or g23018 ( n2984 , n39614 , n22211 );
    or g23019 ( n13210 , n9905 , n22078 );
    or g23020 ( n36088 , n31584 , n23163 );
    xnor g23021 ( n21715 , n37030 , n18866 );
    and g23022 ( n27932 , n40810 , n24794 );
    and g23023 ( n9724 , n39638 , n35066 );
    nor g23024 ( n23321 , n26916 , n16293 );
    or g23025 ( n9407 , n27157 , n28341 );
    and g23026 ( n21747 , n4950 , n42150 );
    nor g23027 ( n16415 , n39410 , n27048 );
    or g23028 ( n30374 , n2227 , n34939 );
    or g23029 ( n17861 , n37339 , n34108 );
    or g23030 ( n1001 , n5795 , n33193 );
    nor g23031 ( n22033 , n13977 , n16317 );
    not g23032 ( n27808 , n25607 );
    and g23033 ( n23253 , n33822 , n16203 );
    or g23034 ( n28906 , n15663 , n31499 );
    or g23035 ( n6238 , n41045 , n24849 );
    or g23036 ( n9483 , n27832 , n32686 );
    nor g23037 ( n17105 , n11057 , n796 );
    nor g23038 ( n29902 , n38802 , n8190 );
    xnor g23039 ( n18744 , n4467 , n13223 );
    xnor g23040 ( n38863 , n14515 , n31619 );
    xnor g23041 ( n20056 , n784 , n3537 );
    xnor g23042 ( n4661 , n26544 , n9672 );
    xnor g23043 ( n32223 , n7320 , n38823 );
    xnor g23044 ( n31884 , n34691 , n37353 );
    or g23045 ( n33560 , n39930 , n21295 );
    not g23046 ( n14048 , n20190 );
    and g23047 ( n10364 , n33783 , n29246 );
    and g23048 ( n16659 , n39167 , n13755 );
    or g23049 ( n32822 , n22764 , n12152 );
    or g23050 ( n20963 , n23745 , n2188 );
    or g23051 ( n27332 , n7142 , n38232 );
    nor g23052 ( n37428 , n30424 , n14984 );
    or g23053 ( n30178 , n19867 , n16688 );
    or g23054 ( n38731 , n21586 , n15900 );
    or g23055 ( n14827 , n29922 , n40419 );
    or g23056 ( n27720 , n42269 , n4075 );
    nor g23057 ( n5633 , n2199 , n40676 );
    or g23058 ( n1557 , n12306 , n31769 );
    or g23059 ( n3968 , n15752 , n13254 );
    nor g23060 ( n17997 , n24617 , n26581 );
    and g23061 ( n746 , n26562 , n22141 );
    not g23062 ( n24061 , n11988 );
    not g23063 ( n12225 , n1866 );
    or g23064 ( n4828 , n11321 , n36862 );
    and g23065 ( n39304 , n19277 , n16423 );
    xnor g23066 ( n30058 , n36009 , n37585 );
    or g23067 ( n1198 , n20728 , n18449 );
    xnor g23068 ( n27129 , n20972 , n27015 );
    not g23069 ( n26794 , n39200 );
    and g23070 ( n19229 , n41951 , n21331 );
    not g23071 ( n19490 , n20879 );
    or g23072 ( n15841 , n34319 , n39819 );
    or g23073 ( n19620 , n11723 , n7395 );
    not g23074 ( n36094 , n25105 );
    or g23075 ( n14747 , n6398 , n11349 );
    and g23076 ( n13122 , n13499 , n7134 );
    nor g23077 ( n40292 , n6145 , n36812 );
    or g23078 ( n23284 , n14471 , n24677 );
    nor g23079 ( n14937 , n5320 , n20354 );
    or g23080 ( n10678 , n21667 , n1243 );
    not g23081 ( n27414 , n19671 );
    or g23082 ( n960 , n18230 , n20315 );
    and g23083 ( n23424 , n15480 , n19979 );
    or g23084 ( n6481 , n32618 , n12580 );
    and g23085 ( n25035 , n12564 , n29086 );
    and g23086 ( n17614 , n19058 , n7898 );
    not g23087 ( n27531 , n3831 );
    not g23088 ( n9161 , n10697 );
    or g23089 ( n37230 , n24394 , n16285 );
    and g23090 ( n7878 , n12474 , n35092 );
    and g23091 ( n7203 , n19274 , n17637 );
    or g23092 ( n8041 , n7429 , n9358 );
    or g23093 ( n32725 , n17980 , n3761 );
    or g23094 ( n8942 , n9125 , n10953 );
    or g23095 ( n38854 , n33824 , n17984 );
    not g23096 ( n10943 , n40136 );
    not g23097 ( n5073 , n8649 );
    or g23098 ( n33906 , n24432 , n37945 );
    not g23099 ( n38261 , n34330 );
    or g23100 ( n17378 , n36264 , n741 );
    or g23101 ( n18034 , n37948 , n5894 );
    xnor g23102 ( n33982 , n13930 , n17193 );
    and g23103 ( n33008 , n25037 , n1736 );
    or g23104 ( n12229 , n35619 , n4776 );
    and g23105 ( n32183 , n24433 , n21435 );
    or g23106 ( n23010 , n42115 , n9601 );
    or g23107 ( n8281 , n26963 , n30820 );
    or g23108 ( n37381 , n21170 , n42677 );
    xnor g23109 ( n30856 , n42064 , n25401 );
    nor g23110 ( n38013 , n7870 , n8808 );
    not g23111 ( n39123 , n19669 );
    or g23112 ( n41054 , n6797 , n42092 );
    and g23113 ( n13314 , n37812 , n28888 );
    and g23114 ( n20825 , n7434 , n41894 );
    or g23115 ( n24888 , n22330 , n4781 );
    xnor g23116 ( n6884 , n18678 , n29008 );
    not g23117 ( n27921 , n30794 );
    nor g23118 ( n6302 , n14375 , n13515 );
    or g23119 ( n5930 , n16052 , n10464 );
    or g23120 ( n14651 , n11955 , n15355 );
    or g23121 ( n6947 , n33262 , n32877 );
    or g23122 ( n20731 , n22276 , n34269 );
    not g23123 ( n21197 , n15004 );
    xnor g23124 ( n11726 , n3462 , n15307 );
    or g23125 ( n34237 , n5017 , n10097 );
    nor g23126 ( n37502 , n21568 , n22261 );
    or g23127 ( n8843 , n31622 , n13293 );
    nor g23128 ( n19055 , n6625 , n20105 );
    or g23129 ( n6896 , n4216 , n23696 );
    not g23130 ( n898 , n16780 );
    or g23131 ( n40072 , n40350 , n7151 );
    and g23132 ( n7826 , n33098 , n3894 );
    and g23133 ( n1151 , n40723 , n21909 );
    and g23134 ( n2671 , n8866 , n39892 );
    not g23135 ( n3264 , n8900 );
    and g23136 ( n42469 , n22822 , n39070 );
    nor g23137 ( n40579 , n1921 , n38983 );
    not g23138 ( n25959 , n11594 );
    not g23139 ( n34584 , n26142 );
    not g23140 ( n29713 , n18519 );
    not g23141 ( n42272 , n42554 );
    and g23142 ( n10690 , n19849 , n35958 );
    xnor g23143 ( n41865 , n37326 , n3844 );
    and g23144 ( n10593 , n21668 , n12114 );
    nor g23145 ( n30273 , n16991 , n7405 );
    not g23146 ( n20070 , n41208 );
    not g23147 ( n4660 , n30993 );
    not g23148 ( n32598 , n787 );
    and g23149 ( n1721 , n41188 , n28016 );
    or g23150 ( n2003 , n30365 , n23533 );
    not g23151 ( n30139 , n25247 );
    or g23152 ( n39231 , n29406 , n40488 );
    or g23153 ( n39028 , n2884 , n37600 );
    or g23154 ( n42155 , n7650 , n19823 );
    or g23155 ( n4072 , n2868 , n9873 );
    or g23156 ( n28843 , n781 , n25449 );
    and g23157 ( n18521 , n7291 , n9639 );
    or g23158 ( n9280 , n5603 , n33455 );
    nor g23159 ( n35188 , n32050 , n42552 );
    or g23160 ( n26468 , n20504 , n38175 );
    or g23161 ( n4146 , n12235 , n19975 );
    and g23162 ( n7070 , n10021 , n35699 );
    xnor g23163 ( n698 , n29644 , n16091 );
    or g23164 ( n4261 , n33289 , n21910 );
    or g23165 ( n12957 , n14791 , n7839 );
    xnor g23166 ( n9486 , n31848 , n19110 );
    xnor g23167 ( n33662 , n32407 , n15953 );
    or g23168 ( n15820 , n40716 , n29856 );
    or g23169 ( n16085 , n13548 , n31326 );
    and g23170 ( n28547 , n27084 , n42155 );
    or g23171 ( n30994 , n29991 , n34478 );
    and g23172 ( n1824 , n22152 , n15008 );
    not g23173 ( n36099 , n36979 );
    xnor g23174 ( n22691 , n35331 , n8354 );
    xnor g23175 ( n4881 , n14315 , n18605 );
    or g23176 ( n23474 , n13868 , n37589 );
    or g23177 ( n11929 , n30674 , n32327 );
    xnor g23178 ( n3456 , n21141 , n41962 );
    nor g23179 ( n42442 , n42465 , n17706 );
    or g23180 ( n21136 , n1294 , n30422 );
    or g23181 ( n13671 , n25180 , n37213 );
    nor g23182 ( n18028 , n17177 , n39978 );
    nor g23183 ( n7136 , n252 , n22205 );
    and g23184 ( n33666 , n40921 , n29706 );
    or g23185 ( n4932 , n34589 , n34623 );
    not g23186 ( n4795 , n36119 );
    not g23187 ( n23168 , n22097 );
    xnor g23188 ( n27724 , n33491 , n30338 );
    and g23189 ( n12175 , n1492 , n1198 );
    or g23190 ( n6740 , n42361 , n22886 );
    or g23191 ( n34266 , n36880 , n7473 );
    nor g23192 ( n37211 , n39320 , n18021 );
    not g23193 ( n34952 , n24478 );
    nor g23194 ( n9222 , n22726 , n42263 );
    and g23195 ( n30691 , n27387 , n35939 );
    nor g23196 ( n4810 , n40617 , n22014 );
    or g23197 ( n16179 , n35483 , n29338 );
    nor g23198 ( n639 , n25588 , n31466 );
    or g23199 ( n27636 , n25006 , n844 );
    and g23200 ( n1640 , n22870 , n15892 );
    nor g23201 ( n34671 , n37241 , n42226 );
    and g23202 ( n38772 , n33317 , n285 );
    or g23203 ( n10311 , n40323 , n26010 );
    or g23204 ( n36129 , n19318 , n22333 );
    nor g23205 ( n27435 , n24762 , n10451 );
    or g23206 ( n2702 , n39003 , n23098 );
    or g23207 ( n27985 , n20781 , n42188 );
    or g23208 ( n20192 , n16562 , n40888 );
    or g23209 ( n26978 , n12198 , n37761 );
    not g23210 ( n6462 , n29179 );
    or g23211 ( n16762 , n23137 , n328 );
    or g23212 ( n13169 , n22832 , n21697 );
    or g23213 ( n15867 , n7872 , n12220 );
    or g23214 ( n13822 , n27352 , n12167 );
    not g23215 ( n5168 , n17426 );
    nor g23216 ( n34764 , n5452 , n4232 );
    or g23217 ( n37886 , n6004 , n34403 );
    and g23218 ( n769 , n35125 , n25995 );
    and g23219 ( n31810 , n27229 , n2487 );
    and g23220 ( n31485 , n4079 , n20238 );
    or g23221 ( n14912 , n1656 , n36915 );
    nor g23222 ( n37275 , n7356 , n4911 );
    xnor g23223 ( n24978 , n34951 , n20767 );
    and g23224 ( n38980 , n29509 , n20965 );
    xnor g23225 ( n22710 , n105 , n8657 );
    not g23226 ( n34880 , n11896 );
    not g23227 ( n32289 , n7086 );
    or g23228 ( n6631 , n36369 , n27300 );
    xnor g23229 ( n38334 , n42725 , n16914 );
    xnor g23230 ( n22847 , n7572 , n657 );
    or g23231 ( n9058 , n36394 , n36425 );
    and g23232 ( n32547 , n13062 , n3413 );
    xnor g23233 ( n8054 , n39279 , n39936 );
    and g23234 ( n2209 , n13650 , n11241 );
    or g23235 ( n5853 , n4630 , n7265 );
    or g23236 ( n3897 , n16808 , n2507 );
    or g23237 ( n33688 , n11327 , n6002 );
    not g23238 ( n36010 , n25936 );
    or g23239 ( n605 , n15655 , n16659 );
    or g23240 ( n2389 , n15282 , n18305 );
    nor g23241 ( n35413 , n6885 , n23743 );
    and g23242 ( n33081 , n5169 , n1844 );
    xnor g23243 ( n14399 , n25426 , n8299 );
    or g23244 ( n16585 , n5910 , n22727 );
    or g23245 ( n6753 , n29832 , n14503 );
    and g23246 ( n5558 , n13399 , n37607 );
    and g23247 ( n12744 , n34395 , n9999 );
    nor g23248 ( n17016 , n6106 , n31030 );
    and g23249 ( n42073 , n8635 , n16300 );
    not g23250 ( n14206 , n14051 );
    or g23251 ( n21403 , n4050 , n15371 );
    or g23252 ( n5331 , n16287 , n3223 );
    nor g23253 ( n27983 , n2391 , n38419 );
    not g23254 ( n22313 , n15177 );
    not g23255 ( n19599 , n30902 );
    xnor g23256 ( n38004 , n28698 , n35540 );
    xnor g23257 ( n4569 , n10011 , n26934 );
    and g23258 ( n8951 , n39062 , n15645 );
    and g23259 ( n34918 , n24914 , n35087 );
    not g23260 ( n327 , n22763 );
    and g23261 ( n41163 , n18670 , n4860 );
    not g23262 ( n42748 , n13471 );
    or g23263 ( n7505 , n36468 , n22268 );
    not g23264 ( n17738 , n10819 );
    not g23265 ( n25143 , n21246 );
    or g23266 ( n31493 , n26196 , n42477 );
    or g23267 ( n15221 , n23619 , n37300 );
    nor g23268 ( n20597 , n41065 , n33504 );
    or g23269 ( n37205 , n38266 , n23872 );
    or g23270 ( n41229 , n4996 , n38379 );
    xnor g23271 ( n35925 , n453 , n410 );
    not g23272 ( n13140 , n7125 );
    or g23273 ( n8725 , n983 , n6117 );
    or g23274 ( n34929 , n8583 , n25475 );
    and g23275 ( n10788 , n38215 , n31743 );
    or g23276 ( n19685 , n9561 , n16377 );
    and g23277 ( n33798 , n9371 , n1603 );
    or g23278 ( n42044 , n40838 , n26409 );
    and g23279 ( n4160 , n21158 , n9650 );
    not g23280 ( n22077 , n1585 );
    or g23281 ( n15558 , n31286 , n22688 );
    and g23282 ( n13384 , n42785 , n21035 );
    xnor g23283 ( n22729 , n32841 , n36011 );
    or g23284 ( n1018 , n29027 , n27337 );
    not g23285 ( n7671 , n40228 );
    xnor g23286 ( n40777 , n16693 , n15212 );
    or g23287 ( n26216 , n7410 , n21399 );
    and g23288 ( n32715 , n20426 , n34977 );
    and g23289 ( n9887 , n18738 , n15521 );
    nor g23290 ( n41290 , n25373 , n41817 );
    xnor g23291 ( n10451 , n26 , n14200 );
    or g23292 ( n12709 , n41611 , n36305 );
    xnor g23293 ( n27928 , n35865 , n31160 );
    and g23294 ( n2129 , n42062 , n42621 );
    nor g23295 ( n1383 , n18866 , n10515 );
    and g23296 ( n33511 , n42878 , n30023 );
    nor g23297 ( n15763 , n4031 , n19681 );
    xnor g23298 ( n10956 , n35653 , n10252 );
    or g23299 ( n34802 , n4550 , n41990 );
    and g23300 ( n5085 , n38027 , n25563 );
    or g23301 ( n26928 , n21985 , n5578 );
    or g23302 ( n20400 , n33624 , n41022 );
    and g23303 ( n4391 , n24914 , n19398 );
    not g23304 ( n27133 , n2007 );
    or g23305 ( n22006 , n23971 , n25436 );
    not g23306 ( n27232 , n16899 );
    nor g23307 ( n14062 , n42692 , n25568 );
    or g23308 ( n12469 , n29633 , n12215 );
    or g23309 ( n18383 , n15342 , n24624 );
    xnor g23310 ( n8944 , n31992 , n31371 );
    or g23311 ( n40596 , n2608 , n38703 );
    and g23312 ( n17975 , n18999 , n4993 );
    or g23313 ( n1564 , n5408 , n20362 );
    or g23314 ( n29818 , n24156 , n4639 );
    nor g23315 ( n25664 , n3837 , n15452 );
    or g23316 ( n19678 , n36217 , n19444 );
    and g23317 ( n2286 , n27075 , n5958 );
    and g23318 ( n25966 , n28108 , n9589 );
    or g23319 ( n11119 , n25956 , n42544 );
    xnor g23320 ( n19330 , n14502 , n21324 );
    or g23321 ( n6721 , n17694 , n5036 );
    and g23322 ( n26212 , n36243 , n20967 );
    or g23323 ( n20943 , n12811 , n4625 );
    xnor g23324 ( n28469 , n784 , n5181 );
    or g23325 ( n34944 , n5861 , n27027 );
    or g23326 ( n32519 , n16684 , n35713 );
    and g23327 ( n25228 , n6941 , n2024 );
    and g23328 ( n10435 , n5393 , n8102 );
    nor g23329 ( n23518 , n19693 , n29851 );
    xnor g23330 ( n40465 , n24180 , n14462 );
    or g23331 ( n3418 , n20141 , n6073 );
    not g23332 ( n10033 , n31472 );
    or g23333 ( n595 , n24224 , n321 );
    or g23334 ( n21285 , n22371 , n248 );
    and g23335 ( n36522 , n39920 , n15201 );
    and g23336 ( n10149 , n17955 , n16303 );
    or g23337 ( n32777 , n27781 , n36205 );
    or g23338 ( n13610 , n36174 , n28556 );
    nor g23339 ( n598 , n33060 , n1055 );
    not g23340 ( n17327 , n39145 );
    nor g23341 ( n9939 , n36290 , n15926 );
    not g23342 ( n15874 , n11268 );
    or g23343 ( n11754 , n42405 , n41661 );
    and g23344 ( n16498 , n38089 , n17661 );
    nor g23345 ( n32329 , n23600 , n24090 );
    nor g23346 ( n13888 , n3109 , n15043 );
    or g23347 ( n34977 , n28294 , n806 );
    and g23348 ( n25107 , n26251 , n31484 );
    and g23349 ( n26432 , n34543 , n37592 );
    not g23350 ( n16745 , n3619 );
    or g23351 ( n37550 , n24828 , n2738 );
    or g23352 ( n2417 , n14209 , n41784 );
    and g23353 ( n40997 , n31189 , n10336 );
    and g23354 ( n31619 , n48 , n11198 );
    not g23355 ( n4725 , n7012 );
    nor g23356 ( n36662 , n23868 , n42221 );
    xnor g23357 ( n40832 , n7538 , n2828 );
    not g23358 ( n37639 , n39068 );
    not g23359 ( n40981 , n42389 );
    not g23360 ( n12823 , n26091 );
    and g23361 ( n32856 , n30133 , n13521 );
    and g23362 ( n27702 , n10388 , n24552 );
    and g23363 ( n18091 , n11991 , n22852 );
    or g23364 ( n10438 , n10447 , n36087 );
    and g23365 ( n34832 , n4385 , n35931 );
    or g23366 ( n22367 , n4535 , n27252 );
    or g23367 ( n18117 , n10284 , n1870 );
    nor g23368 ( n42386 , n38879 , n22832 );
    or g23369 ( n39116 , n8898 , n28005 );
    and g23370 ( n38319 , n25217 , n716 );
    and g23371 ( n22076 , n19668 , n713 );
    and g23372 ( n2216 , n12207 , n35123 );
    xnor g23373 ( n7641 , n19700 , n23005 );
    and g23374 ( n6429 , n16267 , n17541 );
    and g23375 ( n2770 , n17220 , n11994 );
    not g23376 ( n11923 , n28223 );
    and g23377 ( n34621 , n29647 , n8359 );
    xnor g23378 ( n2913 , n10595 , n34565 );
    or g23379 ( n28112 , n32711 , n36842 );
    or g23380 ( n15456 , n24053 , n29111 );
    not g23381 ( n14910 , n18899 );
    xnor g23382 ( n23252 , n42064 , n26399 );
    or g23383 ( n3996 , n1165 , n6088 );
    or g23384 ( n2186 , n14813 , n31371 );
    and g23385 ( n42263 , n25034 , n27672 );
    or g23386 ( n28823 , n36639 , n10704 );
    nor g23387 ( n39096 , n26231 , n28131 );
    or g23388 ( n1746 , n4713 , n30913 );
    or g23389 ( n22694 , n40728 , n3033 );
    nor g23390 ( n14568 , n17971 , n33002 );
    not g23391 ( n4149 , n31222 );
    or g23392 ( n581 , n33035 , n11349 );
    or g23393 ( n7308 , n36438 , n6912 );
    nor g23394 ( n11157 , n16693 , n18786 );
    not g23395 ( n36942 , n4178 );
    nor g23396 ( n29209 , n36996 , n31614 );
    or g23397 ( n30456 , n26038 , n5931 );
    and g23398 ( n35807 , n22309 , n13088 );
    and g23399 ( n21349 , n29622 , n36920 );
    or g23400 ( n19118 , n3018 , n7591 );
    or g23401 ( n26139 , n27503 , n14625 );
    or g23402 ( n6782 , n26686 , n21186 );
    or g23403 ( n4764 , n18376 , n32962 );
    or g23404 ( n19451 , n18988 , n758 );
    or g23405 ( n38798 , n39195 , n30401 );
    xnor g23406 ( n22633 , n33314 , n14913 );
    and g23407 ( n36537 , n6309 , n4765 );
    nor g23408 ( n40118 , n25826 , n5983 );
    nor g23409 ( n9889 , n24393 , n15815 );
    not g23410 ( n28661 , n26097 );
    nor g23411 ( n14822 , n34292 , n18004 );
    or g23412 ( n14744 , n34675 , n14172 );
    and g23413 ( n11764 , n9180 , n35553 );
    or g23414 ( n41075 , n5964 , n3694 );
    not g23415 ( n39182 , n24846 );
    xnor g23416 ( n3067 , n11168 , n28438 );
    or g23417 ( n42865 , n35139 , n12129 );
    or g23418 ( n5968 , n3405 , n4355 );
    or g23419 ( n18658 , n8689 , n40110 );
    or g23420 ( n14426 , n12531 , n25198 );
    or g23421 ( n23288 , n39489 , n18710 );
    or g23422 ( n33805 , n19530 , n35656 );
    or g23423 ( n29557 , n17589 , n38372 );
    or g23424 ( n8148 , n1360 , n19803 );
    or g23425 ( n6616 , n40462 , n41556 );
    or g23426 ( n4903 , n38623 , n9456 );
    xnor g23427 ( n20516 , n42725 , n25909 );
    and g23428 ( n10037 , n42714 , n1486 );
    or g23429 ( n10682 , n3809 , n26147 );
    xnor g23430 ( n4174 , n39722 , n12558 );
    xnor g23431 ( n35993 , n21381 , n25674 );
    and g23432 ( n9212 , n38536 , n25971 );
    xnor g23433 ( n20591 , n2072 , n41467 );
    xnor g23434 ( n23407 , n29854 , n38931 );
    and g23435 ( n17545 , n5560 , n16231 );
    not g23436 ( n19719 , n29319 );
    or g23437 ( n29527 , n2662 , n29977 );
    or g23438 ( n22870 , n2664 , n29439 );
    nor g23439 ( n26533 , n5964 , n1318 );
    nor g23440 ( n14038 , n33981 , n6919 );
    not g23441 ( n39935 , n6589 );
    nor g23442 ( n8056 , n7339 , n32494 );
    and g23443 ( n17706 , n30973 , n18538 );
    or g23444 ( n16667 , n36501 , n1788 );
    xnor g23445 ( n38033 , n21301 , n37232 );
    not g23446 ( n5302 , n32938 );
    not g23447 ( n13616 , n12476 );
    or g23448 ( n42622 , n35269 , n19566 );
    or g23449 ( n187 , n17514 , n6965 );
    or g23450 ( n12825 , n38723 , n2116 );
    or g23451 ( n12815 , n5877 , n1399 );
    or g23452 ( n5520 , n8147 , n40485 );
    not g23453 ( n22892 , n15439 );
    not g23454 ( n9655 , n2192 );
    or g23455 ( n28619 , n7511 , n29140 );
    and g23456 ( n28718 , n39147 , n23347 );
    xnor g23457 ( n5253 , n12487 , n12696 );
    not g23458 ( n32982 , n28269 );
    and g23459 ( n24817 , n19700 , n39824 );
    and g23460 ( n9194 , n41671 , n30966 );
    and g23461 ( n12341 , n16327 , n29871 );
    not g23462 ( n17399 , n37011 );
    nor g23463 ( n7797 , n41517 , n22036 );
    nor g23464 ( n11607 , n19300 , n24955 );
    not g23465 ( n20832 , n2932 );
    and g23466 ( n3097 , n30633 , n36187 );
    or g23467 ( n15774 , n6632 , n32053 );
    or g23468 ( n6017 , n41646 , n21240 );
    or g23469 ( n39371 , n13100 , n39098 );
    nor g23470 ( n34362 , n41534 , n5741 );
    nor g23471 ( n6612 , n17120 , n31552 );
    or g23472 ( n31086 , n25721 , n15748 );
    and g23473 ( n21784 , n34186 , n8566 );
    or g23474 ( n28938 , n13686 , n40871 );
    or g23475 ( n29977 , n30445 , n33537 );
    or g23476 ( n19575 , n42076 , n19163 );
    and g23477 ( n10103 , n27483 , n20828 );
    or g23478 ( n37400 , n39118 , n2732 );
    and g23479 ( n12856 , n39604 , n39211 );
    and g23480 ( n37364 , n17981 , n9028 );
    nor g23481 ( n25650 , n16598 , n34534 );
    or g23482 ( n13692 , n30496 , n26524 );
    or g23483 ( n38619 , n25049 , n9859 );
    or g23484 ( n29431 , n34767 , n18393 );
    not g23485 ( n19401 , n24816 );
    or g23486 ( n14533 , n20092 , n33599 );
    or g23487 ( n19553 , n40770 , n27715 );
    and g23488 ( n30657 , n846 , n16864 );
    nor g23489 ( n28229 , n2183 , n29111 );
    or g23490 ( n33785 , n11117 , n31227 );
    xnor g23491 ( n4673 , n40391 , n17721 );
    or g23492 ( n19816 , n40109 , n19989 );
    or g23493 ( n37203 , n38713 , n39439 );
    nor g23494 ( n8623 , n17647 , n22018 );
    or g23495 ( n34043 , n22615 , n12493 );
    or g23496 ( n27145 , n19942 , n32674 );
    or g23497 ( n18126 , n5419 , n9730 );
    not g23498 ( n542 , n36762 );
    xnor g23499 ( n29003 , n28464 , n16012 );
    not g23500 ( n5379 , n7599 );
    or g23501 ( n16022 , n8847 , n31961 );
    nor g23502 ( n31341 , n31217 , n27 );
    xnor g23503 ( n36824 , n17004 , n21851 );
    xnor g23504 ( n16722 , n32470 , n40853 );
    xnor g23505 ( n23345 , n36009 , n33462 );
    and g23506 ( n12560 , n26413 , n37412 );
    nor g23507 ( n32037 , n38879 , n18668 );
    or g23508 ( n13073 , n1522 , n18378 );
    not g23509 ( n2254 , n15890 );
    or g23510 ( n33939 , n9495 , n26927 );
    and g23511 ( n33646 , n42814 , n28857 );
    not g23512 ( n20487 , n1971 );
    not g23513 ( n29094 , n26706 );
    and g23514 ( n22017 , n7978 , n30221 );
    and g23515 ( n15703 , n17999 , n2281 );
    and g23516 ( n24477 , n41550 , n12644 );
    or g23517 ( n29737 , n19393 , n1906 );
    nor g23518 ( n6654 , n38938 , n26422 );
    nor g23519 ( n13513 , n16701 , n15146 );
    not g23520 ( n5001 , n36119 );
    and g23521 ( n7073 , n10235 , n37003 );
    or g23522 ( n37684 , n33981 , n10737 );
    or g23523 ( n24942 , n15149 , n33122 );
    not g23524 ( n21428 , n20038 );
    and g23525 ( n31664 , n14205 , n15777 );
    nor g23526 ( n29298 , n7339 , n39576 );
    nor g23527 ( n8307 , n38157 , n6544 );
    or g23528 ( n41817 , n15348 , n5556 );
    and g23529 ( n5026 , n4407 , n25807 );
    and g23530 ( n31482 , n5156 , n26894 );
    not g23531 ( n2171 , n4954 );
    and g23532 ( n24624 , n2481 , n5105 );
    and g23533 ( n35540 , n6610 , n5176 );
    nor g23534 ( n6151 , n32992 , n13995 );
    or g23535 ( n38126 , n35915 , n335 );
    xnor g23536 ( n2968 , n59 , n3406 );
    not g23537 ( n26921 , n15435 );
    not g23538 ( n12769 , n22454 );
    not g23539 ( n21134 , n2096 );
    or g23540 ( n2543 , n7086 , n10498 );
    xnor g23541 ( n20676 , n41013 , n7649 );
    and g23542 ( n23786 , n16972 , n24680 );
    not g23543 ( n8759 , n3425 );
    or g23544 ( n35211 , n10371 , n152 );
    not g23545 ( n40245 , n17935 );
    or g23546 ( n40851 , n40254 , n13129 );
    or g23547 ( n3878 , n16967 , n11711 );
    or g23548 ( n10225 , n2233 , n7654 );
    or g23549 ( n21189 , n37131 , n9555 );
    or g23550 ( n4247 , n30481 , n42531 );
    and g23551 ( n3167 , n3757 , n19534 );
    or g23552 ( n2115 , n25382 , n36652 );
    or g23553 ( n35810 , n35096 , n7066 );
    xnor g23554 ( n29855 , n21973 , n41443 );
    or g23555 ( n12376 , n4240 , n26407 );
    nor g23556 ( n33336 , n36435 , n14392 );
    and g23557 ( n22516 , n34832 , n21126 );
    and g23558 ( n26897 , n11564 , n39308 );
    and g23559 ( n38461 , n6463 , n13808 );
    not g23560 ( n39204 , n32999 );
    and g23561 ( n33795 , n13627 , n7910 );
    nor g23562 ( n19560 , n3136 , n2444 );
    or g23563 ( n32583 , n8138 , n2439 );
    not g23564 ( n32698 , n3442 );
    nor g23565 ( n26704 , n11760 , n19719 );
    or g23566 ( n13213 , n41544 , n12198 );
    xnor g23567 ( n1424 , n33413 , n27040 );
    or g23568 ( n1780 , n23122 , n24254 );
    nor g23569 ( n12083 , n2763 , n18837 );
    or g23570 ( n9321 , n23693 , n10165 );
    not g23571 ( n36052 , n41578 );
    not g23572 ( n15205 , n1825 );
    and g23573 ( n11181 , n29565 , n4067 );
    or g23574 ( n25379 , n34819 , n36087 );
    or g23575 ( n34969 , n7537 , n29884 );
    and g23576 ( n22832 , n30421 , n2349 );
    or g23577 ( n41576 , n5932 , n2476 );
    nor g23578 ( n2437 , n1474 , n39628 );
    or g23579 ( n39238 , n8926 , n20259 );
    nor g23580 ( n29378 , n26309 , n39090 );
    and g23581 ( n12783 , n14480 , n29297 );
    or g23582 ( n1212 , n20066 , n27698 );
    or g23583 ( n26703 , n41694 , n36098 );
    xnor g23584 ( n29563 , n11633 , n39802 );
    or g23585 ( n29048 , n34953 , n28118 );
    not g23586 ( n5406 , n33362 );
    not g23587 ( n34330 , n22812 );
    xnor g23588 ( n5469 , n1664 , n20229 );
    xnor g23589 ( n34072 , n9098 , n6071 );
    nor g23590 ( n24559 , n33794 , n13573 );
    or g23591 ( n18738 , n36924 , n28241 );
    not g23592 ( n23902 , n41955 );
    xnor g23593 ( n17913 , n16693 , n18004 );
    nor g23594 ( n25973 , n42104 , n10621 );
    or g23595 ( n33631 , n27162 , n3536 );
    xnor g23596 ( n38694 , n105 , n3975 );
    and g23597 ( n2559 , n34350 , n7487 );
    or g23598 ( n33109 , n27534 , n4355 );
    and g23599 ( n39128 , n10291 , n34168 );
    and g23600 ( n20048 , n40207 , n38746 );
    xnor g23601 ( n24866 , n12146 , n11674 );
    not g23602 ( n16728 , n35238 );
    or g23603 ( n26134 , n19990 , n28887 );
    and g23604 ( n7442 , n9675 , n30709 );
    or g23605 ( n3349 , n34194 , n4717 );
    or g23606 ( n243 , n11721 , n15245 );
    or g23607 ( n8051 , n19168 , n16483 );
    and g23608 ( n22401 , n1601 , n33500 );
    or g23609 ( n8773 , n13384 , n26354 );
    and g23610 ( n17719 , n38285 , n21525 );
    xnor g23611 ( n20223 , n36423 , n20218 );
    xnor g23612 ( n37032 , n25875 , n17754 );
    or g23613 ( n1713 , n27390 , n6244 );
    xnor g23614 ( n36074 , n22263 , n13059 );
    or g23615 ( n39535 , n22161 , n26795 );
    nor g23616 ( n14805 , n40757 , n7041 );
    xnor g23617 ( n25417 , n1762 , n27303 );
    and g23618 ( n26350 , n30151 , n34512 );
    or g23619 ( n24601 , n29135 , n9224 );
    or g23620 ( n27993 , n6110 , n37195 );
    and g23621 ( n9678 , n40631 , n16937 );
    and g23622 ( n10230 , n20421 , n35056 );
    or g23623 ( n30972 , n26116 , n11805 );
    not g23624 ( n8955 , n14302 );
    and g23625 ( n9550 , n36582 , n20336 );
    not g23626 ( n41532 , n40635 );
    xnor g23627 ( n22638 , n19164 , n37229 );
    or g23628 ( n40647 , n41433 , n3537 );
    or g23629 ( n36634 , n39367 , n40909 );
    or g23630 ( n27822 , n1201 , n42395 );
    not g23631 ( n15507 , n1760 );
    and g23632 ( n31419 , n14404 , n21392 );
    or g23633 ( n20000 , n37896 , n23955 );
    and g23634 ( n32688 , n26018 , n40267 );
    or g23635 ( n27882 , n23598 , n7712 );
    not g23636 ( n10448 , n8907 );
    or g23637 ( n40120 , n39489 , n29127 );
    and g23638 ( n20856 , n18512 , n25861 );
    or g23639 ( n3411 , n15657 , n34838 );
    not g23640 ( n28426 , n29245 );
    nor g23641 ( n5201 , n14471 , n13147 );
    or g23642 ( n10618 , n30859 , n2034 );
    not g23643 ( n1197 , n3209 );
    xnor g23644 ( n15241 , n20972 , n23655 );
    or g23645 ( n18440 , n22470 , n38521 );
    or g23646 ( n24392 , n31371 , n18070 );
    nor g23647 ( n41008 , n34419 , n6220 );
    or g23648 ( n38469 , n41497 , n15021 );
    xnor g23649 ( n16704 , n5041 , n42518 );
    and g23650 ( n35856 , n42883 , n41606 );
    or g23651 ( n1135 , n3786 , n1468 );
    xnor g23652 ( n17692 , n33794 , n28722 );
    or g23653 ( n21194 , n31591 , n36087 );
    and g23654 ( n39196 , n38891 , n33195 );
    nor g23655 ( n40094 , n35950 , n7887 );
    or g23656 ( n35237 , n39108 , n30511 );
    nor g23657 ( n25722 , n2753 , n11643 );
    xnor g23658 ( n22149 , n11014 , n9736 );
    xnor g23659 ( n32643 , n36009 , n42476 );
    not g23660 ( n9900 , n10748 );
    and g23661 ( n19058 , n17294 , n18017 );
    nor g23662 ( n33167 , n33227 , n32747 );
    and g23663 ( n37699 , n34291 , n22446 );
    not g23664 ( n5578 , n40246 );
    nor g23665 ( n10606 , n15118 , n4892 );
    and g23666 ( n28786 , n35402 , n2106 );
    nor g23667 ( n39540 , n405 , n27207 );
    and g23668 ( n25061 , n19881 , n6350 );
    xnor g23669 ( n31115 , n6621 , n24953 );
    nor g23670 ( n20418 , n1507 , n24901 );
    and g23671 ( n16256 , n92 , n3753 );
    and g23672 ( n4887 , n5711 , n21429 );
    not g23673 ( n3701 , n39846 );
    or g23674 ( n42500 , n41433 , n33709 );
    nor g23675 ( n19511 , n5896 , n24807 );
    or g23676 ( n21122 , n33648 , n24250 );
    xnor g23677 ( n13919 , n17427 , n28918 );
    and g23678 ( n37578 , n42832 , n32926 );
    not g23679 ( n9686 , n2497 );
    not g23680 ( n29322 , n40655 );
    xnor g23681 ( n1222 , n4334 , n12555 );
    or g23682 ( n31726 , n4750 , n23735 );
    or g23683 ( n34259 , n6004 , n32223 );
    nor g23684 ( n38373 , n4921 , n25800 );
    and g23685 ( n816 , n17047 , n5866 );
    not g23686 ( n9456 , n17327 );
    xnor g23687 ( n31078 , n41098 , n26838 );
    or g23688 ( n13740 , n22243 , n26924 );
    xnor g23689 ( n25076 , n6767 , n38963 );
    or g23690 ( n9296 , n32293 , n31497 );
    and g23691 ( n40959 , n434 , n29775 );
    and g23692 ( n13318 , n24939 , n39229 );
    and g23693 ( n6999 , n13272 , n28394 );
    nor g23694 ( n11522 , n18866 , n31459 );
    or g23695 ( n2019 , n39297 , n42469 );
    or g23696 ( n9805 , n29540 , n9673 );
    or g23697 ( n33116 , n33926 , n38799 );
    or g23698 ( n41798 , n21938 , n16559 );
    or g23699 ( n2544 , n23452 , n13819 );
    not g23700 ( n31356 , n33039 );
    xnor g23701 ( n12648 , n29724 , n6856 );
    xnor g23702 ( n10513 , n42728 , n30755 );
    not g23703 ( n946 , n42273 );
    and g23704 ( n20035 , n34707 , n20869 );
    nor g23705 ( n4273 , n22563 , n29137 );
    or g23706 ( n30156 , n27753 , n13343 );
    not g23707 ( n10548 , n21673 );
    or g23708 ( n7638 , n30346 , n40295 );
    or g23709 ( n24802 , n13955 , n36657 );
    xnor g23710 ( n24984 , n11426 , n9901 );
    or g23711 ( n270 , n21914 , n27522 );
    not g23712 ( n34955 , n263 );
    not g23713 ( n6368 , n22119 );
    and g23714 ( n9277 , n35875 , n15749 );
    and g23715 ( n26276 , n36743 , n13890 );
    or g23716 ( n3144 , n17850 , n41905 );
    or g23717 ( n37458 , n27963 , n8828 );
    or g23718 ( n4739 , n3311 , n12994 );
    not g23719 ( n3539 , n21183 );
    not g23720 ( n17006 , n42904 );
    or g23721 ( n36333 , n2608 , n5266 );
    xnor g23722 ( n33413 , n2339 , n10755 );
    nor g23723 ( n27276 , n9616 , n29778 );
    or g23724 ( n35099 , n31924 , n36082 );
    and g23725 ( n3267 , n2154 , n17778 );
    or g23726 ( n16795 , n519 , n1688 );
    nor g23727 ( n33361 , n25588 , n34676 );
    or g23728 ( n40201 , n34793 , n15702 );
    not g23729 ( n22106 , n25223 );
    or g23730 ( n37587 , n35951 , n13495 );
    or g23731 ( n27229 , n3485 , n32405 );
    nor g23732 ( n30025 , n917 , n35098 );
    nor g23733 ( n23153 , n39110 , n17995 );
    or g23734 ( n561 , n30835 , n9494 );
    or g23735 ( n41224 , n35386 , n10354 );
    xnor g23736 ( n8552 , n21244 , n1212 );
    not g23737 ( n19414 , n37004 );
    and g23738 ( n15212 , n25923 , n8917 );
    nor g23739 ( n841 , n37536 , n20838 );
    and g23740 ( n33705 , n23512 , n40667 );
    and g23741 ( n16966 , n42689 , n9834 );
    not g23742 ( n41280 , n6782 );
    or g23743 ( n35623 , n12950 , n30626 );
    not g23744 ( n16973 , n27257 );
    and g23745 ( n8977 , n42114 , n3631 );
    not g23746 ( n102 , n37595 );
    or g23747 ( n16025 , n2517 , n28067 );
    not g23748 ( n23473 , n40651 );
    not g23749 ( n42186 , n3048 );
    not g23750 ( n41328 , n16797 );
    and g23751 ( n11964 , n23033 , n41542 );
    or g23752 ( n5715 , n40156 , n38211 );
    not g23753 ( n4659 , n31785 );
    xnor g23754 ( n1305 , n36444 , n11834 );
    or g23755 ( n19238 , n24588 , n34172 );
    and g23756 ( n12636 , n9266 , n273 );
    and g23757 ( n19318 , n5777 , n25218 );
    or g23758 ( n36138 , n30612 , n7899 );
    not g23759 ( n38792 , n6646 );
    or g23760 ( n2707 , n7665 , n28551 );
    and g23761 ( n16467 , n40279 , n9169 );
    or g23762 ( n24935 , n23736 , n36652 );
    or g23763 ( n4571 , n19281 , n13256 );
    nor g23764 ( n3917 , n11398 , n24171 );
    nor g23765 ( n2489 , n31187 , n18240 );
    and g23766 ( n1290 , n13266 , n9993 );
    or g23767 ( n37750 , n6957 , n37180 );
    or g23768 ( n42106 , n18860 , n25736 );
    not g23769 ( n30742 , n13002 );
    or g23770 ( n39960 , n40237 , n32970 );
    or g23771 ( n27125 , n13731 , n7862 );
    not g23772 ( n28901 , n15790 );
    nor g23773 ( n38687 , n39700 , n1837 );
    not g23774 ( n10014 , n20053 );
    nor g23775 ( n16224 , n24441 , n30757 );
    and g23776 ( n12520 , n14046 , n5862 );
    or g23777 ( n28764 , n34495 , n36296 );
    not g23778 ( n16573 , n13042 );
    or g23779 ( n16835 , n18775 , n9703 );
    xnor g23780 ( n4192 , n27433 , n36331 );
    not g23781 ( n915 , n3879 );
    and g23782 ( n26120 , n34306 , n39857 );
    and g23783 ( n22119 , n14924 , n30907 );
    and g23784 ( n10476 , n4214 , n15496 );
    and g23785 ( n36771 , n41753 , n18289 );
    and g23786 ( n23849 , n18977 , n20960 );
    nor g23787 ( n38205 , n35361 , n3727 );
    or g23788 ( n27961 , n17313 , n23032 );
    not g23789 ( n11438 , n7158 );
    xnor g23790 ( n12370 , n7425 , n17934 );
    and g23791 ( n11661 , n22232 , n5944 );
    and g23792 ( n14873 , n8166 , n8943 );
    and g23793 ( n7652 , n445 , n37297 );
    or g23794 ( n4078 , n32278 , n14048 );
    or g23795 ( n20713 , n26116 , n30777 );
    not g23796 ( n41300 , n33196 );
    and g23797 ( n13782 , n32492 , n40883 );
    not g23798 ( n29681 , n15526 );
    and g23799 ( n22645 , n36759 , n20125 );
    nor g23800 ( n18753 , n2199 , n13313 );
    nor g23801 ( n19841 , n15070 , n27735 );
    and g23802 ( n1712 , n17178 , n37717 );
    and g23803 ( n1896 , n28512 , n29064 );
    and g23804 ( n40244 , n29900 , n37789 );
    and g23805 ( n121 , n37393 , n5221 );
    nor g23806 ( n11971 , n2467 , n41096 );
    or g23807 ( n37757 , n8494 , n23602 );
    and g23808 ( n9479 , n15174 , n34230 );
    not g23809 ( n38485 , n33639 );
    and g23810 ( n17088 , n28660 , n29624 );
    not g23811 ( n16742 , n246 );
    not g23812 ( n13176 , n9754 );
    or g23813 ( n21664 , n25752 , n39141 );
    or g23814 ( n5703 , n5408 , n6892 );
    or g23815 ( n199 , n33073 , n5163 );
    and g23816 ( n37344 , n18561 , n26007 );
    not g23817 ( n8194 , n28003 );
    nor g23818 ( n20730 , n4442 , n21108 );
    or g23819 ( n4957 , n23988 , n26975 );
    nor g23820 ( n37462 , n22147 , n41165 );
    or g23821 ( n3673 , n27884 , n5678 );
    nor g23822 ( n15320 , n606 , n208 );
    not g23823 ( n13280 , n29006 );
    or g23824 ( n3269 , n328 , n864 );
    and g23825 ( n16711 , n5872 , n36342 );
    and g23826 ( n11205 , n5314 , n10741 );
    and g23827 ( n36485 , n19502 , n36715 );
    and g23828 ( n22551 , n5871 , n16279 );
    nor g23829 ( n31805 , n37830 , n22286 );
    nor g23830 ( n21804 , n22519 , n15948 );
    and g23831 ( n31427 , n32920 , n936 );
    xnor g23832 ( n22400 , n13735 , n38919 );
    or g23833 ( n10446 , n29564 , n11178 );
    not g23834 ( n35857 , n40407 );
    and g23835 ( n34499 , n21649 , n20665 );
    and g23836 ( n33036 , n5235 , n41068 );
    or g23837 ( n27376 , n30820 , n25716 );
    or g23838 ( n29193 , n19744 , n39576 );
    and g23839 ( n26376 , n31615 , n14100 );
    or g23840 ( n24324 , n42706 , n41712 );
    and g23841 ( n40375 , n21459 , n17828 );
    or g23842 ( n32014 , n39941 , n7309 );
    and g23843 ( n18893 , n29746 , n4891 );
    and g23844 ( n24875 , n12901 , n9454 );
    or g23845 ( n30503 , n30825 , n8704 );
    not g23846 ( n40902 , n36119 );
    or g23847 ( n6107 , n32553 , n4043 );
    or g23848 ( n35351 , n36504 , n7321 );
    or g23849 ( n20114 , n30403 , n39603 );
    not g23850 ( n42273 , n4178 );
    xnor g23851 ( n7068 , n26579 , n8169 );
    and g23852 ( n7309 , n17269 , n12360 );
    not g23853 ( n22205 , n22444 );
    or g23854 ( n42257 , n34445 , n25987 );
    nor g23855 ( n33383 , n8968 , n12670 );
    not g23856 ( n8809 , n5776 );
    not g23857 ( n10778 , n19412 );
    nor g23858 ( n3398 , n5964 , n34133 );
    or g23859 ( n16819 , n26849 , n28809 );
    xnor g23860 ( n24999 , n542 , n40859 );
    or g23861 ( n36125 , n981 , n5806 );
    or g23862 ( n42832 , n26500 , n3936 );
    xnor g23863 ( n6345 , n9142 , n22676 );
    and g23864 ( n28360 , n10123 , n19220 );
    or g23865 ( n28121 , n36052 , n642 );
    or g23866 ( n6242 , n15227 , n1747 );
    and g23867 ( n33787 , n18530 , n9965 );
    or g23868 ( n15677 , n20096 , n20001 );
    and g23869 ( n38125 , n39154 , n16361 );
    or g23870 ( n17594 , n2666 , n34652 );
    or g23871 ( n32098 , n28417 , n22379 );
    nor g23872 ( n10067 , n17120 , n23842 );
    not g23873 ( n17828 , n23981 );
    and g23874 ( n32092 , n39339 , n17789 );
    and g23875 ( n11271 , n19797 , n6021 );
    and g23876 ( n4578 , n35974 , n9981 );
    or g23877 ( n3871 , n35732 , n10141 );
    and g23878 ( n39663 , n5612 , n30198 );
    and g23879 ( n5673 , n14636 , n2629 );
    and g23880 ( n14902 , n1313 , n29331 );
    xnor g23881 ( n34957 , n9448 , n13003 );
    not g23882 ( n42699 , n1879 );
    and g23883 ( n10485 , n37079 , n38118 );
    not g23884 ( n3382 , n40354 );
    not g23885 ( n40713 , n27987 );
    or g23886 ( n23887 , n17744 , n7814 );
    or g23887 ( n39971 , n23929 , n25521 );
    or g23888 ( n40905 , n17888 , n42873 );
    and g23889 ( n506 , n13780 , n13894 );
    or g23890 ( n26636 , n25487 , n12081 );
    or g23891 ( n38966 , n13310 , n24114 );
    or g23892 ( n24589 , n13752 , n2034 );
    and g23893 ( n29864 , n1737 , n34408 );
    and g23894 ( n23210 , n21382 , n10474 );
    not g23895 ( n3603 , n16005 );
    or g23896 ( n32569 , n21006 , n752 );
    xnor g23897 ( n3098 , n34329 , n3554 );
    and g23898 ( n7370 , n15273 , n11893 );
    not g23899 ( n39433 , n18331 );
    and g23900 ( n2415 , n25884 , n35400 );
    xnor g23901 ( n9528 , n16693 , n41823 );
    and g23902 ( n32970 , n32393 , n2914 );
    or g23903 ( n12107 , n6950 , n658 );
    or g23904 ( n7036 , n15717 , n25937 );
    xnor g23905 ( n6448 , n330 , n36080 );
    and g23906 ( n26713 , n26294 , n21353 );
    nor g23907 ( n21579 , n27439 , n38980 );
    and g23908 ( n21914 , n24409 , n25823 );
    or g23909 ( n12088 , n10769 , n38467 );
    not g23910 ( n11267 , n8933 );
    or g23911 ( n33503 , n16581 , n25831 );
    nor g23912 ( n1107 , n24064 , n10037 );
    not g23913 ( n33433 , n19651 );
    not g23914 ( n8991 , n8256 );
    nor g23915 ( n32230 , n34565 , n15498 );
    or g23916 ( n27726 , n28482 , n2092 );
    or g23917 ( n40370 , n14948 , n25765 );
    xnor g23918 ( n631 , n18530 , n31697 );
    and g23919 ( n17988 , n14096 , n30933 );
    or g23920 ( n15773 , n9154 , n10865 );
    or g23921 ( n23187 , n21288 , n8049 );
    or g23922 ( n30096 , n26122 , n35688 );
    nor g23923 ( n35445 , n38879 , n10222 );
    xnor g23924 ( n27394 , n16473 , n34688 );
    xnor g23925 ( n13275 , n40852 , n17390 );
    or g23926 ( n4354 , n39966 , n5372 );
    and g23927 ( n15748 , n5950 , n35341 );
    or g23928 ( n10369 , n12130 , n32024 );
    or g23929 ( n29875 , n17747 , n34949 );
    nor g23930 ( n26870 , n18928 , n38665 );
    or g23931 ( n41744 , n19196 , n30090 );
    and g23932 ( n32527 , n36046 , n38012 );
    and g23933 ( n21869 , n22781 , n4104 );
    or g23934 ( n436 , n24656 , n42806 );
    or g23935 ( n1079 , n7406 , n32675 );
    and g23936 ( n29187 , n899 , n41825 );
    not g23937 ( n2015 , n7709 );
    not g23938 ( n3363 , n3997 );
    or g23939 ( n34689 , n28297 , n27311 );
    nor g23940 ( n9066 , n9668 , n27513 );
    or g23941 ( n13097 , n36306 , n36344 );
    or g23942 ( n8553 , n6423 , n34418 );
    nor g23943 ( n35800 , n9276 , n37237 );
    or g23944 ( n20912 , n38568 , n32346 );
    and g23945 ( n34051 , n7629 , n6674 );
    or g23946 ( n24920 , n17941 , n18762 );
    or g23947 ( n5345 , n33170 , n30487 );
    and g23948 ( n27390 , n16539 , n25889 );
    and g23949 ( n29227 , n41965 , n21858 );
    or g23950 ( n26328 , n28103 , n25001 );
    or g23951 ( n39542 , n40554 , n24038 );
    not g23952 ( n9784 , n11697 );
    xnor g23953 ( n28613 , n4537 , n25045 );
    or g23954 ( n2406 , n392 , n2539 );
    xnor g23955 ( n5575 , n42799 , n40030 );
    or g23956 ( n35621 , n21175 , n31676 );
    not g23957 ( n18761 , n34711 );
    and g23958 ( n21225 , n16475 , n11649 );
    or g23959 ( n2273 , n42626 , n4926 );
    or g23960 ( n37618 , n41773 , n18947 );
    or g23961 ( n41737 , n12226 , n21334 );
    nor g23962 ( n29528 , n1448 , n21388 );
    or g23963 ( n10039 , n4288 , n5583 );
    or g23964 ( n10188 , n38119 , n17766 );
    xnor g23965 ( n22192 , n40191 , n42202 );
    not g23966 ( n7410 , n7508 );
    or g23967 ( n34830 , n12377 , n33826 );
    nor g23968 ( n29955 , n15572 , n1496 );
    nor g23969 ( n6924 , n38932 , n36525 );
    or g23970 ( n19312 , n27503 , n3078 );
    not g23971 ( n10320 , n38108 );
    or g23972 ( n18327 , n27825 , n42152 );
    or g23973 ( n5966 , n28713 , n792 );
    or g23974 ( n19031 , n18443 , n2209 );
    nor g23975 ( n8852 , n27718 , n27407 );
    or g23976 ( n3573 , n18747 , n35526 );
    or g23977 ( n13578 , n6078 , n7414 );
    or g23978 ( n35448 , n29752 , n41487 );
    and g23979 ( n13076 , n23083 , n21554 );
    and g23980 ( n17898 , n16091 , n29644 );
    or g23981 ( n28958 , n6929 , n35453 );
    xnor g23982 ( n34056 , n27245 , n15869 );
    and g23983 ( n29218 , n19591 , n3674 );
    xnor g23984 ( n19839 , n10316 , n19900 );
    and g23985 ( n41730 , n36346 , n15856 );
    nor g23986 ( n35899 , n24289 , n13579 );
    and g23987 ( n34070 , n28458 , n32359 );
    not g23988 ( n34739 , n7449 );
    xnor g23989 ( n16604 , n38685 , n7994 );
    and g23990 ( n22553 , n13355 , n16126 );
    not g23991 ( n9203 , n34230 );
    or g23992 ( n40996 , n18921 , n17088 );
    nor g23993 ( n24585 , n1656 , n9263 );
    or g23994 ( n3596 , n25290 , n4718 );
    or g23995 ( n11588 , n16004 , n6851 );
    not g23996 ( n18678 , n41427 );
    or g23997 ( n30231 , n38870 , n36203 );
    and g23998 ( n2639 , n8936 , n17281 );
    or g23999 ( n15853 , n32217 , n21364 );
    or g24000 ( n27768 , n14343 , n29803 );
    xnor g24001 ( n39518 , n7922 , n41605 );
    or g24002 ( n9946 , n35811 , n34551 );
    not g24003 ( n40359 , n1215 );
    not g24004 ( n7139 , n21918 );
    and g24005 ( n31094 , n1528 , n31481 );
    or g24006 ( n12642 , n28528 , n41413 );
    and g24007 ( n11890 , n32948 , n37480 );
    not g24008 ( n31848 , n10614 );
    xnor g24009 ( n18339 , n26412 , n6030 );
    not g24010 ( n19547 , n10779 );
    xnor g24011 ( n42310 , n27064 , n23458 );
    nor g24012 ( n14724 , n13895 , n2456 );
    not g24013 ( n12106 , n42816 );
    nor g24014 ( n17428 , n6573 , n35933 );
    nor g24015 ( n36470 , n32299 , n11195 );
    or g24016 ( n20966 , n13401 , n31597 );
    and g24017 ( n39186 , n23485 , n8884 );
    not g24018 ( n5070 , n2979 );
    or g24019 ( n35136 , n24283 , n10231 );
    or g24020 ( n40336 , n34909 , n28960 );
    or g24021 ( n40917 , n33071 , n17896 );
    nor g24022 ( n32389 , n1507 , n38405 );
    or g24023 ( n34845 , n34329 , n601 );
    or g24024 ( n3407 , n40713 , n20591 );
    or g24025 ( n23391 , n370 , n25647 );
    nor g24026 ( n36211 , n18866 , n29097 );
    and g24027 ( n26903 , n11351 , n11303 );
    or g24028 ( n14852 , n12221 , n35157 );
    or g24029 ( n20859 , n18716 , n39466 );
    or g24030 ( n30553 , n22485 , n7558 );
    and g24031 ( n34703 , n5460 , n33966 );
    or g24032 ( n5690 , n11147 , n5313 );
    or g24033 ( n41134 , n35772 , n6272 );
    or g24034 ( n7514 , n19911 , n33452 );
    or g24035 ( n39838 , n23817 , n41668 );
    not g24036 ( n29538 , n35850 );
    xnor g24037 ( n8827 , n42127 , n40286 );
    and g24038 ( n9487 , n13029 , n1966 );
    nor g24039 ( n33414 , n6011 , n1502 );
    nor g24040 ( n33218 , n23491 , n40252 );
    xnor g24041 ( n34947 , n37922 , n3598 );
    or g24042 ( n26186 , n41938 , n35726 );
    and g24043 ( n15107 , n27288 , n2610 );
    or g24044 ( n24192 , n37380 , n37120 );
    xnor g24045 ( n19994 , n38257 , n38157 );
    or g24046 ( n28948 , n7175 , n2875 );
    and g24047 ( n37439 , n28589 , n34067 );
    or g24048 ( n4026 , n4318 , n7142 );
    not g24049 ( n25420 , n25561 );
    or g24050 ( n39818 , n24745 , n6839 );
    or g24051 ( n33064 , n34101 , n4578 );
    or g24052 ( n35753 , n8847 , n19097 );
    or g24053 ( n37159 , n40529 , n13632 );
    not g24054 ( n28883 , n36151 );
    or g24055 ( n8152 , n31127 , n904 );
    and g24056 ( n632 , n1437 , n29758 );
    or g24057 ( n6058 , n41193 , n5513 );
    or g24058 ( n30791 , n22946 , n39204 );
    and g24059 ( n5933 , n35000 , n19896 );
    or g24060 ( n31369 , n29395 , n9867 );
    xnor g24061 ( n41626 , n18840 , n12284 );
    and g24062 ( n20004 , n39119 , n26138 );
    xnor g24063 ( n34354 , n28083 , n9009 );
    or g24064 ( n16036 , n14769 , n10359 );
    or g24065 ( n7049 , n28074 , n15581 );
    or g24066 ( n27569 , n39296 , n2861 );
    or g24067 ( n22587 , n34877 , n18436 );
    xnor g24068 ( n111 , n40 , n21820 );
    and g24069 ( n36765 , n32615 , n18695 );
    or g24070 ( n1523 , n16967 , n34324 );
    not g24071 ( n56 , n13857 );
    and g24072 ( n32942 , n25894 , n22897 );
    or g24073 ( n700 , n30452 , n38657 );
    not g24074 ( n40811 , n8699 );
    nor g24075 ( n20911 , n29113 , n17943 );
    or g24076 ( n32515 , n16586 , n26423 );
    or g24077 ( n33731 , n40418 , n2999 );
    and g24078 ( n11461 , n38243 , n31735 );
    and g24079 ( n41143 , n18506 , n6416 );
    xnor g24080 ( n39079 , n2837 , n1311 );
    or g24081 ( n42087 , n11079 , n19627 );
    or g24082 ( n32616 , n26354 , n41080 );
    and g24083 ( n8150 , n2778 , n34203 );
    not g24084 ( n2637 , n35871 );
    or g24085 ( n1878 , n5896 , n2781 );
    and g24086 ( n20746 , n7081 , n5172 );
    or g24087 ( n42559 , n17654 , n41924 );
    and g24088 ( n42881 , n27014 , n458 );
    not g24089 ( n40915 , n28880 );
    nor g24090 ( n11272 , n29423 , n33623 );
    not g24091 ( n31263 , n23184 );
    not g24092 ( n31386 , n3973 );
    or g24093 ( n18559 , n15556 , n12831 );
    xnor g24094 ( n13548 , n16960 , n23976 );
    xnor g24095 ( n5490 , n36009 , n8447 );
    and g24096 ( n16007 , n29148 , n27183 );
    not g24097 ( n30035 , n28350 );
    and g24098 ( n37879 , n33570 , n31163 );
    and g24099 ( n26877 , n11086 , n5837 );
    xnor g24100 ( n7262 , n31989 , n36061 );
    or g24101 ( n41422 , n19744 , n16631 );
    and g24102 ( n30067 , n21073 , n33112 );
    not g24103 ( n41657 , n42837 );
    and g24104 ( n14385 , n16907 , n5767 );
    nor g24105 ( n32269 , n41133 , n18943 );
    and g24106 ( n27267 , n4813 , n32989 );
    and g24107 ( n4094 , n12335 , n34064 );
    xnor g24108 ( n39721 , n27245 , n30974 );
    or g24109 ( n13778 , n17728 , n9627 );
    and g24110 ( n41822 , n33420 , n33315 );
    xnor g24111 ( n37905 , n3812 , n34981 );
    and g24112 ( n10979 , n41285 , n17501 );
    or g24113 ( n13591 , n1253 , n22614 );
    or g24114 ( n17147 , n28785 , n449 );
    not g24115 ( n2477 , n26685 );
    xnor g24116 ( n9352 , n34731 , n4766 );
    or g24117 ( n5783 , n38921 , n36459 );
    not g24118 ( n21126 , n22156 );
    and g24119 ( n16306 , n1599 , n40582 );
    nor g24120 ( n15049 , n10489 , n10808 );
    xnor g24121 ( n184 , n26496 , n2749 );
    nor g24122 ( n26101 , n16598 , n30471 );
    nor g24123 ( n38421 , n12878 , n1368 );
    not g24124 ( n14039 , n28857 );
    not g24125 ( n11783 , n4825 );
    or g24126 ( n40666 , n40274 , n12255 );
    and g24127 ( n22723 , n7968 , n8230 );
    not g24128 ( n19936 , n20896 );
    nor g24129 ( n41873 , n228 , n27132 );
    xnor g24130 ( n38323 , n7421 , n38102 );
    xnor g24131 ( n38489 , n16035 , n10767 );
    or g24132 ( n37700 , n34565 , n23582 );
    nor g24133 ( n41494 , n38770 , n3367 );
    not g24134 ( n18519 , n12465 );
    or g24135 ( n28855 , n32503 , n32800 );
    nor g24136 ( n42109 , n34625 , n36822 );
    nor g24137 ( n17581 , n2263 , n20821 );
    xnor g24138 ( n16670 , n1768 , n42704 );
    nor g24139 ( n42069 , n25544 , n24096 );
    or g24140 ( n18340 , n41819 , n2448 );
    and g24141 ( n18861 , n27653 , n20129 );
    and g24142 ( n76 , n31495 , n19216 );
    or g24143 ( n24257 , n21034 , n3705 );
    and g24144 ( n41022 , n40341 , n5929 );
    or g24145 ( n22926 , n37647 , n27006 );
    not g24146 ( n40372 , n27476 );
    or g24147 ( n34550 , n38051 , n39063 );
    and g24148 ( n36195 , n14573 , n18278 );
    nor g24149 ( n38264 , n34565 , n15500 );
    or g24150 ( n19028 , n37259 , n30863 );
    and g24151 ( n34344 , n2173 , n2471 );
    nor g24152 ( n13141 , n2183 , n30976 );
    not g24153 ( n7818 , n37051 );
    nor g24154 ( n36672 , n34566 , n32324 );
    or g24155 ( n3329 , n22836 , n40487 );
    not g24156 ( n23975 , n15043 );
    xnor g24157 ( n6667 , n9992 , n8273 );
    not g24158 ( n1867 , n13052 );
    xnor g24159 ( n13005 , n30415 , n8079 );
    and g24160 ( n8848 , n38796 , n10294 );
    and g24161 ( n33260 , n37001 , n26574 );
    or g24162 ( n16646 , n19525 , n34725 );
    not g24163 ( n26446 , n39742 );
    or g24164 ( n568 , n4117 , n28081 );
    or g24165 ( n2196 , n7534 , n33237 );
    nor g24166 ( n41441 , n13929 , n39588 );
    and g24167 ( n32044 , n12092 , n27944 );
    and g24168 ( n25851 , n21313 , n27948 );
    or g24169 ( n17310 , n37798 , n35267 );
    not g24170 ( n30550 , n5748 );
    or g24171 ( n6487 , n25474 , n18852 );
    or g24172 ( n16644 , n5795 , n38589 );
    and g24173 ( n673 , n16800 , n32383 );
    or g24174 ( n38400 , n8494 , n21665 );
    and g24175 ( n3922 , n4359 , n40262 );
    and g24176 ( n6949 , n18709 , n23905 );
    not g24177 ( n18920 , n33439 );
    or g24178 ( n10388 , n12881 , n28236 );
    nor g24179 ( n18591 , n16445 , n34279 );
    or g24180 ( n37024 , n24452 , n8658 );
    or g24181 ( n31065 , n6592 , n19842 );
    or g24182 ( n9251 , n22044 , n40101 );
    not g24183 ( n15727 , n11232 );
    nor g24184 ( n17695 , n13502 , n15019 );
    not g24185 ( n36295 , n15539 );
    or g24186 ( n38399 , n12924 , n62 );
    not g24187 ( n19594 , n19642 );
    not g24188 ( n8076 , n14194 );
    nor g24189 ( n19883 , n2963 , n17133 );
    nor g24190 ( n10143 , n37163 , n4992 );
    or g24191 ( n3852 , n10014 , n42079 );
    or g24192 ( n1056 , n2213 , n27616 );
    and g24193 ( n7728 , n19161 , n31092 );
    xnor g24194 ( n29184 , n39864 , n32419 );
    nor g24195 ( n21560 , n2411 , n9496 );
    and g24196 ( n14929 , n13219 , n10826 );
    not g24197 ( n2701 , n17327 );
    not g24198 ( n33624 , n12822 );
    and g24199 ( n4580 , n18117 , n10817 );
    not g24200 ( n23430 , n41236 );
    xnor g24201 ( n26425 , n31989 , n7079 );
    or g24202 ( n40211 , n7805 , n33450 );
    or g24203 ( n30244 , n2117 , n5921 );
    not g24204 ( n37465 , n32054 );
    xnor g24205 ( n39843 , n10076 , n24545 );
    or g24206 ( n6140 , n37638 , n33085 );
    or g24207 ( n19483 , n24468 , n18236 );
    not g24208 ( n14407 , n36488 );
    or g24209 ( n491 , n405 , n30362 );
    or g24210 ( n16156 , n12813 , n19173 );
    not g24211 ( n12998 , n4596 );
    or g24212 ( n19997 , n16586 , n38881 );
    or g24213 ( n10099 , n26192 , n3410 );
    and g24214 ( n27945 , n35957 , n40756 );
    not g24215 ( n17665 , n42353 );
    or g24216 ( n7778 , n37247 , n9075 );
    xnor g24217 ( n25795 , n18395 , n18877 );
    nor g24218 ( n7367 , n39356 , n34714 );
    not g24219 ( n41856 , n24273 );
    not g24220 ( n29949 , n31519 );
    or g24221 ( n27000 , n27329 , n7955 );
    and g24222 ( n30470 , n6749 , n3872 );
    not g24223 ( n28979 , n35307 );
    nor g24224 ( n33265 , n32069 , n27037 );
    nor g24225 ( n36782 , n12248 , n37374 );
    xnor g24226 ( n32246 , n34364 , n23927 );
    xnor g24227 ( n26393 , n17019 , n29737 );
    and g24228 ( n1502 , n36648 , n33759 );
    not g24229 ( n9588 , n8066 );
    or g24230 ( n2946 , n4213 , n1289 );
    or g24231 ( n3127 , n36405 , n11746 );
    not g24232 ( n9619 , n40225 );
    nor g24233 ( n29655 , n21762 , n15386 );
    or g24234 ( n11671 , n13419 , n39626 );
    xnor g24235 ( n4260 , n33570 , n2876 );
    or g24236 ( n40436 , n12325 , n14503 );
    and g24237 ( n10111 , n25306 , n20643 );
    or g24238 ( n5626 , n216 , n2647 );
    or g24239 ( n25106 , n4195 , n16220 );
    and g24240 ( n28892 , n41111 , n32186 );
    or g24241 ( n40892 , n11492 , n17923 );
    or g24242 ( n10463 , n26915 , n788 );
    xnor g24243 ( n24008 , n4879 , n12574 );
    or g24244 ( n42028 , n38897 , n37250 );
    xnor g24245 ( n8228 , n33757 , n23486 );
    or g24246 ( n1047 , n33981 , n21545 );
    or g24247 ( n17740 , n38211 , n37737 );
    or g24248 ( n3461 , n35283 , n26495 );
    xnor g24249 ( n32165 , n14758 , n41471 );
    nor g24250 ( n40207 , n13228 , n2257 );
    or g24251 ( n31462 , n38165 , n13826 );
    not g24252 ( n15527 , n34813 );
    or g24253 ( n1590 , n22167 , n37118 );
    or g24254 ( n3620 , n32752 , n12350 );
    and g24255 ( n8322 , n2147 , n3207 );
    or g24256 ( n6404 , n1980 , n15540 );
    not g24257 ( n3396 , n3003 );
    or g24258 ( n8140 , n7356 , n24606 );
    xnor g24259 ( n3430 , n34731 , n1070 );
    or g24260 ( n10328 , n42722 , n30266 );
    and g24261 ( n25986 , n37714 , n13136 );
    not g24262 ( n931 , n6338 );
    or g24263 ( n35135 , n3981 , n18025 );
    and g24264 ( n15525 , n25242 , n6488 );
    or g24265 ( n6099 , n1139 , n21172 );
    and g24266 ( n20750 , n39340 , n36194 );
    or g24267 ( n11430 , n38863 , n8328 );
    nor g24268 ( n42255 , n365 , n3604 );
    xnor g24269 ( n30625 , n17413 , n31504 );
    xnor g24270 ( n30141 , n24258 , n12032 );
    xnor g24271 ( n4773 , n11819 , n34737 );
    not g24272 ( n17314 , n16445 );
    and g24273 ( n26752 , n36709 , n19453 );
    or g24274 ( n38300 , n12786 , n9205 );
    not g24275 ( n37520 , n14224 );
    not g24276 ( n15441 , n35104 );
    nor g24277 ( n8050 , n41662 , n4132 );
    nor g24278 ( n38025 , n40581 , n31767 );
    not g24279 ( n13415 , n24800 );
    or g24280 ( n1887 , n24222 , n28141 );
    nor g24281 ( n26158 , n29113 , n5628 );
    and g24282 ( n25271 , n11334 , n24332 );
    and g24283 ( n33439 , n31183 , n29090 );
    or g24284 ( n33690 , n17204 , n8742 );
    or g24285 ( n38631 , n39810 , n33113 );
    or g24286 ( n8753 , n3248 , n7219 );
    xnor g24287 ( n27011 , n29667 , n37901 );
    xnor g24288 ( n41391 , n5144 , n33010 );
    or g24289 ( n19381 , n35505 , n37660 );
    not g24290 ( n8880 , n38331 );
    and g24291 ( n22009 , n25415 , n21780 );
    or g24292 ( n1213 , n30581 , n24098 );
    nor g24293 ( n39024 , n2199 , n4599 );
    and g24294 ( n35990 , n25760 , n2926 );
    or g24295 ( n4395 , n21752 , n2354 );
    or g24296 ( n25532 , n2692 , n22216 );
    not g24297 ( n3051 , n31183 );
    and g24298 ( n31747 , n32617 , n13442 );
    or g24299 ( n7424 , n7637 , n12402 );
    or g24300 ( n4152 , n29027 , n39794 );
    and g24301 ( n729 , n13218 , n11366 );
    and g24302 ( n7427 , n39013 , n16584 );
    or g24303 ( n1147 , n21817 , n4669 );
    or g24304 ( n23293 , n11928 , n36050 );
    not g24305 ( n26613 , n42707 );
    not g24306 ( n34031 , n32804 );
    nor g24307 ( n1357 , n16257 , n38362 );
    nor g24308 ( n29985 , n2183 , n25928 );
    or g24309 ( n16919 , n33869 , n31321 );
    or g24310 ( n10338 , n16198 , n20147 );
    or g24311 ( n10973 , n30010 , n30263 );
    or g24312 ( n16206 , n1980 , n23523 );
    not g24313 ( n23940 , n24590 );
    or g24314 ( n36175 , n2199 , n39286 );
    not g24315 ( n39287 , n5819 );
    or g24316 ( n7553 , n3583 , n13669 );
    not g24317 ( n25528 , n17301 );
    or g24318 ( n6366 , n15619 , n29464 );
    or g24319 ( n5031 , n10829 , n42786 );
    xnor g24320 ( n17157 , n22296 , n8803 );
    or g24321 ( n33300 , n31924 , n42614 );
    nor g24322 ( n4531 , n10939 , n22744 );
    not g24323 ( n37051 , n34076 );
    nor g24324 ( n24719 , n1448 , n31027 );
    and g24325 ( n31405 , n31565 , n40856 );
    and g24326 ( n19836 , n19752 , n17099 );
    or g24327 ( n34834 , n1505 , n41891 );
    and g24328 ( n25072 , n5563 , n35634 );
    not g24329 ( n41428 , n13420 );
    not g24330 ( n19925 , n9146 );
    or g24331 ( n42741 , n10099 , n27060 );
    and g24332 ( n31075 , n26036 , n2133 );
    or g24333 ( n11123 , n6748 , n32688 );
    nor g24334 ( n33698 , n30736 , n42119 );
    not g24335 ( n36911 , n6483 );
    not g24336 ( n11708 , n18317 );
    or g24337 ( n23091 , n10350 , n3856 );
    not g24338 ( n20804 , n20980 );
    and g24339 ( n22118 , n39059 , n25140 );
    or g24340 ( n15263 , n40874 , n6079 );
    xnor g24341 ( n39704 , n24411 , n10430 );
    not g24342 ( n11986 , n35230 );
    not g24343 ( n25279 , n18510 );
    and g24344 ( n19614 , n6468 , n20998 );
    and g24345 ( n14761 , n25489 , n27475 );
    not g24346 ( n28149 , n28968 );
    not g24347 ( n2855 , n11511 );
    and g24348 ( n10624 , n6800 , n31611 );
    xnor g24349 ( n10989 , n26794 , n21655 );
    nor g24350 ( n33366 , n28884 , n9724 );
    or g24351 ( n40361 , n15149 , n32552 );
    and g24352 ( n8561 , n7744 , n1413 );
    nor g24353 ( n17535 , n30295 , n36802 );
    nor g24354 ( n31150 , n6799 , n30534 );
    nor g24355 ( n19265 , n1507 , n26946 );
    not g24356 ( n27513 , n12638 );
    or g24357 ( n25422 , n3235 , n10045 );
    or g24358 ( n38982 , n41011 , n15186 );
    or g24359 ( n1992 , n31858 , n28461 );
    not g24360 ( n36723 , n37041 );
    nor g24361 ( n36713 , n14475 , n34594 );
    nor g24362 ( n41602 , n25477 , n1612 );
    or g24363 ( n2580 , n28348 , n29299 );
    or g24364 ( n36623 , n6218 , n10332 );
    and g24365 ( n26250 , n15024 , n15949 );
    or g24366 ( n30564 , n19969 , n35213 );
    or g24367 ( n41946 , n1546 , n15803 );
    or g24368 ( n26320 , n7577 , n32619 );
    nor g24369 ( n7985 , n2603 , n20937 );
    not g24370 ( n41424 , n10162 );
    or g24371 ( n34996 , n3695 , n36839 );
    not g24372 ( n34844 , n6442 );
    not g24373 ( n30192 , n10867 );
    and g24374 ( n23946 , n36358 , n21801 );
    or g24375 ( n32482 , n34687 , n37427 );
    or g24376 ( n39092 , n22091 , n25938 );
    nor g24377 ( n17017 , n35590 , n34159 );
    or g24378 ( n6875 , n14491 , n36880 );
    xnor g24379 ( n2551 , n26475 , n38665 );
    or g24380 ( n34645 , n11389 , n17827 );
    and g24381 ( n3818 , n7770 , n359 );
    and g24382 ( n33318 , n40590 , n9139 );
    not g24383 ( n6032 , n11264 );
    and g24384 ( n39746 , n2933 , n22012 );
    and g24385 ( n41784 , n19006 , n38987 );
    or g24386 ( n29372 , n28700 , n439 );
    not g24387 ( n5188 , n2483 );
    or g24388 ( n27470 , n23557 , n27395 );
    nor g24389 ( n37118 , n36667 , n41226 );
    and g24390 ( n39694 , n38471 , n24540 );
    nor g24391 ( n83 , n8494 , n26585 );
    and g24392 ( n14267 , n621 , n19998 );
    nor g24393 ( n42809 , n36547 , n9596 );
    or g24394 ( n32240 , n38879 , n28079 );
    or g24395 ( n15029 , n25453 , n33671 );
    and g24396 ( n38967 , n32865 , n29204 );
    xnor g24397 ( n20044 , n28458 , n10690 );
    nor g24398 ( n29108 , n8787 , n38507 );
    or g24399 ( n28806 , n14501 , n6413 );
    or g24400 ( n42772 , n4374 , n13701 );
    or g24401 ( n20693 , n22428 , n38924 );
    not g24402 ( n12695 , n36767 );
    not g24403 ( n26961 , n5947 );
    or g24404 ( n24462 , n24513 , n25277 );
    or g24405 ( n10407 , n24496 , n17924 );
    not g24406 ( n42058 , n14803 );
    and g24407 ( n35192 , n31181 , n27244 );
    or g24408 ( n35171 , n19437 , n37952 );
    not g24409 ( n12212 , n11903 );
    or g24410 ( n18966 , n23444 , n19918 );
    and g24411 ( n12319 , n27289 , n39763 );
    nor g24412 ( n41829 , n24115 , n17611 );
    and g24413 ( n22757 , n29468 , n531 );
    not g24414 ( n4305 , n9492 );
    or g24415 ( n32310 , n2697 , n16530 );
    xnor g24416 ( n17625 , n40886 , n28847 );
    or g24417 ( n29505 , n301 , n34061 );
    and g24418 ( n1870 , n40117 , n1915 );
    nor g24419 ( n28364 , n35041 , n7481 );
    or g24420 ( n35812 , n178 , n32614 );
    or g24421 ( n37551 , n32309 , n10921 );
    not g24422 ( n25738 , n13054 );
    and g24423 ( n41799 , n13069 , n3808 );
    or g24424 ( n20782 , n23292 , n35275 );
    or g24425 ( n15486 , n15621 , n4997 );
    and g24426 ( n1082 , n4537 , n25045 );
    nor g24427 ( n32109 , n18233 , n11817 );
    or g24428 ( n29768 , n39618 , n30592 );
    not g24429 ( n20288 , n19832 );
    not g24430 ( n3549 , n9331 );
    or g24431 ( n1504 , n32495 , n36024 );
    or g24432 ( n19277 , n34796 , n41485 );
    or g24433 ( n767 , n28745 , n25523 );
    or g24434 ( n33536 , n15477 , n8615 );
    and g24435 ( n41762 , n39465 , n14339 );
    nor g24436 ( n18715 , n24202 , n8485 );
    nor g24437 ( n5506 , n15100 , n15311 );
    not g24438 ( n36939 , n19248 );
    or g24439 ( n39793 , n40671 , n40514 );
    or g24440 ( n41196 , n763 , n5589 );
    and g24441 ( n31741 , n33574 , n1112 );
    not g24442 ( n40554 , n231 );
    not g24443 ( n28029 , n14782 );
    and g24444 ( n27824 , n15252 , n20471 );
    and g24445 ( n23897 , n42869 , n10370 );
    nor g24446 ( n9566 , n1971 , n11192 );
    xnor g24447 ( n34197 , n36677 , n31612 );
    not g24448 ( n29059 , n29588 );
    not g24449 ( n1499 , n18247 );
    or g24450 ( n33928 , n19523 , n12914 );
    xnor g24451 ( n25265 , n41293 , n10561 );
    or g24452 ( n4981 , n13374 , n6456 );
    or g24453 ( n7932 , n38733 , n24844 );
    or g24454 ( n2578 , n8621 , n1808 );
    and g24455 ( n34133 , n31042 , n1976 );
    nor g24456 ( n28452 , n12054 , n5091 );
    or g24457 ( n25244 , n34221 , n22716 );
    not g24458 ( n41457 , n5646 );
    and g24459 ( n16491 , n16147 , n16434 );
    not g24460 ( n30558 , n37559 );
    nor g24461 ( n32210 , n19054 , n22528 );
    and g24462 ( n15757 , n18307 , n9810 );
    nor g24463 ( n2738 , n17744 , n25537 );
    or g24464 ( n34747 , n36826 , n19352 );
    xnor g24465 ( n7924 , n2501 , n13598 );
    or g24466 ( n39124 , n27915 , n9256 );
    nor g24467 ( n17526 , n39266 , n23423 );
    and g24468 ( n2662 , n3826 , n5354 );
    or g24469 ( n596 , n28615 , n42507 );
    or g24470 ( n26770 , n25460 , n17404 );
    or g24471 ( n30643 , n30307 , n23211 );
    or g24472 ( n24005 , n8281 , n13560 );
    or g24473 ( n36448 , n36344 , n7569 );
    and g24474 ( n25785 , n38827 , n16568 );
    not g24475 ( n24691 , n21366 );
    or g24476 ( n13230 , n14161 , n3057 );
    or g24477 ( n31151 , n21283 , n17229 );
    and g24478 ( n27383 , n35648 , n2805 );
    nor g24479 ( n42826 , n32813 , n13847 );
    nor g24480 ( n27065 , n28965 , n4011 );
    and g24481 ( n32825 , n26583 , n1684 );
    or g24482 ( n29425 , n33328 , n29378 );
    or g24483 ( n41106 , n31106 , n27957 );
    or g24484 ( n39465 , n2929 , n41752 );
    xnor g24485 ( n4914 , n41013 , n38845 );
    or g24486 ( n15847 , n11326 , n40445 );
    or g24487 ( n25805 , n1756 , n17529 );
    not g24488 ( n26681 , n26142 );
    or g24489 ( n10580 , n12355 , n24925 );
    xnor g24490 ( n1485 , n28313 , n34217 );
    or g24491 ( n41845 , n41853 , n19769 );
    not g24492 ( n23838 , n26078 );
    nor g24493 ( n29938 , n3574 , n17613 );
    and g24494 ( n14114 , n24460 , n25868 );
    and g24495 ( n19283 , n6360 , n31532 );
    or g24496 ( n31793 , n40512 , n25133 );
    or g24497 ( n6569 , n29344 , n22333 );
    or g24498 ( n26395 , n30708 , n30496 );
    or g24499 ( n28305 , n8778 , n41981 );
    or g24500 ( n25819 , n34609 , n11643 );
    or g24501 ( n39034 , n3815 , n7740 );
    and g24502 ( n24902 , n42724 , n27639 );
    xnor g24503 ( n28255 , n4218 , n2601 );
    or g24504 ( n37354 , n1971 , n33619 );
    or g24505 ( n34784 , n38824 , n15095 );
    or g24506 ( n23124 , n29613 , n27611 );
    or g24507 ( n34770 , n2199 , n18055 );
    and g24508 ( n2493 , n27894 , n15812 );
    not g24509 ( n34091 , n41578 );
    or g24510 ( n4863 , n34241 , n33671 );
    or g24511 ( n37390 , n24441 , n11320 );
    not g24512 ( n15040 , n21918 );
    nor g24513 ( n37857 , n9499 , n33498 );
    or g24514 ( n28761 , n41218 , n35118 );
    or g24515 ( n19881 , n20721 , n19540 );
    and g24516 ( n31277 , n14978 , n11684 );
    nor g24517 ( n11582 , n29640 , n2009 );
    not g24518 ( n23323 , n7779 );
    or g24519 ( n8918 , n21397 , n40419 );
    or g24520 ( n12254 , n37179 , n21636 );
    nor g24521 ( n26431 , n14707 , n34670 );
    not g24522 ( n15176 , n30306 );
    or g24523 ( n8889 , n23921 , n12631 );
    not g24524 ( n29731 , n34076 );
    and g24525 ( n2439 , n25912 , n32629 );
    or g24526 ( n12240 , n14675 , n33540 );
    or g24527 ( n37071 , n8496 , n19950 );
    or g24528 ( n524 , n16682 , n42253 );
    and g24529 ( n42875 , n26642 , n23672 );
    or g24530 ( n3295 , n19362 , n34017 );
    and g24531 ( n171 , n32277 , n27074 );
    or g24532 ( n26370 , n31696 , n12051 );
    or g24533 ( n17543 , n36821 , n31601 );
    xnor g24534 ( n23087 , n1798 , n27883 );
    not g24535 ( n29579 , n25233 );
    or g24536 ( n12320 , n15149 , n28386 );
    or g24537 ( n1031 , n20686 , n38691 );
    and g24538 ( n34117 , n31330 , n3822 );
    or g24539 ( n36903 , n9430 , n5463 );
    or g24540 ( n29976 , n21235 , n42377 );
    or g24541 ( n17074 , n19691 , n32676 );
    and g24542 ( n32024 , n32537 , n26400 );
    or g24543 ( n33534 , n11404 , n14761 );
    not g24544 ( n41400 , n21968 );
    and g24545 ( n32478 , n29088 , n11104 );
    and g24546 ( n12580 , n18530 , n26274 );
    or g24547 ( n886 , n13176 , n25943 );
    or g24548 ( n6235 , n21553 , n23570 );
    xnor g24549 ( n11692 , n4302 , n40660 );
    and g24550 ( n38800 , n35771 , n14269 );
    nor g24551 ( n3055 , n4561 , n11808 );
    or g24552 ( n28558 , n29276 , n42671 );
    or g24553 ( n35565 , n4790 , n20881 );
    xnor g24554 ( n19878 , n6625 , n13599 );
    not g24555 ( n30862 , n32938 );
    not g24556 ( n22699 , n32165 );
    and g24557 ( n25847 , n9507 , n37192 );
    not g24558 ( n6767 , n5842 );
    not g24559 ( n37839 , n31364 );
    xnor g24560 ( n23827 , n20811 , n27392 );
    or g24561 ( n28274 , n18314 , n18838 );
    or g24562 ( n32507 , n39968 , n8172 );
    or g24563 ( n28939 , n15070 , n14260 );
    and g24564 ( n9807 , n24536 , n6849 );
    not g24565 ( n1752 , n19181 );
    not g24566 ( n33375 , n37872 );
    not g24567 ( n2205 , n15693 );
    or g24568 ( n13217 , n26565 , n40186 );
    or g24569 ( n5363 , n24656 , n24848 );
    or g24570 ( n37194 , n10346 , n22800 );
    xnor g24571 ( n36816 , n32534 , n37439 );
    nor g24572 ( n16363 , n17909 , n38492 );
    and g24573 ( n11255 , n18232 , n10280 );
    and g24574 ( n29584 , n6707 , n32987 );
    or g24575 ( n9497 , n38205 , n33766 );
    not g24576 ( n11168 , n37873 );
    nor g24577 ( n11778 , n27733 , n18349 );
    not g24578 ( n27598 , n24000 );
    and g24579 ( n21280 , n37987 , n5967 );
    not g24580 ( n23386 , n17195 );
    or g24581 ( n34452 , n13332 , n40390 );
    xnor g24582 ( n14631 , n28443 , n14623 );
    and g24583 ( n493 , n30337 , n13159 );
    xnor g24584 ( n6116 , n9180 , n33940 );
    or g24585 ( n22150 , n5706 , n17230 );
    xnor g24586 ( n18854 , n5144 , n32411 );
    or g24587 ( n11909 , n33691 , n36116 );
    nor g24588 ( n26403 , n311 , n26912 );
    or g24589 ( n22087 , n25839 , n19062 );
    or g24590 ( n21384 , n19460 , n41649 );
    or g24591 ( n32592 , n23341 , n12772 );
    nor g24592 ( n29648 , n4308 , n5879 );
    or g24593 ( n6485 , n34781 , n18491 );
    or g24594 ( n5635 , n7616 , n13846 );
    xnor g24595 ( n1855 , n71 , n33029 );
    or g24596 ( n985 , n6881 , n33330 );
    or g24597 ( n18760 , n8708 , n6510 );
    not g24598 ( n25402 , n32072 );
    or g24599 ( n22951 , n4816 , n9417 );
    or g24600 ( n6522 , n37707 , n29162 );
    or g24601 ( n26660 , n8470 , n31277 );
    or g24602 ( n41005 , n3602 , n33265 );
    or g24603 ( n13592 , n18314 , n27492 );
    and g24604 ( n12284 , n18957 , n374 );
    not g24605 ( n36148 , n21502 );
    or g24606 ( n21757 , n20932 , n20999 );
    or g24607 ( n40496 , n3010 , n13590 );
    nor g24608 ( n16100 , n12222 , n7972 );
    not g24609 ( n22128 , n40372 );
    not g24610 ( n34436 , n31184 );
    or g24611 ( n29321 , n25317 , n13198 );
    nor g24612 ( n35213 , n15626 , n39514 );
    xnor g24613 ( n41916 , n9630 , n32522 );
    xnor g24614 ( n30220 , n22263 , n11821 );
    and g24615 ( n18349 , n7983 , n16762 );
    xnor g24616 ( n37181 , n5399 , n25595 );
    and g24617 ( n40475 , n34582 , n28054 );
    xnor g24618 ( n9388 , n16105 , n25455 );
    or g24619 ( n12052 , n3443 , n35556 );
    or g24620 ( n14320 , n30896 , n41438 );
    nor g24621 ( n21501 , n34379 , n34541 );
    nor g24622 ( n42007 , n19519 , n572 );
    and g24623 ( n1825 , n23401 , n27038 );
    not g24624 ( n39722 , n26650 );
    and g24625 ( n37809 , n1748 , n29944 );
    and g24626 ( n26369 , n32672 , n27946 );
    or g24627 ( n17156 , n30579 , n42817 );
    or g24628 ( n34147 , n27355 , n23926 );
    or g24629 ( n1846 , n24052 , n32892 );
    not g24630 ( n42003 , n8759 );
    not g24631 ( n14377 , n41992 );
    or g24632 ( n19799 , n24328 , n34187 );
    or g24633 ( n39103 , n11814 , n6252 );
    or g24634 ( n23190 , n3764 , n42815 );
    or g24635 ( n16064 , n29455 , n39306 );
    or g24636 ( n27838 , n19762 , n15448 );
    not g24637 ( n29476 , n40173 );
    and g24638 ( n38874 , n30520 , n20768 );
    or g24639 ( n42230 , n4666 , n4669 );
    or g24640 ( n27317 , n11050 , n42305 );
    or g24641 ( n8519 , n17827 , n5199 );
    or g24642 ( n12211 , n17794 , n740 );
    not g24643 ( n20982 , n25899 );
    nor g24644 ( n28874 , n25619 , n18894 );
    nor g24645 ( n17059 , n5896 , n16426 );
    not g24646 ( n31286 , n3490 );
    and g24647 ( n41026 , n20641 , n2141 );
    and g24648 ( n5248 , n297 , n29196 );
    xnor g24649 ( n5237 , n34945 , n26820 );
    xnor g24650 ( n26012 , n1664 , n11749 );
    or g24651 ( n23967 , n31121 , n19701 );
    or g24652 ( n17711 , n34674 , n1375 );
    not g24653 ( n10848 , n25899 );
    and g24654 ( n31458 , n4890 , n4831 );
    not g24655 ( n7654 , n9223 );
    or g24656 ( n17246 , n9817 , n3796 );
    or g24657 ( n36854 , n25617 , n37500 );
    and g24658 ( n21805 , n39801 , n4867 );
    or g24659 ( n3360 , n345 , n30437 );
    or g24660 ( n7890 , n29038 , n17994 );
    and g24661 ( n32733 , n9992 , n8273 );
    xnor g24662 ( n33014 , n8225 , n6594 );
    or g24663 ( n32924 , n36332 , n19041 );
    not g24664 ( n22523 , n32593 );
    and g24665 ( n21378 , n31985 , n5093 );
    not g24666 ( n19153 , n2539 );
    or g24667 ( n13088 , n24453 , n40885 );
    or g24668 ( n33989 , n35534 , n19747 );
    nor g24669 ( n14558 , n39903 , n16094 );
    or g24670 ( n7676 , n6132 , n30241 );
    nor g24671 ( n6295 , n13657 , n29067 );
    and g24672 ( n6872 , n23660 , n38803 );
    and g24673 ( n37253 , n37531 , n22406 );
    not g24674 ( n228 , n42554 );
    or g24675 ( n13424 , n37636 , n14526 );
    and g24676 ( n35309 , n6144 , n28284 );
    not g24677 ( n34732 , n41741 );
    or g24678 ( n30495 , n33981 , n642 );
    nor g24679 ( n35049 , n14194 , n20795 );
    not g24680 ( n39624 , n10635 );
    xnor g24681 ( n10214 , n20067 , n4933 );
    or g24682 ( n17168 , n21417 , n19698 );
    and g24683 ( n41318 , n7713 , n25767 );
    nor g24684 ( n28322 , n35924 , n41917 );
    or g24685 ( n12289 , n36597 , n29856 );
    or g24686 ( n11872 , n37549 , n16682 );
    not g24687 ( n21245 , n25918 );
    or g24688 ( n26080 , n25547 , n28722 );
    or g24689 ( n32872 , n9456 , n2538 );
    or g24690 ( n16283 , n37808 , n33487 );
    or g24691 ( n29573 , n2608 , n19806 );
    not g24692 ( n39239 , n41905 );
    not g24693 ( n6861 , n29163 );
    and g24694 ( n7603 , n42256 , n10743 );
    or g24695 ( n9059 , n14341 , n32194 );
    xnor g24696 ( n12394 , n21415 , n41461 );
    nor g24697 ( n37007 , n2962 , n381 );
    or g24698 ( n32057 , n2076 , n32020 );
    not g24699 ( n38444 , n41457 );
    nor g24700 ( n16831 , n25242 , n6488 );
    xnor g24701 ( n39106 , n14246 , n28966 );
    or g24702 ( n25688 , n20510 , n22551 );
    or g24703 ( n693 , n34678 , n16978 );
    not g24704 ( n13042 , n12367 );
    or g24705 ( n17060 , n9031 , n11090 );
    or g24706 ( n2590 , n8441 , n14354 );
    xnor g24707 ( n42890 , n105 , n41928 );
    or g24708 ( n663 , n14700 , n31503 );
    or g24709 ( n27509 , n24243 , n13926 );
    and g24710 ( n42769 , n9638 , n37324 );
    xnor g24711 ( n9037 , n5041 , n2198 );
    nor g24712 ( n37271 , n15413 , n28376 );
    or g24713 ( n10309 , n31422 , n8561 );
    or g24714 ( n11400 , n33815 , n13568 );
    or g24715 ( n7658 , n26367 , n33638 );
    nor g24716 ( n11573 , n33706 , n24195 );
    not g24717 ( n23964 , n10748 );
    nor g24718 ( n15577 , n14707 , n30799 );
    and g24719 ( n27180 , n85 , n29838 );
    or g24720 ( n23375 , n396 , n12392 );
    and g24721 ( n21187 , n25421 , n6443 );
    xnor g24722 ( n35771 , n16693 , n29533 );
    and g24723 ( n4121 , n10509 , n15598 );
    not g24724 ( n13690 , n41081 );
    not g24725 ( n37896 , n101 );
    and g24726 ( n19209 , n1901 , n6513 );
    and g24727 ( n6082 , n31358 , n27547 );
    xnor g24728 ( n9208 , n26428 , n5970 );
    or g24729 ( n250 , n19469 , n23841 );
    and g24730 ( n28750 , n24361 , n18721 );
    or g24731 ( n13328 , n37479 , n10136 );
    or g24732 ( n33994 , n29134 , n13368 );
    nor g24733 ( n14641 , n9448 , n39984 );
    not g24734 ( n8793 , n20971 );
    or g24735 ( n24557 , n39442 , n31590 );
    xnor g24736 ( n7717 , n31099 , n38510 );
    or g24737 ( n15270 , n42270 , n3781 );
    and g24738 ( n41344 , n38717 , n9120 );
    xnor g24739 ( n2809 , n5797 , n38972 );
    or g24740 ( n23312 , n28647 , n35149 );
    not g24741 ( n119 , n34030 );
    not g24742 ( n30398 , n4716 );
    or g24743 ( n31172 , n25516 , n36224 );
    xnor g24744 ( n2944 , n29740 , n36883 );
    xnor g24745 ( n13029 , n12007 , n17367 );
    or g24746 ( n23055 , n7222 , n26828 );
    or g24747 ( n22005 , n42439 , n2517 );
    not g24748 ( n36941 , n7155 );
    or g24749 ( n1655 , n23235 , n39252 );
    and g24750 ( n31902 , n11997 , n8855 );
    and g24751 ( n5894 , n26844 , n25244 );
    or g24752 ( n40749 , n14935 , n31575 );
    or g24753 ( n12116 , n15461 , n36940 );
    or g24754 ( n6149 , n2151 , n27060 );
    and g24755 ( n40286 , n28304 , n20298 );
    not g24756 ( n30674 , n21561 );
    and g24757 ( n22987 , n19500 , n6108 );
    and g24758 ( n7635 , n41495 , n9345 );
    xnor g24759 ( n22580 , n5144 , n18273 );
    nor g24760 ( n29791 , n20797 , n7807 );
    or g24761 ( n14150 , n37664 , n8593 );
    or g24762 ( n16000 , n11265 , n5407 );
    or g24763 ( n28227 , n15585 , n35210 );
    and g24764 ( n12956 , n20307 , n6329 );
    or g24765 ( n38866 , n40699 , n40775 );
    xnor g24766 ( n1127 , n27342 , n15844 );
    not g24767 ( n3636 , n4331 );
    or g24768 ( n24184 , n32800 , n21671 );
    not g24769 ( n8539 , n41253 );
    xnor g24770 ( n23918 , n31989 , n12121 );
    or g24771 ( n1498 , n31452 , n27880 );
    and g24772 ( n20032 , n8648 , n8055 );
    not g24773 ( n6454 , n10749 );
    and g24774 ( n34636 , n25226 , n37895 );
    or g24775 ( n15840 , n26792 , n5193 );
    not g24776 ( n20163 , n1929 );
    or g24777 ( n27525 , n2380 , n36687 );
    and g24778 ( n24530 , n9822 , n35668 );
    and g24779 ( n38786 , n15520 , n35630 );
    nor g24780 ( n20077 , n17744 , n41132 );
    and g24781 ( n31781 , n38178 , n3938 );
    or g24782 ( n15756 , n41484 , n33435 );
    or g24783 ( n16977 , n9189 , n42561 );
    or g24784 ( n9717 , n23971 , n40055 );
    or g24785 ( n31243 , n27920 , n1106 );
    or g24786 ( n24552 , n17563 , n16578 );
    or g24787 ( n24465 , n33433 , n21805 );
    and g24788 ( n1468 , n39743 , n30486 );
    or g24789 ( n11179 , n27920 , n2319 );
    or g24790 ( n16061 , n29112 , n19561 );
    nor g24791 ( n13276 , n11703 , n19730 );
    nor g24792 ( n33696 , n5786 , n7459 );
    nor g24793 ( n3974 , n38563 , n40838 );
    and g24794 ( n34326 , n29245 , n33578 );
    and g24795 ( n10694 , n35703 , n42230 );
    and g24796 ( n477 , n12834 , n33097 );
    or g24797 ( n3858 , n1499 , n10603 );
    xnor g24798 ( n33303 , n5891 , n15370 );
    nor g24799 ( n27021 , n13174 , n22145 );
    not g24800 ( n37280 , n8947 );
    not g24801 ( n25671 , n42817 );
    and g24802 ( n34669 , n35181 , n31891 );
    or g24803 ( n33914 , n6893 , n22164 );
    xnor g24804 ( n14538 , n27874 , n3256 );
    and g24805 ( n8465 , n38182 , n15028 );
    nor g24806 ( n11415 , n27780 , n28591 );
    and g24807 ( n14905 , n42355 , n21233 );
    or g24808 ( n6056 , n28143 , n12002 );
    not g24809 ( n22137 , n39161 );
    and g24810 ( n31839 , n35727 , n29878 );
    or g24811 ( n1027 , n25973 , n7242 );
    or g24812 ( n38422 , n7307 , n38266 );
    and g24813 ( n13348 , n28328 , n1899 );
    not g24814 ( n41498 , n14196 );
    nor g24815 ( n4489 , n4330 , n36990 );
    or g24816 ( n12585 , n33972 , n9914 );
    xnor g24817 ( n30505 , n11145 , n10793 );
    xnor g24818 ( n39957 , n15524 , n2113 );
    nor g24819 ( n20317 , n13546 , n4134 );
    not g24820 ( n14052 , n24856 );
    nor g24821 ( n23858 , n39264 , n17819 );
    or g24822 ( n22510 , n40867 , n33186 );
    or g24823 ( n4645 , n5183 , n1865 );
    or g24824 ( n12202 , n19221 , n18677 );
    not g24825 ( n42327 , n42674 );
    xnor g24826 ( n26121 , n11799 , n10009 );
    not g24827 ( n1793 , n9874 );
    and g24828 ( n1390 , n12798 , n20858 );
    and g24829 ( n38588 , n33086 , n22698 );
    and g24830 ( n34896 , n40046 , n3830 );
    or g24831 ( n39054 , n42706 , n31773 );
    or g24832 ( n35602 , n13745 , n12169 );
    and g24833 ( n42290 , n41773 , n17090 );
    or g24834 ( n31411 , n23505 , n41934 );
    or g24835 ( n35589 , n27786 , n4241 );
    xnor g24836 ( n16752 , n3835 , n26588 );
    or g24837 ( n7238 , n17424 , n7795 );
    and g24838 ( n8173 , n5724 , n26243 );
    and g24839 ( n27015 , n9289 , n33319 );
    or g24840 ( n13082 , n11319 , n37730 );
    or g24841 ( n34872 , n6666 , n13417 );
    or g24842 ( n6890 , n42535 , n32509 );
    xnor g24843 ( n19495 , n14649 , n9514 );
    not g24844 ( n10833 , n17567 );
    not g24845 ( n35089 , n9147 );
    and g24846 ( n35495 , n39938 , n14662 );
    or g24847 ( n17917 , n33712 , n35755 );
    or g24848 ( n9822 , n38556 , n20369 );
    not g24849 ( n17804 , n29416 );
    or g24850 ( n42872 , n6671 , n9341 );
    or g24851 ( n19650 , n38998 , n15780 );
    xnor g24852 ( n16411 , n28083 , n21341 );
    nor g24853 ( n30482 , n30818 , n7 );
    not g24854 ( n2959 , n25403 );
    nor g24855 ( n12594 , n23934 , n14759 );
    and g24856 ( n21583 , n32810 , n32420 );
    not g24857 ( n16764 , n27576 );
    nor g24858 ( n14956 , n17659 , n1925 );
    and g24859 ( n9503 , n5104 , n36165 );
    and g24860 ( n18376 , n23275 , n27763 );
    or g24861 ( n16994 , n17313 , n22361 );
    or g24862 ( n40078 , n39929 , n42160 );
    or g24863 ( n689 , n5348 , n16426 );
    and g24864 ( n7835 , n24339 , n20753 );
    or g24865 ( n33605 , n15384 , n23888 );
    not g24866 ( n38640 , n2060 );
    and g24867 ( n980 , n9476 , n36289 );
    xnor g24868 ( n34980 , n450 , n7636 );
    and g24869 ( n31991 , n28271 , n9136 );
    nor g24870 ( n18975 , n2199 , n9749 );
    and g24871 ( n15292 , n37452 , n21168 );
    and g24872 ( n3794 , n24945 , n6735 );
    or g24873 ( n17617 , n24599 , n35207 );
    or g24874 ( n3555 , n39030 , n28241 );
    and g24875 ( n10433 , n27662 , n24280 );
    or g24876 ( n14582 , n24626 , n1064 );
    nor g24877 ( n37768 , n32042 , n37353 );
    nor g24878 ( n22439 , n10209 , n25065 );
    or g24879 ( n2352 , n41566 , n38142 );
    not g24880 ( n15926 , n36944 );
    and g24881 ( n314 , n28321 , n39067 );
    or g24882 ( n16535 , n29610 , n25838 );
    and g24883 ( n17548 , n938 , n9746 );
    xnor g24884 ( n24878 , n35329 , n10746 );
    nor g24885 ( n4856 , n41325 , n39693 );
    not g24886 ( n20799 , n4137 );
    not g24887 ( n22920 , n40954 );
    or g24888 ( n23831 , n18544 , n9621 );
    xnor g24889 ( n8922 , n34226 , n855 );
    xnor g24890 ( n15191 , n39544 , n1043 );
    xnor g24891 ( n27657 , n18192 , n18441 );
    not g24892 ( n3837 , n25893 );
    or g24893 ( n10507 , n25485 , n37250 );
    not g24894 ( n11432 , n6067 );
    or g24895 ( n38137 , n31165 , n37808 );
    or g24896 ( n12779 , n9319 , n12421 );
    and g24897 ( n11806 , n4520 , n8 );
    or g24898 ( n19130 , n10528 , n27385 );
    nor g24899 ( n2657 , n6774 , n40102 );
    not g24900 ( n37055 , n22125 );
    not g24901 ( n8255 , n23681 );
    nor g24902 ( n26505 , n13139 , n6336 );
    or g24903 ( n2760 , n26116 , n12766 );
    xnor g24904 ( n38181 , n19660 , n19929 );
    xnor g24905 ( n17974 , n36998 , n22751 );
    and g24906 ( n41414 , n25386 , n20536 );
    nor g24907 ( n12764 , n6982 , n30784 );
    nor g24908 ( n29309 , n27658 , n9713 );
    and g24909 ( n40270 , n1465 , n16375 );
    not g24910 ( n23588 , n32599 );
    or g24911 ( n39458 , n34089 , n9895 );
    and g24912 ( n25865 , n27170 , n11926 );
    or g24913 ( n39703 , n24632 , n18564 );
    or g24914 ( n36624 , n38857 , n5637 );
    or g24915 ( n14322 , n5341 , n5059 );
    xnor g24916 ( n7844 , n24119 , n17744 );
    not g24917 ( n17130 , n768 );
    or g24918 ( n29597 , n14461 , n3897 );
    xnor g24919 ( n16874 , n21973 , n7719 );
    not g24920 ( n1110 , n426 );
    or g24921 ( n36271 , n20148 , n11987 );
    or g24922 ( n2343 , n40253 , n7213 );
    and g24923 ( n4046 , n16371 , n8728 );
    and g24924 ( n41475 , n2368 , n20793 );
    and g24925 ( n13145 , n19252 , n1981 );
    not g24926 ( n4294 , n9953 );
    or g24927 ( n39591 , n2820 , n20343 );
    or g24928 ( n4943 , n17314 , n30969 );
    or g24929 ( n27239 , n38433 , n12128 );
    and g24930 ( n8817 , n19576 , n42749 );
    or g24931 ( n36317 , n23325 , n41131 );
    not g24932 ( n4063 , n11176 );
    and g24933 ( n20350 , n26160 , n34897 );
    or g24934 ( n14771 , n11404 , n8344 );
    and g24935 ( n41694 , n546 , n10585 );
    xnor g24936 ( n6069 , n10005 , n33440 );
    or g24937 ( n18846 , n17322 , n18165 );
    or g24938 ( n33811 , n17277 , n37852 );
    or g24939 ( n15549 , n22391 , n1580 );
    and g24940 ( n41458 , n4882 , n37619 );
    or g24941 ( n20325 , n22371 , n19652 );
    or g24942 ( n26444 , n27389 , n26888 );
    not g24943 ( n15599 , n2970 );
    and g24944 ( n25989 , n17360 , n18352 );
    and g24945 ( n11254 , n26414 , n23016 );
    not g24946 ( n35483 , n24531 );
    or g24947 ( n34257 , n30879 , n27111 );
    or g24948 ( n31661 , n40182 , n12727 );
    or g24949 ( n39965 , n41705 , n17678 );
    and g24950 ( n31430 , n9629 , n39419 );
    or g24951 ( n2521 , n26421 , n1416 );
    or g24952 ( n16557 , n19744 , n16008 );
    or g24953 ( n19977 , n11809 , n10898 );
    xnor g24954 ( n23025 , n17264 , n41681 );
    or g24955 ( n19938 , n3989 , n27325 );
    xnor g24956 ( n21930 , n29796 , n21695 );
    not g24957 ( n24625 , n34414 );
    xnor g24958 ( n38572 , n28431 , n4482 );
    or g24959 ( n28933 , n28372 , n5722 );
    or g24960 ( n5129 , n12410 , n336 );
    and g24961 ( n39487 , n41023 , n42719 );
    xnor g24962 ( n1275 , n29375 , n18781 );
    or g24963 ( n19534 , n18236 , n15897 );
    not g24964 ( n1554 , n32544 );
    or g24965 ( n19328 , n30060 , n28748 );
    or g24966 ( n15873 , n18754 , n19701 );
    not g24967 ( n28468 , n39226 );
    or g24968 ( n27427 , n34589 , n9059 );
    or g24969 ( n30000 , n24217 , n39260 );
    or g24970 ( n4488 , n9809 , n6158 );
    or g24971 ( n25982 , n36296 , n7031 );
    or g24972 ( n33246 , n28452 , n7374 );
    or g24973 ( n21517 , n6083 , n41555 );
    or g24974 ( n24731 , n17359 , n16140 );
    or g24975 ( n27634 , n12543 , n11346 );
    or g24976 ( n29876 , n1932 , n39268 );
    or g24977 ( n7632 , n31924 , n5265 );
    or g24978 ( n37688 , n38558 , n2597 );
    nor g24979 ( n37191 , n17744 , n32123 );
    and g24980 ( n14791 , n12561 , n41490 );
    not g24981 ( n10437 , n19499 );
    and g24982 ( n37951 , n14399 , n37310 );
    and g24983 ( n22275 , n24541 , n919 );
    and g24984 ( n32707 , n6058 , n18600 );
    or g24985 ( n18336 , n10333 , n19497 );
    and g24986 ( n39972 , n38941 , n24351 );
    or g24987 ( n38716 , n27799 , n34066 );
    not g24988 ( n9245 , n38217 );
    nor g24989 ( n40471 , n1232 , n27556 );
    nor g24990 ( n13999 , n11436 , n34644 );
    not g24991 ( n9635 , n28077 );
    or g24992 ( n5435 , n20175 , n41993 );
    or g24993 ( n3175 , n23769 , n25696 );
    or g24994 ( n25548 , n37119 , n13582 );
    or g24995 ( n41882 , n2781 , n39108 );
    and g24996 ( n35707 , n27843 , n19703 );
    and g24997 ( n29580 , n21459 , n32144 );
    xnor g24998 ( n14823 , n27762 , n25300 );
    nor g24999 ( n8073 , n383 , n5587 );
    not g25000 ( n11844 , n27629 );
    nor g25001 ( n24060 , n35193 , n1454 );
    or g25002 ( n2396 , n9544 , n10378 );
    xnor g25003 ( n25726 , n21534 , n6563 );
    and g25004 ( n36061 , n7846 , n29307 );
    xnor g25005 ( n11992 , n31099 , n34477 );
    nor g25006 ( n33204 , n32277 , n34588 );
    and g25007 ( n40272 , n38134 , n1690 );
    and g25008 ( n33619 , n26135 , n14887 );
    or g25009 ( n2306 , n39236 , n14086 );
    nor g25010 ( n9779 , n41534 , n30587 );
    or g25011 ( n40493 , n29303 , n28453 );
    and g25012 ( n37161 , n26835 , n23481 );
    or g25013 ( n27791 , n34292 , n4797 );
    nor g25014 ( n1381 , n3955 , n6448 );
    nor g25015 ( n15663 , n20285 , n6014 );
    xnor g25016 ( n38668 , n39852 , n13421 );
    and g25017 ( n32483 , n2707 , n1262 );
    xnor g25018 ( n432 , n12304 , n33429 );
    xnor g25019 ( n643 , n18456 , n14471 );
    or g25020 ( n36190 , n41534 , n8951 );
    and g25021 ( n4365 , n25027 , n16269 );
    and g25022 ( n12371 , n16202 , n40134 );
    nor g25023 ( n42184 , n40128 , n35303 );
    and g25024 ( n25670 , n14562 , n33140 );
    and g25025 ( n9087 , n6028 , n39601 );
    nor g25026 ( n19156 , n14467 , n41139 );
    and g25027 ( n5449 , n3018 , n7591 );
    not g25028 ( n8049 , n42051 );
    or g25029 ( n28488 , n2628 , n8533 );
    not g25030 ( n12442 , n7236 );
    or g25031 ( n33818 , n35483 , n33527 );
    and g25032 ( n16692 , n8684 , n27462 );
    nor g25033 ( n3089 , n4340 , n11196 );
    nor g25034 ( n34038 , n37538 , n12275 );
    xnor g25035 ( n5230 , n24218 , n16192 );
    and g25036 ( n39789 , n26415 , n324 );
    not g25037 ( n21592 , n32118 );
    and g25038 ( n22127 , n736 , n33899 );
    or g25039 ( n846 , n22175 , n31313 );
    nor g25040 ( n31832 , n38122 , n30322 );
    or g25041 ( n41792 , n6667 , n20498 );
    and g25042 ( n30225 , n2717 , n24244 );
    nor g25043 ( n4668 , n36993 , n37566 );
    nor g25044 ( n5307 , n17577 , n27605 );
    or g25045 ( n19670 , n42340 , n28561 );
    not g25046 ( n37241 , n14004 );
    or g25047 ( n14106 , n36394 , n7050 );
    or g25048 ( n3450 , n26399 , n29857 );
    or g25049 ( n20002 , n4669 , n32320 );
    or g25050 ( n14163 , n24062 , n41561 );
    and g25051 ( n30362 , n13418 , n32432 );
    not g25052 ( n14441 , n597 );
    not g25053 ( n33797 , n5734 );
    not g25054 ( n14614 , n40725 );
    or g25055 ( n3682 , n11309 , n21770 );
    not g25056 ( n34254 , n12773 );
    xnor g25057 ( n10289 , n14821 , n3564 );
    not g25058 ( n10045 , n28850 );
    or g25059 ( n40564 , n12987 , n7326 );
    xnor g25060 ( n32278 , n36356 , n9683 );
    not g25061 ( n39104 , n40499 );
    nor g25062 ( n4381 , n18866 , n36061 );
    not g25063 ( n37563 , n27953 );
    or g25064 ( n26048 , n38053 , n7373 );
    not g25065 ( n40110 , n17598 );
    nor g25066 ( n472 , n4967 , n31340 );
    not g25067 ( n2445 , n25893 );
    xnor g25068 ( n16062 , n20920 , n21433 );
    not g25069 ( n31992 , n17234 );
    or g25070 ( n38788 , n40074 , n40253 );
    or g25071 ( n33229 , n28725 , n36861 );
    not g25072 ( n19114 , n38562 );
    or g25073 ( n692 , n7370 , n16935 );
    xnor g25074 ( n38503 , n6625 , n35160 );
    xnor g25075 ( n17790 , n29796 , n41858 );
    and g25076 ( n1644 , n23089 , n24335 );
    xnor g25077 ( n6369 , n383 , n16839 );
    or g25078 ( n5314 , n12110 , n33590 );
    not g25079 ( n7339 , n25207 );
    or g25080 ( n1016 , n7882 , n1361 );
    and g25081 ( n12056 , n6285 , n31316 );
    or g25082 ( n6803 , n18625 , n36765 );
    and g25083 ( n2512 , n12261 , n16555 );
    not g25084 ( n9201 , n38399 );
    nor g25085 ( n37207 , n16211 , n14223 );
    or g25086 ( n11187 , n25875 , n16839 );
    xnor g25087 ( n21287 , n16406 , n32418 );
    not g25088 ( n34317 , n34693 );
    nor g25089 ( n31351 , n36062 , n40729 );
    or g25090 ( n1953 , n12577 , n40481 );
    nor g25091 ( n19270 , n26067 , n25320 );
    or g25092 ( n8471 , n4282 , n19069 );
    or g25093 ( n9170 , n41126 , n16216 );
    and g25094 ( n12831 , n10449 , n38137 );
    or g25095 ( n39013 , n19436 , n41565 );
    and g25096 ( n16479 , n25337 , n26890 );
    or g25097 ( n14872 , n16967 , n15671 );
    not g25098 ( n9062 , n20714 );
    or g25099 ( n41593 , n19619 , n39674 );
    or g25100 ( n26629 , n14047 , n837 );
    or g25101 ( n9606 , n16608 , n13885 );
    or g25102 ( n32438 , n41666 , n13912 );
    not g25103 ( n29281 , n15117 );
    or g25104 ( n33894 , n5657 , n11030 );
    or g25105 ( n40490 , n28395 , n9539 );
    and g25106 ( n30318 , n21317 , n9330 );
    nor g25107 ( n29337 , n23727 , n30218 );
    and g25108 ( n16630 , n7439 , n39995 );
    not g25109 ( n19762 , n29713 );
    nor g25110 ( n25553 , n22967 , n7749 );
    and g25111 ( n23241 , n27604 , n36075 );
    or g25112 ( n40835 , n28349 , n40118 );
    not g25113 ( n7922 , n32119 );
    not g25114 ( n27540 , n24810 );
    not g25115 ( n7142 , n7818 );
    or g25116 ( n7161 , n3006 , n20183 );
    xnor g25117 ( n4820 , n6962 , n21364 );
    or g25118 ( n25120 , n37139 , n10265 );
    or g25119 ( n27032 , n5324 , n18412 );
    xnor g25120 ( n13389 , n21973 , n35303 );
    and g25121 ( n41592 , n20389 , n35457 );
    and g25122 ( n4096 , n5822 , n32881 );
    or g25123 ( n33660 , n15388 , n41194 );
    and g25124 ( n19113 , n13072 , n38292 );
    or g25125 ( n10750 , n21207 , n40291 );
    xnor g25126 ( n32841 , n17159 , n1694 );
    and g25127 ( n33806 , n38972 , n5797 );
    not g25128 ( n28887 , n29429 );
    or g25129 ( n10868 , n2381 , n19159 );
    or g25130 ( n15103 , n12113 , n21500 );
    or g25131 ( n13001 , n17744 , n33010 );
    not g25132 ( n10041 , n40987 );
    and g25133 ( n6400 , n31411 , n847 );
    not g25134 ( n10535 , n25370 );
    and g25135 ( n9863 , n37316 , n41978 );
    and g25136 ( n38040 , n11899 , n26285 );
    xnor g25137 ( n7877 , n17225 , n15642 );
    not g25138 ( n32351 , n11879 );
    and g25139 ( n36952 , n42624 , n40430 );
    not g25140 ( n15089 , n32485 );
    or g25141 ( n26310 , n19622 , n15421 );
    not g25142 ( n25988 , n35345 );
    or g25143 ( n34865 , n40146 , n10707 );
    nor g25144 ( n12950 , n5001 , n21143 );
    or g25145 ( n12180 , n26102 , n33804 );
    nor g25146 ( n22616 , n35349 , n17337 );
    or g25147 ( n39437 , n23386 , n1608 );
    and g25148 ( n31051 , n41507 , n23508 );
    or g25149 ( n10538 , n22610 , n7411 );
    and g25150 ( n34204 , n6569 , n5527 );
    or g25151 ( n9834 , n25959 , n1286 );
    and g25152 ( n17602 , n32366 , n16097 );
    or g25153 ( n8833 , n34031 , n13577 );
    not g25154 ( n33974 , n13506 );
    xnor g25155 ( n28730 , n42898 , n22652 );
    not g25156 ( n41629 , n32393 );
    or g25157 ( n9856 , n18390 , n30193 );
    and g25158 ( n11620 , n5276 , n38312 );
    nor g25159 ( n13320 , n22041 , n30551 );
    or g25160 ( n25636 , n32729 , n12684 );
    xnor g25161 ( n33777 , n13224 , n34727 );
    or g25162 ( n14158 , n1896 , n40407 );
    and g25163 ( n18778 , n13382 , n260 );
    and g25164 ( n23380 , n31373 , n9661 );
    nor g25165 ( n11866 , n25588 , n20407 );
    nor g25166 ( n24151 , n18914 , n11305 );
    or g25167 ( n9425 , n38879 , n36379 );
    and g25168 ( n29493 , n24359 , n10607 );
    not g25169 ( n1149 , n30062 );
    not g25170 ( n34225 , n23239 );
    nor g25171 ( n26868 , n40621 , n32631 );
    and g25172 ( n23589 , n29505 , n28504 );
    or g25173 ( n13304 , n34527 , n39550 );
    or g25174 ( n2911 , n24626 , n16563 );
    or g25175 ( n9640 , n15350 , n30235 );
    not g25176 ( n30376 , n41231 );
    or g25177 ( n3182 , n5348 , n30886 );
    or g25178 ( n1364 , n5179 , n35101 );
    not g25179 ( n13174 , n28821 );
    not g25180 ( n41859 , n3265 );
    and g25181 ( n41717 , n3784 , n31642 );
    or g25182 ( n18602 , n33691 , n1910 );
    nor g25183 ( n23844 , n13900 , n5074 );
    and g25184 ( n40741 , n5523 , n10426 );
    or g25185 ( n32292 , n21031 , n3728 );
    or g25186 ( n40627 , n39776 , n25924 );
    and g25187 ( n26755 , n11865 , n30577 );
    and g25188 ( n41479 , n22207 , n26798 );
    and g25189 ( n28249 , n15336 , n41452 );
    or g25190 ( n32692 , n36464 , n37767 );
    not g25191 ( n25423 , n39727 );
    not g25192 ( n4951 , n23193 );
    and g25193 ( n2013 , n30469 , n4894 );
    or g25194 ( n28550 , n27511 , n25449 );
    and g25195 ( n7260 , n8121 , n26936 );
    or g25196 ( n30079 , n21177 , n36511 );
    not g25197 ( n1812 , n40161 );
    or g25198 ( n1802 , n16328 , n38303 );
    or g25199 ( n24932 , n634 , n40702 );
    not g25200 ( n10092 , n23514 );
    or g25201 ( n4759 , n42798 , n1295 );
    or g25202 ( n14073 , n18081 , n12896 );
    or g25203 ( n10357 , n14296 , n26183 );
    nor g25204 ( n40798 , n19630 , n33546 );
    and g25205 ( n38559 , n18530 , n12010 );
    or g25206 ( n95 , n3309 , n28743 );
    not g25207 ( n5941 , n26366 );
    or g25208 ( n39633 , n38993 , n29299 );
    or g25209 ( n9565 , n36217 , n12361 );
    nor g25210 ( n16149 , n27745 , n40656 );
    xnor g25211 ( n2780 , n5041 , n38281 );
    or g25212 ( n9002 , n1670 , n23301 );
    and g25213 ( n21080 , n21522 , n3463 );
    not g25214 ( n24656 , n16075 );
    xnor g25215 ( n23980 , n24163 , n37220 );
    and g25216 ( n40894 , n25197 , n40998 );
    nor g25217 ( n9023 , n6957 , n35032 );
    or g25218 ( n11302 , n15282 , n16734 );
    or g25219 ( n39132 , n14922 , n13992 );
    or g25220 ( n5301 , n2831 , n35178 );
    or g25221 ( n998 , n7589 , n8090 );
    or g25222 ( n15312 , n19129 , n39635 );
    or g25223 ( n16707 , n7826 , n14762 );
    not g25224 ( n19095 , n24646 );
    xnor g25225 ( n4912 , n11436 , n23582 );
    or g25226 ( n15543 , n21328 , n7703 );
    not g25227 ( n37434 , n23595 );
    or g25228 ( n14778 , n10537 , n14301 );
    and g25229 ( n20754 , n24443 , n7684 );
    and g25230 ( n33819 , n14639 , n5020 );
    or g25231 ( n6844 , n17839 , n41521 );
    not g25232 ( n36747 , n35896 );
    or g25233 ( n19823 , n24656 , n33986 );
    or g25234 ( n11372 , n16607 , n24183 );
    and g25235 ( n23872 , n16861 , n19621 );
    or g25236 ( n15901 , n24808 , n32219 );
    and g25237 ( n10472 , n21488 , n20462 );
    and g25238 ( n2617 , n4555 , n10662 );
    or g25239 ( n41751 , n12643 , n35637 );
    or g25240 ( n3399 , n24656 , n25896 );
    or g25241 ( n8236 , n1290 , n11814 );
    not g25242 ( n22563 , n21978 );
    and g25243 ( n26338 , n22168 , n33821 );
    or g25244 ( n15828 , n30483 , n18074 );
    not g25245 ( n5049 , n631 );
    or g25246 ( n28100 , n16199 , n10698 );
    or g25247 ( n8754 , n7020 , n3972 );
    xnor g25248 ( n12860 , n4664 , n17193 );
    and g25249 ( n19496 , n21689 , n21395 );
    and g25250 ( n20925 , n21968 , n25479 );
    not g25251 ( n8427 , n24891 );
    or g25252 ( n20674 , n15959 , n1044 );
    or g25253 ( n36414 , n17256 , n8703 );
    not g25254 ( n12699 , n28459 );
    or g25255 ( n36992 , n39043 , n5984 );
    or g25256 ( n8599 , n31967 , n4854 );
    or g25257 ( n9761 , n26612 , n3868 );
    not g25258 ( n17292 , n9429 );
    and g25259 ( n8498 , n27862 , n31506 );
    xnor g25260 ( n28527 , n9878 , n7600 );
    nor g25261 ( n32869 , n23330 , n39342 );
    not g25262 ( n28424 , n17774 );
    and g25263 ( n5657 , n41419 , n17046 );
    not g25264 ( n35476 , n24875 );
    nor g25265 ( n28961 , n17193 , n13059 );
    xnor g25266 ( n31548 , n37922 , n13122 );
    xnor g25267 ( n4636 , n13444 , n41456 );
    and g25268 ( n35100 , n9323 , n581 );
    xnor g25269 ( n17112 , n8346 , n16598 );
    nor g25270 ( n14793 , n9793 , n38036 );
    nor g25271 ( n32939 , n14091 , n28116 );
    or g25272 ( n20024 , n2548 , n16025 );
    or g25273 ( n31935 , n26122 , n39080 );
    or g25274 ( n30158 , n29552 , n5683 );
    or g25275 ( n41760 , n14252 , n30290 );
    and g25276 ( n26882 , n33050 , n35079 );
    and g25277 ( n9599 , n39069 , n32790 );
    not g25278 ( n26174 , n17825 );
    xnor g25279 ( n11149 , n12440 , n19147 );
    not g25280 ( n12514 , n29560 );
    and g25281 ( n28337 , n2737 , n12678 );
    not g25282 ( n2575 , n24799 );
    and g25283 ( n19871 , n24079 , n12844 );
    not g25284 ( n23204 , n33920 );
    not g25285 ( n1617 , n9637 );
    not g25286 ( n26332 , n32596 );
    or g25287 ( n40266 , n22409 , n27679 );
    nor g25288 ( n35284 , n1197 , n12198 );
    or g25289 ( n12095 , n26634 , n37952 );
    or g25290 ( n32481 , n1381 , n29833 );
    and g25291 ( n26808 , n33395 , n22200 );
    not g25292 ( n40755 , n31072 );
    not g25293 ( n26577 , n23030 );
    and g25294 ( n13478 , n38667 , n37121 );
    and g25295 ( n21857 , n27876 , n13688 );
    not g25296 ( n30463 , n6196 );
    and g25297 ( n36658 , n38774 , n16522 );
    xnor g25298 ( n12785 , n34731 , n11306 );
    and g25299 ( n30795 , n31682 , n10686 );
    not g25300 ( n8015 , n42239 );
    not g25301 ( n10675 , n35344 );
    not g25302 ( n35534 , n3264 );
    and g25303 ( n6458 , n10831 , n30718 );
    buf g25304 ( n27663 , n2495 );
    nor g25305 ( n32635 , n9507 , n37192 );
    or g25306 ( n1635 , n18244 , n24303 );
    or g25307 ( n37382 , n7839 , n3978 );
    or g25308 ( n137 , n16433 , n29545 );
    or g25309 ( n17012 , n25890 , n14281 );
    nor g25310 ( n13496 , n5197 , n33940 );
    or g25311 ( n22936 , n10669 , n23563 );
    and g25312 ( n39993 , n37797 , n25797 );
    or g25313 ( n25718 , n15070 , n28330 );
    and g25314 ( n31858 , n12949 , n36670 );
    or g25315 ( n5943 , n16682 , n9014 );
    and g25316 ( n28401 , n17308 , n12036 );
    nor g25317 ( n32498 , n5964 , n38160 );
    and g25318 ( n16220 , n25815 , n30494 );
    or g25319 ( n36207 , n15392 , n23857 );
    and g25320 ( n15542 , n40549 , n2984 );
    or g25321 ( n38593 , n18181 , n25451 );
    xnor g25322 ( n15700 , n42030 , n33019 );
    or g25323 ( n13211 , n5722 , n37105 );
    or g25324 ( n8634 , n10557 , n367 );
    not g25325 ( n11989 , n29883 );
    and g25326 ( n39775 , n15398 , n3711 );
    and g25327 ( n11511 , n38496 , n27807 );
    xnor g25328 ( n29670 , n11436 , n40984 );
    and g25329 ( n37231 , n14425 , n8456 );
    xnor g25330 ( n27710 , n22799 , n15791 );
    or g25331 ( n7499 , n30321 , n25213 );
    or g25332 ( n25952 , n17910 , n38945 );
    or g25333 ( n25703 , n8661 , n5766 );
    and g25334 ( n12000 , n10876 , n18509 );
    not g25335 ( n24068 , n22953 );
    not g25336 ( n28341 , n1931 );
    or g25337 ( n42839 , n34150 , n42896 );
    not g25338 ( n425 , n22533 );
    or g25339 ( n24311 , n39182 , n10669 );
    nor g25340 ( n4454 , n16620 , n17126 );
    and g25341 ( n41240 , n14594 , n39998 );
    or g25342 ( n22877 , n11336 , n30122 );
    and g25343 ( n17503 , n663 , n4518 );
    or g25344 ( n20358 , n15112 , n16882 );
    or g25345 ( n25327 , n42540 , n1326 );
    and g25346 ( n2833 , n18112 , n11223 );
    or g25347 ( n29554 , n23971 , n9865 );
    not g25348 ( n11413 , n5462 );
    or g25349 ( n40631 , n40024 , n42394 );
    xnor g25350 ( n4481 , n29323 , n16995 );
    not g25351 ( n19880 , n36388 );
    not g25352 ( n7904 , n10943 );
    xnor g25353 ( n42062 , n18880 , n10533 );
    nor g25354 ( n36036 , n18954 , n42841 );
    and g25355 ( n26988 , n7205 , n42075 );
    or g25356 ( n28091 , n24738 , n25440 );
    or g25357 ( n33079 , n14945 , n23590 );
    not g25358 ( n30422 , n19617 );
    or g25359 ( n14947 , n20138 , n8797 );
    nor g25360 ( n4092 , n22161 , n26769 );
    not g25361 ( n20078 , n5578 );
    nor g25362 ( n10664 , n1507 , n33235 );
    and g25363 ( n28891 , n20603 , n13727 );
    nor g25364 ( n25509 , n1507 , n32221 );
    and g25365 ( n5120 , n604 , n37731 );
    or g25366 ( n17834 , n21539 , n1347 );
    xnor g25367 ( n17674 , n32297 , n41331 );
    or g25368 ( n16110 , n41767 , n364 );
    xnor g25369 ( n40754 , n3752 , n15575 );
    and g25370 ( n40102 , n815 , n24921 );
    xnor g25371 ( n29083 , n14932 , n19303 );
    or g25372 ( n40778 , n14155 , n20446 );
    xnor g25373 ( n27667 , n36899 , n41152 );
    or g25374 ( n21699 , n7669 , n22031 );
    xnor g25375 ( n5344 , n41013 , n31109 );
    and g25376 ( n26159 , n16713 , n21161 );
    and g25377 ( n2514 , n23970 , n15785 );
    or g25378 ( n11853 , n38160 , n41487 );
    and g25379 ( n26690 , n18858 , n284 );
    xnor g25380 ( n7540 , n5441 , n6839 );
    xnor g25381 ( n20986 , n24210 , n40036 );
    not g25382 ( n2839 , n32573 );
    nor g25383 ( n34270 , n39266 , n35736 );
    nor g25384 ( n14484 , n10598 , n41331 );
    or g25385 ( n42719 , n18651 , n19608 );
    not g25386 ( n39481 , n36942 );
    not g25387 ( n16211 , n30463 );
    or g25388 ( n11712 , n31491 , n11410 );
    xnor g25389 ( n30311 , n28497 , n30149 );
    and g25390 ( n38031 , n32452 , n21119 );
    nor g25391 ( n33118 , n11531 , n30871 );
    or g25392 ( n38907 , n26690 , n34044 );
    or g25393 ( n7722 , n1314 , n21886 );
    xnor g25394 ( n31538 , n19453 , n36709 );
    or g25395 ( n34538 , n35952 , n39906 );
    or g25396 ( n28641 , n19775 , n1184 );
    or g25397 ( n32816 , n32068 , n39848 );
    and g25398 ( n13099 , n7528 , n22500 );
    or g25399 ( n11055 , n12198 , n21887 );
    or g25400 ( n23390 , n14112 , n13435 );
    and g25401 ( n10199 , n37287 , n4073 );
    or g25402 ( n13705 , n23261 , n839 );
    or g25403 ( n37882 , n5480 , n9617 );
    and g25404 ( n18310 , n5400 , n18054 );
    and g25405 ( n20776 , n14922 , n13992 );
    or g25406 ( n33188 , n3870 , n15505 );
    and g25407 ( n34959 , n16161 , n3400 );
    not g25408 ( n35712 , n23883 );
    and g25409 ( n38909 , n5130 , n5047 );
    and g25410 ( n17341 , n7781 , n34252 );
    or g25411 ( n32166 , n24547 , n19963 );
    xnor g25412 ( n39562 , n35217 , n21393 );
    nor g25413 ( n26696 , n6840 , n27358 );
    and g25414 ( n13640 , n2161 , n5595 );
    or g25415 ( n12073 , n935 , n37784 );
    nor g25416 ( n3472 , n962 , n144 );
    or g25417 ( n42390 , n528 , n21333 );
    and g25418 ( n27675 , n35498 , n20951 );
    and g25419 ( n9901 , n20264 , n22498 );
    or g25420 ( n7519 , n18239 , n23936 );
    not g25421 ( n9210 , n34076 );
    nor g25422 ( n33281 , n42445 , n26200 );
    nor g25423 ( n31982 , n10831 , n30718 );
    or g25424 ( n2023 , n7020 , n24461 );
    and g25425 ( n25304 , n30416 , n37002 );
    and g25426 ( n31473 , n4557 , n10080 );
    and g25427 ( n1756 , n10417 , n38846 );
    or g25428 ( n41638 , n17539 , n2530 );
    not g25429 ( n31973 , n19485 );
    and g25430 ( n16793 , n19945 , n18306 );
    xnor g25431 ( n40012 , n12806 , n28991 );
    or g25432 ( n36847 , n14552 , n9402 );
    nor g25433 ( n14762 , n2387 , n2178 );
    and g25434 ( n5852 , n19739 , n22803 );
    not g25435 ( n36863 , n33702 );
    and g25436 ( n18574 , n10577 , n20903 );
    and g25437 ( n31015 , n15814 , n35496 );
    nor g25438 ( n37948 , n34337 , n40035 );
    or g25439 ( n41659 , n17770 , n5805 );
    and g25440 ( n9468 , n35248 , n25134 );
    nor g25441 ( n29327 , n9528 , n35810 );
    or g25442 ( n19198 , n13061 , n13830 );
    or g25443 ( n17283 , n28143 , n23742 );
    not g25444 ( n21951 , n29836 );
    nor g25445 ( n36820 , n30742 , n13625 );
    or g25446 ( n34367 , n10855 , n19594 );
    xnor g25447 ( n11488 , n20855 , n5964 );
    or g25448 ( n5050 , n1581 , n10801 );
    and g25449 ( n28624 , n26687 , n1964 );
    or g25450 ( n30880 , n28360 , n41868 );
    nor g25451 ( n16559 , n27808 , n1185 );
    xnor g25452 ( n761 , n12146 , n33878 );
    or g25453 ( n36912 , n19892 , n11403 );
    nor g25454 ( n3989 , n4102 , n6718 );
    and g25455 ( n25996 , n5334 , n15407 );
    or g25456 ( n6057 , n11091 , n20932 );
    or g25457 ( n24548 , n24626 , n21791 );
    and g25458 ( n37060 , n243 , n1196 );
    and g25459 ( n35742 , n30740 , n11000 );
    or g25460 ( n14058 , n14362 , n1134 );
    and g25461 ( n13750 , n39549 , n8350 );
    not g25462 ( n12146 , n15070 );
    not g25463 ( n19178 , n25899 );
    or g25464 ( n283 , n34424 , n22991 );
    nor g25465 ( n28002 , n38267 , n33477 );
    not g25466 ( n14594 , n7035 );
    xnor g25467 ( n28781 , n11436 , n22146 );
    or g25468 ( n21227 , n23476 , n17318 );
    or g25469 ( n16275 , n14944 , n40342 );
    or g25470 ( n24703 , n37963 , n42522 );
    and g25471 ( n34720 , n14947 , n22600 );
    xnor g25472 ( n35000 , n34844 , n27275 );
    and g25473 ( n15397 , n36740 , n7038 );
    not g25474 ( n22201 , n15133 );
    and g25475 ( n28392 , n32570 , n786 );
    not g25476 ( n31688 , n27243 );
    or g25477 ( n20380 , n23675 , n37434 );
    or g25478 ( n992 , n18798 , n18978 );
    or g25479 ( n7168 , n22427 , n33748 );
    or g25480 ( n3599 , n32512 , n10295 );
    and g25481 ( n12863 , n41133 , n18943 );
    and g25482 ( n13193 , n4315 , n10841 );
    or g25483 ( n19395 , n10815 , n12220 );
    xnor g25484 ( n27653 , n40 , n23842 );
    or g25485 ( n14543 , n39365 , n30665 );
    not g25486 ( n27968 , n4822 );
    or g25487 ( n22965 , n42140 , n19803 );
    not g25488 ( n14213 , n2587 );
    or g25489 ( n24065 , n19379 , n39108 );
    and g25490 ( n38340 , n7554 , n7431 );
    xnor g25491 ( n6002 , n20489 , n17846 );
    and g25492 ( n10506 , n12569 , n33980 );
    and g25493 ( n11507 , n9262 , n9261 );
    and g25494 ( n25168 , n36480 , n26774 );
    or g25495 ( n21030 , n20740 , n3935 );
    not g25496 ( n41040 , n26242 );
    or g25497 ( n8005 , n32461 , n17170 );
    xnor g25498 ( n89 , n20721 , n16598 );
    not g25499 ( n24876 , n5912 );
    or g25500 ( n28268 , n40509 , n34609 );
    or g25501 ( n10553 , n8031 , n40534 );
    not g25502 ( n22444 , n13234 );
    or g25503 ( n34381 , n15064 , n8002 );
    or g25504 ( n8317 , n7856 , n22516 );
    nor g25505 ( n6074 , n36164 , n13168 );
    nor g25506 ( n34623 , n41761 , n39507 );
    nor g25507 ( n8080 , n17393 , n37289 );
    not g25508 ( n11295 , n38486 );
    not g25509 ( n29346 , n42331 );
    and g25510 ( n23749 , n1526 , n1594 );
    not g25511 ( n8412 , n42197 );
    not g25512 ( n30821 , n8565 );
    xnor g25513 ( n32990 , n31460 , n38223 );
    not g25514 ( n14168 , n29650 );
    or g25515 ( n26302 , n16586 , n16504 );
    or g25516 ( n21508 , n4521 , n18665 );
    nor g25517 ( n38363 , n38879 , n7490 );
    xnor g25518 ( n32738 , n28083 , n40741 );
    or g25519 ( n15407 , n25352 , n18016 );
    not g25520 ( n31864 , n26100 );
    and g25521 ( n29841 , n9180 , n31713 );
    or g25522 ( n40273 , n20092 , n24241 );
    or g25523 ( n36081 , n25964 , n38254 );
    xnor g25524 ( n35525 , n22879 , n35417 );
    not g25525 ( n42333 , n22587 );
    or g25526 ( n17929 , n328 , n15305 );
    nor g25527 ( n33488 , n23115 , n14692 );
    nor g25528 ( n23553 , n13969 , n29869 );
    not g25529 ( n35395 , n21165 );
    or g25530 ( n10189 , n33095 , n18846 );
    not g25531 ( n7289 , n4178 );
    nor g25532 ( n3902 , n24127 , n6114 );
    or g25533 ( n41184 , n10559 , n9390 );
    or g25534 ( n30548 , n35764 , n13742 );
    or g25535 ( n4968 , n2330 , n25440 );
    not g25536 ( n34356 , n6876 );
    not g25537 ( n13388 , n22414 );
    and g25538 ( n7180 , n36004 , n21768 );
    or g25539 ( n3163 , n20901 , n22885 );
    or g25540 ( n29044 , n25499 , n26170 );
    and g25541 ( n6672 , n19704 , n37528 );
    xnor g25542 ( n24822 , n30692 , n12301 );
    nor g25543 ( n39210 , n35653 , n36651 );
    nor g25544 ( n2066 , n17120 , n21098 );
    and g25545 ( n2227 , n8396 , n39103 );
    or g25546 ( n13137 , n5839 , n6290 );
    and g25547 ( n27240 , n13189 , n18972 );
    nor g25548 ( n4994 , n25974 , n17835 );
    or g25549 ( n21383 , n39150 , n25567 );
    not g25550 ( n5320 , n24856 );
    not g25551 ( n30637 , n39807 );
    and g25552 ( n37947 , n38351 , n3328 );
    not g25553 ( n22282 , n36521 );
    or g25554 ( n11590 , n12722 , n19993 );
    not g25555 ( n42697 , n27702 );
    not g25556 ( n1765 , n26575 );
    or g25557 ( n2361 , n30674 , n32745 );
    or g25558 ( n6084 , n5110 , n29634 );
    xnor g25559 ( n5268 , n22263 , n7752 );
    not g25560 ( n21293 , n42915 );
    xnor g25561 ( n20879 , n5891 , n35495 );
    or g25562 ( n13749 , n13961 , n23210 );
    nor g25563 ( n5396 , n15678 , n37753 );
    and g25564 ( n10515 , n42102 , n23223 );
    and g25565 ( n37303 , n26152 , n18336 );
    or g25566 ( n955 , n23749 , n38720 );
    or g25567 ( n23628 , n32663 , n27416 );
    not g25568 ( n5259 , n9210 );
    or g25569 ( n42038 , n20138 , n8358 );
    or g25570 ( n5214 , n3526 , n8732 );
    not g25571 ( n28333 , n27308 );
    or g25572 ( n16356 , n3396 , n31098 );
    and g25573 ( n15065 , n40330 , n12263 );
    xnor g25574 ( n32484 , n23995 , n25588 );
    and g25575 ( n18572 , n36612 , n31767 );
    and g25576 ( n1414 , n18440 , n18397 );
    not g25577 ( n16530 , n2486 );
    or g25578 ( n8789 , n39940 , n25959 );
    or g25579 ( n32653 , n14851 , n32149 );
    and g25580 ( n8586 , n32287 , n40677 );
    nor g25581 ( n11425 , n30262 , n23354 );
    or g25582 ( n42402 , n32217 , n26604 );
    or g25583 ( n5125 , n2517 , n42205 );
    nor g25584 ( n24170 , n34565 , n34896 );
    or g25585 ( n41795 , n4416 , n18243 );
    or g25586 ( n26829 , n24779 , n17468 );
    not g25587 ( n842 , n13111 );
    or g25588 ( n36643 , n33081 , n7290 );
    not g25589 ( n39439 , n41758 );
    xnor g25590 ( n14645 , n35000 , n19896 );
    or g25591 ( n30988 , n41572 , n40987 );
    or g25592 ( n15954 , n2507 , n36383 );
    and g25593 ( n26910 , n13680 , n3110 );
    and g25594 ( n18009 , n236 , n40037 );
    and g25595 ( n35036 , n23705 , n4242 );
    or g25596 ( n3143 , n2404 , n21048 );
    and g25597 ( n21596 , n16422 , n15996 );
    and g25598 ( n12171 , n40463 , n39271 );
    or g25599 ( n12741 , n31265 , n28803 );
    or g25600 ( n22981 , n39986 , n32100 );
    xnor g25601 ( n6552 , n9180 , n13375 );
    not g25602 ( n5009 , n21474 );
    and g25603 ( n2897 , n37311 , n31056 );
    and g25604 ( n30993 , n9954 , n13326 );
    or g25605 ( n17600 , n1372 , n38407 );
    nor g25606 ( n3637 , n14471 , n41493 );
    not g25607 ( n34444 , n19629 );
    or g25608 ( n29632 , n4412 , n20953 );
    or g25609 ( n27104 , n40389 , n8322 );
    xnor g25610 ( n18858 , n11436 , n39753 );
    xnor g25611 ( n31434 , n32760 , n34986 );
    or g25612 ( n23230 , n18770 , n28461 );
    nor g25613 ( n11642 , n7688 , n6983 );
    not g25614 ( n27154 , n39293 );
    and g25615 ( n33248 , n3572 , n3846 );
    and g25616 ( n24670 , n13699 , n30259 );
    or g25617 ( n10148 , n21041 , n36162 );
    xnor g25618 ( n21871 , n42064 , n27640 );
    nor g25619 ( n33334 , n25944 , n36968 );
    and g25620 ( n21698 , n13798 , n38291 );
    or g25621 ( n27814 , n10903 , n32295 );
    or g25622 ( n35600 , n25907 , n8127 );
    nor g25623 ( n17963 , n17744 , n10385 );
    nor g25624 ( n16272 , n30909 , n16234 );
    or g25625 ( n2051 , n12535 , n5183 );
    not g25626 ( n10853 , n1371 );
    not g25627 ( n12822 , n32271 );
    or g25628 ( n17233 , n19067 , n11004 );
    nor g25629 ( n15932 , n15070 , n20381 );
    nor g25630 ( n17926 , n20617 , n41046 );
    nor g25631 ( n42828 , n2199 , n16227 );
    or g25632 ( n18405 , n28393 , n25693 );
    not g25633 ( n22811 , n31021 );
    or g25634 ( n36750 , n7794 , n14278 );
    and g25635 ( n6279 , n14566 , n41991 );
    and g25636 ( n9315 , n24651 , n3825 );
    or g25637 ( n26658 , n9431 , n31415 );
    or g25638 ( n18647 , n19486 , n14707 );
    nor g25639 ( n26684 , n3687 , n32244 );
    or g25640 ( n8268 , n27904 , n21942 );
    or g25641 ( n13026 , n18314 , n33722 );
    not g25642 ( n28530 , n20714 );
    xnor g25643 ( n21995 , n15399 , n1991 );
    or g25644 ( n14924 , n1116 , n4956 );
    not g25645 ( n29858 , n8649 );
    not g25646 ( n33540 , n20857 );
    or g25647 ( n18948 , n35672 , n8275 );
    nor g25648 ( n12429 , n26168 , n37711 );
    xnor g25649 ( n1252 , n26475 , n13587 );
    and g25650 ( n32588 , n11666 , n6700 );
    or g25651 ( n12564 , n14471 , n23742 );
    or g25652 ( n7813 , n18250 , n28241 );
    nor g25653 ( n30 , n34565 , n1436 );
    not g25654 ( n41759 , n29030 );
    or g25655 ( n41708 , n10598 , n6745 );
    xnor g25656 ( n621 , n37829 , n32503 );
    not g25657 ( n21534 , n19221 );
    nor g25658 ( n22944 , n18866 , n16911 );
    not g25659 ( n9586 , n22233 );
    nor g25660 ( n20362 , n26126 , n41255 );
    nor g25661 ( n10609 , n18928 , n724 );
    or g25662 ( n26523 , n13263 , n29825 );
    xnor g25663 ( n5537 , n18990 , n32172 );
    or g25664 ( n1325 , n20817 , n3088 );
    not g25665 ( n35259 , n3693 );
    and g25666 ( n20135 , n10482 , n13015 );
    nor g25667 ( n30060 , n18866 , n15799 );
    or g25668 ( n8154 , n19041 , n12586 );
    or g25669 ( n31064 , n18967 , n23203 );
    not g25670 ( n23585 , n30053 );
    or g25671 ( n20762 , n3131 , n10889 );
    nor g25672 ( n6373 , n39405 , n7830 );
    nor g25673 ( n16208 , n41534 , n20734 );
    not g25674 ( n40225 , n1516 );
    or g25675 ( n33052 , n3238 , n20834 );
    xnor g25676 ( n42687 , n11133 , n33272 );
    and g25677 ( n4593 , n13933 , n18620 );
    not g25678 ( n9971 , n18917 );
    and g25679 ( n10906 , n16080 , n42721 );
    or g25680 ( n21920 , n33115 , n25062 );
    and g25681 ( n25053 , n10640 , n3948 );
    nor g25682 ( n21586 , n14310 , n20397 );
    and g25683 ( n26956 , n33571 , n20480 );
    and g25684 ( n18433 , n28644 , n8811 );
    xnor g25685 ( n35687 , n2799 , n20413 );
    or g25686 ( n37314 , n23882 , n32821 );
    or g25687 ( n10334 , n27924 , n33293 );
    xnor g25688 ( n7812 , n21308 , n24013 );
    or g25689 ( n8112 , n23990 , n29069 );
    or g25690 ( n11856 , n29844 , n29615 );
    or g25691 ( n30965 , n18071 , n16466 );
    or g25692 ( n25663 , n35708 , n9145 );
    or g25693 ( n20335 , n16390 , n31442 );
    not g25694 ( n28896 , n27680 );
    nor g25695 ( n3890 , n28749 , n7873 );
    xnor g25696 ( n38771 , n2350 , n34122 );
    and g25697 ( n12909 , n42583 , n35399 );
    or g25698 ( n41690 , n32159 , n1404 );
    or g25699 ( n10891 , n2698 , n22370 );
    nor g25700 ( n32080 , n5598 , n35150 );
    xnor g25701 ( n15890 , n22753 , n19259 );
    and g25702 ( n30598 , n40012 , n7240 );
    and g25703 ( n34525 , n10920 , n28916 );
    not g25704 ( n23272 , n11047 );
    or g25705 ( n22328 , n3636 , n23632 );
    xnor g25706 ( n29246 , n17137 , n28375 );
    and g25707 ( n1861 , n27828 , n6052 );
    and g25708 ( n24286 , n36160 , n20374 );
    and g25709 ( n30800 , n20944 , n31623 );
    xnor g25710 ( n34427 , n24163 , n4363 );
    not g25711 ( n29404 , n3202 );
    and g25712 ( n19354 , n6226 , n16951 );
    or g25713 ( n24287 , n2303 , n6842 );
    or g25714 ( n36693 , n23673 , n19332 );
    nor g25715 ( n41895 , n20077 , n6208 );
    not g25716 ( n405 , n26959 );
    or g25717 ( n11795 , n18798 , n339 );
    or g25718 ( n17257 , n33152 , n18434 );
    xnor g25719 ( n36450 , n41947 , n16388 );
    or g25720 ( n2676 , n21201 , n28483 );
    nor g25721 ( n12167 , n33981 , n5278 );
    nor g25722 ( n35012 , n4972 , n21833 );
    or g25723 ( n24039 , n38962 , n33151 );
    and g25724 ( n27865 , n33084 , n13427 );
    or g25725 ( n42528 , n40126 , n39481 );
    or g25726 ( n7784 , n798 , n22133 );
    and g25727 ( n4718 , n21281 , n5804 );
    xnor g25728 ( n2161 , n11051 , n23726 );
    nor g25729 ( n42595 , n7870 , n15596 );
    xnor g25730 ( n21895 , n17434 , n38157 );
    xnor g25731 ( n4960 , n40638 , n12540 );
    xnor g25732 ( n24149 , n18678 , n25540 );
    nor g25733 ( n36418 , n5857 , n37301 );
    nor g25734 ( n25410 , n13324 , n41895 );
    and g25735 ( n42302 , n25135 , n4347 );
    not g25736 ( n38479 , n39909 );
    or g25737 ( n12365 , n2800 , n12603 );
    and g25738 ( n9521 , n12503 , n16072 );
    not g25739 ( n30743 , n27308 );
    nor g25740 ( n11523 , n40929 , n27531 );
    or g25741 ( n2621 , n41923 , n6711 );
    or g25742 ( n20244 , n17998 , n37633 );
    not g25743 ( n36998 , n16598 );
    or g25744 ( n31870 , n34738 , n41487 );
    not g25745 ( n27524 , n13002 );
    not g25746 ( n1688 , n14712 );
    and g25747 ( n13446 , n15923 , n3995 );
    or g25748 ( n4093 , n6283 , n34502 );
    nor g25749 ( n14886 , n13801 , n10327 );
    or g25750 ( n6344 , n37031 , n1610 );
    not g25751 ( n37210 , n21246 );
    and g25752 ( n28428 , n35589 , n36611 );
    or g25753 ( n12979 , n12383 , n10194 );
    and g25754 ( n36322 , n30639 , n41842 );
    not g25755 ( n33792 , n1466 );
    not g25756 ( n10666 , n3478 );
    not g25757 ( n13748 , n13951 );
    or g25758 ( n18419 , n35838 , n8518 );
    nor g25759 ( n17339 , n29019 , n24712 );
    or g25760 ( n2291 , n11818 , n36252 );
    or g25761 ( n37283 , n35834 , n16550 );
    or g25762 ( n6973 , n8543 , n25626 );
    xnor g25763 ( n24113 , n24998 , n11405 );
    and g25764 ( n20404 , n33365 , n9670 );
    or g25765 ( n18041 , n1721 , n30575 );
    xnor g25766 ( n6477 , n34731 , n42084 );
    nor g25767 ( n16133 , n17724 , n36501 );
    xnor g25768 ( n33778 , n17200 , n34213 );
    and g25769 ( n3838 , n39713 , n7099 );
    not g25770 ( n40485 , n9146 );
    not g25771 ( n27964 , n19086 );
    or g25772 ( n38516 , n28937 , n20288 );
    xnor g25773 ( n22425 , n12487 , n34241 );
    xnor g25774 ( n27558 , n41695 , n23302 );
    or g25775 ( n32960 , n35068 , n8179 );
    and g25776 ( n16371 , n38985 , n8975 );
    or g25777 ( n21686 , n20561 , n16285 );
    or g25778 ( n38951 , n15282 , n17891 );
    nor g25779 ( n12842 , n31378 , n11645 );
    not g25780 ( n2317 , n27895 );
    or g25781 ( n42271 , n2865 , n10559 );
    nor g25782 ( n13941 , n41859 , n5426 );
    nor g25783 ( n41057 , n23942 , n41252 );
    or g25784 ( n16543 , n22967 , n22914 );
    nor g25785 ( n13324 , n29740 , n31453 );
    or g25786 ( n30146 , n21210 , n28405 );
    nor g25787 ( n13411 , n4869 , n35270 );
    and g25788 ( n21021 , n33840 , n39263 );
    and g25789 ( n13703 , n10594 , n23999 );
    and g25790 ( n11727 , n7960 , n33555 );
    not g25791 ( n8147 , n561 );
    nor g25792 ( n35250 , n40543 , n7251 );
    or g25793 ( n12393 , n19969 , n38473 );
    or g25794 ( n21298 , n18997 , n14547 );
    and g25795 ( n14763 , n26291 , n35812 );
    and g25796 ( n5242 , n36749 , n6922 );
    or g25797 ( n16853 , n2031 , n34948 );
    nor g25798 ( n1348 , n29077 , n17347 );
    not g25799 ( n18891 , n13510 );
    or g25800 ( n29442 , n21095 , n8075 );
    or g25801 ( n34200 , n1507 , n29430 );
    and g25802 ( n40801 , n21537 , n30393 );
    not g25803 ( n5945 , n9206 );
    and g25804 ( n40274 , n23918 , n858 );
    or g25805 ( n22260 , n11307 , n34739 );
    or g25806 ( n25159 , n3930 , n16536 );
    xnor g25807 ( n68 , n10078 , n36186 );
    nor g25808 ( n27806 , n1219 , n40602 );
    not g25809 ( n4732 , n23980 );
    or g25810 ( n15032 , n40978 , n41102 );
    or g25811 ( n23392 , n12383 , n21219 );
    or g25812 ( n29148 , n26354 , n24431 );
    and g25813 ( n13828 , n31568 , n28922 );
    or g25814 ( n27077 , n15577 , n16879 );
    nor g25815 ( n712 , n14471 , n24864 );
    not g25816 ( n11431 , n4165 );
    or g25817 ( n13621 , n35637 , n22912 );
    or g25818 ( n32875 , n13766 , n32980 );
    and g25819 ( n16666 , n26445 , n20101 );
    nor g25820 ( n41740 , n7197 , n41871 );
    or g25821 ( n5233 , n40554 , n20354 );
    xnor g25822 ( n16729 , n23209 , n4226 );
    nor g25823 ( n36136 , n35193 , n24714 );
    or g25824 ( n12689 , n38781 , n36041 );
    not g25825 ( n16466 , n40686 );
    not g25826 ( n10313 , n4354 );
    xnor g25827 ( n35113 , n30139 , n9470 );
    and g25828 ( n21399 , n14730 , n18200 );
    and g25829 ( n34430 , n6259 , n18582 );
    or g25830 ( n21801 , n34997 , n28572 );
    nor g25831 ( n6817 , n27265 , n15358 );
    or g25832 ( n42145 , n14501 , n7053 );
    or g25833 ( n12922 , n19523 , n27645 );
    xnor g25834 ( n6266 , n7922 , n24693 );
    not g25835 ( n15780 , n4999 );
    not g25836 ( n37451 , n33854 );
    not g25837 ( n34429 , n25630 );
    and g25838 ( n30894 , n21988 , n288 );
    xnor g25839 ( n41063 , n23330 , n40477 );
    not g25840 ( n28377 , n34030 );
    and g25841 ( n36320 , n7142 , n24 );
    nor g25842 ( n25862 , n1255 , n5794 );
    xnor g25843 ( n549 , n23322 , n9908 );
    not g25844 ( n5643 , n25069 );
    or g25845 ( n24085 , n17084 , n11510 );
    and g25846 ( n1586 , n12919 , n30289 );
    not g25847 ( n20090 , n33011 );
    or g25848 ( n33459 , n29585 , n40554 );
    or g25849 ( n28496 , n18228 , n16138 );
    and g25850 ( n28646 , n31342 , n4383 );
    or g25851 ( n7713 , n19241 , n10364 );
    or g25852 ( n32012 , n15296 , n15095 );
    or g25853 ( n31225 , n734 , n22512 );
    and g25854 ( n34194 , n9337 , n2123 );
    and g25855 ( n19348 , n35047 , n37459 );
    and g25856 ( n29757 , n20963 , n16612 );
    or g25857 ( n7607 , n40773 , n10696 );
    and g25858 ( n11574 , n36388 , n37820 );
    not g25859 ( n32542 , n9051 );
    or g25860 ( n36705 , n16304 , n24832 );
    not g25861 ( n18393 , n25994 );
    and g25862 ( n36000 , n19684 , n37876 );
    or g25863 ( n11155 , n23510 , n10330 );
    nor g25864 ( n8415 , n34114 , n23174 );
    not g25865 ( n35348 , n19656 );
    not g25866 ( n19493 , n17549 );
    not g25867 ( n26875 , n18228 );
    nor g25868 ( n31652 , n14101 , n41248 );
    xnor g25869 ( n28808 , n41013 , n24157 );
    and g25870 ( n25505 , n18012 , n40843 );
    or g25871 ( n25199 , n19482 , n41590 );
    or g25872 ( n2720 , n20730 , n29856 );
    xnor g25873 ( n27953 , n10913 , n14707 );
    nor g25874 ( n21304 , n37127 , n35484 );
    not g25875 ( n21246 , n18792 );
    nor g25876 ( n28526 , n18866 , n9848 );
    nor g25877 ( n25175 , n27971 , n27906 );
    xnor g25878 ( n41774 , n35741 , n12760 );
    or g25879 ( n37541 , n25466 , n14459 );
    and g25880 ( n34459 , n19914 , n976 );
    and g25881 ( n37938 , n19429 , n35683 );
    or g25882 ( n3756 , n25589 , n29518 );
    xnor g25883 ( n864 , n17652 , n14605 );
    xnor g25884 ( n13780 , n9848 , n18866 );
    nor g25885 ( n826 , n42617 , n15433 );
    and g25886 ( n20877 , n6914 , n11176 );
    xnor g25887 ( n9533 , n28377 , n39306 );
    xnor g25888 ( n10980 , n20850 , n24175 );
    nor g25889 ( n38417 , n41534 , n40449 );
    xnor g25890 ( n38932 , n9619 , n8297 );
    or g25891 ( n39516 , n1289 , n37007 );
    or g25892 ( n35341 , n37616 , n41977 );
    xnor g25893 ( n2715 , n31188 , n30164 );
    xnor g25894 ( n12145 , n34875 , n33930 );
    or g25895 ( n39230 , n6370 , n16772 );
    and g25896 ( n24038 , n37998 , n2621 );
    not g25897 ( n23004 , n5337 );
    or g25898 ( n16978 , n24055 , n28883 );
    not g25899 ( n4165 , n21197 );
    xnor g25900 ( n39440 , n36998 , n4338 );
    and g25901 ( n9238 , n7033 , n9099 );
    not g25902 ( n14863 , n4502 );
    nor g25903 ( n32189 , n2566 , n39777 );
    or g25904 ( n6879 , n34565 , n30251 );
    xnor g25905 ( n18836 , n33706 , n37395 );
    not g25906 ( n37535 , n26351 );
    xnor g25907 ( n16376 , n17476 , n13889 );
    and g25908 ( n18857 , n11788 , n33189 );
    or g25909 ( n36223 , n38142 , n18590 );
    nor g25910 ( n33245 , n29782 , n40043 );
    and g25911 ( n40934 , n39863 , n19685 );
    and g25912 ( n18332 , n26763 , n34971 );
    or g25913 ( n7968 , n782 , n34345 );
    nor g25914 ( n30847 , n10598 , n7465 );
    and g25915 ( n39850 , n3850 , n35576 );
    or g25916 ( n7978 , n10029 , n38456 );
    or g25917 ( n35498 , n20771 , n23732 );
    xnor g25918 ( n25337 , n11220 , n4132 );
    not g25919 ( n7381 , n5196 );
    or g25920 ( n35290 , n4043 , n7557 );
    xnor g25921 ( n31878 , n16297 , n20348 );
    or g25922 ( n31517 , n17950 , n27385 );
    and g25923 ( n5150 , n1229 , n2163 );
    or g25924 ( n36923 , n9844 , n22520 );
    or g25925 ( n24974 , n26071 , n17383 );
    not g25926 ( n32003 , n12132 );
    xnor g25927 ( n22546 , n41013 , n1610 );
    and g25928 ( n38665 , n7718 , n37320 );
    not g25929 ( n6001 , n21787 );
    not g25930 ( n25597 , n11541 );
    xnor g25931 ( n14035 , n4974 , n16071 );
    nor g25932 ( n32025 , n32895 , n31220 );
    or g25933 ( n21056 , n35414 , n24569 );
    nor g25934 ( n40101 , n36667 , n16892 );
    not g25935 ( n3580 , n20832 );
    or g25936 ( n35520 , n38779 , n16627 );
    xnor g25937 ( n16857 , n39178 , n39902 );
    or g25938 ( n42888 , n18622 , n5992 );
    or g25939 ( n16090 , n7551 , n21033 );
    or g25940 ( n38831 , n1806 , n1677 );
    or g25941 ( n16034 , n28634 , n19066 );
    and g25942 ( n4233 , n15618 , n35189 );
    or g25943 ( n19040 , n5964 , n13396 );
    not g25944 ( n2903 , n21998 );
    or g25945 ( n15492 , n34569 , n30390 );
    not g25946 ( n16735 , n21318 );
    xnor g25947 ( n20238 , n42064 , n40004 );
    or g25948 ( n42789 , n7668 , n41724 );
    or g25949 ( n37929 , n32372 , n7928 );
    or g25950 ( n11895 , n28210 , n17576 );
    or g25951 ( n8672 , n16947 , n28562 );
    and g25952 ( n3508 , n1606 , n27696 );
    or g25953 ( n12200 , n33027 , n18515 );
    not g25954 ( n29296 , n29474 );
    or g25955 ( n6060 , n22428 , n8778 );
    not g25956 ( n41084 , n22316 );
    or g25957 ( n23734 , n11909 , n23225 );
    nor g25958 ( n40507 , n9235 , n6178 );
    nor g25959 ( n4875 , n5605 , n18747 );
    or g25960 ( n27288 , n13212 , n32676 );
    not g25961 ( n14275 , n6437 );
    nor g25962 ( n26652 , n34565 , n22146 );
    xnor g25963 ( n42488 , n25211 , n5032 );
    xnor g25964 ( n14979 , n35154 , n35115 );
    or g25965 ( n7733 , n2496 , n23051 );
    or g25966 ( n29392 , n9319 , n249 );
    or g25967 ( n9890 , n19375 , n2802 );
    not g25968 ( n13945 , n37672 );
    or g25969 ( n38159 , n3696 , n27761 );
    and g25970 ( n5508 , n22741 , n5010 );
    or g25971 ( n30246 , n12614 , n39697 );
    xnor g25972 ( n16960 , n6861 , n29231 );
    or g25973 ( n36248 , n5330 , n12290 );
    or g25974 ( n41170 , n5904 , n13532 );
    not g25975 ( n30798 , n33638 );
    xnor g25976 ( n25578 , n28637 , n14212 );
    nor g25977 ( n5942 , n19282 , n3327 );
    not g25978 ( n22242 , n27656 );
    or g25979 ( n25032 , n11186 , n31025 );
    not g25980 ( n11440 , n34323 );
    and g25981 ( n36954 , n21818 , n3717 );
    not g25982 ( n589 , n3209 );
    or g25983 ( n21101 , n42323 , n42899 );
    xnor g25984 ( n23131 , n23061 , n11481 );
    or g25985 ( n37200 , n7020 , n8383 );
    not g25986 ( n40624 , n12857 );
    or g25987 ( n8426 , n17075 , n3410 );
    or g25988 ( n30944 , n8726 , n39072 );
    or g25989 ( n22324 , n9748 , n17222 );
    xnor g25990 ( n17782 , n6625 , n31428 );
    or g25991 ( n12883 , n18634 , n32796 );
    xnor g25992 ( n22492 , n3139 , n39023 );
    or g25993 ( n37023 , n20955 , n41862 );
    and g25994 ( n38783 , n6134 , n827 );
    or g25995 ( n34494 , n31907 , n5258 );
    or g25996 ( n28017 , n42280 , n12867 );
    not g25997 ( n34821 , n18429 );
    nor g25998 ( n18402 , n8769 , n37794 );
    and g25999 ( n6293 , n28303 , n32066 );
    and g26000 ( n3888 , n27619 , n17841 );
    or g26001 ( n24593 , n14454 , n40164 );
    and g26002 ( n15604 , n19076 , n4710 );
    not g26003 ( n16848 , n13106 );
    not g26004 ( n41668 , n12709 );
    not g26005 ( n22942 , n34143 );
    and g26006 ( n15848 , n42435 , n26821 );
    xnor g26007 ( n28396 , n12605 , n7884 );
    nor g26008 ( n7981 , n17049 , n34632 );
    and g26009 ( n32372 , n11671 , n37049 );
    nor g26010 ( n33149 , n21153 , n16122 );
    xnor g26011 ( n31088 , n14096 , n1988 );
    or g26012 ( n4242 , n7897 , n42734 );
    not g26013 ( n7212 , n36909 );
    or g26014 ( n21482 , n19235 , n30413 );
    or g26015 ( n23688 , n13368 , n5529 );
    nor g26016 ( n6533 , n28710 , n30064 );
    not g26017 ( n34212 , n26321 );
    not g26018 ( n4249 , n14190 );
    and g26019 ( n33049 , n30557 , n38231 );
    and g26020 ( n16227 , n6150 , n13365 );
    or g26021 ( n14024 , n26638 , n3728 );
    xnor g26022 ( n31309 , n41826 , n40002 );
    not g26023 ( n15956 , n24716 );
    xnor g26024 ( n17859 , n39053 , n10148 );
    or g26025 ( n34572 , n23739 , n20565 );
    not g26026 ( n16671 , n21606 );
    and g26027 ( n40074 , n21238 , n31414 );
    xnor g26028 ( n32940 , n40320 , n22304 );
    or g26029 ( n3540 , n39910 , n27455 );
    not g26030 ( n25078 , n1853 );
    or g26031 ( n29663 , n8638 , n20773 );
    and g26032 ( n1164 , n24562 , n36985 );
    and g26033 ( n13746 , n25080 , n1593 );
    not g26034 ( n9774 , n4309 );
    nor g26035 ( n28784 , n22482 , n14448 );
    nor g26036 ( n33185 , n5230 , n16036 );
    nor g26037 ( n34227 , n41671 , n30966 );
    or g26038 ( n18538 , n14260 , n17229 );
    nor g26039 ( n1440 , n39739 , n6647 );
    xnor g26040 ( n27886 , n6861 , n26887 );
    or g26041 ( n42628 , n36560 , n40461 );
    not g26042 ( n33095 , n33559 );
    or g26043 ( n33932 , n30739 , n22005 );
    and g26044 ( n13549 , n41212 , n11810 );
    or g26045 ( n1646 , n21481 , n13566 );
    or g26046 ( n7938 , n23221 , n39991 );
    or g26047 ( n447 , n25009 , n15703 );
    and g26048 ( n39337 , n19804 , n5608 );
    not g26049 ( n41505 , n18705 );
    and g26050 ( n8375 , n22656 , n40189 );
    and g26051 ( n42039 , n20080 , n8782 );
    or g26052 ( n8028 , n39327 , n22487 );
    or g26053 ( n16072 , n40322 , n23375 );
    nor g26054 ( n8774 , n13218 , n11366 );
    and g26055 ( n15854 , n30506 , n34438 );
    and g26056 ( n18915 , n30344 , n7891 );
    nor g26057 ( n547 , n26680 , n28128 );
    and g26058 ( n2811 , n9631 , n33327 );
    or g26059 ( n31245 , n17876 , n22858 );
    or g26060 ( n3568 , n14481 , n8444 );
    nor g26061 ( n27512 , n39590 , n27635 );
    or g26062 ( n31602 , n41197 , n4356 );
    xnor g26063 ( n24252 , n41013 , n14949 );
    or g26064 ( n14220 , n11299 , n12768 );
    not g26065 ( n14746 , n20980 );
    not g26066 ( n4909 , n11186 );
    xnor g26067 ( n32427 , n36557 , n18212 );
    xnor g26068 ( n32008 , n27675 , n38879 );
    or g26069 ( n24204 , n29282 , n7244 );
    nor g26070 ( n6311 , n32453 , n1430 );
    xnor g26071 ( n35922 , n39456 , n34974 );
    or g26072 ( n3199 , n36623 , n35441 );
    xnor g26073 ( n34822 , n8837 , n38833 );
    or g26074 ( n1830 , n28788 , n38884 );
    and g26075 ( n9048 , n28026 , n38812 );
    or g26076 ( n10883 , n26168 , n34473 );
    not g26077 ( n12152 , n28403 );
    or g26078 ( n22026 , n41318 , n31918 );
    xnor g26079 ( n34118 , n31857 , n23641 );
    not g26080 ( n9783 , n40225 );
    or g26081 ( n4681 , n5201 , n17230 );
    xnor g26082 ( n10689 , n4124 , n17744 );
    xnor g26083 ( n17603 , n31474 , n40732 );
    nor g26084 ( n624 , n4345 , n10048 );
    nor g26085 ( n33907 , n27994 , n24213 );
    nor g26086 ( n18905 , n10902 , n779 );
    and g26087 ( n16507 , n41364 , n33016 );
    xnor g26088 ( n38914 , n19282 , n30007 );
    or g26089 ( n8629 , n6701 , n23225 );
    or g26090 ( n7964 , n5419 , n11790 );
    or g26091 ( n30015 , n39505 , n41990 );
    and g26092 ( n1900 , n27694 , n33784 );
    xnor g26093 ( n18200 , n13464 , n5964 );
    xnor g26094 ( n23360 , n31989 , n15832 );
    or g26095 ( n25834 , n6085 , n29361 );
    xnor g26096 ( n37356 , n34875 , n38021 );
    or g26097 ( n19827 , n31261 , n16556 );
    or g26098 ( n4215 , n33597 , n36619 );
    not g26099 ( n19355 , n40734 );
    xnor g26100 ( n35033 , n24579 , n2706 );
    nor g26101 ( n20787 , n8167 , n34861 );
    nor g26102 ( n8538 , n27898 , n11883 );
    xnor g26103 ( n27378 , n13038 , n39052 );
    and g26104 ( n19616 , n38971 , n11733 );
    or g26105 ( n15223 , n37671 , n24539 );
    or g26106 ( n27728 , n26987 , n14237 );
    or g26107 ( n675 , n5978 , n28854 );
    and g26108 ( n18635 , n15132 , n25493 );
    or g26109 ( n26979 , n21096 , n16437 );
    not g26110 ( n35133 , n18417 );
    and g26111 ( n4086 , n24914 , n42473 );
    xnor g26112 ( n33876 , n19045 , n2190 );
    or g26113 ( n5008 , n6973 , n10987 );
    or g26114 ( n34067 , n5113 , n27663 );
    and g26115 ( n28701 , n1111 , n2747 );
    xnor g26116 ( n42200 , n34352 , n9840 );
    nor g26117 ( n876 , n32539 , n3595 );
    xnor g26118 ( n32181 , n2950 , n19732 );
    or g26119 ( n4314 , n3664 , n23334 );
    nor g26120 ( n26273 , n18795 , n12447 );
    and g26121 ( n25127 , n11110 , n2398 );
    xnor g26122 ( n39782 , n34352 , n2807 );
    nor g26123 ( n25906 , n27758 , n34495 );
    xnor g26124 ( n27247 , n38886 , n37641 );
    nor g26125 ( n20824 , n36346 , n15856 );
    or g26126 ( n39990 , n4535 , n10719 );
    xnor g26127 ( n21648 , n3549 , n13814 );
    and g26128 ( n41710 , n42853 , n22662 );
    and g26129 ( n29738 , n42348 , n37491 );
    or g26130 ( n25184 , n36844 , n21679 );
    or g26131 ( n6793 , n37031 , n34632 );
    or g26132 ( n26405 , n510 , n14688 );
    not g26133 ( n4166 , n5864 );
    and g26134 ( n14398 , n22425 , n34702 );
    xnor g26135 ( n15194 , n24165 , n12633 );
    and g26136 ( n9494 , n4610 , n6090 );
    or g26137 ( n3326 , n7539 , n4249 );
    nor g26138 ( n14032 , n29395 , n30859 );
    not g26139 ( n4717 , n14008 );
    or g26140 ( n4224 , n9847 , n20600 );
    xnor g26141 ( n24834 , n30103 , n2511 );
    not g26142 ( n1387 , n26925 );
    and g26143 ( n3749 , n19109 , n19050 );
    and g26144 ( n37913 , n26682 , n10401 );
    or g26145 ( n15422 , n40485 , n14130 );
    or g26146 ( n37732 , n33810 , n37674 );
    nor g26147 ( n27389 , n31158 , n3286 );
    or g26148 ( n4794 , n15374 , n20263 );
    and g26149 ( n40602 , n6055 , n26966 );
    not g26150 ( n18024 , n32371 );
    nor g26151 ( n24394 , n3663 , n26847 );
    and g26152 ( n5552 , n3792 , n16755 );
    or g26153 ( n14121 , n25406 , n28214 );
    xnor g26154 ( n12715 , n38658 , n14707 );
    nor g26155 ( n10493 , n8494 , n13786 );
    or g26156 ( n10988 , n14945 , n34119 );
    or g26157 ( n38133 , n8494 , n34906 );
    not g26158 ( n15884 , n26234 );
    not g26159 ( n41604 , n10399 );
    and g26160 ( n38223 , n21775 , n19593 );
    not g26161 ( n7459 , n28195 );
    not g26162 ( n6478 , n24108 );
    or g26163 ( n30149 , n31632 , n8688 );
    xnor g26164 ( n30562 , n40 , n3116 );
    not g26165 ( n9682 , n37760 );
    or g26166 ( n29741 , n9040 , n33287 );
    xnor g26167 ( n19581 , n37436 , n22744 );
    and g26168 ( n38239 , n22679 , n36970 );
    xnor g26169 ( n34685 , n10585 , n546 );
    or g26170 ( n14408 , n22404 , n35695 );
    or g26171 ( n14525 , n16809 , n14641 );
    and g26172 ( n18885 , n17004 , n21851 );
    or g26173 ( n11351 , n7207 , n26855 );
    and g26174 ( n20623 , n11429 , n9899 );
    nor g26175 ( n13075 , n9367 , n8158 );
    or g26176 ( n24256 , n19753 , n14908 );
    not g26177 ( n30150 , n25437 );
    and g26178 ( n32781 , n32506 , n2855 );
    and g26179 ( n28262 , n36487 , n12246 );
    or g26180 ( n32052 , n3487 , n5190 );
    xnor g26181 ( n30275 , n11295 , n853 );
    nor g26182 ( n28946 , n28575 , n11767 );
    or g26183 ( n5710 , n30298 , n42536 );
    not g26184 ( n36514 , n10707 );
    or g26185 ( n29810 , n40114 , n24235 );
    and g26186 ( n20424 , n24525 , n5405 );
    xnor g26187 ( n19705 , n30400 , n16160 );
    nor g26188 ( n32844 , n25273 , n4096 );
    nor g26189 ( n32163 , n27593 , n7213 );
    xnor g26190 ( n32979 , n15051 , n6467 );
    or g26191 ( n31093 , n13726 , n30538 );
    nor g26192 ( n39199 , n27627 , n6467 );
    and g26193 ( n13273 , n33850 , n42285 );
    xnor g26194 ( n21946 , n31099 , n12258 );
    xnor g26195 ( n9698 , n27334 , n488 );
    or g26196 ( n11336 , n14112 , n15070 );
    not g26197 ( n19592 , n36372 );
    xnor g26198 ( n8660 , n31989 , n9710 );
    and g26199 ( n33197 , n18439 , n27864 );
    or g26200 ( n10656 , n23736 , n26079 );
    or g26201 ( n37320 , n18916 , n31727 );
    or g26202 ( n15876 , n19523 , n20004 );
    nor g26203 ( n21049 , n23572 , n19284 );
    and g26204 ( n7740 , n8537 , n10074 );
    or g26205 ( n5072 , n3036 , n38200 );
    or g26206 ( n6700 , n14707 , n4987 );
    or g26207 ( n3086 , n36515 , n21772 );
    not g26208 ( n16693 , n34292 );
    not g26209 ( n24547 , n20072 );
    not g26210 ( n39531 , n18285 );
    or g26211 ( n39684 , n33330 , n19852 );
    not g26212 ( n6132 , n23948 );
    and g26213 ( n26502 , n5339 , n17757 );
    and g26214 ( n4356 , n2638 , n40681 );
    and g26215 ( n13469 , n34251 , n18560 );
    not g26216 ( n20379 , n32661 );
    or g26217 ( n42032 , n13299 , n14635 );
    or g26218 ( n19654 , n29276 , n10207 );
    or g26219 ( n21897 , n24621 , n33453 );
    or g26220 ( n29570 , n20700 , n25780 );
    or g26221 ( n6497 , n22859 , n15676 );
    and g26222 ( n28195 , n33731 , n9744 );
    or g26223 ( n6323 , n3313 , n37777 );
    xnor g26224 ( n20539 , n32632 , n39131 );
    or g26225 ( n21964 , n29521 , n39481 );
    or g26226 ( n33641 , n8626 , n23751 );
    not g26227 ( n3546 , n91 );
    not g26228 ( n14743 , n25883 );
    xnor g26229 ( n12829 , n16547 , n34699 );
    or g26230 ( n27564 , n7857 , n19191 );
    or g26231 ( n26920 , n42811 , n37723 );
    or g26232 ( n40402 , n24658 , n30635 );
    nor g26233 ( n40340 , n3656 , n27193 );
    not g26234 ( n8585 , n4445 );
    xnor g26235 ( n15761 , n41013 , n16426 );
    or g26236 ( n26649 , n26870 , n1576 );
    not g26237 ( n34485 , n42710 );
    or g26238 ( n39417 , n21373 , n20659 );
    nor g26239 ( n42316 , n41629 , n8662 );
    xnor g26240 ( n42326 , n3053 , n42840 );
    or g26241 ( n32286 , n30896 , n5440 );
    or g26242 ( n14425 , n2025 , n12789 );
    or g26243 ( n34983 , n26786 , n7852 );
    and g26244 ( n17353 , n14419 , n4001 );
    xnor g26245 ( n19874 , n41013 , n12417 );
    or g26246 ( n34206 , n30094 , n5818 );
    or g26247 ( n7875 , n7512 , n9983 );
    and g26248 ( n42308 , n1218 , n17863 );
    and g26249 ( n30824 , n12269 , n14514 );
    not g26250 ( n42266 , n30247 );
    and g26251 ( n31254 , n22055 , n8987 );
    not g26252 ( n12226 , n34931 );
    or g26253 ( n923 , n22289 , n37634 );
    and g26254 ( n18770 , n40910 , n3650 );
    and g26255 ( n26340 , n4652 , n12580 );
    or g26256 ( n7709 , n31522 , n31881 );
    and g26257 ( n15013 , n20327 , n30876 );
    or g26258 ( n34966 , n15015 , n25735 );
    or g26259 ( n33247 , n27270 , n14934 );
    or g26260 ( n21769 , n32627 , n8828 );
    xnor g26261 ( n24476 , n41053 , n20616 );
    or g26262 ( n22775 , n15527 , n34048 );
    not g26263 ( n21018 , n35962 );
    nor g26264 ( n36380 , n25588 , n39849 );
    or g26265 ( n31147 , n10717 , n1292 );
    not g26266 ( n21877 , n38898 );
    or g26267 ( n36149 , n2519 , n4607 );
    or g26268 ( n24716 , n683 , n14062 );
    xnor g26269 ( n31849 , n15843 , n33789 );
    not g26270 ( n7196 , n22312 );
    or g26271 ( n7412 , n42396 , n42786 );
    nor g26272 ( n29551 , n38314 , n2258 );
    not g26273 ( n17922 , n42654 );
    or g26274 ( n37629 , n16682 , n40844 );
    not g26275 ( n16243 , n10292 );
    and g26276 ( n14351 , n40013 , n27094 );
    or g26277 ( n38451 , n38157 , n42732 );
    nor g26278 ( n37737 , n15613 , n27805 );
    or g26279 ( n27755 , n17827 , n15011 );
    not g26280 ( n17320 , n37792 );
    xnor g26281 ( n27750 , n378 , n19354 );
    and g26282 ( n6505 , n34047 , n36736 );
    not g26283 ( n29455 , n8569 );
    and g26284 ( n31046 , n7943 , n41568 );
    not g26285 ( n17990 , n5129 );
    nor g26286 ( n14350 , n8494 , n34863 );
    not g26287 ( n28912 , n18746 );
    and g26288 ( n28134 , n21674 , n11281 );
    not g26289 ( n15325 , n22777 );
    xnor g26290 ( n11618 , n5975 , n1655 );
    and g26291 ( n21938 , n11646 , n2925 );
    or g26292 ( n18646 , n7242 , n33696 );
    or g26293 ( n25527 , n1917 , n36082 );
    or g26294 ( n32537 , n16226 , n31527 );
    or g26295 ( n31608 , n11976 , n29016 );
    and g26296 ( n29630 , n12746 , n31618 );
    or g26297 ( n23152 , n35166 , n23694 );
    or g26298 ( n2872 , n13470 , n22701 );
    and g26299 ( n26260 , n15488 , n25791 );
    and g26300 ( n7765 , n14255 , n24144 );
    or g26301 ( n12767 , n40434 , n39433 );
    xnor g26302 ( n40068 , n12781 , n17457 );
    and g26303 ( n26637 , n3791 , n16766 );
    xnor g26304 ( n1524 , n4055 , n34219 );
    not g26305 ( n28028 , n9654 );
    not g26306 ( n4467 , n27419 );
    nor g26307 ( n28281 , n12104 , n5197 );
    nor g26308 ( n38464 , n4443 , n25106 );
    not g26309 ( n9418 , n36627 );
    nor g26310 ( n21533 , n3769 , n30715 );
    nor g26311 ( n4560 , n22437 , n42017 );
    xnor g26312 ( n9118 , n28120 , n11443 );
    or g26313 ( n32550 , n39292 , n7469 );
    not g26314 ( n2279 , n4178 );
    and g26315 ( n27306 , n41010 , n17323 );
    and g26316 ( n41466 , n34454 , n8492 );
    not g26317 ( n29715 , n13054 );
    xnor g26318 ( n10594 , n20557 , n4803 );
    or g26319 ( n21441 , n12562 , n11134 );
    or g26320 ( n16940 , n39416 , n10953 );
    xnor g26321 ( n18995 , n6625 , n38740 );
    xnor g26322 ( n348 , n21559 , n33824 );
    xnor g26323 ( n18526 , n1622 , n42243 );
    not g26324 ( n34165 , n17088 );
    or g26325 ( n5034 , n15095 , n34063 );
    and g26326 ( n41213 , n27286 , n16042 );
    or g26327 ( n4761 , n2043 , n1687 );
    and g26328 ( n9609 , n3833 , n4626 );
    or g26329 ( n9571 , n3879 , n34925 );
    not g26330 ( n13995 , n19571 );
    or g26331 ( n26364 , n10212 , n8304 );
    not g26332 ( n14420 , n27925 );
    or g26333 ( n28871 , n11902 , n20663 );
    and g26334 ( n18868 , n17029 , n19031 );
    xnor g26335 ( n36577 , n38777 , n17181 );
    and g26336 ( n6346 , n34272 , n10062 );
    or g26337 ( n33146 , n35366 , n27455 );
    or g26338 ( n22331 , n30185 , n32967 );
    xnor g26339 ( n41671 , n25884 , n21205 );
    not g26340 ( n4561 , n25105 );
    and g26341 ( n7668 , n33732 , n2953 );
    nor g26342 ( n6043 , n19164 , n15265 );
    or g26343 ( n33565 , n41773 , n10418 );
    or g26344 ( n2057 , n4702 , n29077 );
    or g26345 ( n30927 , n40738 , n30117 );
    or g26346 ( n41087 , n35450 , n9521 );
    nor g26347 ( n23787 , n408 , n22162 );
    and g26348 ( n17432 , n18713 , n37406 );
    and g26349 ( n27050 , n23002 , n30997 );
    nor g26350 ( n29016 , n36341 , n35676 );
    or g26351 ( n27747 , n1814 , n25429 );
    xnor g26352 ( n36053 , n25884 , n17943 );
    or g26353 ( n458 , n39461 , n3993 );
    or g26354 ( n41492 , n30867 , n25303 );
    not g26355 ( n4712 , n246 );
    or g26356 ( n25408 , n9445 , n24607 );
    nor g26357 ( n4318 , n21407 , n10600 );
    not g26358 ( n6628 , n16079 );
    not g26359 ( n22312 , n1794 );
    nor g26360 ( n4965 , n21652 , n31579 );
    and g26361 ( n38993 , n6499 , n33868 );
    and g26362 ( n15550 , n29837 , n18671 );
    xnor g26363 ( n35367 , n10834 , n4336 );
    xnor g26364 ( n33070 , n11383 , n12084 );
    and g26365 ( n33041 , n7343 , n5687 );
    or g26366 ( n15585 , n22991 , n16429 );
    or g26367 ( n20861 , n35772 , n37117 );
    and g26368 ( n28757 , n31024 , n17562 );
    not g26369 ( n15619 , n33343 );
    or g26370 ( n32387 , n40210 , n33197 );
    xnor g26371 ( n18030 , n28614 , n37690 );
    or g26372 ( n24988 , n33291 , n626 );
    nor g26373 ( n40914 , n23770 , n32843 );
    and g26374 ( n36253 , n39655 , n30107 );
    and g26375 ( n10582 , n15825 , n25565 );
    or g26376 ( n29387 , n17654 , n21557 );
    and g26377 ( n38326 , n1089 , n8224 );
    and g26378 ( n23144 , n24860 , n14132 );
    nor g26379 ( n29405 , n6503 , n8571 );
    xnor g26380 ( n21451 , n29113 , n11495 );
    not g26381 ( n2093 , n9174 );
    nor g26382 ( n14500 , n15237 , n40219 );
    or g26383 ( n5745 , n27612 , n40652 );
    nor g26384 ( n42001 , n3704 , n23057 );
    or g26385 ( n31486 , n19609 , n42207 );
    and g26386 ( n29998 , n9773 , n37497 );
    or g26387 ( n31621 , n24690 , n40775 );
    or g26388 ( n5569 , n32230 , n26944 );
    or g26389 ( n9096 , n1933 , n28158 );
    or g26390 ( n42846 , n15493 , n17104 );
    or g26391 ( n16384 , n10576 , n19193 );
    not g26392 ( n38438 , n37434 );
    or g26393 ( n10884 , n36216 , n40486 );
    xnor g26394 ( n34063 , n33405 , n33524 );
    xnor g26395 ( n22233 , n18859 , n9799 );
    xnor g26396 ( n12223 , n5891 , n4824 );
    not g26397 ( n4670 , n42154 );
    and g26398 ( n21860 , n26011 , n42199 );
    not g26399 ( n18807 , n17516 );
    and g26400 ( n34172 , n40788 , n7101 );
    nor g26401 ( n33213 , n20067 , n13552 );
    not g26402 ( n39368 , n38288 );
    and g26403 ( n24770 , n3899 , n3174 );
    xnor g26404 ( n40585 , n11436 , n2838 );
    nor g26405 ( n21624 , n32376 , n35721 );
    not g26406 ( n36689 , n34103 );
    xnor g26407 ( n1319 , n33222 , n37047 );
    or g26408 ( n10159 , n13423 , n18965 );
    xnor g26409 ( n22025 , n15266 , n11782 );
    not g26410 ( n30652 , n34880 );
    not g26411 ( n440 , n2298 );
    or g26412 ( n16561 , n10313 , n21237 );
    nor g26413 ( n7430 , n6490 , n26115 );
    xnor g26414 ( n1667 , n7443 , n28924 );
    or g26415 ( n23086 , n18789 , n24391 );
    or g26416 ( n14931 , n4018 , n40244 );
    not g26417 ( n16214 , n40458 );
    or g26418 ( n5687 , n35301 , n2844 );
    or g26419 ( n8191 , n3583 , n2667 );
    and g26420 ( n22730 , n30377 , n15566 );
    nor g26421 ( n33986 , n13796 , n26248 );
    and g26422 ( n40884 , n21244 , n1212 );
    or g26423 ( n24178 , n18314 , n38933 );
    and g26424 ( n40625 , n26683 , n4168 );
    or g26425 ( n34635 , n18866 , n552 );
    and g26426 ( n34981 , n30518 , n25375 );
    and g26427 ( n26478 , n36209 , n386 );
    or g26428 ( n11112 , n27667 , n23986 );
    and g26429 ( n10020 , n4503 , n25058 );
    and g26430 ( n24643 , n17632 , n19405 );
    nor g26431 ( n37244 , n14471 , n35045 );
    not g26432 ( n11321 , n11594 );
    xnor g26433 ( n37557 , n4844 , n42688 );
    or g26434 ( n1872 , n27908 , n11582 );
    and g26435 ( n2333 , n9648 , n39004 );
    or g26436 ( n41155 , n15314 , n14054 );
    nor g26437 ( n12628 , n27808 , n2410 );
    or g26438 ( n21281 , n23941 , n34917 );
    or g26439 ( n21768 , n34419 , n18973 );
    not g26440 ( n11225 , n39546 );
    xnor g26441 ( n22 , n19680 , n38202 );
    or g26442 ( n30659 , n15317 , n7167 );
    and g26443 ( n18006 , n512 , n7129 );
    nor g26444 ( n18642 , n10810 , n21257 );
    and g26445 ( n19267 , n14214 , n25491 );
    and g26446 ( n18274 , n27885 , n27100 );
    nor g26447 ( n4900 , n12795 , n16979 );
    xnor g26448 ( n37589 , n29359 , n15494 );
    or g26449 ( n7859 , n23773 , n27761 );
    not g26450 ( n41406 , n32849 );
    or g26451 ( n2421 , n29368 , n10045 );
    or g26452 ( n36465 , n3916 , n35192 );
    or g26453 ( n7158 , n16923 , n28045 );
    and g26454 ( n20474 , n10983 , n37409 );
    nor g26455 ( n11553 , n33687 , n3889 );
    and g26456 ( n27112 , n18794 , n28059 );
    and g26457 ( n15014 , n25327 , n16040 );
    or g26458 ( n25192 , n23604 , n31321 );
    not g26459 ( n5978 , n18584 );
    or g26460 ( n37067 , n19214 , n15317 );
    xnor g26461 ( n2915 , n26579 , n34676 );
    and g26462 ( n20687 , n4172 , n35725 );
    or g26463 ( n23238 , n21268 , n10147 );
    or g26464 ( n32581 , n1441 , n14603 );
    xnor g26465 ( n23197 , n6688 , n15986 );
    nor g26466 ( n21371 , n35471 , n10255 );
    and g26467 ( n27401 , n25220 , n29393 );
    or g26468 ( n36665 , n23202 , n36120 );
    xnor g26469 ( n16063 , n11436 , n15498 );
    or g26470 ( n16820 , n18053 , n15175 );
    or g26471 ( n37710 , n39808 , n6000 );
    or g26472 ( n40518 , n13712 , n15405 );
    and g26473 ( n39802 , n40121 , n33078 );
    not g26474 ( n38835 , n17232 );
    or g26475 ( n3601 , n29942 , n20331 );
    xnor g26476 ( n34298 , n11436 , n34505 );
    and g26477 ( n1815 , n29570 , n34340 );
    and g26478 ( n11673 , n35594 , n40131 );
    nor g26479 ( n9473 , n42792 , n38117 );
    or g26480 ( n41377 , n41812 , n34267 );
    or g26481 ( n26163 , n20250 , n1708 );
    or g26482 ( n35048 , n40710 , n11390 );
    nor g26483 ( n40193 , n26255 , n20560 );
    not g26484 ( n42128 , n35311 );
    and g26485 ( n13337 , n6233 , n28569 );
    or g26486 ( n1401 , n30237 , n4564 );
    or g26487 ( n7090 , n17120 , n19068 );
    nor g26488 ( n4504 , n9030 , n20106 );
    not g26489 ( n23703 , n41759 );
    nor g26490 ( n31563 , n7183 , n16062 );
    and g26491 ( n30091 , n31182 , n9598 );
    and g26492 ( n8389 , n1894 , n17350 );
    and g26493 ( n22764 , n39686 , n30828 );
    and g26494 ( n38548 , n18570 , n24791 );
    or g26495 ( n22760 , n15445 , n10233 );
    nor g26496 ( n21690 , n5320 , n3853 );
    or g26497 ( n24095 , n14581 , n34391 );
    not g26498 ( n269 , n29557 );
    or g26499 ( n30990 , n9238 , n35879 );
    or g26500 ( n27655 , n3945 , n2624 );
    not g26501 ( n20425 , n36025 );
    or g26502 ( n11330 , n113 , n32103 );
    and g26503 ( n18639 , n10339 , n5331 );
    and g26504 ( n35253 , n37670 , n11350 );
    not g26505 ( n25029 , n14524 );
    or g26506 ( n3108 , n32194 , n36301 );
    or g26507 ( n27586 , n7139 , n1408 );
    or g26508 ( n9706 , n19058 , n7898 );
    nor g26509 ( n14519 , n9796 , n28935 );
    or g26510 ( n11176 , n6646 , n29363 );
    not g26511 ( n5002 , n20287 );
    or g26512 ( n7556 , n40830 , n7612 );
    and g26513 ( n8505 , n29159 , n14574 );
    xnor g26514 ( n13183 , n21973 , n29381 );
    nor g26515 ( n40670 , n31105 , n17508 );
    or g26516 ( n16065 , n30838 , n5261 );
    or g26517 ( n35724 , n32204 , n31950 );
    xnor g26518 ( n11528 , n39852 , n3727 );
    and g26519 ( n14848 , n32914 , n6853 );
    not g26520 ( n18224 , n34145 );
    not g26521 ( n25206 , n17195 );
    and g26522 ( n37988 , n8596 , n12411 );
    or g26523 ( n34239 , n14718 , n23711 );
    xnor g26524 ( n4692 , n6841 , n37519 );
    or g26525 ( n30260 , n37044 , n24484 );
    or g26526 ( n25267 , n25929 , n5984 );
    xnor g26527 ( n28636 , n36998 , n2394 );
    or g26528 ( n39160 , n15192 , n22355 );
    or g26529 ( n2966 , n10346 , n30678 );
    or g26530 ( n20146 , n54 , n31164 );
    xnor g26531 ( n19383 , n31054 , n5028 );
    or g26532 ( n6143 , n451 , n33262 );
    or g26533 ( n15157 , n13436 , n12771 );
    or g26534 ( n311 , n1994 , n32815 );
    not g26535 ( n40990 , n1412 );
    or g26536 ( n7332 , n40839 , n1280 );
    nor g26537 ( n42566 , n22877 , n40696 );
    or g26538 ( n36748 , n39804 , n14353 );
    or g26539 ( n7643 , n14622 , n16438 );
    nor g26540 ( n1410 , n35678 , n36787 );
    or g26541 ( n7958 , n17830 , n35656 );
    or g26542 ( n10469 , n22759 , n37578 );
    or g26543 ( n29945 , n29294 , n32923 );
    xnor g26544 ( n24088 , n19186 , n16129 );
    xnor g26545 ( n20206 , n31989 , n17856 );
    not g26546 ( n32779 , n28956 );
    or g26547 ( n7208 , n26647 , n39081 );
    or g26548 ( n37608 , n10284 , n18879 );
    or g26549 ( n10145 , n19535 , n17239 );
    not g26550 ( n11039 , n535 );
    xnor g26551 ( n1601 , n36998 , n7977 );
    or g26552 ( n9522 , n28551 , n20382 );
    nor g26553 ( n37854 , n28120 , n2582 );
    or g26554 ( n9929 , n17871 , n36779 );
    or g26555 ( n41785 , n39032 , n17794 );
    or g26556 ( n33836 , n15185 , n2040 );
    or g26557 ( n460 , n42206 , n14153 );
    xnor g26558 ( n8057 , n31928 , n29197 );
    nor g26559 ( n21004 , n12264 , n32111 );
    xnor g26560 ( n41843 , n39760 , n10879 );
    and g26561 ( n6026 , n18732 , n38709 );
    and g26562 ( n7569 , n13898 , n32504 );
    or g26563 ( n18470 , n37813 , n35431 );
    nor g26564 ( n32972 , n33774 , n35467 );
    or g26565 ( n37895 , n4892 , n5813 );
    nor g26566 ( n13503 , n2717 , n24244 );
    and g26567 ( n3978 , n17662 , n9712 );
    and g26568 ( n6537 , n11290 , n27930 );
    or g26569 ( n28676 , n22297 , n19848 );
    not g26570 ( n31965 , n17275 );
    xnor g26571 ( n34376 , n18558 , n31579 );
    or g26572 ( n33277 , n37559 , n27313 );
    xnor g26573 ( n20439 , n22693 , n10239 );
    xnor g26574 ( n12693 , n4341 , n27047 );
    and g26575 ( n29898 , n22166 , n32577 );
    and g26576 ( n9452 , n6822 , n29107 );
    and g26577 ( n15392 , n14270 , n19246 );
    or g26578 ( n38724 , n40072 , n32912 );
    or g26579 ( n18743 , n23082 , n28186 );
    nor g26580 ( n7452 , n39556 , n13797 );
    or g26581 ( n41554 , n5140 , n12579 );
    or g26582 ( n35598 , n16294 , n7773 );
    nor g26583 ( n14991 , n11251 , n15390 );
    and g26584 ( n28607 , n15086 , n11652 );
    nor g26585 ( n25100 , n20516 , n8237 );
    and g26586 ( n29983 , n34686 , n4096 );
    or g26587 ( n38880 , n4893 , n29018 );
    or g26588 ( n28380 , n6686 , n4539 );
    and g26589 ( n16930 , n35406 , n18154 );
    xnor g26590 ( n21727 , n12836 , n40563 );
    nor g26591 ( n12872 , n8494 , n17187 );
    and g26592 ( n33569 , n28948 , n19044 );
    xnor g26593 ( n31723 , n4385 , n39794 );
    and g26594 ( n9651 , n6704 , n6755 );
    or g26595 ( n22668 , n22705 , n12178 );
    xnor g26596 ( n17615 , n25470 , n36117 );
    or g26597 ( n40553 , n11340 , n38354 );
    or g26598 ( n8767 , n2954 , n11732 );
    not g26599 ( n15572 , n22294 );
    or g26600 ( n14970 , n8094 , n39810 );
    and g26601 ( n22693 , n5076 , n17732 );
    and g26602 ( n10821 , n19513 , n21345 );
    xnor g26603 ( n31988 , n23602 , n8494 );
    and g26604 ( n20189 , n8795 , n2553 );
    or g26605 ( n18423 , n6558 , n24708 );
    nor g26606 ( n28366 , n44 , n36746 );
    and g26607 ( n7725 , n36238 , n6523 );
    and g26608 ( n28765 , n25748 , n27218 );
    xnor g26609 ( n32649 , n32470 , n12718 );
    not g26610 ( n13234 , n12069 );
    and g26611 ( n38940 , n24324 , n22663 );
    nor g26612 ( n17461 , n8346 , n16430 );
    or g26613 ( n20569 , n12692 , n24380 );
    and g26614 ( n5799 , n2475 , n31922 );
    and g26615 ( n21976 , n22938 , n25667 );
    nor g26616 ( n11077 , n33981 , n15690 );
    xnor g26617 ( n35358 , n36197 , n38879 );
    or g26618 ( n14734 , n23509 , n17832 );
    or g26619 ( n27318 , n39839 , n28722 );
    and g26620 ( n13698 , n384 , n25997 );
    xnor g26621 ( n33969 , n38886 , n13115 );
    not g26622 ( n5926 , n10279 );
    or g26623 ( n42864 , n16984 , n2565 );
    xnor g26624 ( n25519 , n34226 , n28471 );
    xnor g26625 ( n20023 , n4334 , n26498 );
    or g26626 ( n23515 , n12700 , n4332 );
    nor g26627 ( n42059 , n39303 , n17630 );
    or g26628 ( n34693 , n9228 , n9975 );
    and g26629 ( n730 , n24393 , n24834 );
    and g26630 ( n7066 , n35215 , n24285 );
    xnor g26631 ( n22745 , n7465 , n10598 );
    nor g26632 ( n18611 , n30343 , n38092 );
    not g26633 ( n5614 , n17080 );
    not g26634 ( n14364 , n4424 );
    xnor g26635 ( n23521 , n21585 , n39321 );
    xnor g26636 ( n41924 , n42091 , n25070 );
    or g26637 ( n23229 , n36689 , n26973 );
    xnor g26638 ( n30406 , n552 , n18866 );
    or g26639 ( n6609 , n28301 , n32686 );
    and g26640 ( n16199 , n1513 , n16976 );
    not g26641 ( n894 , n14209 );
    or g26642 ( n34644 , n37715 , n24011 );
    xnor g26643 ( n40187 , n32470 , n19066 );
    not g26644 ( n23783 , n6889 );
    or g26645 ( n12272 , n12288 , n1735 );
    and g26646 ( n23013 , n33443 , n10323 );
    nor g26647 ( n33513 , n7397 , n41048 );
    or g26648 ( n703 , n34434 , n34320 );
    nor g26649 ( n29459 , n1507 , n26984 );
    or g26650 ( n21678 , n34017 , n13957 );
    or g26651 ( n19335 , n30435 , n18398 );
    or g26652 ( n12820 , n18314 , n19280 );
    and g26653 ( n5565 , n31514 , n36314 );
    nor g26654 ( n17241 , n13921 , n15077 );
    not g26655 ( n34226 , n31352 );
    and g26656 ( n28438 , n17554 , n19543 );
    nor g26657 ( n6965 , n25173 , n21761 );
    or g26658 ( n23854 , n11424 , n38196 );
    or g26659 ( n13602 , n25961 , n10742 );
    xnor g26660 ( n40549 , n36998 , n3569 );
    and g26661 ( n2726 , n29657 , n25678 );
    or g26662 ( n36925 , n42405 , n13835 );
    nor g26663 ( n37623 , n1507 , n4366 );
    nor g26664 ( n423 , n4659 , n2434 );
    or g26665 ( n22085 , n12576 , n18393 );
    or g26666 ( n5300 , n31724 , n4363 );
    nor g26667 ( n7934 , n17120 , n4735 );
    nor g26668 ( n2648 , n42585 , n25029 );
    or g26669 ( n12458 , n10804 , n39108 );
    not g26670 ( n33931 , n20542 );
    and g26671 ( n32056 , n42914 , n346 );
    nor g26672 ( n41975 , n17744 , n33316 );
    and g26673 ( n1063 , n41589 , n3184 );
    or g26674 ( n29238 , n6709 , n5036 );
    and g26675 ( n23042 , n12356 , n7102 );
    nor g26676 ( n2506 , n32682 , n29806 );
    not g26677 ( n16810 , n14089 );
    not g26678 ( n38991 , n22212 );
    not g26679 ( n38427 , n27102 );
    and g26680 ( n7899 , n10293 , n10932 );
    not g26681 ( n2786 , n4854 );
    nor g26682 ( n131 , n42272 , n15869 );
    nor g26683 ( n15222 , n34816 , n41327 );
    xnor g26684 ( n2689 , n9443 , n33981 );
    or g26685 ( n34531 , n23563 , n22018 );
    not g26686 ( n42786 , n38282 );
    or g26687 ( n5536 , n3991 , n10760 );
    and g26688 ( n9239 , n10500 , n34452 );
    nor g26689 ( n4627 , n5964 , n3971 );
    nor g26690 ( n3434 , n33219 , n18052 );
    or g26691 ( n40171 , n32842 , n27319 );
    or g26692 ( n22795 , n154 , n6739 );
    or g26693 ( n34116 , n10684 , n42448 );
    or g26694 ( n19579 , n946 , n33431 );
    or g26695 ( n28321 , n38463 , n20565 );
    xnor g26696 ( n22194 , n2127 , n10241 );
    not g26697 ( n22086 , n40006 );
    and g26698 ( n10533 , n6245 , n23833 );
    or g26699 ( n23529 , n24298 , n888 );
    xnor g26700 ( n23495 , n32470 , n37506 );
    or g26701 ( n15682 , n16497 , n38191 );
    or g26702 ( n33161 , n10737 , n42513 );
    or g26703 ( n4584 , n25004 , n12768 );
    and g26704 ( n7827 , n13693 , n5361 );
    or g26705 ( n35419 , n8064 , n25774 );
    nor g26706 ( n3392 , n15727 , n30897 );
    and g26707 ( n5458 , n12230 , n20353 );
    or g26708 ( n4959 , n15976 , n29833 );
    and g26709 ( n11494 , n11170 , n36152 );
    or g26710 ( n22913 , n18273 , n3856 );
    or g26711 ( n7624 , n31391 , n30713 );
    or g26712 ( n25767 , n28375 , n1688 );
    or g26713 ( n38660 , n20835 , n29985 );
    and g26714 ( n15074 , n24323 , n20636 );
    not g26715 ( n41113 , n35038 );
    not g26716 ( n6246 , n40735 );
    not g26717 ( n2320 , n21439 );
    or g26718 ( n9620 , n25195 , n21404 );
    or g26719 ( n13905 , n30358 , n25179 );
    not g26720 ( n38789 , n33989 );
    nor g26721 ( n4789 , n1224 , n41762 );
    and g26722 ( n41655 , n30706 , n15712 );
    and g26723 ( n11310 , n2385 , n22674 );
    or g26724 ( n26719 , n33643 , n9610 );
    and g26725 ( n22964 , n22226 , n2998 );
    or g26726 ( n27608 , n9040 , n9825 );
    not g26727 ( n36585 , n38721 );
    or g26728 ( n16003 , n34575 , n13490 );
    or g26729 ( n7605 , n29669 , n15762 );
    and g26730 ( n30408 , n12590 , n25741 );
    or g26731 ( n14624 , n21712 , n13495 );
    nor g26732 ( n39411 , n37256 , n8825 );
    xnor g26733 ( n31554 , n9155 , n37711 );
    or g26734 ( n17270 , n36864 , n5227 );
    nor g26735 ( n22035 , n4266 , n36972 );
    or g26736 ( n12903 , n15130 , n28264 );
    and g26737 ( n16350 , n29220 , n14190 );
    or g26738 ( n12611 , n3223 , n418 );
    or g26739 ( n4518 , n36965 , n7289 );
    and g26740 ( n40831 , n29400 , n27202 );
    xnor g26741 ( n38791 , n32734 , n10713 );
    not g26742 ( n28726 , n13851 );
    or g26743 ( n20937 , n42045 , n6493 );
    xnor g26744 ( n27134 , n9619 , n22983 );
    xnor g26745 ( n39053 , n40391 , n6035 );
    not g26746 ( n19810 , n34975 );
    xnor g26747 ( n7032 , n31099 , n31322 );
    and g26748 ( n16611 , n13674 , n23495 );
    not g26749 ( n37779 , n11047 );
    and g26750 ( n18817 , n11293 , n38535 );
    not g26751 ( n4223 , n7358 );
    not g26752 ( n4651 , n34173 );
    not g26753 ( n12655 , n40371 );
    or g26754 ( n37069 , n29844 , n18068 );
    not g26755 ( n20292 , n37681 );
    or g26756 ( n36225 , n26471 , n21772 );
    xnor g26757 ( n22292 , n3514 , n34565 );
    xnor g26758 ( n172 , n15972 , n24197 );
    not g26759 ( n20486 , n55 );
    or g26760 ( n19708 , n10317 , n23286 );
    not g26761 ( n13751 , n3547 );
    and g26762 ( n448 , n16815 , n32562 );
    or g26763 ( n36595 , n7857 , n5141 );
    or g26764 ( n6470 , n18203 , n42357 );
    or g26765 ( n18483 , n33412 , n15762 );
    and g26766 ( n23722 , n14159 , n14158 );
    or g26767 ( n6577 , n20317 , n27385 );
    xnor g26768 ( n2669 , n3713 , n19975 );
    or g26769 ( n12622 , n40109 , n11647 );
    not g26770 ( n38944 , n42666 );
    xnor g26771 ( n72 , n41480 , n21239 );
    not g26772 ( n31997 , n23847 );
    xnor g26773 ( n19879 , n34721 , n18092 );
    xnor g26774 ( n12781 , n35273 , n14471 );
    or g26775 ( n312 , n38795 , n5910 );
    or g26776 ( n26603 , n4717 , n40077 );
    nor g26777 ( n38207 , n2323 , n13305 );
    not g26778 ( n14765 , n42541 );
    or g26779 ( n22665 , n12898 , n16465 );
    not g26780 ( n34641 , n39391 );
    xnor g26781 ( n26227 , n13274 , n15764 );
    or g26782 ( n9111 , n38251 , n4436 );
    xnor g26783 ( n40320 , n35477 , n3690 );
    xnor g26784 ( n33348 , n38712 , n13061 );
    nor g26785 ( n35223 , n2445 , n8083 );
    xnor g26786 ( n809 , n7262 , n15502 );
    or g26787 ( n28588 , n14765 , n16449 );
    not g26788 ( n6688 , n3619 );
    xnor g26789 ( n25609 , n5041 , n2582 );
    or g26790 ( n6799 , n11317 , n28736 );
    and g26791 ( n10965 , n5943 , n40620 );
    not g26792 ( n9146 , n7958 );
    or g26793 ( n7866 , n25784 , n2791 );
    nor g26794 ( n21279 , n37109 , n14640 );
    or g26795 ( n25242 , n16533 , n10063 );
    not g26796 ( n7475 , n1615 );
    or g26797 ( n7228 , n9980 , n42645 );
    xnor g26798 ( n6539 , n15972 , n40304 );
    and g26799 ( n3558 , n25551 , n42831 );
    nor g26800 ( n27679 , n99 , n1406 );
    or g26801 ( n30760 , n1169 , n6510 );
    or g26802 ( n30012 , n20978 , n19909 );
    and g26803 ( n31937 , n31291 , n10481 );
    xnor g26804 ( n4974 , n21192 , n26688 );
    or g26805 ( n11878 , n36621 , n8059 );
    not g26806 ( n34949 , n19578 );
    or g26807 ( n9293 , n41218 , n6500 );
    or g26808 ( n40406 , n27554 , n16718 );
    not g26809 ( n39568 , n31097 );
    not g26810 ( n32526 , n3366 );
    and g26811 ( n17482 , n21022 , n9698 );
    not g26812 ( n27213 , n34885 );
    or g26813 ( n36047 , n15096 , n18683 );
    and g26814 ( n19185 , n37807 , n31968 );
    not g26815 ( n38029 , n20761 );
    and g26816 ( n8312 , n25435 , n22399 );
    or g26817 ( n28580 , n41128 , n32259 );
    or g26818 ( n5452 , n9721 , n12621 );
    nor g26819 ( n1673 , n27483 , n20828 );
    or g26820 ( n31281 , n4545 , n8410 );
    or g26821 ( n12474 , n5208 , n39647 );
    xnor g26822 ( n5786 , n34731 , n35013 );
    not g26823 ( n31724 , n38444 );
    and g26824 ( n14414 , n2842 , n3052 );
    or g26825 ( n25268 , n21836 , n36991 );
    or g26826 ( n5725 , n1507 , n22599 );
    or g26827 ( n23493 , n33027 , n2438 );
    and g26828 ( n13493 , n20551 , n21590 );
    nor g26829 ( n7230 , n3735 , n41216 );
    and g26830 ( n9710 , n5954 , n34055 );
    or g26831 ( n23740 , n28080 , n37110 );
    or g26832 ( n40058 , n26129 , n39423 );
    not g26833 ( n7707 , n15042 );
    or g26834 ( n19900 , n1824 , n36662 );
    or g26835 ( n13258 , n15149 , n29182 );
    and g26836 ( n29900 , n39361 , n8776 );
    or g26837 ( n31971 , n14471 , n3501 );
    and g26838 ( n28848 , n13097 , n29597 );
    or g26839 ( n40425 , n26915 , n18984 );
    or g26840 ( n36598 , n13762 , n756 );
    xnor g26841 ( n21230 , n105 , n3971 );
    and g26842 ( n42450 , n21065 , n39841 );
    or g26843 ( n636 , n2223 , n42620 );
    or g26844 ( n23617 , n14559 , n37793 );
    or g26845 ( n22380 , n7375 , n25329 );
    nor g26846 ( n18323 , n34292 , n29240 );
    not g26847 ( n9137 , n28090 );
    or g26848 ( n28826 , n39908 , n22941 );
    or g26849 ( n12335 , n5756 , n37280 );
    or g26850 ( n33368 , n10149 , n6637 );
    or g26851 ( n38445 , n25377 , n30644 );
    and g26852 ( n3166 , n19514 , n2956 );
    nor g26853 ( n7957 , n23439 , n9728 );
    nor g26854 ( n13590 , n5347 , n20235 );
    not g26855 ( n22713 , n36120 );
    or g26856 ( n7261 , n9225 , n8006 );
    and g26857 ( n17770 , n19546 , n23606 );
    xnor g26858 ( n4549 , n16528 , n14197 );
    xnor g26859 ( n34602 , n21534 , n20049 );
    xnor g26860 ( n14405 , n8210 , n12045 );
    not g26861 ( n29780 , n22500 );
    or g26862 ( n28756 , n31485 , n24189 );
    or g26863 ( n8637 , n14454 , n1345 );
    xnor g26864 ( n3909 , n27398 , n18197 );
    or g26865 ( n30077 , n11148 , n3088 );
    or g26866 ( n6420 , n19275 , n15950 );
    and g26867 ( n5848 , n11345 , n39336 );
    not g26868 ( n27131 , n24079 );
    or g26869 ( n18952 , n26081 , n41207 );
    and g26870 ( n18969 , n20136 , n18609 );
    nor g26871 ( n21985 , n34343 , n40510 );
    or g26872 ( n40382 , n17615 , n12086 );
    nor g26873 ( n24697 , n33160 , n11557 );
    or g26874 ( n27639 , n41498 , n12200 );
    not g26875 ( n29504 , n2424 );
    or g26876 ( n35945 , n7826 , n30903 );
    and g26877 ( n24432 , n40064 , n7403 );
    nor g26878 ( n24017 , n15336 , n41452 );
    not g26879 ( n34816 , n30405 );
    or g26880 ( n9273 , n42113 , n42845 );
    or g26881 ( n36779 , n23745 , n5688 );
    not g26882 ( n35452 , n39921 );
    and g26883 ( n34557 , n32012 , n34124 );
    not g26884 ( n14511 , n12935 );
    and g26885 ( n34962 , n35154 , n10187 );
    nor g26886 ( n17556 , n41419 , n17046 );
    not g26887 ( n4727 , n21971 );
    or g26888 ( n12312 , n2493 , n35529 );
    or g26889 ( n11563 , n1231 , n39040 );
    and g26890 ( n8646 , n12342 , n22612 );
    nor g26891 ( n27448 , n40476 , n8127 );
    and g26892 ( n24260 , n6095 , n2344 );
    xnor g26893 ( n9436 , n10639 , n23450 );
    or g26894 ( n3510 , n27022 , n3781 );
    not g26895 ( n42429 , n12767 );
    or g26896 ( n16519 , n29455 , n37229 );
    or g26897 ( n42322 , n5813 , n22815 );
    or g26898 ( n36520 , n37952 , n24318 );
    or g26899 ( n16725 , n27088 , n11026 );
    xnor g26900 ( n26337 , n30672 , n36117 );
    not g26901 ( n22885 , n18024 );
    xnor g26902 ( n10004 , n30768 , n25146 );
    or g26903 ( n28465 , n6423 , n34557 );
    or g26904 ( n4077 , n545 , n4088 );
    nor g26905 ( n39273 , n1555 , n22676 );
    not g26906 ( n15953 , n25193 );
    nor g26907 ( n28998 , n40029 , n33808 );
    or g26908 ( n12118 , n41460 , n10491 );
    xnor g26909 ( n17652 , n836 , n19273 );
    and g26910 ( n13963 , n10461 , n23237 );
    xnor g26911 ( n11554 , n17813 , n4683 );
    not g26912 ( n17980 , n8525 );
    nor g26913 ( n31803 , n35657 , n4632 );
    and g26914 ( n17397 , n40662 , n18649 );
    or g26915 ( n18270 , n10816 , n36087 );
    and g26916 ( n8940 , n12608 , n28983 );
    or g26917 ( n22097 , n19991 , n705 );
    nor g26918 ( n36111 , n39286 , n39368 );
    not g26919 ( n11566 , n9184 );
    nor g26920 ( n18354 , n4228 , n39634 );
    and g26921 ( n25935 , n34401 , n19447 );
    or g26922 ( n15667 , n4085 , n13645 );
    or g26923 ( n16097 , n37599 , n9085 );
    not g26924 ( n2599 , n35221 );
    xnor g26925 ( n15732 , n25143 , n28900 );
    or g26926 ( n38846 , n9503 , n22766 );
    xnor g26927 ( n24002 , n27035 , n16006 );
    not g26928 ( n38119 , n22934 );
    or g26929 ( n1981 , n3630 , n42694 );
    or g26930 ( n6562 , n7701 , n27824 );
    not g26931 ( n30094 , n23715 );
    or g26932 ( n19252 , n40021 , n22728 );
    and g26933 ( n37666 , n21459 , n3602 );
    or g26934 ( n35536 , n12882 , n15293 );
    or g26935 ( n20843 , n36948 , n18019 );
    xnor g26936 ( n3348 , n105 , n22909 );
    nor g26937 ( n18065 , n25306 , n20643 );
    or g26938 ( n31521 , n31498 , n3119 );
    or g26939 ( n10050 , n41705 , n5567 );
    not g26940 ( n34090 , n42338 );
    not g26941 ( n9079 , n9512 );
    xnor g26942 ( n22771 , n39722 , n38727 );
    or g26943 ( n26574 , n28289 , n30285 );
    and g26944 ( n6436 , n24555 , n36351 );
    or g26945 ( n34737 , n2619 , n14721 );
    not g26946 ( n20245 , n28404 );
    and g26947 ( n15504 , n9056 , n5288 );
    and g26948 ( n34423 , n22738 , n7945 );
    or g26949 ( n23543 , n18261 , n26888 );
    and g26950 ( n27610 , n4848 , n40420 );
    or g26951 ( n28693 , n14287 , n18593 );
    and g26952 ( n37468 , n8471 , n31002 );
    nor g26953 ( n29340 , n34565 , n14634 );
    not g26954 ( n33721 , n23966 );
    nor g26955 ( n16020 , n17438 , n21902 );
    nor g26956 ( n30573 , n8974 , n4649 );
    nor g26957 ( n32062 , n13899 , n8040 );
    nor g26958 ( n11837 , n37815 , n53 );
    or g26959 ( n19831 , n13117 , n8662 );
    nor g26960 ( n36896 , n16598 , n28186 );
    and g26961 ( n23225 , n39281 , n13770 );
    and g26962 ( n30863 , n10922 , n42849 );
    not g26963 ( n9423 , n1991 );
    or g26964 ( n5285 , n27350 , n2466 );
    and g26965 ( n42489 , n39597 , n21640 );
    or g26966 ( n9744 , n5964 , n14643 );
    xnor g26967 ( n16647 , n35154 , n29127 );
    nor g26968 ( n1789 , n38597 , n41300 );
    or g26969 ( n13017 , n10306 , n28613 );
    or g26970 ( n19477 , n31704 , n8762 );
    not g26971 ( n2675 , n17406 );
    or g26972 ( n1737 , n22257 , n42124 );
    or g26973 ( n25563 , n38921 , n23396 );
    and g26974 ( n16186 , n4604 , n29085 );
    or g26975 ( n14109 , n12575 , n21703 );
    or g26976 ( n19008 , n37603 , n21864 );
    not g26977 ( n739 , n37515 );
    and g26978 ( n38727 , n24429 , n9186 );
    or g26979 ( n33885 , n39755 , n36193 );
    or g26980 ( n11022 , n34712 , n14569 );
    not g26981 ( n7286 , n14787 );
    and g26982 ( n36186 , n29997 , n16858 );
    and g26983 ( n26076 , n11939 , n30532 );
    or g26984 ( n25596 , n19159 , n30296 );
    and g26985 ( n620 , n37941 , n2653 );
    xnor g26986 ( n2026 , n12223 , n12903 );
    or g26987 ( n21395 , n22540 , n18735 );
    not g26988 ( n29089 , n13095 );
    or g26989 ( n29733 , n40719 , n22569 );
    or g26990 ( n34514 , n23736 , n8526 );
    xnor g26991 ( n38130 , n42203 , n5630 );
    not g26992 ( n35651 , n33418 );
    xnor g26993 ( n41042 , n19116 , n12803 );
    or g26994 ( n1862 , n24008 , n5473 );
    not g26995 ( n26633 , n7389 );
    nor g26996 ( n16029 , n32833 , n16432 );
    nor g26997 ( n20364 , n28363 , n14188 );
    or g26998 ( n7120 , n37016 , n39847 );
    or g26999 ( n5591 , n42476 , n29388 );
    or g27000 ( n23448 , n39679 , n22379 );
    or g27001 ( n2983 , n12700 , n7800 );
    xnor g27002 ( n42356 , n26279 , n25381 );
    and g27003 ( n2269 , n24028 , n42117 );
    or g27004 ( n8121 , n41081 , n11375 );
    and g27005 ( n23876 , n16261 , n7163 );
    not g27006 ( n35337 , n10697 );
    xnor g27007 ( n15509 , n11 , n17744 );
    or g27008 ( n29556 , n22804 , n38525 );
    or g27009 ( n15475 , n472 , n19969 );
    not g27010 ( n36089 , n5821 );
    or g27011 ( n21936 , n23077 , n6170 );
    or g27012 ( n41483 , n24760 , n10156 );
    nor g27013 ( n15544 , n15056 , n19527 );
    xnor g27014 ( n15450 , n21634 , n7815 );
    nor g27015 ( n35328 , n18395 , n1164 );
    nor g27016 ( n20867 , n9319 , n27503 );
    or g27017 ( n3063 , n11286 , n32037 );
    xnor g27018 ( n18013 , n29129 , n11688 );
    not g27019 ( n15524 , n21998 );
    and g27020 ( n26984 , n41378 , n9811 );
    or g27021 ( n29123 , n32068 , n32247 );
    xnor g27022 ( n9244 , n23267 , n33786 );
    and g27023 ( n13824 , n2262 , n38280 );
    and g27024 ( n34682 , n32444 , n40597 );
    or g27025 ( n17023 , n1031 , n4239 );
    or g27026 ( n36321 , n11539 , n24108 );
    nor g27027 ( n7372 , n41995 , n19960 );
    xnor g27028 ( n37758 , n2338 , n30423 );
    or g27029 ( n7819 , n4403 , n21697 );
    not g27030 ( n24610 , n33807 );
    xnor g27031 ( n42686 , n15972 , n27267 );
    or g27032 ( n24446 , n37707 , n19170 );
    or g27033 ( n41937 , n19053 , n574 );
    not g27034 ( n4257 , n23908 );
    or g27035 ( n9836 , n28451 , n37952 );
    and g27036 ( n33022 , n21786 , n28702 );
    and g27037 ( n14585 , n39943 , n18 );
    nor g27038 ( n38098 , n12960 , n6274 );
    or g27039 ( n24628 , n14164 , n2794 );
    or g27040 ( n33006 , n3800 , n31009 );
    not g27041 ( n6812 , n18480 );
    nor g27042 ( n39474 , n32539 , n24826 );
    or g27043 ( n21323 , n16431 , n38293 );
    and g27044 ( n41706 , n6396 , n19507 );
    xnor g27045 ( n6601 , n24527 , n30859 );
    or g27046 ( n25517 , n31960 , n17570 );
    nor g27047 ( n26508 , n26617 , n10447 );
    xnor g27048 ( n36356 , n15524 , n34324 );
    nor g27049 ( n25315 , n41391 , n14520 );
    not g27050 ( n3481 , n40045 );
    not g27051 ( n39226 , n5819 );
    or g27052 ( n25604 , n18812 , n38174 );
    or g27053 ( n22019 , n2937 , n40705 );
    or g27054 ( n8946 , n22348 , n28021 );
    or g27055 ( n28476 , n13041 , n27548 );
    not g27056 ( n26609 , n34173 );
    not g27057 ( n514 , n34298 );
    or g27058 ( n22273 , n12198 , n9812 );
    or g27059 ( n16172 , n2408 , n21600 );
    or g27060 ( n40119 , n25591 , n20068 );
    or g27061 ( n8856 , n37168 , n33827 );
    not g27062 ( n17404 , n29332 );
    not g27063 ( n7039 , n24762 );
    and g27064 ( n14155 , n32704 , n12013 );
    not g27065 ( n36112 , n1572 );
    and g27066 ( n33268 , n26899 , n18820 );
    or g27067 ( n12581 , n32100 , n23775 );
    and g27068 ( n22919 , n36964 , n16037 );
    xnor g27069 ( n13298 , n35259 , n6406 );
    not g27070 ( n25878 , n39987 );
    or g27071 ( n35798 , n41943 , n23422 );
    or g27072 ( n41579 , n38872 , n40854 );
    and g27073 ( n22316 , n26872 , n11341 );
    or g27074 ( n16956 , n15965 , n21788 );
    not g27075 ( n9930 , n1803 );
    and g27076 ( n14909 , n26362 , n36708 );
    nor g27077 ( n9197 , n25789 , n16234 );
    not g27078 ( n1448 , n24273 );
    or g27079 ( n35482 , n22687 , n17881 );
    not g27080 ( n12526 , n21229 );
    xnor g27081 ( n6614 , n25701 , n20729 );
    xnor g27082 ( n36970 , n18530 , n7775 );
    not g27083 ( n2034 , n29332 );
    or g27084 ( n32810 , n38844 , n36078 );
    not g27085 ( n32294 , n13996 );
    or g27086 ( n24663 , n36117 , n13504 );
    and g27087 ( n488 , n25510 , n40143 );
    not g27088 ( n9961 , n12318 );
    and g27089 ( n34288 , n1805 , n31177 );
    not g27090 ( n18798 , n30638 );
    or g27091 ( n3454 , n37131 , n11016 );
    and g27092 ( n21337 , n35645 , n24961 );
    nor g27093 ( n10608 , n28884 , n40218 );
    nor g27094 ( n35262 , n41013 , n5731 );
    or g27095 ( n17857 , n19635 , n3517 );
    or g27096 ( n29503 , n36729 , n29897 );
    xnor g27097 ( n9291 , n10123 , n19220 );
    and g27098 ( n9 , n362 , n32360 );
    and g27099 ( n34246 , n1047 , n26528 );
    nor g27100 ( n29872 , n8494 , n11071 );
    or g27101 ( n36243 , n9264 , n11660 );
    not g27102 ( n15803 , n599 );
    or g27103 ( n3833 , n7666 , n11061 );
    or g27104 ( n35327 , n37965 , n15302 );
    or g27105 ( n40346 , n26888 , n14991 );
    or g27106 ( n409 , n21174 , n36925 );
    xnor g27107 ( n32750 , n35059 , n17368 );
    and g27108 ( n31693 , n40108 , n5955 );
    or g27109 ( n4252 , n28774 , n12982 );
    xnor g27110 ( n2099 , n24892 , n32224 );
    or g27111 ( n21924 , n440 , n33567 );
    or g27112 ( n26465 , n35403 , n41207 );
    or g27113 ( n27041 , n33521 , n290 );
    and g27114 ( n10561 , n10203 , n36262 );
    or g27115 ( n38952 , n10378 , n32698 );
    or g27116 ( n18177 , n133 , n32377 );
    or g27117 ( n3797 , n42793 , n31487 );
    or g27118 ( n26550 , n39413 , n12397 );
    xnor g27119 ( n10245 , n5144 , n34204 );
    nor g27120 ( n6231 , n13269 , n21785 );
    and g27121 ( n14250 , n31723 , n13678 );
    xnor g27122 ( n11281 , n37709 , n40675 );
    not g27123 ( n3385 , n21594 );
    nor g27124 ( n26455 , n21599 , n9723 );
    and g27125 ( n41464 , n40557 , n19709 );
    or g27126 ( n26073 , n29161 , n3692 );
    not g27127 ( n32905 , n30014 );
    or g27128 ( n7010 , n23261 , n18073 );
    not g27129 ( n6024 , n26969 );
    nor g27130 ( n4190 , n41231 , n26623 );
    or g27131 ( n1689 , n26196 , n30025 );
    nor g27132 ( n3057 , n34292 , n41777 );
    xnor g27133 ( n13793 , n36998 , n4222 );
    xnor g27134 ( n8213 , n9316 , n40731 );
    xnor g27135 ( n10025 , n39104 , n11163 );
    and g27136 ( n31901 , n23382 , n18942 );
    or g27137 ( n10175 , n11898 , n31949 );
    or g27138 ( n28975 , n2608 , n41637 );
    xnor g27139 ( n7200 , n36938 , n41717 );
    not g27140 ( n31519 , n14206 );
    not g27141 ( n2338 , n8504 );
    and g27142 ( n14659 , n299 , n39886 );
    not g27143 ( n17441 , n17722 );
    nor g27144 ( n41006 , n27142 , n26808 );
    or g27145 ( n24094 , n21535 , n28500 );
    xnor g27146 ( n36882 , n15860 , n35187 );
    nor g27147 ( n2056 , n35125 , n25995 );
    xnor g27148 ( n40965 , n29450 , n1553 );
    and g27149 ( n21427 , n26692 , n42 );
    xnor g27150 ( n41991 , n35727 , n15107 );
    or g27151 ( n21651 , n20381 , n12867 );
    and g27152 ( n31217 , n27536 , n34083 );
    nor g27153 ( n9579 , n30505 , n28284 );
    nor g27154 ( n2384 , n5869 , n32838 );
    or g27155 ( n4053 , n33902 , n17084 );
    nor g27156 ( n3816 , n38782 , n18744 );
    and g27157 ( n42899 , n15736 , n29132 );
    or g27158 ( n17799 , n41521 , n27136 );
    or g27159 ( n12164 , n7839 , n15084 );
    or g27160 ( n37846 , n18660 , n11432 );
    or g27161 ( n27005 , n14844 , n31321 );
    or g27162 ( n12368 , n34169 , n14053 );
    and g27163 ( n38955 , n21593 , n9111 );
    or g27164 ( n20806 , n23277 , n22551 );
    and g27165 ( n27673 , n16570 , n38187 );
    not g27166 ( n9754 , n5582 );
    and g27167 ( n705 , n28688 , n11950 );
    or g27168 ( n15521 , n500 , n2470 );
    nor g27169 ( n4221 , n41040 , n40668 );
    xnor g27170 ( n737 , n7943 , n10751 );
    or g27171 ( n20423 , n31375 , n18772 );
    or g27172 ( n37753 , n40576 , n245 );
    not g27173 ( n29261 , n7380 );
    and g27174 ( n38623 , n31040 , n21110 );
    nor g27175 ( n10852 , n34651 , n19036 );
    and g27176 ( n34169 , n29238 , n12454 );
    xnor g27177 ( n11003 , n3683 , n6417 );
    and g27178 ( n18750 , n11951 , n20267 );
    and g27179 ( n629 , n39718 , n19094 );
    and g27180 ( n37559 , n31058 , n7586 );
    not g27181 ( n22263 , n17193 );
    or g27182 ( n23299 , n4775 , n5692 );
    or g27183 ( n30121 , n42321 , n35866 );
    or g27184 ( n37627 , n42032 , n12754 );
    and g27185 ( n27863 , n40962 , n35128 );
    or g27186 ( n4419 , n7549 , n18342 );
    nor g27187 ( n40538 , n11938 , n17288 );
    or g27188 ( n31003 , n27241 , n32594 );
    or g27189 ( n34914 , n38426 , n22554 );
    nor g27190 ( n28390 , n20727 , n2804 );
    or g27191 ( n17839 , n21000 , n30652 );
    not g27192 ( n13714 , n13138 );
    or g27193 ( n32075 , n22862 , n32646 );
    or g27194 ( n18560 , n10521 , n33926 );
    xnor g27195 ( n38824 , n42209 , n26856 );
    and g27196 ( n2434 , n9246 , n5209 );
    xnor g27197 ( n20526 , n25676 , n36963 );
    nor g27198 ( n16825 , n17744 , n3563 );
    not g27199 ( n10953 , n3361 );
    nor g27200 ( n17311 , n7158 , n19108 );
    nor g27201 ( n22925 , n26534 , n4198 );
    or g27202 ( n40802 , n20446 , n10272 );
    and g27203 ( n28689 , n37702 , n5070 );
    or g27204 ( n1076 , n42649 , n17758 );
    and g27205 ( n22178 , n23193 , n40493 );
    not g27206 ( n18696 , n6984 );
    and g27207 ( n24885 , n42527 , n17600 );
    or g27208 ( n39996 , n734 , n6886 );
    nor g27209 ( n35751 , n29019 , n31213 );
    or g27210 ( n23768 , n4414 , n3190 );
    or g27211 ( n36888 , n37883 , n5178 );
    not g27212 ( n16952 , n13753 );
    not g27213 ( n31681 , n27759 );
    and g27214 ( n34164 , n19671 , n31915 );
    or g27215 ( n33215 , n5558 , n36936 );
    or g27216 ( n16084 , n37980 , n10736 );
    nor g27217 ( n33034 , n12222 , n22628 );
    nor g27218 ( n26359 , n34292 , n36716 );
    or g27219 ( n19161 , n18645 , n12022 );
    or g27220 ( n7179 , n28643 , n39575 );
    not g27221 ( n28544 , n3468 );
    and g27222 ( n29788 , n13876 , n31381 );
    nor g27223 ( n19690 , n27398 , n5423 );
    or g27224 ( n28450 , n2512 , n28136 );
    not g27225 ( n566 , n35394 );
    and g27226 ( n24841 , n25502 , n19588 );
    and g27227 ( n23561 , n25979 , n10750 );
    not g27228 ( n26911 , n32817 );
    or g27229 ( n39623 , n19980 , n4107 );
    nor g27230 ( n5330 , n5768 , n8078 );
    and g27231 ( n28953 , n19088 , n41273 );
    or g27232 ( n29045 , n22950 , n38438 );
    not g27233 ( n38749 , n41623 );
    or g27234 ( n33984 , n24146 , n39991 );
    nor g27235 ( n12119 , n13899 , n38647 );
    and g27236 ( n34359 , n27055 , n30723 );
    and g27237 ( n19421 , n1137 , n42716 );
    and g27238 ( n22061 , n21633 , n25311 );
    or g27239 ( n17820 , n3051 , n32875 );
    or g27240 ( n7944 , n28883 , n2882 );
    not g27241 ( n41992 , n40372 );
    nor g27242 ( n36242 , n20345 , n29069 );
    nor g27243 ( n12727 , n5808 , n24704 );
    and g27244 ( n10781 , n3087 , n12572 );
    nor g27245 ( n2922 , n19855 , n30995 );
    or g27246 ( n39339 , n30502 , n25104 );
    or g27247 ( n20214 , n35770 , n23548 );
    not g27248 ( n23926 , n31294 );
    and g27249 ( n14967 , n2751 , n13975 );
    not g27250 ( n14489 , n9290 );
    nor g27251 ( n6292 , n34975 , n25625 );
    or g27252 ( n4407 , n25781 , n23589 );
    or g27253 ( n1306 , n9245 , n5150 );
    nor g27254 ( n35091 , n41309 , n10725 );
    and g27255 ( n3537 , n22248 , n30335 );
    or g27256 ( n5820 , n15070 , n36524 );
    or g27257 ( n17927 , n19748 , n27280 );
    and g27258 ( n35882 , n1477 , n42078 );
    or g27259 ( n9346 , n6098 , n26384 );
    nor g27260 ( n39674 , n25173 , n8254 );
    xnor g27261 ( n34049 , n29800 , n15953 );
    and g27262 ( n8338 , n32665 , n10774 );
    nor g27263 ( n2309 , n16780 , n25446 );
    or g27264 ( n85 , n4394 , n4637 );
    or g27265 ( n11261 , n19803 , n3263 );
    and g27266 ( n30720 , n35059 , n17368 );
    not g27267 ( n5227 , n12247 );
    and g27268 ( n16599 , n2681 , n29405 );
    or g27269 ( n24351 , n1960 , n19847 );
    and g27270 ( n7692 , n23715 , n28326 );
    not g27271 ( n30538 , n36674 );
    xnor g27272 ( n20803 , n27734 , n35859 );
    or g27273 ( n13572 , n31703 , n7242 );
    or g27274 ( n3821 , n41530 , n27127 );
    and g27275 ( n5033 , n7352 , n4019 );
    and g27276 ( n38110 , n24411 , n36006 );
    and g27277 ( n13507 , n36055 , n23923 );
    and g27278 ( n27730 , n41529 , n36655 );
    and g27279 ( n36536 , n16933 , n11973 );
    and g27280 ( n13747 , n2955 , n40939 );
    not g27281 ( n9370 , n21306 );
    or g27282 ( n26282 , n37959 , n16046 );
    nor g27283 ( n39583 , n25917 , n22250 );
    not g27284 ( n32967 , n16857 );
    nor g27285 ( n21660 , n26503 , n9440 );
    nor g27286 ( n32011 , n3524 , n42742 );
    not g27287 ( n33837 , n28224 );
    or g27288 ( n19657 , n3077 , n18185 );
    nor g27289 ( n12692 , n13151 , n29197 );
    or g27290 ( n35363 , n33522 , n13566 );
    or g27291 ( n30245 , n8087 , n4551 );
    or g27292 ( n37570 , n7127 , n12926 );
    xnor g27293 ( n6908 , n34731 , n8468 );
    not g27294 ( n10160 , n8834 );
    and g27295 ( n1783 , n16953 , n4986 );
    not g27296 ( n1658 , n17156 );
    or g27297 ( n8205 , n991 , n40862 );
    nor g27298 ( n35359 , n38836 , n27624 );
    xnor g27299 ( n4034 , n9550 , n39266 );
    xnor g27300 ( n29359 , n30830 , n34842 );
    or g27301 ( n8394 , n16848 , n25129 );
    and g27302 ( n33431 , n7135 , n25363 );
    not g27303 ( n26274 , n4276 );
    and g27304 ( n42654 , n7064 , n26738 );
    or g27305 ( n36354 , n29058 , n36073 );
    and g27306 ( n36793 , n24397 , n9575 );
    or g27307 ( n36231 , n17002 , n11178 );
    or g27308 ( n40953 , n3706 , n2429 );
    not g27309 ( n3949 , n38571 );
    xnor g27310 ( n21851 , n40638 , n42855 );
    or g27311 ( n37375 , n8156 , n17633 );
    not g27312 ( n21998 , n38992 );
    and g27313 ( n33468 , n4615 , n15839 );
    or g27314 ( n29502 , n28685 , n41424 );
    and g27315 ( n34544 , n36051 , n31819 );
    xnor g27316 ( n32843 , n6767 , n39055 );
    or g27317 ( n30292 , n42732 , n31503 );
    and g27318 ( n28847 , n29055 , n16283 );
    or g27319 ( n23058 , n712 , n40319 );
    xnor g27320 ( n28981 , n42064 , n24012 );
    nor g27321 ( n14591 , n2199 , n18978 );
    and g27322 ( n4768 , n22030 , n21302 );
    or g27323 ( n15225 , n5795 , n12829 );
    xnor g27324 ( n27517 , n6067 , n36102 );
    not g27325 ( n39861 , n11881 );
    not g27326 ( n37237 , n32657 );
    or g27327 ( n21261 , n38584 , n12199 );
    nor g27328 ( n39881 , n28694 , n36058 );
    or g27329 ( n20655 , n14048 , n17433 );
    or g27330 ( n19739 , n4241 , n1735 );
    nor g27331 ( n32390 , n3299 , n16946 );
    and g27332 ( n24103 , n24914 , n3387 );
    and g27333 ( n20227 , n4393 , n34339 );
    or g27334 ( n12708 , n1518 , n26789 );
    not g27335 ( n34594 , n3178 );
    or g27336 ( n32381 , n3580 , n37816 );
    not g27337 ( n7001 , n38080 );
    or g27338 ( n3872 , n17903 , n32167 );
    or g27339 ( n39020 , n33474 , n20856 );
    and g27340 ( n3901 , n1473 , n31423 );
    not g27341 ( n41239 , n40721 );
    or g27342 ( n23033 , n25507 , n34535 );
    and g27343 ( n15299 , n1081 , n214 );
    or g27344 ( n30291 , n36036 , n41543 );
    not g27345 ( n1 , n2358 );
    and g27346 ( n24805 , n26318 , n31362 );
    not g27347 ( n18736 , n8747 );
    nor g27348 ( n34166 , n13845 , n6298 );
    or g27349 ( n25916 , n30844 , n1884 );
    or g27350 ( n24059 , n20549 , n35155 );
    or g27351 ( n2553 , n34184 , n14983 );
    not g27352 ( n31777 , n17346 );
    or g27353 ( n42235 , n26120 , n9418 );
    or g27354 ( n384 , n36051 , n31819 );
    or g27355 ( n17294 , n11431 , n24440 );
    or g27356 ( n31338 , n33289 , n31101 );
    not g27357 ( n861 , n34277 );
    not g27358 ( n36993 , n35238 );
    or g27359 ( n32713 , n22864 , n22476 );
    or g27360 ( n27216 , n23906 , n30367 );
    not g27361 ( n11724 , n14478 );
    and g27362 ( n18662 , n20966 , n41190 );
    nor g27363 ( n37906 , n10011 , n7144 );
    nor g27364 ( n32797 , n33433 , n30118 );
    and g27365 ( n11257 , n21383 , n12548 );
    or g27366 ( n39268 , n22349 , n37647 );
    and g27367 ( n42084 , n7419 , n7052 );
    or g27368 ( n17269 , n38576 , n34785 );
    or g27369 ( n41033 , n31216 , n9417 );
    or g27370 ( n42075 , n24212 , n12958 );
    and g27371 ( n2713 , n42276 , n1543 );
    nor g27372 ( n6665 , n16403 , n24317 );
    or g27373 ( n38252 , n18827 , n28028 );
    or g27374 ( n25103 , n81 , n14044 );
    or g27375 ( n4596 , n24754 , n32973 );
    or g27376 ( n27481 , n36143 , n40795 );
    and g27377 ( n30212 , n32058 , n27185 );
    or g27378 ( n39224 , n35866 , n2991 );
    or g27379 ( n28260 , n17585 , n41540 );
    not g27380 ( n31665 , n3898 );
    nor g27381 ( n4258 , n9557 , n31640 );
    or g27382 ( n18799 , n9647 , n28985 );
    and g27383 ( n38412 , n36510 , n14477 );
    or g27384 ( n12977 , n18817 , n40235 );
    xnor g27385 ( n22407 , n898 , n11510 );
    not g27386 ( n41616 , n7820 );
    xnor g27387 ( n28605 , n12982 , n4140 );
    or g27388 ( n42296 , n543 , n12198 );
    or g27389 ( n42239 , n35197 , n2179 );
    or g27390 ( n1438 , n34184 , n9801 );
    or g27391 ( n31624 , n42826 , n28021 );
    or g27392 ( n19410 , n34539 , n14944 );
    not g27393 ( n13195 , n6365 );
    and g27394 ( n22253 , n36011 , n32841 );
    nor g27395 ( n1175 , n14382 , n39091 );
    nor g27396 ( n8262 , n2849 , n32110 );
    not g27397 ( n12745 , n13009 );
    or g27398 ( n38654 , n13435 , n25862 );
    xnor g27399 ( n4425 , n6885 , n33680 );
    or g27400 ( n13259 , n5964 , n16197 );
    nor g27401 ( n22971 , n38879 , n38510 );
    or g27402 ( n19420 , n9873 , n11178 );
    not g27403 ( n28314 , n14924 );
    nor g27404 ( n23855 , n10510 , n35106 );
    and g27405 ( n28508 , n25724 , n42470 );
    nor g27406 ( n39948 , n12054 , n27945 );
    not g27407 ( n34728 , n30929 );
    xnor g27408 ( n7178 , n24306 , n23628 );
    or g27409 ( n6474 , n27335 , n34634 );
    or g27410 ( n2001 , n22043 , n32623 );
    nor g27411 ( n24402 , n34565 , n26244 );
    and g27412 ( n11318 , n26699 , n32357 );
    or g27413 ( n18478 , n14471 , n6371 );
    not g27414 ( n18495 , n39543 );
    not g27415 ( n12098 , n42707 );
    and g27416 ( n22156 , n27509 , n23269 );
    not g27417 ( n38563 , n366 );
    or g27418 ( n113 , n32985 , n16285 );
    or g27419 ( n45 , n40212 , n7593 );
    or g27420 ( n13404 , n41684 , n21132 );
    not g27421 ( n7378 , n26515 );
    or g27422 ( n18991 , n10435 , n23017 );
    or g27423 ( n40700 , n39493 , n7815 );
    nor g27424 ( n23427 , n39174 , n14345 );
    nor g27425 ( n7794 , n19260 , n10804 );
    or g27426 ( n18351 , n34651 , n31902 );
    and g27427 ( n9935 , n10652 , n8153 );
    or g27428 ( n31840 , n35548 , n30340 );
    or g27429 ( n36357 , n26500 , n26006 );
    not g27430 ( n14667 , n30728 );
    nor g27431 ( n8594 , n16039 , n7275 );
    not g27432 ( n40237 , n28518 );
    and g27433 ( n12298 , n27847 , n14795 );
    and g27434 ( n17849 , n21616 , n32737 );
    or g27435 ( n30817 , n1788 , n41639 );
    or g27436 ( n37287 , n23637 , n15256 );
    or g27437 ( n42545 , n2272 , n33321 );
    or g27438 ( n39325 , n32405 , n21516 );
    or g27439 ( n23660 , n15492 , n12904 );
    or g27440 ( n37097 , n26652 , n3135 );
    or g27441 ( n39751 , n11068 , n1970 );
    or g27442 ( n30806 , n29322 , n42088 );
    and g27443 ( n15540 , n20619 , n9842 );
    or g27444 ( n13907 , n440 , n3149 );
    xnor g27445 ( n32004 , n23686 , n27186 );
    and g27446 ( n15487 , n17879 , n39469 );
    not g27447 ( n22604 , n26358 );
    or g27448 ( n9593 , n12315 , n20921 );
    xnor g27449 ( n13781 , n4481 , n9320 );
    and g27450 ( n18984 , n32073 , n6986 );
    or g27451 ( n18128 , n10926 , n3994 );
    xnor g27452 ( n16298 , n37896 , n15893 );
    nor g27453 ( n40262 , n38640 , n34188 );
    and g27454 ( n10733 , n33229 , n10006 );
    or g27455 ( n14421 , n668 , n12382 );
    or g27456 ( n32365 , n42421 , n13099 );
    xnor g27457 ( n42373 , n8502 , n39506 );
    and g27458 ( n3100 , n6364 , n16162 );
    not g27459 ( n13529 , n38262 );
    xnor g27460 ( n7639 , n26542 , n25202 );
    and g27461 ( n14450 , n8435 , n33309 );
    or g27462 ( n9188 , n18026 , n2983 );
    nor g27463 ( n22748 , n15070 , n17545 );
    or g27464 ( n25013 , n29658 , n13165 );
    xnor g27465 ( n13449 , n10303 , n31868 );
    and g27466 ( n17107 , n26303 , n21989 );
    or g27467 ( n10209 , n35706 , n6445 );
    or g27468 ( n32251 , n20978 , n38409 );
    not g27469 ( n28010 , n30210 );
    and g27470 ( n29118 , n8962 , n31296 );
    or g27471 ( n8271 , n16648 , n27079 );
    or g27472 ( n12771 , n24972 , n30590 );
    and g27473 ( n27562 , n42239 , n34683 );
    and g27474 ( n3213 , n10271 , n38660 );
    not g27475 ( n12851 , n29575 );
    not g27476 ( n39539 , n36151 );
    and g27477 ( n29979 , n27795 , n41843 );
    or g27478 ( n13062 , n30046 , n39345 );
    or g27479 ( n34243 , n7849 , n25233 );
    not g27480 ( n30979 , n348 );
    and g27481 ( n27033 , n42051 , n24663 );
    and g27482 ( n1774 , n39453 , n26249 );
    or g27483 ( n7843 , n4501 , n38058 );
    or g27484 ( n2613 , n3415 , n26545 );
    nor g27485 ( n2267 , n34761 , n22164 );
    or g27486 ( n38182 , n28596 , n14585 );
    nor g27487 ( n14750 , n1971 , n24238 );
    and g27488 ( n3521 , n10887 , n30468 );
    or g27489 ( n8286 , n15070 , n33878 );
    nor g27490 ( n3786 , n1301 , n23607 );
    nor g27491 ( n13702 , n23485 , n8884 );
    xnor g27492 ( n27343 , n11133 , n5812 );
    xnor g27493 ( n22213 , n14419 , n4001 );
    nor g27494 ( n38872 , n35289 , n33036 );
    or g27495 ( n10403 , n34114 , n40277 );
    or g27496 ( n11382 , n27081 , n14216 );
    or g27497 ( n30248 , n20069 , n35879 );
    not g27498 ( n21199 , n14394 );
    not g27499 ( n14070 , n40297 );
    or g27500 ( n23631 , n42650 , n31569 );
    xnor g27501 ( n26537 , n17264 , n41710 );
    nor g27502 ( n24542 , n17476 , n9659 );
    nor g27503 ( n4724 , n28407 , n23254 );
    nor g27504 ( n40568 , n16977 , n29721 );
    nor g27505 ( n30810 , n9272 , n6515 );
    or g27506 ( n27361 , n29054 , n17102 );
    xnor g27507 ( n5857 , n18530 , n9709 );
    and g27508 ( n16601 , n41125 , n36686 );
    not g27509 ( n17567 , n11830 );
    or g27510 ( n42353 , n36724 , n24088 );
    nor g27511 ( n26461 , n16489 , n34225 );
    not g27512 ( n18873 , n26724 );
    xnor g27513 ( n37245 , n20015 , n9873 );
    or g27514 ( n31855 , n27380 , n38459 );
    and g27515 ( n18121 , n40780 , n23687 );
    not g27516 ( n6728 , n41256 );
    or g27517 ( n17248 , n2160 , n22325 );
    xnor g27518 ( n5655 , n20487 , n38354 );
    and g27519 ( n9563 , n24176 , n41804 );
    or g27520 ( n12834 , n42376 , n1120 );
    or g27521 ( n25489 , n37565 , n23130 );
    xnor g27522 ( n4200 , n36562 , n26049 );
    or g27523 ( n27696 , n30358 , n35260 );
    nor g27524 ( n39823 , n17909 , n13549 );
    nor g27525 ( n31520 , n16244 , n4653 );
    and g27526 ( n13815 , n42224 , n27652 );
    xnor g27527 ( n26535 , n13444 , n12515 );
    or g27528 ( n38599 , n29913 , n40381 );
    not g27529 ( n5311 , n11437 );
    or g27530 ( n2975 , n25322 , n10111 );
    nor g27531 ( n16383 , n25155 , n35956 );
    or g27532 ( n16963 , n22641 , n42479 );
    nor g27533 ( n1597 , n38256 , n13664 );
    not g27534 ( n34651 , n478 );
    or g27535 ( n27304 , n25587 , n8988 );
    or g27536 ( n36015 , n8731 , n31656 );
    or g27537 ( n28170 , n39275 , n34608 );
    xnor g27538 ( n14946 , n7922 , n12807 );
    nor g27539 ( n5264 , n34565 , n17657 );
    xnor g27540 ( n34102 , n19519 , n39844 );
    xnor g27541 ( n22259 , n41695 , n15671 );
    or g27542 ( n20284 , n5308 , n24535 );
    xnor g27543 ( n37049 , n38749 , n10685 );
    or g27544 ( n20805 , n5166 , n26295 );
    and g27545 ( n41354 , n21726 , n21271 );
    or g27546 ( n4237 , n22622 , n21807 );
    or g27547 ( n5548 , n10208 , n10308 );
    or g27548 ( n10787 , n20191 , n28461 );
    and g27549 ( n37549 , n22038 , n14204 );
    and g27550 ( n37591 , n20527 , n26146 );
    or g27551 ( n21135 , n25279 , n17629 );
    not g27552 ( n24105 , n16350 );
    nor g27553 ( n14666 , n27960 , n21747 );
    or g27554 ( n10401 , n6574 , n33691 );
    xnor g27555 ( n40498 , n14034 , n16632 );
    or g27556 ( n31085 , n6358 , n10241 );
    xnor g27557 ( n6519 , n40 , n27580 );
    nor g27558 ( n32290 , n11784 , n20359 );
    or g27559 ( n27607 , n21212 , n32194 );
    and g27560 ( n7466 , n16740 , n9004 );
    nor g27561 ( n30167 , n27324 , n26826 );
    nor g27562 ( n25581 , n34565 , n17291 );
    or g27563 ( n15864 , n22159 , n22987 );
    not g27564 ( n3490 , n20416 );
    nor g27565 ( n7331 , n17744 , n34549 );
    xnor g27566 ( n11542 , n31989 , n16911 );
    xnor g27567 ( n18912 , n29786 , n18030 );
    nor g27568 ( n40877 , n39604 , n39211 );
    or g27569 ( n36287 , n36831 , n16485 );
    nor g27570 ( n28129 , n20115 , n20399 );
    or g27571 ( n22083 , n11798 , n6571 );
    nor g27572 ( n5012 , n5896 , n23 );
    or g27573 ( n16898 , n6201 , n22733 );
    not g27574 ( n33750 , n26467 );
    or g27575 ( n28717 , n15384 , n24765 );
    and g27576 ( n17919 , n25834 , n17487 );
    nor g27577 ( n16338 , n6303 , n11443 );
    or g27578 ( n29152 , n14308 , n35401 );
    not g27579 ( n16532 , n9051 );
    or g27580 ( n20679 , n22561 , n3077 );
    and g27581 ( n2600 , n11635 , n582 );
    nor g27582 ( n37402 , n23407 , n41149 );
    and g27583 ( n12907 , n35038 , n40385 );
    or g27584 ( n20326 , n40944 , n37263 );
    or g27585 ( n14518 , n39560 , n8092 );
    and g27586 ( n37968 , n16120 , n40125 );
    xnor g27587 ( n42047 , n34731 , n5278 );
    or g27588 ( n41742 , n35423 , n22942 );
    not g27589 ( n19796 , n5213 );
    not g27590 ( n3080 , n17234 );
    xnor g27591 ( n34156 , n35727 , n20341 );
    or g27592 ( n15977 , n22372 , n16957 );
    not g27593 ( n20370 , n22424 );
    or g27594 ( n12006 , n27450 , n30383 );
    not g27595 ( n10929 , n6260 );
    nor g27596 ( n28451 , n35588 , n28654 );
    nor g27597 ( n7021 , n31771 , n7251 );
    or g27598 ( n20182 , n26476 , n31910 );
    and g27599 ( n36915 , n35836 , n30934 );
    or g27600 ( n25411 , n937 , n2089 );
    xnor g27601 ( n17349 , n32731 , n37728 );
    or g27602 ( n6095 , n16784 , n33755 );
    or g27603 ( n100 , n40109 , n6837 );
    and g27604 ( n6418 , n37400 , n35816 );
    not g27605 ( n11799 , n15356 );
    and g27606 ( n23513 , n34193 , n27889 );
    or g27607 ( n30459 , n40456 , n9708 );
    or g27608 ( n5590 , n7962 , n15095 );
    or g27609 ( n17701 , n5745 , n1256 );
    or g27610 ( n5104 , n28554 , n40547 );
    or g27611 ( n17409 , n36585 , n24322 );
    or g27612 ( n38468 , n28407 , n18315 );
    and g27613 ( n33869 , n42526 , n14858 );
    or g27614 ( n33083 , n241 , n6374 );
    not g27615 ( n9377 , n23347 );
    xnor g27616 ( n27784 , n3885 , n39266 );
    nor g27617 ( n18115 , n39927 , n33985 );
    and g27618 ( n1584 , n21146 , n10264 );
    not g27619 ( n30005 , n13335 );
    xnor g27620 ( n28974 , n21973 , n5039 );
    and g27621 ( n11324 , n5067 , n23713 );
    or g27622 ( n20308 , n25573 , n25239 );
    or g27623 ( n41507 , n6480 , n16460 );
    nor g27624 ( n37103 , n17744 , n15550 );
    or g27625 ( n30526 , n5498 , n22791 );
    and g27626 ( n38374 , n38476 , n21936 );
    or g27627 ( n9380 , n26155 , n40194 );
    or g27628 ( n26206 , n39583 , n25036 );
    nor g27629 ( n23762 , n35743 , n6985 );
    not g27630 ( n1761 , n7693 );
    nor g27631 ( n27001 , n35310 , n16563 );
    or g27632 ( n22880 , n35140 , n39536 );
    and g27633 ( n13504 , n18752 , n39691 );
    or g27634 ( n22869 , n31600 , n24254 );
    xnor g27635 ( n25788 , n6650 , n33857 );
    or g27636 ( n9086 , n42006 , n4842 );
    or g27637 ( n1310 , n10598 , n2227 );
    or g27638 ( n10550 , n8847 , n25614 );
    and g27639 ( n3925 , n41805 , n22493 );
    xnor g27640 ( n33466 , n16866 , n11774 );
    and g27641 ( n36492 , n31788 , n6225 );
    not g27642 ( n28490 , n33397 );
    nor g27643 ( n29149 , n25172 , n41425 );
    xnor g27644 ( n16171 , n1768 , n23313 );
    xnor g27645 ( n18751 , n38777 , n4360 );
    xnor g27646 ( n27138 , n15972 , n10447 );
    or g27647 ( n21990 , n18257 , n21327 );
    or g27648 ( n24384 , n42901 , n6478 );
    and g27649 ( n27091 , n4572 , n33975 );
    or g27650 ( n25336 , n36235 , n20352 );
    or g27651 ( n14086 , n25600 , n20440 );
    and g27652 ( n33128 , n13844 , n40706 );
    and g27653 ( n15531 , n32953 , n8629 );
    and g27654 ( n2735 , n26724 , n5817 );
    not g27655 ( n33053 , n39139 );
    not g27656 ( n11269 , n39378 );
    and g27657 ( n24784 , n26105 , n37358 );
    not g27658 ( n40390 , n8642 );
    and g27659 ( n16401 , n37727 , n26608 );
    xnor g27660 ( n16622 , n14978 , n11684 );
    or g27661 ( n2097 , n18242 , n27378 );
    or g27662 ( n29509 , n1185 , n6273 );
    nor g27663 ( n9885 , n27762 , n583 );
    and g27664 ( n33637 , n24911 , n4960 );
    or g27665 ( n38925 , n37776 , n34167 );
    nor g27666 ( n18806 , n13811 , n686 );
    or g27667 ( n41279 , n4405 , n38142 );
    and g27668 ( n33658 , n9561 , n16377 );
    not g27669 ( n4008 , n34911 );
    or g27670 ( n31655 , n15526 , n3701 );
    or g27671 ( n29145 , n40109 , n39455 );
    or g27672 ( n34369 , n29932 , n39146 );
    nor g27673 ( n20249 , n8194 , n37867 );
    nor g27674 ( n41340 , n39700 , n24653 );
    and g27675 ( n35606 , n31553 , n6850 );
    or g27676 ( n15878 , n24627 , n17321 );
    or g27677 ( n15041 , n31579 , n9040 );
    or g27678 ( n39890 , n20215 , n1326 );
    nor g27679 ( n11066 , n5236 , n41177 );
    not g27680 ( n31009 , n384 );
    and g27681 ( n23035 , n16672 , n36 );
    xnor g27682 ( n23145 , n24750 , n37468 );
    nor g27683 ( n29074 , n20158 , n42032 );
    or g27684 ( n9073 , n38837 , n26684 );
    or g27685 ( n25712 , n34093 , n16986 );
    and g27686 ( n20409 , n32164 , n1813 );
    or g27687 ( n18813 , n40970 , n34029 );
    nor g27688 ( n22866 , n33730 , n19936 );
    and g27689 ( n24782 , n17018 , n27437 );
    or g27690 ( n1745 , n4854 , n17926 );
    or g27691 ( n32915 , n28247 , n11731 );
    nor g27692 ( n26357 , n17100 , n4119 );
    and g27693 ( n42758 , n42564 , n30548 );
    or g27694 ( n22390 , n20116 , n34533 );
    or g27695 ( n19430 , n6651 , n30184 );
    or g27696 ( n25086 , n28286 , n38325 );
    or g27697 ( n15497 , n2277 , n23895 );
    and g27698 ( n35511 , n33651 , n6804 );
    not g27699 ( n32751 , n15401 );
    and g27700 ( n38379 , n4174 , n18253 );
    or g27701 ( n32304 , n7609 , n8752 );
    or g27702 ( n38502 , n5847 , n41819 );
    or g27703 ( n28957 , n623 , n10302 );
    or g27704 ( n26311 , n23244 , n17914 );
    and g27705 ( n36401 , n31476 , n18001 );
    or g27706 ( n6204 , n803 , n6537 );
    and g27707 ( n32398 , n32870 , n6491 );
    and g27708 ( n12811 , n24293 , n18824 );
    and g27709 ( n14985 , n18994 , n29618 );
    xnor g27710 ( n40911 , n35897 , n33622 );
    or g27711 ( n22049 , n11693 , n25221 );
    or g27712 ( n36390 , n17644 , n1908 );
    or g27713 ( n38521 , n8952 , n18805 );
    not g27714 ( n37577 , n392 );
    or g27715 ( n10982 , n30423 , n29857 );
    not g27716 ( n25964 , n37694 );
    or g27717 ( n6664 , n122 , n31678 );
    or g27718 ( n12529 , n38443 , n12153 );
    nor g27719 ( n18373 , n16018 , n31877 );
    xnor g27720 ( n2483 , n15796 , n20406 );
    xnor g27721 ( n15480 , n17476 , n42874 );
    nor g27722 ( n19370 , n34813 , n39314 );
    xnor g27723 ( n38580 , n784 , n816 );
    not g27724 ( n19396 , n17893 );
    nor g27725 ( n34353 , n39036 , n21263 );
    xnor g27726 ( n19591 , n35727 , n813 );
    not g27727 ( n41471 , n21933 );
    or g27728 ( n36121 , n34743 , n9145 );
    nor g27729 ( n10569 , n25817 , n34984 );
    or g27730 ( n23578 , n39182 , n42894 );
    nor g27731 ( n6566 , n7443 , n21341 );
    or g27732 ( n916 , n42895 , n32267 );
    or g27733 ( n23255 , n18401 , n27621 );
    and g27734 ( n16357 , n19040 , n38298 );
    not g27735 ( n9819 , n4058 );
    or g27736 ( n32907 , n20488 , n14099 );
    or g27737 ( n24529 , n9703 , n7737 );
    and g27738 ( n24026 , n17588 , n15539 );
    xnor g27739 ( n40008 , n32506 , n24755 );
    or g27740 ( n4826 , n15806 , n38632 );
    and g27741 ( n143 , n12282 , n14651 );
    not g27742 ( n23173 , n25031 );
    or g27743 ( n2779 , n14704 , n31995 );
    xnor g27744 ( n34978 , n9669 , n12917 );
    or g27745 ( n7618 , n22146 , n26409 );
    and g27746 ( n12610 , n15993 , n6882 );
    or g27747 ( n14293 , n4084 , n8088 );
    nor g27748 ( n33256 , n3098 , n23263 );
    and g27749 ( n17844 , n9170 , n40408 );
    or g27750 ( n22893 , n5426 , n36687 );
    nor g27751 ( n42519 , n25703 , n21952 );
    or g27752 ( n23570 , n41601 , n18931 );
    nor g27753 ( n3185 , n10152 , n4787 );
    or g27754 ( n26155 , n356 , n31950 );
    or g27755 ( n29825 , n15315 , n16410 );
    not g27756 ( n41670 , n16536 );
    not g27757 ( n7673 , n35391 );
    not g27758 ( n6430 , n14186 );
    nor g27759 ( n39563 , n36749 , n6922 );
    not g27760 ( n15391 , n41063 );
    or g27761 ( n14030 , n32410 , n42365 );
    or g27762 ( n22308 , n34281 , n8946 );
    nor g27763 ( n41987 , n5099 , n35280 );
    not g27764 ( n6152 , n8084 );
    xnor g27765 ( n8631 , n13353 , n22908 );
    not g27766 ( n28947 , n33951 );
    xnor g27767 ( n15195 , n18696 , n8322 );
    xnor g27768 ( n19926 , n34731 , n15958 );
    or g27769 ( n41421 , n10090 , n21867 );
    not g27770 ( n22863 , n3198 );
    xnor g27771 ( n5043 , n10906 , n16160 );
    not g27772 ( n37707 , n25592 );
    not g27773 ( n38262 , n33843 );
    and g27774 ( n32730 , n36138 , n3456 );
    nor g27775 ( n39626 , n15281 , n16060 );
    xnor g27776 ( n10316 , n6625 , n12931 );
    not g27777 ( n25247 , n39861 );
    nor g27778 ( n19731 , n3795 , n38461 );
    not g27779 ( n36619 , n4280 );
    not g27780 ( n2943 , n411 );
    not g27781 ( n37722 , n434 );
    or g27782 ( n25096 , n35386 , n22703 );
    xnor g27783 ( n7888 , n711 , n38879 );
    or g27784 ( n25606 , n13132 , n37578 );
    nor g27785 ( n12554 , n33312 , n9120 );
    or g27786 ( n3266 , n1669 , n12177 );
    or g27787 ( n26326 , n19009 , n22932 );
    or g27788 ( n19060 , n11069 , n29194 );
    and g27789 ( n975 , n11240 , n31668 );
    or g27790 ( n40573 , n27431 , n34972 );
    not g27791 ( n24183 , n17598 );
    xnor g27792 ( n25357 , n784 , n15278 );
    not g27793 ( n31415 , n5811 );
    or g27794 ( n14893 , n36604 , n29974 );
    or g27795 ( n17622 , n1581 , n41298 );
    or g27796 ( n22486 , n638 , n3031 );
    and g27797 ( n5906 , n24573 , n22111 );
    and g27798 ( n35227 , n39028 , n18626 );
    not g27799 ( n12804 , n35112 );
    xnor g27800 ( n39305 , n17264 , n19379 );
    and g27801 ( n1199 , n7990 , n24462 );
    and g27802 ( n32549 , n30385 , n2879 );
    not g27803 ( n21826 , n5842 );
    nor g27804 ( n1577 , n28593 , n1251 );
    or g27805 ( n26948 , n5380 , n27127 );
    or g27806 ( n35913 , n560 , n30329 );
    not g27807 ( n24115 , n33632 );
    or g27808 ( n25463 , n39501 , n29918 );
    and g27809 ( n23675 , n1421 , n12929 );
    and g27810 ( n14431 , n28092 , n27247 );
    and g27811 ( n36842 , n7091 , n706 );
    or g27812 ( n12496 , n29214 , n17901 );
    or g27813 ( n16122 , n22078 , n5100 );
    and g27814 ( n32153 , n6625 , n20105 );
    or g27815 ( n13695 , n40710 , n30004 );
    xnor g27816 ( n41291 , n34731 , n15690 );
    and g27817 ( n22784 , n8266 , n32421 );
    and g27818 ( n25481 , n954 , n33947 );
    nor g27819 ( n18025 , n37044 , n31603 );
    or g27820 ( n28685 , n29278 , n40157 );
    or g27821 ( n16288 , n16780 , n13428 );
    nor g27822 ( n35562 , n21229 , n7386 );
    not g27823 ( n1970 , n9964 );
    or g27824 ( n26741 , n25628 , n17104 );
    not g27825 ( n31956 , n11409 );
    not g27826 ( n41086 , n27257 );
    or g27827 ( n3731 , n1110 , n37759 );
    or g27828 ( n6128 , n30635 , n10471 );
    xnor g27829 ( n4762 , n9219 , n30904 );
    xnor g27830 ( n34375 , n18678 , n42263 );
    and g27831 ( n16223 , n179 , n2480 );
    or g27832 ( n929 , n19486 , n42327 );
    and g27833 ( n18399 , n13107 , n29364 );
    nor g27834 ( n3196 , n14707 , n27709 );
    not g27835 ( n12085 , n42032 );
    or g27836 ( n15126 , n32125 , n8847 );
    and g27837 ( n30775 , n39623 , n22356 );
    and g27838 ( n3359 , n14946 , n6682 );
    or g27839 ( n2326 , n19391 , n27562 );
    xnor g27840 ( n32536 , n23663 , n11943 );
    nor g27841 ( n36443 , n40080 , n4483 );
    or g27842 ( n6561 , n28149 , n37030 );
    and g27843 ( n40422 , n25160 , n18304 );
    xnor g27844 ( n41303 , n34731 , n32884 );
    not g27845 ( n21175 , n27506 );
    xnor g27846 ( n36633 , n32643 , n22960 );
    and g27847 ( n8595 , n39985 , n20537 );
    not g27848 ( n19217 , n16097 );
    and g27849 ( n38348 , n28232 , n26960 );
    xnor g27850 ( n24355 , n32850 , n20377 );
    or g27851 ( n32946 , n40489 , n34569 );
    or g27852 ( n16673 , n39556 , n33973 );
    not g27853 ( n32090 , n25665 );
    or g27854 ( n23843 , n6558 , n32483 );
    and g27855 ( n15265 , n7272 , n23536 );
    and g27856 ( n30316 , n13855 , n22192 );
    not g27857 ( n41439 , n20322 );
    not g27858 ( n35752 , n3749 );
    not g27859 ( n34293 , n12986 );
    or g27860 ( n14045 , n13123 , n15479 );
    not g27861 ( n12487 , n40499 );
    and g27862 ( n1930 , n31297 , n11502 );
    not g27863 ( n15133 , n25067 );
    xnor g27864 ( n10376 , n18466 , n19224 );
    not g27865 ( n32534 , n9062 );
    nor g27866 ( n19865 , n31378 , n37565 );
    and g27867 ( n15484 , n11226 , n26465 );
    or g27868 ( n3341 , n6182 , n31927 );
    not g27869 ( n29117 , n41457 );
    and g27870 ( n35758 , n2318 , n16038 );
    xnor g27871 ( n6647 , n24998 , n25460 );
    not g27872 ( n4416 , n1419 );
    or g27873 ( n32717 , n33383 , n28986 );
    not g27874 ( n39120 , n27516 );
    not g27875 ( n39752 , n36290 );
    xnor g27876 ( n32206 , n21051 , n21549 );
    nor g27877 ( n5194 , n32327 , n16234 );
    nor g27878 ( n35082 , n14471 , n12008 );
    nor g27879 ( n17560 , n16866 , n42202 );
    not g27880 ( n5258 , n36809 );
    and g27881 ( n27603 , n31126 , n7680 );
    and g27882 ( n35115 , n24769 , n7420 );
    xnor g27883 ( n35897 , n23944 , n12395 );
    xnor g27884 ( n26422 , n10612 , n31828 );
    or g27885 ( n21394 , n32147 , n13386 );
    or g27886 ( n17873 , n14707 , n8881 );
    or g27887 ( n6226 , n4807 , n21578 );
    not g27888 ( n17609 , n27479 );
    or g27889 ( n480 , n1938 , n33243 );
    not g27890 ( n24732 , n24659 );
    or g27891 ( n27248 , n33623 , n13866 );
    not g27892 ( n21514 , n18811 );
    and g27893 ( n16379 , n34003 , n32936 );
    or g27894 ( n41912 , n34565 , n22919 );
    nor g27895 ( n39288 , n20039 , n5847 );
    or g27896 ( n37068 , n30472 , n34728 );
    or g27897 ( n27479 , n34481 , n5188 );
    or g27898 ( n39010 , n14023 , n31660 );
    nor g27899 ( n41 , n35711 , n40473 );
    xnor g27900 ( n13224 , n25042 , n26654 );
    nor g27901 ( n39001 , n18924 , n690 );
    and g27902 ( n11196 , n42005 , n24458 );
    not g27903 ( n11798 , n1214 );
    or g27904 ( n36262 , n11404 , n42518 );
    and g27905 ( n25478 , n6475 , n25276 );
    or g27906 ( n17133 , n14049 , n34338 );
    or g27907 ( n41125 , n33904 , n42002 );
    nor g27908 ( n14689 , n25172 , n20901 );
    and g27909 ( n12379 , n9052 , n16135 );
    and g27910 ( n39276 , n6821 , n8509 );
    nor g27911 ( n20590 , n22904 , n5206 );
    or g27912 ( n25894 , n42885 , n31489 );
    or g27913 ( n40365 , n35915 , n34096 );
    not g27914 ( n16620 , n1681 );
    and g27915 ( n17394 , n23729 , n35354 );
    or g27916 ( n16445 , n38309 , n42911 );
    xnor g27917 ( n3141 , n11023 , n7878 );
    or g27918 ( n5738 , n14471 , n6110 );
    or g27919 ( n9236 , n550 , n2899 );
    xnor g27920 ( n26181 , n37176 , n39152 );
    nor g27921 ( n3464 , n18218 , n2243 );
    and g27922 ( n23140 , n4988 , n28124 );
    or g27923 ( n24795 , n16096 , n4979 );
    not g27924 ( n8559 , n25381 );
    or g27925 ( n33126 , n1075 , n1608 );
    or g27926 ( n23037 , n28143 , n34172 );
    or g27927 ( n27790 , n31524 , n32241 );
    not g27928 ( n27907 , n25247 );
    or g27929 ( n40906 , n27784 , n31753 );
    or g27930 ( n35894 , n1452 , n34368 );
    or g27931 ( n33952 , n16109 , n15863 );
    and g27932 ( n37015 , n1919 , n2716 );
    and g27933 ( n6044 , n36829 , n19187 );
    not g27934 ( n2655 , n37630 );
    and g27935 ( n12606 , n18739 , n3041 );
    or g27936 ( n13878 , n4085 , n13528 );
    nor g27937 ( n2341 , n31256 , n22797 );
    not g27938 ( n4470 , n30738 );
    or g27939 ( n24430 , n15282 , n17166 );
    not g27940 ( n6510 , n20832 );
    or g27941 ( n17607 , n11612 , n31475 );
    xnor g27942 ( n33898 , n32779 , n7094 );
    xnor g27943 ( n24748 , n174 , n38763 );
    or g27944 ( n39857 , n1971 , n25522 );
    and g27945 ( n20287 , n25619 , n10089 );
    not g27946 ( n29395 , n6065 );
    and g27947 ( n21442 , n28811 , n11659 );
    and g27948 ( n2055 , n5387 , n34940 );
    not g27949 ( n29968 , n27063 );
    nor g27950 ( n19825 , n39874 , n3942 );
    or g27951 ( n23023 , n35866 , n29381 );
    not g27952 ( n21178 , n25853 );
    not g27953 ( n20103 , n41680 );
    not g27954 ( n23031 , n14252 );
    not g27955 ( n33815 , n16397 );
    or g27956 ( n21389 , n25782 , n18056 );
    and g27957 ( n21393 , n16859 , n24570 );
    and g27958 ( n30051 , n31116 , n16026 );
    and g27959 ( n36504 , n25548 , n17402 );
    nor g27960 ( n30373 , n37868 , n20003 );
    not g27961 ( n10405 , n40896 );
    or g27962 ( n12246 , n29968 , n26914 );
    nor g27963 ( n3037 , n27031 , n21688 );
    not g27964 ( n35727 , n14471 );
    or g27965 ( n38259 , n22427 , n27601 );
    xnor g27966 ( n10221 , n29740 , n15167 );
    nor g27967 ( n33625 , n4084 , n32051 );
    nor g27968 ( n7933 , n32783 , n34129 );
    or g27969 ( n2960 , n41752 , n13501 );
    not g27970 ( n41789 , n2133 );
    or g27971 ( n12502 , n4492 , n26934 );
    and g27972 ( n11144 , n24485 , n12076 );
    or g27973 ( n26584 , n1459 , n31156 );
    or g27974 ( n41934 , n7430 , n32194 );
    or g27975 ( n32434 , n32610 , n25425 );
    or g27976 ( n21540 , n9185 , n21278 );
    or g27977 ( n5505 , n7410 , n40412 );
    nor g27978 ( n3528 , n39622 , n23316 );
    nor g27979 ( n30533 , n19515 , n30697 );
    nor g27980 ( n30585 , n19547 , n13381 );
    nor g27981 ( n1159 , n562 , n17304 );
    or g27982 ( n1587 , n25566 , n11601 );
    and g27983 ( n3477 , n12093 , n30609 );
    and g27984 ( n7647 , n767 , n27617 );
    and g27985 ( n24479 , n9132 , n12533 );
    or g27986 ( n34350 , n29049 , n34034 );
    and g27987 ( n28989 , n10663 , n29277 );
    or g27988 ( n22644 , n30168 , n12414 );
    or g27989 ( n4721 , n4803 , n17229 );
    and g27990 ( n32857 , n4834 , n19238 );
    xnor g27991 ( n1539 , n12885 , n13528 );
    or g27992 ( n11606 , n13174 , n2592 );
    not g27993 ( n8012 , n25987 );
    nor g27994 ( n28256 , n5896 , n5567 );
    and g27995 ( n23540 , n4250 , n31404 );
    and g27996 ( n12676 , n31295 , n5503 );
    or g27997 ( n5361 , n32801 , n25310 );
    and g27998 ( n4829 , n8096 , n2422 );
    not g27999 ( n37569 , n23195 );
    or g28000 ( n27688 , n5928 , n3659 );
    not g28001 ( n32245 , n6557 );
    not g28002 ( n31822 , n11828 );
    not g28003 ( n23878 , n19757 );
    or g28004 ( n9294 , n34565 , n20492 );
    or g28005 ( n29819 , n24758 , n41259 );
    or g28006 ( n1979 , n4854 , n29318 );
    nor g28007 ( n26040 , n18866 , n14894 );
    nor g28008 ( n31199 , n36117 , n2811 );
    and g28009 ( n9918 , n17058 , n40285 );
    or g28010 ( n27638 , n975 , n8238 );
    not g28011 ( n3432 , n17354 );
    and g28012 ( n36946 , n31039 , n40647 );
    and g28013 ( n18844 , n2695 , n2775 );
    xnor g28014 ( n42698 , n21888 , n19376 );
    or g28015 ( n556 , n1404 , n31252 );
    and g28016 ( n4131 , n26213 , n636 );
    and g28017 ( n31109 , n10158 , n8961 );
    not g28018 ( n24023 , n9682 );
    nor g28019 ( n35767 , n34886 , n39239 );
    and g28020 ( n13482 , n5289 , n39809 );
    or g28021 ( n13875 , n21898 , n41813 );
    or g28022 ( n35410 , n18032 , n1995 );
    and g28023 ( n6431 , n2083 , n32634 );
    or g28024 ( n31645 , n30086 , n10045 );
    and g28025 ( n35208 , n21459 , n3363 );
    and g28026 ( n16390 , n5751 , n41700 );
    and g28027 ( n12425 , n30260 , n18147 );
    or g28028 ( n18783 , n24438 , n11655 );
    or g28029 ( n7905 , n14258 , n21123 );
    nor g28030 ( n22463 , n24115 , n33473 );
    or g28031 ( n30736 , n16598 , n8205 );
    or g28032 ( n25835 , n23204 , n42372 );
    nor g28033 ( n12751 , n31969 , n41798 );
    or g28034 ( n26148 , n34825 , n16751 );
    nor g28035 ( n41544 , n14753 , n34736 );
    and g28036 ( n3943 , n31749 , n19439 );
    and g28037 ( n14847 , n13812 , n21651 );
    or g28038 ( n14866 , n16211 , n11890 );
    xnor g28039 ( n35967 , n1464 , n27080 );
    and g28040 ( n30090 , n30111 , n39574 );
    and g28041 ( n2178 , n27838 , n20930 );
    and g28042 ( n3170 , n22403 , n18356 );
    not g28043 ( n10810 , n41025 );
    nor g28044 ( n14354 , n36823 , n35275 );
    xnor g28045 ( n5266 , n40958 , n10683 );
    or g28046 ( n4591 , n31932 , n36453 );
    or g28047 ( n37651 , n40713 , n38402 );
    not g28048 ( n16885 , n23004 );
    or g28049 ( n7353 , n20338 , n1975 );
    or g28050 ( n20651 , n1524 , n35915 );
    or g28051 ( n41680 , n16271 , n41178 );
    not g28052 ( n8901 , n14463 );
    or g28053 ( n1883 , n5071 , n11364 );
    or g28054 ( n1392 , n33485 , n19329 );
    or g28055 ( n42592 , n14539 , n14398 );
    nor g28056 ( n21469 , n21286 , n6904 );
    or g28057 ( n42380 , n12700 , n40097 );
    not g28058 ( n3747 , n16796 );
    or g28059 ( n14619 , n2684 , n25324 );
    and g28060 ( n35019 , n5919 , n40234 );
    not g28061 ( n35145 , n9614 );
    not g28062 ( n27241 , n38918 );
    or g28063 ( n39916 , n20351 , n34910 );
    nor g28064 ( n19755 , n16598 , n3518 );
    nor g28065 ( n10070 , n30076 , n19403 );
    or g28066 ( n33186 , n32974 , n440 );
    xnor g28067 ( n19345 , n25354 , n28277 );
    nor g28068 ( n17513 , n21476 , n2732 );
    and g28069 ( n22436 , n32106 , n29167 );
    or g28070 ( n32565 , n18028 , n42479 );
    or g28071 ( n21763 , n28565 , n1415 );
    and g28072 ( n14137 , n29523 , n8923 );
    or g28073 ( n40364 , n32800 , n42511 );
    nor g28074 ( n3338 , n27011 , n39370 );
    xnor g28075 ( n1466 , n22842 , n32247 );
    xnor g28076 ( n30180 , n38679 , n3302 );
    and g28077 ( n13343 , n2706 , n24579 );
    or g28078 ( n4774 , n38861 , n21628 );
    or g28079 ( n24728 , n34287 , n10646 );
    and g28080 ( n8772 , n1350 , n40890 );
    or g28081 ( n30981 , n11629 , n8740 );
    not g28082 ( n9702 , n8133 );
    xnor g28083 ( n28497 , n27907 , n14998 );
    or g28084 ( n33554 , n30406 , n40393 );
    or g28085 ( n5392 , n32711 , n23607 );
    or g28086 ( n4035 , n19020 , n28471 );
    or g28087 ( n2158 , n32652 , n10125 );
    xnor g28088 ( n20485 , n19183 , n30328 );
    and g28089 ( n1274 , n32297 , n12507 );
    xnor g28090 ( n36337 , n31840 , n4140 );
    nor g28091 ( n41286 , n8648 , n8055 );
    and g28092 ( n24070 , n9041 , n28478 );
    and g28093 ( n21545 , n17263 , n1545 );
    xnor g28094 ( n35865 , n6625 , n13212 );
    not g28095 ( n29271 , n8463 );
    and g28096 ( n34490 , n35154 , n32296 );
    or g28097 ( n42089 , n20788 , n39579 );
    nor g28098 ( n385 , n8894 , n13922 );
    not g28099 ( n6527 , n10793 );
    and g28100 ( n8674 , n33246 , n3607 );
    and g28101 ( n42766 , n28511 , n32392 );
    xnor g28102 ( n36093 , n8638 , n2312 );
    and g28103 ( n35140 , n14230 , n6630 );
    and g28104 ( n39184 , n36321 , n664 );
    nor g28105 ( n38296 , n19328 , n16708 );
    xnor g28106 ( n23063 , n36615 , n1330 );
    not g28107 ( n11391 , n25795 );
    not g28108 ( n41601 , n3315 );
    not g28109 ( n14280 , n5819 );
    not g28110 ( n26194 , n24026 );
    not g28111 ( n12814 , n30158 );
    and g28112 ( n32237 , n30339 , n400 );
    or g28113 ( n6918 , n3818 , n41990 );
    and g28114 ( n21413 , n33413 , n27040 );
    nor g28115 ( n35639 , n11812 , n4327 );
    or g28116 ( n5838 , n37009 , n25141 );
    or g28117 ( n34680 , n28920 , n15342 );
    xnor g28118 ( n29331 , n9180 , n38633 );
    nor g28119 ( n24644 , n6727 , n34613 );
    xnor g28120 ( n1797 , n32463 , n25608 );
    or g28121 ( n8841 , n24068 , n10263 );
    xnor g28122 ( n34932 , n9619 , n25689 );
    or g28123 ( n11141 , n41601 , n42651 );
    or g28124 ( n22769 , n1507 , n39310 );
    nor g28125 ( n30206 , n3015 , n5726 );
    nor g28126 ( n34238 , n13773 , n29739 );
    or g28127 ( n28466 , n32609 , n11327 );
    and g28128 ( n35715 , n41511 , n19022 );
    not g28129 ( n59 , n41992 );
    or g28130 ( n3938 , n26538 , n29588 );
    not g28131 ( n42803 , n29271 );
    nor g28132 ( n20928 , n13173 , n17861 );
    or g28133 ( n9872 , n17001 , n37828 );
    and g28134 ( n37384 , n30431 , n13950 );
    or g28135 ( n26026 , n11969 , n26570 );
    or g28136 ( n17274 , n29329 , n27131 );
    and g28137 ( n26495 , n42373 , n33799 );
    or g28138 ( n33501 , n35294 , n27164 );
    nor g28139 ( n36774 , n31934 , n41016 );
    or g28140 ( n36589 , n27123 , n12768 );
    or g28141 ( n26682 , n17086 , n39347 );
    not g28142 ( n36238 , n20982 );
    xnor g28143 ( n42679 , n19700 , n37340 );
    or g28144 ( n30105 , n5195 , n23494 );
    and g28145 ( n1210 , n13636 , n2300 );
    or g28146 ( n9446 , n32325 , n14489 );
    or g28147 ( n33339 , n25448 , n19788 );
    or g28148 ( n13719 , n16106 , n12627 );
    and g28149 ( n20382 , n194 , n38628 );
    or g28150 ( n13387 , n35336 , n35695 );
    or g28151 ( n26450 , n9044 , n803 );
    or g28152 ( n35092 , n41717 , n31497 );
    or g28153 ( n28409 , n37662 , n27827 );
    nor g28154 ( n33616 , n20952 , n36417 );
    not g28155 ( n8099 , n30939 );
    or g28156 ( n28037 , n28590 , n42645 );
    or g28157 ( n4888 , n30470 , n30822 );
    or g28158 ( n12819 , n4778 , n4874 );
    or g28159 ( n33651 , n15748 , n12867 );
    not g28160 ( n12162 , n23718 );
    nor g28161 ( n2967 , n42468 , n32528 );
    or g28162 ( n31804 , n7142 , n15875 );
    xnor g28163 ( n15183 , n18066 , n129 );
    nor g28164 ( n1025 , n33051 , n10397 );
    or g28165 ( n29678 , n14945 , n2559 );
    or g28166 ( n13321 , n31307 , n34195 );
    or g28167 ( n8259 , n14407 , n41916 );
    or g28168 ( n42795 , n35732 , n28216 );
    and g28169 ( n42491 , n13023 , n32162 );
    or g28170 ( n2908 , n36396 , n22427 );
    or g28171 ( n19528 , n19494 , n26161 );
    not g28172 ( n41526 , n33626 );
    xnor g28173 ( n7948 , n11845 , n33996 );
    not g28174 ( n8103 , n38258 );
    and g28175 ( n40229 , n29443 , n12849 );
    xnor g28176 ( n18341 , n31099 , n23924 );
    not g28177 ( n27762 , n1568 );
    and g28178 ( n1266 , n31251 , n9220 );
    nor g28179 ( n25010 , n18997 , n8234 );
    nor g28180 ( n11117 , n1691 , n18614 );
    xnor g28181 ( n26712 , n36932 , n39825 );
    or g28182 ( n21198 , n29058 , n29240 );
    not g28183 ( n42204 , n18524 );
    nor g28184 ( n31132 , n14707 , n11048 );
    xnor g28185 ( n18095 , n33100 , n9386 );
    nor g28186 ( n18789 , n22538 , n3690 );
    and g28187 ( n35989 , n39217 , n18098 );
    and g28188 ( n21155 , n19125 , n36830 );
    xnor g28189 ( n31325 , n24390 , n26030 );
    or g28190 ( n15760 , n38463 , n17340 );
    or g28191 ( n24596 , n17193 , n39731 );
    or g28192 ( n31167 , n11128 , n15337 );
    not g28193 ( n28403 , n13994 );
    and g28194 ( n20629 , n37391 , n19821 );
    xnor g28195 ( n32033 , n32160 , n37996 );
    and g28196 ( n743 , n31707 , n33720 );
    or g28197 ( n35508 , n38192 , n21028 );
    nor g28198 ( n37273 , n36667 , n28044 );
    not g28199 ( n29323 , n32485 );
    or g28200 ( n11858 , n5140 , n19962 );
    not g28201 ( n11713 , n1842 );
    or g28202 ( n13693 , n36313 , n14955 );
    and g28203 ( n20243 , n3966 , n35837 );
    and g28204 ( n11650 , n2030 , n16749 );
    and g28205 ( n19963 , n38602 , n38832 );
    and g28206 ( n28737 , n32251 , n22621 );
    and g28207 ( n17385 , n12889 , n30257 );
    not g28208 ( n34972 , n25594 );
    xnor g28209 ( n30285 , n19037 , n9613 );
    xnor g28210 ( n32807 , n11023 , n8086 );
    xnor g28211 ( n7187 , n13461 , n32806 );
    or g28212 ( n16937 , n5140 , n12831 );
    xnor g28213 ( n19448 , n25619 , n14700 );
    or g28214 ( n25006 , n37853 , n4552 );
    or g28215 ( n23690 , n18083 , n26760 );
    and g28216 ( n3642 , n23580 , n35979 );
    and g28217 ( n35275 , n38439 , n38480 );
    or g28218 ( n16571 , n27669 , n26922 );
    nor g28219 ( n25590 , n30764 , n19963 );
    and g28220 ( n6730 , n41763 , n25734 );
    and g28221 ( n36379 , n30803 , n23647 );
    or g28222 ( n18241 , n17464 , n11814 );
    or g28223 ( n10702 , n24917 , n6019 );
    xnor g28224 ( n34115 , n6957 , n37180 );
    and g28225 ( n35554 , n7095 , n13956 );
    xnor g28226 ( n11046 , n20245 , n22517 );
    or g28227 ( n22700 , n12375 , n6170 );
    and g28228 ( n30355 , n7208 , n97 );
    or g28229 ( n18229 , n7439 , n39995 );
    or g28230 ( n42009 , n41433 , n4853 );
    or g28231 ( n22933 , n1619 , n15900 );
    xnor g28232 ( n30338 , n29395 , n34371 );
    and g28233 ( n19737 , n18760 , n23257 );
    not g28234 ( n20416 , n27476 );
    or g28235 ( n20266 , n42615 , n15006 );
    or g28236 ( n19357 , n23902 , n3417 );
    or g28237 ( n984 , n9876 , n35531 );
    and g28238 ( n37289 , n9699 , n6207 );
    nor g28239 ( n23331 , n5187 , n4592 );
    nor g28240 ( n30460 , n1526 , n1594 );
    nor g28241 ( n27488 , n40210 , n26330 );
    or g28242 ( n23485 , n16208 , n12149 );
    not g28243 ( n10558 , n38661 );
    or g28244 ( n39565 , n41923 , n23013 );
    nor g28245 ( n28061 , n16598 , n3569 );
    or g28246 ( n20758 , n8713 , n29270 );
    or g28247 ( n5691 , n40102 , n5910 );
    not g28248 ( n6268 , n31604 );
    or g28249 ( n6964 , n31261 , n23641 );
    not g28250 ( n4706 , n24860 );
    xnor g28251 ( n40500 , n15010 , n40714 );
    or g28252 ( n2413 , n14775 , n1558 );
    or g28253 ( n26184 , n14939 , n23489 );
    nor g28254 ( n21487 , n9482 , n26430 );
    or g28255 ( n29894 , n19036 , n28239 );
    or g28256 ( n25731 , n6743 , n41938 );
    or g28257 ( n16755 , n2164 , n41885 );
    or g28258 ( n12313 , n7704 , n5332 );
    not g28259 ( n23732 , n9546 );
    not g28260 ( n41117 , n13409 );
    not g28261 ( n30264 , n26919 );
    not g28262 ( n40662 , n29640 );
    and g28263 ( n6686 , n19155 , n32649 );
    not g28264 ( n7471 , n32055 );
    not g28265 ( n6490 , n33692 );
    or g28266 ( n11345 , n23614 , n42734 );
    not g28267 ( n14882 , n37186 );
    or g28268 ( n39677 , n16491 , n37779 );
    or g28269 ( n10261 , n14192 , n32032 );
    nor g28270 ( n20478 , n29296 , n41820 );
    xnor g28271 ( n35786 , n6625 , n25803 );
    not g28272 ( n35966 , n18142 );
    or g28273 ( n40535 , n22253 , n40111 );
    not g28274 ( n39058 , n37336 );
    or g28275 ( n29887 , n16791 , n27053 );
    or g28276 ( n18370 , n15487 , n21250 );
    not g28277 ( n31950 , n7069 );
    or g28278 ( n18569 , n5808 , n17340 );
    xnor g28279 ( n802 , n13444 , n36796 );
    not g28280 ( n38424 , n12967 );
    and g28281 ( n5220 , n33258 , n40034 );
    or g28282 ( n31392 , n42425 , n29653 );
    nor g28283 ( n24759 , n14381 , n39394 );
    nor g28284 ( n22235 , n34387 , n42160 );
    or g28285 ( n11174 , n20701 , n29856 );
    and g28286 ( n18426 , n26266 , n22284 );
    or g28287 ( n2931 , n10247 , n34174 );
    and g28288 ( n1790 , n36066 , n18015 );
    nor g28289 ( n31185 , n38251 , n7719 );
    and g28290 ( n1429 , n23010 , n7729 );
    or g28291 ( n316 , n1317 , n33464 );
    or g28292 ( n38027 , n10118 , n3691 );
    or g28293 ( n37649 , n1575 , n7860 );
    or g28294 ( n42027 , n35651 , n7689 );
    or g28295 ( n7770 , n38727 , n14053 );
    xnor g28296 ( n7883 , n40543 , n34292 );
    not g28297 ( n8044 , n26432 );
    not g28298 ( n26825 , n21154 );
    not g28299 ( n40323 , n29711 );
    not g28300 ( n14796 , n6341 );
    and g28301 ( n23648 , n1778 , n17710 );
    and g28302 ( n35515 , n39374 , n39670 );
    or g28303 ( n14253 , n13790 , n15561 );
    not g28304 ( n31674 , n37811 );
    or g28305 ( n40089 , n14262 , n38196 );
    or g28306 ( n18570 , n26481 , n42328 );
    or g28307 ( n3793 , n3433 , n20458 );
    not g28308 ( n39571 , n26902 );
    or g28309 ( n16790 , n9931 , n12198 );
    or g28310 ( n21191 , n29295 , n21966 );
    or g28311 ( n39207 , n8774 , n25704 );
    or g28312 ( n41836 , n20932 , n4112 );
    nor g28313 ( n9303 , n8611 , n38931 );
    or g28314 ( n6626 , n15899 , n36904 );
    or g28315 ( n18545 , n5507 , n17704 );
    not g28316 ( n22224 , n8190 );
    or g28317 ( n17732 , n41439 , n30136 );
    nor g28318 ( n11299 , n22433 , n33001 );
    and g28319 ( n35286 , n13900 , n5074 );
    and g28320 ( n27837 , n4334 , n28639 );
    nor g28321 ( n26885 , n2199 , n24012 );
    xnor g28322 ( n25556 , n13261 , n34720 );
    nor g28323 ( n26270 , n32710 , n15862 );
    and g28324 ( n28707 , n21379 , n6386 );
    and g28325 ( n813 , n8528 , n12571 );
    and g28326 ( n8318 , n19292 , n23816 );
    or g28327 ( n7247 , n10778 , n23022 );
    xnor g28328 ( n41652 , n6625 , n16784 );
    and g28329 ( n12582 , n33605 , n40552 );
    not g28330 ( n3003 , n3178 );
    and g28331 ( n17230 , n4093 , n25400 );
    xnor g28332 ( n33219 , n21877 , n1414 );
    not g28333 ( n33253 , n6161 );
    or g28334 ( n15139 , n37304 , n3410 );
    and g28335 ( n40206 , n30870 , n34125 );
    or g28336 ( n35064 , n40718 , n38293 );
    and g28337 ( n37742 , n16795 , n15767 );
    nor g28338 ( n31648 , n11845 , n33996 );
    xnor g28339 ( n33455 , n40428 , n1971 );
    or g28340 ( n20197 , n6578 , n40877 );
    or g28341 ( n37345 , n39553 , n36641 );
    nor g28342 ( n18897 , n23033 , n41542 );
    and g28343 ( n2021 , n9731 , n37499 );
    or g28344 ( n4445 , n12251 , n20457 );
    or g28345 ( n28753 , n19700 , n39587 );
    not g28346 ( n22773 , n402 );
    xnor g28347 ( n15296 , n42062 , n42621 );
    and g28348 ( n28088 , n32760 , n34986 );
    nor g28349 ( n41702 , n30420 , n37758 );
    and g28350 ( n8469 , n20223 , n1101 );
    or g28351 ( n10286 , n21558 , n13075 );
    xnor g28352 ( n26294 , n34731 , n8198 );
    or g28353 ( n8695 , n29135 , n16481 );
    nor g28354 ( n163 , n11460 , n39413 );
    xnor g28355 ( n17577 , n25042 , n7547 );
    or g28356 ( n830 , n16338 , n24867 );
    nor g28357 ( n36419 , n32589 , n38623 );
    nor g28358 ( n16648 , n35301 , n41581 );
    or g28359 ( n36987 , n26331 , n7073 );
    and g28360 ( n38222 , n39547 , n35972 );
    and g28361 ( n37867 , n18151 , n6047 );
    nor g28362 ( n29015 , n11448 , n16647 );
    xnor g28363 ( n41190 , n22773 , n31858 );
    or g28364 ( n13039 , n33185 , n37952 );
    and g28365 ( n26708 , n4490 , n23827 );
    and g28366 ( n41072 , n33518 , n23144 );
    nor g28367 ( n13600 , n34686 , n4333 );
    xnor g28368 ( n30883 , n31099 , n4171 );
    or g28369 ( n27991 , n39511 , n10553 );
    nor g28370 ( n15472 , n20345 , n5113 );
    and g28371 ( n42416 , n1474 , n39628 );
    and g28372 ( n16948 , n34820 , n10446 );
    or g28373 ( n11170 , n38149 , n18964 );
    and g28374 ( n36446 , n2598 , n28914 );
    or g28375 ( n21693 , n14806 , n30379 );
    xnor g28376 ( n16351 , n37410 , n7550 );
    or g28377 ( n20187 , n35661 , n31447 );
    nor g28378 ( n13187 , n33314 , n18492 );
    and g28379 ( n38518 , n22178 , n36882 );
    xnor g28380 ( n1530 , n21141 , n38772 );
    and g28381 ( n7373 , n13871 , n24060 );
    and g28382 ( n38876 , n16585 , n39231 );
    or g28383 ( n7108 , n17432 , n39481 );
    nor g28384 ( n36583 , n12808 , n32743 );
    or g28385 ( n6159 , n37785 , n16586 );
    or g28386 ( n27650 , n38186 , n22557 );
    xnor g28387 ( n2816 , n32154 , n23965 );
    nor g28388 ( n30115 , n24443 , n7684 );
    xnor g28389 ( n15275 , n31099 , n866 );
    xnor g28390 ( n18592 , n2488 , n38409 );
    or g28391 ( n607 , n19221 , n33630 );
    or g28392 ( n11161 , n16161 , n14791 );
    and g28393 ( n42540 , n11544 , n20022 );
    not g28394 ( n39714 , n33995 );
    or g28395 ( n12800 , n1882 , n20225 );
    and g28396 ( n8402 , n40453 , n41412 );
    xnor g28397 ( n15386 , n28225 , n13100 );
    or g28398 ( n2681 , n6876 , n5656 );
    not g28399 ( n23234 , n12657 );
    not g28400 ( n17081 , n39337 );
    or g28401 ( n5497 , n39326 , n31156 );
    and g28402 ( n30757 , n38396 , n36691 );
    or g28403 ( n39708 , n18244 , n28168 );
    or g28404 ( n18360 , n37763 , n30356 );
    not g28405 ( n1778 , n39831 );
    not g28406 ( n479 , n3579 );
    not g28407 ( n36868 , n42760 );
    or g28408 ( n34757 , n36998 , n60 );
    not g28409 ( n15035 , n16399 );
    and g28410 ( n855 , n25192 , n26382 );
    and g28411 ( n15729 , n32963 , n38169 );
    and g28412 ( n3538 , n30615 , n37612 );
    nor g28413 ( n37447 , n31256 , n36099 );
    xnor g28414 ( n33162 , n38243 , n31735 );
    not g28415 ( n33002 , n33302 );
    not g28416 ( n41197 , n30555 );
    not g28417 ( n34337 , n21306 );
    or g28418 ( n25269 , n9369 , n5564 );
    not g28419 ( n37616 , n18123 );
    or g28420 ( n26255 , n32498 , n12853 );
    or g28421 ( n23659 , n25964 , n12014 );
    not g28422 ( n16473 , n6984 );
    or g28423 ( n31778 , n2600 , n20338 );
    nor g28424 ( n9438 , n32143 , n4764 );
    or g28425 ( n29248 , n25954 , n36975 );
    not g28426 ( n6547 , n25308 );
    xnor g28427 ( n24191 , n16983 , n8494 );
    or g28428 ( n6144 , n7582 , n8438 );
    not g28429 ( n32667 , n38466 );
    and g28430 ( n38751 , n31541 , n35872 );
    not g28431 ( n25924 , n7156 );
    or g28432 ( n4352 , n15505 , n3220 );
    or g28433 ( n19038 , n38748 , n12706 );
    and g28434 ( n1049 , n14034 , n16632 );
    nor g28435 ( n37304 , n695 , n6601 );
    nor g28436 ( n38273 , n21385 , n26804 );
    not g28437 ( n41468 , n6310 );
    and g28438 ( n34324 , n14914 , n9531 );
    or g28439 ( n5165 , n7226 , n3226 );
    and g28440 ( n23718 , n3716 , n5725 );
    not g28441 ( n39503 , n29415 );
    or g28442 ( n40524 , n40109 , n21217 );
    or g28443 ( n3760 , n36697 , n36536 );
    and g28444 ( n8645 , n36370 , n4707 );
    and g28445 ( n27606 , n10728 , n3017 );
    not g28446 ( n37263 , n26969 );
    and g28447 ( n19526 , n5748 , n8932 );
    not g28448 ( n8401 , n34383 );
    not g28449 ( n7088 , n20055 );
    and g28450 ( n18296 , n12211 , n4284 );
    not g28451 ( n29328 , n25511 );
    or g28452 ( n13596 , n14252 , n21740 );
    or g28453 ( n11095 , n20932 , n32126 );
    and g28454 ( n31374 , n24136 , n30574 );
    nor g28455 ( n23556 , n45 , n31874 );
    not g28456 ( n14954 , n20360 );
    or g28457 ( n30771 , n40350 , n22471 );
    or g28458 ( n30966 , n2748 , n37461 );
    and g28459 ( n36002 , n19611 , n13671 );
    not g28460 ( n14316 , n35838 );
    or g28461 ( n415 , n8619 , n15444 );
    xnor g28462 ( n11379 , n8787 , n9067 );
    xnor g28463 ( n25373 , n40 , n13014 );
    nor g28464 ( n24488 , n7342 , n21791 );
    or g28465 ( n41552 , n33321 , n36103 );
    or g28466 ( n36259 , n19390 , n28554 );
    xnor g28467 ( n34503 , n32865 , n29204 );
    not g28468 ( n28643 , n13105 );
    and g28469 ( n23015 , n4721 , n5870 );
    nor g28470 ( n5672 , n22263 , n6786 );
    or g28471 ( n10426 , n20232 , n27781 );
    xnor g28472 ( n17772 , n5240 , n5263 );
    nor g28473 ( n10380 , n6503 , n14733 );
    xnor g28474 ( n30662 , n33342 , n12134 );
    or g28475 ( n39522 , n3580 , n19344 );
    or g28476 ( n505 , n6451 , n1611 );
    or g28477 ( n27012 , n41534 , n30336 );
    or g28478 ( n16551 , n4139 , n13920 );
    or g28479 ( n36064 , n1078 , n31147 );
    and g28480 ( n12645 , n41154 , n13624 );
    and g28481 ( n40459 , n31610 , n20047 );
    or g28482 ( n2120 , n433 , n12265 );
    not g28483 ( n24352 , n33916 );
    and g28484 ( n26330 , n17711 , n10458 );
    xnor g28485 ( n5642 , n41218 , n28624 );
    not g28486 ( n29884 , n15956 );
    xnor g28487 ( n36452 , n39104 , n14618 );
    not g28488 ( n41487 , n23168 );
    and g28489 ( n23882 , n11578 , n24111 );
    or g28490 ( n21626 , n16837 , n39951 );
    or g28491 ( n24347 , n19358 , n33173 );
    nor g28492 ( n39423 , n28333 , n2559 );
    or g28493 ( n33555 , n11798 , n41888 );
    and g28494 ( n38647 , n17892 , n21441 );
    not g28495 ( n11974 , n25519 );
    and g28496 ( n7646 , n15393 , n39792 );
    and g28497 ( n35179 , n7624 , n31971 );
    or g28498 ( n29213 , n13332 , n24993 );
    xnor g28499 ( n24754 , n21634 , n9913 );
    or g28500 ( n35281 , n37029 , n681 );
    or g28501 ( n33296 , n31032 , n17249 );
    or g28502 ( n30848 , n42906 , n17703 );
    nor g28503 ( n37878 , n24892 , n8150 );
    xnor g28504 ( n23000 , n16055 , n7062 );
    not g28505 ( n39217 , n29163 );
    or g28506 ( n5213 , n5205 , n22224 );
    and g28507 ( n10554 , n14648 , n13289 );
    not g28508 ( n13916 , n29762 );
    and g28509 ( n30610 , n25051 , n25171 );
    nor g28510 ( n20913 , n37124 , n24249 );
    and g28511 ( n27902 , n16352 , n25181 );
    or g28512 ( n28371 , n18214 , n39811 );
    or g28513 ( n32394 , n17370 , n16799 );
    and g28514 ( n31614 , n13210 , n2652 );
    or g28515 ( n37834 , n14707 , n10913 );
    or g28516 ( n20297 , n11786 , n11791 );
    or g28517 ( n29828 , n7841 , n13191 );
    not g28518 ( n28735 , n32713 );
    or g28519 ( n3617 , n5475 , n14088 );
    and g28520 ( n39696 , n39721 , n3127 );
    or g28521 ( n41255 , n21044 , n16239 );
    or g28522 ( n2695 , n36099 , n25394 );
    nor g28523 ( n33703 , n13828 , n35634 );
    nor g28524 ( n40351 , n14144 , n25918 );
    not g28525 ( n6863 , n23167 );
    or g28526 ( n27183 , n20021 , n28763 );
    xnor g28527 ( n15541 , n2868 , n7219 );
    xnor g28528 ( n17228 , n9133 , n1837 );
    not g28529 ( n13994 , n6744 );
    or g28530 ( n20262 , n24114 , n41385 );
    nor g28531 ( n35313 , n37488 , n16903 );
    and g28532 ( n29454 , n30420 , n37758 );
    nor g28533 ( n20517 , n34565 , n88 );
    and g28534 ( n20191 , n6070 , n32227 );
    or g28535 ( n9506 , n16990 , n25959 );
    not g28536 ( n13825 , n13203 );
    and g28537 ( n19687 , n34238 , n26918 );
    and g28538 ( n610 , n5883 , n16044 );
    or g28539 ( n10723 , n7879 , n7711 );
    or g28540 ( n39075 , n6834 , n40651 );
    xnor g28541 ( n31772 , n33231 , n42592 );
    or g28542 ( n31972 , n11798 , n38904 );
    xnor g28543 ( n17443 , n105 , n9876 );
    xnor g28544 ( n38497 , n30752 , n13860 );
    not g28545 ( n25839 , n14584 );
    nor g28546 ( n40235 , n34628 , n29898 );
    or g28547 ( n22483 , n14474 , n21612 );
    nor g28548 ( n8454 , n16662 , n21591 );
    not g28549 ( n25915 , n586 );
    or g28550 ( n38215 , n17101 , n26326 );
    and g28551 ( n11118 , n25884 , n16650 );
    and g28552 ( n2466 , n1781 , n27364 );
    not g28553 ( n38892 , n30548 );
    nor g28554 ( n26807 , n22538 , n34023 );
    and g28555 ( n35224 , n29066 , n34812 );
    and g28556 ( n14201 , n2072 , n41467 );
    xnor g28557 ( n1552 , n37175 , n42787 );
    and g28558 ( n1817 , n19314 , n27991 );
    not g28559 ( n35915 , n36811 );
    not g28560 ( n19262 , n14004 );
    and g28561 ( n20654 , n2157 , n28327 );
    or g28562 ( n18919 , n655 , n1758 );
    or g28563 ( n12346 , n22409 , n8675 );
    and g28564 ( n38857 , n502 , n38859 );
    or g28565 ( n24457 , n16833 , n1404 );
    or g28566 ( n16183 , n37149 , n5529 );
    not g28567 ( n19890 , n36863 );
    and g28568 ( n19619 , n5175 , n10445 );
    and g28569 ( n28598 , n9506 , n40060 );
    and g28570 ( n292 , n28272 , n12339 );
    xnor g28571 ( n17154 , n14242 , n34539 );
    nor g28572 ( n41878 , n28584 , n28977 );
    xnor g28573 ( n16437 , n10564 , n29235 );
    not g28574 ( n17198 , n22454 );
    or g28575 ( n15415 , n17250 , n16873 );
    nor g28576 ( n30364 , n39569 , n9392 );
    xnor g28577 ( n8489 , n36712 , n42755 );
    and g28578 ( n22998 , n21135 , n18890 );
    nor g28579 ( n42135 , n34212 , n38826 );
    xnor g28580 ( n4387 , n31329 , n26703 );
    and g28581 ( n8496 , n21228 , n42277 );
    or g28582 ( n31492 , n10778 , n15400 );
    xnor g28583 ( n39323 , n105 , n42588 );
    or g28584 ( n39637 , n17977 , n4926 );
    or g28585 ( n10753 , n42510 , n21372 );
    or g28586 ( n17076 , n24352 , n11242 );
    nor g28587 ( n29264 , n5416 , n24116 );
    nor g28588 ( n12187 , n9240 , n25109 );
    not g28589 ( n169 , n11867 );
    xnor g28590 ( n38228 , n20811 , n11092 );
    or g28591 ( n17809 , n4842 , n30871 );
    nor g28592 ( n30917 , n1178 , n35515 );
    or g28593 ( n2481 , n14390 , n29045 );
    nor g28594 ( n31782 , n9742 , n16290 );
    or g28595 ( n6008 , n36958 , n31829 );
    and g28596 ( n8381 , n36471 , n29105 );
    nor g28597 ( n38913 , n17744 , n36741 );
    or g28598 ( n578 , n26964 , n21060 );
    or g28599 ( n20346 , n9955 , n40052 );
    and g28600 ( n18826 , n21077 , n13945 );
    and g28601 ( n26065 , n14264 , n12785 );
    and g28602 ( n42537 , n36278 , n38270 );
    or g28603 ( n26034 , n4934 , n14346 );
    not g28604 ( n37664 , n20224 );
    and g28605 ( n23860 , n28773 , n31990 );
    or g28606 ( n5622 , n38412 , n27453 );
    and g28607 ( n3287 , n34376 , n6737 );
    or g28608 ( n17910 , n33877 , n37771 );
    or g28609 ( n10502 , n14763 , n10289 );
    or g28610 ( n37412 , n1788 , n21157 );
    and g28611 ( n36856 , n2417 , n11427 );
    not g28612 ( n22993 , n36950 );
    nor g28613 ( n18155 , n18954 , n17221 );
    or g28614 ( n22494 , n23509 , n13897 );
    nor g28615 ( n19145 , n30734 , n32176 );
    or g28616 ( n29081 , n8021 , n17602 );
    and g28617 ( n33590 , n20128 , n42687 );
    xnor g28618 ( n26742 , n30103 , n32748 );
    nor g28619 ( n4106 , n8494 , n870 );
    xnor g28620 ( n3686 , n12109 , n6089 );
    or g28621 ( n38208 , n5495 , n15573 );
    and g28622 ( n18973 , n12309 , n1876 );
    and g28623 ( n7988 , n35553 , n36761 );
    and g28624 ( n34260 , n7000 , n33845 );
    not g28625 ( n37128 , n36841 );
    xnor g28626 ( n24966 , n15111 , n7279 );
    not g28627 ( n35538 , n29565 );
    not g28628 ( n14821 , n28821 );
    nor g28629 ( n2845 , n13707 , n23132 );
    or g28630 ( n2010 , n10624 , n1540 );
    or g28631 ( n16474 , n18937 , n9569 );
    nor g28632 ( n41540 , n14941 , n30011 );
    or g28633 ( n18044 , n21249 , n31401 );
    or g28634 ( n2926 , n26188 , n16628 );
    or g28635 ( n31476 , n7483 , n13074 );
    or g28636 ( n20253 , n31722 , n34608 );
    not g28637 ( n19248 , n39309 );
    and g28638 ( n10179 , n11929 , n2211 );
    nor g28639 ( n31306 , n6671 , n41385 );
    not g28640 ( n32118 , n2562 );
    or g28641 ( n891 , n33046 , n28913 );
    not g28642 ( n19693 , n17714 );
    or g28643 ( n16750 , n24401 , n319 );
    and g28644 ( n37264 , n17668 , n32524 );
    nor g28645 ( n17456 , n17193 , n42913 );
    or g28646 ( n31893 , n27675 , n2012 );
    and g28647 ( n33719 , n19968 , n42350 );
    or g28648 ( n1528 , n8494 , n15106 );
    xnor g28649 ( n33100 , n1216 , n23675 );
    not g28650 ( n13559 , n28473 );
    and g28651 ( n31697 , n14163 , n8071 );
    not g28652 ( n30822 , n8422 );
    or g28653 ( n22366 , n12807 , n25451 );
    or g28654 ( n26954 , n2575 , n39745 );
    and g28655 ( n13862 , n4925 , n32127 );
    or g28656 ( n24779 , n18576 , n10760 );
    or g28657 ( n4429 , n29645 , n34106 );
    or g28658 ( n37592 , n36090 , n25434 );
    nor g28659 ( n34192 , n5768 , n16472 );
    not g28660 ( n23365 , n20608 );
    or g28661 ( n15408 , n8757 , n33543 );
    and g28662 ( n29354 , n30320 , n25168 );
    or g28663 ( n31638 , n9003 , n1825 );
    nor g28664 ( n11877 , n27762 , n4495 );
    xnor g28665 ( n37137 , n7625 , n4811 );
    or g28666 ( n28384 , n13797 , n25907 );
    or g28667 ( n6607 , n28093 , n38306 );
    or g28668 ( n953 , n19880 , n9805 );
    or g28669 ( n3597 , n5670 , n40314 );
    or g28670 ( n32629 , n19190 , n29526 );
    xnor g28671 ( n34054 , n42022 , n3153 );
    or g28672 ( n38916 , n31781 , n27765 );
    not g28673 ( n22577 , n41969 );
    xnor g28674 ( n19577 , n31099 , n18668 );
    or g28675 ( n24747 , n28488 , n17344 );
    and g28676 ( n41591 , n18066 , n129 );
    or g28677 ( n36236 , n31982 , n29856 );
    or g28678 ( n7472 , n22376 , n37851 );
    and g28679 ( n5555 , n26452 , n25099 );
    and g28680 ( n5482 , n11454 , n5586 );
    xnor g28681 ( n30322 , n29740 , n39093 );
    or g28682 ( n29190 , n15775 , n33467 );
    nor g28683 ( n33210 , n36702 , n33379 );
    or g28684 ( n22377 , n12796 , n22412 );
    nor g28685 ( n3520 , n41856 , n38348 );
    and g28686 ( n20054 , n7025 , n10159 );
    or g28687 ( n14663 , n31841 , n31326 );
    and g28688 ( n7516 , n17213 , n6634 );
    nor g28689 ( n24405 , n25727 , n9012 );
    and g28690 ( n39553 , n26695 , n5801 );
    or g28691 ( n41797 , n9622 , n19442 );
    and g28692 ( n13741 , n37456 , n23578 );
    not g28693 ( n14091 , n32558 );
    or g28694 ( n1187 , n8494 , n31129 );
    and g28695 ( n11478 , n4748 , n17209 );
    nor g28696 ( n14406 , n38742 , n16086 );
    or g28697 ( n26092 , n20280 , n31475 );
    or g28698 ( n40860 , n518 , n25504 );
    and g28699 ( n25215 , n8499 , n14679 );
    and g28700 ( n38633 , n18460 , n14620 );
    xnor g28701 ( n26033 , n12146 , n646 );
    and g28702 ( n7811 , n24439 , n34665 );
    or g28703 ( n40920 , n27020 , n34371 );
    or g28704 ( n11463 , n35294 , n34437 );
    and g28705 ( n28326 , n20151 , n14124 );
    or g28706 ( n11689 , n30979 , n26999 );
    not g28707 ( n16924 , n41523 );
    xnor g28708 ( n28350 , n9079 , n30687 );
    and g28709 ( n5090 , n6939 , n40355 );
    not g28710 ( n42405 , n28517 );
    or g28711 ( n41308 , n17842 , n10306 );
    and g28712 ( n33254 , n11699 , n31800 );
    and g28713 ( n37415 , n33656 , n36601 );
    not g28714 ( n3502 , n21503 );
    not g28715 ( n36369 , n7103 );
    or g28716 ( n23616 , n42870 , n24012 );
    nor g28717 ( n14297 , n30941 , n4740 );
    or g28718 ( n41580 , n33989 , n2057 );
    xnor g28719 ( n32101 , n465 , n33453 );
    or g28720 ( n14020 , n4995 , n29581 );
    nor g28721 ( n30793 , n9793 , n10727 );
    or g28722 ( n11956 , n3242 , n41348 );
    nor g28723 ( n38183 , n19221 , n24305 );
    not g28724 ( n12761 , n34501 );
    nor g28725 ( n13787 , n2292 , n7884 );
    and g28726 ( n18100 , n35011 , n1590 );
    and g28727 ( n27926 , n11020 , n14510 );
    and g28728 ( n1707 , n25872 , n18746 );
    and g28729 ( n18173 , n21384 , n14891 );
    or g28730 ( n8337 , n28228 , n15861 );
    not g28731 ( n35713 , n36942 );
    nor g28732 ( n26529 , n7715 , n31767 );
    not g28733 ( n16251 , n36196 );
    xnor g28734 ( n9630 , n965 , n23138 );
    or g28735 ( n29400 , n14587 , n13031 );
    xnor g28736 ( n2532 , n42515 , n36306 );
    or g28737 ( n18656 , n10852 , n4578 );
    and g28738 ( n2268 , n17154 , n19944 );
    not g28739 ( n19054 , n22426 );
    and g28740 ( n3255 , n37097 , n32218 );
    nor g28741 ( n26237 , n29511 , n317 );
    or g28742 ( n21734 , n15941 , n8500 );
    and g28743 ( n26836 , n13859 , n36286 );
    or g28744 ( n21530 , n4829 , n32661 );
    not g28745 ( n34778 , n42814 );
    or g28746 ( n23639 , n38138 , n21709 );
    and g28747 ( n30034 , n33172 , n9046 );
    not g28748 ( n29308 , n26448 );
    nor g28749 ( n10864 , n19792 , n13999 );
    and g28750 ( n29510 , n8744 , n28268 );
    or g28751 ( n12041 , n25991 , n20853 );
    not g28752 ( n12382 , n7587 );
    not g28753 ( n36539 , n40006 );
    not g28754 ( n12671 , n753 );
    and g28755 ( n39293 , n35062 , n28820 );
    and g28756 ( n32271 , n2238 , n3631 );
    or g28757 ( n5923 , n37843 , n16999 );
    and g28758 ( n39050 , n1494 , n10174 );
    or g28759 ( n41202 , n6373 , n33612 );
    or g28760 ( n30421 , n40311 , n3586 );
    xnor g28761 ( n14613 , n21332 , n11389 );
    not g28762 ( n2846 , n27756 );
    and g28763 ( n9962 , n3732 , n40765 );
    nor g28764 ( n20519 , n164 , n28564 );
    or g28765 ( n8878 , n28013 , n33063 );
    xnor g28766 ( n10465 , n40296 , n24006 );
    nor g28767 ( n2337 , n35711 , n42511 );
    nor g28768 ( n17916 , n25410 , n3814 );
    or g28769 ( n12321 , n16412 , n3001 );
    nor g28770 ( n9581 , n19127 , n9502 );
    or g28771 ( n41716 , n33900 , n41649 );
    xnor g28772 ( n37341 , n13504 , n36117 );
    nor g28773 ( n38881 , n1674 , n38121 );
    or g28774 ( n5060 , n27924 , n34284 );
    nor g28775 ( n37956 , n21424 , n24858 );
    and g28776 ( n5764 , n36581 , n27692 );
    nor g28777 ( n18343 , n35646 , n7324 );
    and g28778 ( n25689 , n4317 , n14576 );
    and g28779 ( n8418 , n32343 , n13874 );
    or g28780 ( n3649 , n27233 , n27921 );
    or g28781 ( n6581 , n39425 , n36975 );
    or g28782 ( n37915 , n37162 , n8938 );
    or g28783 ( n32334 , n16738 , n20722 );
    or g28784 ( n7746 , n39783 , n14489 );
    nor g28785 ( n25672 , n1308 , n26451 );
    and g28786 ( n27178 , n7261 , n12536 );
    or g28787 ( n29274 , n24329 , n15169 );
    nor g28788 ( n27019 , n16106 , n18080 );
    not g28789 ( n2478 , n23279 );
    or g28790 ( n34372 , n17719 , n20589 );
    not g28791 ( n15147 , n10428 );
    or g28792 ( n30619 , n28021 , n3350 );
    and g28793 ( n21365 , n12667 , n29175 );
    and g28794 ( n16101 , n17282 , n40953 );
    nor g28795 ( n15206 , n39266 , n3943 );
    and g28796 ( n5484 , n3725 , n21514 );
    xnor g28797 ( n23117 , n18702 , n3818 );
    and g28798 ( n15690 , n3390 , n26062 );
    and g28799 ( n20168 , n27574 , n20764 );
    or g28800 ( n41808 , n5718 , n18225 );
    and g28801 ( n36858 , n18810 , n17761 );
    and g28802 ( n20098 , n19819 , n5553 );
    not g28803 ( n30961 , n10890 );
    or g28804 ( n28072 , n18889 , n35834 );
    or g28805 ( n39513 , n31731 , n19478 );
    xnor g28806 ( n32006 , n26185 , n7356 );
    xnor g28807 ( n29418 , n7311 , n24707 );
    xnor g28808 ( n32361 , n34731 , n17620 );
    and g28809 ( n15277 , n29157 , n24019 );
    xnor g28810 ( n10811 , n6138 , n13642 );
    or g28811 ( n39492 , n41752 , n11618 );
    xnor g28812 ( n33377 , n39713 , n7099 );
    and g28813 ( n14010 , n39415 , n6721 );
    not g28814 ( n36234 , n12933 );
    xnor g28815 ( n34401 , n36046 , n14836 );
    and g28816 ( n21550 , n11058 , n24601 );
    or g28817 ( n14007 , n13441 , n1586 );
    or g28818 ( n42303 , n1567 , n32036 );
    nor g28819 ( n27698 , n9020 , n14218 );
    and g28820 ( n2394 , n3921 , n39729 );
    or g28821 ( n37514 , n6400 , n12011 );
    or g28822 ( n13691 , n15572 , n23598 );
    and g28823 ( n40431 , n29262 , n16154 );
    or g28824 ( n34940 , n10483 , n31585 );
    or g28825 ( n25518 , n18007 , n8650 );
    or g28826 ( n35846 , n20138 , n27708 );
    not g28827 ( n8167 , n13662 );
    xnor g28828 ( n33415 , n35727 , n37143 );
    or g28829 ( n29171 , n4106 , n37885 );
    or g28830 ( n22323 , n34865 , n1636 );
    not g28831 ( n21969 , n22537 );
    or g28832 ( n11452 , n8401 , n1723 );
    not g28833 ( n18043 , n25482 );
    or g28834 ( n38049 , n34472 , n38331 );
    and g28835 ( n25316 , n37190 , n36273 );
    not g28836 ( n19443 , n33249 );
    or g28837 ( n41504 , n34985 , n42694 );
    xnor g28838 ( n23906 , n27627 , n32483 );
    nor g28839 ( n11142 , n16894 , n9791 );
    or g28840 ( n22549 , n23971 , n23593 );
    or g28841 ( n38357 , n25619 , n28115 );
    nor g28842 ( n8260 , n30347 , n6114 );
    nor g28843 ( n33835 , n14264 , n12785 );
    and g28844 ( n27113 , n23789 , n14778 );
    or g28845 ( n20562 , n10953 , n15601 );
    and g28846 ( n2276 , n18854 , n35542 );
    or g28847 ( n20743 , n35866 , n17499 );
    or g28848 ( n19112 , n6742 , n16129 );
    nor g28849 ( n927 , n17120 , n26276 );
    xnor g28850 ( n9356 , n7621 , n22814 );
    nor g28851 ( n7559 , n8494 , n16948 );
    xnor g28852 ( n30692 , n11220 , n12811 );
    or g28853 ( n1800 , n40127 , n42557 );
    nor g28854 ( n27554 , n36996 , n28737 );
    and g28855 ( n20239 , n6896 , n11605 );
    xnor g28856 ( n14638 , n7489 , n26317 );
    or g28857 ( n23193 , n39331 , n33846 );
    or g28858 ( n12743 , n21697 , n29067 );
    or g28859 ( n42781 , n24949 , n31076 );
    and g28860 ( n26563 , n15412 , n3908 );
    and g28861 ( n13777 , n8872 , n37866 );
    xnor g28862 ( n15022 , n29347 , n31166 );
    nor g28863 ( n25820 , n17120 , n4563 );
    nor g28864 ( n1299 , n22140 , n6695 );
    or g28865 ( n6670 , n5065 , n28042 );
    xnor g28866 ( n17568 , n39887 , n4509 );
    or g28867 ( n40767 , n34799 , n14389 );
    or g28868 ( n4186 , n6419 , n11156 );
    not g28869 ( n16741 , n40466 );
    or g28870 ( n28914 , n6358 , n33184 );
    or g28871 ( n24830 , n37457 , n17696 );
    nor g28872 ( n32228 , n38879 , n20934 );
    or g28873 ( n21786 , n19484 , n24309 );
    not g28874 ( n11220 , n28051 );
    not g28875 ( n16987 , n42707 );
    not g28876 ( n7667 , n29374 );
    not g28877 ( n14272 , n23083 );
    and g28878 ( n35170 , n17100 , n25646 );
    and g28879 ( n32885 , n9270 , n7828 );
    xnor g28880 ( n33577 , n2037 , n28609 );
    or g28881 ( n23207 , n4272 , n37779 );
    or g28882 ( n5882 , n14454 , n20013 );
    xnor g28883 ( n9688 , n25143 , n15011 );
    nor g28884 ( n33465 , n33745 , n7504 );
    not g28885 ( n26116 , n21106 );
    or g28886 ( n9408 , n18010 , n25626 );
    or g28887 ( n25680 , n37136 , n1373 );
    nor g28888 ( n36580 , n33981 , n35503 );
    not g28889 ( n42331 , n2093 );
    and g28890 ( n3414 , n32338 , n28588 );
    nor g28891 ( n8781 , n38390 , n6868 );
    xnor g28892 ( n21595 , n11436 , n24308 );
    or g28893 ( n12079 , n2199 , n15904 );
    nor g28894 ( n35004 , n25334 , n3031 );
    or g28895 ( n5720 , n18866 , n17120 );
    or g28896 ( n30236 , n20588 , n11961 );
    or g28897 ( n24132 , n24496 , n8420 );
    xnor g28898 ( n192 , n12808 , n14980 );
    and g28899 ( n37380 , n15938 , n12469 );
    or g28900 ( n31203 , n19170 , n21023 );
    or g28901 ( n9968 , n15144 , n28711 );
    not g28902 ( n6992 , n33052 );
    or g28903 ( n36916 , n17744 , n8703 );
    not g28904 ( n17275 , n13506 );
    nor g28905 ( n9192 , n19164 , n18758 );
    nor g28906 ( n18465 , n13041 , n1217 );
    nor g28907 ( n170 , n38430 , n27401 );
    not g28908 ( n40366 , n7748 );
    not g28909 ( n6138 , n7999 );
    xnor g28910 ( n26053 , n17378 , n19221 );
    or g28911 ( n15744 , n2379 , n35834 );
    nor g28912 ( n342 , n17427 , n9277 );
    or g28913 ( n7134 , n3781 , n18815 );
    not g28914 ( n10962 , n19248 );
    not g28915 ( n33589 , n26737 );
    not g28916 ( n3248 , n13696 );
    nor g28917 ( n13756 , n22109 , n38864 );
    or g28918 ( n5560 , n36883 , n35713 );
    and g28919 ( n30011 , n10134 , n29678 );
    not g28920 ( n19535 , n1398 );
    xnor g28921 ( n40279 , n16215 , n6521 );
    nor g28922 ( n37677 , n25170 , n38847 );
    or g28923 ( n2480 , n17947 , n40292 );
    xnor g28924 ( n12599 , n25118 , n40401 );
    and g28925 ( n5218 , n7495 , n7819 );
    or g28926 ( n22152 , n21804 , n17542 );
    or g28927 ( n4253 , n38111 , n26149 );
    or g28928 ( n20530 , n25043 , n7845 );
    xnor g28929 ( n4938 , n11436 , n5599 );
    not g28930 ( n15705 , n23166 );
    or g28931 ( n16228 , n18865 , n38024 );
    xnor g28932 ( n17658 , n4021 , n31609 );
    and g28933 ( n24531 , n39500 , n1592 );
    or g28934 ( n6871 , n6828 , n22091 );
    not g28935 ( n34831 , n21166 );
    not g28936 ( n8734 , n6744 );
    or g28937 ( n32613 , n3441 , n40766 );
    and g28938 ( n10249 , n40863 , n26526 );
    xnor g28939 ( n24439 , n22263 , n13327 );
    nor g28940 ( n36432 , n38879 , n866 );
    and g28941 ( n13938 , n36579 , n40672 );
    and g28942 ( n2813 , n30425 , n26929 );
    or g28943 ( n12649 , n5826 , n6881 );
    or g28944 ( n14269 , n40904 , n33363 );
    not g28945 ( n31497 , n23168 );
    or g28946 ( n27583 , n42623 , n23289 );
    or g28947 ( n34219 , n15846 , n14019 );
    nor g28948 ( n4112 , n33656 , n36601 );
    not g28949 ( n28081 , n2543 );
    and g28950 ( n8421 , n37469 , n40187 );
    xnor g28951 ( n13624 , n7980 , n16692 );
    and g28952 ( n10597 , n20805 , n36454 );
    not g28953 ( n19300 , n27086 );
    and g28954 ( n37703 , n15697 , n10547 );
    xnor g28955 ( n9061 , n18338 , n33909 );
    and g28956 ( n35057 , n20289 , n34121 );
    or g28957 ( n28592 , n41534 , n21555 );
    or g28958 ( n21311 , n37064 , n13215 );
    or g28959 ( n33023 , n32798 , n10045 );
    xnor g28960 ( n21034 , n30764 , n39702 );
    or g28961 ( n15463 , n26800 , n32341 );
    and g28962 ( n15080 , n16959 , n37887 );
    nor g28963 ( n6283 , n14707 , n31428 );
    not g28964 ( n1841 , n24876 );
    or g28965 ( n40219 , n10912 , n9918 );
    not g28966 ( n12841 , n30628 );
    xnor g28967 ( n25355 , n11295 , n13603 );
    or g28968 ( n39641 , n10941 , n15514 );
    or g28969 ( n8359 , n7443 , n3415 );
    or g28970 ( n39192 , n18866 , n25061 );
    and g28971 ( n1070 , n6752 , n5222 );
    not g28972 ( n36823 , n31785 );
    not g28973 ( n5940 , n21515 );
    and g28974 ( n41667 , n25469 , n37831 );
    xnor g28975 ( n35055 , n38378 , n24582 );
    xnor g28976 ( n34323 , n9180 , n12972 );
    xnor g28977 ( n30221 , n7943 , n4928 );
    and g28978 ( n20341 , n4678 , n15570 );
    nor g28979 ( n16436 , n28477 , n34263 );
    xnor g28980 ( n30693 , n11103 , n15834 );
    xnor g28981 ( n18614 , n11436 , n12676 );
    or g28982 ( n28669 , n36585 , n12778 );
    and g28983 ( n40168 , n5515 , n20356 );
    or g28984 ( n29391 , n28769 , n15573 );
    or g28985 ( n2810 , n40272 , n14944 );
    and g28986 ( n18811 , n34932 , n31923 );
    or g28987 ( n20738 , n4398 , n27416 );
    nor g28988 ( n12948 , n31873 , n22205 );
    and g28989 ( n22021 , n28582 , n32921 );
    and g28990 ( n8297 , n37145 , n7876 );
    not g28991 ( n22915 , n5915 );
    xnor g28992 ( n35889 , n9250 , n42384 );
    or g28993 ( n40107 , n4552 , n33162 );
    not g28994 ( n41595 , n31267 );
    not g28995 ( n32009 , n7125 );
    or g28996 ( n8800 , n41968 , n11298 );
    or g28997 ( n35383 , n40079 , n17449 );
    and g28998 ( n17469 , n9079 , n21227 );
    and g28999 ( n839 , n2725 , n24080 );
    not g29000 ( n36636 , n32118 );
    or g29001 ( n40290 , n107 , n21565 );
    not g29002 ( n38581 , n28871 );
    not g29003 ( n20735 , n15519 );
    or g29004 ( n18052 , n7201 , n17982 );
    nor g29005 ( n8160 , n34892 , n8287 );
    or g29006 ( n40103 , n21707 , n29028 );
    or g29007 ( n3289 , n7356 , n28869 );
    not g29008 ( n2902 , n33971 );
    or g29009 ( n33325 , n21201 , n2838 );
    not g29010 ( n4404 , n28202 );
    and g29011 ( n21092 , n3012 , n9385 );
    not g29012 ( n4736 , n14022 );
    nor g29013 ( n35803 , n27499 , n8200 );
    or g29014 ( n16014 , n7330 , n28197 );
    and g29015 ( n5911 , n26311 , n32207 );
    or g29016 ( n17519 , n38712 , n18458 );
    or g29017 ( n22902 , n17291 , n30071 );
    xnor g29018 ( n20202 , n14469 , n13806 );
    and g29019 ( n5772 , n36897 , n16721 );
    nor g29020 ( n9107 , n41446 , n4695 );
    xnor g29021 ( n1551 , n13151 , n26204 );
    and g29022 ( n9299 , n37160 , n5489 );
    not g29023 ( n23741 , n3066 );
    not g29024 ( n1743 , n22378 );
    nor g29025 ( n8107 , n5946 , n11442 );
    nor g29026 ( n41162 , n34565 , n30349 );
    or g29027 ( n38971 , n19459 , n30216 );
    not g29028 ( n11897 , n32086 );
    xnor g29029 ( n40388 , n26146 , n20527 );
    not g29030 ( n18962 , n38403 );
    and g29031 ( n3415 , n31630 , n23413 );
    not g29032 ( n34352 , n17131 );
    xnor g29033 ( n40974 , n36998 , n23897 );
    or g29034 ( n20091 , n38266 , n12783 );
    and g29035 ( n12178 , n3081 , n37022 );
    and g29036 ( n16914 , n32541 , n16259 );
    not g29037 ( n9557 , n35093 );
    and g29038 ( n13524 , n14713 , n42237 );
    nor g29039 ( n8506 , n40698 , n32125 );
    xnor g29040 ( n19598 , n28458 , n14687 );
    xnor g29041 ( n19168 , n23744 , n14707 );
    not g29042 ( n39491 , n33379 );
    and g29043 ( n37708 , n25307 , n12749 );
    or g29044 ( n3090 , n25136 , n31730 );
    or g29045 ( n938 , n4506 , n30394 );
    not g29046 ( n5649 , n8646 );
    not g29047 ( n26998 , n23986 );
    and g29048 ( n42672 , n31062 , n5827 );
    or g29049 ( n28828 , n20168 , n7832 );
    not g29050 ( n35005 , n369 );
    nor g29051 ( n7170 , n15070 , n24740 );
    and g29052 ( n32741 , n14330 , n28493 );
    or g29053 ( n32524 , n12956 , n13112 );
    and g29054 ( n5217 , n5762 , n14118 );
    not g29055 ( n21479 , n3272 );
    and g29056 ( n8593 , n2128 , n41806 );
    or g29057 ( n16145 , n23745 , n31473 );
    or g29058 ( n14066 , n37466 , n3378 );
    or g29059 ( n15872 , n848 , n6970 );
    xnor g29060 ( n28039 , n21823 , n32158 );
    or g29061 ( n28802 , n40346 , n8459 );
    or g29062 ( n5040 , n36044 , n38020 );
    not g29063 ( n25219 , n14064 );
    xnor g29064 ( n36700 , n13358 , n24994 );
    or g29065 ( n7552 , n31214 , n21064 );
    and g29066 ( n452 , n34100 , n27664 );
    not g29067 ( n15004 , n34653 );
    nor g29068 ( n29550 , n7648 , n24116 );
    or g29069 ( n40117 , n29712 , n34728 );
    xnor g29070 ( n25274 , n6625 , n24022 );
    or g29071 ( n35924 , n29026 , n34862 );
    not g29072 ( n13261 , n29457 );
    or g29073 ( n14786 , n4768 , n26631 );
    nor g29074 ( n7436 , n17999 , n2281 );
    not g29075 ( n39408 , n2320 );
    and g29076 ( n22104 , n24963 , n36086 );
    nor g29077 ( n24463 , n23594 , n10335 );
    and g29078 ( n36425 , n9106 , n5333 );
    nor g29079 ( n23806 , n25898 , n8072 );
    or g29080 ( n10442 , n25827 , n11796 );
    xnor g29081 ( n38893 , n41218 , n27017 );
    and g29082 ( n5760 , n10937 , n42106 );
    or g29083 ( n7301 , n28745 , n27978 );
    and g29084 ( n4428 , n32441 , n24980 );
    or g29085 ( n22712 , n26759 , n22952 );
    nor g29086 ( n41757 , n10456 , n15545 );
    or g29087 ( n22939 , n5927 , n39122 );
    not g29088 ( n38466 , n3137 );
    nor g29089 ( n10202 , n38789 , n29348 );
    not g29090 ( n1656 , n17426 );
    or g29091 ( n29888 , n26910 , n34311 );
    nor g29092 ( n14134 , n16211 , n18073 );
    not g29093 ( n26068 , n41416 );
    and g29094 ( n25669 , n10762 , n15057 );
    or g29095 ( n33737 , n30116 , n5984 );
    or g29096 ( n22794 , n14281 , n14716 );
    and g29097 ( n3222 , n4641 , n11046 );
    and g29098 ( n4130 , n35886 , n15060 );
    xnor g29099 ( n16268 , n5073 , n22090 );
    nor g29100 ( n2907 , n35769 , n4562 );
    and g29101 ( n4979 , n33405 , n33524 );
    or g29102 ( n10805 , n20141 , n7442 );
    nor g29103 ( n9610 , n3966 , n35837 );
    and g29104 ( n25486 , n38342 , n1836 );
    and g29105 ( n26582 , n42833 , n1727 );
    not g29106 ( n30857 , n9316 );
    and g29107 ( n35153 , n41115 , n28506 );
    not g29108 ( n39068 , n7125 );
    and g29109 ( n20532 , n29193 , n3779 );
    or g29110 ( n42670 , n14454 , n6387 );
    or g29111 ( n6882 , n40462 , n26250 );
    or g29112 ( n29224 , n22871 , n37633 );
    or g29113 ( n1595 , n37683 , n3916 );
    or g29114 ( n33062 , n38157 , n17434 );
    and g29115 ( n31114 , n14210 , n35537 );
    or g29116 ( n14555 , n31769 , n24653 );
    xnor g29117 ( n29701 , n12806 , n4639 );
    or g29118 ( n29643 , n41526 , n6808 );
    or g29119 ( n39646 , n40710 , n30024 );
    not g29120 ( n33803 , n2279 );
    or g29121 ( n31285 , n31552 , n7172 );
    or g29122 ( n14193 , n36269 , n30225 );
    not g29123 ( n8920 , n13649 );
    or g29124 ( n9914 , n25142 , n8781 );
    and g29125 ( n15996 , n37822 , n5856 );
    nor g29126 ( n7252 , n15232 , n18723 );
    and g29127 ( n40329 , n41537 , n25866 );
    and g29128 ( n37143 , n15829 , n515 );
    or g29129 ( n41610 , n23146 , n24233 );
    nor g29130 ( n26041 , n13336 , n6078 );
    nor g29131 ( n31596 , n41447 , n34853 );
    not g29132 ( n41977 , n14233 );
    xnor g29133 ( n25212 , n105 , n24300 );
    or g29134 ( n32937 , n32818 , n24445 );
    or g29135 ( n13972 , n5795 , n35808 );
    or g29136 ( n20598 , n41325 , n35633 );
    and g29137 ( n2244 , n26084 , n390 );
    nor g29138 ( n18528 , n40163 , n37749 );
    or g29139 ( n41115 , n3914 , n39134 );
    or g29140 ( n28804 , n4352 , n21225 );
    or g29141 ( n9590 , n37539 , n9913 );
    or g29142 ( n11078 , n33847 , n21268 );
    and g29143 ( n36849 , n10711 , n36147 );
    xnor g29144 ( n10176 , n30397 , n21547 );
    or g29145 ( n1276 , n8809 , n33121 );
    or g29146 ( n10444 , n1389 , n3311 );
    not g29147 ( n14365 , n14725 );
    or g29148 ( n13089 , n978 , n42544 );
    or g29149 ( n3250 , n20932 , n40397 );
    not g29150 ( n26902 , n23541 );
    or g29151 ( n24500 , n24656 , n5485 );
    not g29152 ( n2586 , n31433 );
    or g29153 ( n10547 , n40668 , n33671 );
    and g29154 ( n7327 , n3718 , n15673 );
    xnor g29155 ( n3783 , n36094 , n20474 );
    xnor g29156 ( n15983 , n17877 , n26157 );
    not g29157 ( n8021 , n40875 );
    or g29158 ( n33945 , n11735 , n5904 );
    or g29159 ( n25092 , n35287 , n36467 );
    and g29160 ( n6797 , n25764 , n40906 );
    or g29161 ( n37556 , n10460 , n26755 );
    and g29162 ( n9541 , n5272 , n26499 );
    not g29163 ( n25451 , n40600 );
    or g29164 ( n35860 , n19762 , n4766 );
    or g29165 ( n10344 , n328 , n23490 );
    not g29166 ( n21347 , n41969 );
    or g29167 ( n7390 , n40934 , n18363 );
    or g29168 ( n14741 , n31501 , n31361 );
    xnor g29169 ( n15156 , n7004 , n18300 );
    not g29170 ( n29844 , n40861 );
    not g29171 ( n19313 , n12704 );
    or g29172 ( n26404 , n21170 , n20780 );
    xnor g29173 ( n23910 , n9841 , n42294 );
    nor g29174 ( n3959 , n29684 , n21517 );
    not g29175 ( n1516 , n17738 );
    or g29176 ( n27889 , n16910 , n25011 );
    or g29177 ( n39473 , n29233 , n10889 );
    and g29178 ( n15792 , n18896 , n26628 );
    not g29179 ( n18408 , n26858 );
    or g29180 ( n18445 , n10756 , n30293 );
    or g29181 ( n39435 , n2132 , n21764 );
    and g29182 ( n13453 , n41727 , n5157 );
    and g29183 ( n39616 , n17986 , n16184 );
    not g29184 ( n2647 , n4280 );
    not g29185 ( n32794 , n11409 );
    or g29186 ( n39725 , n33744 , n32732 );
    or g29187 ( n3875 , n11957 , n39142 );
    nor g29188 ( n30785 , n5964 , n6613 );
    or g29189 ( n14892 , n32446 , n42183 );
    not g29190 ( n22352 , n32406 );
    not g29191 ( n15537 , n41942 );
    nor g29192 ( n33476 , n3961 , n38503 );
    and g29193 ( n40239 , n15241 , n4184 );
    or g29194 ( n7173 , n11410 , n16840 );
    or g29195 ( n17792 , n13380 , n32290 );
    or g29196 ( n4513 , n21025 , n15550 );
    xnor g29197 ( n38670 , n23090 , n10516 );
    or g29198 ( n22286 , n9457 , n40039 );
    or g29199 ( n37285 , n898 , n22875 );
    or g29200 ( n22317 , n29046 , n29454 );
    not g29201 ( n20498 , n9312 );
    xnor g29202 ( n14212 , n7904 , n26479 );
    xnor g29203 ( n24749 , n33058 , n9095 );
    or g29204 ( n10841 , n41325 , n12198 );
    not g29205 ( n545 , n34931 );
    or g29206 ( n16800 , n16856 , n13687 );
    and g29207 ( n27670 , n1119 , n29415 );
    nor g29208 ( n413 , n2232 , n8146 );
    nor g29209 ( n16799 , n40090 , n34738 );
    and g29210 ( n2172 , n35504 , n953 );
    or g29211 ( n20841 , n14472 , n23096 );
    or g29212 ( n22421 , n29422 , n7229 );
    or g29213 ( n11164 , n19803 , n17502 );
    or g29214 ( n32305 , n36511 , n19411 );
    nor g29215 ( n36719 , n21680 , n8110 );
    not g29216 ( n1470 , n30892 );
    or g29217 ( n35626 , n22272 , n27921 );
    and g29218 ( n16319 , n4749 , n20639 );
    xnor g29219 ( n42301 , n17872 , n34135 );
    or g29220 ( n11888 , n20699 , n24418 );
    and g29221 ( n2152 , n22760 , n19213 );
    not g29222 ( n4937 , n39139 );
    or g29223 ( n16922 , n32170 , n10827 );
    or g29224 ( n7871 , n39059 , n8146 );
    and g29225 ( n12665 , n15142 , n22420 );
    or g29226 ( n20744 , n3004 , n15522 );
    or g29227 ( n35906 , n6011 , n940 );
    or g29228 ( n8304 , n3034 , n9577 );
    or g29229 ( n14906 , n4154 , n22568 );
    or g29230 ( n36758 , n25547 , n34052 );
    nor g29231 ( n39267 , n36117 , n33869 );
    nor g29232 ( n19275 , n10902 , n24840 );
    xnor g29233 ( n29499 , n27789 , n24383 );
    nor g29234 ( n1950 , n9638 , n37324 );
    or g29235 ( n14008 , n36584 , n17756 );
    or g29236 ( n29704 , n4843 , n11305 );
    not g29237 ( n16789 , n10884 );
    or g29238 ( n39227 , n10770 , n39811 );
    or g29239 ( n35316 , n30583 , n25073 );
    or g29240 ( n25513 , n41444 , n21602 );
    not g29241 ( n31300 , n29709 );
    or g29242 ( n41122 , n3954 , n36416 );
    xnor g29243 ( n16965 , n42064 , n12104 );
    or g29244 ( n32275 , n5491 , n10268 );
    or g29245 ( n32196 , n41691 , n29884 );
    and g29246 ( n6745 , n27366 , n3079 );
    and g29247 ( n20406 , n26677 , n26711 );
    and g29248 ( n13565 , n3117 , n23298 );
    or g29249 ( n10262 , n33164 , n6335 );
    or g29250 ( n31297 , n21396 , n30720 );
    or g29251 ( n14344 , n5729 , n33333 );
    xnor g29252 ( n22307 , n5484 , n35264 );
    and g29253 ( n27530 , n21170 , n12507 );
    or g29254 ( n8490 , n9617 , n35731 );
    or g29255 ( n16005 , n19933 , n36917 );
    not g29256 ( n234 , n28565 );
    xnor g29257 ( n17281 , n37953 , n27551 );
    not g29258 ( n8903 , n28839 );
    xnor g29259 ( n19 , n42656 , n39498 );
    or g29260 ( n17684 , n25419 , n2675 );
    or g29261 ( n35659 , n28982 , n21307 );
    or g29262 ( n36978 , n7516 , n30525 );
    and g29263 ( n42665 , n11024 , n4496 );
    or g29264 ( n39876 , n12392 , n24357 );
    or g29265 ( n27846 , n4227 , n33321 );
    and g29266 ( n22003 , n41464 , n25988 );
    not g29267 ( n42871 , n14258 );
    or g29268 ( n12870 , n5910 , n38569 );
    or g29269 ( n29223 , n37434 , n8234 );
    not g29270 ( n40709 , n18147 );
    not g29271 ( n21771 , n42444 );
    or g29272 ( n37743 , n33314 , n9766 );
    not g29273 ( n41048 , n21661 );
    nor g29274 ( n25661 , n36814 , n14249 );
    or g29275 ( n13440 , n21907 , n24506 );
    or g29276 ( n24174 , n35748 , n24614 );
    not g29277 ( n29720 , n23069 );
    or g29278 ( n26390 , n19784 , n24597 );
    and g29279 ( n16247 , n204 , n11043 );
    xnor g29280 ( n6300 , n31099 , n7490 );
    or g29281 ( n22459 , n21705 , n22409 );
    xnor g29282 ( n35808 , n25828 , n28280 );
    not g29283 ( n35289 , n34151 );
    or g29284 ( n3685 , n26317 , n28407 );
    or g29285 ( n15797 , n14707 , n3028 );
    not g29286 ( n32637 , n8093 );
    not g29287 ( n34606 , n34098 );
    not g29288 ( n17659 , n10395 );
    or g29289 ( n32421 , n20728 , n23523 );
    or g29290 ( n31599 , n23073 , n27238 );
    and g29291 ( n40495 , n25717 , n30990 );
    and g29292 ( n14211 , n16297 , n20348 );
    not g29293 ( n15050 , n28836 );
    not g29294 ( n15435 , n29271 );
    not g29295 ( n27780 , n32693 );
    xnor g29296 ( n22051 , n29928 , n2974 );
    or g29297 ( n37701 , n8628 , n23146 );
    or g29298 ( n4521 , n33345 , n29962 );
    or g29299 ( n37036 , n1997 , n29700 );
    or g29300 ( n28459 , n30314 , n7422 );
    or g29301 ( n16726 , n36210 , n35276 );
    or g29302 ( n39041 , n40082 , n12669 );
    xnor g29303 ( n1819 , n669 , n27688 );
    nor g29304 ( n42806 , n30873 , n41077 );
    xnor g29305 ( n4248 , n36009 , n12354 );
    and g29306 ( n11739 , n32625 , n22937 );
    or g29307 ( n19819 , n26948 , n28689 );
    not g29308 ( n27917 , n16690 );
    or g29309 ( n33591 , n38879 , n39216 );
    not g29310 ( n41066 , n9403 );
    and g29311 ( n30371 , n2920 , n6461 );
    nor g29312 ( n42335 , n18951 , n29864 );
    and g29313 ( n17685 , n19037 , n9613 );
    not g29314 ( n4109 , n7984 );
    and g29315 ( n31759 , n14994 , n35299 );
    and g29316 ( n37234 , n38383 , n32052 );
    and g29317 ( n23566 , n14021 , n18461 );
    xnor g29318 ( n19342 , n31177 , n1805 );
    and g29319 ( n12046 , n38788 , n20300 );
    not g29320 ( n30490 , n3265 );
    not g29321 ( n31352 , n19119 );
    or g29322 ( n25752 , n12392 , n27341 );
    or g29323 ( n21830 , n3821 , n4768 );
    or g29324 ( n24208 , n33318 , n13116 );
    or g29325 ( n18617 , n7682 , n38416 );
    nor g29326 ( n25004 , n32900 , n34304 );
    xnor g29327 ( n41164 , n32048 , n7053 );
    not g29328 ( n17680 , n3214 );
    or g29329 ( n31820 , n5896 , n23011 );
    xnor g29330 ( n14653 , n41013 , n27367 );
    or g29331 ( n27901 , n14550 , n3278 );
    xnor g29332 ( n27263 , n38256 , n17548 );
    or g29333 ( n8327 , n7696 , n24254 );
    not g29334 ( n10118 , n42696 );
    xnor g29335 ( n25655 , n42715 , n42908 );
    or g29336 ( n32805 , n30674 , n27947 );
    xnor g29337 ( n16482 , n34731 , n10737 );
    and g29338 ( n30467 , n42031 , n33083 );
    or g29339 ( n8452 , n36424 , n42431 );
    xnor g29340 ( n37830 , n36998 , n3518 );
    or g29341 ( n3064 , n19476 , n37632 );
    or g29342 ( n7744 , n19402 , n12702 );
    or g29343 ( n42324 , n6915 , n31618 );
    or g29344 ( n18943 , n17560 , n30316 );
    not g29345 ( n11881 , n36843 );
    or g29346 ( n13717 , n27914 , n15880 );
    not g29347 ( n27140 , n30033 );
    and g29348 ( n34670 , n28099 , n12323 );
    or g29349 ( n28763 , n35915 , n18823 );
    xnor g29350 ( n39091 , n12007 , n14607 );
    or g29351 ( n41281 , n12232 , n3130 );
    or g29352 ( n19334 , n35922 , n15401 );
    or g29353 ( n15643 , n14287 , n35378 );
    not g29354 ( n4796 , n478 );
    and g29355 ( n21265 , n3163 , n39107 );
    or g29356 ( n3445 , n34565 , n38428 );
    nor g29357 ( n15202 , n9215 , n38907 );
    nor g29358 ( n8701 , n13103 , n39611 );
    or g29359 ( n30989 , n32455 , n40255 );
    or g29360 ( n42579 , n11199 , n6469 );
    and g29361 ( n21377 , n33646 , n7820 );
    nor g29362 ( n42309 , n19772 , n33592 );
    and g29363 ( n16550 , n11249 , n24683 );
    not g29364 ( n28482 , n31827 );
    not g29365 ( n16736 , n16397 );
    nor g29366 ( n27335 , n35780 , n22352 );
    nor g29367 ( n35769 , n5980 , n5287 );
    or g29368 ( n40812 , n34847 , n42160 );
    or g29369 ( n19472 , n36235 , n16103 );
    or g29370 ( n28876 , n31707 , n18006 );
    or g29371 ( n22636 , n23761 , n40961 );
    or g29372 ( n22958 , n42312 , n30142 );
    or g29373 ( n12262 , n4885 , n25924 );
    or g29374 ( n16669 , n30714 , n12456 );
    xnor g29375 ( n21328 , n451 , n32277 );
    nor g29376 ( n32724 , n17182 , n20191 );
    or g29377 ( n18502 , n15388 , n29813 );
    not g29378 ( n15806 , n40263 );
    or g29379 ( n1140 , n14099 , n33354 );
    or g29380 ( n35050 , n40109 , n25778 );
    or g29381 ( n24519 , n16223 , n22981 );
    xnor g29382 ( n28898 , n15058 , n42640 );
    or g29383 ( n21168 , n18748 , n31601 );
    or g29384 ( n31272 , n37980 , n10058 );
    or g29385 ( n26648 , n35294 , n41375 );
    xnor g29386 ( n21797 , n27035 , n14218 );
    nor g29387 ( n17992 , n14707 , n33910 );
    nor g29388 ( n681 , n5334 , n15407 );
    or g29389 ( n37170 , n1451 , n28817 );
    xnor g29390 ( n23908 , n33745 , n5277 );
    xnor g29391 ( n19773 , n39222 , n36614 );
    not g29392 ( n40481 , n27666 );
    nor g29393 ( n22092 , n1338 , n5631 );
    nor g29394 ( n15880 , n36117 , n36244 );
    not g29395 ( n242 , n25164 );
    nor g29396 ( n34019 , n34292 , n8151 );
    and g29397 ( n34148 , n36567 , n34375 );
    and g29398 ( n41736 , n31661 , n19268 );
    and g29399 ( n14077 , n19662 , n29911 );
    or g29400 ( n8488 , n41400 , n14065 );
    and g29401 ( n11951 , n11759 , n4940 );
    or g29402 ( n9993 , n27712 , n23670 );
    not g29403 ( n28283 , n20154 );
    not g29404 ( n24227 , n13355 );
    or g29405 ( n30411 , n3102 , n21788 );
    not g29406 ( n17598 , n7958 );
    or g29407 ( n8129 , n27424 , n39675 );
    and g29408 ( n13255 , n17003 , n34550 );
    not g29409 ( n7706 , n13279 );
    or g29410 ( n18039 , n36897 , n16721 );
    or g29411 ( n29921 , n23931 , n37195 );
    nor g29412 ( n1938 , n3812 , n25909 );
    xnor g29413 ( n70 , n40233 , n38030 );
    nor g29414 ( n24598 , n13345 , n11376 );
    or g29415 ( n21033 , n15078 , n18393 );
    xnor g29416 ( n4217 , n10108 , n17193 );
    or g29417 ( n21917 , n6507 , n18281 );
    not g29418 ( n13054 , n9774 );
    or g29419 ( n36761 , n37849 , n13496 );
    or g29420 ( n23899 , n5645 , n38954 );
    not g29421 ( n35361 , n31785 );
    and g29422 ( n10229 , n35433 , n32188 );
    or g29423 ( n38997 , n42299 , n35216 );
    not g29424 ( n33313 , n12367 );
    nor g29425 ( n38706 , n21253 , n7338 );
    or g29426 ( n21716 , n34762 , n28680 );
    or g29427 ( n3815 , n15050 , n4494 );
    xnor g29428 ( n6241 , n26033 , n23639 );
    nor g29429 ( n7841 , n17120 , n23888 );
    nor g29430 ( n23796 , n5302 , n13709 );
    and g29431 ( n4183 , n40814 , n1035 );
    or g29432 ( n21493 , n25558 , n12058 );
    or g29433 ( n15684 , n27330 , n27540 );
    xnor g29434 ( n31808 , n12787 , n34292 );
    or g29435 ( n11450 , n6806 , n7810 );
    and g29436 ( n14238 , n5626 , n15885 );
    and g29437 ( n33955 , n22231 , n22323 );
    xnor g29438 ( n28303 , n42064 , n6571 );
    or g29439 ( n5825 , n3925 , n21905 );
    or g29440 ( n21161 , n15611 , n35459 );
    nor g29441 ( n2936 , n9796 , n23675 );
    xnor g29442 ( n27883 , n29740 , n924 );
    and g29443 ( n11928 , n17158 , n3321 );
    or g29444 ( n38062 , n31542 , n5265 );
    or g29445 ( n13812 , n14650 , n21170 );
    and g29446 ( n21584 , n8229 , n13831 );
    not g29447 ( n10622 , n29516 );
    not g29448 ( n1455 , n9716 );
    xnor g29449 ( n15394 , n25619 , n10832 );
    not g29450 ( n19845 , n13910 );
    and g29451 ( n34953 , n26045 , n5699 );
    and g29452 ( n32902 , n25926 , n16463 );
    not g29453 ( n6993 , n12178 );
    and g29454 ( n36483 , n9301 , n12080 );
    not g29455 ( n31378 , n8949 );
    xnor g29456 ( n31102 , n20506 , n13543 );
    and g29457 ( n2355 , n16215 , n28638 );
    and g29458 ( n11451 , n492 , n31560 );
    not g29459 ( n12054 , n16582 );
    or g29460 ( n2716 , n17141 , n27891 );
    not g29461 ( n32212 , n25592 );
    and g29462 ( n3635 , n21755 , n29025 );
    or g29463 ( n4418 , n23709 , n34269 );
    or g29464 ( n21566 , n9035 , n5153 );
    and g29465 ( n5204 , n22139 , n7501 );
    or g29466 ( n14221 , n13851 , n18667 );
    or g29467 ( n19875 , n34994 , n29173 );
    or g29468 ( n25217 , n14707 , n1956 );
    not g29469 ( n4543 , n10277 );
    or g29470 ( n28368 , n23141 , n6842 );
    and g29471 ( n31426 , n1232 , n27556 );
    not g29472 ( n33495 , n32509 );
    or g29473 ( n37609 , n15483 , n39924 );
    not g29474 ( n40393 , n24920 );
    not g29475 ( n4296 , n38125 );
    or g29476 ( n41476 , n18102 , n38729 );
    or g29477 ( n10428 , n24152 , n18525 );
    xnor g29478 ( n1623 , n28415 , n11695 );
    or g29479 ( n28455 , n29092 , n7787 );
    or g29480 ( n23814 , n41788 , n17511 );
    or g29481 ( n42176 , n27761 , n343 );
    or g29482 ( n8332 , n14198 , n31736 );
    or g29483 ( n42426 , n21050 , n35216 );
    not g29484 ( n27714 , n14639 );
    and g29485 ( n10769 , n20962 , n42257 );
    xnor g29486 ( n18185 , n16934 , n2266 );
    and g29487 ( n21791 , n28903 , n21622 );
    nor g29488 ( n9795 , n14202 , n42697 );
    nor g29489 ( n5189 , n5964 , n8657 );
    or g29490 ( n20395 , n21096 , n41768 );
    xnor g29491 ( n16677 , n36009 , n1203 );
    not g29492 ( n34153 , n26930 );
    xnor g29493 ( n2118 , n13444 , n12913 );
    nor g29494 ( n41339 , n37494 , n42540 );
    nor g29495 ( n14494 , n25908 , n28237 );
    or g29496 ( n1699 , n27142 , n20054 );
    and g29497 ( n14089 , n10084 , n20309 );
    and g29498 ( n3677 , n25922 , n34808 );
    or g29499 ( n6862 , n28617 , n24416 );
    not g29500 ( n31923 , n2301 );
    and g29501 ( n39152 , n40199 , n8334 );
    nor g29502 ( n14784 , n33935 , n29156 );
    xnor g29503 ( n15150 , n4795 , n2112 );
    and g29504 ( n21746 , n23270 , n28513 );
    or g29505 ( n37748 , n37131 , n41600 );
    or g29506 ( n29352 , n21947 , n1387 );
    or g29507 ( n10705 , n413 , n6192 );
    or g29508 ( n24097 , n25777 , n5341 );
    or g29509 ( n33093 , n25802 , n23695 );
    and g29510 ( n1747 , n3221 , n25809 );
    not g29511 ( n9234 , n14962 );
    xnor g29512 ( n21823 , n22888 , n10068 );
    and g29513 ( n3083 , n3293 , n8985 );
    xnor g29514 ( n16201 , n2339 , n39988 );
    nor g29515 ( n11572 , n36345 , n5509 );
    nor g29516 ( n21854 , n34565 , n15935 );
    xnor g29517 ( n30306 , n19082 , n17120 );
    not g29518 ( n22753 , n1572 );
    or g29519 ( n39987 , n1478 , n12638 );
    or g29520 ( n24896 , n27191 , n41342 );
    not g29521 ( n38511 , n2593 );
    nor g29522 ( n20621 , n3420 , n31858 );
    or g29523 ( n42829 , n38538 , n23201 );
    nor g29524 ( n2614 , n34787 , n14378 );
    or g29525 ( n35613 , n6510 , n29421 );
    not g29526 ( n18622 , n4961 );
    not g29527 ( n21183 , n18807 );
    not g29528 ( n23301 , n21462 );
    not g29529 ( n37625 , n26232 );
    not g29530 ( n32087 , n23369 );
    not g29531 ( n27384 , n26086 );
    or g29532 ( n6668 , n18220 , n37736 );
    or g29533 ( n14510 , n3252 , n23733 );
    xnor g29534 ( n10774 , n17198 , n21319 );
    or g29535 ( n24517 , n7827 , n2012 );
    or g29536 ( n27496 , n9048 , n33206 );
    or g29537 ( n6855 , n36117 , n21217 );
    not g29538 ( n15681 , n3315 );
    xnor g29539 ( n5606 , n35727 , n4666 );
    xnor g29540 ( n4123 , n24210 , n34392 );
    and g29541 ( n11316 , n45 , n31874 );
    nor g29542 ( n2092 , n32793 , n1006 );
    or g29543 ( n12504 , n3939 , n40032 );
    or g29544 ( n8959 , n19469 , n20405 );
    or g29545 ( n21835 , n24292 , n9213 );
    not g29546 ( n2687 , n24603 );
    or g29547 ( n34399 , n38218 , n14764 );
    or g29548 ( n23869 , n36498 , n16838 );
    xnor g29549 ( n4897 , n6355 , n15286 );
    or g29550 ( n19552 , n13620 , n27761 );
    or g29551 ( n36772 , n13948 , n25078 );
    and g29552 ( n22370 , n15536 , n16781 );
    nor g29553 ( n18118 , n40369 , n24783 );
    not g29554 ( n974 , n37239 );
    or g29555 ( n27168 , n35450 , n28561 );
    and g29556 ( n41732 , n38664 , n38375 );
    or g29557 ( n12753 , n32762 , n13647 );
    and g29558 ( n7623 , n24464 , n38540 );
    not g29559 ( n6602 , n19227 );
    or g29560 ( n22141 , n6094 , n23213 );
    nor g29561 ( n31437 , n605 , n41341 );
    not g29562 ( n11346 , n18862 );
    or g29563 ( n15129 , n2992 , n29930 );
    or g29564 ( n9368 , n12566 , n32671 );
    and g29565 ( n6309 , n5414 , n18127 );
    or g29566 ( n30303 , n29826 , n31176 );
    and g29567 ( n33873 , n22963 , n17639 );
    or g29568 ( n537 , n38653 , n17280 );
    and g29569 ( n23348 , n24406 , n795 );
    or g29570 ( n5603 , n5859 , n28207 );
    or g29571 ( n32336 , n21068 , n29776 );
    not g29572 ( n29658 , n21816 );
    and g29573 ( n14223 , n34366 , n41043 );
    or g29574 ( n20996 , n12452 , n439 );
    not g29575 ( n1913 , n38642 );
    and g29576 ( n22751 , n35561 , n33816 );
    or g29577 ( n30501 , n34204 , n34960 );
    not g29578 ( n24441 , n25630 );
    and g29579 ( n18865 , n18813 , n15420 );
    or g29580 ( n20012 , n25725 , n16281 );
    or g29581 ( n7330 , n21558 , n9489 );
    xnor g29582 ( n29611 , n14502 , n12607 );
    nor g29583 ( n33252 , n15823 , n38772 );
    not g29584 ( n6684 , n15541 );
    xnor g29585 ( n12537 , n2338 , n38507 );
    not g29586 ( n27745 , n40912 );
    not g29587 ( n28801 , n9279 );
    xnor g29588 ( n32552 , n40150 , n6579 );
    and g29589 ( n9799 , n37426 , n23100 );
    not g29590 ( n29049 , n8566 );
    and g29591 ( n28345 , n12905 , n40089 );
    or g29592 ( n16976 , n12650 , n19848 );
    and g29593 ( n41676 , n34518 , n31876 );
    or g29594 ( n27870 , n29104 , n23520 );
    and g29595 ( n27490 , n20490 , n22736 );
    or g29596 ( n20119 , n4762 , n7378 );
    and g29597 ( n4088 , n35546 , n34814 );
    or g29598 ( n32205 , n27232 , n8418 );
    or g29599 ( n33358 , n24289 , n12768 );
    and g29600 ( n42682 , n6767 , n6675 );
    nor g29601 ( n20613 , n7236 , n17922 );
    or g29602 ( n31233 , n28932 , n11475 );
    and g29603 ( n25448 , n29639 , n18849 );
    and g29604 ( n19955 , n12693 , n39667 );
    nor g29605 ( n32848 , n3437 , n27260 );
    or g29606 ( n11045 , n37968 , n26348 );
    or g29607 ( n9672 , n26889 , n10503 );
    and g29608 ( n23067 , n14080 , n33565 );
    or g29609 ( n35125 , n3700 , n34715 );
    nor g29610 ( n10534 , n5961 , n22432 );
    not g29611 ( n38777 , n16994 );
    or g29612 ( n4205 , n15096 , n29808 );
    and g29613 ( n27109 , n6508 , n30503 );
    xnor g29614 ( n40771 , n24159 , n39316 );
    and g29615 ( n22628 , n13602 , n41912 );
    nor g29616 ( n38560 , n18866 , n7079 );
    or g29617 ( n30947 , n3954 , n23332 );
    or g29618 ( n4684 , n10625 , n25116 );
    and g29619 ( n36022 , n23072 , n42480 );
    or g29620 ( n32331 , n11818 , n7075 );
    or g29621 ( n11831 , n1190 , n21697 );
    xnor g29622 ( n42191 , n13290 , n21358 );
    or g29623 ( n12626 , n15185 , n20880 );
    nor g29624 ( n42437 , n2223 , n23300 );
    not g29625 ( n27595 , n14240 );
    or g29626 ( n17282 , n32087 , n10878 );
    or g29627 ( n4626 , n27712 , n4735 );
    or g29628 ( n37298 , n34292 , n40543 );
    or g29629 ( n31152 , n13837 , n38013 );
    not g29630 ( n27915 , n35705 );
    or g29631 ( n42051 , n5899 , n37341 );
    or g29632 ( n36879 , n25033 , n36485 );
    and g29633 ( n39350 , n38760 , n39272 );
    xnor g29634 ( n8897 , n38836 , n42125 );
    nor g29635 ( n29252 , n10598 , n31681 );
    and g29636 ( n39634 , n16380 , n19458 );
    xnor g29637 ( n21436 , n29120 , n24539 );
    or g29638 ( n15676 , n10714 , n34959 );
    not g29639 ( n39924 , n31184 );
    or g29640 ( n12602 , n29815 , n18337 );
    not g29641 ( n40785 , n38555 );
    or g29642 ( n24777 , n5341 , n12665 );
    xnor g29643 ( n14390 , n35347 , n41172 );
    and g29644 ( n31553 , n40399 , n38410 );
    not g29645 ( n16826 , n38819 );
    xnor g29646 ( n3301 , n25942 , n27591 );
    or g29647 ( n12217 , n9673 , n31465 );
    not g29648 ( n8952 , n32078 );
    not g29649 ( n26344 , n15354 );
    and g29650 ( n14800 , n9846 , n42412 );
    and g29651 ( n11092 , n28842 , n35183 );
    xnor g29652 ( n10875 , n31275 , n6763 );
    not g29653 ( n11460 , n6054 );
    or g29654 ( n19458 , n23907 , n1416 );
    or g29655 ( n7057 , n3571 , n3851 );
    not g29656 ( n19014 , n42844 );
    or g29657 ( n18147 , n36793 , n19007 );
    or g29658 ( n39046 , n36257 , n16683 );
    not g29659 ( n39609 , n28259 );
    and g29660 ( n14875 , n8493 , n15065 );
    or g29661 ( n1204 , n5274 , n21282 );
    not g29662 ( n37961 , n26655 );
    or g29663 ( n33384 , n7127 , n37238 );
    nor g29664 ( n23359 , n12954 , n34256 );
    nor g29665 ( n15349 , n16604 , n29793 );
    not g29666 ( n18236 , n29047 );
    nor g29667 ( n24909 , n21786 , n28702 );
    not g29668 ( n15822 , n38112 );
    xnor g29669 ( n12682 , n36998 , n38401 );
    or g29670 ( n31934 , n40521 , n29311 );
    and g29671 ( n22692 , n3655 , n29453 );
    xnor g29672 ( n24912 , n41218 , n37419 );
    xnor g29673 ( n40454 , n28648 , n28430 );
    or g29674 ( n37782 , n18763 , n10636 );
    not g29675 ( n15807 , n1166 );
    or g29676 ( n24362 , n35899 , n12768 );
    not g29677 ( n16980 , n36224 );
    xnor g29678 ( n39611 , n24734 , n26048 );
    xnor g29679 ( n9126 , n16442 , n38301 );
    or g29680 ( n21511 , n34262 , n7276 );
    not g29681 ( n14363 , n40125 );
    xnor g29682 ( n5533 , n41652 , n42400 );
    and g29683 ( n11186 , n33591 , n41189 );
    or g29684 ( n37187 , n1867 , n26737 );
    not g29685 ( n7999 , n32526 );
    and g29686 ( n30853 , n16731 , n3371 );
    and g29687 ( n10447 , n25166 , n42590 );
    xnor g29688 ( n15088 , n11657 , n10715 );
    xnor g29689 ( n35939 , n30549 , n25133 );
    or g29690 ( n20248 , n1404 , n32782 );
    not g29691 ( n30045 , n41165 );
    not g29692 ( n15771 , n36769 );
    or g29693 ( n42323 , n19469 , n36631 );
    or g29694 ( n16933 , n27092 , n21650 );
    xnor g29695 ( n19263 , n19463 , n7768 );
    or g29696 ( n5669 , n20612 , n4592 );
    or g29697 ( n19940 , n33142 , n18086 );
    and g29698 ( n21527 , n3145 , n25747 );
    or g29699 ( n1886 , n10406 , n18102 );
    nor g29700 ( n12963 , n5319 , n37691 );
    not g29701 ( n19494 , n637 );
    or g29702 ( n24385 , n32245 , n23388 );
    and g29703 ( n40484 , n20890 , n31993 );
    or g29704 ( n30749 , n20394 , n31361 );
    or g29705 ( n41786 , n4492 , n27306 );
    and g29706 ( n34993 , n34936 , n10185 );
    or g29707 ( n23317 , n22437 , n34007 );
    or g29708 ( n41731 , n11628 , n14553 );
    xnor g29709 ( n37841 , n2130 , n32214 );
    xnor g29710 ( n17636 , n36568 , n33981 );
    not g29711 ( n17914 , n18017 );
    or g29712 ( n37861 , n10967 , n14000 );
    xnor g29713 ( n33043 , n34248 , n1971 );
    xnor g29714 ( n3500 , n26579 , n5377 );
    xnor g29715 ( n9226 , n5457 , n32873 );
    nor g29716 ( n33847 , n29681 , n39846 );
    not g29717 ( n10978 , n3190 );
    or g29718 ( n18150 , n3982 , n28933 );
    and g29719 ( n25522 , n14359 , n41324 );
    xnor g29720 ( n32055 , n24677 , n14471 );
    or g29721 ( n17879 , n1110 , n9521 );
    nor g29722 ( n683 , n14457 , n38056 );
    or g29723 ( n8692 , n38761 , n11052 );
    xnor g29724 ( n14477 , n29452 , n6393 );
    or g29725 ( n42727 , n20932 , n37218 );
    or g29726 ( n30486 , n37062 , n13101 );
    xnor g29727 ( n10207 , n921 , n19338 );
    or g29728 ( n24244 , n11053 , n30750 );
    and g29729 ( n21060 , n15928 , n20906 );
    xnor g29730 ( n10173 , n7425 , n9459 );
    or g29731 ( n34342 , n32770 , n30614 );
    not g29732 ( n42431 , n21455 );
    and g29733 ( n8587 , n9927 , n31929 );
    xnor g29734 ( n29721 , n20204 , n30908 );
    or g29735 ( n20886 , n18927 , n11960 );
    xnor g29736 ( n16547 , n4511 , n26769 );
    nor g29737 ( n6788 , n32542 , n37425 );
    or g29738 ( n2490 , n40881 , n24124 );
    and g29739 ( n27193 , n11185 , n35640 );
    and g29740 ( n37027 , n12213 , n22650 );
    or g29741 ( n22001 , n18005 , n21919 );
    nor g29742 ( n19131 , n33745 , n38067 );
    or g29743 ( n6674 , n11239 , n3560 );
    xnor g29744 ( n17664 , n1907 , n18256 );
    or g29745 ( n18896 , n32920 , n936 );
    or g29746 ( n4891 , n16205 , n7468 );
    or g29747 ( n11545 , n32100 , n7573 );
    xnor g29748 ( n28658 , n4334 , n12610 );
    not g29749 ( n29513 , n15399 );
    and g29750 ( n42105 , n34295 , n40290 );
    nor g29751 ( n22023 , n16391 , n10387 );
    nor g29752 ( n5849 , n247 , n35482 );
    or g29753 ( n3452 , n1173 , n21893 );
    nor g29754 ( n42466 , n22577 , n5364 );
    or g29755 ( n36881 , n35274 , n14166 );
    or g29756 ( n6289 , n22866 , n2507 );
    or g29757 ( n8670 , n18314 , n20452 );
    not g29758 ( n27900 , n31626 );
    and g29759 ( n11955 , n6164 , n27521 );
    nor g29760 ( n32458 , n36993 , n10582 );
    and g29761 ( n34256 , n29733 , n5433 );
    nor g29762 ( n31090 , n31310 , n19951 );
    nor g29763 ( n7872 , n4205 , n300 );
    xnor g29764 ( n30838 , n6 , n22927 );
    or g29765 ( n30047 , n29443 , n12849 );
    xnor g29766 ( n30855 , n40191 , n41820 );
    not g29767 ( n30103 , n40299 );
    not g29768 ( n32110 , n744 );
    not g29769 ( n1829 , n8132 );
    not g29770 ( n39827 , n31 );
    xnor g29771 ( n5182 , n105 , n1318 );
    and g29772 ( n36490 , n6888 , n23317 );
    or g29773 ( n4136 , n27081 , n35401 );
    or g29774 ( n5682 , n33694 , n1006 );
    and g29775 ( n39393 , n38415 , n7505 );
    or g29776 ( n1543 , n22273 , n31469 );
    or g29777 ( n34598 , n19666 , n23749 );
    and g29778 ( n17640 , n27927 , n24274 );
    or g29779 ( n13079 , n15095 , n28039 );
    or g29780 ( n15235 , n1980 , n30974 );
    or g29781 ( n24633 , n32410 , n42464 );
    not g29782 ( n18679 , n12467 );
    or g29783 ( n17520 , n19762 , n33813 );
    xnor g29784 ( n5793 , n33444 , n11491 );
    and g29785 ( n41689 , n32260 , n8690 );
    and g29786 ( n7418 , n20143 , n6471 );
    or g29787 ( n33412 , n32329 , n21856 );
    or g29788 ( n12703 , n6904 , n22767 );
    or g29789 ( n31162 , n31702 , n27950 );
    or g29790 ( n35254 , n29677 , n37877 );
    and g29791 ( n29255 , n22798 , n21617 );
    or g29792 ( n33270 , n21955 , n12910 );
    or g29793 ( n41835 , n15900 , n6484 );
    nor g29794 ( n12017 , n41302 , n33735 );
    xnor g29795 ( n5890 , n19592 , n21563 );
    xnor g29796 ( n10732 , n6703 , n2199 );
    nor g29797 ( n5742 , n41112 , n9065 );
    xnor g29798 ( n30861 , n12146 , n28653 );
    nor g29799 ( n40761 , n28658 , n5388 );
    and g29800 ( n33623 , n18255 , n40609 );
    nor g29801 ( n18590 , n25402 , n24106 );
    and g29802 ( n27561 , n41218 , n27595 );
    and g29803 ( n14704 , n16385 , n6803 );
    not g29804 ( n35898 , n32588 );
    and g29805 ( n24033 , n13697 , n31163 );
    not g29806 ( n25775 , n10587 );
    nor g29807 ( n26567 , n38173 , n10755 );
    nor g29808 ( n15997 , n13674 , n23495 );
    or g29809 ( n13090 , n39266 , n13509 );
    or g29810 ( n41550 , n37685 , n21364 );
    or g29811 ( n126 , n18798 , n40195 );
    not g29812 ( n2086 , n29349 );
    or g29813 ( n37160 , n16212 , n16159 );
    or g29814 ( n23129 , n13453 , n15780 );
    and g29815 ( n5299 , n16431 , n14017 );
    not g29816 ( n27407 , n10308 );
    not g29817 ( n33135 , n30220 );
    nor g29818 ( n32918 , n26916 , n16538 );
    xnor g29819 ( n31161 , n21457 , n21791 );
    not g29820 ( n2105 , n23032 );
    xnor g29821 ( n8868 , n17198 , n13944 );
    nor g29822 ( n29773 , n33434 , n40868 );
    or g29823 ( n40975 , n1186 , n23821 );
    and g29824 ( n25741 , n8336 , n28496 );
    xnor g29825 ( n31136 , n29670 , n29676 );
    not g29826 ( n35468 , n1134 );
    or g29827 ( n11206 , n23728 , n17911 );
    or g29828 ( n6354 , n41591 , n31531 );
    nor g29829 ( n32425 , n14707 , n748 );
    or g29830 ( n42606 , n16381 , n5342 );
    not g29831 ( n15101 , n10297 );
    or g29832 ( n39969 , n5978 , n24822 );
    xnor g29833 ( n31291 , n1464 , n41332 );
    xnor g29834 ( n9421 , n25619 , n33604 );
    nor g29835 ( n34695 , n40472 , n24049 );
    or g29836 ( n24908 , n32605 , n4090 );
    and g29837 ( n21904 , n27263 , n36955 );
    or g29838 ( n28660 , n22342 , n39789 );
    nor g29839 ( n25282 , n32701 , n2180 );
    not g29840 ( n30030 , n37770 );
    not g29841 ( n24549 , n25607 );
    and g29842 ( n19809 , n11540 , n14915 );
    or g29843 ( n24182 , n17067 , n37371 );
    not g29844 ( n28894 , n39587 );
    and g29845 ( n32358 , n8187 , n33047 );
    xnor g29846 ( n14718 , n11784 , n10790 );
    or g29847 ( n17350 , n39391 , n39508 );
    xnor g29848 ( n41338 , n31226 , n42014 );
    and g29849 ( n20992 , n18530 , n14300 );
    or g29850 ( n34374 , n33528 , n22289 );
    xnor g29851 ( n6 , n25118 , n13635 );
    or g29852 ( n5172 , n31918 , n38690 );
    nor g29853 ( n14788 , n4922 , n16234 );
    or g29854 ( n22929 , n30313 , n32892 );
    nor g29855 ( n34730 , n3074 , n1302 );
    nor g29856 ( n40550 , n10414 , n32296 );
    and g29857 ( n21217 , n17543 , n22913 );
    not g29858 ( n28317 , n2418 );
    or g29859 ( n14333 , n789 , n31986 );
    not g29860 ( n42392 , n38341 );
    or g29861 ( n4175 , n34547 , n31964 );
    or g29862 ( n42876 , n6020 , n42220 );
    nor g29863 ( n3796 , n16598 , n34228 );
    or g29864 ( n22155 , n31482 , n9508 );
    nor g29865 ( n36527 , n20952 , n38021 );
    nor g29866 ( n18133 , n4451 , n34490 );
    nor g29867 ( n26963 , n15530 , n4263 );
    xnor g29868 ( n6329 , n41013 , n24326 );
    and g29869 ( n20312 , n18887 , n25054 );
    and g29870 ( n5454 , n33509 , n1135 );
    xnor g29871 ( n39247 , n11436 , n22919 );
    nor g29872 ( n40547 , n17744 , n12582 );
    or g29873 ( n16242 , n29118 , n41649 );
    and g29874 ( n15375 , n6640 , n19291 );
    and g29875 ( n14274 , n2635 , n6704 );
    and g29876 ( n16808 , n2532 , n13903 );
    or g29877 ( n42262 , n20288 , n29965 );
    not g29878 ( n17561 , n2919 );
    or g29879 ( n40199 , n28643 , n6353 );
    or g29880 ( n27467 , n16509 , n22355 );
    xnor g29881 ( n19566 , n34947 , n39074 );
    and g29882 ( n27910 , n20236 , n14113 );
    not g29883 ( n22398 , n32148 );
    and g29884 ( n40035 , n15316 , n533 );
    xnor g29885 ( n10984 , n37026 , n82 );
    not g29886 ( n27612 , n39289 );
    or g29887 ( n23765 , n25677 , n42380 );
    and g29888 ( n6039 , n26074 , n2928 );
    or g29889 ( n890 , n22427 , n1288 );
    not g29890 ( n877 , n8504 );
    and g29891 ( n2694 , n28835 , n21040 );
    and g29892 ( n25567 , n12107 , n23932 );
    and g29893 ( n15759 , n21311 , n39800 );
    or g29894 ( n4005 , n8551 , n26577 );
    and g29895 ( n5198 , n24703 , n25431 );
    or g29896 ( n38091 , n2193 , n4014 );
    not g29897 ( n11549 , n11423 );
    or g29898 ( n42619 , n34105 , n25200 );
    xnor g29899 ( n25610 , n21476 , n25038 );
    or g29900 ( n23029 , n35023 , n14434 );
    or g29901 ( n1271 , n26651 , n34793 );
    or g29902 ( n30629 , n16586 , n600 );
    not g29903 ( n25025 , n31222 );
    or g29904 ( n7377 , n12538 , n14012 );
    or g29905 ( n33309 , n17946 , n1036 );
    or g29906 ( n30758 , n29164 , n6156 );
    not g29907 ( n11784 , n25738 );
    or g29908 ( n7217 , n1267 , n10465 );
    nor g29909 ( n25926 , n35606 , n6114 );
    and g29910 ( n42420 , n16431 , n40680 );
    and g29911 ( n7474 , n39473 , n1845 );
    or g29912 ( n38280 , n5991 , n28027 );
    not g29913 ( n34762 , n36811 );
    nor g29914 ( n40489 , n8089 , n6206 );
    not g29915 ( n3610 , n21875 );
    not g29916 ( n16489 , n3209 );
    and g29917 ( n3042 , n25655 , n13522 );
    or g29918 ( n18347 , n38098 , n6359 );
    and g29919 ( n17539 , n34727 , n13224 );
    xnor g29920 ( n40155 , n11434 , n10141 );
    or g29921 ( n27094 , n10460 , n26841 );
    or g29922 ( n6816 , n2893 , n7896 );
    xnor g29923 ( n33642 , n35322 , n36659 );
    xnor g29924 ( n7198 , n27968 , n3677 );
    or g29925 ( n23277 , n31535 , n17321 );
    not g29926 ( n20252 , n1086 );
    nor g29927 ( n12730 , n22387 , n41088 );
    nor g29928 ( n29199 , n31126 , n7680 );
    or g29929 ( n18110 , n12906 , n22756 );
    not g29930 ( n40405 , n25111 );
    or g29931 ( n42175 , n6170 , n12121 );
    xnor g29932 ( n42833 , n32160 , n23013 );
    nor g29933 ( n15310 , n26256 , n36089 );
    nor g29934 ( n25466 , n7987 , n31530 );
    or g29935 ( n40503 , n32683 , n33742 );
    or g29936 ( n8743 , n22955 , n12867 );
    or g29937 ( n16114 , n12947 , n19565 );
    or g29938 ( n7565 , n254 , n14622 );
    and g29939 ( n42867 , n5296 , n10734 );
    or g29940 ( n14964 , n27518 , n42544 );
    or g29941 ( n21238 , n36142 , n40484 );
    not g29942 ( n10579 , n3060 );
    nor g29943 ( n14603 , n26394 , n30820 );
    or g29944 ( n30120 , n36117 , n30447 );
    nor g29945 ( n40055 , n10104 , n35353 );
    nor g29946 ( n6255 , n7598 , n11407 );
    nor g29947 ( n6380 , n39827 , n30150 );
    or g29948 ( n32760 , n12628 , n12044 );
    or g29949 ( n35552 , n5551 , n40178 );
    and g29950 ( n39550 , n4078 , n1523 );
    not g29951 ( n38283 , n7760 );
    or g29952 ( n22453 , n11774 , n34267 );
    and g29953 ( n29809 , n20533 , n25645 );
    and g29954 ( n18608 , n17430 , n270 );
    and g29955 ( n11651 , n33641 , n11665 );
    not g29956 ( n27542 , n31571 );
    xnor g29957 ( n18972 , n2632 , n1640 );
    or g29958 ( n27196 , n4679 , n12484 );
    or g29959 ( n32995 , n11553 , n21721 );
    or g29960 ( n32337 , n1954 , n41854 );
    xnor g29961 ( n2751 , n36998 , n17021 );
    or g29962 ( n29725 , n5812 , n34796 );
    not g29963 ( n5947 , n39364 );
    xnor g29964 ( n37595 , n9030 , n7335 );
    or g29965 ( n10124 , n33982 , n36483 );
    or g29966 ( n35447 , n10496 , n18170 );
    nor g29967 ( n33461 , n5302 , n39988 );
    or g29968 ( n20906 , n34466 , n31213 );
    xnor g29969 ( n17118 , n31018 , n31880 );
    and g29970 ( n33704 , n26208 , n1855 );
    or g29971 ( n23603 , n24495 , n6394 );
    or g29972 ( n41796 , n15125 , n23444 );
    or g29973 ( n16444 , n40109 , n35739 );
    and g29974 ( n15245 , n11131 , n4973 );
    and g29975 ( n33588 , n19822 , n37424 );
    xnor g29976 ( n33435 , n2292 , n24614 );
    not g29977 ( n18345 , n25972 );
    or g29978 ( n3628 , n19416 , n9896 );
    and g29979 ( n23559 , n139 , n8448 );
    or g29980 ( n8909 , n29942 , n42792 );
    and g29981 ( n10106 , n8633 , n188 );
    not g29982 ( n1921 , n7391 );
    or g29983 ( n40633 , n37664 , n7283 );
    or g29984 ( n13896 , n25174 , n14040 );
    xnor g29985 ( n6403 , n12977 , n39701 );
    xnor g29986 ( n18272 , n38899 , n20035 );
    not g29987 ( n26196 , n5305 );
    not g29988 ( n26089 , n172 );
    not g29989 ( n28608 , n30297 );
    or g29990 ( n37329 , n2052 , n31156 );
    nor g29991 ( n30417 , n27961 , n2780 );
    or g29992 ( n38584 , n25142 , n30733 );
    not g29993 ( n30140 , n4782 );
    xnor g29994 ( n38571 , n16418 , n38713 );
    or g29995 ( n17745 , n3720 , n8736 );
    or g29996 ( n24838 , n34810 , n41326 );
    not g29997 ( n20323 , n26613 );
    not g29998 ( n10226 , n28956 );
    and g29999 ( n41347 , n1471 , n2406 );
    nor g30000 ( n22968 , n37708 , n42036 );
    and g30001 ( n25520 , n2961 , n15568 );
    or g30002 ( n30642 , n23082 , n29434 );
    or g30003 ( n359 , n11135 , n17104 );
    or g30004 ( n34307 , n35559 , n9862 );
    nor g30005 ( n9576 , n32802 , n17110 );
    or g30006 ( n34593 , n12658 , n32707 );
    or g30007 ( n31985 , n9534 , n17475 );
    or g30008 ( n8961 , n12964 , n3657 );
    or g30009 ( n38779 , n16466 , n9938 );
    not g30010 ( n17264 , n12514 );
    or g30011 ( n42849 , n1444 , n29637 );
    or g30012 ( n10287 , n20831 , n39839 );
    or g30013 ( n18355 , n9474 , n34027 );
    and g30014 ( n14949 , n28829 , n4622 );
    and g30015 ( n13733 , n15279 , n13800 );
    or g30016 ( n33943 , n31452 , n35416 );
    or g30017 ( n35241 , n39571 , n11092 );
    not g30018 ( n6732 , n3907 );
    xnor g30019 ( n2952 , n33917 , n25238 );
    and g30020 ( n25719 , n12145 , n5937 );
    and g30021 ( n8989 , n23019 , n35756 );
    or g30022 ( n41091 , n23026 , n36573 );
    or g30023 ( n18255 , n42408 , n33926 );
    and g30024 ( n19359 , n31424 , n30580 );
    and g30025 ( n28554 , n32753 , n20905 );
    xnor g30026 ( n35709 , n11383 , n13310 );
    xnor g30027 ( n39384 , n26579 , n30152 );
    or g30028 ( n39525 , n34869 , n40561 );
    or g30029 ( n9909 , n42220 , n15210 );
    not g30030 ( n9652 , n32175 );
    and g30031 ( n19782 , n15050 , n40474 );
    or g30032 ( n15825 , n27831 , n36344 );
    not g30033 ( n6054 , n26032 );
    nor g30034 ( n17491 , n35771 , n14269 );
    or g30035 ( n28478 , n32070 , n26797 );
    or g30036 ( n15749 , n34462 , n2785 );
    xnor g30037 ( n978 , n31293 , n1434 );
    or g30038 ( n3219 , n5458 , n21299 );
    nor g30039 ( n18116 , n20759 , n4483 );
    or g30040 ( n18754 , n19486 , n16058 );
    and g30041 ( n37843 , n34540 , n23992 );
    and g30042 ( n19387 , n32937 , n16626 );
    xnor g30043 ( n40889 , n15495 , n15607 );
    nor g30044 ( n18607 , n35030 , n28659 );
    and g30045 ( n19766 , n24420 , n21889 );
    or g30046 ( n1124 , n37706 , n23563 );
    xnor g30047 ( n38714 , n105 , n6613 );
    xnor g30048 ( n38905 , n20966 , n41190 );
    or g30049 ( n39035 , n2909 , n34993 );
    nor g30050 ( n34807 , n20948 , n29654 );
    and g30051 ( n21546 , n25452 , n29908 );
    not g30052 ( n22675 , n23629 );
    or g30053 ( n21206 , n26625 , n21268 );
    or g30054 ( n18640 , n18607 , n25178 );
    and g30055 ( n39697 , n7320 , n38823 );
    nor g30056 ( n39898 , n5398 , n36962 );
    nor g30057 ( n23198 , n26483 , n22269 );
    nor g30058 ( n18587 , n5170 , n13313 );
    not g30059 ( n11530 , n22525 );
    and g30060 ( n21977 , n13432 , n26450 );
    or g30061 ( n37537 , n35320 , n13514 );
    or g30062 ( n3527 , n33873 , n29388 );
    or g30063 ( n849 , n15905 , n23834 );
    or g30064 ( n31926 , n37980 , n19825 );
    and g30065 ( n26488 , n12353 , n34178 );
    or g30066 ( n21659 , n12722 , n30968 );
    nor g30067 ( n16083 , n29103 , n33400 );
    not g30068 ( n15281 , n16582 );
    or g30069 ( n3176 , n7443 , n36902 );
    or g30070 ( n39219 , n7196 , n19359 );
    nor g30071 ( n1967 , n33981 , n21283 );
    not g30072 ( n15403 , n1879 );
    or g30073 ( n22873 , n28495 , n13282 );
    and g30074 ( n11476 , n14310 , n20397 );
    nor g30075 ( n29994 , n35112 , n31356 );
    not g30076 ( n26339 , n35831 );
    xnor g30077 ( n8484 , n3068 , n34908 );
    not g30078 ( n28638 , n38533 );
    xnor g30079 ( n41343 , n6760 , n17149 );
    not g30080 ( n33401 , n686 );
    or g30081 ( n4122 , n42442 , n826 );
    and g30082 ( n18196 , n26691 , n25618 );
    nor g30083 ( n40056 , n32949 , n34826 );
    or g30084 ( n15794 , n7142 , n16383 );
    or g30085 ( n23368 , n2883 , n21772 );
    nor g30086 ( n36105 , n7001 , n6037 );
    or g30087 ( n19127 , n23982 , n33320 );
    xnor g30088 ( n41814 , n36009 , n9000 );
    xnor g30089 ( n35617 , n25231 , n20725 );
    and g30090 ( n80 , n26073 , n41607 );
    or g30091 ( n17424 , n42637 , n23211 );
    nor g30092 ( n30700 , n35055 , n4932 );
    nor g30093 ( n38910 , n33751 , n42784 );
    and g30094 ( n38942 , n33663 , n34425 );
    or g30095 ( n22930 , n33556 , n3368 );
    or g30096 ( n28739 , n10789 , n9753 );
    nor g30097 ( n32628 , n10152 , n1581 );
    nor g30098 ( n741 , n23745 , n42342 );
    not g30099 ( n26168 , n1681 );
    or g30100 ( n13652 , n18866 , n7307 );
    or g30101 ( n9659 , n15552 , n7831 );
    or g30102 ( n22479 , n2296 , n2363 );
    and g30103 ( n40473 , n18079 , n2771 );
    or g30104 ( n14430 , n25526 , n33557 );
    or g30105 ( n13792 , n15780 , n36101 );
    or g30106 ( n25585 , n13530 , n30239 );
    xnor g30107 ( n6176 , n27900 , n27827 );
    or g30108 ( n25208 , n4619 , n16669 );
    or g30109 ( n42700 , n37139 , n31606 );
    xnor g30110 ( n736 , n12146 , n20215 );
    or g30111 ( n41838 , n15370 , n13074 );
    or g30112 ( n12451 , n30053 , n1757 );
    not g30113 ( n27765 , n35869 );
    or g30114 ( n28176 , n11800 , n1536 );
    not g30115 ( n23369 , n1287 );
    nor g30116 ( n25576 , n39266 , n7775 );
    xnor g30117 ( n29438 , n28377 , n33260 );
    or g30118 ( n10627 , n7482 , n20446 );
    or g30119 ( n38225 , n35308 , n15658 );
    not g30120 ( n4424 , n21183 );
    or g30121 ( n24343 , n27631 , n9717 );
    not g30122 ( n24016 , n39854 );
    not g30123 ( n15685 , n40013 );
    or g30124 ( n23113 , n42864 , n14659 );
    and g30125 ( n21364 , n28834 , n14729 );
    or g30126 ( n37735 , n13687 , n36573 );
    or g30127 ( n21750 , n22197 , n15246 );
    not g30128 ( n1338 , n19629 );
    not g30129 ( n23080 , n4109 );
    nor g30130 ( n35941 , n23546 , n3774 );
    not g30131 ( n15675 , n11398 );
    nor g30132 ( n14248 , n812 , n24561 );
    nor g30133 ( n20638 , n40275 , n18043 );
    not g30134 ( n112 , n28577 );
    and g30135 ( n18486 , n34399 , n8095 );
    not g30136 ( n32341 , n23326 );
    or g30137 ( n30059 , n3767 , n24395 );
    not g30138 ( n42567 , n29457 );
    or g30139 ( n24451 , n21170 , n30772 );
    or g30140 ( n14933 , n39954 , n15743 );
    xnor g30141 ( n38462 , n31989 , n7307 );
    and g30142 ( n2593 , n33340 , n7380 );
    and g30143 ( n18758 , n25606 , n10407 );
    or g30144 ( n31729 , n20075 , n1911 );
    or g30145 ( n5492 , n9673 , n37677 );
    not g30146 ( n19574 , n12260 );
    not g30147 ( n41114 , n18566 );
    and g30148 ( n18499 , n29034 , n2687 );
    or g30149 ( n30913 , n23971 , n26516 );
    or g30150 ( n6995 , n10979 , n2657 );
    and g30151 ( n19332 , n25205 , n9120 );
    nor g30152 ( n10717 , n18749 , n1252 );
    not g30153 ( n30237 , n4873 );
    not g30154 ( n35158 , n16075 );
    or g30155 ( n20212 , n27092 , n22924 );
    or g30156 ( n4303 , n26632 , n7616 );
    and g30157 ( n24168 , n27423 , n32626 );
    or g30158 ( n20637 , n6452 , n18332 );
    and g30159 ( n21817 , n11266 , n36281 );
    not g30160 ( n25673 , n11879 );
    or g30161 ( n10795 , n24248 , n29229 );
    and g30162 ( n4954 , n10061 , n13542 );
    and g30163 ( n23270 , n41013 , n42064 );
    or g30164 ( n21070 , n9893 , n16803 );
    xnor g30165 ( n10324 , n14302 , n10661 );
    or g30166 ( n590 , n4130 , n1053 );
    not g30167 ( n22310 , n38271 );
    or g30168 ( n23642 , n41614 , n13025 );
    nor g30169 ( n9772 , n22915 , n8014 );
    nor g30170 ( n36507 , n31256 , n14139 );
    or g30171 ( n40328 , n15771 , n36463 );
    or g30172 ( n41707 , n17919 , n39481 );
    or g30173 ( n11501 , n21564 , n1970 );
    or g30174 ( n17683 , n31580 , n36774 );
    or g30175 ( n7757 , n41532 , n22568 );
    and g30176 ( n18458 , n20109 , n9853 );
    xnor g30177 ( n33808 , n35727 , n364 );
    and g30178 ( n41216 , n12082 , n24995 );
    not g30179 ( n20554 , n12652 );
    not g30180 ( n23082 , n17918 );
    or g30181 ( n14961 , n23880 , n17218 );
    nor g30182 ( n19225 , n30743 , n28624 );
    or g30183 ( n1019 , n13732 , n42447 );
    not g30184 ( n13265 , n13345 );
    and g30185 ( n13744 , n22302 , n24796 );
    or g30186 ( n36469 , n33530 , n18612 );
    and g30187 ( n12028 , n33716 , n37554 );
    or g30188 ( n37004 , n20749 , n32516 );
    not g30189 ( n31372 , n31461 );
    and g30190 ( n39153 , n40717 , n18776 );
    or g30191 ( n25248 , n40485 , n32232 );
    and g30192 ( n32353 , n19001 , n24126 );
    xnor g30193 ( n12015 , n20016 , n10732 );
    or g30194 ( n40657 , n36349 , n37640 );
    and g30195 ( n414 , n39157 , n15170 );
    xnor g30196 ( n14759 , n24159 , n31218 );
    xnor g30197 ( n17789 , n31099 , n6092 );
    and g30198 ( n6288 , n30158 , n35634 );
    and g30199 ( n30767 , n13915 , n37613 );
    xnor g30200 ( n24027 , n7118 , n34565 );
    or g30201 ( n10478 , n1702 , n36717 );
    or g30202 ( n29342 , n17538 , n26369 );
    and g30203 ( n40014 , n39864 , n32419 );
    nor g30204 ( n38014 , n39556 , n16388 );
    or g30205 ( n40828 , n14244 , n24104 );
    nor g30206 ( n4306 , n34926 , n14011 );
    xnor g30207 ( n9228 , n20851 , n8530 );
    xnor g30208 ( n33202 , n19700 , n8864 );
    not g30209 ( n13282 , n30845 );
    and g30210 ( n21440 , n41618 , n38567 );
    xnor g30211 ( n22027 , n34562 , n40154 );
    not g30212 ( n25030 , n23018 );
    or g30213 ( n4520 , n7427 , n30668 );
    or g30214 ( n40595 , n6836 , n41891 );
    or g30215 ( n7610 , n4373 , n31580 );
    xnor g30216 ( n29727 , n5041 , n22464 );
    not g30217 ( n8694 , n35238 );
    and g30218 ( n5294 , n22725 , n42403 );
    or g30219 ( n24292 , n14622 , n41523 );
    xnor g30220 ( n29709 , n41129 , n14707 );
    or g30221 ( n15933 , n24482 , n37202 );
    xnor g30222 ( n588 , n12524 , n7732 );
    not g30223 ( n23942 , n7975 );
    not g30224 ( n25781 , n29715 );
    or g30225 ( n12999 , n25440 , n28329 );
    or g30226 ( n24794 , n37615 , n19470 );
    not g30227 ( n37167 , n5448 );
    or g30228 ( n25538 , n39661 , n41532 );
    or g30229 ( n3579 , n38228 , n21562 );
    nor g30230 ( n21528 , n36117 , n15540 );
    nor g30231 ( n18961 , n25930 , n10412 );
    not g30232 ( n18667 , n32990 );
    not g30233 ( n4173 , n31138 );
    not g30234 ( n29896 , n18438 );
    or g30235 ( n22255 , n12991 , n2499 );
    or g30236 ( n5397 , n34565 , n4680 );
    or g30237 ( n31058 , n33733 , n4806 );
    or g30238 ( n16035 , n10423 , n19487 );
    xnor g30239 ( n719 , n41053 , n9986 );
    not g30240 ( n20617 , n38323 );
    and g30241 ( n22735 , n18184 , n16770 );
    and g30242 ( n5091 , n39607 , n17806 );
    and g30243 ( n30653 , n24181 , n31659 );
    xnor g30244 ( n33058 , n34562 , n5199 );
    xnor g30245 ( n33629 , n11884 , n23212 );
    or g30246 ( n14439 , n30552 , n13044 );
    or g30247 ( n39605 , n804 , n10103 );
    not g30248 ( n28564 , n34754 );
    or g30249 ( n999 , n9329 , n18096 );
    or g30250 ( n28936 , n9532 , n32956 );
    not g30251 ( n4089 , n32696 );
    or g30252 ( n24520 , n6009 , n11988 );
    or g30253 ( n3771 , n1292 , n24193 );
    or g30254 ( n36351 , n16373 , n35048 );
    not g30255 ( n29474 , n3425 );
    and g30256 ( n21065 , n20463 , n22972 );
    not g30257 ( n42245 , n34479 );
    or g30258 ( n35239 , n7273 , n5096 );
    and g30259 ( n16197 , n7913 , n42768 );
    or g30260 ( n40123 , n27546 , n41532 );
    xnor g30261 ( n32576 , n8279 , n28670 );
    and g30262 ( n28148 , n15691 , n1761 );
    not g30263 ( n36953 , n18915 );
    nor g30264 ( n38093 , n6331 , n42284 );
    and g30265 ( n6694 , n25404 , n17628 );
    not g30266 ( n22946 , n25321 );
    or g30267 ( n6705 , n41249 , n25504 );
    and g30268 ( n31679 , n35905 , n17594 );
    not g30269 ( n28884 , n12098 );
    and g30270 ( n27416 , n5611 , n28905 );
    or g30271 ( n35940 , n38484 , n16188 );
    and g30272 ( n33274 , n33904 , n42002 );
    xnor g30273 ( n11884 , n7564 , n5677 );
    or g30274 ( n14717 , n31849 , n23859 );
    or g30275 ( n28973 , n33981 , n5411 );
    nor g30276 ( n19931 , n25076 , n41166 );
    xnor g30277 ( n1478 , n5341 , n38135 );
    nor g30278 ( n20688 , n42018 , n10452 );
    and g30279 ( n23547 , n39895 , n3513 );
    xnor g30280 ( n17162 , n40922 , n35609 );
    or g30281 ( n10798 , n9031 , n3245 );
    or g30282 ( n16969 , n26044 , n21225 );
    or g30283 ( n9396 , n87 , n24482 );
    and g30284 ( n7058 , n41773 , n27246 );
    not g30285 ( n15857 , n21257 );
    or g30286 ( n8385 , n32744 , n14184 );
    or g30287 ( n28315 , n40588 , n11615 );
    or g30288 ( n13164 , n26961 , n40400 );
    or g30289 ( n5553 , n11960 , n503 );
    and g30290 ( n20748 , n25052 , n33021 );
    xnor g30291 ( n5074 , n31099 , n39660 );
    xnor g30292 ( n13764 , n3232 , n13342 );
    or g30293 ( n13874 , n36815 , n11192 );
    or g30294 ( n9345 , n17827 , n15211 );
    or g30295 ( n26322 , n23232 , n36930 );
    or g30296 ( n20385 , n35732 , n2113 );
    not g30297 ( n34120 , n31847 );
    not g30298 ( n9513 , n36954 );
    nor g30299 ( n11234 , n4796 , n24611 );
    and g30300 ( n21481 , n23950 , n12183 );
    nor g30301 ( n26945 , n5823 , n5607 );
    or g30302 ( n28929 , n37183 , n17365 );
    or g30303 ( n15362 , n16530 , n4755 );
    and g30304 ( n28116 , n25120 , n28465 );
    or g30305 ( n30686 , n37399 , n19104 );
    not g30306 ( n32520 , n17107 );
    or g30307 ( n23484 , n34091 , n41258 );
    and g30308 ( n38152 , n17226 , n11041 );
    and g30309 ( n32901 , n2714 , n8065 );
    nor g30310 ( n19437 , n33596 , n10419 );
    or g30311 ( n37066 , n28400 , n36514 );
    or g30312 ( n15672 , n10818 , n6114 );
    nor g30313 ( n24189 , n2199 , n40004 );
    or g30314 ( n2683 , n22867 , n35269 );
    or g30315 ( n42222 , n28149 , n40577 );
    or g30316 ( n25452 , n27490 , n33075 );
    and g30317 ( n31354 , n41067 , n40684 );
    and g30318 ( n24699 , n12420 , n41417 );
    and g30319 ( n555 , n39682 , n7179 );
    and g30320 ( n15781 , n28280 , n25828 );
    not g30321 ( n22339 , n3366 );
    or g30322 ( n10109 , n26567 , n21413 );
    or g30323 ( n24763 , n22271 , n3210 );
    nor g30324 ( n27149 , n23914 , n39919 );
    not g30325 ( n17342 , n27223 );
    or g30326 ( n28574 , n15116 , n38392 );
    not g30327 ( n37176 , n18285 );
    and g30328 ( n18703 , n30698 , n41983 );
    or g30329 ( n20537 , n17714 , n757 );
    nor g30330 ( n22217 , n26617 , n12122 );
    or g30331 ( n0 , n3302 , n2802 );
    or g30332 ( n39424 , n27439 , n4752 );
    or g30333 ( n2028 , n34805 , n19618 );
    not g30334 ( n25784 , n22310 );
    or g30335 ( n29966 , n2095 , n34493 );
    and g30336 ( n33184 , n41377 , n30994 );
    and g30337 ( n25164 , n8137 , n10246 );
    and g30338 ( n41950 , n1942 , n19776 );
    xnor g30339 ( n5187 , n11029 , n3474 );
    not g30340 ( n41208 , n11524 );
    not g30341 ( n34363 , n34021 );
    nor g30342 ( n15436 , n10598 , n4580 );
    or g30343 ( n37343 , n4717 , n12610 );
    not g30344 ( n6865 , n25521 );
    or g30345 ( n33140 , n5356 , n23835 );
    or g30346 ( n33601 , n25675 , n11225 );
    not g30347 ( n16564 , n29987 );
    or g30348 ( n31908 , n42706 , n15639 );
    not g30349 ( n28956 , n37222 );
    not g30350 ( n25603 , n20124 );
    nor g30351 ( n34773 , n31582 , n18118 );
    or g30352 ( n33980 , n37891 , n14053 );
    or g30353 ( n29925 , n17124 , n8942 );
    nor g30354 ( n31491 , n38388 , n13161 );
    nor g30355 ( n9007 , n12885 , n7843 );
    nor g30356 ( n3024 , n7806 , n16111 );
    or g30357 ( n24865 , n423 , n2416 );
    xnor g30358 ( n7450 , n6767 , n10048 );
    or g30359 ( n31149 , n17814 , n14438 );
    and g30360 ( n41440 , n10004 , n7594 );
    or g30361 ( n17334 , n24635 , n10559 );
    xnor g30362 ( n12500 , n10814 , n16589 );
    xnor g30363 ( n36173 , n35377 , n22123 );
    not g30364 ( n34999 , n35873 );
    and g30365 ( n32070 , n24951 , n24969 );
    not g30366 ( n4911 , n23725 );
    xnor g30367 ( n8549 , n29886 , n18136 );
    or g30368 ( n4783 , n10724 , n41413 );
    or g30369 ( n14499 , n12152 , n5134 );
    and g30370 ( n18162 , n19060 , n17913 );
    nor g30371 ( n20476 , n33028 , n41831 );
    or g30372 ( n6752 , n35554 , n31271 );
    nor g30373 ( n24727 , n27722 , n4850 );
    or g30374 ( n26692 , n20723 , n34607 );
    and g30375 ( n25125 , n11009 , n15189 );
    or g30376 ( n22000 , n18165 , n14820 );
    or g30377 ( n35851 , n42115 , n5298 );
    and g30378 ( n31879 , n28104 , n4519 );
    or g30379 ( n36668 , n2958 , n35267 );
    and g30380 ( n39455 , n1423 , n37741 );
    or g30381 ( n12736 , n18798 , n36431 );
    or g30382 ( n18400 , n32173 , n11273 );
    or g30383 ( n39419 , n25996 , n25829 );
    nor g30384 ( n29013 , n41285 , n17501 );
    or g30385 ( n22384 , n23040 , n18593 );
    xnor g30386 ( n36391 , n9017 , n3075 );
    or g30387 ( n35690 , n11075 , n22472 );
    xnor g30388 ( n16883 , n36998 , n13852 );
    and g30389 ( n12322 , n37298 , n16716 );
    not g30390 ( n41641 , n39487 );
    and g30391 ( n21324 , n31817 , n6495 );
    and g30392 ( n25579 , n40893 , n24706 );
    or g30393 ( n18439 , n29514 , n3802 );
    or g30394 ( n608 , n19081 , n29147 );
    or g30395 ( n40079 , n39245 , n11456 );
    or g30396 ( n5244 , n24187 , n13951 );
    and g30397 ( n21655 , n2273 , n25980 );
    or g30398 ( n39638 , n425 , n9908 );
    xnor g30399 ( n38703 , n31314 , n7583 );
    or g30400 ( n29569 , n32792 , n35978 );
    nor g30401 ( n41349 , n1847 , n26838 );
    not g30402 ( n14635 , n2682 );
    nor g30403 ( n1337 , n19813 , n16912 );
    nor g30404 ( n38509 , n7723 , n32437 );
    and g30405 ( n7129 , n41050 , n21394 );
    or g30406 ( n29999 , n466 , n33330 );
    or g30407 ( n810 , n12700 , n16415 );
    or g30408 ( n10420 , n21150 , n999 );
    not g30409 ( n17137 , n28051 );
    and g30410 ( n12906 , n21635 , n33011 );
    not g30411 ( n5061 , n23059 );
    or g30412 ( n22679 , n37013 , n26359 );
    not g30413 ( n10910 , n14552 );
    not g30414 ( n38837 , n7362 );
    or g30415 ( n28557 , n15906 , n742 );
    or g30416 ( n7629 , n25602 , n41401 );
    not g30417 ( n2868 , n34414 );
    nor g30418 ( n42668 , n34292 , n25575 );
    or g30419 ( n7155 , n37808 , n11932 );
    or g30420 ( n7662 , n34294 , n41891 );
    xnor g30421 ( n26341 , n12146 , n23802 );
    or g30422 ( n2579 , n1827 , n22746 );
    or g30423 ( n27280 , n13974 , n5310 );
    or g30424 ( n29749 , n2088 , n41436 );
    and g30425 ( n34862 , n9664 , n13648 );
    not g30426 ( n15410 , n19895 );
    not g30427 ( n35287 , n16797 );
    xnor g30428 ( n574 , n2971 , n41062 );
    not g30429 ( n37805 , n16058 );
    nor g30430 ( n34881 , n5964 , n35375 );
    and g30431 ( n30251 , n42829 , n41198 );
    or g30432 ( n36825 , n36092 , n38404 );
    xnor g30433 ( n13045 , n39531 , n7873 );
    nor g30434 ( n27023 , n20860 , n11468 );
    or g30435 ( n28178 , n3664 , n11189 );
    not g30436 ( n41309 , n27162 );
    or g30437 ( n40935 , n29488 , n2586 );
    or g30438 ( n2346 , n23528 , n17455 );
    and g30439 ( n12549 , n31158 , n3286 );
    or g30440 ( n3653 , n6264 , n22797 );
    nor g30441 ( n7634 , n20429 , n7842 );
    nor g30442 ( n32347 , n7605 , n17391 );
    or g30443 ( n26057 , n10107 , n30820 );
    or g30444 ( n20079 , n15064 , n3380 );
    or g30445 ( n39888 , n5082 , n12030 );
    not g30446 ( n9271 , n36327 );
    or g30447 ( n34141 , n27377 , n28241 );
    xnor g30448 ( n22521 , n33341 , n1971 );
    or g30449 ( n26679 , n36275 , n7902 );
    xnor g30450 ( n17629 , n30200 , n21066 );
    nor g30451 ( n24698 , n15717 , n12366 );
    or g30452 ( n34046 , n24614 , n7220 );
    xnor g30453 ( n38413 , n39432 , n39553 );
    not g30454 ( n11702 , n33220 );
    xnor g30455 ( n34379 , n34945 , n29998 );
    or g30456 ( n35832 , n33546 , n41487 );
    not g30457 ( n21934 , n39429 );
    not g30458 ( n12332 , n33807 );
    xnor g30459 ( n6538 , n22543 , n19221 );
    nor g30460 ( n38167 , n22588 , n4841 );
    not g30461 ( n10278 , n36026 );
    nor g30462 ( n39690 , n26609 , n4701 );
    nor g30463 ( n9038 , n24567 , n2906 );
    or g30464 ( n31424 , n24656 , n35342 );
    or g30465 ( n6526 , n28887 , n8751 );
    xnor g30466 ( n40514 , n4538 , n20054 );
    xnor g30467 ( n8288 , n32930 , n7524 );
    or g30468 ( n12686 , n40259 , n21838 );
    and g30469 ( n1820 , n28957 , n23527 );
    or g30470 ( n12473 , n13685 , n36983 );
    nor g30471 ( n41031 , n10223 , n21019 );
    or g30472 ( n17440 , n217 , n38293 );
    and g30473 ( n22464 , n16458 , n29283 );
    and g30474 ( n41539 , n24084 , n1145 );
    or g30475 ( n37632 , n1792 , n6415 );
    not g30476 ( n2429 , n11473 );
    nor g30477 ( n37112 , n39266 , n31776 );
    xnor g30478 ( n31137 , n20376 , n21619 );
    or g30479 ( n33037 , n39292 , n2165 );
    xnor g30480 ( n37193 , n22577 , n36915 );
    or g30481 ( n12214 , n9061 , n27840 );
    xnor g30482 ( n36594 , n4302 , n14844 );
    not g30483 ( n22289 , n24453 );
    nor g30484 ( n15078 , n18843 , n25347 );
    or g30485 ( n26977 , n29761 , n27965 );
    nor g30486 ( n11412 , n22726 , n41405 );
    or g30487 ( n2071 , n23151 , n19152 );
    nor g30488 ( n42477 , n22490 , n29432 );
    xnor g30489 ( n28243 , n28864 , n36493 );
    and g30490 ( n36368 , n11501 , n30885 );
    or g30491 ( n35830 , n20412 , n15997 );
    and g30492 ( n6807 , n21927 , n27209 );
    nor g30493 ( n41849 , n1507 , n4403 );
    and g30494 ( n14894 , n18714 , n39653 );
    and g30495 ( n30165 , n27751 , n12965 );
    xnor g30496 ( n36017 , n784 , n13244 );
    and g30497 ( n10430 , n19272 , n13302 );
    and g30498 ( n33985 , n544 , n24548 );
    or g30499 ( n17734 , n15753 , n12443 );
    or g30500 ( n34601 , n3749 , n403 );
    not g30501 ( n39532 , n31764 );
    not g30502 ( n22538 , n101 );
    or g30503 ( n35609 , n22299 , n26070 );
    not g30504 ( n22340 , n9882 );
    or g30505 ( n37307 , n26713 , n31663 );
    not g30506 ( n29834 , n24976 );
    or g30507 ( n35071 , n20883 , n27127 );
    and g30508 ( n24565 , n25354 , n28277 );
    or g30509 ( n8929 , n1685 , n25722 );
    or g30510 ( n32561 , n39118 , n21080 );
    and g30511 ( n31702 , n5144 , n21551 );
    or g30512 ( n13803 , n8861 , n16471 );
    or g30513 ( n29802 , n34520 , n14672 );
    nor g30514 ( n33042 , n15936 , n30974 );
    and g30515 ( n34711 , n16580 , n20929 );
    or g30516 ( n1428 , n17277 , n26132 );
    not g30517 ( n10625 , n4404 );
    xnor g30518 ( n7694 , n4795 , n31303 );
    xnor g30519 ( n25319 , n35786 , n4878 );
    xnor g30520 ( n13924 , n2338 , n8963 );
    xnor g30521 ( n9072 , n22781 , n4104 );
    not g30522 ( n25043 , n40225 );
    not g30523 ( n5415 , n35987 );
    or g30524 ( n38675 , n42369 , n13032 );
    nor g30525 ( n15033 , n33840 , n39263 );
    xnor g30526 ( n7693 , n28319 , n9601 );
    xnor g30527 ( n27529 , n35246 , n16003 );
    and g30528 ( n33287 , n2634 , n11521 );
    or g30529 ( n23596 , n1414 , n23031 );
    or g30530 ( n34657 , n41601 , n29469 );
    or g30531 ( n25287 , n30599 , n38345 );
    or g30532 ( n23836 , n3038 , n34569 );
    or g30533 ( n41204 , n42055 , n39528 );
    and g30534 ( n17900 , n26958 , n19042 );
    not g30535 ( n29777 , n33702 );
    or g30536 ( n371 , n11078 , n27116 );
    or g30537 ( n25880 , n30358 , n21324 );
    or g30538 ( n38018 , n6989 , n12668 );
    not g30539 ( n3856 , n35221 );
    xnor g30540 ( n24199 , n509 , n34532 );
    not g30541 ( n34939 , n6032 );
    xnor g30542 ( n36290 , n34951 , n37957 );
    xnor g30543 ( n42196 , n784 , n15012 );
    nor g30544 ( n19218 , n37671 , n14985 );
    nor g30545 ( n39277 , n8953 , n6732 );
    or g30546 ( n39934 , n32892 , n17536 );
    or g30547 ( n39179 , n11472 , n21216 );
    and g30548 ( n38986 , n16252 , n27456 );
    or g30549 ( n22386 , n28935 , n20633 );
    xnor g30550 ( n27694 , n41013 , n19163 );
    nor g30551 ( n8053 , n8271 , n42281 );
    or g30552 ( n3624 , n28344 , n9045 );
    or g30553 ( n42493 , n12803 , n3728 );
    or g30554 ( n14777 , n34594 , n34893 );
    or g30555 ( n12280 , n38565 , n23272 );
    and g30556 ( n26874 , n11304 , n4419 );
    not g30557 ( n20574 , n42169 );
    xnor g30558 ( n25724 , n1651 , n15070 );
    nor g30559 ( n12372 , n33269 , n31223 );
    or g30560 ( n35788 , n39828 , n5033 );
    nor g30561 ( n6168 , n8494 , n15639 );
    or g30562 ( n18932 , n19479 , n29325 );
    or g30563 ( n13263 , n29942 , n33973 );
    and g30564 ( n32179 , n12774 , n17603 );
    or g30565 ( n27212 , n26974 , n34974 );
    and g30566 ( n39825 , n29133 , n41185 );
    nor g30567 ( n3655 , n32446 , n13670 );
    nor g30568 ( n12830 , n24264 , n24480 );
    or g30569 ( n9100 , n29841 , n30350 );
    not g30570 ( n6545 , n33701 );
    or g30571 ( n35007 , n33022 , n3623 );
    or g30572 ( n14015 , n26885 , n33609 );
    xnor g30573 ( n5640 , n2921 , n24840 );
    and g30574 ( n32258 , n28178 , n33805 );
    and g30575 ( n6837 , n35196 , n16855 );
    or g30576 ( n4603 , n8033 , n24219 );
    or g30577 ( n1106 , n20051 , n33556 );
    and g30578 ( n24238 , n11802 , n41222 );
    xnor g30579 ( n30721 , n4334 , n30269 );
    not g30580 ( n17596 , n16811 );
    and g30581 ( n30395 , n38236 , n536 );
    not g30582 ( n19701 , n17252 );
    xnor g30583 ( n39462 , n27904 , n18866 );
    nor g30584 ( n28997 , n35796 , n31719 );
    and g30585 ( n12652 , n4445 , n38452 );
    xnor g30586 ( n18334 , n38140 , n28323 );
    and g30587 ( n41897 , n13472 , n8060 );
    or g30588 ( n9143 , n26269 , n33285 );
    and g30589 ( n3033 , n17541 , n38903 );
    xnor g30590 ( n2988 , n23746 , n874 );
    or g30591 ( n29641 , n34202 , n34638 );
    not g30592 ( n19665 , n17454 );
    or g30593 ( n16549 , n34433 , n7335 );
    not g30594 ( n13857 , n40586 );
    or g30595 ( n2955 , n5299 , n23258 );
    or g30596 ( n22995 , n1390 , n26041 );
    xnor g30597 ( n17058 , n9133 , n34041 );
    xnor g30598 ( n31868 , n4385 , n839 );
    or g30599 ( n9013 , n28605 , n32235 );
    or g30600 ( n32268 , n3951 , n25863 );
    not g30601 ( n2486 , n24825 );
    xnor g30602 ( n42317 , n32779 , n823 );
    not g30603 ( n35265 , n14041 );
    xnor g30604 ( n21935 , n12146 , n23558 );
    or g30605 ( n11946 , n27103 , n34939 );
    nor g30606 ( n7263 , n38566 , n12763 );
    not g30607 ( n37337 , n32530 );
    nor g30608 ( n26758 , n36117 , n23453 );
    or g30609 ( n34240 , n13619 , n33542 );
    or g30610 ( n11983 , n23895 , n3845 );
    and g30611 ( n36553 , n31906 , n25772 );
    not g30612 ( n22409 , n41669 );
    xnor g30613 ( n27364 , n23686 , n22911 );
    xnor g30614 ( n39336 , n19592 , n7435 );
    nor g30615 ( n37761 , n14131 , n24419 );
    nor g30616 ( n13391 , n19813 , n23042 );
    and g30617 ( n32224 , n1739 , n38619 );
    not g30618 ( n10555 , n37187 );
    or g30619 ( n24987 , n41767 , n33864 );
    xnor g30620 ( n23649 , n13133 , n16419 );
    or g30621 ( n39162 , n5635 , n27857 );
    or g30622 ( n27887 , n9673 , n14987 );
    and g30623 ( n30008 , n6223 , n41918 );
    or g30624 ( n25675 , n40350 , n26696 );
    not g30625 ( n42110 , n25505 );
    and g30626 ( n7118 , n33018 , n4042 );
    nor g30627 ( n37778 , n5964 , n31399 );
    nor g30628 ( n29832 , n40590 , n9139 );
    not g30629 ( n40090 , n26056 );
    or g30630 ( n18234 , n23085 , n7912 );
    xnor g30631 ( n19855 , n21598 , n40885 );
    not g30632 ( n40588 , n41321 );
    not g30633 ( n32470 , n7125 );
    nor g30634 ( n22299 , n6742 , n23253 );
    or g30635 ( n35873 , n9382 , n39188 );
    or g30636 ( n17487 , n27712 , n10007 );
    nor g30637 ( n40223 , n18997 , n22988 );
    nor g30638 ( n18425 , n27613 , n24051 );
    or g30639 ( n30009 , n30235 , n40498 );
    xnor g30640 ( n3075 , n71 , n4119 );
    or g30641 ( n36940 , n14433 , n35193 );
    or g30642 ( n41330 , n16915 , n436 );
    or g30643 ( n39874 , n15482 , n35572 );
    and g30644 ( n42730 , n2947 , n715 );
    or g30645 ( n29146 , n14407 , n28336 );
    or g30646 ( n10216 , n19890 , n5707 );
    and g30647 ( n38218 , n24209 , n26833 );
    and g30648 ( n10081 , n21042 , n22601 );
    or g30649 ( n21625 , n32645 , n15573 );
    and g30650 ( n13396 , n30324 , n41151 );
    not g30651 ( n29636 , n34624 );
    or g30652 ( n1132 , n15191 , n31244 );
    not g30653 ( n11376 , n2654 );
    and g30654 ( n27878 , n1958 , n20108 );
    nor g30655 ( n27929 , n34761 , n37384 );
    and g30656 ( n30020 , n35194 , n7449 );
    or g30657 ( n27307 , n3992 , n20219 );
    and g30658 ( n10987 , n38542 , n9152 );
    and g30659 ( n38038 , n32400 , n24916 );
    xnor g30660 ( n2068 , n14226 , n13883 );
    xnor g30661 ( n25482 , n1110 , n26795 );
    or g30662 ( n18886 , n28863 , n23760 );
    xnor g30663 ( n34346 , n24278 , n11152 );
    or g30664 ( n33713 , n38556 , n26479 );
    not g30665 ( n29423 , n19508 );
    and g30666 ( n19682 , n3849 , n9963 );
    nor g30667 ( n5934 , n27572 , n9424 );
    nor g30668 ( n36926 , n26371 , n27706 );
    not g30669 ( n36365 , n41847 );
    xnor g30670 ( n30958 , n39237 , n5964 );
    and g30671 ( n2814 , n3151 , n12241 );
    or g30672 ( n13898 , n2592 , n7737 );
    or g30673 ( n33983 , n1790 , n32551 );
    nor g30674 ( n2499 , n5964 , n17678 );
    nor g30675 ( n29126 , n1219 , n2039 );
    or g30676 ( n35084 , n9680 , n29930 );
    or g30677 ( n21425 , n27836 , n14807 );
    or g30678 ( n28694 , n39332 , n42595 );
    or g30679 ( n11088 , n13635 , n27179 );
    and g30680 ( n24953 , n29923 , n8388 );
    and g30681 ( n5282 , n6424 , n27491 );
    nor g30682 ( n16663 , n29087 , n15859 );
    or g30683 ( n36035 , n12252 , n17972 );
    or g30684 ( n15885 , n28406 , n24560 );
    and g30685 ( n36575 , n26434 , n16130 );
    xnor g30686 ( n37734 , n12876 , n27819 );
    and g30687 ( n19478 , n18755 , n21921 );
    and g30688 ( n22652 , n31718 , n27845 );
    or g30689 ( n373 , n11942 , n14281 );
    not g30690 ( n10163 , n32399 );
    and g30691 ( n16925 , n33266 , n8802 );
    and g30692 ( n13955 , n12079 , n33125 );
    nor g30693 ( n33853 , n32412 , n41232 );
    or g30694 ( n17357 , n994 , n24996 );
    not g30695 ( n30611 , n14206 );
    or g30696 ( n15380 , n36845 , n11981 );
    xnor g30697 ( n6840 , n39532 , n13645 );
    and g30698 ( n27632 , n2918 , n41041 );
    or g30699 ( n38220 , n23763 , n10299 );
    xnor g30700 ( n40717 , n40 , n26276 );
    and g30701 ( n29367 , n40156 , n39562 );
    or g30702 ( n19656 , n34489 , n12340 );
    or g30703 ( n17375 , n35051 , n25704 );
    and g30704 ( n5543 , n24129 , n4142 );
    nor g30705 ( n21082 , n4872 , n4550 );
    and g30706 ( n7547 , n26852 , n23967 );
    and g30707 ( n37073 , n17283 , n25712 );
    not g30708 ( n22530 , n34239 );
    and g30709 ( n9302 , n38769 , n33913 );
    not g30710 ( n25364 , n852 );
    not g30711 ( n39760 , n41208 );
    xnor g30712 ( n25995 , n32624 , n25543 );
    xnor g30713 ( n8335 , n33617 , n7209 );
    and g30714 ( n30214 , n6248 , n37744 );
    xnor g30715 ( n3973 , n4872 , n28505 );
    nor g30716 ( n30935 , n21286 , n1261 );
    and g30717 ( n10028 , n30411 , n40758 );
    xnor g30718 ( n36828 , n1863 , n15751 );
    or g30719 ( n6146 , n22619 , n23138 );
    or g30720 ( n16778 , n28732 , n12210 );
    and g30721 ( n19371 , n33564 , n31272 );
    or g30722 ( n27826 , n34537 , n6024 );
    or g30723 ( n40029 , n29033 , n23738 );
    or g30724 ( n30191 , n35386 , n21624 );
    and g30725 ( n3290 , n20357 , n21890 );
    not g30726 ( n32256 , n2253 );
    or g30727 ( n18759 , n20112 , n35677 );
    and g30728 ( n9794 , n8278 , n29953 );
    and g30729 ( n36383 , n8912 , n39454 );
    and g30730 ( n3151 , n33044 , n2238 );
    xnor g30731 ( n7164 , n5041 , n20375 );
    and g30732 ( n39203 , n30475 , n9830 );
    not g30733 ( n21192 , n14870 );
    not g30734 ( n31073 , n30487 );
    or g30735 ( n20664 , n2199 , n27640 );
    xnor g30736 ( n9507 , n11436 , n9823 );
    not g30737 ( n11581 , n32945 );
    nor g30738 ( n37581 , n6278 , n2156 );
    or g30739 ( n12485 , n3719 , n35531 );
    and g30740 ( n39781 , n8877 , n6998 );
    not g30741 ( n5408 , n13886 );
    or g30742 ( n20097 , n5981 , n37806 );
    not g30743 ( n35657 , n26782 );
    or g30744 ( n42853 , n16052 , n40333 );
    and g30745 ( n35306 , n14881 , n30195 );
    or g30746 ( n7451 , n34208 , n1551 );
    or g30747 ( n34923 , n13367 , n21923 );
    xnor g30748 ( n31224 , n2903 , n29051 );
    or g30749 ( n29871 , n5793 , n12456 );
    or g30750 ( n42355 , n6702 , n13383 );
    or g30751 ( n24364 , n968 , n29361 );
    and g30752 ( n30613 , n30996 , n23737 );
    xnor g30753 ( n20870 , n32160 , n5298 );
    or g30754 ( n35504 , n2012 , n17788 );
    and g30755 ( n23009 , n32349 , n662 );
    and g30756 ( n6635 , n29882 , n3285 );
    or g30757 ( n32582 , n7410 , n22552 );
    or g30758 ( n28603 , n36284 , n34006 );
    and g30759 ( n37294 , n39656 , n39716 );
    not g30760 ( n23389 , n36917 );
    not g30761 ( n31785 , n21975 );
    nor g30762 ( n22505 , n23311 , n25543 );
    or g30763 ( n3478 , n32599 , n28825 );
    not g30764 ( n28174 , n27760 );
    and g30765 ( n4786 , n654 , n15022 );
    not g30766 ( n30592 , n36912 );
    or g30767 ( n18713 , n17244 , n29242 );
    or g30768 ( n7545 , n14988 , n11314 );
    not g30769 ( n32898 , n23106 );
    or g30770 ( n41189 , n7543 , n25612 );
    or g30771 ( n32306 , n41001 , n7868 );
    xnor g30772 ( n9843 , n9783 , n33903 );
    or g30773 ( n21674 , n868 , n25506 );
    not g30774 ( n21300 , n21734 );
    or g30775 ( n41801 , n13820 , n17425 );
    and g30776 ( n4006 , n12380 , n16322 );
    xnor g30777 ( n38609 , n14740 , n7647 );
    or g30778 ( n5636 , n8826 , n26854 );
    or g30779 ( n4380 , n15780 , n5997 );
    xnor g30780 ( n31194 , n39798 , n35161 );
    xnor g30781 ( n14517 , n14502 , n33502 );
    or g30782 ( n8917 , n41433 , n39849 );
    or g30783 ( n6513 , n35968 , n28220 );
    or g30784 ( n31872 , n13450 , n28599 );
    not g30785 ( n24810 , n30826 );
    or g30786 ( n34405 , n38249 , n4801 );
    or g30787 ( n10264 , n20135 , n19461 );
    xnor g30788 ( n38785 , n42127 , n42631 );
    nor g30789 ( n754 , n15070 , n23802 );
    not g30790 ( n38621 , n38545 );
    or g30791 ( n39871 , n4535 , n40951 );
    and g30792 ( n9766 , n7195 , n3329 );
    or g30793 ( n21878 , n5168 , n27303 );
    or g30794 ( n23506 , n28488 , n9206 );
    or g30795 ( n26263 , n1971 , n6436 );
    nor g30796 ( n13143 , n37148 , n29727 );
    or g30797 ( n28138 , n2437 , n25178 );
    and g30798 ( n23555 , n14670 , n10933 );
    and g30799 ( n27320 , n25384 , n9976 );
    xnor g30800 ( n21291 , n29476 , n35374 );
    nor g30801 ( n7229 , n25588 , n7256 );
    xnor g30802 ( n36875 , n32254 , n41486 );
    or g30803 ( n36254 , n13704 , n40872 );
    or g30804 ( n19932 , n40578 , n13467 );
    and g30805 ( n2516 , n16961 , n21056 );
    or g30806 ( n13485 , n7413 , n27210 );
    and g30807 ( n33291 , n110 , n26662 );
    xnor g30808 ( n2998 , n26691 , n10073 );
    or g30809 ( n25749 , n30273 , n1404 );
    or g30810 ( n1221 , n13147 , n41487 );
    and g30811 ( n33828 , n22710 , n24208 );
    and g30812 ( n18772 , n42354 , n19757 );
    or g30813 ( n33329 , n8398 , n24020 );
    or g30814 ( n5609 , n14298 , n32942 );
    and g30815 ( n1895 , n3479 , n41771 );
    or g30816 ( n8356 , n4670 , n24835 );
    or g30817 ( n24632 , n28167 , n14153 );
    or g30818 ( n13153 , n40804 , n33797 );
    not g30819 ( n38506 , n12249 );
    or g30820 ( n5676 , n11880 , n173 );
    and g30821 ( n41099 , n19943 , n35335 );
    or g30822 ( n9707 , n2011 , n19768 );
    and g30823 ( n17620 , n31462 , n42219 );
    nor g30824 ( n26427 , n25679 , n6519 );
    or g30825 ( n23188 , n21258 , n17680 );
    nor g30826 ( n10945 , n1935 , n11002 );
    or g30827 ( n3319 , n6575 , n31693 );
    not g30828 ( n2892 , n11264 );
    nor g30829 ( n41061 , n41704 , n2590 );
    or g30830 ( n37488 , n7601 , n21019 );
    and g30831 ( n26193 , n30249 , n37775 );
    and g30832 ( n19206 , n39989 , n36188 );
    or g30833 ( n494 , n33624 , n6859 );
    not g30834 ( n8758 , n5623 );
    nor g30835 ( n29216 , n39367 , n21221 );
    and g30836 ( n21430 , n12734 , n11836 );
    not g30837 ( n26739 , n22782 );
    xnor g30838 ( n4566 , n11147 , n33923 );
    xnor g30839 ( n19610 , n42761 , n36170 );
    or g30840 ( n28523 , n14386 , n31756 );
    or g30841 ( n9101 , n2032 , n37296 );
    and g30842 ( n39702 , n33962 , n15312 );
    and g30843 ( n8613 , n2001 , n34531 );
    or g30844 ( n29606 , n8187 , n33047 );
    nor g30845 ( n26631 , n27137 , n36795 );
    or g30846 ( n24688 , n4169 , n39059 );
    and g30847 ( n35747 , n11509 , n23444 );
    not g30848 ( n27098 , n23516 );
    not g30849 ( n14515 , n31785 );
    or g30850 ( n13776 , n37498 , n24516 );
    xnor g30851 ( n13483 , n31239 , n28703 );
    nor g30852 ( n39245 , n35573 , n35314 );
    nor g30853 ( n3212 , n11782 , n15266 );
    and g30854 ( n17924 , n27104 , n33507 );
    xnor g30855 ( n36704 , n6625 , n18567 );
    or g30856 ( n10995 , n42307 , n39839 );
    or g30857 ( n30076 , n13756 , n31527 );
    nor g30858 ( n20575 , n27159 , n42242 );
    or g30859 ( n30716 , n18144 , n33537 );
    and g30860 ( n1294 , n30729 , n28972 );
    not g30861 ( n16215 , n7221 );
    not g30862 ( n32701 , n23004 );
    or g30863 ( n30497 , n26736 , n29750 );
    or g30864 ( n31904 , n9952 , n18629 );
    and g30865 ( n39672 , n38566 , n12763 );
    and g30866 ( n9722 , n15682 , n10441 );
    not g30867 ( n18496 , n26201 );
    or g30868 ( n21590 , n6628 , n10360 );
    nor g30869 ( n12782 , n7356 , n11478 );
    not g30870 ( n39790 , n31118 );
    xnor g30871 ( n7644 , n6625 , n6550 );
    or g30872 ( n27190 , n42131 , n32586 );
    xnor g30873 ( n23205 , n34352 , n21535 );
    nor g30874 ( n40293 , n19547 , n35489 );
    not g30875 ( n14388 , n35195 );
    or g30876 ( n16291 , n7714 , n19104 );
    or g30877 ( n19859 , n5041 , n29392 );
    not g30878 ( n1339 , n35984 );
    or g30879 ( n39711 , n21703 , n18788 );
    or g30880 ( n37359 , n34704 , n30114 );
    and g30881 ( n38387 , n14332 , n15275 );
    and g30882 ( n4550 , n31755 , n7274 );
    not g30883 ( n33027 , n7986 );
    or g30884 ( n38664 , n24547 , n8111 );
    or g30885 ( n696 , n18666 , n17249 );
    or g30886 ( n11869 , n21373 , n10009 );
    xnor g30887 ( n42653 , n1499 , n29969 );
    xnor g30888 ( n29891 , n9264 , n14791 );
    xnor g30889 ( n39080 , n23945 , n27339 );
    not g30890 ( n11380 , n11353 );
    or g30891 ( n40583 , n23426 , n9456 );
    nor g30892 ( n39126 , n22173 , n17343 );
    or g30893 ( n14921 , n28468 , n9891 );
    or g30894 ( n41212 , n25149 , n1289 );
    xnor g30895 ( n3335 , n29056 , n18639 );
    or g30896 ( n40797 , n14013 , n40310 );
    xnor g30897 ( n11154 , n2130 , n7213 );
    or g30898 ( n370 , n15763 , n37029 );
    or g30899 ( n36257 , n440 , n28856 );
    or g30900 ( n5939 , n12968 , n7196 );
    nor g30901 ( n6445 , n22100 , n12778 );
    or g30902 ( n27043 , n3902 , n8636 );
    or g30903 ( n3059 , n11229 , n23895 );
    and g30904 ( n18016 , n9367 , n8158 );
    and g30905 ( n32124 , n34591 , n23838 );
    and g30906 ( n40539 , n41803 , n40778 );
    or g30907 ( n3342 , n35337 , n15481 );
    and g30908 ( n23059 , n31086 , n24730 );
    or g30909 ( n37594 , n13281 , n15505 );
    xnor g30910 ( n26763 , n26 , n30371 );
    and g30911 ( n35890 , n42212 , n21986 );
    not g30912 ( n19079 , n13741 );
    nor g30913 ( n2982 , n35331 , n8354 );
    not g30914 ( n19282 , n41208 );
    xnor g30915 ( n5180 , n26892 , n7519 );
    not g30916 ( n5585 , n33803 );
    or g30917 ( n26289 , n22427 , n7513 );
    not g30918 ( n18190 , n28940 );
    xnor g30919 ( n15830 , n13929 , n39588 );
    xnor g30920 ( n6005 , n17038 , n23876 );
    or g30921 ( n29242 , n12101 , n12484 );
    or g30922 ( n34513 , n10496 , n36023 );
    not g30923 ( n15495 , n246 );
    or g30924 ( n4568 , n41475 , n41100 );
    nor g30925 ( n15625 , n24264 , n10068 );
    not g30926 ( n19540 , n42652 );
    or g30927 ( n11429 , n29120 , n1173 );
    and g30928 ( n9085 , n38108 , n607 );
    and g30929 ( n25507 , n13936 , n33009 );
    nor g30930 ( n38011 , n28650 , n32140 );
    or g30931 ( n22329 , n5964 , n15277 );
    or g30932 ( n38341 , n20093 , n2013 );
    not g30933 ( n33285 , n13960 );
    or g30934 ( n15459 , n40512 , n27211 );
    or g30935 ( n11062 , n6900 , n21048 );
    xnor g30936 ( n32634 , n7980 , n38078 );
    or g30937 ( n41219 , n38591 , n37749 );
    xnor g30938 ( n38290 , n29740 , n18788 );
    nor g30939 ( n18767 , n41715 , n5952 );
    or g30940 ( n11207 , n39478 , n27240 );
    or g30941 ( n27244 , n34485 , n35160 );
    nor g30942 ( n14646 , n24819 , n7359 );
    not g30943 ( n24546 , n37873 );
    and g30944 ( n5335 , n9228 , n9975 );
    or g30945 ( n26437 , n10051 , n10953 );
    and g30946 ( n35936 , n28458 , n4382 );
    and g30947 ( n38433 , n852 , n32838 );
    nor g30948 ( n21453 , n23792 , n24116 );
    not g30949 ( n19613 , n30579 );
    or g30950 ( n30656 , n32277 , n27363 );
    or g30951 ( n26267 , n25313 , n30383 );
    and g30952 ( n30471 , n22418 , n23544 );
    and g30953 ( n18988 , n26047 , n36841 );
    or g30954 ( n8237 , n24849 , n2827 );
    xnor g30955 ( n41826 , n40 , n31186 );
    and g30956 ( n29403 , n39969 , n20943 );
    nor g30957 ( n20270 , n7479 , n21019 );
    or g30958 ( n32272 , n1133 , n41148 );
    or g30959 ( n19677 , n36296 , n33036 );
    or g30960 ( n32504 , n15362 , n9419 );
    not g30961 ( n27627 , n21480 );
    nor g30962 ( n39274 , n17945 , n18913 );
    not g30963 ( n17970 , n22607 );
    or g30964 ( n34321 , n35807 , n9958 );
    or g30965 ( n33682 , n42515 , n16287 );
    and g30966 ( n20283 , n20342 , n393 );
    or g30967 ( n38759 , n40266 , n24072 );
    nor g30968 ( n39258 , n36561 , n11724 );
    and g30969 ( n5365 , n28196 , n14 );
    not g30970 ( n972 , n38555 );
    not g30971 ( n8625 , n32291 );
    or g30972 ( n7762 , n9678 , n36222 );
    not g30973 ( n34826 , n3045 );
    not g30974 ( n15406 , n15331 );
    xnor g30975 ( n12208 , n5144 , n32877 );
    and g30976 ( n17145 , n8269 , n17329 );
    nor g30977 ( n677 , n3080 , n9851 );
    nor g30978 ( n33710 , n11847 , n21324 );
    or g30979 ( n12719 , n2768 , n2047 );
    and g30980 ( n17215 , n11283 , n31388 );
    or g30981 ( n25476 , n35452 , n20759 );
    xnor g30982 ( n7445 , n36362 , n18223 );
    and g30983 ( n35577 , n10949 , n4966 );
    or g30984 ( n17801 , n1067 , n36344 );
    nor g30985 ( n6685 , n36117 , n10958 );
    not g30986 ( n16108 , n41937 );
    and g30987 ( n42454 , n19219 , n4471 );
    not g30988 ( n30738 , n1986 );
    xnor g30989 ( n3429 , n41718 , n5256 );
    and g30990 ( n28535 , n23291 , n28676 );
    not g30991 ( n24172 , n42092 );
    xnor g30992 ( n19576 , n34444 , n27340 );
    or g30993 ( n37215 , n11306 , n12669 );
    not g30994 ( n16109 , n20393 );
    and g30995 ( n1267 , n35579 , n40704 );
    and g30996 ( n38618 , n12649 , n8197 );
    and g30997 ( n10665 , n22324 , n40166 );
    or g30998 ( n41368 , n6247 , n22213 );
    not g30999 ( n40053 , n3783 );
    or g31000 ( n32596 , n28488 , n42850 );
    nor g31001 ( n33104 , n2482 , n2930 );
    and g31002 ( n19327 , n4418 , n16201 );
    or g31003 ( n6202 , n22821 , n27507 );
    and g31004 ( n25561 , n33351 , n23564 );
    and g31005 ( n26342 , n15643 , n21573 );
    nor g31006 ( n30296 , n40875 , n36890 );
    or g31007 ( n22626 , n19247 , n38691 );
    and g31008 ( n2304 , n35400 , n32838 );
    not g31009 ( n23683 , n15543 );
    nor g31010 ( n17952 , n19292 , n23816 );
    and g31011 ( n17204 , n41281 , n36126 );
    or g31012 ( n15754 , n35046 , n20021 );
    not g31013 ( n42706 , n30845 );
    or g31014 ( n30321 , n30820 , n22033 );
    or g31015 ( n16011 , n31641 , n33670 );
    and g31016 ( n23354 , n25369 , n36668 );
    and g31017 ( n34917 , n37936 , n8575 );
    or g31018 ( n38172 , n30235 , n27195 );
    xnor g31019 ( n10831 , n27371 , n38547 );
    and g31020 ( n37680 , n38551 , n337 );
    not g31021 ( n23311 , n19508 );
    and g31022 ( n32606 , n20316 , n24928 );
    nor g31023 ( n37367 , n16998 , n35300 );
    not g31024 ( n9312 , n25835 );
    and g31025 ( n9089 , n38148 , n36586 );
    and g31026 ( n13859 , n37544 , n30794 );
    and g31027 ( n40420 , n37377 , n15939 );
    not g31028 ( n14611 , n6840 );
    xnor g31029 ( n26839 , n27843 , n19703 );
    or g31030 ( n23089 , n18778 , n37243 );
    xnor g31031 ( n10443 , n37437 , n40252 );
    and g31032 ( n28900 , n3205 , n4162 );
    and g31033 ( n29533 , n13089 , n30015 );
    or g31034 ( n18994 , n12149 , n31248 );
    or g31035 ( n30441 , n19264 , n12672 );
    or g31036 ( n3576 , n25259 , n38691 );
    not g31037 ( n36019 , n34940 );
    not g31038 ( n1375 , n17117 );
    not g31039 ( n17234 , n26032 );
    or g31040 ( n8939 , n33755 , n21176 );
    or g31041 ( n6556 , n38157 , n9750 );
    or g31042 ( n40026 , n36687 , n14218 );
    not g31043 ( n7109 , n40152 );
    xnor g31044 ( n34736 , n29740 , n35339 );
    xnor g31045 ( n26123 , n26 , n16318 );
    not g31046 ( n16661 , n13256 );
    xnor g31047 ( n9992 , n32160 , n41848 );
    and g31048 ( n33137 , n42071 , n20689 );
    not g31049 ( n24482 , n27654 );
    nor g31050 ( n10119 , n16431 , n14017 );
    and g31051 ( n31436 , n28895 , n40530 );
    nor g31052 ( n8192 , n40156 , n35449 );
    not g31053 ( n154 , n13871 );
    or g31054 ( n41172 , n13185 , n22118 );
    or g31055 ( n5616 , n30919 , n39499 );
    not g31056 ( n38288 , n14810 );
    or g31057 ( n11571 , n11696 , n10704 );
    and g31058 ( n35023 , n4581 , n13972 );
    and g31059 ( n6911 , n7937 , n32304 );
    xnor g31060 ( n36541 , n41013 , n22618 );
    and g31061 ( n35883 , n30415 , n8079 );
    xnor g31062 ( n2079 , n27418 , n24619 );
    xnor g31063 ( n9891 , n30562 , n12815 );
    and g31064 ( n10346 , n4977 , n32862 );
    nor g31065 ( n30116 , n20307 , n6329 );
    and g31066 ( n33129 , n3797 , n30819 );
    and g31067 ( n24992 , n42475 , n39726 );
    or g31068 ( n35039 , n37645 , n6612 );
    or g31069 ( n35668 , n27563 , n14137 );
    not g31070 ( n7863 , n21466 );
    and g31071 ( n16067 , n29109 , n15535 );
    and g31072 ( n30153 , n40861 , n26048 );
    xnor g31073 ( n24952 , n23180 , n31384 );
    or g31074 ( n37267 , n6168 , n25194 );
    not g31075 ( n27189 , n21389 );
    not g31076 ( n4758 , n17085 );
    or g31077 ( n23512 , n19371 , n20078 );
    or g31078 ( n5283 , n11050 , n38956 );
    and g31079 ( n37105 , n20749 , n32516 );
    nor g31080 ( n21679 , n13243 , n13422 );
    and g31081 ( n15866 , n42445 , n26200 );
    or g31082 ( n12855 , n21269 , n41494 );
    and g31083 ( n15370 , n12384 , n34342 );
    and g31084 ( n27205 , n42808 , n5521 );
    xnor g31085 ( n21742 , n28252 , n16657 );
    nor g31086 ( n20200 , n17170 , n14260 );
    or g31087 ( n606 , n31845 , n14600 );
    and g31088 ( n32111 , n40802 , n10357 );
    not g31089 ( n34474 , n6651 );
    not g31090 ( n3101 , n7946 );
    and g31091 ( n21882 , n41611 , n36305 );
    and g31092 ( n27210 , n19718 , n34077 );
    not g31093 ( n5246 , n26358 );
    or g31094 ( n14396 , n32785 , n1289 );
    or g31095 ( n27651 , n41923 , n23450 );
    not g31096 ( n6023 , n29582 );
    xnor g31097 ( n11657 , n784 , n22480 );
    nor g31098 ( n24331 , n6116 , n40977 );
    or g31099 ( n7174 , n14616 , n11986 );
    or g31100 ( n32788 , n26921 , n2988 );
    and g31101 ( n32007 , n12701 , n31448 );
    nor g31102 ( n1012 , n38879 , n12258 );
    nor g31103 ( n27453 , n42115 , n6393 );
    nor g31104 ( n23748 , n1781 , n27364 );
    and g31105 ( n5161 , n5319 , n37691 );
    or g31106 ( n40217 , n32578 , n26149 );
    xnor g31107 ( n12946 , n27035 , n2992 );
    or g31108 ( n5765 , n3317 , n18877 );
    or g31109 ( n18867 , n42537 , n39828 );
    and g31110 ( n31573 , n10102 , n14846 );
    and g31111 ( n203 , n22241 , n28017 );
    or g31112 ( n37518 , n20243 , n1959 );
    and g31113 ( n20763 , n31935 , n8845 );
    and g31114 ( n29571 , n40179 , n2640 );
    or g31115 ( n2452 , n38196 , n41099 );
    not g31116 ( n4592 , n22444 );
    xnor g31117 ( n42907 , n4492 , n37902 );
    and g31118 ( n24157 , n17136 , n42690 );
    nor g31119 ( n9415 , n24742 , n7926 );
    and g31120 ( n6092 , n12613 , n33161 );
    or g31121 ( n38499 , n25964 , n24697 );
    and g31122 ( n20821 , n22084 , n23596 );
    nor g31123 ( n21828 , n32289 , n42164 );
    or g31124 ( n7718 , n7056 , n9398 );
    or g31125 ( n25235 , n27578 , n19843 );
    or g31126 ( n2123 , n27379 , n42264 );
    not g31127 ( n36445 , n127 );
    or g31128 ( n14850 , n10098 , n1631 );
    xnor g31129 ( n39406 , n6625 , n17297 );
    or g31130 ( n35543 , n1507 , n42779 );
    xnor g31131 ( n21366 , n11051 , n9357 );
    and g31132 ( n18353 , n11228 , n8377 );
    and g31133 ( n27941 , n8260 , n27655 );
    and g31134 ( n971 , n7881 , n11634 );
    or g31135 ( n38915 , n1995 , n11631 );
    xnor g31136 ( n8428 , n35727 , n31049 );
    and g31137 ( n19898 , n14135 , n31063 );
    or g31138 ( n39868 , n7511 , n14238 );
    or g31139 ( n25761 , n9724 , n37890 );
    or g31140 ( n33244 , n15429 , n31458 );
    or g31141 ( n16329 , n29135 , n10647 );
    or g31142 ( n24285 , n38152 , n33849 );
    and g31143 ( n15746 , n28466 , n37431 );
    or g31144 ( n38415 , n19221 , n26250 );
    or g31145 ( n16506 , n10213 , n11284 );
    or g31146 ( n29102 , n26417 , n19205 );
    xnor g31147 ( n15237 , n21957 , n15192 );
    and g31148 ( n30786 , n33180 , n31670 );
    nor g31149 ( n84 , n29414 , n5123 );
    or g31150 ( n32039 , n9470 , n41007 );
    and g31151 ( n674 , n26123 , n21443 );
    xnor g31152 ( n22136 , n18874 , n19170 );
    or g31153 ( n10318 , n2586 , n28598 );
    nor g31154 ( n9892 , n10143 , n40945 );
    or g31155 ( n25397 , n24612 , n39491 );
    and g31156 ( n11824 , n105 , n25585 );
    not g31157 ( n24064 , n24023 );
    and g31158 ( n28576 , n20786 , n9978 );
    or g31159 ( n35794 , n42693 , n35707 );
    nor g31160 ( n41869 , n17724 , n3291 );
    nor g31161 ( n37572 , n13444 , n21994 );
    nor g31162 ( n42344 , n1153 , n40539 );
    or g31163 ( n7224 , n35138 , n26008 );
    not g31164 ( n17814 , n18246 );
    or g31165 ( n5809 , n7040 , n14955 );
    or g31166 ( n7456 , n40703 , n12729 );
    not g31167 ( n3812 , n40297 );
    and g31168 ( n37484 , n35580 , n32192 );
    and g31169 ( n31575 , n34049 , n6609 );
    not g31170 ( n42556 , n11667 );
    not g31171 ( n38256 , n13106 );
    or g31172 ( n9705 , n37552 , n30681 );
    and g31173 ( n13582 , n5034 , n29032 );
    or g31174 ( n9578 , n20821 , n40554 );
    or g31175 ( n9186 , n21341 , n29930 );
    and g31176 ( n9798 , n40288 , n18658 );
    or g31177 ( n35643 , n1647 , n14622 );
    or g31178 ( n35723 , n14822 , n18162 );
    or g31179 ( n38539 , n29027 , n4132 );
    and g31180 ( n35679 , n26180 , n12473 );
    or g31181 ( n3691 , n34584 , n29994 );
    and g31182 ( n29071 , n24029 , n13171 );
    and g31183 ( n17398 , n38353 , n6591 );
    or g31184 ( n28811 , n39934 , n10163 );
    or g31185 ( n4809 , n4258 , n32446 );
    and g31186 ( n39331 , n3760 , n41512 );
    or g31187 ( n11110 , n32181 , n27683 );
    or g31188 ( n30557 , n34927 , n3751 );
    or g31189 ( n5664 , n10168 , n20383 );
    not g31190 ( n3571 , n34880 );
    nor g31191 ( n4379 , n40974 , n8995 );
    nor g31192 ( n16195 , n17272 , n980 );
    or g31193 ( n4048 , n27271 , n33537 );
    not g31194 ( n13868 , n11559 );
    xnor g31195 ( n308 , n36212 , n16015 );
    or g31196 ( n30541 , n41752 , n42211 );
    xnor g31197 ( n20708 , n35727 , n13446 );
    and g31198 ( n9894 , n6071 , n9098 );
    or g31199 ( n25197 , n3192 , n25451 );
    not g31200 ( n35314 , n40505 );
    and g31201 ( n31399 , n6846 , n35988 );
    and g31202 ( n14448 , n8905 , n36339 );
    or g31203 ( n33897 , n25236 , n33640 );
    and g31204 ( n20626 , n34964 , n31646 );
    and g31205 ( n12228 , n31274 , n28146 );
    or g31206 ( n3412 , n28571 , n5258 );
    and g31207 ( n12598 , n4527 , n198 );
    nor g31208 ( n14952 , n1448 , n29381 );
    or g31209 ( n20988 , n22371 , n25315 );
    xnor g31210 ( n17525 , n8591 , n39786 );
    xnor g31211 ( n17741 , n19052 , n7167 );
    or g31212 ( n19896 , n6431 , n14754 );
    or g31213 ( n7911 , n19029 , n9586 );
    or g31214 ( n7343 , n39689 , n12494 );
    and g31215 ( n22884 , n18980 , n26497 );
    or g31216 ( n16581 , n3583 , n5791 );
    nor g31217 ( n40349 , n5896 , n20004 );
    and g31218 ( n25101 , n40846 , n21669 );
    or g31219 ( n16606 , n26984 , n16216 );
    and g31220 ( n14683 , n5370 , n28868 );
    nor g31221 ( n29492 , n38157 , n12555 );
    or g31222 ( n40018 , n1569 , n2675 );
    or g31223 ( n13675 , n4839 , n31345 );
    or g31224 ( n22806 , n2792 , n4753 );
    nor g31225 ( n33865 , n15668 , n41291 );
    or g31226 ( n22541 , n17815 , n29726 );
    and g31227 ( n30360 , n41563 , n41791 );
    and g31228 ( n35242 , n32650 , n40135 );
    and g31229 ( n33744 , n15947 , n29180 );
    or g31230 ( n30372 , n35850 , n9997 );
    or g31231 ( n30323 , n37671 , n10733 );
    or g31232 ( n7017 , n22409 , n33387 );
    or g31233 ( n1973 , n26785 , n32606 );
    and g31234 ( n26288 , n22936 , n6871 );
    or g31235 ( n29629 , n24626 , n36417 );
    or g31236 ( n17211 , n16149 , n29092 );
    or g31237 ( n6639 , n18212 , n15633 );
    or g31238 ( n10061 , n32447 , n41223 );
    and g31239 ( n36410 , n15413 , n28376 );
    or g31240 ( n23780 , n19084 , n20003 );
    or g31241 ( n35298 , n21611 , n6415 );
    not g31242 ( n7564 , n21197 );
    and g31243 ( n3645 , n42759 , n11552 );
    or g31244 ( n24414 , n33624 , n314 );
    or g31245 ( n13292 , n22751 , n18236 );
    and g31246 ( n6240 , n32462 , n17484 );
    nor g31247 ( n39662 , n3437 , n11093 );
    nor g31248 ( n11180 , n23839 , n6200 );
    or g31249 ( n3107 , n35706 , n1728 );
    or g31250 ( n6350 , n34987 , n9510 );
    not g31251 ( n6440 , n30109 );
    or g31252 ( n2961 , n8455 , n37460 );
    or g31253 ( n12039 , n12166 , n9321 );
    or g31254 ( n13679 , n37389 , n2270 );
    or g31255 ( n4295 , n15064 , n22706 );
    nor g31256 ( n12953 , n4937 , n26478 );
    not g31257 ( n37873 , n19086 );
    not g31258 ( n18796 , n11781 );
    or g31259 ( n3589 , n28643 , n15202 );
    and g31260 ( n2432 , n37620 , n19198 );
    or g31261 ( n21454 , n13204 , n36848 );
    xnor g31262 ( n23371 , n25631 , n11105 );
    not g31263 ( n14279 , n39462 );
    not g31264 ( n25468 , n39966 );
    and g31265 ( n35131 , n27581 , n36353 );
    xnor g31266 ( n32963 , n6547 , n6411 );
    and g31267 ( n12026 , n18530 , n13444 );
    and g31268 ( n930 , n16913 , n3613 );
    or g31269 ( n42156 , n7927 , n13364 );
    or g31270 ( n41790 , n22091 , n16860 );
    xnor g31271 ( n20230 , n1762 , n21442 );
    and g31272 ( n26767 , n25212 , n14005 );
    or g31273 ( n22792 , n13338 , n28034 );
    xnor g31274 ( n17226 , n12146 , n14245 );
    nor g31275 ( n1503 , n37 , n33550 );
    xnor g31276 ( n18641 , n10592 , n30786 );
    nor g31277 ( n15109 , n6761 , n16896 );
    nor g31278 ( n10508 , n21088 , n6512 );
    nor g31279 ( n13477 , n7475 , n34819 );
    or g31280 ( n6977 , n14853 , n3715 );
    not g31281 ( n7836 , n5940 );
    or g31282 ( n30177 , n8219 , n31038 );
    nor g31283 ( n13724 , n25775 , n18441 );
    or g31284 ( n35205 , n15889 , n1692 );
    or g31285 ( n5965 , n18798 , n35673 );
    or g31286 ( n36180 , n28135 , n22609 );
    and g31287 ( n3026 , n15634 , n23018 );
    or g31288 ( n40047 , n5124 , n41750 );
    and g31289 ( n37774 , n2347 , n11209 );
    or g31290 ( n12271 , n16605 , n31012 );
    nor g31291 ( n18723 , n35105 , n31073 );
    or g31292 ( n33608 , n34413 , n32820 );
    not g31293 ( n15096 , n3264 );
    not g31294 ( n22161 , n36776 );
    not g31295 ( n16830 , n33795 );
    or g31296 ( n9246 , n40462 , n29522 );
    or g31297 ( n6551 , n17753 , n38258 );
    xnor g31298 ( n9281 , n28612 , n15809 );
    or g31299 ( n15657 , n2708 , n36962 );
    or g31300 ( n8013 , n22659 , n35745 );
    not g31301 ( n26706 , n28755 );
    or g31302 ( n39471 , n25526 , n22696 );
    or g31303 ( n33249 , n28511 , n32392 );
    or g31304 ( n16246 , n26321 , n42907 );
    and g31305 ( n33048 , n36121 , n36310 );
    or g31306 ( n667 , n39677 , n39015 );
    or g31307 ( n5662 , n6560 , n19133 );
    or g31308 ( n1885 , n14471 , n8924 );
    or g31309 ( n6696 , n2213 , n7814 );
    not g31310 ( n14465 , n14375 );
    nor g31311 ( n3444 , n29113 , n21947 );
    or g31312 ( n34211 , n1110 , n23498 );
    xnor g31313 ( n18983 , n40296 , n5472 );
    nor g31314 ( n5629 , n28252 , n2113 );
    and g31315 ( n38447 , n40851 , n9770 );
    xnor g31316 ( n36928 , n18561 , n26007 );
    not g31317 ( n34787 , n25630 );
    and g31318 ( n14854 , n23863 , n10124 );
    and g31319 ( n12721 , n26067 , n25320 );
    nor g31320 ( n18264 , n10833 , n35571 );
    xnor g31321 ( n21339 , n6625 , n29403 );
    not g31322 ( n25233 , n41457 );
    xnor g31323 ( n23886 , n40698 , n28566 );
    nor g31324 ( n4062 , n6257 , n37423 );
    nor g31325 ( n22404 , n31260 , n17089 );
    and g31326 ( n178 , n16399 , n19564 );
    xnor g31327 ( n28841 , n18858 , n284 );
    or g31328 ( n41195 , n22529 , n8421 );
    or g31329 ( n15490 , n42302 , n3728 );
    or g31330 ( n18699 , n29811 , n17448 );
    and g31331 ( n39095 , n20592 , n14912 );
    or g31332 ( n19006 , n33535 , n630 );
    xnor g31333 ( n34268 , n23896 , n34548 );
    and g31334 ( n24793 , n3436 , n31643 );
    nor g31335 ( n2530 , n34698 , n26654 );
    or g31336 ( n20955 , n27039 , n29936 );
    or g31337 ( n13526 , n3693 , n1514 );
    or g31338 ( n19588 , n29487 , n3229 );
    or g31339 ( n6308 , n24294 , n632 );
    or g31340 ( n5902 , n39115 , n1223 );
    nor g31341 ( n7759 , n15118 , n37996 );
    and g31342 ( n33930 , n16531 , n1777 );
    or g31343 ( n42635 , n23201 , n33539 );
    or g31344 ( n14108 , n16586 , n13360 );
    not g31345 ( n29041 , n14120 );
    xnor g31346 ( n39599 , n22054 , n9122 );
    or g31347 ( n36 , n14847 , n29579 );
    not g31348 ( n10681 , n19772 );
    nor g31349 ( n6815 , n18599 , n595 );
    xnor g31350 ( n40236 , n16651 , n18064 );
    and g31351 ( n1269 , n9925 , n13152 );
    or g31352 ( n40542 , n9820 , n11976 );
    or g31353 ( n20768 , n23942 , n35533 );
    or g31354 ( n16813 , n34960 , n13504 );
    nor g31355 ( n24303 , n960 , n11690 );
    or g31356 ( n16259 , n38980 , n41767 );
    or g31357 ( n36736 , n22840 , n25704 );
    nor g31358 ( n21979 , n17561 , n42297 );
    or g31359 ( n36122 , n2608 , n20045 );
    and g31360 ( n26654 , n20839 , n34367 );
    or g31361 ( n8395 , n29927 , n35386 );
    and g31362 ( n42300 , n23861 , n24455 );
    nor g31363 ( n29358 , n20202 , n5684 );
    or g31364 ( n10016 , n29978 , n26927 );
    and g31365 ( n11301 , n40975 , n4030 );
    or g31366 ( n32900 , n26672 , n19476 );
    or g31367 ( n42790 , n19084 , n5764 );
    or g31368 ( n1426 , n18244 , n37225 );
    or g31369 ( n16983 , n36952 , n36320 );
    not g31370 ( n18364 , n11112 );
    and g31371 ( n5893 , n5648 , n7530 );
    and g31372 ( n41015 , n13661 , n27139 );
    or g31373 ( n11742 , n13533 , n37848 );
    or g31374 ( n8364 , n14434 , n11507 );
    not g31375 ( n294 , n13251 );
    or g31376 ( n29753 , n83 , n35852 );
    or g31377 ( n14261 , n13354 , n24506 );
    not g31378 ( n37455 , n42458 );
    nor g31379 ( n4056 , n5896 , n24157 );
    and g31380 ( n15906 , n19846 , n23846 );
    and g31381 ( n30369 , n27077 , n37413 );
    not g31382 ( n18825 , n7401 );
    or g31383 ( n32831 , n14457 , n36540 );
    nor g31384 ( n35384 , n29088 , n11104 );
    and g31385 ( n9539 , n8787 , n26930 );
    or g31386 ( n6903 , n39539 , n34002 );
    or g31387 ( n6412 , n42881 , n4013 );
    or g31388 ( n7444 , n15879 , n21272 );
    nor g31389 ( n42067 , n40401 , n28407 );
    or g31390 ( n27230 , n27594 , n25164 );
    xnor g31391 ( n23773 , n21991 , n4399 );
    nor g31392 ( n36734 , n39025 , n30717 );
    or g31393 ( n16739 , n36815 , n24993 );
    xnor g31394 ( n35261 , n27129 , n5374 );
    and g31395 ( n34284 , n41269 , n9662 );
    and g31396 ( n15084 , n13114 , n7533 );
    nor g31397 ( n19122 , n20115 , n26971 );
    and g31398 ( n345 , n10148 , n39053 );
    not g31399 ( n8904 , n42803 );
    and g31400 ( n31468 , n13358 , n24994 );
    and g31401 ( n23341 , n25869 , n24717 );
    nor g31402 ( n4737 , n3438 , n12160 );
    not g31403 ( n33199 , n22980 );
    or g31404 ( n17616 , n38837 , n10869 );
    and g31405 ( n32432 , n1556 , n41936 );
    xnor g31406 ( n2724 , n16693 , n37564 );
    or g31407 ( n16360 , n24864 , n25959 );
    or g31408 ( n29935 , n14945 , n6515 );
    xnor g31409 ( n7315 , n28548 , n36596 );
    xnor g31410 ( n4917 , n9827 , n41689 );
    or g31411 ( n38272 , n3656 , n11978 );
    nor g31412 ( n33567 , n20685 , n37541 );
    xnor g31413 ( n25697 , n2488 , n38530 );
    or g31414 ( n18959 , n26927 , n21607 );
    and g31415 ( n29587 , n30656 , n613 );
    or g31416 ( n29680 , n16598 , n20721 );
    and g31417 ( n11405 , n32039 , n31398 );
    or g31418 ( n5645 , n10248 , n10496 );
    nor g31419 ( n42453 , n26649 , n5659 );
    or g31420 ( n14473 , n34486 , n12050 );
    and g31421 ( n39260 , n34354 , n28687 );
    and g31422 ( n41590 , n39386 , n15870 );
    and g31423 ( n4021 , n36683 , n36268 );
    nor g31424 ( n12880 , n14471 , n33337 );
    not g31425 ( n28202 , n32831 );
    and g31426 ( n28139 , n26327 , n8370 );
    not g31427 ( n8075 , n42347 );
    xnor g31428 ( n42638 , n34426 , n31197 );
    and g31429 ( n9474 , n16604 , n29793 );
    or g31430 ( n31236 , n9145 , n14623 );
    or g31431 ( n28589 , n4192 , n5110 );
    or g31432 ( n4813 , n32800 , n29510 );
    and g31433 ( n8254 , n5710 , n23768 );
    and g31434 ( n23203 , n4722 , n2969 );
    xnor g31435 ( n17925 , n27093 , n4957 );
    not g31436 ( n13832 , n4873 );
    not g31437 ( n527 , n9331 );
    xnor g31438 ( n36451 , n7004 , n12840 );
    not g31439 ( n30530 , n17617 );
    not g31440 ( n34609 , n24747 );
    or g31441 ( n31104 , n36747 , n27069 );
    or g31442 ( n6906 , n6370 , n11125 );
    nor g31443 ( n6326 , n32793 , n23444 );
    or g31444 ( n854 , n11181 , n25665 );
    or g31445 ( n15291 , n1432 , n22566 );
    or g31446 ( n29114 , n15064 , n15190 );
    or g31447 ( n21728 , n39962 , n16319 );
    xnor g31448 ( n33971 , n11531 , n30186 );
    or g31449 ( n13377 , n34373 , n30186 );
    or g31450 ( n14031 , n1917 , n36535 );
    or g31451 ( n17495 , n40323 , n27482 );
    and g31452 ( n22610 , n42298 , n12151 );
    or g31453 ( n18781 , n16997 , n729 );
    xnor g31454 ( n38295 , n12146 , n14142 );
    or g31455 ( n37797 , n5493 , n23366 );
    xnor g31456 ( n28573 , n17299 , n38088 );
    or g31457 ( n982 , n39768 , n29141 );
    nor g31458 ( n14579 , n14338 , n28848 );
    or g31459 ( n21053 , n31108 , n23936 );
    and g31460 ( n12802 , n38091 , n14495 );
    or g31461 ( n3184 , n15208 , n18102 );
    and g31462 ( n22157 , n40654 , n1147 );
    or g31463 ( n2518 , n33643 , n14694 );
    not g31464 ( n14112 , n3264 );
    or g31465 ( n42291 , n18404 , n33686 );
    or g31466 ( n33959 , n30958 , n32457 );
    or g31467 ( n1624 , n6536 , n33547 );
    and g31468 ( n18366 , n27251 , n4287 );
    or g31469 ( n14911 , n19143 , n15780 );
    or g31470 ( n25832 , n9987 , n18158 );
    not g31471 ( n21503 , n42844 );
    or g31472 ( n28560 , n24417 , n18548 );
    and g31473 ( n18828 , n40233 , n38030 );
    or g31474 ( n13107 , n14225 , n8171 );
    or g31475 ( n13688 , n40462 , n41461 );
    not g31476 ( n18290 , n36315 );
    xnor g31477 ( n37322 , n34731 , n161 );
    and g31478 ( n16911 , n41368 , n32083 );
    or g31479 ( n11850 , n20899 , n21023 );
    or g31480 ( n23260 , n39024 , n38358 );
    xnor g31481 ( n24056 , n30742 , n41539 );
    nor g31482 ( n14179 , n6147 , n19966 );
    xnor g31483 ( n4427 , n8928 , n38238 );
    or g31484 ( n6248 , n18771 , n11246 );
    or g31485 ( n16723 , n2036 , n5117 );
    or g31486 ( n25980 , n37439 , n27028 );
    not g31487 ( n24846 , n32526 );
    xnor g31488 ( n2230 , n32212 , n38993 );
    nor g31489 ( n1393 , n14515 , n555 );
    or g31490 ( n18307 , n23653 , n2658 );
    not g31491 ( n32573 , n39870 );
    and g31492 ( n21460 , n10483 , n31585 );
    xnor g31493 ( n8282 , n105 , n519 );
    xnor g31494 ( n11356 , n7621 , n30212 );
    or g31495 ( n37508 , n38054 , n19590 );
    xnor g31496 ( n41791 , n31099 , n13199 );
    not g31497 ( n31313 , n17593 );
    and g31498 ( n23641 , n5755 , n25864 );
    not g31499 ( n900 , n23507 );
    and g31500 ( n27305 , n34142 , n34630 );
    not g31501 ( n32079 , n6519 );
    or g31502 ( n36808 , n8067 , n17535 );
    nor g31503 ( n23928 , n22109 , n4368 );
    xnor g31504 ( n27093 , n15972 , n40643 );
    or g31505 ( n23156 , n11476 , n895 );
    not g31506 ( n16664 , n40496 );
    nor g31507 ( n23576 , n5964 , n28731 );
    not g31508 ( n32624 , n23681 );
    and g31509 ( n16594 , n34836 , n18573 );
    nor g31510 ( n22469 , n34936 , n10185 );
    not g31511 ( n26202 , n34229 );
    or g31512 ( n15061 , n11838 , n14805 );
    not g31513 ( n21284 , n42854 );
    or g31514 ( n2126 , n18330 , n25010 );
    and g31515 ( n32673 , n19203 , n30363 );
    or g31516 ( n10877 , n38147 , n12322 );
    xnor g31517 ( n24282 , n19501 , n6222 );
    nor g31518 ( n22188 , n10448 , n25357 );
    nor g31519 ( n7096 , n40866 , n14627 );
    or g31520 ( n26316 , n2489 , n7616 );
    and g31521 ( n30462 , n15842 , n14367 );
    xnor g31522 ( n42104 , n842 , n448 );
    nor g31523 ( n13585 , n16691 , n13995 );
    not g31524 ( n26476 , n37046 );
    nor g31525 ( n40940 , n38617 , n11781 );
    not g31526 ( n39710 , n34577 );
    or g31527 ( n20029 , n28860 , n27683 );
    or g31528 ( n32287 , n13066 , n27025 );
    or g31529 ( n13443 , n3812 , n30112 );
    or g31530 ( n42617 , n6019 , n13539 );
    or g31531 ( n9106 , n25246 , n15868 );
    and g31532 ( n41940 , n11060 , n27138 );
    and g31533 ( n14025 , n542 , n5301 );
    or g31534 ( n20515 , n40321 , n32980 );
    xnor g31535 ( n2603 , n8255 , n9851 );
    not g31536 ( n26024 , n27247 );
    xnor g31537 ( n32460 , n36539 , n22004 );
    or g31538 ( n33194 , n36344 , n19496 );
    not g31539 ( n32998 , n23348 );
    or g31540 ( n25321 , n25721 , n29580 );
    xnor g31541 ( n38742 , n36009 , n24901 );
    and g31542 ( n14152 , n42064 , n29168 );
    xnor g31543 ( n20170 , n39256 , n16598 );
    or g31544 ( n23240 , n20169 , n32687 );
    not g31545 ( n9673 , n35604 );
    and g31546 ( n3754 , n33779 , n7416 );
    or g31547 ( n20162 , n12700 , n41824 );
    nor g31548 ( n634 , n18759 , n2402 );
    or g31549 ( n18164 , n5782 , n8352 );
    nor g31550 ( n41194 , n20060 , n37082 );
    or g31551 ( n15207 , n22063 , n16214 );
    or g31552 ( n22072 , n22205 , n10129 );
    xnor g31553 ( n41637 , n29285 , n33832 );
    and g31554 ( n34300 , n33634 , n24427 );
    not g31555 ( n3664 , n9641 );
    not g31556 ( n33858 , n33345 );
    or g31557 ( n42329 , n41134 , n37521 );
    or g31558 ( n12897 , n29020 , n41532 );
    and g31559 ( n27611 , n16670 , n30177 );
    or g31560 ( n20624 , n31322 , n550 );
    nor g31561 ( n32796 , n7648 , n26253 );
    and g31562 ( n17167 , n18493 , n16871 );
    xnor g31563 ( n10744 , n31474 , n13170 );
    and g31564 ( n42856 , n38104 , n17779 );
    or g31565 ( n10545 , n19924 , n34338 );
    not g31566 ( n17119 , n26469 );
    nor g31567 ( n245 , n25588 , n7498 );
    nor g31568 ( n30348 , n15070 , n13337 );
    or g31569 ( n24126 , n22554 , n27228 );
    or g31570 ( n33967 , n33289 , n25464 );
    not g31571 ( n21048 , n19928 );
    not g31572 ( n6277 , n36043 );
    nor g31573 ( n35632 , n2199 , n6571 );
    and g31574 ( n18130 , n37260 , n38334 );
    or g31575 ( n29351 , n28775 , n16316 );
    not g31576 ( n15467 , n3759 );
    xnor g31577 ( n24141 , n2317 , n20231 );
    and g31578 ( n23459 , n26337 , n38338 );
    or g31579 ( n27235 , n14408 , n42569 );
    or g31580 ( n37712 , n22091 , n4711 );
    or g31581 ( n24884 , n29980 , n28969 );
    xnor g31582 ( n41450 , n34735 , n31403 );
    not g31583 ( n9997 , n26165 );
    or g31584 ( n26473 , n19084 , n18458 );
    and g31585 ( n21314 , n25497 , n19751 );
    or g31586 ( n10384 , n15470 , n28343 );
    and g31587 ( n5588 , n26255 , n20560 );
    nor g31588 ( n34718 , n29523 , n8923 );
    and g31589 ( n15478 , n22474 , n4958 );
    not g31590 ( n6663 , n9671 );
    nor g31591 ( n30940 , n16649 , n19258 );
    nor g31592 ( n17921 , n15070 , n20215 );
    or g31593 ( n32280 , n25573 , n11203 );
    not g31594 ( n2435 , n42421 );
    not g31595 ( n5684 , n29310 );
    not g31596 ( n24372 , n2093 );
    xnor g31597 ( n27285 , n4302 , n28525 );
    or g31598 ( n34175 , n18711 , n11279 );
    not g31599 ( n31247 , n31094 );
    or g31600 ( n20121 , n15010 , n7732 );
    or g31601 ( n40723 , n29056 , n3548 );
    or g31602 ( n4992 , n8755 , n3882 );
    and g31603 ( n12050 , n5213 , n42359 );
    not g31604 ( n17865 , n10102 );
    or g31605 ( n11810 , n6501 , n29388 );
    not g31606 ( n41990 , n9654 );
    xnor g31607 ( n26428 , n12190 , n9468 );
    or g31608 ( n17028 , n11798 , n3167 );
    and g31609 ( n10329 , n35950 , n7887 );
    or g31610 ( n13092 , n12198 , n38736 );
    and g31611 ( n30802 , n176 , n28145 );
    or g31612 ( n38496 , n1075 , n2993 );
    or g31613 ( n30256 , n12046 , n29884 );
    nor g31614 ( n7900 , n26194 , n31386 );
    or g31615 ( n8515 , n43 , n38855 );
    xnor g31616 ( n14581 , n37708 , n42036 );
    and g31617 ( n25277 , n42063 , n15394 );
    xnor g31618 ( n5892 , n2241 , n4415 );
    or g31619 ( n30960 , n35799 , n41752 );
    nor g31620 ( n1540 , n17087 , n22718 );
    xnor g31621 ( n41864 , n6625 , n14868 );
    and g31622 ( n22419 , n14496 , n2843 );
    and g31623 ( n14939 , n18111 , n18113 );
    or g31624 ( n21685 , n35463 , n23886 );
    or g31625 ( n39484 , n37630 , n11970 );
    and g31626 ( n5541 , n33661 , n15628 );
    nor g31627 ( n22766 , n36117 , n39781 );
    or g31628 ( n26105 , n103 , n8097 );
    or g31629 ( n41531 , n37180 , n34955 );
    or g31630 ( n32231 , n26379 , n35267 );
    or g31631 ( n20447 , n8375 , n8442 );
    or g31632 ( n36966 , n9764 , n31999 );
    or g31633 ( n20264 , n12607 , n34949 );
    nor g31634 ( n42365 , n7782 , n36008 );
    or g31635 ( n21762 , n4515 , n34511 );
    not g31636 ( n17551 , n41788 );
    not g31637 ( n17583 , n17454 );
    and g31638 ( n8908 , n16128 , n37338 );
    or g31639 ( n13931 , n1971 , n6252 );
    nor g31640 ( n12296 , n36034 , n22555 );
    not g31641 ( n17767 , n29188 );
    or g31642 ( n2823 , n7357 , n34793 );
    nor g31643 ( n1924 , n27588 , n39163 );
    nor g31644 ( n986 , n28104 , n4519 );
    and g31645 ( n31444 , n19721 , n4294 );
    or g31646 ( n24711 , n13684 , n33291 );
    xnor g31647 ( n31685 , n15003 , n8375 );
    and g31648 ( n3028 , n21089 , n29830 );
    or g31649 ( n8883 , n24518 , n32726 );
    not g31650 ( n27704 , n246 );
    or g31651 ( n9121 , n16826 , n41052 );
    and g31652 ( n392 , n30148 , n2192 );
    xnor g31653 ( n37876 , n2903 , n33768 );
    or g31654 ( n11680 , n37197 , n26635 );
    not g31655 ( n28982 , n11397 );
    xnor g31656 ( n10510 , n18678 , n7874 );
    and g31657 ( n15244 , n1258 , n32248 );
    nor g31658 ( n28772 , n20817 , n23127 );
    xnor g31659 ( n12786 , n31542 , n35787 );
    nor g31660 ( n28854 , n23731 , n41164 );
    or g31661 ( n16855 , n19866 , n10028 );
    xnor g31662 ( n7591 , n562 , n41131 );
    nor g31663 ( n19536 , n3769 , n28025 );
    or g31664 ( n17757 , n40512 , n24308 );
    and g31665 ( n21803 , n33906 , n18061 );
    not g31666 ( n31786 , n26415 );
    or g31667 ( n1821 , n750 , n40464 );
    not g31668 ( n31278 , n9215 );
    nor g31669 ( n39383 , n2199 , n17473 );
    xnor g31670 ( n28503 , n21156 , n34035 );
    or g31671 ( n11669 , n3642 , n20030 );
    or g31672 ( n40051 , n10927 , n24295 );
    or g31673 ( n12433 , n24845 , n32752 );
    and g31674 ( n17425 , n38787 , n31933 );
    or g31675 ( n42669 , n31618 , n25444 );
    or g31676 ( n11191 , n37648 , n38149 );
    not g31677 ( n35829 , n22634 );
    and g31678 ( n42010 , n12398 , n41123 );
    and g31679 ( n39461 , n25905 , n3547 );
    and g31680 ( n20521 , n25124 , n3394 );
    and g31681 ( n11825 , n20732 , n16847 );
    and g31682 ( n20199 , n27728 , n2665 );
    and g31683 ( n2587 , n33991 , n35054 );
    not g31684 ( n20345 , n24687 );
    not g31685 ( n14074 , n9814 );
    not g31686 ( n28036 , n3794 );
    not g31687 ( n29115 , n33548 );
    and g31688 ( n40845 , n18220 , n37736 );
    or g31689 ( n1625 , n14234 , n5978 );
    or g31690 ( n9289 , n8031 , n9291 );
    and g31691 ( n34132 , n12517 , n32816 );
    nor g31692 ( n8444 , n12305 , n9626 );
    and g31693 ( n29708 , n15344 , n24935 );
    nor g31694 ( n38595 , n42679 , n15824 );
    nor g31695 ( n28418 , n21366 , n1598 );
    or g31696 ( n29867 , n17796 , n25975 );
    nor g31697 ( n5318 , n17201 , n5383 );
    nor g31698 ( n18398 , n42250 , n38726 );
    or g31699 ( n20863 , n550 , n1203 );
    or g31700 ( n9266 , n15423 , n30169 );
    not g31701 ( n354 , n13805 );
    not g31702 ( n10275 , n29196 );
    and g31703 ( n14601 , n28346 , n41725 );
    nor g31704 ( n25276 , n25230 , n27115 );
    or g31705 ( n1146 , n9961 , n33700 );
    and g31706 ( n37901 , n36803 , n42136 );
    xnor g31707 ( n22381 , n22787 , n13672 );
    or g31708 ( n13678 , n34905 , n30953 );
    and g31709 ( n29183 , n9394 , n13402 );
    nor g31710 ( n19138 , n33981 , n1070 );
    not g31711 ( n11453 , n4141 );
    or g31712 ( n25869 , n32534 , n21777 );
    or g31713 ( n4494 , n13974 , n5310 );
    xnor g31714 ( n10924 , n11436 , n17291 );
    xnor g31715 ( n24428 , n17377 , n18412 );
    or g31716 ( n40019 , n25254 , n33464 );
    or g31717 ( n21600 , n39149 , n2149 );
    and g31718 ( n264 , n11213 , n6854 );
    or g31719 ( n167 , n21720 , n1149 );
    or g31720 ( n18038 , n17193 , n35163 );
    nor g31721 ( n10129 , n18799 , n19598 );
    or g31722 ( n7006 , n1077 , n10645 );
    or g31723 ( n9132 , n39266 , n9550 );
    and g31724 ( n29508 , n28603 , n1912 );
    not g31725 ( n3462 , n9051 );
    not g31726 ( n22170 , n37776 );
    or g31727 ( n12420 , n27682 , n27589 );
    xnor g31728 ( n29017 , n36394 , n22896 );
    or g31729 ( n3953 , n4717 , n36571 );
    not g31730 ( n31480 , n34918 );
    or g31731 ( n9603 , n30896 , n3587 );
    or g31732 ( n40794 , n14494 , n29322 );
    nor g31733 ( n32671 , n34358 , n19110 );
    not g31734 ( n19183 , n27764 );
    not g31735 ( n9829 , n35854 );
    or g31736 ( n39469 , n18287 , n26117 );
    or g31737 ( n31110 , n20010 , n439 );
    nor g31738 ( n36291 , n24420 , n21889 );
    or g31739 ( n14403 , n35890 , n35004 );
    not g31740 ( n31888 , n41140 );
    not g31741 ( n38411 , n7334 );
    not g31742 ( n28650 , n36141 );
    and g31743 ( n5351 , n41161 , n20365 );
    xnor g31744 ( n33069 , n24163 , n33032 );
    xnor g31745 ( n17733 , n26794 , n35629 );
    or g31746 ( n5916 , n8852 , n13486 );
    not g31747 ( n26871 , n34363 );
    and g31748 ( n24581 , n41630 , n22657 );
    not g31749 ( n13006 , n7141 );
    not g31750 ( n31927 , n5345 );
    xnor g31751 ( n6849 , n32297 , n29165 );
    or g31752 ( n6439 , n25547 , n21535 );
    not g31753 ( n38545 , n21197 );
    or g31754 ( n7333 , n20699 , n16927 );
    and g31755 ( n21166 , n39953 , n33277 );
    or g31756 ( n17981 , n13832 , n13783 );
    or g31757 ( n25270 , n13074 , n40286 );
    or g31758 ( n34065 , n10645 , n21854 );
    and g31759 ( n10616 , n5404 , n37649 );
    or g31760 ( n19712 , n40281 , n16357 );
    or g31761 ( n12089 , n29227 , n39578 );
    not g31762 ( n11760 , n19269 );
    nor g31763 ( n2064 , n42558 , n42546 );
    and g31764 ( n4366 , n23702 , n24685 );
    xnor g31765 ( n42822 , n105 , n6006 );
    xnor g31766 ( n12873 , n7282 , n11424 );
    and g31767 ( n23665 , n5018 , n13698 );
    or g31768 ( n3722 , n2199 , n10861 );
    or g31769 ( n28369 , n29300 , n14668 );
    and g31770 ( n3854 , n13173 , n17861 );
    nor g31771 ( n39875 , n41380 , n33561 );
    and g31772 ( n12565 , n35135 , n18187 );
    xnor g31773 ( n23461 , n36046 , n39459 );
    or g31774 ( n33176 , n4430 , n18622 );
    or g31775 ( n18629 , n37763 , n17997 );
    nor g31776 ( n26481 , n33796 , n11834 );
    nor g31777 ( n28741 , n37044 , n5386 );
    not g31778 ( n35394 , n13301 );
    not g31779 ( n35323 , n40748 );
    and g31780 ( n6723 , n31225 , n24269 );
    and g31781 ( n4767 , n38579 , n10550 );
    nor g31782 ( n35350 , n20728 , n42787 );
    or g31783 ( n1361 , n40710 , n26853 );
    not g31784 ( n6692 , n3811 );
    nor g31785 ( n39061 , n3447 , n18742 );
    and g31786 ( n18851 , n2573 , n2301 );
    or g31787 ( n9398 , n7410 , n19756 );
    nor g31788 ( n39830 , n15506 , n5293 );
    nor g31789 ( n37924 , n29313 , n12205 );
    nor g31790 ( n18018 , n19581 , n39840 );
    not g31791 ( n7604 , n33811 );
    or g31792 ( n19939 , n6419 , n7759 );
    xnor g31793 ( n4801 , n40687 , n36287 );
    and g31794 ( n10958 , n33862 , n30501 );
    and g31795 ( n16089 , n1996 , n32378 );
    xnor g31796 ( n33189 , n34731 , n35503 );
    xnor g31797 ( n6727 , n26406 , n38245 );
    or g31798 ( n18741 , n35193 , n5534 );
    and g31799 ( n19303 , n17028 , n16090 );
    and g31800 ( n29316 , n39739 , n6647 );
    nor g31801 ( n11311 , n16952 , n8997 );
    nor g31802 ( n486 , n9664 , n13648 );
    or g31803 ( n36069 , n8816 , n32484 );
    nor g31804 ( n13957 , n33960 , n27154 );
    not g31805 ( n983 , n12088 );
    and g31806 ( n27017 , n27737 , n32211 );
    or g31807 ( n1282 , n25588 , n17706 );
    not g31808 ( n17906 , n33313 );
    not g31809 ( n19435 , n15441 );
    not g31810 ( n35653 , n36012 );
    xnor g31811 ( n37807 , n18880 , n33427 );
    or g31812 ( n5360 , n21697 , n16293 );
    not g31813 ( n27955 , n26994 );
    not g31814 ( n32679 , n36521 );
    not g31815 ( n30685 , n29715 );
    or g31816 ( n14815 , n27637 , n16930 );
    not g31817 ( n26214 , n5098 );
    and g31818 ( n15399 , n37285 , n16288 );
    nor g31819 ( n40769 , n36112 , n41361 );
    or g31820 ( n40198 , n3677 , n5728 );
    and g31821 ( n19142 , n19315 , n23197 );
    and g31822 ( n28269 , n21997 , n12078 );
    not g31823 ( n21972 , n23849 );
    nor g31824 ( n3876 , n10416 , n39816 );
    or g31825 ( n2187 , n3034 , n1819 );
    nor g31826 ( n27553 , n20186 , n20230 );
    nor g31827 ( n18368 , n4447 , n37093 );
    or g31828 ( n32440 , n36422 , n14122 );
    or g31829 ( n7287 , n14481 , n27249 );
    and g31830 ( n29402 , n38357 , n5002 );
    or g31831 ( n6045 , n9616 , n41877 );
    or g31832 ( n34935 , n22135 , n12863 );
    and g31833 ( n20018 , n28877 , n30484 );
    or g31834 ( n37602 , n3487 , n27403 );
    or g31835 ( n41911 , n23292 , n11821 );
    not g31836 ( n4546 , n31694 );
    or g31837 ( n5724 , n7232 , n18826 );
    or g31838 ( n28096 , n32477 , n22201 );
    not g31839 ( n7716 , n27299 );
    xnor g31840 ( n35102 , n10639 , n41385 );
    or g31841 ( n23622 , n29459 , n25001 );
    xnor g31842 ( n15613 , n38749 , n20746 );
    xnor g31843 ( n42873 , n14631 , n37132 );
    or g31844 ( n39620 , n14019 , n3122 );
    or g31845 ( n31853 , n23445 , n37628 );
    not g31846 ( n23610 , n32448 );
    or g31847 ( n10734 , n10756 , n13018 );
    xnor g31848 ( n37607 , n19700 , n33709 );
    or g31849 ( n18446 , n38879 , n25694 );
    not g31850 ( n16603 , n14759 );
    not g31851 ( n39262 , n11948 );
    and g31852 ( n17468 , n4673 , n22793 );
    not g31853 ( n22415 , n28577 );
    not g31854 ( n19767 , n41283 );
    or g31855 ( n628 , n19345 , n31475 );
    or g31856 ( n32401 , n20049 , n7864 );
    or g31857 ( n14528 , n24077 , n17925 );
    and g31858 ( n9837 , n23190 , n39965 );
    xnor g31859 ( n7347 , n26000 , n19221 );
    not g31860 ( n30166 , n3539 );
    or g31861 ( n18280 , n24782 , n4271 );
    or g31862 ( n3324 , n17495 , n19140 );
    and g31863 ( n9182 , n22062 , n21315 );
    and g31864 ( n5960 , n31504 , n17413 );
    and g31865 ( n20102 , n11367 , n25572 );
    xnor g31866 ( n25070 , n37437 , n39984 );
    or g31867 ( n22451 , n14702 , n21 );
    not g31868 ( n42340 , n14954 );
    and g31869 ( n15062 , n15031 , n19904 );
    and g31870 ( n22040 , n28612 , n42297 );
    nor g31871 ( n28695 , n14393 , n9359 );
    or g31872 ( n24550 , n3785 , n14958 );
    and g31873 ( n12647 , n14719 , n30341 );
    nor g31874 ( n3504 , n14471 , n15922 );
    not g31875 ( n32867 , n29953 );
    or g31876 ( n284 , n30591 , n10212 );
    or g31877 ( n30712 , n31265 , n19270 );
    not g31878 ( n22426 , n8573 );
    and g31879 ( n42547 , n764 , n27125 );
    and g31880 ( n31111 , n4459 , n28224 );
    not g31881 ( n36904 , n16579 );
    or g31882 ( n2048 , n17262 , n10398 );
    or g31883 ( n40589 , n38266 , n4675 );
    not g31884 ( n550 , n15196 );
    or g31885 ( n29272 , n23922 , n32894 );
    or g31886 ( n41085 , n13985 , n34195 );
    or g31887 ( n30952 , n5450 , n11183 );
    not g31888 ( n5096 , n5406 );
    and g31889 ( n1837 , n6466 , n42410 );
    not g31890 ( n966 , n18212 );
    or g31891 ( n8208 , n4543 , n1069 );
    nor g31892 ( n11091 , n21022 , n9698 );
    and g31893 ( n336 , n4472 , n40796 );
    xnor g31894 ( n31013 , n41218 , n12592 );
    xnor g31895 ( n11654 , n3713 , n6039 );
    xnor g31896 ( n8578 , n29858 , n27699 );
    nor g31897 ( n20405 , n32651 , n17333 );
    and g31898 ( n7283 , n34700 , n18355 );
    nor g31899 ( n37171 , n2199 , n6703 );
    xnor g31900 ( n34282 , n31848 , n1934 );
    and g31901 ( n9428 , n33703 , n18331 );
    not g31902 ( n1630 , n26233 );
    or g31903 ( n33856 , n36016 , n12504 );
    or g31904 ( n5561 , n13237 , n9884 );
    or g31905 ( n14752 , n26357 , n37912 );
    not g31906 ( n26401 , n21208 );
    and g31907 ( n32873 , n31754 , n10049 );
    not g31908 ( n5441 , n21710 );
    nor g31909 ( n30850 , n40862 , n40918 );
    or g31910 ( n18695 , n39790 , n491 );
    or g31911 ( n13869 , n39988 , n39098 );
    or g31912 ( n7486 , n6370 , n13562 );
    or g31913 ( n30038 , n21893 , n24416 );
    or g31914 ( n1170 , n41920 , n2268 );
    or g31915 ( n10196 , n23623 , n31357 );
    or g31916 ( n10312 , n21814 , n22355 );
    and g31917 ( n22816 , n7182 , n14397 );
    xnor g31918 ( n38128 , n33416 , n27711 );
    nor g31919 ( n26625 , n18417 , n12671 );
    or g31920 ( n2377 , n31440 , n18381 );
    or g31921 ( n29761 , n27738 , n25792 );
    and g31922 ( n25774 , n38911 , n35618 );
    or g31923 ( n4289 , n1657 , n1231 );
    and g31924 ( n12199 , n14476 , n11365 );
    or g31925 ( n2141 , n36238 , n38276 );
    xnor g31926 ( n4284 , n40191 , n19005 );
    xnor g31927 ( n26492 , n2897 , n34565 );
    or g31928 ( n18547 , n1980 , n13601 );
    or g31929 ( n40791 , n1735 , n15690 );
    or g31930 ( n5414 , n9264 , n6592 );
    not g31931 ( n36844 , n29429 );
    or g31932 ( n33833 , n23444 , n7764 );
    or g31933 ( n1150 , n9901 , n8442 );
    or g31934 ( n32158 , n24267 , n21803 );
    not g31935 ( n23374 , n32727 );
    xnor g31936 ( n30315 , n29740 , n10958 );
    xnor g31937 ( n16396 , n42725 , n3632 );
    nor g31938 ( n5467 , n34651 , n16832 );
    or g31939 ( n7799 , n10536 , n11164 );
    or g31940 ( n10589 , n20141 , n6371 );
    and g31941 ( n7867 , n26182 , n6420 );
    and g31942 ( n34523 , n2898 , n26320 );
    or g31943 ( n19951 , n24402 , n14366 );
    or g31944 ( n23212 , n13782 , n29549 );
    nor g31945 ( n36367 , n21733 , n6757 );
    and g31946 ( n17340 , n28704 , n26679 );
    xnor g31947 ( n18907 , n21448 , n17611 );
    or g31948 ( n38635 , n14465 , n33481 );
    xnor g31949 ( n13345 , n21534 , n33630 );
    not g31950 ( n25471 , n41512 );
    not g31951 ( n23431 , n2135 );
    or g31952 ( n32182 , n20288 , n9863 );
    and g31953 ( n9381 , n14371 , n11169 );
    or g31954 ( n4976 , n31914 , n34267 );
    or g31955 ( n32927 , n4660 , n12574 );
    or g31956 ( n28506 , n8042 , n2701 );
    nor g31957 ( n3217 , n29844 , n26549 );
    not g31958 ( n3625 , n19121 );
    and g31959 ( n4132 , n5590 , n41434 );
    or g31960 ( n21081 , n17656 , n37626 );
    not g31961 ( n18954 , n19667 );
    and g31962 ( n10048 , n16474 , n10830 );
    xnor g31963 ( n16191 , n38774 , n16522 );
    nor g31964 ( n37288 , n40156 , n39562 );
    nor g31965 ( n17446 , n8494 , n38039 );
    or g31966 ( n30484 , n25526 , n10170 );
    not g31967 ( n20120 , n7100 );
    or g31968 ( n34612 , n7321 , n11433 );
    and g31969 ( n7053 , n9380 , n10140 );
    nor g31970 ( n34138 , n8434 , n30622 );
    nor g31971 ( n35914 , n15289 , n22666 );
    or g31972 ( n28815 , n23807 , n23261 );
    or g31973 ( n12996 , n36251 , n29779 );
    not g31974 ( n40868 , n1828 );
    and g31975 ( n576 , n18856 , n38159 );
    not g31976 ( n12519 , n7316 );
    not g31977 ( n14096 , n28347 );
    and g31978 ( n6310 , n3206 , n38286 );
    or g31979 ( n33732 , n22388 , n30842 );
    and g31980 ( n5794 , n34793 , n41471 );
    or g31981 ( n4930 , n34796 , n8536 );
    and g31982 ( n15998 , n11670 , n6004 );
    or g31983 ( n11313 , n6762 , n31218 );
    and g31984 ( n40623 , n26898 , n12462 );
    not g31985 ( n4784 , n12367 );
    xnor g31986 ( n15896 , n13296 , n13469 );
    not g31987 ( n35189 , n12135 );
    and g31988 ( n8430 , n31180 , n1376 );
    or g31989 ( n19748 , n35301 , n17193 );
    xnor g31990 ( n5146 , n33416 , n19133 );
    or g31991 ( n14512 , n3487 , n27259 );
    not g31992 ( n5781 , n28023 );
    or g31993 ( n1028 , n6632 , n781 );
    and g31994 ( n17135 , n27564 , n18821 );
    and g31995 ( n11714 , n14382 , n39091 );
    or g31996 ( n18386 , n29495 , n37981 );
    not g31997 ( n6529 , n1303 );
    not g31998 ( n30554 , n23711 );
    and g31999 ( n1358 , n22060 , n26441 );
    nor g32000 ( n35717 , n27905 , n1602 );
    not g32001 ( n40703 , n23184 );
    or g32002 ( n39658 , n34400 , n30704 );
    or g32003 ( n18894 , n29480 , n10094 );
    not g32004 ( n4091 , n17736 );
    and g32005 ( n9122 , n4204 , n33723 );
    nor g32006 ( n30309 , n291 , n2257 );
    xnor g32007 ( n4411 , n5275 , n40214 );
    or g32008 ( n32364 , n12059 , n13369 );
    or g32009 ( n42363 , n18157 , n37237 );
    and g32010 ( n30794 , n6755 , n35204 );
    xnor g32011 ( n20126 , n7724 , n3489 );
    nor g32012 ( n15005 , n42258 , n10392 );
    or g32013 ( n38812 , n28555 , n16146 );
    or g32014 ( n20282 , n1155 , n516 );
    or g32015 ( n3376 , n37585 , n19866 );
    xnor g32016 ( n27323 , n35925 , n26614 );
    or g32017 ( n42189 , n21776 , n23566 );
    nor g32018 ( n24288 , n14863 , n24715 );
    and g32019 ( n26272 , n41173 , n10641 );
    and g32020 ( n14856 , n32927 , n16760 );
    and g32021 ( n24506 , n33359 , n30077 );
    not g32022 ( n15317 , n19531 );
    and g32023 ( n21574 , n27433 , n36331 );
    and g32024 ( n26791 , n7597 , n19820 );
    not g32025 ( n2407 , n35158 );
    or g32026 ( n18357 , n30358 , n13980 );
    and g32027 ( n21047 , n42198 , n685 );
    and g32028 ( n21691 , n20637 , n24725 );
    not g32029 ( n25343 , n36025 );
    and g32030 ( n16012 , n11013 , n4068 );
    xnor g32031 ( n1291 , n10367 , n24968 );
    nor g32032 ( n24230 , n33187 , n25603 );
    or g32033 ( n34708 , n34569 , n11490 );
    xnor g32034 ( n29201 , n36667 , n32942 );
    and g32035 ( n29608 , n1798 , n27883 );
    not g32036 ( n14125 , n9051 );
    or g32037 ( n42714 , n17086 , n6555 );
    or g32038 ( n40112 , n1456 , n5154 );
    nor g32039 ( n33748 , n3762 , n34706 );
    and g32040 ( n25770 , n14197 , n16528 );
    or g32041 ( n39472 , n38276 , n28500 );
    or g32042 ( n29657 , n42096 , n19812 );
    and g32043 ( n34418 , n676 , n30162 );
    not g32044 ( n11383 , n38661 );
    xnor g32045 ( n42022 , n40 , n5403 );
    or g32046 ( n31560 , n20411 , n28894 );
    or g32047 ( n3687 , n38879 , n1028 );
    and g32048 ( n11264 , n17669 , n5389 );
    not g32049 ( n40191 , n22454 );
    and g32050 ( n28417 , n15162 , n14319 );
    xnor g32051 ( n27677 , n31989 , n29097 );
    or g32052 ( n15367 , n33115 , n18502 );
    or g32053 ( n30396 , n21260 , n20169 );
    or g32054 ( n15710 , n9024 , n23954 );
    not g32055 ( n23425 , n30608 );
    and g32056 ( n14590 , n36656 , n31980 );
    not g32057 ( n24496 , n14454 );
    nor g32058 ( n18183 , n785 , n15448 );
    or g32059 ( n15824 , n38014 , n3020 );
    or g32060 ( n30452 , n42753 , n27385 );
    nor g32061 ( n38613 , n30058 , n7722 );
    or g32062 ( n1547 , n13830 , n30312 );
    or g32063 ( n36144 , n36848 , n17973 );
    or g32064 ( n26371 , n38945 , n42520 );
    or g32065 ( n38875 , n29058 , n32580 );
    nor g32066 ( n35714 , n29784 , n9940 );
    and g32067 ( n28817 , n22301 , n3202 );
    and g32068 ( n7417 , n17745 , n19875 );
    or g32069 ( n29769 , n26533 , n7663 );
    xnor g32070 ( n12523 , n19577 , n13822 );
    xnor g32071 ( n40256 , n24190 , n10598 );
    or g32072 ( n37433 , n11629 , n7675 );
    nor g32073 ( n7500 , n35195 , n22982 );
    not g32074 ( n31989 , n18866 );
    or g32075 ( n20549 , n41290 , n41147 );
    and g32076 ( n1352 , n36006 , n18401 );
    xnor g32077 ( n10686 , n36009 , n13582 );
    not g32078 ( n32895 , n31318 );
    and g32079 ( n23604 , n37125 , n30476 );
    or g32080 ( n25059 , n12700 , n9860 );
    and g32081 ( n13044 , n3958 , n28354 );
    not g32082 ( n28617 , n34414 );
    and g32083 ( n27671 , n32177 , n15833 );
    xnor g32084 ( n15330 , n9250 , n33954 );
    or g32085 ( n5834 , n1329 , n8506 );
    nor g32086 ( n12430 , n37335 , n18050 );
    and g32087 ( n39731 , n13177 , n21672 );
    xnor g32088 ( n34489 , n21555 , n41534 );
    and g32089 ( n2366 , n13519 , n23075 );
    xnor g32090 ( n26232 , n19385 , n9703 );
    or g32091 ( n12518 , n33838 , n5997 );
    or g32092 ( n17662 , n22597 , n11695 );
    nor g32093 ( n26917 , n6663 , n32430 );
    and g32094 ( n14721 , n24306 , n23628 );
    xnor g32095 ( n14595 , n22874 , n41362 );
    not g32096 ( n42794 , n36754 );
    or g32097 ( n2106 , n4366 , n24108 );
    nor g32098 ( n20495 , n20086 , n27275 );
    or g32099 ( n21578 , n31905 , n36203 );
    or g32100 ( n8349 , n21563 , n30071 );
    or g32101 ( n42685 , n31751 , n24053 );
    or g32102 ( n31241 , n13222 , n42021 );
    or g32103 ( n28790 , n38120 , n29930 );
    nor g32104 ( n6751 , n11032 , n5051 );
    nor g32105 ( n31004 , n6457 , n40525 );
    and g32106 ( n41159 , n39094 , n32738 );
    xnor g32107 ( n16432 , n1622 , n42620 );
    xnor g32108 ( n17050 , n26996 , n10626 );
    or g32109 ( n39907 , n30499 , n19590 );
    or g32110 ( n2376 , n15014 , n31634 );
    not g32111 ( n32042 , n36137 );
    nor g32112 ( n19968 , n3558 , n21019 );
    and g32113 ( n23774 , n6644 , n8801 );
    and g32114 ( n29258 , n16829 , n14517 );
    or g32115 ( n34839 , n9009 , n25033 );
    or g32116 ( n12951 , n2213 , n8479 );
    or g32117 ( n5804 , n42604 , n4185 );
    or g32118 ( n23291 , n17810 , n313 );
    xnor g32119 ( n37794 , n527 , n31902 );
    and g32120 ( n9406 , n1770 , n34599 );
    or g32121 ( n7906 , n16996 , n13285 );
    and g32122 ( n7340 , n17051 , n16775 );
    or g32123 ( n14444 , n2412 , n34695 );
    or g32124 ( n16697 , n29782 , n36832 );
    or g32125 ( n35583 , n40607 , n23760 );
    and g32126 ( n19786 , n23219 , n32838 );
    and g32127 ( n6676 , n38801 , n36421 );
    xnor g32128 ( n7712 , n6634 , n17213 );
    or g32129 ( n25156 , n19639 , n13258 );
    or g32130 ( n14191 , n22673 , n8409 );
    xnor g32131 ( n5708 , n25552 , n30199 );
    or g32132 ( n4377 , n6048 , n12129 );
    nor g32133 ( n17550 , n24393 , n24834 );
    and g32134 ( n26924 , n33831 , n14191 );
    not g32135 ( n1051 , n16308 );
    and g32136 ( n9399 , n24101 , n8365 );
    or g32137 ( n38244 , n38604 , n4786 );
    and g32138 ( n1908 , n31273 , n38716 );
    nor g32139 ( n25346 , n1507 , n25116 );
    not g32140 ( n4861 , n38298 );
    and g32141 ( n3514 , n27993 , n38979 );
    xnor g32142 ( n16548 , n18529 , n25235 );
    xnor g32143 ( n33028 , n898 , n9928 );
    or g32144 ( n37918 , n34686 , n42489 );
    not g32145 ( n23963 , n4206 );
    and g32146 ( n6550 , n33282 , n35507 );
    and g32147 ( n35952 , n32806 , n13461 );
    not g32148 ( n34253 , n4060 );
    nor g32149 ( n14657 , n42142 , n12089 );
    or g32150 ( n32881 , n21995 , n38423 );
    not g32151 ( n28241 , n23365 );
    or g32152 ( n21200 , n17013 , n3196 );
    or g32153 ( n1382 , n23880 , n20767 );
    or g32154 ( n41503 , n21531 , n30140 );
    nor g32155 ( n27108 , n9264 , n8707 );
    or g32156 ( n13726 , n22427 , n33472 );
    or g32157 ( n3060 , n3026 , n22722 );
    or g32158 ( n16077 , n14340 , n26637 );
    not g32159 ( n2972 , n25288 );
    not g32160 ( n38992 , n1977 );
    not g32161 ( n15003 , n38486 );
    nor g32162 ( n17826 , n32475 , n15809 );
    nor g32163 ( n5844 , n35974 , n9981 );
    not g32164 ( n17589 , n6038 );
    or g32165 ( n8551 , n2507 , n14804 );
    nor g32166 ( n34006 , n39266 , n3498 );
    or g32167 ( n41408 , n41002 , n36810 );
    nor g32168 ( n31900 , n19221 , n20049 );
    and g32169 ( n20075 , n31064 , n41989 );
    and g32170 ( n27079 , n26496 , n2749 );
    and g32171 ( n38743 , n23419 , n28799 );
    and g32172 ( n41201 , n27279 , n6005 );
    xnor g32173 ( n37914 , n15089 , n11645 );
    and g32174 ( n24807 , n3064 , n13463 );
    nor g32175 ( n20027 , n7315 , n4592 );
    or g32176 ( n21505 , n11431 , n814 );
    xnor g32177 ( n21766 , n41013 , n30101 );
    or g32178 ( n11377 , n39106 , n26888 );
    or g32179 ( n12412 , n17120 , n27580 );
    nor g32180 ( n33111 , n25041 , n19233 );
    xnor g32181 ( n9304 , n31048 , n33635 );
    or g32182 ( n33711 , n6414 , n12081 );
    nor g32183 ( n33144 , n26377 , n21319 );
    xnor g32184 ( n10588 , n21332 , n39083 );
    not g32185 ( n31626 , n31510 );
    or g32186 ( n3479 , n21777 , n4660 );
    nor g32187 ( n6158 , n31115 , n35088 );
    or g32188 ( n9149 , n13197 , n24566 );
    or g32189 ( n13990 , n27840 , n36905 );
    or g32190 ( n29386 , n30348 , n22365 );
    or g32191 ( n38655 , n40978 , n15607 );
    or g32192 ( n41803 , n34268 , n39924 );
    and g32193 ( n5790 , n32742 , n42876 );
    or g32194 ( n6031 , n7242 , n13823 );
    not g32195 ( n25222 , n1112 );
    nor g32196 ( n11631 , n20732 , n16847 );
    or g32197 ( n22803 , n4048 , n15989 );
    not g32198 ( n40786 , n16057 );
    nor g32199 ( n2884 , n19054 , n775 );
    or g32200 ( n12635 , n41394 , n28335 );
    or g32201 ( n11167 , n33027 , n79 );
    or g32202 ( n23477 , n42340 , n6411 );
    and g32203 ( n21602 , n14277 , n28952 );
    xnor g32204 ( n35185 , n2127 , n9646 );
    nor g32205 ( n32858 , n13947 , n25957 );
    xnor g32206 ( n30575 , n2183 , n36717 );
    xnor g32207 ( n9551 , n39418 , n24039 );
    not g32208 ( n17667 , n18318 );
    not g32209 ( n22788 , n25255 );
    nor g32210 ( n11593 , n10131 , n9776 );
    or g32211 ( n38459 , n15681 , n20306 );
    xnor g32212 ( n5190 , n19203 , n30363 );
    nor g32213 ( n18221 , n14471 , n37143 );
    and g32214 ( n13475 , n36557 , n26441 );
    or g32215 ( n10487 , n16786 , n42544 );
    and g32216 ( n790 , n30515 , n4917 );
    and g32217 ( n41691 , n40524 , n22015 );
    xnor g32218 ( n38736 , n25428 , n982 );
    not g32219 ( n25709 , n31266 );
    and g32220 ( n38039 , n21418 , n25854 );
    or g32221 ( n9028 , n15696 , n20630 );
    or g32222 ( n37257 , n12757 , n12527 );
    not g32223 ( n39526 , n33171 );
    not g32224 ( n2822 , n31244 );
    and g32225 ( n42817 , n28546 , n30286 );
    xnor g32226 ( n33308 , n35727 , n30511 );
    and g32227 ( n14809 , n450 , n7636 );
    or g32228 ( n31526 , n14471 , n29700 );
    not g32229 ( n4012 , n9604 );
    not g32230 ( n12051 , n22863 );
    or g32231 ( n29946 , n29328 , n38520 );
    or g32232 ( n29124 , n8926 , n15670 );
    not g32233 ( n26641 , n12465 );
    or g32234 ( n34946 , n38777 , n17181 );
    not g32235 ( n3893 , n41847 );
    nor g32236 ( n22064 , n14475 , n4567 );
    or g32237 ( n31057 , n42529 , n24449 );
    or g32238 ( n19886 , n10513 , n7637 );
    not g32239 ( n5531 , n31111 );
    or g32240 ( n4350 , n20546 , n8035 );
    xnor g32241 ( n7997 , n10293 , n10932 );
    or g32242 ( n11985 , n32168 , n12721 );
    or g32243 ( n21035 , n29281 , n12717 );
    nor g32244 ( n31000 , n20487 , n29899 );
    xnor g32245 ( n23373 , n27705 , n35245 );
    nor g32246 ( n31678 , n22173 , n18962 );
    xnor g32247 ( n4686 , n4800 , n40649 );
    and g32248 ( n35165 , n23517 , n8116 );
    xnor g32249 ( n14550 , n41856 , n33527 );
    and g32250 ( n38565 , n19169 , n28123 );
    and g32251 ( n17165 , n2287 , n7241 );
    xnor g32252 ( n33086 , n29034 , n9801 );
    or g32253 ( n32702 , n1997 , n10620 );
    xnor g32254 ( n25388 , n16693 , n17005 );
    not g32255 ( n14146 , n11777 );
    xnor g32256 ( n42211 , n38901 , n8854 );
    or g32257 ( n28972 , n14813 , n15942 );
    xnor g32258 ( n27779 , n26899 , n18820 );
    or g32259 ( n3321 , n36600 , n32835 );
    xnor g32260 ( n17306 , n34040 , n32270 );
    or g32261 ( n38841 , n4306 , n10760 );
    or g32262 ( n29997 , n36780 , n39072 );
    nor g32263 ( n29313 , n40 , n37991 );
    or g32264 ( n37198 , n550 , n37558 );
    or g32265 ( n10187 , n3639 , n40137 );
    not g32266 ( n31271 , n19002 );
    not g32267 ( n22057 , n478 );
    nor g32268 ( n32512 , n7723 , n16748 );
    not g32269 ( n17082 , n25930 );
    and g32270 ( n18328 , n16701 , n15146 );
    or g32271 ( n26611 , n41977 , n2980 );
    or g32272 ( n29168 , n11111 , n24387 );
    and g32273 ( n18482 , n35820 , n11795 );
    or g32274 ( n40093 , n22358 , n6359 );
    or g32275 ( n18262 , n9048 , n20277 );
    and g32276 ( n18228 , n10362 , n22684 );
    or g32277 ( n21621 , n29574 , n13703 );
    and g32278 ( n1738 , n39620 , n40659 );
    or g32279 ( n14116 , n18971 , n38674 );
    and g32280 ( n21665 , n40960 , n15231 );
    or g32281 ( n7403 , n31994 , n32700 );
    or g32282 ( n35128 , n25389 , n38646 );
    or g32283 ( n39414 , n7433 , n29009 );
    or g32284 ( n26383 , n28258 , n30035 );
    and g32285 ( n36511 , n4601 , n37530 );
    or g32286 ( n27971 , n41263 , n18841 );
    or g32287 ( n10303 , n37217 , n26376 );
    or g32288 ( n20493 , n21752 , n39694 );
    and g32289 ( n14170 , n39148 , n9074 );
    or g32290 ( n32417 , n35320 , n18842 );
    nor g32291 ( n897 , n31542 , n33963 );
    nor g32292 ( n15852 , n37577 , n19153 );
    or g32293 ( n18256 , n33665 , n7750 );
    nor g32294 ( n28087 , n36636 , n23233 );
    or g32295 ( n36864 , n38207 , n4552 );
    or g32296 ( n24641 , n27567 , n11321 );
    not g32297 ( n41578 , n21870 );
    nor g32298 ( n42260 , n22112 , n7587 );
    or g32299 ( n8667 , n29857 , n26946 );
    xnor g32300 ( n37248 , n2631 , n22350 );
    xnor g32301 ( n6297 , n12405 , n29828 );
    xnor g32302 ( n15381 , n4796 , n16730 );
    and g32303 ( n7219 , n22632 , n40812 );
    or g32304 ( n35642 , n14903 , n6728 );
    xnor g32305 ( n1133 , n41065 , n6080 );
    and g32306 ( n10925 , n39643 , n633 );
    or g32307 ( n7571 , n1980 , n28624 );
    or g32308 ( n17661 , n5454 , n41574 );
    or g32309 ( n2307 , n29183 , n7767 );
    and g32310 ( n24283 , n20368 , n10034 );
    and g32311 ( n11820 , n15124 , n22682 );
    or g32312 ( n23294 , n26310 , n30316 );
    and g32313 ( n41205 , n37012 , n26543 );
    not g32314 ( n4491 , n928 );
    not g32315 ( n16842 , n31140 );
    not g32316 ( n40710 , n25700 );
    xnor g32317 ( n11497 , n22263 , n23808 );
    xnor g32318 ( n21633 , n31099 , n10506 );
    and g32319 ( n24042 , n32929 , n3440 );
    and g32320 ( n34003 , n5249 , n41708 );
    not g32321 ( n37094 , n30638 );
    and g32322 ( n33904 , n6611 , n2779 );
    not g32323 ( n18138 , n19735 );
    or g32324 ( n41146 , n33981 , n18521 );
    xnor g32325 ( n42521 , n17788 , n5896 );
    or g32326 ( n2550 , n5660 , n34728 );
    or g32327 ( n41059 , n21201 , n10958 );
    and g32328 ( n29605 , n36069 , n9737 );
    xnor g32329 ( n39733 , n38535 , n11293 );
    nor g32330 ( n5683 , n38356 , n38348 );
    and g32331 ( n31509 , n30987 , n27397 );
    xnor g32332 ( n11029 , n12146 , n15080 );
    or g32333 ( n4003 , n16996 , n38658 );
    nor g32334 ( n1454 , n5061 , n11561 );
    not g32335 ( n21476 , n39068 );
    or g32336 ( n27066 , n14129 , n2904 );
    and g32337 ( n787 , n36127 , n32399 );
    and g32338 ( n25230 , n12557 , n12832 );
    and g32339 ( n15569 , n20852 , n19245 );
    nor g32340 ( n35944 , n40441 , n17782 );
    and g32341 ( n22279 , n39648 , n26762 );
    not g32342 ( n7404 , n12725 );
    nor g32343 ( n41035 , n36117 , n17057 );
    or g32344 ( n37387 , n41943 , n15734 );
    or g32345 ( n20871 , n32339 , n37014 );
    or g32346 ( n19776 , n22344 , n33106 );
    and g32347 ( n29228 , n73 , n26109 );
    not g32348 ( n10858 , n30143 );
    xnor g32349 ( n17964 , n4304 , n32798 );
    or g32350 ( n3850 , n37903 , n36663 );
    and g32351 ( n22158 , n40707 , n31280 );
    or g32352 ( n27828 , n6097 , n22819 );
    or g32353 ( n401 , n10473 , n3728 );
    and g32354 ( n9279 , n721 , n22917 );
    not g32355 ( n22954 , n22212 );
    or g32356 ( n22514 , n10844 , n41683 );
    nor g32357 ( n24764 , n40406 , n4054 );
    xnor g32358 ( n2667 , n39077 , n31080 );
    nor g32359 ( n31700 , n30409 , n24947 );
    nor g32360 ( n26793 , n27590 , n26151 );
    or g32361 ( n33242 , n12001 , n27058 );
    not g32362 ( n27782 , n36513 );
    nor g32363 ( n20107 , n16695 , n37563 );
    and g32364 ( n11577 , n34659 , n5691 );
    and g32365 ( n31145 , n21255 , n33424 );
    not g32366 ( n15499 , n10505 );
    and g32367 ( n36644 , n15988 , n19016 );
    or g32368 ( n29600 , n11346 , n4100 );
    or g32369 ( n31757 , n21692 , n21436 );
    or g32370 ( n6516 , n40940 , n30068 );
    and g32371 ( n21898 , n5041 , n12883 );
    or g32372 ( n20584 , n16598 , n23140 );
    xnor g32373 ( n1722 , n15089 , n23604 );
    and g32374 ( n11177 , n20282 , n19970 );
    nor g32375 ( n40122 , n1890 , n34465 );
    or g32376 ( n6873 , n1668 , n13368 );
    nor g32377 ( n13102 , n13769 , n27186 );
    nor g32378 ( n36988 , n2375 , n14119 );
    or g32379 ( n41109 , n16151 , n3234 );
    nor g32380 ( n41726 , n8971 , n29280 );
    xnor g32381 ( n19121 , n30832 , n10172 );
    or g32382 ( n4080 , n9904 , n18100 );
    xnor g32383 ( n24031 , n33678 , n13953 );
    nor g32384 ( n17953 , n29739 , n506 );
    nor g32385 ( n41294 , n14105 , n28629 );
    or g32386 ( n4469 , n9297 , n35634 );
    or g32387 ( n5803 , n34105 , n29477 );
    xnor g32388 ( n4508 , n5246 , n17466 );
    or g32389 ( n34026 , n33680 , n29299 );
    and g32390 ( n39765 , n33219 , n18052 );
    or g32391 ( n38070 , n42755 , n28253 );
    xnor g32392 ( n17372 , n18530 , n21280 );
    nor g32393 ( n18379 , n5413 , n869 );
    nor g32394 ( n22270 , n18176 , n5053 );
    or g32395 ( n26029 , n3703 , n35362 );
    or g32396 ( n29718 , n1638 , n28881 );
    or g32397 ( n7755 , n27319 , n29191 );
    or g32398 ( n21958 , n10066 , n30070 );
    or g32399 ( n23833 , n23394 , n26488 );
    and g32400 ( n9763 , n12977 , n39701 );
    and g32401 ( n31388 , n219 , n37507 );
    xnor g32402 ( n22457 , n19348 , n16752 );
    and g32403 ( n24195 , n3419 , n8349 );
    nor g32404 ( n17608 , n14707 , n23933 );
    or g32405 ( n33148 , n2784 , n29508 );
    nor g32406 ( n14790 , n5938 , n32090 );
    nor g32407 ( n24310 , n10142 , n29356 );
    or g32408 ( n15246 , n20699 , n11816 );
    or g32409 ( n40641 , n8474 , n34841 );
    or g32410 ( n7915 , n31235 , n5281 );
    not g32411 ( n35021 , n16138 );
    xnor g32412 ( n11917 , n31821 , n34538 );
    and g32413 ( n31981 , n11535 , n37550 );
    or g32414 ( n5887 , n21069 , n29058 );
    and g32415 ( n28444 , n17749 , n33004 );
    nor g32416 ( n41244 , n6750 , n10452 );
    or g32417 ( n771 , n40404 , n32922 );
    and g32418 ( n1023 , n26425 , n11089 );
    and g32419 ( n7406 , n34341 , n26029 );
    and g32420 ( n38658 , n37704 , n40806 );
    or g32421 ( n7731 , n4189 , n29614 );
    and g32422 ( n16908 , n14415 , n41276 );
    or g32423 ( n42389 , n13917 , n25732 );
    or g32424 ( n4111 , n4378 , n31925 );
    or g32425 ( n7438 , n36105 , n11979 );
    not g32426 ( n17742 , n22576 );
    not g32427 ( n25377 , n19451 );
    nor g32428 ( n33810 , n17193 , n23808 );
    not g32429 ( n896 , n27134 );
    and g32430 ( n12522 , n476 , n33717 );
    or g32431 ( n9074 , n26542 , n22924 );
    or g32432 ( n37328 , n26927 , n17550 );
    and g32433 ( n33462 , n15603 , n28980 );
    not g32434 ( n22333 , n29731 );
    or g32435 ( n39060 , n1535 , n24044 );
    or g32436 ( n38851 , n19777 , n7616 );
    or g32437 ( n35886 , n28961 , n1100 );
    or g32438 ( n12770 , n3884 , n32029 );
    or g32439 ( n10281 , n27687 , n11574 );
    xnor g32440 ( n33676 , n18521 , n33981 );
    not g32441 ( n11483 , n22987 );
    and g32442 ( n20971 , n14584 , n15297 );
    and g32443 ( n5496 , n4493 , n35620 );
    or g32444 ( n41432 , n21686 , n14348 );
    nor g32445 ( n420 , n17563 , n6073 );
    not g32446 ( n29077 , n13859 );
    and g32447 ( n16189 , n36538 , n25611 );
    and g32448 ( n11411 , n15334 , n26440 );
    or g32449 ( n29529 , n1971 , n12075 );
    or g32450 ( n17781 , n25137 , n24661 );
    not g32451 ( n5841 , n13119 );
    or g32452 ( n20228 , n7916 , n23893 );
    nor g32453 ( n37715 , n35928 , n16234 );
    and g32454 ( n4709 , n21459 , n19494 );
    nor g32455 ( n23519 , n9083 , n21576 );
    or g32456 ( n36281 , n26354 , n16508 );
    and g32457 ( n16610 , n38694 , n29342 );
    or g32458 ( n7253 , n19791 , n33216 );
    or g32459 ( n11212 , n24677 , n38996 );
    and g32460 ( n24611 , n38928 , n13349 );
    xnor g32461 ( n5596 , n13444 , n17500 );
    or g32462 ( n12857 , n13612 , n22784 );
    nor g32463 ( n28311 , n25417 , n36620 );
    or g32464 ( n37442 , n12522 , n33213 );
    xnor g32465 ( n2188 , n24590 , n33936 );
    or g32466 ( n33286 , n9225 , n8840 );
    or g32467 ( n1836 , n36887 , n34882 );
    or g32468 ( n18801 , n22691 , n14806 );
    not g32469 ( n22343 , n22854 );
    or g32470 ( n40453 , n36788 , n6771 );
    not g32471 ( n16896 , n20087 );
    or g32472 ( n22959 , n23778 , n33369 );
    nor g32473 ( n26175 , n6573 , n20118 );
    xnor g32474 ( n21688 , n25041 , n19000 );
    or g32475 ( n32050 , n1192 , n2943 );
    and g32476 ( n32020 , n1755 , n15713 );
    or g32477 ( n14160 , n7795 , n9172 );
    or g32478 ( n40567 , n40612 , n34995 );
    or g32479 ( n11870 , n33954 , n30616 );
    not g32480 ( n18862 , n9182 );
    nor g32481 ( n9032 , n39330 , n20229 );
    and g32482 ( n12621 , n21705 , n21845 );
    xnor g32483 ( n6375 , n42064 , n34423 );
    or g32484 ( n2718 , n11995 , n6265 );
    or g32485 ( n20619 , n32123 , n2647 );
    or g32486 ( n8326 , n3697 , n15507 );
    nor g32487 ( n8685 , n6354 , n22397 );
    or g32488 ( n2974 , n135 , n29291 );
    not g32489 ( n20250 , n42154 );
    or g32490 ( n7387 , n23998 , n22767 );
    or g32491 ( n11075 , n29942 , n2769 );
    or g32492 ( n9214 , n41892 , n24077 );
    not g32493 ( n15423 , n7702 );
    and g32494 ( n5428 , n5129 , n21271 );
    nor g32495 ( n35740 , n31541 , n38475 );
    or g32496 ( n5005 , n40178 , n12341 );
    nor g32497 ( n21848 , n14188 , n34179 );
    or g32498 ( n19022 , n39805 , n6832 );
    not g32499 ( n14901 , n9956 );
    or g32500 ( n5226 , n16586 , n34385 );
    xnor g32501 ( n23243 , n17944 , n17120 );
    not g32502 ( n40995 , n10848 );
    or g32503 ( n9286 , n20086 , n20390 );
    or g32504 ( n13327 , n33102 , n4799 );
    xnor g32505 ( n12501 , n6914 , n18068 );
    nor g32506 ( n32594 , n29698 , n20702 );
    or g32507 ( n17632 , n32673 , n18264 );
    and g32508 ( n12149 , n27613 , n24051 );
    and g32509 ( n23777 , n38671 , n42825 );
    or g32510 ( n6687 , n26939 , n29979 );
    and g32511 ( n20229 , n4863 , n31594 );
    or g32512 ( n16380 , n21388 , n36687 );
    or g32513 ( n34890 , n10839 , n21289 );
    xnor g32514 ( n19063 , n29347 , n2303 );
    and g32515 ( n22489 , n3944 , n7164 );
    or g32516 ( n31670 , n6693 , n35732 );
    xnor g32517 ( n40814 , n28313 , n20759 );
    not g32518 ( n39700 , n8182 );
    or g32519 ( n23544 , n27298 , n9690 );
    or g32520 ( n36608 , n37481 , n35193 );
    and g32521 ( n12260 , n14522 , n20645 );
    and g32522 ( n31322 , n10642 , n27046 );
    or g32523 ( n15559 , n34565 , n34505 );
    or g32524 ( n3921 , n37065 , n25303 );
    or g32525 ( n17806 , n9991 , n42446 );
    nor g32526 ( n27504 , n14471 , n22499 );
    and g32527 ( n26162 , n27212 , n19334 );
    not g32528 ( n35310 , n13042 );
    not g32529 ( n1853 , n41236 );
    and g32530 ( n42490 , n32084 , n26773 );
    not g32531 ( n16430 , n3442 );
    not g32532 ( n30818 , n38991 );
    not g32533 ( n21597 , n21742 );
    or g32534 ( n31695 , n24766 , n27045 );
    nor g32535 ( n27088 , n7467 , n41713 );
    and g32536 ( n41820 , n19018 , n27360 );
    or g32537 ( n12231 , n20522 , n12220 );
    or g32538 ( n1260 , n30748 , n27221 );
    or g32539 ( n29295 , n34260 , n16575 );
    and g32540 ( n40494 , n21940 , n37527 );
    or g32541 ( n16407 , n35516 , n22628 );
    and g32542 ( n11597 , n38161 , n17518 );
    and g32543 ( n23106 , n9686 , n40636 );
    nor g32544 ( n11827 , n13849 , n12750 );
    or g32545 ( n4126 , n9958 , n15661 );
    xnor g32546 ( n19983 , n719 , n6520 );
    xnor g32547 ( n41747 , n29740 , n1738 );
    nor g32548 ( n3935 , n8494 , n10665 );
    nor g32549 ( n1589 , n33674 , n39803 );
    xnor g32550 ( n8718 , n33172 , n9046 );
    and g32551 ( n32093 , n4638 , n16266 );
    or g32552 ( n34462 , n18018 , n39811 );
    nor g32553 ( n4679 , n29781 , n21658 );
    not g32554 ( n23962 , n40934 );
    or g32555 ( n28071 , n27295 , n876 );
    or g32556 ( n25027 , n4397 , n15919 );
    or g32557 ( n497 , n14448 , n37808 );
    nor g32558 ( n12410 , n4102 , n7961 );
    nor g32559 ( n16341 , n18866 , n35518 );
    not g32560 ( n24386 , n33000 );
    nor g32561 ( n11076 , n19155 , n32649 );
    and g32562 ( n11683 , n36045 , n40595 );
    nor g32563 ( n16785 , n30280 , n2758 );
    or g32564 ( n35762 , n32943 , n651 );
    xnor g32565 ( n2222 , n30139 , n16563 );
    not g32566 ( n23154 , n36452 );
    and g32567 ( n23096 , n15677 , n42767 );
    and g32568 ( n2327 , n5734 , n8753 );
    and g32569 ( n6722 , n35733 , n33823 );
    not g32570 ( n16075 , n13713 );
    or g32571 ( n38383 , n32800 , n35571 );
    not g32572 ( n35874 , n478 );
    xnor g32573 ( n42799 , n20070 , n16538 );
    and g32574 ( n21542 , n24057 , n20670 );
    nor g32575 ( n42229 , n30605 , n6542 );
    xnor g32576 ( n16600 , n4692 , n16228 );
    and g32577 ( n24319 , n7427 , n30668 );
    nor g32578 ( n22886 , n41850 , n17537 );
    or g32579 ( n26571 , n34606 , n42357 );
    nor g32580 ( n37368 , n24186 , n13607 );
    and g32581 ( n2125 , n8330 , n26441 );
    nor g32582 ( n34322 , n2375 , n27788 );
    or g32583 ( n12755 , n14250 , n18691 );
    or g32584 ( n15772 , n6132 , n37505 );
    not g32585 ( n21491 , n22875 );
    nor g32586 ( n18096 , n14826 , n8794 );
    and g32587 ( n3927 , n30916 , n4164 );
    xnor g32588 ( n21557 , n10173 , n6927 );
    xnor g32589 ( n41067 , n23322 , n27816 );
    or g32590 ( n29390 , n12112 , n13889 );
    and g32591 ( n25280 , n13592 , n39471 );
    nor g32592 ( n26806 , n2841 , n10475 );
    and g32593 ( n27310 , n31191 , n19669 );
    xnor g32594 ( n16787 , n28101 , n36350 );
    not g32595 ( n18027 , n16709 );
    or g32596 ( n14199 , n10082 , n12051 );
    and g32597 ( n4239 , n2134 , n21412 );
    or g32598 ( n33119 , n323 , n19890 );
    or g32599 ( n3766 , n16479 , n8050 );
    nor g32600 ( n36201 , n21929 , n1064 );
    or g32601 ( n9526 , n13074 , n12284 );
    not g32602 ( n34190 , n20645 );
    or g32603 ( n29022 , n22851 , n18085 );
    and g32604 ( n8891 , n28238 , n37278 );
    and g32605 ( n37220 , n29289 , n12108 );
    nor g32606 ( n37897 , n2795 , n29739 );
    not g32607 ( n24509 , n12530 );
    or g32608 ( n25034 , n7982 , n10579 );
    not g32609 ( n40799 , n2533 );
    or g32610 ( n41568 , n11140 , n12550 );
    and g32611 ( n23202 , n42249 , n1519 );
    or g32612 ( n7664 , n37288 , n37029 );
    or g32613 ( n14028 , n36995 , n24314 );
    and g32614 ( n38887 , n36302 , n31938 );
    and g32615 ( n11215 , n13317 , n31547 );
    not g32616 ( n186 , n34500 );
    or g32617 ( n12143 , n31791 , n21655 );
    or g32618 ( n8652 , n26730 , n40831 );
    not g32619 ( n20700 , n33512 );
    xnor g32620 ( n18644 , n39899 , n490 );
    xnor g32621 ( n42831 , n36491 , n2199 );
    xnor g32622 ( n23816 , n22263 , n27431 );
    nor g32623 ( n41530 , n22030 , n21302 );
    and g32624 ( n8130 , n40608 , n8335 );
    or g32625 ( n29211 , n25964 , n20099 );
    or g32626 ( n25331 , n4839 , n6971 );
    xnor g32627 ( n27620 , n13677 , n18706 );
    or g32628 ( n27445 , n34232 , n17104 );
    or g32629 ( n35457 , n17574 , n34972 );
    nor g32630 ( n14846 , n4190 , n3036 );
    xnor g32631 ( n42242 , n31474 , n4098 );
    and g32632 ( n36488 , n32999 , n10052 );
    and g32633 ( n27703 , n10631 , n36781 );
    or g32634 ( n15148 , n16127 , n26351 );
    or g32635 ( n14367 , n33403 , n8329 );
    and g32636 ( n37330 , n32823 , n7292 );
    and g32637 ( n31514 , n18996 , n1862 );
    or g32638 ( n38449 , n20018 , n35216 );
    or g32639 ( n5873 , n21166 , n16124 );
    nor g32640 ( n8742 , n25348 , n35249 );
    or g32641 ( n21188 , n19580 , n23067 );
    or g32642 ( n21179 , n42896 , n33874 );
    xnor g32643 ( n14760 , n36998 , n30471 );
    nor g32644 ( n16343 , n35720 , n16642 );
    or g32645 ( n38832 , n25483 , n36682 );
    or g32646 ( n8890 , n14707 , n4936 );
    and g32647 ( n19927 , n16958 , n36783 );
    nor g32648 ( n24309 , n42003 , n1609 );
    not g32649 ( n39811 , n9078 );
    or g32650 ( n34233 , n36007 , n12129 );
    nor g32651 ( n11763 , n14828 , n35186 );
    or g32652 ( n28668 , n4924 , n27410 );
    or g32653 ( n16361 , n3573 , n13428 );
    or g32654 ( n33602 , n26518 , n333 );
    or g32655 ( n41050 , n11445 , n18279 );
    or g32656 ( n24762 , n11854 , n41440 );
    or g32657 ( n11070 , n37108 , n21024 );
    not g32658 ( n2571 , n8944 );
    and g32659 ( n29924 , n34563 , n39900 );
    or g32660 ( n3340 , n11340 , n11255 );
    or g32661 ( n40404 , n6779 , n35911 );
    not g32662 ( n32603 , n1294 );
    and g32663 ( n40315 , n24393 , n15815 );
    and g32664 ( n34458 , n36406 , n9050 );
    xnor g32665 ( n58 , n105 , n35375 );
    and g32666 ( n18292 , n15971 , n2046 );
    not g32667 ( n36701 , n23746 );
    or g32668 ( n40815 , n6891 , n2675 );
    and g32669 ( n15026 , n20093 , n2013 );
    or g32670 ( n29055 , n37806 , n12816 );
    and g32671 ( n10650 , n2678 , n38893 );
    or g32672 ( n42029 , n20030 , n38063 );
    or g32673 ( n1760 , n23455 , n32055 );
    xnor g32674 ( n39512 , n36046 , n29100 );
    and g32675 ( n4045 , n2722 , n38792 );
    or g32676 ( n3207 , n16738 , n12839 );
    xnor g32677 ( n3911 , n6914 , n35304 );
    or g32678 ( n32904 , n3602 , n30134 );
    and g32679 ( n20033 , n25374 , n24837 );
    nor g32680 ( n42228 , n16352 , n25181 );
    not g32681 ( n28055 , n34183 );
    not g32682 ( n31970 , n13718 );
    and g32683 ( n40696 , n21222 , n21719 );
    or g32684 ( n42524 , n29782 , n27401 );
    or g32685 ( n32612 , n24734 , n29172 );
    or g32686 ( n29883 , n6683 , n16182 );
    and g32687 ( n16521 , n24225 , n6884 );
    or g32688 ( n28903 , n18407 , n17122 );
    and g32689 ( n20164 , n31193 , n30815 );
    xnor g32690 ( n12704 , n33053 , n10069 );
    and g32691 ( n11688 , n21743 , n28574 );
    or g32692 ( n9429 , n4540 , n9080 );
    and g32693 ( n4185 , n20917 , n4136 );
    xnor g32694 ( n28752 , n35477 , n26601 );
    xnor g32695 ( n40928 , n35727 , n35045 );
    and g32696 ( n23802 , n21701 , n14464 );
    or g32697 ( n25273 , n18929 , n26226 );
    and g32698 ( n27857 , n21520 , n40976 );
    xnor g32699 ( n2241 , n21133 , n28359 );
    or g32700 ( n21121 , n34373 , n3867 );
    not g32701 ( n36561 , n26162 );
    xnor g32702 ( n36007 , n10319 , n40469 );
    nor g32703 ( n6690 , n25917 , n503 );
    or g32704 ( n29972 , n27242 , n31389 );
    nor g32705 ( n5901 , n15647 , n10039 );
    or g32706 ( n15928 , n16590 , n35751 );
    or g32707 ( n108 , n14957 , n11455 );
    or g32708 ( n10876 , n38638 , n26189 );
    or g32709 ( n2390 , n42852 , n40507 );
    or g32710 ( n38298 , n32693 , n42217 );
    xnor g32711 ( n11268 , n22103 , n12046 );
    not g32712 ( n32323 , n23886 );
    and g32713 ( n38112 , n20334 , n5461 );
    nor g32714 ( n20716 , n38879 , n39660 );
    or g32715 ( n37313 , n41865 , n12129 );
    or g32716 ( n34761 , n27477 , n36671 );
    nor g32717 ( n8387 , n1143 , n13309 );
    or g32718 ( n2678 , n27568 , n730 );
    and g32719 ( n7507 , n12273 , n34322 );
    or g32720 ( n4704 , n36618 , n23828 );
    nor g32721 ( n32808 , n19060 , n17913 );
    xnor g32722 ( n7234 , n4385 , n338 );
    or g32723 ( n13266 , n42220 , n11211 );
    and g32724 ( n25202 , n32880 , n40357 );
    or g32725 ( n42681 , n26235 , n23154 );
    or g32726 ( n29180 , n29236 , n38958 );
    or g32727 ( n6591 , n25017 , n17238 );
    not g32728 ( n4511 , n6161 );
    not g32729 ( n13667 , n21291 );
    xnor g32730 ( n8055 , n31099 , n6807 );
    not g32731 ( n26941 , n17722 );
    and g32732 ( n24083 , n185 , n36766 );
    nor g32733 ( n37784 , n29783 , n24456 );
    and g32734 ( n32689 , n13353 , n22908 );
    or g32735 ( n6802 , n3338 , n17321 );
    and g32736 ( n15192 , n23794 , n8603 );
    or g32737 ( n11308 , n14309 , n15787 );
    xnor g32738 ( n23564 , n34875 , n10620 );
    not g32739 ( n3178 , n8430 );
    or g32740 ( n39607 , n14944 , n22676 );
    xnor g32741 ( n19829 , n11537 , n23242 );
    not g32742 ( n19630 , n1615 );
    or g32743 ( n41264 , n19769 , n28254 );
    or g32744 ( n612 , n38060 , n34303 );
    or g32745 ( n36412 , n16909 , n2705 );
    not g32746 ( n12885 , n32118 );
    or g32747 ( n4297 , n25055 , n30906 );
    not g32748 ( n28917 , n11677 );
    xnor g32749 ( n36273 , n25631 , n17341 );
    not g32750 ( n35294 , n41253 );
    and g32751 ( n10742 , n34990 , n3187 );
    nor g32752 ( n33887 , n16728 , n30690 );
    or g32753 ( n25932 , n32684 , n18393 );
    and g32754 ( n29259 , n11250 , n7160 );
    nor g32755 ( n5832 , n25588 , n8169 );
    not g32756 ( n37790 , n10556 );
    and g32757 ( n13889 , n42222 , n11224 );
    not g32758 ( n30176 , n1133 );
    and g32759 ( n11978 , n7906 , n21896 );
    nor g32760 ( n24758 , n39544 , n40598 );
    and g32761 ( n31911 , n2718 , n19420 );
    or g32762 ( n37002 , n2584 , n22767 );
    or g32763 ( n23658 , n34292 , n18606 );
    xnor g32764 ( n10563 , n22903 , n20803 );
    or g32765 ( n11370 , n6170 , n1969 );
    not g32766 ( n2555 , n23020 );
    or g32767 ( n14715 , n25263 , n13121 );
    or g32768 ( n26723 , n37751 , n39635 );
    or g32769 ( n23638 , n36052 , n27132 );
    xnor g32770 ( n42071 , n31099 , n25762 );
    not g32771 ( n36671 , n3428 );
    not g32772 ( n7700 , n21349 );
    or g32773 ( n8895 , n40688 , n26991 );
    not g32774 ( n4447 , n30902 );
    and g32775 ( n8541 , n31533 , n17375 );
    nor g32776 ( n41720 , n33856 , n7786 );
    or g32777 ( n14772 , n222 , n5096 );
    or g32778 ( n2403 , n13516 , n30182 );
    or g32779 ( n16068 , n28503 , n41684 );
    or g32780 ( n24746 , n9787 , n12152 );
    not g32781 ( n34673 , n26957 );
    or g32782 ( n29244 , n29515 , n4421 );
    and g32783 ( n3883 , n784 , n27922 );
    or g32784 ( n18148 , n16464 , n10022 );
    or g32785 ( n9984 , n40018 , n5828 );
    nor g32786 ( n8020 , n5896 , n30666 );
    xnor g32787 ( n14681 , n18624 , n38220 );
    and g32788 ( n3705 , n18941 , n8027 );
    or g32789 ( n3482 , n28243 , n42152 );
    and g32790 ( n12505 , n8878 , n9091 );
    or g32791 ( n22994 , n23472 , n41238 );
    and g32792 ( n22417 , n25020 , n17417 );
    not g32793 ( n14575 , n24504 );
    nor g32794 ( n40430 , n18083 , n10593 );
    not g32795 ( n9691 , n40979 );
    and g32796 ( n24363 , n35067 , n34233 );
    or g32797 ( n20155 , n31037 , n31937 );
    or g32798 ( n17376 , n20682 , n17009 );
    or g32799 ( n15984 , n42083 , n17812 );
    and g32800 ( n21333 , n33093 , n7969 );
    and g32801 ( n32214 , n20203 , n9761 );
    and g32802 ( n15063 , n10573 , n28073 );
    or g32803 ( n33872 , n1488 , n35492 );
    xnor g32804 ( n8256 , n35005 , n16166 );
    or g32805 ( n30516 , n24625 , n23183 );
    not g32806 ( n31734 , n14158 );
    or g32807 ( n26958 , n14471 , n15474 );
    xnor g32808 ( n15067 , n784 , n17460 );
    not g32809 ( n40001 , n7255 );
    or g32810 ( n40923 , n20242 , n41990 );
    nor g32811 ( n34332 , n33422 , n42059 );
    or g32812 ( n26685 , n5552 , n22318 );
    not g32813 ( n40950 , n39112 );
    or g32814 ( n20525 , n12427 , n8401 );
    or g32815 ( n16187 , n37329 , n42851 );
    or g32816 ( n3453 , n9634 , n38164 );
    and g32817 ( n1283 , n29044 , n20676 );
    not g32818 ( n17871 , n8839 );
    or g32819 ( n25883 , n31266 , n31685 );
    xnor g32820 ( n11557 , n26579 , n42195 );
    not g32821 ( n11576 , n38288 );
    or g32822 ( n41651 , n26908 , n22278 );
    nor g32823 ( n27533 , n3769 , n32971 );
    not g32824 ( n20547 , n17157 );
    and g32825 ( n17881 , n26307 , n18615 );
    and g32826 ( n9738 , n27596 , n19893 );
    or g32827 ( n38587 , n34202 , n5085 );
    or g32828 ( n7045 , n10341 , n5578 );
    nor g32829 ( n35302 , n5964 , n41460 );
    nor g32830 ( n12361 , n16598 , n3155 );
    nor g32831 ( n10909 , n31113 , n13995 );
    xnor g32832 ( n30740 , n26475 , n37365 );
    or g32833 ( n14295 , n15544 , n122 );
    nor g32834 ( n9980 , n34787 , n36929 );
    or g32835 ( n407 , n17393 , n3985 );
    or g32836 ( n8231 , n32536 , n40157 );
    nor g32837 ( n3476 , n3348 , n21030 );
    nor g32838 ( n27271 , n31742 , n19351 );
    nor g32839 ( n2746 , n31917 , n944 );
    or g32840 ( n36185 , n39306 , n25784 );
    or g32841 ( n747 , n25577 , n12581 );
    and g32842 ( n17445 , n8827 , n26206 );
    or g32843 ( n11823 , n4667 , n41413 );
    or g32844 ( n11169 , n33267 , n11972 );
    nor g32845 ( n24845 , n29435 , n3341 );
    or g32846 ( n26062 , n25562 , n27738 );
    or g32847 ( n17102 , n6578 , n34073 );
    or g32848 ( n20753 , n38235 , n25787 );
    not g32849 ( n31843 , n18688 );
    or g32850 ( n14660 , n41534 , n9941 );
    or g32851 ( n23432 , n31326 , n30099 );
    not g32852 ( n18131 , n31694 );
    nor g32853 ( n13555 , n10235 , n37003 );
    not g32854 ( n34500 , n41117 );
    nor g32855 ( n5766 , n15800 , n17145 );
    nor g32856 ( n28038 , n20707 , n9802 );
    not g32857 ( n25592 , n17738 );
    xnor g32858 ( n5540 , n5246 , n7030 );
    or g32859 ( n39144 , n9673 , n31913 );
    and g32860 ( n27237 , n5876 , n7584 );
    nor g32861 ( n34684 , n12468 , n7332 );
    and g32862 ( n12758 , n27886 , n23112 );
    or g32863 ( n18643 , n24454 , n7854 );
    or g32864 ( n11043 , n3248 , n9067 );
    nor g32865 ( n20505 , n18681 , n33371 );
    or g32866 ( n23417 , n32740 , n17109 );
    or g32867 ( n21177 , n4097 , n32341 );
    or g32868 ( n5883 , n4660 , n26204 );
    or g32869 ( n42130 , n34636 , n20978 );
    xnor g32870 ( n28600 , n32506 , n41914 );
    and g32871 ( n26391 , n19552 , n35065 );
    or g32872 ( n14446 , n40428 , n21172 );
    or g32873 ( n26050 , n9031 , n10966 );
    and g32874 ( n41319 , n31941 , n28463 );
    or g32875 ( n5274 , n21956 , n27127 );
    nor g32876 ( n18628 , n5964 , n2244 );
    and g32877 ( n17504 , n38047 , n10096 );
    nor g32878 ( n23834 , n1178 , n134 );
    not g32879 ( n42361 , n39226 );
    or g32880 ( n26118 , n7356 , n31114 );
    and g32881 ( n2096 , n28762 , n17463 );
    not g32882 ( n33216 , n7818 );
    and g32883 ( n38529 , n26420 , n2409 );
    or g32884 ( n23217 , n17667 , n4942 );
    nor g32885 ( n1792 , n39692 , n16685 );
    nor g32886 ( n37859 , n10021 , n35699 );
    or g32887 ( n8985 , n39635 , n41676 );
    or g32888 ( n37764 , n25959 , n24776 );
    and g32889 ( n7391 , n28592 , n19656 );
    not g32890 ( n14139 , n4231 );
    not g32891 ( n27450 , n10700 );
    not g32892 ( n26172 , n37478 );
    nor g32893 ( n26408 , n15590 , n12061 );
    xnor g32894 ( n32219 , n35553 , n36761 );
    or g32895 ( n38604 , n33297 , n30999 );
    or g32896 ( n22084 , n39765 , n14460 );
    or g32897 ( n2053 , n8035 , n31543 );
    not g32898 ( n38712 , n38080 );
    or g32899 ( n10824 , n36849 , n17827 );
    or g32900 ( n29535 , n7792 , n25250 );
    or g32901 ( n15637 , n15595 , n21152 );
    or g32902 ( n29260 , n12383 , n31511 );
    not g32903 ( n27434 , n25605 );
    or g32904 ( n33492 , n11480 , n36962 );
    or g32905 ( n9139 , n6835 , n27320 );
    not g32906 ( n3259 , n28095 );
    or g32907 ( n14205 , n8876 , n23361 );
    and g32908 ( n21661 , n40693 , n12810 );
    nor g32909 ( n30284 , n14332 , n15275 );
    or g32910 ( n25720 , n3311 , n18456 );
    nor g32911 ( n7995 , n12476 , n17429 );
    not g32912 ( n26115 , n6337 );
    or g32913 ( n32374 , n11311 , n290 );
    xnor g32914 ( n35603 , n27886 , n23112 );
    nor g32915 ( n7800 , n17387 , n9500 );
    not g32916 ( n35427 , n24931 );
    not g32917 ( n6147 , n11075 );
    or g32918 ( n3044 , n21866 , n3231 );
    and g32919 ( n404 , n27909 , n34012 );
    or g32920 ( n42624 , n21668 , n12114 );
    xnor g32921 ( n33367 , n11596 , n31011 );
    and g32922 ( n12351 , n25944 , n36968 );
    nor g32923 ( n8048 , n22117 , n28396 );
    or g32924 ( n6988 , n36258 , n1223 );
    or g32925 ( n13008 , n564 , n3626 );
    or g32926 ( n12680 , n33692 , n6337 );
    xnor g32927 ( n3970 , n9180 , n42763 );
    or g32928 ( n20524 , n17949 , n22427 );
    or g32929 ( n2874 , n14471 , n16134 );
    or g32930 ( n3718 , n8129 , n18453 );
    xnor g32931 ( n10764 , n40638 , n30118 );
    or g32932 ( n15193 , n19647 , n4238 );
    nor g32933 ( n21352 , n4937 , n41714 );
    not g32934 ( n18477 , n15173 );
    and g32935 ( n33773 , n39266 , n14570 );
    or g32936 ( n41851 , n4560 , n35478 );
    nor g32937 ( n33099 , n17843 , n23001 );
    not g32938 ( n17301 , n20131 );
    and g32939 ( n18490 , n19923 , n6880 );
    and g32940 ( n23328 , n21653 , n30291 );
    not g32941 ( n9814 , n34880 );
    or g32942 ( n6645 , n2801 , n19570 );
    and g32943 ( n17267 , n12908 , n10454 );
    or g32944 ( n27592 , n39526 , n25742 );
    or g32945 ( n11120 , n28454 , n30791 );
    or g32946 ( n32851 , n14471 , n18542 );
    or g32947 ( n31690 , n40295 , n36559 );
    or g32948 ( n13519 , n10902 , n19123 );
    or g32949 ( n25627 , n299 , n33892 );
    nor g32950 ( n35500 , n20707 , n23555 );
    nor g32951 ( n31738 , n34045 , n19705 );
    nor g32952 ( n27973 , n27250 , n34701 );
    and g32953 ( n4705 , n41220 , n4342 );
    and g32954 ( n8560 , n23664 , n25330 );
    and g32955 ( n36827 , n38226 , n40338 );
    and g32956 ( n6035 , n9656 , n37976 );
    and g32957 ( n28236 , n10422 , n10 );
    nor g32958 ( n28045 , n38157 , n42023 );
    not g32959 ( n2645 , n28003 );
    or g32960 ( n6659 , n17258 , n30822 );
    and g32961 ( n13709 , n32993 , n35203 );
    nor g32962 ( n27056 , n29354 , n39675 );
    not g32963 ( n32001 , n25899 );
    or g32964 ( n16219 , n41284 , n24053 );
    nor g32965 ( n20631 , n34565 , n27701 );
    xnor g32966 ( n32232 , n32660 , n33352 );
    or g32967 ( n8687 , n16414 , n439 );
    or g32968 ( n4643 , n28596 , n24603 );
    xnor g32969 ( n1599 , n4334 , n21314 );
    or g32970 ( n21149 , n4305 , n30173 );
    nor g32971 ( n12713 , n15393 , n39792 );
    or g32972 ( n11729 , n32263 , n38352 );
    not g32973 ( n1289 , n9312 );
    or g32974 ( n30545 , n28823 , n37179 );
    and g32975 ( n30998 , n3429 , n23156 );
    or g32976 ( n8517 , n3213 , n1442 );
    and g32977 ( n19723 , n9794 , n4569 );
    or g32978 ( n37920 , n11340 , n41594 );
    nor g32979 ( n40591 , n39456 , n33776 );
    not g32980 ( n1351 , n20230 );
    or g32981 ( n16262 , n34565 , n16441 );
    xnor g32982 ( n18240 , n22346 , n27871 );
    not g32983 ( n2339 , n33130 );
    or g32984 ( n4931 , n24197 , n26992 );
    xnor g32985 ( n30389 , n4304 , n35856 );
    nor g32986 ( n1749 , n1507 , n7833 );
    and g32987 ( n17475 , n38382 , n38477 );
    or g32988 ( n12824 , n13605 , n19890 );
    or g32989 ( n32695 , n37980 , n2392 );
    nor g32990 ( n25353 , n36532 , n802 );
    or g32991 ( n3040 , n15751 , n12669 );
    or g32992 ( n14564 , n792 , n20508 );
    or g32993 ( n5179 , n30068 , n9919 );
    not g32994 ( n22159 , n39384 );
    nor g32995 ( n17183 , n4389 , n24253 );
    or g32996 ( n36801 , n28143 , n799 );
    xnor g32997 ( n13136 , n11436 , n9207 );
    not g32998 ( n22187 , n28177 );
    or g32999 ( n35806 , n21037 , n37381 );
    or g33000 ( n16295 , n23880 , n6492 );
    or g33001 ( n23905 , n39502 , n39098 );
    nor g33002 ( n3806 , n18427 , n14120 );
    and g33003 ( n22554 , n12921 , n11990 );
    xnor g33004 ( n7791 , n37969 , n8908 );
    or g33005 ( n35595 , n36527 , n31070 );
    and g33006 ( n40999 , n29413 , n7614 );
    nor g33007 ( n13254 , n1197 , n30068 );
    not g33008 ( n16398 , n32474 );
    not g33009 ( n19521 , n27776 );
    xnor g33010 ( n31329 , n37074 , n20626 );
    or g33011 ( n19289 , n40192 , n38376 );
    or g33012 ( n27345 , n26965 , n38662 );
    or g33013 ( n3772 , n13063 , n12979 );
    and g33014 ( n29051 , n24580 , n18205 );
    and g33015 ( n4490 , n21370 , n8764 );
    and g33016 ( n13100 , n3615 , n21196 );
    or g33017 ( n6854 , n1048 , n39136 );
    and g33018 ( n20175 , n32076 , n15609 );
    or g33019 ( n41743 , n16736 , n21280 );
    and g33020 ( n2217 , n17873 , n1037 );
    and g33021 ( n24847 , n29377 , n28476 );
    nor g33022 ( n22841 , n16598 , n24521 );
    and g33023 ( n33707 , n37269 , n35164 );
    and g33024 ( n6397 , n10526 , n18177 );
    xnor g33025 ( n12155 , n21765 , n23540 );
    not g33026 ( n24171 , n14669 );
    not g33027 ( n2573 , n34932 );
    nor g33028 ( n28538 , n27762 , n27859 );
    not g33029 ( n25547 , n30510 );
    or g33030 ( n5114 , n5151 , n32826 );
    xnor g33031 ( n1899 , n21559 , n15359 );
    xnor g33032 ( n36426 , n105 , n26342 );
    or g33033 ( n17818 , n4335 , n35332 );
    or g33034 ( n38861 , n21913 , n38175 );
    nor g33035 ( n41566 , n12394 , n24689 );
    or g33036 ( n21061 , n11378 , n36201 );
    or g33037 ( n22698 , n30917 , n28583 );
    and g33038 ( n10395 , n32236 , n21834 );
    or g33039 ( n37140 , n24037 , n40389 );
    not g33040 ( n28389 , n40906 );
    or g33041 ( n22601 , n972 , n27500 );
    or g33042 ( n32522 , n19917 , n15250 );
    and g33043 ( n22670 , n17309 , n3710 );
    or g33044 ( n21447 , n38436 , n18981 );
    and g33045 ( n1200 , n14971 , n19711 );
    nor g33046 ( n41958 , n16323 , n20297 );
    not g33047 ( n30222 , n27622 );
    nor g33048 ( n41600 , n6473 , n8793 );
    xnor g33049 ( n41018 , n8502 , n25464 );
    nor g33050 ( n13774 , n33061 , n39362 );
    and g33051 ( n42623 , n33357 , n807 );
    or g33052 ( n36603 , n37910 , n17756 );
    not g33053 ( n34129 , n10373 );
    or g33054 ( n5088 , n14420 , n33910 );
    or g33055 ( n379 , n33664 , n3854 );
    xnor g33056 ( n96 , n41013 , n39612 );
    nor g33057 ( n7426 , n34349 , n21182 );
    not g33058 ( n35932 , n10010 );
    xnor g33059 ( n22424 , n7567 , n31401 );
    and g33060 ( n232 , n15501 , n1833 );
    xnor g33061 ( n14978 , n26579 , n13384 );
    and g33062 ( n19452 , n15985 , n9352 );
    nor g33063 ( n16805 , n25196 , n12694 );
    or g33064 ( n36127 , n15423 , n30381 );
    or g33065 ( n4832 , n14851 , n35153 );
    and g33066 ( n23957 , n25492 , n3667 );
    xnor g33067 ( n34183 , n13444 , n8545 );
    nor g33068 ( n14879 , n17744 , n2896 );
    or g33069 ( n38209 , n22091 , n27724 );
    not g33070 ( n40222 , n33295 );
    xnor g33071 ( n20082 , n12146 , n16591 );
    xnor g33072 ( n39088 , n27100 , n27885 );
    and g33073 ( n10373 , n30951 , n38642 );
    or g33074 ( n29369 , n29005 , n42758 );
    or g33075 ( n19324 , n33563 , n27016 );
    nor g33076 ( n7952 , n29392 , n31767 );
    nor g33077 ( n5138 , n5896 , n16643 );
    nor g33078 ( n9684 , n27758 , n28885 );
    and g33079 ( n22321 , n8638 , n20773 );
    nor g33080 ( n32510 , n27750 , n34050 );
    not g33081 ( n20111 , n38431 );
    not g33082 ( n3036 , n13668 );
    not g33083 ( n15196 , n19521 );
    nor g33084 ( n25801 , n28874 , n20968 );
    xnor g33085 ( n8045 , n6861 , n37730 );
    xnor g33086 ( n17484 , n2205 , n25125 );
    xnor g33087 ( n24684 , n8437 , n13934 );
    or g33088 ( n97 , n550 , n34981 );
    not g33089 ( n4756 , n11867 );
    not g33090 ( n25145 , n16893 );
    and g33091 ( n19379 , n18276 , n1984 );
    nor g33092 ( n23258 , n19630 , n37913 );
    nor g33093 ( n27018 , n17182 , n37290 );
    or g33094 ( n38051 , n35267 , n16515 );
    xnor g33095 ( n27713 , n35727 , n4312 );
    nor g33096 ( n7011 , n21674 , n11281 );
    or g33097 ( n18452 , n38815 , n22278 );
    nor g33098 ( n2615 , n4027 , n19947 );
    and g33099 ( n13237 , n10775 , n10162 );
    and g33100 ( n28922 , n24425 , n1172 );
    not g33101 ( n18072 , n7156 );
    not g33102 ( n32705 , n2931 );
    or g33103 ( n7705 , n31497 , n15596 );
    xnor g33104 ( n18352 , n4937 , n25790 );
    xnor g33105 ( n28433 , n14331 , n31787 );
    or g33106 ( n22927 , n42381 , n12228 );
    or g33107 ( n32296 , n17642 , n19687 );
    and g33108 ( n32611 , n21061 , n17762 );
    not g33109 ( n25755 , n24472 );
    not g33110 ( n42086 , n24794 );
    nor g33111 ( n19647 , n37216 , n39944 );
    or g33112 ( n36049 , n4212 , n16705 );
    and g33113 ( n16804 , n9286 , n14852 );
    or g33114 ( n35665 , n18767 , n18404 );
    nor g33115 ( n10992 , n39223 , n20572 );
    or g33116 ( n40147 , n35829 , n4273 );
    and g33117 ( n26317 , n27882 , n42194 );
    and g33118 ( n39936 , n39780 , n14173 );
    or g33119 ( n25695 , n14684 , n38605 );
    and g33120 ( n30909 , n1570 , n5223 );
    and g33121 ( n13034 , n26715 , n16945 );
    or g33122 ( n11811 , n31824 , n21109 );
    or g33123 ( n6564 , n21702 , n40551 );
    or g33124 ( n9152 , n10997 , n42387 );
    or g33125 ( n41104 , n21893 , n4933 );
    nor g33126 ( n22949 , n1466 , n40811 );
    or g33127 ( n28367 , n6638 , n39159 );
    nor g33128 ( n34123 , n35301 , n41456 );
    or g33129 ( n23344 , n19882 , n42544 );
    nor g33130 ( n11395 , n22022 , n29412 );
    nor g33131 ( n1472 , n30818 , n24015 );
    or g33132 ( n11265 , n8665 , n2565 );
    or g33133 ( n7630 , n8145 , n7306 );
    nor g33134 ( n31534 , n6952 , n40402 );
    and g33135 ( n12075 , n33886 , n3638 );
    not g33136 ( n25582 , n28632 );
    or g33137 ( n8702 , n38900 , n41317 );
    and g33138 ( n24193 , n1840 , n5851 );
    xnor g33139 ( n40701 , n22604 , n10669 );
    or g33140 ( n4322 , n12812 , n38767 );
    or g33141 ( n30394 , n16586 , n35491 );
    and g33142 ( n39679 , n12824 , n20912 );
    or g33143 ( n27242 , n910 , n5183 );
    not g33144 ( n34697 , n21405 );
    xnor g33145 ( n9615 , n2005 , n9424 );
    and g33146 ( n30948 , n21389 , n31706 );
    and g33147 ( n6571 , n39629 , n30925 );
    nor g33148 ( n13247 , n2370 , n35992 );
    and g33149 ( n21970 , n3360 , n15745 );
    nor g33150 ( n21260 , n35301 , n12515 );
    or g33151 ( n20576 , n27761 , n35858 );
    and g33152 ( n8912 , n34487 , n40098 );
    not g33153 ( n18219 , n27481 );
    xnor g33154 ( n39427 , n6962 , n6501 );
    not g33155 ( n38463 , n24737 );
    not g33156 ( n10850 , n20435 );
    and g33157 ( n1181 , n27793 , n17900 );
    not g33158 ( n7386 , n31045 );
    nor g33159 ( n14546 , n37616 , n9037 );
    and g33160 ( n14266 , n24550 , n16370 );
    or g33161 ( n2640 , n26922 , n17503 );
    or g33162 ( n5601 , n39681 , n39715 );
    nor g33163 ( n11040 , n35876 , n24188 );
    nor g33164 ( n15187 , n7744 , n1413 );
    not g33165 ( n6106 , n369 );
    and g33166 ( n40139 , n18258 , n38434 );
    nor g33167 ( n15233 , n14471 , n23795 );
    or g33168 ( n14632 , n282 , n7460 );
    nor g33169 ( n32386 , n39705 , n9470 );
    nor g33170 ( n1859 , n40472 , n23998 );
    or g33171 ( n13479 , n28745 , n18141 );
    nor g33172 ( n1704 , n25468 , n20172 );
    nor g33173 ( n11347 , n4228 , n30802 );
    not g33174 ( n22966 , n17696 );
    and g33175 ( n35635 , n41901 , n39007 );
    and g33176 ( n32803 , n10540 , n6513 );
    or g33177 ( n28976 , n36117 , n25470 );
    xnor g33178 ( n11481 , n15706 , n34194 );
    and g33179 ( n36839 , n35783 , n25044 );
    xnor g33180 ( n32920 , n5042 , n19580 );
    nor g33181 ( n7727 , n38879 , n10506 );
    or g33182 ( n35862 , n3034 , n38677 );
    or g33183 ( n22416 , n11993 , n26830 );
    or g33184 ( n40508 , n2230 , n30523 );
    and g33185 ( n20451 , n22085 , n25720 );
    or g33186 ( n14151 , n40832 , n40110 );
    xnor g33187 ( n8689 , n1544 , n3241 );
    xnor g33188 ( n21740 , n10443 , n33221 );
    or g33189 ( n2433 , n31441 , n35268 );
    not g33190 ( n18093 , n23948 );
    nor g33191 ( n38820 , n30743 , n23717 );
    or g33192 ( n21422 , n3331 , n1631 );
    nor g33193 ( n38333 , n27786 , n16966 );
    nor g33194 ( n24146 , n32084 , n25609 );
    or g33195 ( n685 , n21950 , n7319 );
    xnor g33196 ( n19706 , n20986 , n17289 );
    or g33197 ( n20203 , n40261 , n15726 );
    and g33198 ( n133 , n21991 , n4399 );
    or g33199 ( n21993 , n9673 , n20107 );
    not g33200 ( n32949 , n23259 );
    nor g33201 ( n5805 , n21907 , n6845 );
    or g33202 ( n6447 , n11667 , n6813 );
    and g33203 ( n26132 , n14033 , n16557 );
    xnor g33204 ( n27002 , n2551 , n25385 );
    not g33205 ( n1254 , n16890 );
    and g33206 ( n15267 , n14418 , n561 );
    nor g33207 ( n28700 , n36017 , n20466 );
    or g33208 ( n35079 , n7687 , n40805 );
    or g33209 ( n35252 , n30276 , n4923 );
    xnor g33210 ( n14606 , n5441 , n34523 );
    or g33211 ( n30436 , n11410 , n16142 );
    nor g33212 ( n41898 , n37149 , n34392 );
    not g33213 ( n141 , n7999 );
    xnor g33214 ( n26662 , n28443 , n4946 );
    not g33215 ( n22437 , n17426 );
    or g33216 ( n33364 , n20302 , n17404 );
    not g33217 ( n7221 , n40136 );
    or g33218 ( n41612 , n7027 , n34009 );
    and g33219 ( n23335 , n1362 , n18040 );
    or g33220 ( n18790 , n31580 , n8391 );
    nor g33221 ( n6576 , n5926 , n32856 );
    or g33222 ( n3746 , n38250 , n31618 );
    not g33223 ( n33345 , n30826 );
    or g33224 ( n11018 , n35516 , n7972 );
    or g33225 ( n42835 , n32375 , n22282 );
    or g33226 ( n13799 , n40852 , n29234 );
    nor g33227 ( n7973 , n20890 , n31993 );
    or g33228 ( n25490 , n39539 , n15606 );
    xnor g33229 ( n7105 , n22888 , n32051 );
    not g33230 ( n12198 , n22074 );
    nor g33231 ( n27502 , n5964 , n37752 );
    and g33232 ( n40041 , n30109 , n2670 );
    and g33233 ( n4970 , n26529 , n37551 );
    not g33234 ( n29854 , n6660 );
    or g33235 ( n41910 , n7250 , n41215 );
    xnor g33236 ( n37908 , n38749 , n10680 );
    xnor g33237 ( n2953 , n26579 , n2124 );
    or g33238 ( n42158 , n31805 , n33537 );
    nor g33239 ( n3561 , n40067 , n18072 );
    xnor g33240 ( n4007 , n9336 , n10568 );
    nor g33241 ( n2319 , n4879 , n27673 );
    and g33242 ( n32221 , n35220 , n998 );
    or g33243 ( n34904 , n31516 , n1006 );
    or g33244 ( n4194 , n36633 , n20498 );
    and g33245 ( n31527 , n20847 , n12855 );
    or g33246 ( n34280 , n35856 , n29930 );
    not g33247 ( n6331 , n16033 );
    nor g33248 ( n23289 , n34698 , n36219 );
    or g33249 ( n34450 , n11234 , n16852 );
    or g33250 ( n14655 , n42425 , n17187 );
    not g33251 ( n20548 , n28404 );
    not g33252 ( n41699 , n17880 );
    not g33253 ( n2956 , n28347 );
    or g33254 ( n20295 , n32508 , n11455 );
    nor g33255 ( n12489 , n12773 , n24148 );
    nor g33256 ( n23438 , n14658 , n37519 );
    or g33257 ( n14592 , n28443 , n35747 );
    not g33258 ( n26345 , n16582 );
    nor g33259 ( n21220 , n5964 , n21375 );
    nor g33260 ( n39837 , n3735 , n20616 );
    or g33261 ( n36737 , n38882 , n40481 );
    or g33262 ( n42551 , n20684 , n22075 );
    nor g33263 ( n11126 , n21911 , n1530 );
    or g33264 ( n2367 , n28015 , n15900 );
    nor g33265 ( n26192 , n26195 , n20329 );
    not g33266 ( n28395 , n25691 );
    or g33267 ( n13131 , n28647 , n29172 );
    or g33268 ( n16017 , n24656 , n36291 );
    xnor g33269 ( n29963 , n36625 , n32488 );
    not g33270 ( n2213 , n22310 );
    or g33271 ( n17384 , n7822 , n35364 );
    not g33272 ( n27179 , n23667 );
    and g33273 ( n34273 , n20396 , n6668 );
    and g33274 ( n14157 , n11081 , n13739 );
    xnor g33275 ( n31310 , n784 , n40431 );
    xnor g33276 ( n35826 , n5144 , n4441 );
    or g33277 ( n26453 , n9329 , n21224 );
    xnor g33278 ( n10003 , n22346 , n39507 );
    not g33279 ( n5528 , n10769 );
    or g33280 ( n9136 , n780 , n28273 );
    not g33281 ( n31736 , n5985 );
    or g33282 ( n42599 , n2854 , n17640 );
    nor g33283 ( n39869 , n7421 , n14844 );
    nor g33284 ( n37138 , n32964 , n29252 );
    or g33285 ( n7470 , n18268 , n8276 );
    or g33286 ( n21322 , n11725 , n35442 );
    xnor g33287 ( n9367 , n11436 , n20825 );
    and g33288 ( n10060 , n3453 , n17571 );
    or g33289 ( n35181 , n9049 , n14668 );
    and g33290 ( n29913 , n25076 , n41166 );
    or g33291 ( n18616 , n34750 , n34447 );
    or g33292 ( n1531 , n21953 , n20473 );
    not g33293 ( n24753 , n33428 );
    nor g33294 ( n8806 , n25060 , n2765 );
    or g33295 ( n16252 , n10045 , n42171 );
    and g33296 ( n40656 , n31672 , n35136 );
    or g33297 ( n23546 , n32708 , n38264 );
    and g33298 ( n37698 , n334 , n8139 );
    nor g33299 ( n16447 , n18320 , n33328 );
    and g33300 ( n4033 , n41303 , n33956 );
    and g33301 ( n8178 , n14833 , n13406 );
    not g33302 ( n37233 , n13372 );
    not g33303 ( n40271 , n14975 );
    or g33304 ( n37986 , n5964 , n42588 );
    or g33305 ( n32833 , n33407 , n22363 );
    or g33306 ( n14674 , n18866 , n17856 );
    or g33307 ( n36555 , n5419 , n6302 );
    xnor g33308 ( n35030 , n2921 , n17504 );
    nor g33309 ( n15653 , n10652 , n8153 );
    xnor g33310 ( n25714 , n32452 , n21119 );
    or g33311 ( n42107 , n21048 , n42894 );
    not g33312 ( n33643 , n7986 );
    not g33313 ( n1757 , n957 );
    and g33314 ( n36096 , n39202 , n104 );
    not g33315 ( n22835 , n3033 );
    nor g33316 ( n18058 , n2199 , n26399 );
    nor g33317 ( n25252 , n35497 , n13493 );
    not g33318 ( n6557 , n35932 );
    xnor g33319 ( n24642 , n42181 , n15817 );
    and g33320 ( n26777 , n38260 , n16213 );
    xnor g33321 ( n12221 , n21929 , n20390 );
    or g33322 ( n8531 , n27145 , n8034 );
    or g33323 ( n23358 , n29214 , n27269 );
    or g33324 ( n22865 , n5153 , n14668 );
    not g33325 ( n227 , n39851 );
    or g33326 ( n2002 , n21771 , n3481 );
    not g33327 ( n40720 , n39287 );
    not g33328 ( n38494 , n21106 );
    nor g33329 ( n32965 , n14707 , n24609 );
    not g33330 ( n24483 , n32229 );
    or g33331 ( n2997 , n4236 , n9617 );
    and g33332 ( n20352 , n37832 , n27113 );
    or g33333 ( n14044 , n28423 , n1995 );
    or g33334 ( n13289 , n40818 , n20146 );
    nor g33335 ( n5796 , n8494 , n10880 );
    and g33336 ( n4815 , n20340 , n11536 );
    and g33337 ( n12121 , n40542 , n11386 );
    or g33338 ( n8448 , n13833 , n10032 );
    not g33339 ( n29614 , n350 );
    nor g33340 ( n6122 , n33981 , n34315 );
    or g33341 ( n38948 , n22821 , n31779 );
    and g33342 ( n5109 , n22263 , n4664 );
    not g33343 ( n12866 , n7110 );
    xnor g33344 ( n30154 , n21954 , n36322 );
    or g33345 ( n37246 , n29388 , n37690 );
    or g33346 ( n41755 , n11024 , n4496 );
    or g33347 ( n10807 , n12495 , n39702 );
    not g33348 ( n14870 , n27744 );
    xnor g33349 ( n10117 , n12161 , n3750 );
    nor g33350 ( n4412 , n35005 , n3941 );
    or g33351 ( n12472 , n29043 , n26664 );
    or g33352 ( n30518 , n28774 , n32719 );
    not g33353 ( n2408 , n21195 );
    or g33354 ( n22627 , n41728 , n16553 );
    not g33355 ( n17971 , n24957 );
    or g33356 ( n38891 , n24975 , n31671 );
    and g33357 ( n39483 , n14347 , n14372 );
    and g33358 ( n12096 , n25880 , n22541 );
    and g33359 ( n40342 , n25495 , n7301 );
    not g33360 ( n3231 , n5655 );
    not g33361 ( n30189 , n39068 );
    nor g33362 ( n13057 , n21309 , n32027 );
    not g33363 ( n39558 , n7067 );
    xnor g33364 ( n25149 , n39994 , n39427 );
    nor g33365 ( n30860 , n1507 , n16095 );
    not g33366 ( n17647 , n8759 );
    nor g33367 ( n32670 , n21371 , n2907 );
    not g33368 ( n40472 , n35871 );
    or g33369 ( n17751 , n3487 , n26840 );
    or g33370 ( n3492 , n15070 , n6769 );
    and g33371 ( n5181 , n19708 , n40470 );
    xnor g33372 ( n23550 , n36697 , n21334 );
    or g33373 ( n20577 , n41940 , n26508 );
    not g33374 ( n5430 , n42672 );
    xnor g33375 ( n15647 , n28867 , n13671 );
    xnor g33376 ( n29088 , n31539 , n6418 );
    or g33377 ( n31400 , n19969 , n25157 );
    or g33378 ( n27646 , n13486 , n41966 );
    xnor g33379 ( n14908 , n34968 , n25287 );
    not g33380 ( n40398 , n26494 );
    not g33381 ( n23088 , n19316 );
    and g33382 ( n11920 , n39296 , n2861 );
    or g33383 ( n24228 , n30652 , n21276 );
    or g33384 ( n35110 , n5229 , n40147 );
    or g33385 ( n16584 , n32277 , n33940 );
    and g33386 ( n2878 , n2267 , n20530 );
    not g33387 ( n37697 , n26472 );
    xnor g33388 ( n31546 , n35035 , n33431 );
    xnor g33389 ( n34294 , n20956 , n1446 );
    or g33390 ( n11042 , n35301 , n17410 );
    not g33391 ( n9402 , n28183 );
    not g33392 ( n14129 , n3940 );
    or g33393 ( n18201 , n39105 , n27434 );
    nor g33394 ( n15990 , n18275 , n15014 );
    and g33395 ( n28475 , n2391 , n38419 );
    or g33396 ( n3899 , n26337 , n38338 );
    not g33397 ( n16605 , n23963 );
    and g33398 ( n13689 , n32283 , n38447 );
    or g33399 ( n28023 , n5818 , n30529 );
    or g33400 ( n37221 , n36162 , n42080 );
    or g33401 ( n6091 , n17345 , n24020 );
    or g33402 ( n12992 , n9031 , n10854 );
    or g33403 ( n16713 , n25877 , n5841 );
    or g33404 ( n16326 , n2472 , n25820 );
    nor g33405 ( n18085 , n10539 , n30703 );
    or g33406 ( n1486 , n6574 , n20412 );
    not g33407 ( n9319 , n3264 );
    not g33408 ( n8611 , n13140 );
    or g33409 ( n6534 , n13381 , n14944 );
    xnor g33410 ( n28299 , n41013 , n6254 );
    not g33411 ( n34009 , n40878 );
    xnor g33412 ( n18295 , n2338 , n32258 );
    or g33413 ( n11608 , n18452 , n27393 );
    or g33414 ( n15554 , n38524 , n32233 );
    and g33415 ( n42894 , n7128 , n2122 );
    or g33416 ( n15234 , n277 , n4259 );
    or g33417 ( n28218 , n2213 , n11674 );
    not g33418 ( n37953 , n4746 );
    or g33419 ( n350 , n13511 , n17634 );
    or g33420 ( n9123 , n28979 , n37576 );
    xnor g33421 ( n10782 , n23686 , n7283 );
    nor g33422 ( n41971 , n589 , n38119 );
    not g33423 ( n20015 , n13696 );
    or g33424 ( n14742 , n26444 , n12549 );
    or g33425 ( n30584 , n23085 , n24664 );
    or g33426 ( n22596 , n41534 , n2584 );
    xnor g33427 ( n18251 , n2862 , n20189 );
    or g33428 ( n5235 , n38791 , n328 );
    or g33429 ( n19794 , n2256 , n34225 );
    and g33430 ( n9947 , n6687 , n23403 );
    not g33431 ( n18637 , n21303 );
    or g33432 ( n18955 , n21304 , n30652 );
    or g33433 ( n29198 , n935 , n41536 );
    xnor g33434 ( n16391 , n5144 , n25537 );
    and g33435 ( n31299 , n18370 , n33736 );
    xnor g33436 ( n42474 , n32632 , n24251 );
    or g33437 ( n9830 , n4802 , n25007 );
    and g33438 ( n25458 , n17265 , n37681 );
    or g33439 ( n6466 , n9748 , n37703 );
    or g33440 ( n40648 , n1673 , n24068 );
    or g33441 ( n20396 , n3893 , n28989 );
    not g33442 ( n29388 , n37446 );
    and g33443 ( n30266 , n39031 , n652 );
    and g33444 ( n42787 , n29078 , n17068 );
    or g33445 ( n26804 , n33088 , n6554 );
    and g33446 ( n3351 , n28431 , n5973 );
    xnor g33447 ( n37543 , n32794 , n3919 );
    not g33448 ( n9448 , n40912 );
    or g33449 ( n9517 , n24471 , n8226 );
    and g33450 ( n20413 , n41830 , n20655 );
    and g33451 ( n36115 , n6600 , n16668 );
    or g33452 ( n12390 , n23819 , n25530 );
    nor g33453 ( n6349 , n12372 , n11040 );
    or g33454 ( n15629 , n13832 , n34941 );
    nor g33455 ( n34740 , n41220 , n4342 );
    nor g33456 ( n39215 , n17120 , n12756 );
    xnor g33457 ( n31585 , n33473 , n16598 );
    or g33458 ( n33335 , n37805 , n10477 );
    not g33459 ( n17746 , n16335 );
    not g33460 ( n2857 , n1 );
    or g33461 ( n3819 , n8004 , n30602 );
    not g33462 ( n13063 , n215 );
    and g33463 ( n6154 , n26668 , n12827 );
    or g33464 ( n40034 , n33743 , n42153 );
    or g33465 ( n11803 , n42514 , n34467 );
    or g33466 ( n30337 , n34373 , n4933 );
    or g33467 ( n19481 , n28725 , n34473 );
    or g33468 ( n3400 , n11511 , n7220 );
    or g33469 ( n13845 , n23503 , n14195 );
    or g33470 ( n15393 , n16970 , n37992 );
    or g33471 ( n30755 , n14422 , n547 );
    and g33472 ( n40867 , n16011 , n2378 );
    or g33473 ( n17014 , n5500 , n42479 );
    or g33474 ( n26819 , n25802 , n23172 );
    xnor g33475 ( n17716 , n15089 , n33582 );
    or g33476 ( n24522 , n41426 , n31493 );
    and g33477 ( n21850 , n15613 , n27805 );
    or g33478 ( n38446 , n5896 , n20302 );
    or g33479 ( n10849 , n24895 , n34634 );
    xnor g33480 ( n20685 , n527 , n37947 );
    and g33481 ( n29625 , n17081 , n1775 );
    nor g33482 ( n4357 , n34387 , n13468 );
    or g33483 ( n29923 , n3242 , n2465 );
    or g33484 ( n504 , n26863 , n41922 );
    and g33485 ( n1334 , n5592 , n26148 );
    and g33486 ( n6110 , n18150 , n17791 );
    not g33487 ( n37500 , n29723 );
    and g33488 ( n36082 , n33347 , n10478 );
    and g33489 ( n25250 , n17319 , n36609 );
    or g33490 ( n21643 , n1940 , n42119 );
    nor g33491 ( n28705 , n14021 , n18461 );
    nor g33492 ( n40839 , n12837 , n9485 );
    and g33493 ( n22911 , n37701 , n34612 );
    not g33494 ( n17383 , n11151 );
    not g33495 ( n5582 , n2101 );
    and g33496 ( n39651 , n18540 , n26937 );
    or g33497 ( n30494 , n36253 , n25640 );
    not g33498 ( n9275 , n31138 );
    and g33499 ( n14036 , n41652 , n42400 );
    nor g33500 ( n4899 , n35005 , n3521 );
    nor g33501 ( n41472 , n10434 , n15359 );
    nor g33502 ( n11129 , n41187 , n25443 );
    xnor g33503 ( n38906 , n6625 , n38940 );
    or g33504 ( n31328 , n39213 , n36915 );
    or g33505 ( n31240 , n34128 , n34561 );
    nor g33506 ( n23925 , n38242 , n4256 );
    and g33507 ( n36745 , n25691 , n27794 );
    and g33508 ( n14081 , n22835 , n35167 );
    and g33509 ( n24957 , n30217 , n4110 );
    not g33510 ( n35144 , n12873 );
    or g33511 ( n30761 , n22401 , n29539 );
    not g33512 ( n35269 , n2535 );
    or g33513 ( n34833 , n25108 , n13649 );
    or g33514 ( n13978 , n34224 , n5554 );
    and g33515 ( n2181 , n36042 , n35821 );
    or g33516 ( n27350 , n23748 , n25626 );
    not g33517 ( n37040 , n13577 );
    and g33518 ( n21156 , n12247 , n37556 );
    xnor g33519 ( n11942 , n40025 , n24970 );
    or g33520 ( n490 , n2216 , n778 );
    or g33521 ( n188 , n40057 , n28740 );
    or g33522 ( n13537 , n35266 , n25210 );
    not g33523 ( n13523 , n33974 );
    or g33524 ( n18416 , n22172 , n223 );
    and g33525 ( n26638 , n4953 , n35130 );
    or g33526 ( n2527 , n36272 , n3798 );
    xnor g33527 ( n27107 , n5177 , n11363 );
    not g33528 ( n6442 , n25025 );
    not g33529 ( n25348 , n31665 );
    not g33530 ( n10902 , n7702 );
    and g33531 ( n17717 , n38310 , n3500 );
    nor g33532 ( n11930 , n36028 , n13995 );
    xnor g33533 ( n36655 , n39217 , n12072 );
    or g33534 ( n19368 , n11057 , n28235 );
    or g33535 ( n6608 , n33755 , n12258 );
    and g33536 ( n17367 , n9483 , n7284 );
    and g33537 ( n7977 , n4846 , n27254 );
    not g33538 ( n35142 , n29610 );
    or g33539 ( n21401 , n17707 , n35057 );
    or g33540 ( n9323 , n14944 , n25488 );
    or g33541 ( n32758 , n35879 , n35503 );
    and g33542 ( n36767 , n33007 , n26469 );
    and g33543 ( n17026 , n68 , n9756 );
    and g33544 ( n32812 , n13969 , n29869 );
    and g33545 ( n14998 , n27602 , n36714 );
    not g33546 ( n5022 , n1430 );
    or g33547 ( n6853 , n2175 , n1257 );
    nor g33548 ( n21211 , n19471 , n38245 );
    not g33549 ( n14562 , n10918 );
    or g33550 ( n16372 , n37763 , n16625 );
    or g33551 ( n3725 , n16910 , n25689 );
    or g33552 ( n13879 , n1020 , n7996 );
    not g33553 ( n3574 , n30958 );
    or g33554 ( n34805 , n37633 , n26728 );
    and g33555 ( n18293 , n4920 , n16386 );
    not g33556 ( n12984 , n426 );
    or g33557 ( n23605 , n42782 , n42860 );
    nor g33558 ( n32451 , n36117 , n36155 );
    or g33559 ( n214 , n30130 , n42701 );
    and g33560 ( n24535 , n14815 , n17115 );
    or g33561 ( n38096 , n28623 , n3543 );
    nor g33562 ( n7711 , n6885 , n5131 );
    not g33563 ( n14972 , n40916 );
    nor g33564 ( n26374 , n16333 , n30297 );
    nor g33565 ( n35251 , n2971 , n6848 );
    or g33566 ( n13729 , n12590 , n25741 );
    or g33567 ( n3419 , n35029 , n20498 );
    not g33568 ( n1664 , n12224 );
    or g33569 ( n20365 , n10728 , n3017 );
    nor g33570 ( n11390 , n8084 , n36978 );
    or g33571 ( n26043 , n18811 , n9558 );
    nor g33572 ( n9130 , n31480 , n21470 );
    or g33573 ( n6081 , n5605 , n15238 );
    or g33574 ( n34580 , n12711 , n38152 );
    xnor g33575 ( n10445 , n22346 , n8254 );
    nor g33576 ( n42618 , n22877 , n21825 );
    not g33577 ( n3134 , n35126 );
    not g33578 ( n272 , n26422 );
    or g33579 ( n33908 , n34594 , n42255 );
    or g33580 ( n17593 , n37842 , n4724 );
    and g33581 ( n18107 , n3550 , n41029 );
    or g33582 ( n37626 , n20932 , n372 );
    or g33583 ( n20918 , n3637 , n31692 );
    nor g33584 ( n22171 , n31050 , n26055 );
    or g33585 ( n24686 , n3521 , n23472 );
    not g33586 ( n9196 , n20471 );
    nor g33587 ( n36739 , n25588 , n4478 );
    nor g33588 ( n16833 , n31906 , n25772 );
    or g33589 ( n11309 , n17249 , n26470 );
    or g33590 ( n11625 , n6754 , n30113 );
    or g33591 ( n7304 , n18753 , n18533 );
    nor g33592 ( n28827 , n10929 , n35100 );
    nor g33593 ( n26099 , n4651 , n25865 );
    not g33594 ( n5824 , n5393 );
    and g33595 ( n25329 , n24132 , n30890 );
    xnor g33596 ( n2442 , n3840 , n35598 );
    or g33597 ( n24562 , n14384 , n19356 );
    nor g33598 ( n22075 , n34835 , n2010 );
    and g33599 ( n40637 , n32120 , n13233 );
    or g33600 ( n14858 , n29932 , n17544 );
    or g33601 ( n35003 , n22964 , n19953 );
    and g33602 ( n42577 , n41773 , n38012 );
    or g33603 ( n23676 , n26325 , n40612 );
    and g33604 ( n21725 , n35030 , n28659 );
    or g33605 ( n40606 , n7615 , n151 );
    and g33606 ( n37106 , n19306 , n18547 );
    or g33607 ( n34742 , n2368 , n29462 );
    xnor g33608 ( n36058 , n11534 , n39679 );
    xnor g33609 ( n40942 , n14638 , n8161 );
    not g33610 ( n2130 , n28956 );
    not g33611 ( n35352 , n10619 );
    or g33612 ( n28 , n30796 , n14199 );
    or g33613 ( n10551 , n29027 , n25928 );
    xnor g33614 ( n14078 , n4784 , n40598 );
    nor g33615 ( n14410 , n34090 , n12807 );
    or g33616 ( n23387 , n8494 , n816 );
    or g33617 ( n5108 , n20201 , n26935 );
    or g33618 ( n8678 , n31918 , n37742 );
    or g33619 ( n4399 , n27019 , n41954 );
    nor g33620 ( n30092 , n38382 , n38477 );
    not g33621 ( n27499 , n28444 );
    or g33622 ( n6321 , n17911 , n41776 );
    or g33623 ( n35054 , n19599 , n39299 );
    not g33624 ( n15186 , n28662 );
    and g33625 ( n10605 , n19967 , n42499 );
    or g33626 ( n29130 , n41466 , n24830 );
    or g33627 ( n8933 , n34192 , n41376 );
    and g33628 ( n7747 , n22994 , n3374 );
    nor g33629 ( n28674 , n4671 , n13559 );
    xnor g33630 ( n13977 , n36009 , n19015 );
    or g33631 ( n9905 , n28035 , n23211 );
    not g33632 ( n4029 , n19351 );
    and g33633 ( n12766 , n36680 , n23854 );
    or g33634 ( n9965 , n35250 , n38052 );
    not g33635 ( n24114 , n14575 );
    not g33636 ( n12057 , n40927 );
    not g33637 ( n10587 , n35766 );
    or g33638 ( n1257 , n40785 , n14874 );
    or g33639 ( n13268 , n34954 , n8482 );
    and g33640 ( n1168 , n32469 , n7705 );
    and g33641 ( n24701 , n17811 , n15309 );
    or g33642 ( n42812 , n18314 , n12961 );
    or g33643 ( n27451 , n8626 , n41226 );
    and g33644 ( n29268 , n15324 , n37267 );
    and g33645 ( n13256 , n23147 , n4466 );
    and g33646 ( n26269 , n4196 , n34145 );
    not g33647 ( n40214 , n17055 );
    xnor g33648 ( n23938 , n32470 , n20232 );
    not g33649 ( n25681 , n13895 );
    nor g33650 ( n19930 , n42529 , n22745 );
    or g33651 ( n15030 , n32084 , n2284 );
    or g33652 ( n42014 , n28472 , n23065 );
    xnor g33653 ( n20673 , n31099 , n21976 );
    not g33654 ( n8442 , n112 );
    nor g33655 ( n17538 , n8494 , n26502 );
    not g33656 ( n38105 , n7673 );
    and g33657 ( n40170 , n13017 , n41379 );
    or g33658 ( n2509 , n39383 , n27863 );
    or g33659 ( n34702 , n38688 , n391 );
    not g33660 ( n34039 , n9006 );
    and g33661 ( n36466 , n10924 , n1392 );
    not g33662 ( n22649 , n9843 );
    nor g33663 ( n33107 , n7342 , n338 );
    and g33664 ( n5654 , n8437 , n13934 );
    nor g33665 ( n17642 , n14188 , n22814 );
    and g33666 ( n25424 , n38543 , n14376 );
    not g33667 ( n3715 , n36809 );
    or g33668 ( n26283 , n1560 , n21899 );
    and g33669 ( n20749 , n27800 , n39132 );
    or g33670 ( n2920 , n3690 , n27666 );
    or g33671 ( n22881 , n38865 , n33297 );
    or g33672 ( n8445 , n6636 , n42796 );
    and g33673 ( n1456 , n18233 , n11817 );
    or g33674 ( n22931 , n19753 , n13128 );
    not g33675 ( n21248 , n14550 );
    or g33676 ( n5479 , n17742 , n9010 );
    and g33677 ( n26710 , n4367 , n23603 );
    or g33678 ( n31890 , n40066 , n15186 );
    or g33679 ( n39499 , n38359 , n14776 );
    not g33680 ( n27223 , n40153 );
    or g33681 ( n32107 , n41767 , n13552 );
    and g33682 ( n22250 , n27668 , n22258 );
    not g33683 ( n23772 , n6176 );
    nor g33684 ( n31998 , n32480 , n5046 );
    nor g33685 ( n20810 , n28132 , n30883 );
    and g33686 ( n40626 , n10000 , n36634 );
    not g33687 ( n27081 , n37478 );
    xnor g33688 ( n40130 , n11633 , n5131 );
    xnor g33689 ( n5907 , n41218 , n33653 );
    not g33690 ( n39632 , n11160 );
    or g33691 ( n15715 , n19518 , n34569 );
    nor g33692 ( n31703 , n7029 , n39380 );
    nor g33693 ( n19790 , n2199 , n32320 );
    xnor g33694 ( n26855 , n13785 , n36492 );
    and g33695 ( n5847 , n18189 , n3507 );
    and g33696 ( n14836 , n2443 , n14437 );
    or g33697 ( n41931 , n3090 , n42702 );
    nor g33698 ( n558 , n17625 , n6368 );
    and g33699 ( n38512 , n25 , n19583 );
    or g33700 ( n42371 , n18020 , n27111 );
    and g33701 ( n25485 , n24630 , n30057 );
    or g33702 ( n7578 , n41313 , n10740 );
    nor g33703 ( n4982 , n9060 , n7198 );
    or g33704 ( n24706 , n36787 , n29388 );
    not g33705 ( n3276 , n14187 );
    and g33706 ( n5350 , n31536 , n15081 );
    or g33707 ( n17185 , n26961 , n29755 );
    xnor g33708 ( n28463 , n784 , n16948 );
    or g33709 ( n37396 , n15512 , n52 );
    or g33710 ( n29035 , n15513 , n14503 );
    and g33711 ( n3330 , n34530 , n6485 );
    or g33712 ( n27405 , n19135 , n42137 );
    and g33713 ( n33182 , n31969 , n41798 );
    or g33714 ( n37214 , n7542 , n21268 );
    not g33715 ( n21404 , n20967 );
    or g33716 ( n14071 , n7057 , n10022 );
    and g33717 ( n4824 , n24987 , n14482 );
    and g33718 ( n19509 , n32584 , n10938 );
    and g33719 ( n32242 , n22300 , n28628 );
    and g33720 ( n16222 , n33935 , n31442 );
    or g33721 ( n12030 , n8487 , n9103 );
    nor g33722 ( n42723 , n14614 , n15719 );
    nor g33723 ( n33727 , n4821 , n15290 );
    and g33724 ( n28416 , n17852 , n14667 );
    and g33725 ( n20896 , n35854 , n20000 );
    and g33726 ( n32509 , n32861 , n1187 );
    not g33727 ( n10576 , n38894 );
    not g33728 ( n13300 , n16075 );
    nor g33729 ( n25897 , n14707 , n29909 );
    and g33730 ( n24682 , n15796 , n35295 );
    nor g33731 ( n21831 , n34566 , n20337 );
    or g33732 ( n33076 , n6864 , n17888 );
    or g33733 ( n7865 , n5605 , n22776 );
    nor g33734 ( n39138 , n24216 , n34371 );
    or g33735 ( n20807 , n18868 , n41767 );
    not g33736 ( n7278 , n2076 );
    xnor g33737 ( n20258 , n26103 , n12800 );
    not g33738 ( n4226 , n5211 );
    and g33739 ( n38021 , n23912 , n15251 );
    or g33740 ( n25859 , n26876 , n36296 );
    and g33741 ( n1522 , n24814 , n8201 );
    nor g33742 ( n20150 , n19087 , n13995 );
    and g33743 ( n35210 , n19211 , n35475 );
    and g33744 ( n32348 , n37534 , n33499 );
    or g33745 ( n37571 , n8486 , n19836 );
    xnor g33746 ( n36334 , n42558 , n28863 );
    or g33747 ( n28331 , n18897 , n37647 );
    not g33748 ( n13296 , n36012 );
    or g33749 ( n29853 , n26834 , n12125 );
    not g33750 ( n2427 , n27476 );
    or g33751 ( n39067 , n32294 , n38090 );
    not g33752 ( n24692 , n29599 );
    or g33753 ( n11555 , n22544 , n28796 );
    not g33754 ( n25917 , n10779 );
    nor g33755 ( n28528 , n27543 , n8045 );
    not g33756 ( n20349 , n38114 );
    or g33757 ( n12921 , n19409 , n32688 );
    and g33758 ( n40671 , n40458 , n41828 );
    and g33759 ( n9817 , n17592 , n26355 );
    or g33760 ( n23428 , n1342 , n5894 );
    and g33761 ( n42533 , n1143 , n13309 );
    or g33762 ( n4536 , n5408 , n7626 );
    or g33763 ( n27850 , n12477 , n19104 );
    not g33764 ( n21902 , n2290 );
    or g33765 ( n34971 , n27008 , n22353 );
    xnor g33766 ( n8984 , n21935 , n15826 );
    not g33767 ( n881 , n4820 );
    and g33768 ( n38864 , n7456 , n22295 );
    xnor g33769 ( n1450 , n36009 , n27260 );
    or g33770 ( n36031 , n2259 , n37960 );
    or g33771 ( n15687 , n36913 , n11455 );
    not g33772 ( n36996 , n37335 );
    or g33773 ( n5433 , n18070 , n6672 );
    or g33774 ( n14059 , n15152 , n25622 );
    not g33775 ( n20529 , n36411 );
    and g33776 ( n10529 , n14445 , n2291 );
    nor g33777 ( n24206 , n5528 , n530 );
    xnor g33778 ( n12573 , n9535 , n18372 );
    not g33779 ( n41396 , n38603 );
    xnor g33780 ( n11337 , n19441 , n32840 );
    nor g33781 ( n5420 , n17049 , n33223 );
    or g33782 ( n28653 , n31490 , n24770 );
    not g33783 ( n2375 , n42803 );
    not g33784 ( n32178 , n8747 );
    or g33785 ( n1519 , n33518 , n23144 );
    or g33786 ( n3633 , n27302 , n8830 );
    and g33787 ( n37059 , n17246 , n18365 );
    not g33788 ( n22151 , n42409 );
    not g33789 ( n37335 , n17131 );
    nor g33790 ( n38767 , n27762 , n41750 );
    not g33791 ( n27818 , n30341 );
    or g33792 ( n41692 , n35382 , n5198 );
    or g33793 ( n3142 , n981 , n7426 );
    and g33794 ( n13797 , n28037 , n36544 );
    or g33795 ( n17534 , n7935 , n5338 );
    or g33796 ( n6200 , n3029 , n19419 );
    and g33797 ( n30919 , n13550 , n22059 );
    and g33798 ( n35868 , n41773 , n16637 );
    nor g33799 ( n22504 , n22086 , n29510 );
    and g33800 ( n3994 , n16572 , n27293 );
    not g33801 ( n40765 , n6676 );
    xnor g33802 ( n13363 , n6625 , n1820 );
    or g33803 ( n26677 , n35483 , n42125 );
    or g33804 ( n19093 , n39781 , n39098 );
    and g33805 ( n9709 , n25517 , n6528 );
    and g33806 ( n22502 , n22326 , n41731 );
    nor g33807 ( n23068 , n33783 , n29246 );
    or g33808 ( n19641 , n18622 , n1904 );
    not g33809 ( n19045 , n13042 );
    or g33810 ( n40548 , n18496 , n19596 );
    or g33811 ( n24491 , n14823 , n7042 );
    not g33812 ( n4877 , n42204 );
    not g33813 ( n31452 , n2529 );
    or g33814 ( n30695 , n23969 , n7340 );
    or g33815 ( n35670 , n29269 , n24771 );
    or g33816 ( n35219 , n6636 , n14532 );
    nor g33817 ( n17352 , n17672 , n36013 );
    not g33818 ( n1637 , n29154 );
    nor g33819 ( n18032 , n37800 , n27150 );
    xnor g33820 ( n31155 , n42898 , n19737 );
    and g33821 ( n18004 , n6036 , n32519 );
    not g33822 ( n31928 , n35307 );
    xnor g33823 ( n20045 , n7245 , n29961 );
    xnor g33824 ( n17201 , n27334 , n10925 );
    or g33825 ( n34126 , n23259 , n3045 );
    or g33826 ( n5700 , n22639 , n19497 );
    xnor g33827 ( n16490 , n38441 , n4760 );
    or g33828 ( n15720 , n7026 , n22201 );
    not g33829 ( n17104 , n32371 );
    or g33830 ( n39374 , n32683 , n25351 );
    nor g33831 ( n38200 , n23588 , n36552 );
    xnor g33832 ( n33695 , n16370 , n24550 );
    and g33833 ( n39413 , n10501 , n35357 );
    xnor g33834 ( n15510 , n6314 , n39925 );
    xnor g33835 ( n26773 , n2338 , n34819 );
    or g33836 ( n11913 , n22631 , n15692 );
    and g33837 ( n26686 , n8394 , n20841 );
    or g33838 ( n3716 , n34254 , n34459 );
    xnor g33839 ( n21250 , n15743 , n14707 );
    not g33840 ( n26407 , n39289 );
    xnor g33841 ( n29091 , n295 , n16553 );
    or g33842 ( n30980 , n31850 , n3754 );
    and g33843 ( n17388 , n14358 , n38549 );
    or g33844 ( n38054 , n17888 , n7176 );
    xnor g33845 ( n25612 , n39216 , n38879 );
    not g33846 ( n23563 , n13759 );
    or g33847 ( n41463 , n12777 , n39585 );
    and g33848 ( n14104 , n7524 , n32930 );
    and g33849 ( n19149 , n33622 , n35897 );
    and g33850 ( n26090 , n18034 , n25380 );
    or g33851 ( n27089 , n19969 , n11583 );
    or g33852 ( n38950 , n20218 , n25440 );
    and g33853 ( n9614 , n41095 , n40614 );
    not g33854 ( n29176 , n33280 );
    xnor g33855 ( n6653 , n25631 , n24452 );
    nor g33856 ( n14775 , n22625 , n34133 );
    xnor g33857 ( n25211 , n15089 , n33129 );
    or g33858 ( n37716 , n12713 , n35695 );
    or g33859 ( n31722 , n18585 , n35695 );
    and g33860 ( n10483 , n31349 , n36412 );
    or g33861 ( n1690 , n33451 , n8956 );
    nor g33862 ( n8830 , n20115 , n16256 );
    or g33863 ( n20014 , n7356 , n26185 );
    or g33864 ( n32578 , n40259 , n26319 );
    xnor g33865 ( n37410 , n36998 , n21900 );
    or g33866 ( n32579 , n15980 , n33328 );
    or g33867 ( n27959 , n12495 , n3316 );
    and g33868 ( n35417 , n27068 , n26037 );
    or g33869 ( n16880 , n23085 , n9644 );
    and g33870 ( n1215 , n37684 , n40119 );
    not g33871 ( n1588 , n5010 );
    or g33872 ( n13982 , n37119 , n5532 );
    and g33873 ( n7279 , n20007 , n16125 );
    xnor g33874 ( n22650 , n30768 , n34804 );
    or g33875 ( n7766 , n5455 , n9417 );
    or g33876 ( n37076 , n14622 , n21676 );
    xnor g33877 ( n18619 , n18530 , n16315 );
    or g33878 ( n21971 , n27545 , n31540 );
    xnor g33879 ( n21585 , n36998 , n28186 );
    or g33880 ( n22309 , n3281 , n9196 );
    xnor g33881 ( n3807 , n38350 , n15082 );
    or g33882 ( n19285 , n39483 , n35031 );
    not g33883 ( n26201 , n34922 );
    or g33884 ( n7583 , n11911 , n32878 );
    and g33885 ( n39470 , n36427 , n7686 );
    or g33886 ( n33965 , n31265 , n17303 );
    or g33887 ( n3895 , n26349 , n22031 );
    xnor g33888 ( n9594 , n33251 , n12770 );
    nor g33889 ( n32684 , n8810 , n42087 );
    not g33890 ( n18863 , n25531 );
    not g33891 ( n5353 , n22492 );
    nor g33892 ( n20658 , n37582 , n11494 );
    or g33893 ( n33125 , n4823 , n27406 );
    xnor g33894 ( n3168 , n27704 , n25865 );
    or g33895 ( n26020 , n2464 , n25303 );
    and g33896 ( n29762 , n13459 , n2424 );
    and g33897 ( n42646 , n12894 , n26271 );
    not g33898 ( n35035 , n42204 );
    nor g33899 ( n35559 , n36117 , n4816 );
    nor g33900 ( n18035 , n17193 , n27669 );
    xnor g33901 ( n27984 , n16201 , n4418 );
    or g33902 ( n23789 , n26542 , n2404 );
    and g33903 ( n39919 , n26571 , n16698 );
    or g33904 ( n10947 , n27376 , n15895 );
    xnor g33905 ( n29838 , n26579 , n3439 );
    or g33906 ( n5399 , n27956 , n2299 );
    not g33907 ( n21367 , n40932 );
    and g33908 ( n134 , n2376 , n40880 );
    and g33909 ( n6755 , n31099 , n36865 );
    or g33910 ( n32871 , n41346 , n20446 );
    or g33911 ( n1686 , n16223 , n36649 );
    and g33912 ( n8455 , n25908 , n28237 );
    or g33913 ( n40113 , n31302 , n3154 );
    xnor g33914 ( n4339 , n4127 , n42389 );
    and g33915 ( n5599 , n14792 , n9011 );
    and g33916 ( n3518 , n41101 , n17023 );
    nor g33917 ( n22475 , n1990 , n18314 );
    or g33918 ( n35822 , n18165 , n24882 );
    and g33919 ( n29121 , n16506 , n27283 );
    not g33920 ( n40752 , n39208 );
    or g33921 ( n35585 , n22920 , n33082 );
    xnor g33922 ( n27896 , n37403 , n13985 );
    and g33923 ( n32499 , n35727 , n37547 );
    and g33924 ( n22004 , n13557 , n24076 );
    not g33925 ( n2513 , n18800 );
    and g33926 ( n18525 , n5676 , n36572 );
    nor g33927 ( n12408 , n1765 , n5079 );
    or g33928 ( n25748 , n8004 , n12648 );
    not g33929 ( n27148 , n31510 );
    nor g33930 ( n34002 , n25145 , n28255 );
    or g33931 ( n32059 , n38959 , n10557 );
    not g33932 ( n13336 , n24273 );
    and g33933 ( n4169 , n11543 , n28815 );
    xnor g33934 ( n10271 , n9775 , n27337 );
    nor g33935 ( n13551 , n38242 , n21671 );
    not g33936 ( n29056 , n11525 );
    nor g33937 ( n17976 , n39645 , n34011 );
    and g33938 ( n39399 , n25599 , n36064 );
    nor g33939 ( n19374 , n5086 , n39238 );
    or g33940 ( n20128 , n5991 , n17212 );
    not g33941 ( n14520 , n24786 );
    not g33942 ( n9883 , n20544 );
    xnor g33943 ( n37921 , n11702 , n7569 );
    xnor g33944 ( n1108 , n36998 , n21164 );
    and g33945 ( n7856 , n35931 , n22409 );
    and g33946 ( n18712 , n37091 , n32659 );
    and g33947 ( n9000 , n25658 , n5164 );
    and g33948 ( n10406 , n37631 , n21329 );
    or g33949 ( n30330 , n15283 , n23228 );
    nor g33950 ( n4812 , n27524 , n23989 );
    or g33951 ( n35446 , n41887 , n33926 );
    and g33952 ( n20001 , n32757 , n27182 );
    or g33953 ( n8925 , n42870 , n16359 );
    or g33954 ( n15995 , n37516 , n29201 );
    and g33955 ( n41682 , n19990 , n27520 );
    or g33956 ( n41028 , n6278 , n14155 );
    not g33957 ( n30438 , n33807 );
    nor g33958 ( n2767 , n6823 , n14456 );
    or g33959 ( n39816 , n11678 , n36376 );
    xnor g33960 ( n7285 , n36364 , n39193 );
    nor g33961 ( n33454 , n30189 , n12683 );
    or g33962 ( n963 , n2095 , n24355 );
    nor g33963 ( n8751 , n25668 , n29682 );
    nor g33964 ( n22206 , n167 , n14513 );
    or g33965 ( n40677 , n41534 , n42299 );
    or g33966 ( n31968 , n31525 , n29149 );
    or g33967 ( n38651 , n6138 , n19632 );
    xnor g33968 ( n31385 , n38749 , n33985 );
    or g33969 ( n2914 , n9719 , n40482 );
    not g33970 ( n38274 , n8514 );
    and g33971 ( n15401 , n4047 , n6777 );
    not g33972 ( n4553 , n4359 );
    or g33973 ( n33060 , n5262 , n12334 );
    or g33974 ( n33800 , n37802 , n10145 );
    or g33975 ( n26365 , n32256 , n42020 );
    nor g33976 ( n18179 , n10812 , n29401 );
    or g33977 ( n25465 , n41136 , n20296 );
    and g33978 ( n30521 , n5702 , n40767 );
    xnor g33979 ( n7741 , n20548 , n33036 );
    or g33980 ( n6523 , n25646 , n20260 );
    not g33981 ( n35098 , n39188 );
    and g33982 ( n7504 , n31912 , n19743 );
    xnor g33983 ( n718 , n13677 , n1418 );
    not g33984 ( n26394 , n5675 );
    xnor g33985 ( n2247 , n7943 , n41568 );
    or g33986 ( n14842 , n41131 , n41207 );
    or g33987 ( n34488 , n31641 , n41295 );
    and g33988 ( n8363 , n39265 , n34982 );
    xnor g33989 ( n5851 , n39757 , n34172 );
    or g33990 ( n5066 , n18165 , n21123 );
    and g33991 ( n13511 , n19741 , n18351 );
    nor g33992 ( n19389 , n21741 , n21262 );
    or g33993 ( n37228 , n12482 , n36052 );
    or g33994 ( n26771 , n5497 , n1385 );
    or g33995 ( n28102 , n33057 , n34010 );
    or g33996 ( n23697 , n12794 , n13391 );
    and g33997 ( n21341 , n2393 , n24821 );
    not g33998 ( n1292 , n28517 );
    and g33999 ( n41404 , n18855 , n29225 );
    or g34000 ( n24600 , n40431 , n23489 );
    or g34001 ( n36538 , n16284 , n41431 );
    and g34002 ( n4639 , n41482 , n25103 );
    or g34003 ( n20585 , n24031 , n12129 );
    or g34004 ( n3002 , n18798 , n8541 );
    or g34005 ( n14936 , n3573 , n8945 );
    or g34006 ( n12617 , n27267 , n7265 );
    xnor g34007 ( n27693 , n24814 , n8201 );
    or g34008 ( n17565 , n11340 , n8178 );
    xnor g34009 ( n42735 , n41587 , n3191 );
    and g34010 ( n37871 , n37482 , n2915 );
    and g34011 ( n9413 , n4123 , n35744 );
    and g34012 ( n34119 , n6910 , n18733 );
    xnor g34013 ( n31529 , n35650 , n31512 );
    not g34014 ( n277 , n28798 );
    not g34015 ( n20998 , n31578 );
    nor g34016 ( n6280 , n27644 , n16484 );
    xnor g34017 ( n12100 , n6800 , n31611 );
    or g34018 ( n40727 , n25627 , n32244 );
    not g34019 ( n16076 , n36488 );
    or g34020 ( n19974 , n10915 , n40475 );
    or g34021 ( n17189 , n41631 , n15268 );
    not g34022 ( n2668 , n26368 );
    or g34023 ( n1754 , n18853 , n39924 );
    and g34024 ( n15045 , n15499 , n22856 );
    nor g34025 ( n11016 , n6715 , n35898 );
    not g34026 ( n25475 , n1130 );
    xnor g34027 ( n32981 , n25426 , n41136 );
    nor g34028 ( n42033 , n17744 , n4883 );
    or g34029 ( n32238 , n2105 , n24923 );
    and g34030 ( n13108 , n26967 , n9267 );
    not g34031 ( n24291 , n10008 );
    and g34032 ( n11643 , n39770 , n8720 );
    and g34033 ( n4766 , n32723 , n31488 );
    nor g34034 ( n23922 , n5964 , n33522 );
    and g34035 ( n14200 , n24345 , n8321 );
    and g34036 ( n7152 , n30315 , n25941 );
    or g34037 ( n12542 , n10220 , n33691 );
    not g34038 ( n12754 , n27050 );
    or g34039 ( n34860 , n2507 , n10404 );
    xnor g34040 ( n10135 , n16745 , n4598 );
    and g34041 ( n25091 , n25188 , n31117 );
    not g34042 ( n5110 , n2495 );
    nor g34043 ( n8788 , n30742 , n16497 );
    and g34044 ( n1694 , n39871 , n8754 );
    or g34045 ( n15072 , n19186 , n6154 );
    or g34046 ( n11940 , n31366 , n19702 );
    not g34047 ( n32632 , n42550 );
    xnor g34048 ( n21863 , n39295 , n26187 );
    or g34049 ( n4635 , n35717 , n11026 );
    or g34050 ( n32601 , n23261 , n10638 );
    and g34051 ( n41148 , n21120 , n5600 );
    not g34052 ( n40141 , n25978 );
    xnor g34053 ( n15576 , n20086 , n6693 );
    and g34054 ( n2880 , n20053 , n20977 );
    or g34055 ( n26962 , n21779 , n5881 );
    nor g34056 ( n22592 , n8494 , n24497 );
    or g34057 ( n26209 , n38436 , n4384 );
    not g34058 ( n20496 , n9256 );
    and g34059 ( n5671 , n39798 , n35161 );
    or g34060 ( n5238 , n2972 , n7647 );
    not g34061 ( n42192 , n4047 );
    or g34062 ( n37812 , n15809 , n22920 );
    not g34063 ( n13236 , n26620 );
    or g34064 ( n13806 , n27537 , n34962 );
    xnor g34065 ( n7937 , n24278 , n5628 );
    nor g34066 ( n39022 , n5605 , n25280 );
    or g34067 ( n33739 , n942 , n11814 );
    or g34068 ( n22458 , n18647 , n30442 );
    or g34069 ( n5119 , n30085 , n27127 );
    and g34070 ( n30926 , n3266 , n27422 );
    xnor g34071 ( n34437 , n29718 , n3929 );
    or g34072 ( n42644 , n25588 , n28113 );
    not g34073 ( n14105 , n24023 );
    and g34074 ( n39208 , n41805 , n25291 );
    not g34075 ( n39897 , n18998 );
    xnor g34076 ( n27981 , n38035 , n22757 );
    xnor g34077 ( n18599 , n24093 , n7537 );
    and g34078 ( n1280 , n15068 , n28767 );
    and g34079 ( n40607 , n17400 , n42147 );
    and g34080 ( n11008 , n24364 , n23461 );
    not g34081 ( n35255 , n4424 );
    or g34082 ( n13376 , n7196 , n17022 );
    xnor g34083 ( n13743 , n33570 , n13051 );
    or g34084 ( n24631 , n25945 , n22379 );
    or g34085 ( n6390 , n1292 , n30080 );
    nor g34086 ( n28191 , n34565 , n5599 );
    or g34087 ( n1142 , n21815 , n42517 );
    or g34088 ( n4225 , n20893 , n20969 );
    and g34089 ( n9097 , n9002 , n26388 );
    and g34090 ( n2285 , n38607 , n42571 );
    nor g34091 ( n9364 , n4084 , n2867 );
    xnor g34092 ( n106 , n12190 , n26132 );
    nor g34093 ( n23620 , n33981 , n31979 );
    nor g34094 ( n13228 , n36337 , n20392 );
    xnor g34095 ( n26753 , n26683 , n4168 );
    and g34096 ( n17174 , n36910 , n35113 );
    or g34097 ( n14678 , n42076 , n41605 );
    and g34098 ( n15863 , n14336 , n15612 );
    or g34099 ( n35844 , n18627 , n37155 );
    nor g34100 ( n35412 , n27733 , n15044 );
    not g34101 ( n7338 , n40514 );
    and g34102 ( n29660 , n14189 , n28094 );
    not g34103 ( n31294 , n29711 );
    and g34104 ( n5864 , n21136 , n32129 );
    nor g34105 ( n14535 , n17120 , n29173 );
    or g34106 ( n15306 , n30017 , n41374 );
    and g34107 ( n18053 , n40632 , n42542 );
    nor g34108 ( n21496 , n40067 , n30821 );
    xnor g34109 ( n11394 , n25927 , n31558 );
    nor g34110 ( n8726 , n27960 , n12845 );
    and g34111 ( n34241 , n15649 , n22965 );
    xnor g34112 ( n31353 , n453 , n28625 );
    or g34113 ( n4910 , n36852 , n36844 );
    not g34114 ( n41715 , n19014 );
    or g34115 ( n10343 , n27711 , n8658 );
    nor g34116 ( n16625 , n25660 , n38975 );
    nor g34117 ( n36172 , n35508 , n23482 );
    or g34118 ( n24081 , n17827 , n2870 );
    or g34119 ( n42854 , n41261 , n39203 );
    xnor g34120 ( n13770 , n10558 , n17065 );
    and g34121 ( n19525 , n42366 , n4420 );
    nor g34122 ( n10355 , n33938 , n16326 );
    not g34123 ( n7891 , n28809 );
    and g34124 ( n19986 , n29333 , n41105 );
    and g34125 ( n5663 , n6409 , n15459 );
    or g34126 ( n19684 , n24374 , n41869 );
    and g34127 ( n18668 , n3903 , n21861 );
    or g34128 ( n6600 , n23268 , n1351 );
    not g34129 ( n22726 , n27086 );
    and g34130 ( n14271 , n255 , n1751 );
    not g34131 ( n20437 , n35547 );
    or g34132 ( n31171 , n12543 , n22797 );
    not g34133 ( n3315 , n31519 );
    xnor g34134 ( n27265 , n39760 , n24037 );
    or g34135 ( n4780 , n20733 , n28289 );
    and g34136 ( n8907 , n3445 , n13037 );
    not g34137 ( n21703 , n28177 );
    not g34138 ( n7611 , n29708 );
    xnor g34139 ( n8797 , n5593 , n14400 );
    xnor g34140 ( n23159 , n24218 , n24123 );
    and g34141 ( n37296 , n5384 , n31577 );
    and g34142 ( n30282 , n12520 , n22847 );
    not g34143 ( n17756 , n30016 );
    nor g34144 ( n17355 , n10390 , n27291 );
    xnor g34145 ( n25554 , n7980 , n8180 );
    or g34146 ( n16346 , n19625 , n39997 );
    and g34147 ( n28220 , n2396 , n31486 );
    or g34148 ( n27563 , n29803 , n34718 );
    nor g34149 ( n9490 , n28695 , n22595 );
    or g34150 ( n33697 , n9937 , n14784 );
    or g34151 ( n18374 , n36576 , n12129 );
    or g34152 ( n8877 , n23509 , n6297 );
    or g34153 ( n16300 , n10967 , n35467 );
    and g34154 ( n25437 , n25411 , n30384 );
    nor g34155 ( n17836 , n25588 , n22948 );
    nor g34156 ( n12813 , n36539 , n20767 );
    or g34157 ( n35827 , n18775 , n33066 );
    or g34158 ( n13030 , n40259 , n18373 );
    nor g34159 ( n1074 , n6300 , n17705 );
    and g34160 ( n8212 , n14652 , n39513 );
    or g34161 ( n25734 , n34404 , n18031 );
    nor g34162 ( n4637 , n15070 , n42020 );
    nor g34163 ( n37090 , n25421 , n6443 );
    or g34164 ( n4064 , n15584 , n35227 );
    or g34165 ( n10500 , n30657 , n39756 );
    or g34166 ( n3364 , n21330 , n31068 );
    or g34167 ( n3662 , n9415 , n21019 );
    xnor g34168 ( n36721 , n12274 , n7588 );
    or g34169 ( n7407 , n9734 , n24279 );
    or g34170 ( n28716 , n20243 , n26719 );
    not g34171 ( n39218 , n34185 );
    xnor g34172 ( n24554 , n7937 , n32304 );
    and g34173 ( n35197 , n27797 , n25013 );
    or g34174 ( n21729 , n26156 , n21552 );
    or g34175 ( n29019 , n27729 , n37627 );
    and g34176 ( n39515 , n19276 , n1676 );
    not g34177 ( n12543 , n24103 );
    or g34178 ( n42589 , n14442 , n12896 );
    and g34179 ( n4323 , n3984 , n4125 );
    nor g34180 ( n34496 , n7567 , n25743 );
    not g34181 ( n20468 , n32444 );
    or g34182 ( n27757 , n10019 , n8432 );
    or g34183 ( n8114 , n39526 , n25742 );
    nor g34184 ( n40133 , n23612 , n37366 );
    nor g34185 ( n6181 , n12344 , n22542 );
    and g34186 ( n39617 , n11356 , n19688 );
    and g34187 ( n9974 , n33715 , n12135 );
    or g34188 ( n26674 , n5211 , n25751 );
    or g34189 ( n17077 , n41286 , n2597 );
    or g34190 ( n15833 , n7801 , n6730 );
    and g34191 ( n11317 , n32916 , n36969 );
    not g34192 ( n26670 , n39642 );
    nor g34193 ( n3078 , n24951 , n24969 );
    nor g34194 ( n14737 , n28691 , n9076 );
    not g34195 ( n28253 , n19531 );
    nor g34196 ( n17540 , n38738 , n41593 );
    and g34197 ( n42289 , n28387 , n23937 );
    or g34198 ( n34299 , n24358 , n23199 );
    and g34199 ( n13013 , n32006 , n18206 );
    and g34200 ( n6156 , n14537 , n11729 );
    and g34201 ( n11674 , n15680 , n2700 );
    and g34202 ( n20337 , n19388 , n5662 );
    not g34203 ( n785 , n32558 );
    and g34204 ( n21983 , n18526 , n26878 );
    and g34205 ( n21283 , n41174 , n6157 );
    not g34206 ( n8504 , n37760 );
    or g34207 ( n10366 , n34448 , n41079 );
    and g34208 ( n34974 , n41599 , n24342 );
    or g34209 ( n22261 , n12909 , n38219 );
    and g34210 ( n21151 , n15916 , n14322 );
    nor g34211 ( n31838 , n7817 , n2196 );
    or g34212 ( n15670 , n11459 , n8087 );
    not g34213 ( n37667 , n36216 );
    not g34214 ( n26689 , n16987 );
    or g34215 ( n17816 , n5258 , n5079 );
    and g34216 ( n12684 , n35664 , n36692 );
    or g34217 ( n23339 , n37671 , n33462 );
    or g34218 ( n30384 , n31542 , n41809 );
    or g34219 ( n1245 , n26507 , n520 );
    and g34220 ( n23674 , n19891 , n25393 );
    or g34221 ( n24489 , n7003 , n6195 );
    nor g34222 ( n28788 , n34292 , n29343 );
    xnor g34223 ( n34789 , n21534 , n26250 );
    not g34224 ( n4271 , n36661 );
    or g34225 ( n24921 , n28098 , n21767 );
    or g34226 ( n36855 , n12910 , n13694 );
    not g34227 ( n1208 , n33801 );
    or g34228 ( n29205 , n40624 , n8283 );
    xnor g34229 ( n16364 , n38314 , n5313 );
    xnor g34230 ( n11885 , n19305 , n4985 );
    or g34231 ( n14118 , n8494 , n36091 );
    and g34232 ( n4052 , n42250 , n38726 );
    and g34233 ( n14688 , n27129 , n5374 );
    or g34234 ( n33822 , n12071 , n256 );
    or g34235 ( n525 , n14481 , n40816 );
    or g34236 ( n18409 , n20138 , n30711 );
    not g34237 ( n16500 , n7916 );
    or g34238 ( n17128 , n21131 , n18494 );
    and g34239 ( n15946 , n35315 , n29641 );
    not g34240 ( n42554 , n41623 );
    or g34241 ( n14498 , n20283 , n34972 );
    or g34242 ( n19462 , n2765 , n11708 );
    xnor g34243 ( n30668 , n20604 , n5605 );
    or g34244 ( n42673 , n40462 , n39171 );
    not g34245 ( n38704 , n19326 );
    not g34246 ( n1917 , n11682 );
    xnor g34247 ( n39115 , n8457 , n36629 );
    or g34248 ( n42413 , n8669 , n16170 );
    nor g34249 ( n1871 , n14471 , n42308 );
    and g34250 ( n19840 , n14239 , n13036 );
    xnor g34251 ( n17178 , n11436 , n1436 );
    xnor g34252 ( n14984 , n34731 , n14126 );
    or g34253 ( n35475 , n41907 , n27515 );
    or g34254 ( n1773 , n41915 , n33681 );
    xnor g34255 ( n40284 , n13160 , n4028 );
    not g34256 ( n12724 , n24106 );
    and g34257 ( n23590 , n12589 , n39181 );
    or g34258 ( n14060 , n5037 , n10530 );
    or g34259 ( n353 , n38256 , n24197 );
    and g34260 ( n39366 , n23308 , n31348 );
    and g34261 ( n33635 , n28893 , n26473 );
    or g34262 ( n42468 , n35040 , n34085 );
    or g34263 ( n2008 , n35429 , n37633 );
    and g34264 ( n31176 , n15361 , n37846 );
    not g34265 ( n24713 , n29967 );
    nor g34266 ( n7232 , n33981 , n42321 );
    not g34267 ( n4743 , n25108 );
    or g34268 ( n38289 , n19871 , n10797 );
    and g34269 ( n7322 , n25381 , n20462 );
    and g34270 ( n42732 , n25112 , n17524 );
    or g34271 ( n10190 , n3954 , n39334 );
    or g34272 ( n18189 , n12366 , n26789 );
    xnor g34273 ( n41363 , n34795 , n17760 );
    and g34274 ( n2515 , n29905 , n20715 );
    not g34275 ( n29764 , n27824 );
    and g34276 ( n39557 , n7538 , n2828 );
    and g34277 ( n41493 , n4741 , n13016 );
    nor g34278 ( n15959 , n34341 , n26029 );
    not g34279 ( n2789 , n23831 );
    nor g34280 ( n11246 , n15717 , n1273 );
    xnor g34281 ( n4557 , n9941 , n41534 );
    not g34282 ( n19651 , n36762 );
    or g34283 ( n15231 , n11656 , n3133 );
    nor g34284 ( n41622 , n10601 , n1895 );
    and g34285 ( n11339 , n26145 , n13156 );
    or g34286 ( n22449 , n218 , n23583 );
    xnor g34287 ( n27418 , n6625 , n41678 );
    or g34288 ( n41417 , n12112 , n10626 );
    and g34289 ( n15130 , n20539 , n14893 );
    or g34290 ( n702 , n13689 , n1292 );
    nor g34291 ( n11771 , n17330 , n41042 );
    nor g34292 ( n16533 , n17724 , n33179 );
    nor g34293 ( n42862 , n41408 , n31548 );
    or g34294 ( n28644 , n10674 , n16597 );
    nor g34295 ( n1910 , n30396 , n5268 );
    and g34296 ( n18184 , n28742 , n9158 );
    or g34297 ( n20752 , n40313 , n36962 );
    or g34298 ( n2546 , n15666 , n4402 );
    or g34299 ( n7225 , n2296 , n41399 );
    or g34300 ( n36632 , n23214 , n39724 );
    and g34301 ( n2666 , n8791 , n31508 );
    nor g34302 ( n5928 , n15429 , n42634 );
    nor g34303 ( n18291 , n18951 , n20158 );
    and g34304 ( n7682 , n11644 , n31908 );
    nor g34305 ( n42859 , n455 , n18517 );
    xnor g34306 ( n11247 , n3065 , n31802 );
    or g34307 ( n5158 , n22578 , n41274 );
    or g34308 ( n25687 , n9372 , n30679 );
    xnor g34309 ( n28849 , n37908 , n31212 );
    and g34310 ( n33638 , n33158 , n32448 );
    or g34311 ( n5156 , n34391 , n7254 );
    xnor g34312 ( n11691 , n7836 , n18349 );
    or g34313 ( n8744 , n23859 , n32608 );
    not g34314 ( n34628 , n1681 );
    and g34315 ( n1687 , n1213 , n33517 );
    nor g34316 ( n16843 , n30743 , n33728 );
    or g34317 ( n37426 , n6003 , n5212 );
    and g34318 ( n15445 , n3067 , n40112 );
    and g34319 ( n27871 , n17123 , n11934 );
    and g34320 ( n13416 , n6091 , n11421 );
    or g34321 ( n39560 , n147 , n21466 );
    xnor g34322 ( n13120 , n33310 , n14116 );
    and g34323 ( n42563 , n8643 , n234 );
    and g34324 ( n12574 , n19415 , n23579 );
    and g34325 ( n39951 , n29827 , n38131 );
    xnor g34326 ( n27793 , n11436 , n5563 );
    xnor g34327 ( n21003 , n1863 , n8083 );
    not g34328 ( n17377 , n3334 );
    not g34329 ( n38964 , n1721 );
    xnor g34330 ( n40992 , n41515 , n18758 );
    or g34331 ( n37601 , n15020 , n13584 );
    or g34332 ( n41379 , n30192 , n6029 );
    nor g34333 ( n40636 , n27572 , n38313 );
    or g34334 ( n29905 , n25589 , n15957 );
    and g34335 ( n38689 , n8638 , n10813 );
    nor g34336 ( n970 , n9272 , n42691 );
    nor g34337 ( n7441 , n27762 , n14586 );
    xnor g34338 ( n12892 , n34105 , n29477 );
    and g34339 ( n28186 , n29335 , n42594 );
    xnor g34340 ( n32936 , n25789 , n32277 );
    xnor g34341 ( n30930 , n15590 , n23547 );
    not g34342 ( n17170 , n18901 );
    and g34343 ( n42419 , n15102 , n5569 );
    nor g34344 ( n23988 , n2722 , n35807 );
    nor g34345 ( n22388 , n15070 , n41639 );
    xnor g34346 ( n5404 , n37709 , n12306 );
    not g34347 ( n10993 , n4045 );
    not g34348 ( n907 , n12425 );
    or g34349 ( n18001 , n5125 , n2576 );
    nor g34350 ( n38669 , n38712 , n19919 );
    or g34351 ( n13723 , n10986 , n42535 );
    and g34352 ( n5780 , n23106 , n35470 );
    or g34353 ( n6206 , n15485 , n41069 );
    or g34354 ( n4259 , n34584 , n28311 );
    xnor g34355 ( n17544 , n32583 , n5922 );
    and g34356 ( n13190 , n35318 , n1672 );
    nor g34357 ( n19413 , n1197 , n19260 );
    or g34358 ( n35015 , n8022 , n4036 );
    not g34359 ( n9084 , n41357 );
    not g34360 ( n27161 , n23219 );
    or g34361 ( n33257 , n6041 , n40689 );
    xnor g34362 ( n1336 , n23873 , n11777 );
    nor g34363 ( n15758 , n21476 , n3598 );
    not g34364 ( n22972 , n22956 );
    or g34365 ( n18958 , n20778 , n34225 );
    and g34366 ( n7255 , n12697 , n12933 );
    not g34367 ( n37969 , n9331 );
    or g34368 ( n7910 , n41086 , n12002 );
    xnor g34369 ( n40312 , n21097 , n24842 );
    nor g34370 ( n15594 , n10595 , n4483 );
    or g34371 ( n41840 , n20164 , n24033 );
    not g34372 ( n37403 , n12514 );
    or g34373 ( n5145 , n13366 , n32545 );
    not g34374 ( n3817 , n34933 );
    and g34375 ( n37756 , n25397 , n19505 );
    not g34376 ( n35901 , n6674 );
    or g34377 ( n3658 , n41891 , n34177 );
    or g34378 ( n10055 , n36967 , n42491 );
    and g34379 ( n37182 , n8124 , n10660 );
    xnor g34380 ( n16814 , n24892 , n36107 );
    not g34381 ( n10057 , n19914 );
    or g34382 ( n39389 , n35431 , n24371 );
    and g34383 ( n34085 , n32423 , n33402 );
    and g34384 ( n18514 , n17019 , n29737 );
    not g34385 ( n33044 , n34206 );
    or g34386 ( n19715 , n41328 , n12500 );
    or g34387 ( n21949 , n26916 , n37728 );
    and g34388 ( n197 , n19900 , n10316 );
    and g34389 ( n29811 , n11363 , n5177 );
    or g34390 ( n21720 , n9137 , n586 );
    or g34391 ( n15135 , n34994 , n42787 );
    xnor g34392 ( n30138 , n12386 , n3152 );
    not g34393 ( n21862 , n16495 );
    or g34394 ( n6416 , n7361 , n19955 );
    or g34395 ( n23393 , n25623 , n25482 );
    or g34396 ( n16931 , n10592 , n10620 );
    or g34397 ( n18609 , n14457 , n4276 );
    xnor g34398 ( n23090 , n24210 , n2436 );
    nor g34399 ( n34639 , n37241 , n24310 );
    or g34400 ( n36502 , n6004 , n32607 );
    and g34401 ( n19805 , n21570 , n24047 );
    or g34402 ( n25272 , n42706 , n28848 );
    and g34403 ( n35672 , n2342 , n4458 );
    or g34404 ( n25362 , n26162 , n14478 );
    not g34405 ( n14583 , n42024 );
    and g34406 ( n17009 , n37394 , n35826 );
    and g34407 ( n8601 , n22839 , n6239 );
    nor g34408 ( n19455 , n41179 , n41576 );
    nor g34409 ( n17797 , n25588 , n42280 );
    not g34410 ( n3801 , n5254 );
    or g34411 ( n14251 , n23040 , n16166 );
    not g34412 ( n25299 , n21675 );
    and g34413 ( n19005 , n1532 , n23785 );
    or g34414 ( n38830 , n17149 , n26922 );
    xnor g34415 ( n9157 , n27741 , n31859 );
    or g34416 ( n26894 , n16967 , n32811 );
    not g34417 ( n3209 , n14656 );
    or g34418 ( n1388 , n38735 , n9387 );
    not g34419 ( n15796 , n21998 );
    xnor g34420 ( n16055 , n28225 , n21812 );
    and g34421 ( n670 , n42643 , n12154 );
    or g34422 ( n5827 , n31401 , n25407 );
    and g34423 ( n32743 , n21139 , n20470 );
    not g34424 ( n26409 , n28057 );
    or g34425 ( n37463 , n23292 , n23466 );
    or g34426 ( n22496 , n36368 , n34267 );
    not g34427 ( n7737 , n30555 );
    or g34428 ( n27347 , n19969 , n40933 );
    or g34429 ( n21196 , n37664 , n39033 );
    and g34430 ( n3473 , n11856 , n39737 );
    or g34431 ( n34729 , n21128 , n36836 );
    and g34432 ( n41102 , n10567 , n3871 );
    or g34433 ( n4996 , n42220 , n20916 );
    nor g34434 ( n27841 , n31135 , n15813 );
    or g34435 ( n9739 , n22833 , n42437 );
    nor g34436 ( n38327 , n9796 , n18412 );
    nor g34437 ( n17477 , n3769 , n37683 );
    or g34438 ( n35582 , n32044 , n42425 );
    nor g34439 ( n28960 , n5896 , n1610 );
    or g34440 ( n7745 , n11346 , n3528 );
    or g34441 ( n9726 , n4836 , n2366 );
    not g34442 ( n19832 , n3361 );
    or g34443 ( n36013 , n42646 , n34134 );
    or g34444 ( n8113 , n12700 , n28789 );
    xnor g34445 ( n20543 , n8906 , n22923 );
    nor g34446 ( n42034 , n589 , n328 );
    not g34447 ( n10601 , n19508 );
    not g34448 ( n5615 , n282 );
    not g34449 ( n21840 , n14763 );
    and g34450 ( n1716 , n6056 , n7051 );
    xnor g34451 ( n35733 , n25884 , n20497 );
    and g34452 ( n18877 , n26723 , n25518 );
    or g34453 ( n8598 , n25146 , n1735 );
    or g34454 ( n27141 , n21537 , n30393 );
    not g34455 ( n69 , n13159 );
    nor g34456 ( n5680 , n36117 , n31098 );
    or g34457 ( n22612 , n21347 , n36368 );
    and g34458 ( n19273 , n7112 , n12609 );
    not g34459 ( n20513 , n34880 );
    not g34460 ( n26419 , n1439 );
    or g34461 ( n30589 , n20633 , n23558 );
    xnor g34462 ( n42277 , n31099 , n29407 );
    or g34463 ( n35494 , n27533 , n7953 );
    or g34464 ( n5374 , n24168 , n19679 );
    or g34465 ( n39737 , n24177 , n22110 );
    or g34466 ( n16042 , n20428 , n8302 );
    or g34467 ( n36610 , n38689 , n24437 );
    not g34468 ( n1986 , n39766 );
    not g34469 ( n1244 , n4313 );
    and g34470 ( n24677 , n35278 , n9924 );
    nor g34471 ( n27120 , n15261 , n41605 );
    or g34472 ( n13068 , n33330 , n19632 );
    xnor g34473 ( n17395 , n34875 , n6220 );
    or g34474 ( n42415 , n25602 , n22115 );
    or g34475 ( n37573 , n3636 , n410 );
    and g34476 ( n32274 , n14834 , n9890 );
    or g34477 ( n21522 , n5647 , n3715 );
    or g34478 ( n13060 , n34485 , n6039 );
    xnor g34479 ( n27403 , n21609 , n39916 );
    and g34480 ( n3853 , n5325 , n2788 );
    or g34481 ( n19846 , n42600 , n4730 );
    and g34482 ( n23 , n6608 , n28521 );
    or g34483 ( n41398 , n22619 , n33482 );
    xnor g34484 ( n20581 , n20791 , n27460 );
    xnor g34485 ( n26275 , n35727 , n11727 );
    nor g34486 ( n6851 , n4469 , n41813 );
    nor g34487 ( n9411 , n21201 , n38067 );
    not g34488 ( n30066 , n34258 );
    or g34489 ( n24092 , n972 , n6141 );
    or g34490 ( n10379 , n4161 , n42769 );
    nor g34491 ( n39043 , n17668 , n32524 );
    or g34492 ( n15214 , n41819 , n27803 );
    nor g34493 ( n15528 , n13306 , n8103 );
    and g34494 ( n8209 , n40063 , n34514 );
    xnor g34495 ( n23179 , n14377 , n22487 );
    or g34496 ( n26248 , n8212 , n3947 );
    or g34497 ( n32647 , n12495 , n34726 );
    xnor g34498 ( n18506 , n25043 , n41594 );
    or g34499 ( n27225 , n3977 , n40157 );
    or g34500 ( n42512 , n31738 , n26888 );
    or g34501 ( n4114 , n27553 , n2565 );
    and g34502 ( n25540 , n30699 , n26822 );
    or g34503 ( n24422 , n31999 , n28058 );
    nor g34504 ( n32188 , n17393 , n16757 );
    nor g34505 ( n12413 , n14471 , n38538 );
    not g34506 ( n952 , n6894 );
    xnor g34507 ( n22179 , n17439 , n6877 );
    or g34508 ( n16665 , n42908 , n30822 );
    nor g34509 ( n11936 , n14989 , n31438 );
    or g34510 ( n22029 , n27663 , n3406 );
    nor g34511 ( n9696 , n2080 , n32860 );
    or g34512 ( n13850 , n28725 , n2601 );
    nor g34513 ( n39358 , n38730 , n19320 );
    or g34514 ( n35916 , n3783 , n34422 );
    or g34515 ( n40433 , n29664 , n35557 );
    nor g34516 ( n35373 , n33662 , n34450 );
    or g34517 ( n1346 , n36365 , n24910 );
    xnor g34518 ( n27114 , n25556 , n11207 );
    and g34519 ( n16912 , n27214 , n33753 );
    and g34520 ( n24299 , n39795 , n27336 );
    or g34521 ( n15870 , n41996 , n19781 );
    or g34522 ( n11602 , n30065 , n33103 );
    or g34523 ( n10371 , n27375 , n2675 );
    and g34524 ( n5868 , n32143 , n4764 );
    xnor g34525 ( n8597 , n542 , n41999 );
    xnor g34526 ( n37909 , n7881 , n11634 );
    xnor g34527 ( n18204 , n5144 , n9609 );
    xnor g34528 ( n31273 , n31099 , n22832 );
    nor g34529 ( n8731 , n19471 , n7623 );
    not g34530 ( n32119 , n3137 );
    and g34531 ( n32241 , n11563 , n19199 );
    and g34532 ( n41283 , n10989 , n447 );
    or g34533 ( n41135 , n40824 , n2699 );
    or g34534 ( n28645 , n20996 , n29660 );
    or g34535 ( n40899 , n23569 , n12419 );
    or g34536 ( n25922 , n15545 , n29980 );
    not g34537 ( n9020 , n38545 );
    or g34538 ( n33516 , n22513 , n15932 );
    xnor g34539 ( n12576 , n24695 , n643 );
    xnor g34540 ( n3857 , n13415 , n13065 );
    nor g34541 ( n23250 , n8494 , n5181 );
    and g34542 ( n42018 , n8816 , n32484 );
    nor g34543 ( n37689 , n24180 , n21722 );
    or g34544 ( n12901 , n20485 , n10373 );
    and g34545 ( n37972 , n36259 , n13246 );
    xnor g34546 ( n29375 , n21448 , n13991 );
    and g34547 ( n18834 , n29845 , n9363 );
    or g34548 ( n8855 , n42370 , n29360 );
    or g34549 ( n26950 , n3396 , n28525 );
    and g34550 ( n19888 , n41876 , n11940 );
    or g34551 ( n9780 , n41113 , n5505 );
    or g34552 ( n36434 , n29322 , n36171 );
    or g34553 ( n28066 , n40819 , n15232 );
    and g34554 ( n3443 , n39605 , n32917 );
    or g34555 ( n40719 , n39408 , n18809 );
    or g34556 ( n1918 , n2834 , n41181 );
    not g34557 ( n1794 , n27776 );
    not g34558 ( n33807 , n4278 );
    and g34559 ( n40182 , n15984 , n21495 );
    and g34560 ( n30430 , n39908 , n22941 );
    not g34561 ( n20186 , n23268 );
    or g34562 ( n36041 , n661 , n24183 );
    and g34563 ( n35101 , n4914 , n34453 );
    xnor g34564 ( n20702 , n36938 , n6082 );
    or g34565 ( n1982 , n7084 , n4150 );
    not g34566 ( n7637 , n25624 );
    and g34567 ( n42299 , n18554 , n34431 );
    and g34568 ( n21612 , n8853 , n12398 );
    or g34569 ( n35996 , n42084 , n21172 );
    and g34570 ( n31045 , n8189 , n615 );
    or g34571 ( n23554 , n27584 , n3234 );
    and g34572 ( n9485 , n8705 , n30688 );
    or g34573 ( n3041 , n25588 , n38008 );
    not g34574 ( n9804 , n35201 );
    or g34575 ( n22168 , n41317 , n34850 );
    and g34576 ( n23776 , n28233 , n40601 );
    or g34577 ( n7515 , n4535 , n1895 );
    and g34578 ( n36244 , n33471 , n23575 );
    and g34579 ( n18564 , n15217 , n18204 );
    xnor g34580 ( n17965 , n32297 , n20033 );
    and g34581 ( n34311 , n33729 , n10783 );
    or g34582 ( n33882 , n36249 , n41130 );
    xnor g34583 ( n21591 , n10558 , n15009 );
    not g34584 ( n11515 , n7911 );
    xnor g34585 ( n30506 , n36444 , n19765 );
    and g34586 ( n27325 , n21419 , n40115 );
    and g34587 ( n16558 , n38906 , n24988 );
    nor g34588 ( n40461 , n15118 , n33260 );
    or g34589 ( n13581 , n41280 , n18613 );
    not g34590 ( n12189 , n29402 );
    xnor g34591 ( n34325 , n36009 , n6413 );
    and g34592 ( n11237 , n21153 , n16122 );
    or g34593 ( n3466 , n28837 , n18082 );
    or g34594 ( n38842 , n34905 , n33660 );
    or g34595 ( n21892 , n41032 , n32786 );
    and g34596 ( n32551 , n4814 , n29717 );
    or g34597 ( n5557 , n36506 , n18236 );
    nor g34598 ( n27135 , n7834 , n1487 );
    xnor g34599 ( n40903 , n9412 , n28495 );
    not g34600 ( n29158 , n20114 );
    nor g34601 ( n26133 , n2445 , n16007 );
    xnor g34602 ( n32159 , n28307 , n35599 );
    not g34603 ( n22120 , n38559 );
    not g34604 ( n24858 , n6227 );
    and g34605 ( n30715 , n1754 , n34888 );
    xnor g34606 ( n27635 , n784 , n2600 );
    nor g34607 ( n40213 , n14039 , n41616 );
    or g34608 ( n27443 , n11974 , n32474 );
    or g34609 ( n26410 , n40710 , n35409 );
    or g34610 ( n17743 , n24665 , n32465 );
    xnor g34611 ( n16406 , n41013 , n23467 );
    nor g34612 ( n39981 , n32874 , n7665 );
    nor g34613 ( n34463 , n33815 , n8451 );
    xnor g34614 ( n23801 , n33148 , n11289 );
    and g34615 ( n36741 , n41735 , n34902 );
    or g34616 ( n27948 , n26588 , n11417 );
    xnor g34617 ( n39859 , n19876 , n19716 );
    or g34618 ( n7428 , n39759 , n35772 );
    not g34619 ( n40419 , n9290 );
    and g34620 ( n13594 , n27755 , n37555 );
    not g34621 ( n15470 , n1702 );
    and g34622 ( n39686 , n29470 , n19854 );
    and g34623 ( n23224 , n20034 , n7553 );
    nor g34624 ( n4474 , n41065 , n16594 );
    and g34625 ( n37544 , n5780 , n14274 );
    not g34626 ( n29668 , n8595 );
    and g34627 ( n20450 , n42802 , n13527 );
    not g34628 ( n39432 , n7673 );
    xnor g34629 ( n18033 , n14370 , n503 );
    and g34630 ( n10718 , n29710 , n31467 );
    xnor g34631 ( n31366 , n17989 , n10552 );
    xnor g34632 ( n908 , n42837 , n41867 );
    and g34633 ( n29054 , n13717 , n20082 );
    and g34634 ( n7336 , n27770 , n35961 );
    or g34635 ( n18676 , n32087 , n36446 );
    and g34636 ( n572 , n18959 , n31257 );
    nor g34637 ( n3678 , n36899 , n11648 );
    and g34638 ( n32681 , n14633 , n24133 );
    xnor g34639 ( n2293 , n25619 , n40449 );
    or g34640 ( n28627 , n32157 , n34436 );
    or g34641 ( n34694 , n4567 , n33133 );
    xnor g34642 ( n16537 , n24064 , n15748 );
    or g34643 ( n18112 , n5203 , n41312 );
    or g34644 ( n3426 , n8494 , n4094 );
    or g34645 ( n5222 , n7383 , n39993 );
    xnor g34646 ( n17158 , n12146 , n38904 );
    and g34647 ( n22647 , n7029 , n39380 );
    or g34648 ( n2192 , n18604 , n37799 );
    or g34649 ( n39011 , n27101 , n29345 );
    and g34650 ( n26788 , n8922 , n14544 );
    or g34651 ( n8693 , n29771 , n28335 );
    and g34652 ( n9543 , n34280 , n29448 );
    and g34653 ( n21446 , n26901 , n12996 );
    not g34654 ( n27331 , n25457 );
    or g34655 ( n23402 , n32890 , n30191 );
    nor g34656 ( n9378 , n13338 , n36758 );
    nor g34657 ( n37524 , n35595 , n29003 );
    or g34658 ( n34370 , n15064 , n36241 );
    and g34659 ( n8143 , n7270 , n39375 );
    or g34660 ( n9949 , n23842 , n31271 );
    xnor g34661 ( n24668 , n11436 , n38038 );
    and g34662 ( n26351 , n5846 , n19357 );
    or g34663 ( n28615 , n31958 , n28230 );
    and g34664 ( n4267 , n10659 , n2305 );
    xnor g34665 ( n17835 , n15111 , n23523 );
    nor g34666 ( n28423 , n11391 , n23741 );
    or g34667 ( n14832 , n16952 , n33700 );
    xnor g34668 ( n19077 , n24265 , n15968 );
    and g34669 ( n5211 , n18318 , n8404 );
    xnor g34670 ( n6508 , n29667 , n33082 );
    or g34671 ( n22200 , n16492 , n6554 );
    not g34672 ( n10361 , n34174 );
    xnor g34673 ( n28875 , n33642 , n33442 );
    and g34674 ( n26828 , n29455 , n39943 );
    xnor g34675 ( n7365 , n32625 , n22937 );
    nor g34676 ( n29776 , n36117 , n29842 );
    or g34677 ( n6932 , n8475 , n15120 );
    xnor g34678 ( n31615 , n32253 , n10638 );
    xnor g34679 ( n42048 , n12146 , n17545 );
    not g34680 ( n7570 , n6825 );
    not g34681 ( n10206 , n14329 );
    not g34682 ( n14826 , n20705 );
    or g34683 ( n3118 , n2183 , n2858 );
    or g34684 ( n25947 , n624 , n27676 );
    xnor g34685 ( n139 , n19700 , n35270 );
    or g34686 ( n38032 , n41159 , n39806 );
    or g34687 ( n36841 , n2864 , n16889 );
    nor g34688 ( n23192 , n21512 , n26091 );
    nor g34689 ( n31710 , n34686 , n21965 );
    or g34690 ( n3724 , n25909 , n2802 );
    or g34691 ( n16196 , n17845 , n25176 );
    or g34692 ( n40688 , n12416 , n28241 );
    nor g34693 ( n37379 , n36993 , n34842 );
    and g34694 ( n2410 , n21588 , n29544 );
    or g34695 ( n19849 , n26743 , n24652 );
    not g34696 ( n33227 , n22291 );
    and g34697 ( n8353 , n25508 , n31457 );
    xnor g34698 ( n12551 , n9441 , n42399 );
    or g34699 ( n35969 , n5795 , n14067 );
    or g34700 ( n34408 , n26177 , n25206 );
    or g34701 ( n22241 , n33020 , n27332 );
    not g34702 ( n17188 , n1670 );
    and g34703 ( n33479 , n41488 , n36725 );
    and g34704 ( n13710 , n33654 , n23852 );
    or g34705 ( n35980 , n4552 , n18642 );
    or g34706 ( n34938 , n7797 , n28643 );
    and g34707 ( n1928 , n39996 , n26812 );
    or g34708 ( n7524 , n30253 , n27234 );
    nor g34709 ( n12452 , n14189 , n28094 );
    xnor g34710 ( n26615 , n6348 , n26239 );
    and g34711 ( n35027 , n9287 , n11406 );
    or g34712 ( n21139 , n871 , n25451 );
    and g34713 ( n37238 , n24392 , n15964 );
    nor g34714 ( n6435 , n35255 , n35779 );
    or g34715 ( n30300 , n25407 , n8254 );
    or g34716 ( n28059 , n33815 , n27947 );
    nor g34717 ( n25652 , n17299 , n30728 );
    or g34718 ( n16123 , n30069 , n12220 );
    and g34719 ( n2910 , n32298 , n27747 );
    or g34720 ( n6823 , n39288 , n10604 );
    not g34721 ( n27874 , n35455 );
    or g34722 ( n28664 , n42486 , n27410 );
    or g34723 ( n9016 , n6504 , n15186 );
    xnor g34724 ( n3017 , n38485 , n30875 );
    nor g34725 ( n22369 , n16821 , n10314 );
    or g34726 ( n28835 , n23808 , n40245 );
    and g34727 ( n34838 , n33586 , n22503 );
    or g34728 ( n40087 , n27884 , n1694 );
    and g34729 ( n20494 , n39606 , n21335 );
    xnor g34730 ( n27370 , n34875 , n1389 );
    nor g34731 ( n30002 , n6131 , n27542 );
    not g34732 ( n5912 , n56 );
    xnor g34733 ( n42164 , n35553 , n15238 );
    or g34734 ( n30773 , n9809 , n1349 );
    nor g34735 ( n15438 , n25895 , n8371 );
    nor g34736 ( n25275 , n29973 , n28594 );
    or g34737 ( n42598 , n29631 , n6000 );
    nor g34738 ( n35257 , n37284 , n28756 );
    and g34739 ( n16509 , n7917 , n4763 );
    nor g34740 ( n34218 , n17471 , n24865 );
    and g34741 ( n33766 , n18616 , n11528 );
    xnor g34742 ( n33005 , n25143 , n24965 );
    or g34743 ( n6230 , n35144 , n27671 );
    not g34744 ( n19788 , n7289 );
    not g34745 ( n8200 , n15733 );
    and g34746 ( n20116 , n14993 , n12321 );
    or g34747 ( n19044 , n23292 , n12726 );
    not g34748 ( n256 , n17342 );
    nor g34749 ( n30957 , n15391 , n29754 );
    or g34750 ( n26221 , n36587 , n30616 );
    or g34751 ( n5953 , n3601 , n20512 );
    not g34752 ( n33745 , n24498 );
    or g34753 ( n33881 , n34411 , n38299 );
    or g34754 ( n5979 , n31355 , n10760 );
    not g34755 ( n17427 , n16987 );
    or g34756 ( n3117 , n20601 , n27380 );
    or g34757 ( n9033 , n6839 , n21942 );
    or g34758 ( n31587 , n33417 , n2107 );
    xnor g34759 ( n25198 , n33652 , n26869 );
    or g34760 ( n7095 , n21473 , n27996 );
    or g34761 ( n9575 , n29844 , n37047 );
    or g34762 ( n1570 , n5170 , n37290 );
    not g34763 ( n4138 , n17397 );
    and g34764 ( n4283 , n1003 , n8431 );
    xnor g34765 ( n18815 , n26513 , n2371 );
    not g34766 ( n19769 , n20111 );
    and g34767 ( n12340 , n32968 , n40996 );
    and g34768 ( n35277 , n11623 , n10352 );
    not g34769 ( n18654 , n31521 );
    xnor g34770 ( n35406 , n26972 , n32274 );
    nor g34771 ( n32987 , n24917 , n6019 );
    not g34772 ( n12059 , n4961 );
    and g34773 ( n15268 , n23284 , n1760 );
    or g34774 ( n25564 , n35690 , n7914 );
    or g34775 ( n26375 , n32611 , n33616 );
    or g34776 ( n19556 , n17702 , n36203 );
    or g34777 ( n32135 , n4532 , n2565 );
    nor g34778 ( n7003 , n15717 , n23468 );
    and g34779 ( n6832 , n408 , n22162 );
    or g34780 ( n13632 , n27503 , n16336 );
    or g34781 ( n19507 , n20446 , n23127 );
    not g34782 ( n34874 , n31164 );
    and g34783 ( n27122 , n12809 , n21632 );
    not g34784 ( n2127 , n38080 );
    and g34785 ( n5455 , n28391 , n23036 );
    or g34786 ( n33672 , n31734 , n37387 );
    nor g34787 ( n6637 , n7339 , n25298 );
    not g34788 ( n7467 , n39461 );
    or g34789 ( n42030 , n7646 , n22743 );
    not g34790 ( n18880 , n20416 );
    nor g34791 ( n39416 , n31429 , n35877 );
    or g34792 ( n237 , n31350 , n15064 );
    or g34793 ( n28652 , n19159 , n17646 );
    and g34794 ( n3971 , n9342 , n8548 );
    and g34795 ( n32826 , n15754 , n33851 );
    or g34796 ( n29523 , n4361 , n15434 );
    xnor g34797 ( n40159 , n39217 , n28164 );
    or g34798 ( n37976 , n11417 , n11648 );
    or g34799 ( n21523 , n28433 , n22282 );
    or g34800 ( n36683 , n16598 , n28139 );
    and g34801 ( n39002 , n37026 , n82 );
    not g34802 ( n27311 , n26673 );
    or g34803 ( n42659 , n3583 , n17010 );
    or g34804 ( n6150 , n22373 , n29579 );
    or g34805 ( n24961 , n25238 , n14420 );
    xnor g34806 ( n19891 , n9448 , n32715 );
    not g34807 ( n23330 , n13720 );
    or g34808 ( n1548 , n12432 , n34222 );
    and g34809 ( n24652 , n26371 , n27706 );
    and g34810 ( n42165 , n1722 , n849 );
    not g34811 ( n13041 , n38752 );
    or g34812 ( n25617 , n10581 , n41413 );
    or g34813 ( n16428 , n35182 , n18697 );
    nor g34814 ( n17032 , n23619 , n32975 );
    nor g34815 ( n13556 , n6671 , n33410 );
    or g34816 ( n28290 , n12198 , n30924 );
    or g34817 ( n14577 , n33094 , n1006 );
    not g34818 ( n14675 , n23678 );
    nor g34819 ( n16679 , n38041 , n30398 );
    not g34820 ( n34931 , n23541 );
    or g34821 ( n3221 , n13187 , n38031 );
    or g34822 ( n31435 , n19221 , n24286 );
    not g34823 ( n25137 , n26445 );
    and g34824 ( n23146 , n10828 , n20964 );
    or g34825 ( n31413 , n40785 , n9582 );
    or g34826 ( n38928 , n6503 , n3483 );
    or g34827 ( n5898 , n35438 , n31926 );
    nor g34828 ( n26797 , n29053 , n3556 );
    and g34829 ( n31140 , n10116 , n4135 );
    not g34830 ( n17654 , n22934 );
    or g34831 ( n12759 , n32638 , n25626 );
    or g34832 ( n9741 , n36316 , n987 );
    or g34833 ( n30705 , n24907 , n42563 );
    not g34834 ( n27801 , n29091 );
    xnor g34835 ( n22840 , n3179 , n39714 );
    and g34836 ( n23012 , n14990 , n18164 );
    not g34837 ( n28003 , n42844 );
    and g34838 ( n7453 , n23900 , n36414 );
    or g34839 ( n6172 , n34008 , n3355 );
    xnor g34840 ( n8923 , n26210 , n20369 );
    or g34841 ( n21792 , n14707 , n17165 );
    or g34842 ( n36961 , n14986 , n36251 );
    and g34843 ( n17573 , n2468 , n35517 );
    and g34844 ( n912 , n41299 , n6219 );
    xnor g34845 ( n15190 , n34848 , n13073 );
    and g34846 ( n28696 , n38202 , n19680 );
    and g34847 ( n14075 , n28979 , n3859 );
    nor g34848 ( n40439 , n9848 , n16430 );
    or g34849 ( n15068 , n12236 , n36943 );
    not g34850 ( n36806 , n27555 );
    and g34851 ( n23931 , n9861 , n33056 );
    not g34852 ( n2501 , n27148 );
    or g34853 ( n21658 , n16133 , n3049 );
    or g34854 ( n40163 , n13998 , n32395 );
    and g34855 ( n7019 , n24631 , n5835 );
    and g34856 ( n17542 , n945 , n42401 );
    not g34857 ( n13352 , n41608 );
    and g34858 ( n19404 , n42900 , n8668 );
    and g34859 ( n20740 , n15442 , n8425 );
    not g34860 ( n1580 , n15583 );
    or g34861 ( n39545 , n24180 , n22123 );
    or g34862 ( n31148 , n29214 , n37232 );
    and g34863 ( n30182 , n19071 , n32257 );
    or g34864 ( n31528 , n36355 , n8209 );
    nor g34865 ( n12182 , n31865 , n4444 );
    or g34866 ( n20480 , n15030 , n41789 );
    and g34867 ( n20106 , n10981 , n39567 );
    not g34868 ( n2612 , n8854 );
    xnor g34869 ( n18149 , n24750 , n28629 );
    xnor g34870 ( n34886 , n25849 , n31095 );
    and g34871 ( n26746 , n2974 , n29928 );
    and g34872 ( n38963 , n4754 , n13462 );
    and g34873 ( n39391 , n25365 , n22779 );
    or g34874 ( n42102 , n32919 , n37787 );
    not g34875 ( n14348 , n1843 );
    and g34876 ( n31026 , n24388 , n13788 );
    or g34877 ( n571 , n24656 , n4624 );
    xnor g34878 ( n37824 , n7190 , n28085 );
    nor g34879 ( n27489 , n23554 , n27285 );
    xnor g34880 ( n5370 , n40176 , n22448 );
    or g34881 ( n11684 , n32640 , n21802 );
    or g34882 ( n23691 , n33152 , n20085 );
    and g34883 ( n12868 , n19620 , n11235 );
    xnor g34884 ( n2411 , n29034 , n189 );
    and g34885 ( n2020 , n38561 , n12753 );
    or g34886 ( n33341 , n28246 , n9298 );
    nor g34887 ( n1726 , n32277 , n38237 );
    or g34888 ( n42695 , n15138 , n28274 );
    or g34889 ( n31477 , n10625 , n32040 );
    and g34890 ( n20020 , n7685 , n32061 );
    xnor g34891 ( n27833 , n20952 , n34179 );
    nor g34892 ( n15418 , n18131 , n42908 );
    or g34893 ( n29561 , n643 , n24695 );
    and g34894 ( n30440 , n38301 , n16442 );
    xnor g34895 ( n18831 , n13597 , n23183 );
    not g34896 ( n11976 , n29892 );
    and g34897 ( n10404 , n2698 , n22370 );
    nor g34898 ( n2748 , n41040 , n26688 );
    and g34899 ( n8916 , n16874 , n6979 );
    xnor g34900 ( n10885 , n19172 , n15679 );
    and g34901 ( n32072 , n15667 , n39546 );
    nor g34902 ( n2449 , n12146 , n21354 );
    nor g34903 ( n12186 , n11702 , n29127 );
    or g34904 ( n33007 , n36117 , n39093 );
    not g34905 ( n41944 , n34057 );
    not g34906 ( n27346 , n26816 );
    xnor g34907 ( n11145 , n2413 , n33981 );
    or g34908 ( n32669 , n40184 , n16825 );
    or g34909 ( n9496 , n833 , n9426 );
    nor g34910 ( n15726 , n26058 , n30496 );
    or g34911 ( n40756 , n328 , n10602 );
    and g34912 ( n19989 , n18653 , n7432 );
    or g34913 ( n10786 , n6834 , n12625 );
    and g34914 ( n11044 , n26121 , n29843 );
    or g34915 ( n33396 , n24588 , n30212 );
    not g34916 ( n4545 , n32376 );
    or g34917 ( n2349 , n40175 , n37263 );
    nor g34918 ( n36377 , n18866 , n6595 );
    or g34919 ( n3965 , n16514 , n1044 );
    not g34920 ( n4326 , n16537 );
    or g34921 ( n7487 , n29076 , n2972 );
    or g34922 ( n13656 , n42792 , n31442 );
    and g34923 ( n37780 , n6498 , n21321 );
    or g34924 ( n9899 , n21427 , n1605 );
    not g34925 ( n41433 , n38431 );
    not g34926 ( n31138 , n20714 );
    or g34927 ( n1914 , n41546 , n20719 );
    or g34928 ( n18804 , n6503 , n39205 );
    or g34929 ( n30359 , n22333 , n35981 );
    or g34930 ( n32889 , n9995 , n42479 );
    xnor g34931 ( n25245 , n6870 , n11697 );
    xnor g34932 ( n18488 , n1464 , n34703 );
    or g34933 ( n5858 , n34039 , n407 );
    xnor g34934 ( n13020 , n11436 , n3477 );
    nor g34935 ( n37995 , n14471 , n25969 );
    and g34936 ( n31525 , n23267 , n33786 );
    or g34937 ( n12583 , n36585 , n13115 );
    not g34938 ( n5478 , n9774 );
    not g34939 ( n30929 , n18519 );
    and g34940 ( n4816 , n8247 , n13575 );
    and g34941 ( n28499 , n5548 , n78 );
    nor g34942 ( n20830 , n28872 , n42755 );
    xnor g34943 ( n29445 , n30454 , n11680 );
    and g34944 ( n27351 , n9334 , n29801 );
    and g34945 ( n21334 , n11627 , n35583 );
    nor g34946 ( n14088 , n17744 , n32877 );
    or g34947 ( n11699 , n33683 , n28139 );
    nor g34948 ( n26027 , n9084 , n42185 );
    and g34949 ( n40195 , n29527 , n23064 );
    nor g34950 ( n9515 , n38580 , n1341 );
    or g34951 ( n38313 , n38058 , n23902 );
    or g34952 ( n11891 , n7146 , n11026 );
    not g34953 ( n6959 , n1519 );
    not g34954 ( n34875 , n40372 );
    or g34955 ( n1145 , n28745 , n31014 );
    or g34956 ( n21215 , n41597 , n14481 );
    or g34957 ( n24886 , n41025 , n15857 );
    not g34958 ( n34173 , n22212 );
    not g34959 ( n49 , n31058 );
    and g34960 ( n22669 , n38322 , n4354 );
    nor g34961 ( n11722 , n17120 , n9452 );
    or g34962 ( n34583 , n5896 , n19496 );
    or g34963 ( n35977 , n6628 , n29266 );
    and g34964 ( n33504 , n20559 , n29152 );
    or g34965 ( n26378 , n9229 , n21259 );
    and g34966 ( n29650 , n34693 , n41875 );
    or g34967 ( n381 , n42675 , n6122 );
    and g34968 ( n33630 , n9907 , n28793 );
    not g34969 ( n38922 , n23004 );
    or g34970 ( n36516 , n12138 , n18828 );
    and g34971 ( n20938 , n24742 , n7926 );
    and g34972 ( n39689 , n3008 , n27495 );
    or g34973 ( n26541 , n19469 , n25190 );
    or g34974 ( n32535 , n24820 , n38022 );
    not g34975 ( n8097 , n19745 );
    nor g34976 ( n30418 , n15010 , n17341 );
    and g34977 ( n26801 , n21052 , n10380 );
    or g34978 ( n42696 , n12804 , n33039 );
    xnor g34979 ( n10937 , n21654 , n23774 );
    and g34980 ( n20666 , n36512 , n36475 );
    nor g34981 ( n42138 , n22089 , n7417 );
    or g34982 ( n20063 , n37061 , n15714 );
    and g34983 ( n4619 , n30563 , n9340 );
    nor g34984 ( n36343 , n2645 , n12395 );
    and g34985 ( n259 , n12324 , n36065 );
    xnor g34986 ( n20376 , n26579 , n16768 );
    nor g34987 ( n18321 , n589 , n10778 );
    nor g34988 ( n17284 , n13216 , n30571 );
    and g34989 ( n6794 , n12281 , n34979 );
    or g34990 ( n9806 , n28947 , n432 );
    or g34991 ( n11656 , n16436 , n36962 );
    and g34992 ( n35466 , n5622 , n8850 );
    or g34993 ( n125 , n22460 , n15531 );
    or g34994 ( n40842 , n8973 , n8568 );
    xnor g34995 ( n757 , n14338 , n12315 );
    or g34996 ( n4935 , n21048 , n20855 );
    nor g34997 ( n41371 , n33697 , n13791 );
    and g34998 ( n39817 , n497 , n9274 );
    nor g34999 ( n12927 , n24200 , n14114 );
    nor g35000 ( n26664 , n34292 , n25702 );
    not g35001 ( n7613 , n13140 );
    and g35002 ( n8664 , n6522 , n3262 );
    or g35003 ( n9404 , n6358 , n18908 );
    or g35004 ( n22248 , n28298 , n27292 );
    not g35005 ( n29859 , n41992 );
    not g35006 ( n4847 , n19616 );
    not g35007 ( n13373 , n11713 );
    nor g35008 ( n37467 , n38957 , n38876 );
    not g35009 ( n13515 , n33481 );
    or g35010 ( n15916 , n37098 , n22845 );
    or g35011 ( n1560 , n17279 , n37633 );
    or g35012 ( n11287 , n1581 , n22153 );
    or g35013 ( n35484 , n107 , n22755 );
    or g35014 ( n7432 , n351 , n9042 );
    not g35015 ( n39810 , n38262 );
    xnor g35016 ( n7535 , n29740 , n7453 );
    or g35017 ( n21228 , n394 , n2121 );
    or g35018 ( n16431 , n19486 , n25123 );
    or g35019 ( n34599 , n24454 , n21781 );
    or g35020 ( n5501 , n31227 , n19394 );
    not g35021 ( n26959 , n5819 );
    or g35022 ( n28552 , n17244 , n22335 );
    nor g35023 ( n39078 , n13785 , n34965 );
    or g35024 ( n3377 , n16817 , n38249 );
    and g35025 ( n11952 , n24970 , n40025 );
    and g35026 ( n375 , n29573 , n34923 );
    xnor g35027 ( n5247 , n6625 , n24609 );
    and g35028 ( n30010 , n18630 , n4362 );
    and g35029 ( n10136 , n15100 , n15311 );
    and g35030 ( n42174 , n29195 , n7193 );
    or g35031 ( n13914 , n41360 , n32994 );
    and g35032 ( n14393 , n28579 , n3332 );
    nor g35033 ( n723 , n4388 , n33597 );
    or g35034 ( n33734 , n9544 , n28400 );
    and g35035 ( n2239 , n41795 , n811 );
    or g35036 ( n24155 , n38428 , n28143 );
    nor g35037 ( n39354 , n2199 , n35801 );
    and g35038 ( n7031 , n19038 , n30905 );
    and g35039 ( n6570 , n23870 , n1508 );
    not g35040 ( n32144 , n38920 );
    or g35041 ( n32203 , n42361 , n18420 );
    and g35042 ( n33527 , n40782 , n28049 );
    nor g35043 ( n23533 , n38806 , n36431 );
    nor g35044 ( n2697 , n23930 , n41944 );
    or g35045 ( n8791 , n13470 , n34676 );
    nor g35046 ( n10263 , n2651 , n3617 );
    or g35047 ( n39225 , n39266 , n7961 );
    or g35048 ( n27937 , n7864 , n18428 );
    xnor g35049 ( n26247 , n8255 , n18984 );
    and g35050 ( n3116 , n1034 , n6561 );
    or g35051 ( n3584 , n19030 , n23493 );
    or g35052 ( n34186 , n20015 , n29076 );
    and g35053 ( n3446 , n8286 , n7103 );
    xnor g35054 ( n15742 , n4334 , n42052 );
    or g35055 ( n26599 , n12191 , n17249 );
    xnor g35056 ( n25066 , n14530 , n2272 );
    xnor g35057 ( n39713 , n5891 , n9813 );
    xnor g35058 ( n25827 , n4510 , n34565 );
    xnor g35059 ( n32553 , n34768 , n35794 );
    and g35060 ( n40605 , n13736 , n19988 );
    or g35061 ( n35542 , n7934 , n11061 );
    and g35062 ( n36733 , n41120 , n32531 );
    or g35063 ( n24570 , n8005 , n40696 );
    or g35064 ( n32354 , n3385 , n611 );
    or g35065 ( n27289 , n15689 , n4020 );
    and g35066 ( n25806 , n27159 , n42242 );
    or g35067 ( n37575 , n27865 , n8658 );
    and g35068 ( n26820 , n5667 , n38966 );
    or g35069 ( n36336 , n38563 , n11435 );
    and g35070 ( n10730 , n31766 , n7147 );
    or g35071 ( n20909 , n23445 , n9012 );
    or g35072 ( n24861 , n32053 , n39113 );
    nor g35073 ( n36227 , n14334 , n26709 );
    or g35074 ( n38843 , n40287 , n11708 );
    or g35075 ( n1962 , n21142 , n27532 );
    or g35076 ( n16522 , n14610 , n27527 );
    not g35077 ( n41014 , n21234 );
    not g35078 ( n12742 , n31043 );
    and g35079 ( n10269 , n5979 , n14950 );
    nor g35080 ( n42100 , n6077 , n21811 );
    not g35081 ( n22625 , n33632 );
    not g35082 ( n34305 , n13595 );
    or g35083 ( n33393 , n22821 , n22145 );
    or g35084 ( n8799 , n24323 , n20636 );
    or g35085 ( n15119 , n2703 , n37027 );
    nor g35086 ( n25873 , n25826 , n27062 );
    or g35087 ( n31589 , n33981 , n29023 );
    xnor g35088 ( n31837 , n16473 , n17362 );
    nor g35089 ( n41868 , n16505 , n28086 );
    nor g35090 ( n15976 , n10110 , n22233 );
    or g35091 ( n1916 , n10926 , n4901 );
    nor g35092 ( n20682 , n17744 , n4441 );
    or g35093 ( n29716 , n29056 , n8344 );
    or g35094 ( n17523 , n29256 , n36701 );
    and g35095 ( n8372 , n3968 , n13691 );
    and g35096 ( n7435 , n28804 , n37205 );
    or g35097 ( n12900 , n2260 , n23171 );
    xnor g35098 ( n30982 , n8638 , n5653 );
    and g35099 ( n10643 , n34953 , n28118 );
    not g35100 ( n1730 , n4131 );
    or g35101 ( n19921 , n28383 , n15000 );
    xnor g35102 ( n181 , n2139 , n2509 );
    xnor g35103 ( n12250 , n6625 , n10081 );
    or g35104 ( n2606 , n37806 , n25442 );
    and g35105 ( n36251 , n2851 , n24239 );
    and g35106 ( n26439 , n31363 , n5224 );
    and g35107 ( n27515 , n5788 , n41204 );
    not g35108 ( n26803 , n6869 );
    and g35109 ( n42610 , n17597 , n26671 );
    or g35110 ( n3665 , n29346 , n34567 );
    xnor g35111 ( n2547 , n31456 , n41638 );
    or g35112 ( n3984 , n9760 , n12129 );
    or g35113 ( n16906 , n9375 , n31567 );
    and g35114 ( n7094 , n38072 , n3352 );
    or g35115 ( n1556 , n42516 , n23940 );
    or g35116 ( n21107 , n4599 , n36880 );
    nor g35117 ( n39347 , n5398 , n29717 );
    and g35118 ( n42451 , n25321 , n23384 );
    nor g35119 ( n42439 , n16544 , n20252 );
    xnor g35120 ( n21532 , n17603 , n12774 );
    not g35121 ( n21772 , n1853 );
    or g35122 ( n16125 , n39213 , n19517 );
    and g35123 ( n17848 , n24182 , n17716 );
    xnor g35124 ( n13669 , n28925 , n35698 );
    or g35125 ( n41727 , n23933 , n41981 );
    nor g35126 ( n18981 , n25172 , n24765 );
    or g35127 ( n20094 , n943 , n22892 );
    nor g35128 ( n35454 , n10903 , n7979 );
    or g35129 ( n8431 , n39215 , n41108 );
    and g35130 ( n34080 , n38968 , n13803 );
    or g35131 ( n4950 , n20518 , n36891 );
    or g35132 ( n7983 , n12666 , n21221 );
    or g35133 ( n16769 , n8210 , n41676 );
    not g35134 ( n11340 , n29117 );
    and g35135 ( n6554 , n1531 , n40682 );
    not g35136 ( n10284 , n13300 );
    or g35137 ( n36752 , n20862 , n33216 );
    not g35138 ( n5973 , n13722 );
    and g35139 ( n17877 , n18137 , n19011 );
    xnor g35140 ( n29610 , n42779 , n1507 );
    and g35141 ( n13000 , n20640 , n332 );
    xnor g35142 ( n29247 , n8881 , n14707 );
    not g35143 ( n21881 , n3084 );
    and g35144 ( n16838 , n42686 , n14752 );
    and g35145 ( n4713 , n12521 , n23364 );
    and g35146 ( n25653 , n25041 , n38778 );
    nor g35147 ( n38710 , n19602 , n9840 );
    or g35148 ( n30230 , n2675 , n986 );
    not g35149 ( n7235 , n39148 );
    not g35150 ( n2804 , n12137 );
    not g35151 ( n21813 , n41946 );
    and g35152 ( n9601 , n21757 , n23699 );
    not g35153 ( n5144 , n17744 );
    nor g35154 ( n41920 , n33026 , n34539 );
    not g35155 ( n19311 , n10536 );
    not g35156 ( n3993 , n41713 );
    not g35157 ( n35193 , n5259 );
    or g35158 ( n8776 , n14707 , n18567 );
    xnor g35159 ( n4408 , n24791 , n18570 );
    not g35160 ( n28673 , n30738 );
    and g35161 ( n26953 , n40545 , n20226 );
    or g35162 ( n34857 , n4745 , n10657 );
    or g35163 ( n666 , n41705 , n3927 );
    or g35164 ( n21717 , n24745 , n29021 );
    nor g35165 ( n35166 , n6198 , n8012 );
    or g35166 ( n12201 , n4936 , n6316 );
    not g35167 ( n29885 , n40435 );
    nor g35168 ( n24246 , n34292 , n1177 );
    nor g35169 ( n42065 , n1507 , n37065 );
    or g35170 ( n31105 , n40209 , n8459 );
    nor g35171 ( n16515 , n357 , n39782 );
    and g35172 ( n35249 , n29665 , n36357 );
    or g35173 ( n11532 , n36285 , n24696 );
    not g35174 ( n27016 , n42742 );
    nor g35175 ( n6399 , n17120 , n40930 );
    not g35176 ( n22219 , n41477 );
    and g35177 ( n6252 , n3644 , n18579 );
    not g35178 ( n27220 , n8604 );
    or g35179 ( n40893 , n19853 , n40807 );
    or g35180 ( n28509 , n11600 , n30834 );
    xnor g35181 ( n26126 , n24943 , n17959 );
    or g35182 ( n39800 , n36508 , n27566 );
    or g35183 ( n41719 , n32605 , n36177 );
    and g35184 ( n12315 , n35383 , n12422 );
    and g35185 ( n12653 , n4481 , n9320 );
    not g35186 ( n30448 , n8277 );
    xnor g35187 ( n29428 , n37403 , n22528 );
    or g35188 ( n15168 , n9695 , n37718 );
    or g35189 ( n22302 , n9655 , n27607 );
    or g35190 ( n9712 , n35523 , n34821 );
    or g35191 ( n28435 , n17161 , n22611 );
    or g35192 ( n20095 , n31123 , n34316 );
    nor g35193 ( n2863 , n25777 , n6716 );
    not g35194 ( n15658 , n27569 );
    or g35195 ( n34869 , n7410 , n33322 );
    xnor g35196 ( n36106 , n11436 , n33539 );
    and g35197 ( n31142 , n33305 , n15557 );
    or g35198 ( n16864 , n34253 , n6923 );
    and g35199 ( n14449 , n19572 , n13068 );
    or g35200 ( n41866 , n19273 , n27781 );
    and g35201 ( n7775 , n27911 , n21629 );
    or g35202 ( n25799 , n35834 , n39184 );
    or g35203 ( n40562 , n5896 , n21157 );
    nor g35204 ( n39326 , n2235 , n9667 );
    or g35205 ( n14264 , n18834 , n24138 );
    not g35206 ( n29511 , n13919 );
    or g35207 ( n11303 , n24745 , n36492 );
    and g35208 ( n31955 , n33171 , n31768 );
    not g35209 ( n14454 , n37540 );
    and g35210 ( n34475 , n5535 , n20552 );
    nor g35211 ( n7176 , n9436 , n38765 );
    or g35212 ( n13126 , n24251 , n12210 );
    or g35213 ( n18171 , n20288 , n12558 );
    xnor g35214 ( n23309 , n8971 , n19129 );
    not g35215 ( n6742 , n24510 );
    or g35216 ( n20533 , n8494 , n15287 );
    and g35217 ( n20939 , n42009 , n17186 );
    not g35218 ( n42133 , n39381 );
    or g35219 ( n13436 , n41534 , n7356 );
    not g35220 ( n15020 , n16257 );
    nor g35221 ( n32768 , n14364 , n29051 );
    or g35222 ( n5755 , n20726 , n28166 );
    not g35223 ( n4870 , n33125 );
    and g35224 ( n30367 , n39545 , n23279 );
    or g35225 ( n24634 , n5633 , n40724 );
    not g35226 ( n1759 , n41963 );
    xnor g35227 ( n9945 , n21301 , n31443 );
    and g35228 ( n2785 , n19581 , n39840 );
    and g35229 ( n5952 , n36551 , n36986 );
    or g35230 ( n35545 , n31016 , n24854 );
    not g35231 ( n37590 , n16898 );
    or g35232 ( n28467 , n33695 , n42152 );
    or g35233 ( n35791 , n2731 , n6478 );
    or g35234 ( n7402 , n2683 , n38340 );
    or g35235 ( n20656 , n15700 , n28341 );
    or g35236 ( n265 , n35772 , n40351 );
    not g35237 ( n1903 , n7561 );
    xnor g35238 ( n16255 , n36759 , n20125 );
    xnor g35239 ( n23636 , n17206 , n11945 );
    or g35240 ( n42658 , n39118 , n24049 );
    or g35241 ( n2041 , n41641 , n19389 );
    nor g35242 ( n22181 , n16598 , n4222 );
    and g35243 ( n19662 , n14527 , n29590 );
    nor g35244 ( n38311 , n23561 , n7251 );
    not g35245 ( n20684 , n14925 );
    or g35246 ( n1727 , n10166 , n33414 );
    or g35247 ( n32584 , n39843 , n313 );
    nor g35248 ( n4534 , n24331 , n26921 );
    not g35249 ( n19861 , n19435 );
    and g35250 ( n20273 , n9281 , n35020 );
    not g35251 ( n7082 , n26329 );
    or g35252 ( n30890 , n37960 , n39428 );
    or g35253 ( n361 , n28395 , n21249 );
    xnor g35254 ( n32424 , n9990 , n4037 );
    not g35255 ( n18997 , n6790 );
    xnor g35256 ( n21066 , n42509 , n15070 );
    not g35257 ( n39536 , n29777 );
    xnor g35258 ( n15843 , n6969 , n28128 );
    or g35259 ( n20101 , n4492 , n40226 );
    or g35260 ( n26802 , n41401 , n31724 );
    or g35261 ( n31365 , n18793 , n21721 );
    and g35262 ( n37903 , n20685 , n37541 );
    or g35263 ( n28410 , n8611 , n12677 );
    or g35264 ( n12147 , n12734 , n36941 );
    xnor g35265 ( n17056 , n7943 , n38876 );
    or g35266 ( n5751 , n11855 , n1696 );
    not g35267 ( n13668 , n5646 );
    not g35268 ( n12734 , n28150 );
    or g35269 ( n6590 , n39883 , n5424 );
    and g35270 ( n33312 , n8145 , n7306 );
    and g35271 ( n40194 , n21256 , n15783 );
    nor g35272 ( n39735 , n39266 , n5790 );
    and g35273 ( n28114 , n33551 , n8100 );
    or g35274 ( n23879 , n21904 , n35829 );
    or g35275 ( n42198 , n39974 , n17827 );
    xnor g35276 ( n37530 , n24218 , n40422 );
    and g35277 ( n19608 , n28443 , n31701 );
    not g35278 ( n25150 , n6617 );
    or g35279 ( n37352 , n18623 , n12846 );
    or g35280 ( n24284 , n13193 , n21703 );
    and g35281 ( n23233 , n18463 , n13070 );
    or g35282 ( n16932 , n22020 , n29382 );
    or g35283 ( n42193 , n14726 , n3728 );
    xnor g35284 ( n15043 , n36009 , n29430 );
    or g35285 ( n18074 , n33865 , n12947 );
    not g35286 ( n15051 , n31089 );
    or g35287 ( n29931 , n825 , n35002 );
    or g35288 ( n4915 , n6628 , n26374 );
    and g35289 ( n15888 , n2103 , n4400 );
    not g35290 ( n42016 , n30014 );
    nor g35291 ( n15053 , n39655 , n30107 );
    or g35292 ( n13048 , n20888 , n5183 );
    not g35293 ( n29303 , n40301 );
    nor g35294 ( n35994 , n14840 , n28765 );
    or g35295 ( n19554 , n24547 , n29156 );
    xnor g35296 ( n25340 , n24165 , n20942 );
    and g35297 ( n17222 , n39644 , n41524 );
    nor g35298 ( n33403 , n23708 , n9214 );
    and g35299 ( n25317 , n311 , n26912 );
    and g35300 ( n15877 , n7519 , n26892 );
    xnor g35301 ( n32706 , n4877 , n14699 );
    and g35302 ( n37339 , n17201 , n5383 );
    not g35303 ( n37300 , n31765 );
    not g35304 ( n4798 , n5696 );
    nor g35305 ( n147 , n22921 , n6614 );
    or g35306 ( n1645 , n24670 , n18622 );
    xnor g35307 ( n32248 , n34731 , n1520 );
    nor g35308 ( n36892 , n2038 , n18876 );
    nor g35309 ( n10562 , n34240 , n41491 );
    xnor g35310 ( n42650 , n19068 , n17120 );
    and g35311 ( n7 , n12272 , n10678 );
    nor g35312 ( n34650 , n6138 , n12733 );
    or g35313 ( n12019 , n36235 , n19210 );
    and g35314 ( n9232 , n20992 , n27837 );
    and g35315 ( n28777 , n7252 , n5345 );
    or g35316 ( n14706 , n31958 , n50 );
    xnor g35317 ( n25912 , n40 , n27582 );
    and g35318 ( n19288 , n28636 , n34663 );
    xnor g35319 ( n34078 , n18530 , n23423 );
    or g35320 ( n40537 , n34559 , n39660 );
    or g35321 ( n10479 , n6118 , n4625 );
    and g35322 ( n31077 , n9552 , n38575 );
    and g35323 ( n37371 , n12646 , n31406 );
    or g35324 ( n24944 , n19969 , n34072 );
    or g35325 ( n11148 , n18728 , n25064 );
    and g35326 ( n38562 , n16583 , n36912 );
    not g35327 ( n33417 , n18896 );
    or g35328 ( n4410 , n22428 , n38230 );
    nor g35329 ( n8275 , n39025 , n9524 );
    or g35330 ( n34064 , n30251 , n14955 );
    or g35331 ( n33857 , n17142 , n21187 );
    xnor g35332 ( n13501 , n12300 , n10257 );
    and g35333 ( n21722 , n40519 , n31977 );
    not g35334 ( n15591 , n36939 );
    and g35335 ( n41259 , n7444 , n14078 );
    not g35336 ( n34478 , n35392 );
    not g35337 ( n38041 , n13275 );
    not g35338 ( n35965 , n23004 );
    or g35339 ( n40451 , n33859 , n304 );
    or g35340 ( n42692 , n38559 , n19240 );
    and g35341 ( n5812 , n25208 , n26150 );
    xnor g35342 ( n2469 , n11060 , n27138 );
    xnor g35343 ( n3389 , n42475 , n39726 );
    not g35344 ( n9078 , n39452 );
    or g35345 ( n41935 , n9544 , n11495 );
    nor g35346 ( n30233 , n6885 , n31006 );
    or g35347 ( n30050 , n26067 , n23462 );
    or g35348 ( n27856 , n40579 , n25573 );
    or g35349 ( n21458 , n22489 , n11565 );
    nor g35350 ( n16926 , n12954 , n10680 );
    xnor g35351 ( n12864 , n784 , n9212 );
    or g35352 ( n6709 , n35941 , n256 );
    or g35353 ( n523 , n2710 , n42384 );
    and g35354 ( n6135 , n39074 , n34947 );
    and g35355 ( n37957 , n33942 , n27356 );
    not g35356 ( n18874 , n6660 );
    and g35357 ( n7683 , n37542 , n28580 );
    nor g35358 ( n34234 , n19221 , n2335 );
    xnor g35359 ( n7393 , n35813 , n30658 );
    and g35360 ( n30218 , n42750 , n31572 );
    or g35361 ( n19378 , n13236 , n8971 );
    nor g35362 ( n12400 , n21184 , n4675 );
    or g35363 ( n38302 , n1457 , n37439 );
    or g35364 ( n13349 , n22440 , n2525 );
    or g35365 ( n23329 , n32446 , n23310 );
    nor g35366 ( n7590 , n35605 , n42744 );
    and g35367 ( n21214 , n6961 , n32086 );
    xnor g35368 ( n12071 , n27972 , n20577 );
    and g35369 ( n1975 , n41748 , n17693 );
    or g35370 ( n11266 , n8941 , n24415 );
    or g35371 ( n20088 , n24156 , n28924 );
    or g35372 ( n7780 , n16609 , n5984 );
    nor g35373 ( n31676 , n25438 , n26477 );
    not g35374 ( n3656 , n17567 );
    xnor g35375 ( n41709 , n35553 , n21113 );
    not g35376 ( n39456 , n9691 );
    or g35377 ( n1218 , n12923 , n17229 );
    nor g35378 ( n23181 , n22782 , n36352 );
    or g35379 ( n2485 , n11321 , n1820 );
    and g35380 ( n28153 , n2669 , n42628 );
    or g35381 ( n23408 , n8997 , n10967 );
    and g35382 ( n14184 , n2594 , n1094 );
    nor g35383 ( n11053 , n14707 , n10488 );
    and g35384 ( n5059 , n10658 , n29863 );
    and g35385 ( n30423 , n22573 , n39034 );
    not g35386 ( n3366 , n8627 );
    xnor g35387 ( n10667 , n7922 , n10187 );
    or g35388 ( n23103 , n38157 , n41534 );
    or g35389 ( n23172 , n26270 , n15934 );
    or g35390 ( n10615 , n4043 , n30073 );
    not g35391 ( n32108 , n6997 );
    and g35392 ( n9206 , n39971 , n19072 );
    not g35393 ( n33438 , n24747 );
    or g35394 ( n39853 , n4535 , n18399 );
    xnor g35395 ( n40233 , n8873 , n27661 );
    and g35396 ( n34608 , n41844 , n22689 );
    nor g35397 ( n29903 , n18520 , n15624 );
    nor g35398 ( n5295 , n7358 , n6322 );
    and g35399 ( n3845 , n8773 , n501 );
    not g35400 ( n38084 , n31965 );
    or g35401 ( n35357 , n5031 , n18933 );
    and g35402 ( n37065 , n26702 , n39313 );
    xnor g35403 ( n17268 , n1573 , n36123 );
    or g35404 ( n27322 , n37642 , n30263 );
    not g35405 ( n36319 , n41784 );
    nor g35406 ( n2054 , n31542 , n13310 );
    not g35407 ( n14953 , n37306 );
    nor g35408 ( n1763 , n29702 , n38044 );
    nor g35409 ( n18250 , n27173 , n10261 );
    nor g35410 ( n37853 , n16788 , n40903 );
    xnor g35411 ( n23608 , n21941 , n3521 );
    not g35412 ( n9951 , n21503 );
    or g35413 ( n8176 , n31946 , n7707 );
    or g35414 ( n38757 , n22091 , n1129 );
    or g35415 ( n16099 , n15379 , n6236 );
    xnor g35416 ( n9674 , n22773 , n24143 );
    xnor g35417 ( n21736 , n21192 , n36501 );
    nor g35418 ( n31994 , n14840 , n6346 );
    and g35419 ( n25768 , n6855 , n29557 );
    nor g35420 ( n17979 , n33981 , n40175 );
    nor g35421 ( n7679 , n29303 , n40495 );
    and g35422 ( n41560 , n16493 , n30154 );
    not g35423 ( n31460 , n40173 );
    or g35424 ( n11457 , n22553 , n2215 );
    or g35425 ( n9169 , n31026 , n12674 );
    not g35426 ( n29452 , n34202 );
    xnor g35427 ( n28376 , n31099 , n24723 );
    or g35428 ( n10828 , n38896 , n29316 );
    or g35429 ( n37979 , n40253 , n19682 );
    nor g35430 ( n32532 , n24898 , n23015 );
    and g35431 ( n26769 , n33155 , n34334 );
    or g35432 ( n27204 , n6988 , n13414 );
    not g35433 ( n105 , n5964 );
    or g35434 ( n20314 , n41013 , n17332 );
    not g35435 ( n22967 , n14394 );
    not g35436 ( n1126 , n38037 );
    and g35437 ( n29381 , n14451 , n8702 );
    not g35438 ( n231 , n12942 );
    or g35439 ( n41915 , n29011 , n25504 );
    or g35440 ( n1397 , n29027 , n36563 );
    not g35441 ( n19360 , n28873 );
    or g35442 ( n41988 , n23271 , n17109 );
    or g35443 ( n26484 , n13785 , n37902 );
    or g35444 ( n6680 , n6101 , n7243 );
    or g35445 ( n26074 , n15215 , n38564 );
    and g35446 ( n2885 , n6927 , n10173 );
    nor g35447 ( n20324 , n39544 , n16136 );
    not g35448 ( n16998 , n38898 );
    nor g35449 ( n5704 , n21652 , n19733 );
    or g35450 ( n23395 , n19221 , n15759 );
    not g35451 ( n40635 , n4296 );
    nor g35452 ( n31367 , n38879 , n22762 );
    and g35453 ( n26634 , n33348 , n21708 );
    nor g35454 ( n27466 , n30262 , n18882 );
    nor g35455 ( n36245 , n25261 , n14554 );
    not g35456 ( n15179 , n24153 );
    nor g35457 ( n10722 , n40995 , n1024 );
    xnor g35458 ( n1128 , n35727 , n31420 );
    not g35459 ( n21108 , n9328 );
    and g35460 ( n16545 , n27932 , n16921 );
    or g35461 ( n2560 , n28883 , n30194 );
    or g35462 ( n4426 , n7502 , n30939 );
    and g35463 ( n2781 , n29804 , n26954 );
    xnor g35464 ( n34388 , n9180 , n31713 );
    or g35465 ( n13168 , n8594 , n29750 );
    xnor g35466 ( n35805 , n10195 , n6833 );
    not g35467 ( n18143 , n13955 );
    or g35468 ( n4647 , n26845 , n17930 );
    xnor g35469 ( n30615 , n11220 , n6765 );
    xnor g35470 ( n17558 , n37074 , n18073 );
    and g35471 ( n10121 , n8393 , n35560 );
    xnor g35472 ( n11886 , n26579 , n4478 );
    not g35473 ( n23028 , n31209 );
    or g35474 ( n25403 , n36734 , n40014 );
    or g35475 ( n5384 , n7356 , n29259 );
    xnor g35476 ( n7990 , n7489 , n25304 );
    and g35477 ( n35571 , n27731 , n42371 );
    and g35478 ( n18300 , n20782 , n679 );
    and g35479 ( n41854 , n7390 , n3492 );
    and g35480 ( n41788 , n31087 , n42139 );
    xnor g35481 ( n24339 , n12146 , n35673 );
    not g35482 ( n41124 , n6242 );
    or g35483 ( n2890 , n13887 , n12293 );
    xnor g35484 ( n8437 , n24998 , n9012 );
    xnor g35485 ( n20791 , n41013 , n5567 );
    or g35486 ( n22897 , n20750 , n42694 );
    and g35487 ( n29011 , n14466 , n11233 );
    or g35488 ( n42094 , n31049 , n3715 );
    and g35489 ( n26780 , n3383 , n2115 );
    not g35490 ( n38862 , n11881 );
    xnor g35491 ( n32013 , n40 , n29173 );
    nor g35492 ( n12480 , n36117 , n26391 );
    not g35493 ( n31025 , n31419 );
    or g35494 ( n14277 , n25383 , n23492 );
    and g35495 ( n38036 , n25082 , n20690 );
    and g35496 ( n3271 , n37325 , n32482 );
    and g35497 ( n22864 , n26484 , n16246 );
    not g35498 ( n24504 , n24447 );
    and g35499 ( n10719 , n9922 , n8181 );
    or g35500 ( n3243 , n3698 , n35369 );
    and g35501 ( n12588 , n5874 , n40091 );
    and g35502 ( n29172 , n34913 , n33818 );
    nor g35503 ( n4955 , n20554 , n7032 );
    xnor g35504 ( n39693 , n2338 , n32038 );
    nor g35505 ( n6701 , n42553 , n17065 );
    or g35506 ( n11360 , n14825 , n42033 );
    xnor g35507 ( n39356 , n6625 , n16115 );
    not g35508 ( n22635 , n41054 );
    or g35509 ( n31687 , n15040 , n1225 );
    or g35510 ( n26552 , n1226 , n6273 );
    not g35511 ( n31609 , n3517 );
    or g35512 ( n6076 , n7907 , n32535 );
    or g35513 ( n13267 , n40760 , n2972 );
    not g35514 ( n34414 , n8504 );
    or g35515 ( n21270 , n36718 , n10399 );
    xnor g35516 ( n16323 , n23944 , n21265 );
    or g35517 ( n32559 , n5175 , n22289 );
    xnor g35518 ( n34611 , n17038 , n34829 );
    or g35519 ( n28042 , n26858 , n6051 );
    or g35520 ( n42091 , n35773 , n41553 );
    xnor g35521 ( n25014 , n22093 , n27118 );
    or g35522 ( n25502 , n20106 , n3311 );
    or g35523 ( n1377 , n4379 , n1289 );
    or g35524 ( n11300 , n16780 , n38123 );
    or g35525 ( n15993 , n30254 , n34297 );
    or g35526 ( n26901 , n28774 , n12379 );
    or g35527 ( n18818 , n5931 , n32768 );
    or g35528 ( n7317 , n32472 , n20625 );
    or g35529 ( n3 , n24554 , n14407 );
    not g35530 ( n41301 , n32526 );
    or g35531 ( n33471 , n4283 , n40396 );
    nor g35532 ( n29063 , n15732 , n21477 );
    xnor g35533 ( n17259 , n13743 , n30100 );
    xnor g35534 ( n29285 , n26 , n18269 );
    not g35535 ( n14871 , n7360 );
    xnor g35536 ( n10276 , n26579 , n42537 );
    and g35537 ( n24993 , n34116 , n3104 );
    or g35538 ( n7767 , n14973 , n20145 );
    xnor g35539 ( n1494 , n41013 , n19691 );
    or g35540 ( n11744 , n39991 , n35710 );
    and g35541 ( n16412 , n33687 , n3889 );
    or g35542 ( n41123 , n5964 , n4767 );
    or g35543 ( n9008 , n5941 , n21292 );
    or g35544 ( n25645 , n31278 , n34744 );
    nor g35545 ( n36604 , n34419 , n24953 );
    nor g35546 ( n11568 , n30606 , n7993 );
    or g35547 ( n32533 , n14143 , n40140 );
    and g35548 ( n13645 , n21623 , n29910 );
    nor g35549 ( n9821 , n7968 , n8230 );
    nor g35550 ( n15434 , n14467 , n12783 );
    and g35551 ( n25024 , n15772 , n38194 );
    or g35552 ( n20500 , n28706 , n40713 );
    nor g35553 ( n2035 , n7074 , n30572 );
    or g35554 ( n2287 , n39632 , n1745 );
    or g35555 ( n13641 , n30608 , n2239 );
    and g35556 ( n274 , n32624 , n4704 );
    or g35557 ( n22138 , n34516 , n33297 );
    xnor g35558 ( n4496 , n3769 , n1210 );
    xnor g35559 ( n20508 , n32209 , n37988 );
    and g35560 ( n32811 , n27939 , n8227 );
    or g35561 ( n40739 , n38776 , n31804 );
    or g35562 ( n34507 , n33951 , n15216 );
    and g35563 ( n41333 , n23875 , n18592 );
    xnor g35564 ( n22805 , n30631 , n35789 );
    nor g35565 ( n543 , n41529 , n36655 );
    or g35566 ( n13864 , n12105 , n38544 );
    not g35567 ( n13305 , n28570 );
    or g35568 ( n6127 , n18798 , n7 );
    or g35569 ( n843 , n32068 , n27237 );
    not g35570 ( n12837 , n31694 );
    xnor g35571 ( n40407 , n11614 , n18541 );
    or g35572 ( n19713 , n3306 , n6903 );
    or g35573 ( n10642 , n4033 , n29920 );
    and g35574 ( n9009 , n37386 , n37293 );
    and g35575 ( n24855 , n34532 , n509 );
    and g35576 ( n16556 , n25268 , n26134 );
    or g35577 ( n30729 , n37364 , n39813 );
    nor g35578 ( n8433 , n27681 , n4437 );
    and g35579 ( n32708 , n26412 , n6030 );
    xnor g35580 ( n33263 , n17562 , n31024 );
    xnor g35581 ( n39808 , n38789 , n16268 );
    or g35582 ( n19544 , n12193 , n27561 );
    or g35583 ( n34811 , n6593 , n38800 );
    or g35584 ( n17496 , n34684 , n560 );
    or g35585 ( n8261 , n14899 , n17404 );
    or g35586 ( n31586 , n7743 , n17881 );
    or g35587 ( n9093 , n5549 , n1906 );
    nor g35588 ( n32933 , n26597 , n28184 );
    or g35589 ( n19139 , n19808 , n41681 );
    nor g35590 ( n17063 , n38157 , n34415 );
    or g35591 ( n37268 , n4686 , n15095 );
    xnor g35592 ( n33518 , n27237 , n33981 );
    or g35593 ( n40991 , n41411 , n16876 );
    or g35594 ( n2771 , n9451 , n10071 );
    and g35595 ( n42023 , n11100 , n200 );
    and g35596 ( n40062 , n12948 , n14852 );
    nor g35597 ( n21118 , n35965 , n9514 );
    or g35598 ( n2391 , n5017 , n22592 );
    nor g35599 ( n27146 , n8251 , n11654 );
    and g35600 ( n9199 , n35741 , n12760 );
    or g35601 ( n8935 , n38150 , n1511 );
    nor g35602 ( n5063 , n35264 , n5484 );
    nor g35603 ( n31059 , n2261 , n4298 );
    and g35604 ( n32473 , n3722 , n17338 );
    or g35605 ( n40511 , n17167 , n21715 );
    not g35606 ( n20261 , n27604 );
    or g35607 ( n36797 , n15438 , n31361 );
    or g35608 ( n9453 , n24650 , n6043 );
    nor g35609 ( n8006 , n42272 , n6937 );
    or g35610 ( n35061 , n14927 , n2597 );
    and g35611 ( n5025 , n34494 , n12862 );
    and g35612 ( n17057 , n18724 , n24343 );
    or g35613 ( n25264 , n4670 , n34227 );
    nor g35614 ( n462 , n38157 , n38465 );
    and g35615 ( n16115 , n7720 , n6384 );
    xnor g35616 ( n36542 , n14125 , n9692 );
    and g35617 ( n18494 , n38267 , n33477 );
    and g35618 ( n15580 , n12358 , n25229 );
    not g35619 ( n22799 , n42550 );
    and g35620 ( n15144 , n17300 , n29315 );
    not g35621 ( n9005 , n33978 );
    nor g35622 ( n35046 , n20804 , n24431 );
    nor g35623 ( n16452 , n16500 , n40227 );
    not g35624 ( n14976 , n8892 );
    not g35625 ( n42844 , n27476 );
    and g35626 ( n1520 , n10085 , n40937 );
    not g35627 ( n19578 , n36521 );
    nor g35628 ( n31954 , n9326 , n7438 );
    nor g35629 ( n20504 , n27279 , n6005 );
    nor g35630 ( n34066 , n17267 , n35124 );
    or g35631 ( n27061 , n38761 , n26025 );
    and g35632 ( n18606 , n29995 , n612 );
    not g35633 ( n17344 , n9069 );
    xnor g35634 ( n5922 , n5144 , n34549 );
    xnor g35635 ( n21385 , n39531 , n39596 );
    or g35636 ( n28245 , n24909 , n30652 );
    not g35637 ( n35320 , n37451 );
    or g35638 ( n1179 , n40999 , n425 );
    or g35639 ( n25023 , n26067 , n41288 );
    nor g35640 ( n11466 , n18839 , n31230 );
    not g35641 ( n25882 , n5990 );
    not g35642 ( n13904 , n20309 );
    nor g35643 ( n21276 , n7228 , n36450 );
    and g35644 ( n23756 , n4640 , n36768 );
    or g35645 ( n23725 , n32902 , n38552 );
    or g35646 ( n38513 , n26522 , n27037 );
    not g35647 ( n6179 , n36137 );
    or g35648 ( n7788 , n22667 , n15079 );
    or g35649 ( n2030 , n36117 , n23411 );
    or g35650 ( n4409 , n4228 , n8451 );
    not g35651 ( n19400 , n288 );
    or g35652 ( n18434 , n8361 , n28959 );
    and g35653 ( n14380 , n38458 , n9006 );
    nor g35654 ( n39297 , n16848 , n3508 );
    and g35655 ( n37096 , n34273 , n29893 );
    not g35656 ( n24626 , n40078 );
    or g35657 ( n36386 , n9122 , n12011 );
    or g35658 ( n2475 , n21871 , n22794 );
    or g35659 ( n3159 , n8409 , n33754 );
    or g35660 ( n11700 , n1153 , n14001 );
    or g35661 ( n19716 , n21438 , n16577 );
    xnor g35662 ( n34677 , n14070 , n19750 );
    and g35663 ( n8511 , n0 , n23721 );
    or g35664 ( n16230 , n5197 , n7783 );
    xnor g35665 ( n10536 , n42064 , n35949 );
    or g35666 ( n38229 , n10030 , n6545 );
    or g35667 ( n42883 , n31271 , n35544 );
    not g35668 ( n8122 , n25024 );
    xnor g35669 ( n27588 , n27035 , n26193 );
    or g35670 ( n21486 , n2786 , n40746 );
    or g35671 ( n16526 , n20752 , n26943 );
    not g35672 ( n32312 , n18062 );
    xnor g35673 ( n23180 , n5891 , n35275 );
    and g35674 ( n41909 , n14024 , n505 );
    and g35675 ( n5075 , n10905 , n15041 );
    or g35676 ( n8480 , n39039 , n34949 );
    or g35677 ( n8411 , n12233 , n42201 );
    xnor g35678 ( n13461 , n23080 , n24528 );
    nor g35679 ( n6109 , n35074 , n23466 );
    xnor g35680 ( n36215 , n32048 , n944 );
    and g35681 ( n9049 , n33534 , n41808 );
    and g35682 ( n10168 , n23134 , n233 );
    nor g35683 ( n41049 , n21134 , n11530 );
    and g35684 ( n26783 , n14471 , n11101 );
    and g35685 ( n15911 , n6729 , n42681 );
    or g35686 ( n16616 , n42392 , n4703 );
    and g35687 ( n2818 , n13201 , n21949 );
    or g35688 ( n25071 , n19619 , n11159 );
    and g35689 ( n14386 , n6913 , n20462 );
    not g35690 ( n18910 , n30017 );
    or g35691 ( n2940 , n27952 , n8959 );
    and g35692 ( n20604 , n42684 , n10334 );
    not g35693 ( n37980 , n29949 );
    not g35694 ( n9697 , n15344 );
    nor g35695 ( n5151 , n33190 , n9089 );
    xnor g35696 ( n25239 , n42866 , n9587 );
    or g35697 ( n16531 , n457 , n5701 );
    xnor g35698 ( n29823 , n36938 , n4169 );
    not g35699 ( n37540 , n14008 );
    not g35700 ( n33220 , n38466 );
    or g35701 ( n1720 , n20790 , n12220 );
    not g35702 ( n35025 , n22339 );
    and g35703 ( n10537 , n2498 , n17587 );
    or g35704 ( n901 , n29051 , n3728 );
    nor g35705 ( n9439 , n31596 , n25289 );
    or g35706 ( n31034 , n19015 , n34652 );
    or g35707 ( n3173 , n22350 , n38196 );
    nor g35708 ( n26853 , n20479 , n14123 );
    or g35709 ( n11280 , n2356 , n29126 );
    xnor g35710 ( n4983 , n25043 , n40317 );
    and g35711 ( n37751 , n16853 , n33460 );
    and g35712 ( n7942 , n16750 , n32595 );
    not g35713 ( n25591 , n16482 );
    or g35714 ( n127 , n6115 , n20914 );
    not g35715 ( n11679 , n36468 );
    and g35716 ( n30381 , n19817 , n24678 );
    or g35717 ( n40081 , n635 , n6024 );
    nor g35718 ( n20969 , n6179 , n448 );
    or g35719 ( n27429 , n122 , n24839 );
    and g35720 ( n16495 , n33751 , n42784 );
    and g35721 ( n5529 , n30359 , n21189 );
    or g35722 ( n29882 , n991 , n34590 );
    or g35723 ( n36109 , n18532 , n29118 );
    or g35724 ( n25203 , n34633 , n32194 );
    not g35725 ( n11109 , n31089 );
    not g35726 ( n22545 , n27230 );
    and g35727 ( n225 , n26768 , n40142 );
    and g35728 ( n9920 , n9845 , n23240 );
    not g35729 ( n12600 , n7786 );
    and g35730 ( n13303 , n4007 , n3261 );
    nor g35731 ( n32832 , n33706 , n40607 );
    or g35732 ( n42382 , n23665 , n38006 );
    or g35733 ( n41984 , n29803 , n25578 );
    or g35734 ( n35532 , n39635 , n20054 );
    or g35735 ( n15316 , n33768 , n32256 );
    nor g35736 ( n8486 , n25588 , n3506 );
    and g35737 ( n42913 , n30277 , n33470 );
    or g35738 ( n29002 , n4702 , n16410 );
    and g35739 ( n35781 , n19592 , n9378 );
    or g35740 ( n42443 , n14831 , n21630 );
    and g35741 ( n38674 , n28573 , n29802 );
    nor g35742 ( n36400 , n38654 , n17837 );
    and g35743 ( n27226 , n31934 , n41016 );
    or g35744 ( n39270 , n35738 , n16891 );
    not g35745 ( n10874 , n6926 );
    and g35746 ( n7807 , n31631 , n10862 );
    or g35747 ( n1835 , n39076 , n17152 );
    or g35748 ( n35537 , n13734 , n25277 );
    or g35749 ( n26231 , n36370 , n39393 );
    xnor g35750 ( n23196 , n21652 , n14982 );
    nor g35751 ( n36498 , n26617 , n27267 );
    nor g35752 ( n24658 , n18625 , n23009 );
    xnor g35753 ( n3413 , n37163 , n23743 );
    and g35754 ( n41973 , n21959 , n31118 );
    nor g35755 ( n10391 , n4173 , n19421 );
    or g35756 ( n21222 , n38512 , n20459 );
    xnor g35757 ( n41855 , n24634 , n37063 );
    not g35758 ( n27666 , n22533 );
    and g35759 ( n7314 , n38295 , n25232 );
    and g35760 ( n20814 , n10466 , n13570 );
    not g35761 ( n8784 , n21104 );
    nor g35762 ( n39768 , n39456 , n1190 );
    not g35763 ( n27756 , n21870 );
    and g35764 ( n13124 , n42283 , n24066 );
    not g35765 ( n15505 , n41253 );
    or g35766 ( n38248 , n22440 , n37220 );
    or g35767 ( n9664 , n36919 , n12904 );
    not g35768 ( n11995 , n25533 );
    and g35769 ( n5456 , n9742 , n16290 );
    not g35770 ( n37640 , n716 );
    not g35771 ( n9290 , n2279 );
    and g35772 ( n18279 , n9849 , n602 );
    and g35773 ( n15642 , n40691 , n13914 );
    not g35774 ( n28154 , n36337 );
    or g35775 ( n26022 , n40206 , n22240 );
    or g35776 ( n24354 , n18587 , n39128 );
    and g35777 ( n20294 , n11848 , n1443 );
    or g35778 ( n39280 , n584 , n34939 );
    and g35779 ( n21390 , n15 , n22394 );
    nor g35780 ( n4885 , n39950 , n31505 );
    or g35781 ( n5032 , n28962 , n39138 );
    not g35782 ( n33917 , n11409 );
    xnor g35783 ( n38827 , n4558 , n33048 );
    not g35784 ( n36134 , n21517 );
    and g35785 ( n28924 , n29279 , n25086 );
    and g35786 ( n9067 , n32322 , n41219 );
    and g35787 ( n9044 , n1239 , n11776 );
    not g35788 ( n13637 , n4697 );
    nor g35789 ( n28046 , n2387 , n39904 );
    or g35790 ( n36711 , n5359 , n21510 );
    or g35791 ( n32454 , n134 , n22885 );
    or g35792 ( n34719 , n30432 , n17383 );
    xnor g35793 ( n25074 , n22263 , n11597 );
    or g35794 ( n3497 , n8808 , n6290 );
    xnor g35795 ( n11622 , n6714 , n40572 );
    not g35796 ( n15823 , n14962 );
    or g35797 ( n21477 , n41930 , n11617 );
    not g35798 ( n6831 , n42539 );
    and g35799 ( n9633 , n4260 , n14007 );
    not g35800 ( n10996 , n19925 );
    nor g35801 ( n38557 , n35289 , n39373 );
    or g35802 ( n3122 , n20932 , n23806 );
    or g35803 ( n8867 , n10823 , n34317 );
    or g35804 ( n33786 , n25040 , n30392 );
    and g35805 ( n26491 , n1323 , n18743 );
    and g35806 ( n27739 , n16549 , n22754 );
    and g35807 ( n3428 , n39947 , n41023 );
    or g35808 ( n29639 , n22920 , n42913 );
    and g35809 ( n6363 , n38668 , n19761 );
    and g35810 ( n614 , n9736 , n11014 );
    not g35811 ( n5921 , n8995 );
    xnor g35812 ( n16850 , n11972 , n33267 );
    not g35813 ( n3657 , n22185 );
    or g35814 ( n6981 , n34863 , n19842 );
    and g35815 ( n31591 , n24005 , n33841 );
    or g35816 ( n14438 , n6503 , n30533 );
    nor g35817 ( n28736 , n41761 , n19333 );
    or g35818 ( n8974 , n12955 , n3305 );
    not g35819 ( n17669 , n3573 );
    not g35820 ( n9120 , n36315 );
    or g35821 ( n989 , n36531 , n22143 );
    xnor g35822 ( n21308 , n17159 , n18399 );
    or g35823 ( n5178 , n35386 , n39875 );
    or g35824 ( n20074 , n14756 , n30676 );
    or g35825 ( n30363 , n2288 , n5023 );
    nor g35826 ( n8765 , n17372 , n18302 );
    and g35827 ( n11800 , n8894 , n13922 );
    xnor g35828 ( n26665 , n8439 , n572 );
    and g35829 ( n31159 , n41883 , n30797 );
    or g35830 ( n31002 , n38591 , n35432 );
    or g35831 ( n11107 , n8219 , n33782 );
    xnor g35832 ( n18853 , n35733 , n33823 );
    nor g35833 ( n25890 , n6640 , n19291 );
    not g35834 ( n26996 , n366 );
    not g35835 ( n33715 , n15618 );
    and g35836 ( n7768 , n27467 , n1898 );
    or g35837 ( n16570 , n42512 , n27315 );
    not g35838 ( n26 , n19607 );
    or g35839 ( n39564 , n19221 , n40405 );
    or g35840 ( n8137 , n26005 , n6001 );
    and g35841 ( n34029 , n36451 , n21062 );
    xnor g35842 ( n38666 , n34731 , n6946 );
    xnor g35843 ( n31881 , n29858 , n26604 );
    and g35844 ( n9344 , n10630 , n1929 );
    and g35845 ( n1996 , n19368 , n38195 );
    and g35846 ( n17221 , n38871 , n26550 );
    nor g35847 ( n26965 , n5622 , n8850 );
    or g35848 ( n10590 , n12852 , n5148 );
    or g35849 ( n28271 , n20033 , n34972 );
    or g35850 ( n31344 , n9181 , n33145 );
    and g35851 ( n31228 , n14704 , n31995 );
    or g35852 ( n4618 , n10598 , n37484 );
    nor g35853 ( n20246 , n6843 , n7733 );
    or g35854 ( n28657 , n33012 , n29996 );
    not g35855 ( n28595 , n19120 );
    and g35856 ( n13665 , n24576 , n4605 );
    and g35857 ( n36930 , n38730 , n19320 );
    or g35858 ( n22330 , n14545 , n27127 );
    not g35859 ( n38852 , n18983 );
    and g35860 ( n27121 , n9769 , n9469 );
    not g35861 ( n42702 , n6820 );
    and g35862 ( n4797 , n38722 , n27442 );
    xnor g35863 ( n13148 , n17155 , n38625 );
    or g35864 ( n31663 , n33556 , n7329 );
    and g35865 ( n9873 , n14497 , n16819 );
    and g35866 ( n29043 , n37571 , n9985 );
    or g35867 ( n16991 , n26626 , n10268 );
    not g35868 ( n8588 , n31364 );
    or g35869 ( n2206 , n23509 , n3227 );
    or g35870 ( n42362 , n4669 , n159 );
    or g35871 ( n9056 , n4154 , n3554 );
    nor g35872 ( n8347 , n17193 , n7442 );
    xnor g35873 ( n36083 , n18736 , n3853 );
    and g35874 ( n13767 , n28443 , n23442 );
    and g35875 ( n37395 , n22362 , n42040 );
    or g35876 ( n12986 , n1439 , n23236 );
    and g35877 ( n6945 , n41235 , n4620 );
    and g35878 ( n8792 , n18773 , n19216 );
    not g35879 ( n23948 , n35766 );
    and g35880 ( n5623 , n30391 , n41155 );
    and g35881 ( n10571 , n18013 , n31053 );
    and g35882 ( n9862 , n22140 , n6695 );
    or g35883 ( n39555 , n38119 , n40424 );
    not g35884 ( n39098 , n15956 );
    nor g35885 ( n24276 , n20289 , n34121 );
    and g35886 ( n25470 , n6947 , n12793 );
    not g35887 ( n962 , n15504 );
    nor g35888 ( n19027 , n11380 , n33431 );
    not g35889 ( n14732 , n11506 );
    and g35890 ( n7703 , n27736 , n21734 );
    not g35891 ( n35322 , n12224 );
    or g35892 ( n1037 , n29247 , n26824 );
    nor g35893 ( n24904 , n5441 , n3138 );
    nor g35894 ( n31768 , n34778 , n18679 );
    nor g35895 ( n16164 , n32042 , n24383 );
    xnor g35896 ( n28356 , n5144 , n4883 );
    or g35897 ( n42860 , n122 , n12688 );
    or g35898 ( n14303 , n28231 , n10304 );
    nor g35899 ( n6136 , n13697 , n42809 );
    or g35900 ( n34823 , n5204 , n17032 );
    or g35901 ( n42078 , n4492 , n23435 );
    and g35902 ( n12994 , n1109 , n22749 );
    or g35903 ( n10944 , n40742 , n20064 );
    or g35904 ( n9347 , n20932 , n4243 );
    or g35905 ( n30833 , n9885 , n4738 );
    xnor g35906 ( n23066 , n31989 , n6595 );
    not g35907 ( n29545 , n9312 );
    or g35908 ( n39261 , n9817 , n5421 );
    and g35909 ( n40909 , n15260 , n8867 );
    or g35910 ( n38527 , n1799 , n6288 );
    not g35911 ( n928 , n13857 );
    and g35912 ( n10728 , n24474 , n34062 );
    or g35913 ( n20929 , n18546 , n26229 );
    and g35914 ( n36754 , n38198 , n18041 );
    xnor g35915 ( n25939 , n8499 , n14679 );
    not g35916 ( n35695 , n9312 );
    xnor g35917 ( n17430 , n21133 , n27538 );
    nor g35918 ( n18378 , n30754 , n23807 );
    or g35919 ( n36340 , n40978 , n23743 );
    or g35920 ( n15180 , n33026 , n13665 );
    or g35921 ( n11056 , n15979 , n30931 );
    nor g35922 ( n21426 , n19599 , n1583 );
    or g35923 ( n39750 , n16939 , n31883 );
    xnor g35924 ( n13502 , n1464 , n20901 );
    xnor g35925 ( n33198 , n28458 , n22203 );
    or g35926 ( n42170 , n23179 , n8175 );
    xnor g35927 ( n4392 , n38749 , n32681 );
    or g35928 ( n37528 , n9829 , n26370 );
    or g35929 ( n40469 , n11411 , n34749 );
    not g35930 ( n383 , n2135 );
    and g35931 ( n9561 , n11740 , n22264 );
    or g35932 ( n6758 , n4926 , n36577 );
    nor g35933 ( n7860 , n19045 , n2190 );
    nor g35934 ( n2776 , n21248 , n35587 );
    xnor g35935 ( n39249 , n27213 , n17120 );
    not g35936 ( n41619 , n42738 );
    nor g35937 ( n7670 , n23572 , n27936 );
    or g35938 ( n13672 , n7885 , n15375 );
    and g35939 ( n11233 , n12869 , n11112 );
    and g35940 ( n26823 , n21386 , n40511 );
    or g35941 ( n29119 , n8009 , n25059 );
    not g35942 ( n19813 , n13523 );
    or g35943 ( n29728 , n30965 , n36348 );
    nor g35944 ( n31223 , n34759 , n27973 );
    and g35945 ( n22350 , n2975 , n29284 );
    not g35946 ( n1768 , n6442 );
    or g35947 ( n19916 , n42469 , n12732 );
    xnor g35948 ( n12491 , n2896 , n17744 );
    xnor g35949 ( n25359 , n5344 , n33207 );
    and g35950 ( n36528 , n17374 , n9522 );
    not g35951 ( n14242 , n41603 );
    nor g35952 ( n24044 , n39174 , n36169 );
    and g35953 ( n40838 , n22873 , n27636 );
    nor g35954 ( n3403 , n3581 , n28468 );
    or g35955 ( n10583 , n1507 , n32668 );
    xnor g35956 ( n10043 , n9180 , n22696 );
    nor g35957 ( n31551 , n24156 , n14998 );
    nor g35958 ( n15692 , n29538 , n26165 );
    and g35959 ( n19784 , n4443 , n25106 );
    and g35960 ( n30887 , n28973 , n36773 );
    not g35961 ( n42379 , n40959 );
    nor g35962 ( n42613 , n2199 , n39502 );
    or g35963 ( n18191 , n27984 , n37733 );
    and g35964 ( n29775 , n33570 , n4875 );
    xnor g35965 ( n31363 , n38105 , n16631 );
    or g35966 ( n25698 , n14022 , n5462 );
    and g35967 ( n21500 , n19725 , n18325 );
    or g35968 ( n26539 , n37520 , n40228 );
    or g35969 ( n35622 , n2183 , n37803 );
    and g35970 ( n33151 , n31633 , n9565 );
    or g35971 ( n19505 , n35452 , n31747 );
    xnor g35972 ( n20999 , n39639 , n21507 );
    or g35973 ( n8417 , n21760 , n27127 );
    or g35974 ( n34867 , n31575 , n11762 );
    or g35975 ( n21124 , n28991 , n10646 );
    or g35976 ( n35196 , n11106 , n24887 );
    or g35977 ( n15735 , n5419 , n32839 );
    and g35978 ( n10155 , n23104 , n34903 );
    and g35979 ( n2476 , n18487 , n30559 );
    or g35980 ( n2522 , n7196 , n18567 );
    or g35981 ( n22234 , n38293 , n8029 );
    and g35982 ( n30247 , n5447 , n17257 );
    and g35983 ( n15172 , n3494 , n18213 );
    xnor g35984 ( n19887 , n3769 , n8601 );
    or g35985 ( n15142 , n9208 , n4355 );
    and g35986 ( n26737 , n12131 , n16005 );
    and g35987 ( n7665 , n5062 , n4720 );
    nor g35988 ( n36075 , n23745 , n10468 );
    not g35989 ( n33222 , n40006 );
    or g35990 ( n16812 , n19535 , n28746 );
    xnor g35991 ( n42203 , n18696 , n32437 );
    xnor g35992 ( n2076 , n4501 , n9390 );
    or g35993 ( n9871 , n1507 , n38554 );
    and g35994 ( n12937 , n32703 , n15073 );
    xnor g35995 ( n19835 , n20310 , n19318 );
    not g35996 ( n21721 , n27987 );
    or g35997 ( n21247 , n35750 , n22802 );
    and g35998 ( n38884 , n10120 , n32955 );
    or g35999 ( n23850 , n24626 , n10680 );
    nor g36000 ( n14474 , n4767 , n4483 );
    or g36001 ( n26967 , n15403 , n18197 );
    and g36002 ( n40153 , n26036 , n41680 );
    or g36003 ( n25497 , n21025 , n13750 );
    or g36004 ( n37821 , n25704 , n24232 );
    and g36005 ( n11805 , n32556 , n3183 );
    and g36006 ( n11229 , n38631 , n34405 );
    xnor g36007 ( n6939 , n40337 , n31211 );
    or g36008 ( n219 , n33981 , n3062 );
    or g36009 ( n5056 , n31903 , n14278 );
    or g36010 ( n42129 , n25721 , n20654 );
    nor g36011 ( n34447 , n10460 , n16092 );
    nor g36012 ( n8064 , n33620 , n29134 );
    or g36013 ( n8266 , n28373 , n18311 );
    or g36014 ( n26392 , n3694 , n26789 );
    nor g36015 ( n591 , n35301 , n3235 );
    or g36016 ( n36141 , n25323 , n38758 );
    not g36017 ( n24588 , n11682 );
    not g36018 ( n10687 , n28529 );
    not g36019 ( n38362 , n13584 );
    or g36020 ( n7656 , n4086 , n399 );
    xnor g36021 ( n30512 , n40 , n40930 );
    and g36022 ( n23528 , n5776 , n29626 );
    not g36023 ( n3980 , n9421 );
    or g36024 ( n29050 , n1355 , n36671 );
    or g36025 ( n40234 , n8466 , n792 );
    and g36026 ( n30184 , n32057 , n2557 );
    and g36027 ( n17013 , n33937 , n42341 );
    nor g36028 ( n37445 , n32589 , n28216 );
    or g36029 ( n38809 , n4717 , n29829 );
    nor g36030 ( n20306 , n21339 , n3766 );
    or g36031 ( n31835 , n19337 , n17802 );
    nor g36032 ( n26173 , n23040 , n37365 );
    xnor g36033 ( n10282 , n35727 , n12746 );
    nor g36034 ( n38254 , n6176 , n21159 );
    or g36035 ( n27550 , n25066 , n27739 );
    or g36036 ( n8632 , n34955 , n39294 );
    nor g36037 ( n35407 , n24549 , n11507 );
    nor g36038 ( n31794 , n36932 , n4824 );
    not g36039 ( n19531 , n3084 );
    xnor g36040 ( n17413 , n34731 , n29065 );
    not g36041 ( n122 , n13805 );
    or g36042 ( n12707 , n21542 , n34070 );
    or g36043 ( n36124 , n11930 , n32439 );
    nor g36044 ( n36751 , n15611 , n38729 );
    not g36045 ( n39279 , n29163 );
    not g36046 ( n9171 , n13512 );
    or g36047 ( n25841 , n27735 , n35382 );
    not g36048 ( n21095 , n38469 );
    xnor g36049 ( n31318 , n31323 , n34292 );
    not g36050 ( n19104 , n32982 );
    nor g36051 ( n41263 , n32408 , n16509 );
    nor g36052 ( n9297 , n29392 , n42236 );
    nor g36053 ( n36934 , n26844 , n25244 );
    or g36054 ( n37407 , n33432 , n19848 );
    xnor g36055 ( n22041 , n4511 , n18482 );
    or g36056 ( n7923 , n36296 , n18501 );
    or g36057 ( n16193 , n39769 , n8318 );
    and g36058 ( n7582 , n41773 , n3860 );
    and g36059 ( n22584 , n37907 , n31714 );
    or g36060 ( n10466 , n39388 , n4039 );
    and g36061 ( n10700 , n29074 , n27050 );
    or g36062 ( n18714 , n12498 , n36859 );
    not g36063 ( n26548 , n31376 );
    or g36064 ( n10777 , n18388 , n18511 );
    and g36065 ( n31569 , n34635 , n33554 );
    or g36066 ( n31774 , n15000 , n41265 );
    not g36067 ( n14813 , n32001 );
    not g36068 ( n11468 , n26976 );
    or g36069 ( n25984 , n11487 , n31503 );
    and g36070 ( n20985 , n29729 , n20253 );
    not g36071 ( n30582 , n25960 );
    or g36072 ( n16386 , n37916 , n33575 );
    and g36073 ( n18002 , n27697 , n3499 );
    or g36074 ( n33966 , n36956 , n23444 );
    nor g36075 ( n17418 , n12990 , n2483 );
    and g36076 ( n14061 , n762 , n27839 );
    or g36077 ( n29642 , n17084 , n12395 );
    not g36078 ( n29306 , n7535 );
    xnor g36079 ( n9175 , n18466 , n5847 );
    or g36080 ( n17335 , n28241 , n33149 );
    or g36081 ( n29444 , n11527 , n13235 );
    or g36082 ( n23866 , n26699 , n32357 );
    nor g36083 ( n25792 , n4644 , n11473 );
    not g36084 ( n15740 , n11611 );
    nor g36085 ( n7912 , n15858 , n20113 );
    not g36086 ( n4304 , n5940 );
    or g36087 ( n4059 , n21038 , n22032 );
    or g36088 ( n9211 , n34575 , n18725 );
    or g36089 ( n16157 , n8494 , n21031 );
    or g36090 ( n42197 , n6773 , n32456 );
    not g36091 ( n31471 , n24000 );
    or g36092 ( n3365 , n12495 , n3028 );
    and g36093 ( n15353 , n20314 , n34583 );
    not g36094 ( n24163 , n1903 );
    xnor g36095 ( n13893 , n14649 , n13594 );
    or g36096 ( n33911 , n10070 , n21006 );
    nor g36097 ( n22144 , n9533 , n15205 );
    or g36098 ( n25135 , n19523 , n5216 );
    xnor g36099 ( n2949 , n111 , n30526 );
    not g36100 ( n6161 , n426 );
    or g36101 ( n18740 , n39559 , n24539 );
    nor g36102 ( n17725 , n7001 , n20816 );
    or g36103 ( n36885 , n13580 , n9752 );
    and g36104 ( n2867 , n1427 , n5784 );
    xnor g36105 ( n6455 , n42614 , n29346 );
    or g36106 ( n33177 , n23261 , n8908 );
    or g36107 ( n16154 , n39810 , n40722 );
    or g36108 ( n42252 , n8427 , n4910 );
    xnor g36109 ( n20564 , n26279 , n1144 );
    not g36110 ( n23026 , n22954 );
    or g36111 ( n28338 , n14139 , n1709 );
    xnor g36112 ( n12470 , n31442 , n40128 );
    or g36113 ( n5523 , n328 , n38136 );
    and g36114 ( n41225 , n2431 , n14940 );
    or g36115 ( n20127 , n35767 , n29833 );
    and g36116 ( n5437 , n13507 , n26024 );
    and g36117 ( n10610 , n16396 , n8804 );
    nor g36118 ( n29539 , n16598 , n7977 );
    and g36119 ( n6515 , n31654 , n19410 );
    or g36120 ( n7970 , n37763 , n11572 );
    xnor g36121 ( n24791 , n34735 , n5587 );
    nor g36122 ( n27539 , n16311 , n16430 );
    nor g36123 ( n30815 , n8904 , n13260 );
    not g36124 ( n14988 , n39249 );
    or g36125 ( n41093 , n14407 , n30250 );
    nor g36126 ( n20313 , n35044 , n27115 );
    nor g36127 ( n36919 , n27524 , n34703 );
    or g36128 ( n31846 , n16161 , n37656 );
    or g36129 ( n19417 , n23049 , n1416 );
    or g36130 ( n2351 , n39218 , n419 );
    or g36131 ( n13452 , n30490 , n39902 );
    and g36132 ( n8770 , n24634 , n37063 );
    and g36133 ( n27859 , n10787 , n3249 );
    and g36134 ( n2316 , n18161 , n10551 );
    or g36135 ( n39745 , n17215 , n2507 );
    and g36136 ( n40380 , n11323 , n1276 );
    not g36137 ( n17750 , n10942 );
    nor g36138 ( n30078 , n26831 , n9585 );
    or g36139 ( n35774 , n40697 , n27171 );
    and g36140 ( n41038 , n36791 , n40081 );
    xnor g36141 ( n5659 , n9900 , n24893 );
    nor g36142 ( n30170 , n31565 , n40856 );
    nor g36143 ( n8223 , n33508 , n42372 );
    or g36144 ( n41444 , n27503 , n10768 );
    and g36145 ( n32051 , n10668 , n36440 );
    and g36146 ( n32393 , n35154 , n22465 );
    and g36147 ( n41556 , n14655 , n38394 );
    or g36148 ( n9768 , n40110 , n30419 );
    or g36149 ( n20058 , n40761 , n3583 );
    or g36150 ( n32626 , n27785 , n13146 );
    xnor g36151 ( n8499 , n32632 , n32743 );
    or g36152 ( n25435 , n11445 , n6643 );
    nor g36153 ( n35416 , n37469 , n40187 );
    not g36154 ( n42337 , n8137 );
    not g36155 ( n27954 , n3442 );
    or g36156 ( n13927 , n9807 , n16340 );
    not g36157 ( n1510 , n6491 );
    xnor g36158 ( n8464 , n27836 , n14807 );
    xnor g36159 ( n4662 , n1841 , n3291 );
    or g36160 ( n2986 , n39118 , n5377 );
    and g36161 ( n14422 , n33789 , n15843 );
    xnor g36162 ( n25138 , n38378 , n28732 );
    and g36163 ( n42202 , n32182 , n30387 );
    or g36164 ( n25185 , n8173 , n28096 );
    or g36165 ( n13684 , n37583 , n12220 );
    not g36166 ( n15936 , n34500 );
    or g36167 ( n16878 , n6863 , n11630 );
    or g36168 ( n18573 , n19339 , n24371 );
    not g36169 ( n4301 , n26669 );
    not g36170 ( n25721 , n877 );
    not g36171 ( n31763 , n25807 );
    xnor g36172 ( n22501 , n15219 , n38739 );
    not g36173 ( n41968 , n8197 );
    not g36174 ( n10100 , n17406 );
    not g36175 ( n28464 , n36012 );
    or g36176 ( n15609 , n13603 , n14287 );
    or g36177 ( n29229 , n39699 , n16043 );
    and g36178 ( n42509 , n7368 , n5923 );
    and g36179 ( n3247 , n40251 , n40344 );
    or g36180 ( n41393 , n9939 , n31156 );
    xnor g36181 ( n33517 , n24505 , n24038 );
    nor g36182 ( n7146 , n2318 , n16038 );
    or g36183 ( n18764 , n4140 , n36076 );
    or g36184 ( n9010 , n1292 , n7466 );
    xnor g36185 ( n12848 , n15597 , n17590 );
    xnor g36186 ( n599 , n20237 , n3083 );
    not g36187 ( n36486 , n25607 );
    or g36188 ( n30424 , n25755 , n33997 );
    xnor g36189 ( n39774 , n2839 , n23468 );
    nor g36190 ( n27535 , n5896 , n6254 );
    or g36191 ( n24456 , n7269 , n2269 );
    not g36192 ( n37977 , n40572 );
    xnor g36193 ( n329 , n28979 , n12620 );
    and g36194 ( n8284 , n34929 , n41246 );
    or g36195 ( n26085 , n19259 , n19540 );
    nor g36196 ( n9202 , n36031 , n28340 );
    or g36197 ( n7522 , n9798 , n13701 );
    not g36198 ( n35163 , n13327 );
    nor g36199 ( n36316 , n16598 , n22751 );
    or g36200 ( n33531 , n39665 , n34858 );
    or g36201 ( n11238 , n5298 , n33858 );
    and g36202 ( n15085 , n18864 , n33079 );
    or g36203 ( n40338 , n18775 , n26228 );
    or g36204 ( n39964 , n30007 , n36687 );
    and g36205 ( n31518 , n25174 , n14040 );
    not g36206 ( n39292 , n8565 );
    or g36207 ( n13432 , n1637 , n42584 );
    nor g36208 ( n35177 , n18454 , n41775 );
    or g36209 ( n36614 , n35510 , n20388 );
    and g36210 ( n33768 , n29486 , n35954 );
    or g36211 ( n7666 , n10953 , n8738 );
    not g36212 ( n39412 , n39139 );
    and g36213 ( n12633 , n30079 , n6511 );
    and g36214 ( n17570 , n30145 , n13882 );
    and g36215 ( n41157 , n10047 , n17083 );
    or g36216 ( n30866 , n37840 , n17104 );
    not g36217 ( n15134 , n9651 );
    or g36218 ( n104 , n21170 , n9397 );
    and g36219 ( n6105 , n3777 , n36706 );
    not g36220 ( n31083 , n25734 );
    nor g36221 ( n12511 , n4102 , n17944 );
    xnor g36222 ( n20479 , n16693 , n23035 );
    or g36223 ( n3999 , n32935 , n7667 );
    or g36224 ( n7939 , n11404 , n27673 );
    or g36225 ( n25338 , n35732 , n15869 );
    or g36226 ( n6619 , n21102 , n41913 );
    or g36227 ( n17136 , n14706 , n32566 );
    nor g36228 ( n9489 , n24514 , n38984 );
    or g36229 ( n36471 , n24021 , n33080 );
    not g36230 ( n30446 , n4231 );
    or g36231 ( n33402 , n28666 , n42046 );
    and g36232 ( n27669 , n41492 , n38534 );
    or g36233 ( n8795 , n31434 , n2095 );
    or g36234 ( n23279 , n21214 , n36173 );
    or g36235 ( n13460 , n31677 , n37680 );
    or g36236 ( n33121 , n25536 , n41147 );
    xnor g36237 ( n16721 , n5650 , n24708 );
    not g36238 ( n15565 , n26673 );
    or g36239 ( n32888 , n39443 , n34033 );
    or g36240 ( n19567 , n40643 , n9958 );
    or g36241 ( n29594 , n31459 , n23489 );
    nor g36242 ( n11459 , n26521 , n16171 );
    xnor g36243 ( n665 , n11639 , n5964 );
    or g36244 ( n679 , n24952 , n5408 );
    and g36245 ( n15808 , n25703 , n21952 );
    or g36246 ( n8562 , n13325 , n2034 );
    xnor g36247 ( n4855 , n20323 , n18305 );
    and g36248 ( n42749 , n7377 , n8264 );
    nor g36249 ( n778 , n38922 , n477 );
    not g36250 ( n5656 , n32016 );
    and g36251 ( n26285 , n17308 , n4409 );
    and g36252 ( n16892 , n10344 , n14447 );
    nor g36253 ( n26104 , n15947 , n29180 );
    and g36254 ( n27869 , n35301 , n37773 );
    not g36255 ( n39064 , n8799 );
    or g36256 ( n28012 , n24114 , n19064 );
    or g36257 ( n29992 , n29327 , n14153 );
    and g36258 ( n25395 , n19649 , n19195 );
    or g36259 ( n15850 , n35526 , n25653 );
    not g36260 ( n18174 , n13729 );
    or g36261 ( n4687 , n3511 , n39168 );
    or g36262 ( n11924 , n25136 , n33323 );
    not g36263 ( n21598 , n27964 );
    or g36264 ( n13971 , n28516 , n14931 );
    and g36265 ( n18808 , n33711 , n36775 );
    not g36266 ( n12010 , n38056 );
    or g36267 ( n20434 , n39399 , n7737 );
    nor g36268 ( n9410 , n41234 , n32234 );
    or g36269 ( n29377 , n26791 , n18796 );
    and g36270 ( n36795 , n5747 , n10318 );
    and g36271 ( n37663 , n19381 , n114 );
    xnor g36272 ( n30627 , n7489 , n28425 );
    and g36273 ( n28859 , n42056 , n42718 );
    or g36274 ( n17117 , n7012 , n22608 );
    not g36275 ( n25794 , n23285 );
    or g36276 ( n19013 , n27511 , n34159 );
    not g36277 ( n34184 , n3457 );
    not g36278 ( n32614 , n9138 );
    xnor g36279 ( n31350 , n6147 , n18149 );
    or g36280 ( n20794 , n24183 , n37181 );
    xnor g36281 ( n28388 , n36778 , n19940 );
    not g36282 ( n7127 , n3490 );
    not g36283 ( n20699 , n25700 );
    not g36284 ( n16623 , n22009 );
    xnor g36285 ( n39146 , n15061 , n10744 );
    or g36286 ( n28054 , n10260 , n30325 );
    nor g36287 ( n28448 , n42196 , n36554 );
    or g36288 ( n36821 , n9327 , n15900 );
    not g36289 ( n13540 , n12418 );
    not g36290 ( n30739 , n11882 );
    or g36291 ( n36398 , n9145 , n40480 );
    not g36292 ( n33854 , n17107 );
    not g36293 ( n1356 , n26686 );
    and g36294 ( n18282 , n28548 , n36596 );
    xnor g36295 ( n19862 , n39300 , n5605 );
    xnor g36296 ( n41745 , n784 , n26585 );
    or g36297 ( n26721 , n2905 , n34793 );
    nor g36298 ( n12961 , n4079 , n20238 );
    or g36299 ( n5095 , n14707 , n26953 );
    xnor g36300 ( n25094 , n1338 , n34567 );
    or g36301 ( n5638 , n30226 , n20391 );
    or g36302 ( n25629 , n21631 , n6159 );
    nor g36303 ( n37583 , n110 , n26662 );
    or g36304 ( n4439 , n2713 , n36880 );
    or g36305 ( n38567 , n34565 , n2897 );
    or g36306 ( n19941 , n36770 , n27278 );
    or g36307 ( n32250 , n26933 , n13733 );
    not g36308 ( n40374 , n2235 );
    nor g36309 ( n16744 , n23962 , n26240 );
    nor g36310 ( n29266 , n17276 , n19624 );
    or g36311 ( n42643 , n6550 , n6358 );
    xnor g36312 ( n3299 , n21534 , n23756 );
    and g36313 ( n24607 , n36828 , n18765 );
    or g36314 ( n20105 , n37075 , n5526 );
    or g36315 ( n40452 , n34565 , n8381 );
    and g36316 ( n23453 , n2049 , n5501 );
    and g36317 ( n11183 , n18909 , n15099 );
    nor g36318 ( n3318 , n18520 , n30786 );
    or g36319 ( n17113 , n39489 , n17078 );
    nor g36320 ( n32352 , n18051 , n40669 );
    xnor g36321 ( n5086 , n34875 , n12575 );
    xnor g36322 ( n39165 , n3456 , n36138 );
    or g36323 ( n23078 , n20900 , n11743 );
    or g36324 ( n11635 , n30358 , n39753 );
    or g36325 ( n195 , n5896 , n29619 );
    or g36326 ( n19201 , n37790 , n38007 );
    nor g36327 ( n23151 , n15429 , n25540 );
    and g36328 ( n24786 , n33214 , n12412 );
    xnor g36329 ( n32450 , n19700 , n31603 );
    xor g36330 ( n33436 , n11118 , n16865 );
    or g36331 ( n29356 , n38110 , n34578 );
    not g36332 ( n35355 , n22694 );
    or g36333 ( n39554 , n27540 , n36795 );
    xnor g36334 ( n4001 , n36998 , n26675 );
    xnor g36335 ( n30037 , n35823 , n33981 );
    nor g36336 ( n16520 , n9880 , n23632 );
    or g36337 ( n39826 , n33464 , n36395 );
    xnor g36338 ( n19461 , n9825 , n41534 );
    or g36339 ( n14971 , n42565 , n2997 );
    or g36340 ( n8436 , n38023 , n32829 );
    or g36341 ( n42498 , n42447 , n34574 );
    and g36342 ( n28991 , n9442 , n42622 );
    or g36343 ( n18022 , n26455 , n31580 );
    and g36344 ( n32327 , n35753 , n7578 );
    not g36345 ( n20420 , n26034 );
    or g36346 ( n14164 , n42100 , n12153 );
    nor g36347 ( n38232 , n9355 , n33516 );
    or g36348 ( n13836 , n5882 , n8710 );
    not g36349 ( n11559 , n8465 );
    not g36350 ( n36702 , n24612 );
    and g36351 ( n13212 , n6107 , n24192 );
    and g36352 ( n40746 , n36254 , n1600 );
    not g36353 ( n40024 , n11469 );
    nor g36354 ( n21252 , n41818 , n37442 );
    or g36355 ( n31627 , n25754 , n27385 );
    nor g36356 ( n20443 , n4345 , n21857 );
    and g36357 ( n16008 , n38010 , n28927 );
    nor g36358 ( n12920 , n7796 , n28446 );
    and g36359 ( n22344 , n29959 , n21717 );
    nor g36360 ( n26728 , n21816 , n34024 );
    nor g36361 ( n25735 , n35005 , n41914 );
    and g36362 ( n23476 , n27338 , n36136 );
    xnor g36363 ( n15001 , n40391 , n16325 );
    xnor g36364 ( n15125 , n34112 , n21540 );
    nor g36365 ( n29813 , n8054 , n12755 );
    or g36366 ( n29785 , n41827 , n20633 );
    or g36367 ( n8252 , n24053 , n18522 );
    not g36368 ( n28143 , n26673 );
    xnor g36369 ( n4967 , n16693 , n19397 );
    and g36370 ( n38150 , n9869 , n23117 );
    and g36371 ( n11961 , n20948 , n29654 );
    nor g36372 ( n153 , n19221 , n22721 );
    or g36373 ( n33753 , n121 , n32680 );
    and g36374 ( n11111 , n17151 , n39290 );
    or g36375 ( n42285 , n41730 , n42630 );
    and g36376 ( n25831 , n26323 , n34282 );
    or g36377 ( n34242 , n16532 , n21691 );
    or g36378 ( n38796 , n11498 , n28165 );
    nor g36379 ( n27897 , n11277 , n42807 );
    nor g36380 ( n19193 , n5953 , n30383 );
    or g36381 ( n6895 , n34292 , n39455 );
    nor g36382 ( n17422 , n11070 , n30588 );
    xnor g36383 ( n11135 , n22771 , n18932 );
    or g36384 ( n6928 , n23860 , n16605 );
    or g36385 ( n3652 , n41699 , n28566 );
    and g36386 ( n17218 , n3673 , n34381 );
    xnor g36387 ( n38089 , n42060 , n11200 );
    or g36388 ( n22938 , n28007 , n42447 );
    or g36389 ( n34303 , n23509 , n12784 );
    or g36390 ( n5446 , n11789 , n19510 );
    xnor g36391 ( n27072 , n6090 , n4610 );
    xnor g36392 ( n27195 , n1599 , n40582 );
    or g36393 ( n30885 , n7861 , n30504 );
    or g36394 ( n15218 , n32799 , n21466 );
    or g36395 ( n19236 , n26154 , n39400 );
    nor g36396 ( n32339 , n32408 , n13122 );
    nor g36397 ( n31595 , n18489 , n8165 );
    nor g36398 ( n33670 , n6106 , n1200 );
    nor g36399 ( n21962 , n27134 , n41468 );
    xnor g36400 ( n38346 , n37738 , n1851 );
    or g36401 ( n21374 , n38879 , n25021 );
    xnor g36402 ( n20502 , n105 , n14848 );
    xnor g36403 ( n33258 , n6969 , n4675 );
    and g36404 ( n39216 , n75 , n31984 );
    or g36405 ( n35464 , n35049 , n7616 );
    xnor g36406 ( n34348 , n5144 , n17388 );
    or g36407 ( n13618 , n17451 , n16440 );
    or g36408 ( n38072 , n40673 , n26224 );
    nor g36409 ( n7083 , n14506 , n38409 );
    not g36410 ( n16702 , n37051 );
    or g36411 ( n42182 , n39771 , n33530 );
    not g36412 ( n5917 , n33558 );
    and g36413 ( n11667 , n27230 , n40242 );
    not g36414 ( n29930 , n18800 );
    xnor g36415 ( n21154 , n18335 , n6643 );
    or g36416 ( n20661 , n34996 , n41337 );
    and g36417 ( n37752 , n34237 , n33968 );
    nor g36418 ( n10331 , n36667 , n1211 );
    and g36419 ( n17370 , n12960 , n6274 );
    and g36420 ( n21563 , n9560 , n41316 );
    nor g36421 ( n32656 , n32277 , n38633 );
    not g36422 ( n18102 , n20513 );
    xnor g36423 ( n4649 , n35727 , n2077 );
    not g36424 ( n5197 , n40725 );
    or g36425 ( n13016 , n23118 , n32410 );
    nor g36426 ( n19899 , n785 , n13255 );
    or g36427 ( n34377 , n26098 , n8768 );
    or g36428 ( n33933 , n15282 , n34080 );
    or g36429 ( n37093 , n4492 , n14707 );
    and g36430 ( n15011 , n18409 , n33404 );
    and g36431 ( n29982 , n3204 , n31171 );
    not g36432 ( n28654 , n26855 );
    or g36433 ( n23394 , n7408 , n35269 );
    or g36434 ( n21859 , n10505 , n18589 );
    and g36435 ( n9789 , n25691 , n40403 );
    and g36436 ( n30455 , n4389 , n24253 );
    nor g36437 ( n8293 , n38251 , n32149 );
    nor g36438 ( n2834 , n34698 , n32771 );
    not g36439 ( n21448 , n28051 );
    not g36440 ( n23199 , n37822 );
    not g36441 ( n17739 , n15647 );
    not g36442 ( n9116 , n9174 );
    or g36443 ( n20725 , n12399 , n29384 );
    or g36444 ( n38180 , n16150 , n10161 );
    or g36445 ( n25075 , n25637 , n37623 );
    xnor g36446 ( n6866 , n4284 , n12211 );
    or g36447 ( n11826 , n28535 , n5728 );
    not g36448 ( n13885 , n9432 );
    not g36449 ( n39194 , n19685 );
    xnor g36450 ( n21475 , n38911 , n35618 );
    and g36451 ( n37645 , n2038 , n18876 );
    or g36452 ( n24102 , n11188 , n16137 );
    or g36453 ( n14802 , n23475 , n1416 );
    or g36454 ( n20635 , n24806 , n33798 );
    nor g36455 ( n10027 , n32422 , n16175 );
    or g36456 ( n19075 , n35815 , n24114 );
    and g36457 ( n18884 , n22337 , n35622 );
    xnor g36458 ( n27064 , n10527 , n27624 );
    nor g36459 ( n7931 , n18953 , n25458 );
    or g36460 ( n7697 , n283 , n28882 );
    or g36461 ( n1894 , n33981 , n6946 );
    or g36462 ( n24150 , n40348 , n41860 );
    or g36463 ( n40632 , n15364 , n20409 );
    xnor g36464 ( n3227 , n18942 , n23382 );
    and g36465 ( n40885 , n14403 , n22486 );
    nor g36466 ( n29251 , n36302 , n31938 );
    nor g36467 ( n27678 , n12543 , n1858 );
    or g36468 ( n10052 , n21014 , n14089 );
    and g36469 ( n35207 , n27704 , n16637 );
    nor g36470 ( n42911 , n29052 , n33557 );
    or g36471 ( n11665 , n3454 , n6991 );
    or g36472 ( n27139 , n14707 , n36459 );
    and g36473 ( n32587 , n41199 , n14165 );
    or g36474 ( n32192 , n35763 , n27931 );
    xnor g36475 ( n33875 , n16693 , n3845 );
    not g36476 ( n446 , n26287 );
    or g36477 ( n15019 , n8023 , n10053 );
    xnor g36478 ( n14720 , n18192 , n16892 );
    nor g36479 ( n25266 , n6994 , n29428 );
    and g36480 ( n10816 , n28381 , n6099 );
    or g36481 ( n17962 , n32245 , n42422 );
    or g36482 ( n21163 , n15359 , n24108 );
    nor g36483 ( n31464 , n26722 , n717 );
    not g36484 ( n20632 , n29048 );
    and g36485 ( n9719 , n10084 , n20358 );
    xnor g36486 ( n7898 , n35377 , n16955 );
    nor g36487 ( n7842 , n6867 , n14152 );
    not g36488 ( n13643 , n28531 );
    and g36489 ( n24475 , n11419 , n23645 );
    or g36490 ( n35729 , n25003 , n32892 );
    xnor g36491 ( n28567 , n11383 , n24653 );
    xnor g36492 ( n9886 , n32351 , n17829 );
    or g36493 ( n11912 , n18169 , n639 );
    or g36494 ( n7581 , n28079 , n36393 );
    or g36495 ( n28866 , n42143 , n39646 );
    xnor g36496 ( n15400 , n29956 , n26324 );
    or g36497 ( n21331 , n10674 , n17407 );
    xnor g36498 ( n24404 , n34875 , n37567 );
    or g36499 ( n15502 , n40837 , n37517 );
    not g36500 ( n4948 , n22904 );
    and g36501 ( n42021 , n30933 , n27 );
    not g36502 ( n33561 , n399 );
    or g36503 ( n24558 , n9961 , n23771 );
    and g36504 ( n3885 , n34811 , n5162 );
    and g36505 ( n35374 , n21897 , n20739 );
    or g36506 ( n7720 , n20748 , n41079 );
    or g36507 ( n40619 , n1497 , n26888 );
    not g36508 ( n14143 , n25660 );
    not g36509 ( n33264 , n24954 );
    or g36510 ( n21120 , n39327 , n14450 );
    or g36511 ( n3228 , n7493 , n20446 );
    or g36512 ( n17905 , n17005 , n8220 );
    xnor g36513 ( n19319 , n39722 , n29627 );
    not g36514 ( n32356 , n31701 );
    and g36515 ( n7681 , n26540 , n12437 );
    or g36516 ( n3496 , n11813 , n23545 );
    or g36517 ( n29420 , n22869 , n20090 );
    not g36518 ( n38818 , n36654 );
    not g36519 ( n24371 , n24221 );
    or g36520 ( n17096 , n30864 , n16955 );
    xnor g36521 ( n30380 , n36451 , n21062 );
    or g36522 ( n1849 , n30255 , n36213 );
    xnor g36523 ( n14843 , n330 , n27269 );
    or g36524 ( n1394 , n17909 , n3622 );
    not g36525 ( n8949 , n13138 );
    or g36526 ( n19948 , n30126 , n25768 );
    not g36527 ( n19867 , n6623 );
    and g36528 ( n37213 , n30203 , n31063 );
    not g36529 ( n8777 , n38106 );
    xnor g36530 ( n28357 , n16418 , n33964 );
    and g36531 ( n17390 , n22768 , n42318 );
    or g36532 ( n9828 , n12520 , n22847 );
    or g36533 ( n37316 , n35271 , n2269 );
    not g36534 ( n5175 , n18119 );
    or g36535 ( n18194 , n20295 , n12317 );
    or g36536 ( n37039 , n32277 , n12972 );
    and g36537 ( n13773 , n29831 , n9356 );
    or g36538 ( n5339 , n28426 , n32579 );
    or g36539 ( n31574 , n2276 , n26438 );
    not g36540 ( n36894 , n2221 );
    nor g36541 ( n33322 , n26067 , n28810 );
    or g36542 ( n424 , n3212 , n34360 );
    not g36543 ( n13811 , n1584 );
    or g36544 ( n41894 , n2710 , n38840 );
    nor g36545 ( n34516 , n22027 , n13351 );
    and g36546 ( n36831 , n4055 , n34219 );
    or g36547 ( n28792 , n22450 , n8037 );
    or g36548 ( n17251 , n19400 , n182 );
    not g36549 ( n29120 , n25893 );
    xnor g36550 ( n24798 , n24093 , n27252 );
    not g36551 ( n7574 , n14008 );
    or g36552 ( n12643 , n20 , n10332 );
    not g36553 ( n29299 , n31157 );
    xnor g36554 ( n21978 , n12876 , n28235 );
    or g36555 ( n18949 , n7196 , n18313 );
    or g36556 ( n25189 , n16601 , n12463 );
    or g36557 ( n11701 , n20940 , n1631 );
    or g36558 ( n14069 , n39495 , n25528 );
    or g36559 ( n11792 , n27276 , n31238 );
    not g36560 ( n35156 , n20132 );
    and g36561 ( n18889 , n2014 , n38950 );
    or g36562 ( n32880 , n36659 , n41007 );
    or g36563 ( n31079 , n39538 , n1386 );
    not g36564 ( n25884 , n1287 );
    or g36565 ( n4728 , n27372 , n39481 );
    xnor g36566 ( n179 , n24163 , n21446 );
    or g36567 ( n25363 , n29882 , n42220 );
    or g36568 ( n1542 , n1666 , n22633 );
    not g36569 ( n34625 , n6432 );
    or g36570 ( n20645 , n23908 , n18870 );
    and g36571 ( n26005 , n19324 , n660 );
    not g36572 ( n13106 , n42915 );
    or g36573 ( n37459 , n10674 , n32040 );
    or g36574 ( n8943 , n26927 , n11586 );
    or g36575 ( n28232 , n19808 , n30404 );
    and g36576 ( n9405 , n25068 , n14121 );
    or g36577 ( n860 , n28491 , n23515 );
    nor g36578 ( n30301 , n8827 , n26206 );
    and g36579 ( n5142 , n42528 , n15197 );
    or g36580 ( n22663 , n28898 , n1013 );
    not g36581 ( n10012 , n6542 );
    or g36582 ( n34948 , n12383 , n26873 );
    xnor g36583 ( n1098 , n4392 , n10288 );
    or g36584 ( n11626 , n7751 , n4369 );
    and g36585 ( n18553 , n15924 , n1237 );
    xnor g36586 ( n13648 , n32132 , n33432 );
    xnor g36587 ( n35126 , n6625 , n26953 );
    xnor g36588 ( n16846 , n6242 , n14885 );
    not g36589 ( n21078 , n30988 );
    xnor g36590 ( n24399 , n13624 , n41154 );
    or g36591 ( n12569 , n5207 , n12319 );
    not g36592 ( n26647 , n16107 );
    not g36593 ( n32345 , n1831 );
    or g36594 ( n35884 , n41439 , n15883 );
    or g36595 ( n1040 , n35127 , n19842 );
    or g36596 ( n5336 , n40237 , n42316 );
    or g36597 ( n23251 , n28634 , n24369 );
    or g36598 ( n42330 , n17744 , n7417 );
    and g36599 ( n13951 , n11633 , n41538 );
    and g36600 ( n16734 , n25294 , n34026 );
    xnor g36601 ( n18561 , n10024 , n28935 );
    and g36602 ( n42908 , n7078 , n19301 );
    or g36603 ( n16337 , n22167 , n36752 );
    and g36604 ( n1190 , n24287 , n4300 );
    and g36605 ( n1576 , n25385 , n2551 );
    nor g36606 ( n42304 , n31273 , n38716 );
    nor g36607 ( n26639 , n25775 , n24662 );
    or g36608 ( n28282 , n20509 , n20924 );
    or g36609 ( n29786 , n3089 , n6999 );
    nor g36610 ( n37348 , n42553 , n36038 );
    or g36611 ( n33351 , n38074 , n34571 );
    not g36612 ( n29743 , n24102 );
    nor g36613 ( n2108 , n2851 , n24239 );
    or g36614 ( n31815 , n10395 , n16141 );
    or g36615 ( n16184 , n4430 , n13486 );
    or g36616 ( n19157 , n22730 , n27365 );
    and g36617 ( n15659 , n15429 , n19072 );
    or g36618 ( n14404 , n41013 , n743 );
    xnor g36619 ( n30809 , n2956 , n23314 );
    nor g36620 ( n7408 , n12353 , n34178 );
    or g36621 ( n544 , n41328 , n29559 );
    not g36622 ( n24264 , n7975 );
    xnor g36623 ( n10688 , n42360 , n38495 );
    and g36624 ( n28909 , n33181 , n24941 );
    or g36625 ( n24242 , n24062 , n27062 );
    or g36626 ( n36692 , n20387 , n18553 );
    or g36627 ( n368 , n2140 , n9508 );
    not g36628 ( n1636 , n22195 );
    or g36629 ( n38304 , n15752 , n3403 );
    or g36630 ( n16478 , n4431 , n21970 );
    or g36631 ( n23661 , n550 , n22998 );
    or g36632 ( n30922 , n34428 , n29230 );
    or g36633 ( n31463 , n22765 , n867 );
    nor g36634 ( n7593 , n4340 , n16192 );
    xnor g36635 ( n13736 , n31848 , n1296 );
    and g36636 ( n9538 , n29174 , n6535 );
    not g36637 ( n32253 , n20553 );
    and g36638 ( n10274 , n35563 , n1914 );
    or g36639 ( n24964 , n20444 , n24426 );
    and g36640 ( n6916 , n23754 , n27684 );
    xnor g36641 ( n18186 , n38428 , n34565 );
    and g36642 ( n17386 , n22402 , n8351 );
    xnor g36643 ( n30711 , n13245 , n16156 );
    not g36644 ( n4509 , n8389 );
    or g36645 ( n10267 , n32885 , n26992 );
    and g36646 ( n24224 , n6520 , n719 );
    not g36647 ( n28825 , n36552 );
    or g36648 ( n17312 , n30284 , n31618 );
    or g36649 ( n33634 , n2972 , n29197 );
    and g36650 ( n27951 , n18948 , n32979 );
    and g36651 ( n21781 , n22410 , n4613 );
    not g36652 ( n4013 , n6421 );
    not g36653 ( n6770 , n36267 );
    or g36654 ( n22262 , n18628 , n14010 );
    or g36655 ( n32415 , n33685 , n31156 );
    or g36656 ( n40809 , n34722 , n32243 );
    or g36657 ( n36487 , n28074 , n33897 );
    xnor g36658 ( n27664 , n2419 , n474 );
    and g36659 ( n24308 , n26364 , n18643 );
    nor g36660 ( n15655 , n5679 , n19460 );
    or g36661 ( n24448 , n3944 , n10702 );
    xnor g36662 ( n9435 , n27077 , n37413 );
    or g36663 ( n3471 , n38879 , n26638 );
    and g36664 ( n18841 , n38328 , n31304 );
    nor g36665 ( n34328 , n13863 , n31745 );
    or g36666 ( n4320 , n41319 , n7559 );
    or g36667 ( n10659 , n6082 , n20383 );
    xnor g36668 ( n3296 , n30271 , n18166 );
    nor g36669 ( n28513 , n20173 , n18532 );
    or g36670 ( n27890 , n8288 , n36848 );
    nor g36671 ( n1892 , n29759 , n27778 );
    or g36672 ( n32236 , n9057 , n28816 );
    or g36673 ( n25124 , n17870 , n30597 );
    nor g36674 ( n4400 , n37017 , n35373 );
    and g36675 ( n20646 , n36677 , n31612 );
    and g36676 ( n6946 , n16944 , n41660 );
    and g36677 ( n7337 , n34690 , n9251 );
    xnor g36678 ( n15812 , n25041 , n6669 );
    or g36679 ( n23713 , n16912 , n41007 );
    or g36680 ( n30270 , n5910 , n26931 );
    or g36681 ( n1695 , n37617 , n8784 );
    and g36682 ( n41108 , n4800 , n40649 );
    or g36683 ( n13315 , n6410 , n4394 );
    or g36684 ( n27182 , n10310 , n2650 );
    or g36685 ( n24950 , n2965 , n7981 );
    or g36686 ( n10210 , n6756 , n38926 );
    nor g36687 ( n30676 , n2199 , n13277 );
    or g36688 ( n3529 , n5292 , n24593 );
    or g36689 ( n40069 , n28200 , n9040 );
    not g36690 ( n37829 , n4109 );
    not g36691 ( n4822 , n11524 );
    and g36692 ( n26183 , n36047 , n11342 );
    and g36693 ( n6845 , n12364 , n24237 );
    or g36694 ( n40862 , n24917 , n23355 );
    not g36695 ( n7457 , n7972 );
    xnor g36696 ( n10127 , n42064 , n33900 );
    or g36697 ( n26257 , n2881 , n41007 );
    or g36698 ( n1350 , n28780 , n10996 );
    not g36699 ( n40253 , n25642 );
    and g36700 ( n21886 , n30856 , n23909 );
    and g36701 ( n11859 , n32279 , n8834 );
    or g36702 ( n38644 , n13524 , n37247 );
    or g36703 ( n24756 , n12262 , n10900 );
    or g36704 ( n16641 , n25543 , n2599 );
    not g36705 ( n18665 , n12276 );
    and g36706 ( n1369 , n4818 , n1391 );
    or g36707 ( n33214 , n18199 , n32079 );
    not g36708 ( n41565 , n40977 );
    or g36709 ( n2520 , n31471 , n26204 );
    or g36710 ( n26521 , n1049 , n10391 );
    or g36711 ( n42287 , n26197 , n35216 );
    or g36712 ( n1537 , n2204 , n11967 );
    or g36713 ( n35900 , n35460 , n27087 );
    and g36714 ( n25146 , n34969 , n42182 );
    not g36715 ( n15342 , n1793 );
    and g36716 ( n26838 , n18171 , n41229 );
    xnor g36717 ( n14026 , n7836 , n5075 );
    or g36718 ( n33603 , n31201 , n38944 );
    and g36719 ( n3595 , n34660 , n29881 );
    xnor g36720 ( n9695 , n5144 , n852 );
    and g36721 ( n36288 , n24744 , n20019 );
    nor g36722 ( n15350 , n18813 , n15420 );
    or g36723 ( n12342 , n11367 , n25572 );
    and g36724 ( n31379 , n20823 , n5316 );
    and g36725 ( n2448 , n14109 , n39099 );
    or g36726 ( n18019 , n12051 , n15048 );
    and g36727 ( n22353 , n21824 , n16869 );
    or g36728 ( n32199 , n20804 , n16615 );
    xnor g36729 ( n20124 , n13181 , n6588 );
    and g36730 ( n29156 , n31774 , n27997 );
    or g36731 ( n19257 , n8608 , n37734 );
    and g36732 ( n12904 , n18488 , n19974 );
    not g36733 ( n39289 , n5097 );
    and g36734 ( n35013 , n4095 , n18617 );
    nor g36735 ( n30932 , n24191 , n7555 );
    xnor g36736 ( n8556 , n37932 , n21058 );
    or g36737 ( n31358 , n33338 , n29744 );
    nor g36738 ( n37796 , n4448 , n5089 );
    and g36739 ( n28349 , n17698 , n12195 );
    nor g36740 ( n1959 , n12156 , n7747 );
    nor g36741 ( n21396 , n38157 , n21378 );
    not g36742 ( n42247 , n34427 );
    or g36743 ( n24169 , n19782 , n32909 );
    or g36744 ( n32720 , n31886 , n23321 );
    not g36745 ( n11327 , n13615 );
    xnor g36746 ( n4729 , n18506 , n6416 );
    or g36747 ( n28022 , n15152 , n26211 );
    not g36748 ( n41654 , n4719 );
    not g36749 ( n41728 , n34151 );
    not g36750 ( n12193 , n9293 );
    or g36751 ( n30973 , n32231 , n35756 );
    and g36752 ( n41962 , n25284 , n41686 );
    and g36753 ( n32693 , n41477 , n16157 );
    or g36754 ( n2797 , n42375 , n30435 );
    and g36755 ( n7473 , n23820 , n15114 );
    or g36756 ( n9994 , n26681 , n33099 );
    or g36757 ( n24667 , n19753 , n3132 );
    or g36758 ( n4070 , n6640 , n12826 );
    or g36759 ( n24237 , n13190 , n31687 );
    and g36760 ( n20497 , n42729 , n38397 );
    nor g36761 ( n6244 , n37685 , n8355 );
    nor g36762 ( n5020 , n6503 , n1240 );
    nor g36763 ( n28758 , n33617 , n10531 );
    or g36764 ( n32791 , n19488 , n2095 );
    or g36765 ( n17590 , n17898 , n36672 );
    not g36766 ( n24000 , n26871 );
    or g36767 ( n29746 , n36335 , n38191 );
    not g36768 ( n41558 , n10549 );
    nor g36769 ( n20422 , n11668 , n11715 );
    or g36770 ( n2805 , n22530 , n29643 );
    nor g36771 ( n25110 , n34292 , n23035 );
    nor g36772 ( n15768 , n14298 , n36401 );
    xnor g36773 ( n7461 , n5144 , n39972 );
    or g36774 ( n34357 , n38493 , n23701 );
    nor g36775 ( n22595 , n4334 , n1883 );
    not g36776 ( n6088 , n8477 );
    or g36777 ( n20043 , n22021 , n6024 );
    or g36778 ( n33092 , n6247 , n26839 );
    nor g36779 ( n13766 , n20222 , n18251 );
    nor g36780 ( n6484 , n15194 , n3461 );
    xnor g36781 ( n12673 , n35035 , n22815 );
    or g36782 ( n8226 , n15681 , n7957 );
    xnor g36783 ( n19181 , n10535 , n28535 );
    not g36784 ( n5982 , n26063 );
    nor g36785 ( n7034 , n25588 , n6570 );
    not g36786 ( n25477 , n41631 );
    or g36787 ( n57 , n11431 , n40736 );
    not g36788 ( n17438 , n28545 );
    nor g36789 ( n12040 , n23431 , n15294 );
    not g36790 ( n16106 , n34931 );
    or g36791 ( n20563 , n30754 , n28847 );
    not g36792 ( n27891 , n14046 );
    not g36793 ( n6991 , n38490 );
    or g36794 ( n8822 , n25711 , n39311 );
    nor g36795 ( n2299 , n9607 , n2671 );
    nor g36796 ( n38227 , n37165 , n19063 );
    and g36797 ( n13625 , n42819 , n18682 );
    or g36798 ( n6856 , n17513 , n28727 );
    xnor g36799 ( n28212 , n10601 , n6772 );
    xnor g36800 ( n20536 , n16693 , n11208 );
    or g36801 ( n12760 , n32724 , n27464 );
    and g36802 ( n36342 , n3144 , n40007 );
    xnor g36803 ( n21145 , n7407 , n41534 );
    nor g36804 ( n25896 , n6330 , n31620 );
    or g36805 ( n25666 , n28468 , n41980 );
    not g36806 ( n16636 , n23353 );
    not g36807 ( n7853 , n6698 );
    not g36808 ( n4671 , n22230 );
    or g36809 ( n32870 , n17744 , n24162 );
    not g36810 ( n17435 , n40585 );
    or g36811 ( n10436 , n28566 , n41197 );
    nor g36812 ( n34916 , n38879 , n10851 );
    and g36813 ( n24828 , n16391 , n10387 );
    and g36814 ( n1113 , n36705 , n17866 );
    and g36815 ( n28309 , n34245 , n25162 );
    and g36816 ( n28539 , n3233 , n29007 );
    and g36817 ( n39576 , n20166 , n35327 );
    or g36818 ( n12259 , n36296 , n40741 );
    or g36819 ( n21684 , n29937 , n8170 );
    or g36820 ( n33266 , n21478 , n17656 );
    and g36821 ( n13528 , n24884 , n24604 );
    or g36822 ( n2969 , n31542 , n40714 );
    or g36823 ( n9685 , n20268 , n9487 );
    not g36824 ( n15979 , n36610 );
    and g36825 ( n16439 , n29506 , n10782 );
    or g36826 ( n18661 , n35483 , n37862 );
    or g36827 ( n29666 , n30030 , n30786 );
    or g36828 ( n12398 , n5217 , n16301 );
    xnor g36829 ( n15783 , n4467 , n10296 );
    nor g36830 ( n14343 , n15372 , n19992 );
    and g36831 ( n11968 , n25759 , n38644 );
    not g36832 ( n34774 , n7382 );
    and g36833 ( n8042 , n17701 , n13126 );
    not g36834 ( n37169 , n1985 );
    or g36835 ( n31395 , n4492 , n38102 );
    or g36836 ( n16169 , n35915 , n2615 );
    or g36837 ( n19943 , n13419 , n32791 );
    or g36838 ( n1739 , n40961 , n16996 );
    xnor g36839 ( n18600 , n20958 , n10087 );
    or g36840 ( n23508 , n41923 , n31664 );
    xnor g36841 ( n10065 , n19268 , n31661 );
    or g36842 ( n32806 , n14271 , n21049 );
    or g36843 ( n362 , n2226 , n5860 );
    and g36844 ( n7742 , n31683 , n21081 );
    and g36845 ( n18779 , n11121 , n37710 );
    or g36846 ( n28862 , n23446 , n27738 );
    nor g36847 ( n14291 , n3502 , n37567 );
    nor g36848 ( n11331 , n23026 , n33048 );
    or g36849 ( n14083 , n18622 , n41072 );
    nor g36850 ( n6050 , n14226 , n1296 );
    not g36851 ( n19166 , n22514 );
    and g36852 ( n3598 , n13359 , n35973 );
    and g36853 ( n25090 , n20135 , n19461 );
    xnor g36854 ( n18588 , n37083 , n30812 );
    and g36855 ( n32233 , n29304 , n29805 );
    or g36856 ( n35397 , n20932 , n16351 );
    or g36857 ( n19648 , n5445 , n10745 );
    and g36858 ( n30152 , n27361 , n3123 );
    not g36859 ( n8220 , n38262 );
    not g36860 ( n10714 , n1832 );
    nor g36861 ( n24395 , n8494 , n17460 );
    or g36862 ( n38291 , n11756 , n11871 );
    and g36863 ( n4533 , n18229 , n31983 );
    and g36864 ( n14617 , n37151 , n17315 );
    xnor g36865 ( n26949 , n38749 , n30113 );
    and g36866 ( n22709 , n10927 , n24295 );
    not g36867 ( n19337 , n36392 );
    nor g36868 ( n24797 , n23089 , n24335 );
    or g36869 ( n20471 , n30677 , n30119 );
    or g36870 ( n22560 , n9329 , n35562 );
    xnor g36871 ( n1411 , n33570 , n6187 );
    xnor g36872 ( n20800 , n12146 , n32151 );
    nor g36873 ( n36533 , n24950 , n14538 );
    or g36874 ( n29798 , n23531 , n3583 );
    or g36875 ( n8367 , n6247 , n17325 );
    not g36876 ( n32019 , n29030 );
    or g36877 ( n36840 , n22841 , n14590 );
    or g36878 ( n37479 , n15900 , n5506 );
    xnor g36879 ( n13721 , n39412 , n29020 );
    and g36880 ( n41887 , n2433 , n22865 );
    or g36881 ( n20303 , n22172 , n38199 );
    and g36882 ( n14726 , n23892 , n10538 );
    or g36883 ( n34271 , n17984 , n25833 );
    and g36884 ( n64 , n41241 , n21920 );
    or g36885 ( n5963 , n2370 , n26740 );
    or g36886 ( n19474 , n3333 , n28204 );
    or g36887 ( n8296 , n8004 , n20907 );
    and g36888 ( n39502 , n19575 , n1628 );
    xnor g36889 ( n14243 , n7922 , n40195 );
    or g36890 ( n21386 , n18866 , n37030 );
    and g36891 ( n28379 , n15363 , n7147 );
    nor g36892 ( n6618 , n10806 , n9896 );
    xnor g36893 ( n39436 , n6774 , n32348 );
    or g36894 ( n16448 , n24454 , n20659 );
    or g36895 ( n34032 , n37233 , n31249 );
    nor g36896 ( n22423 , n13474 , n17747 );
    not g36897 ( n18473 , n19735 );
    or g36898 ( n1868 , n10192 , n4742 );
    nor g36899 ( n20440 , n7130 , n8604 );
    nor g36900 ( n13737 , n10277 , n3339 );
    or g36901 ( n12268 , n23522 , n28239 );
    and g36902 ( n31120 , n21830 , n39554 );
    or g36903 ( n30537 , n21393 , n18473 );
    or g36904 ( n25565 , n40570 , n42101 );
    not g36905 ( n42898 , n29475 );
    or g36906 ( n22114 , n22724 , n18104 );
    or g36907 ( n29954 , n13078 , n26426 );
    nor g36908 ( n16765 , n5964 , n519 );
    or g36909 ( n29329 , n21487 , n37633 );
    or g36910 ( n15155 , n8847 , n15907 );
    xnor g36911 ( n37126 , n12024 , n12925 );
    or g36912 ( n12276 , n28223 , n9881 );
    or g36913 ( n721 , n4492 , n40879 );
    and g36914 ( n32878 , n33832 , n29285 );
    xnor g36915 ( n40726 , n32470 , n34632 );
    not g36916 ( n26933 , n4404 );
    and g36917 ( n21846 , n28840 , n14685 );
    not g36918 ( n15693 , n19119 );
    or g36919 ( n28945 , n6114 , n28520 );
    and g36920 ( n7544 , n23730 , n22113 );
    xnor g36921 ( n41001 , n34090 , n29757 );
    xnor g36922 ( n12763 , n898 , n25446 );
    nor g36923 ( n11529 , n39449 , n7356 );
    nor g36924 ( n10518 , n6106 , n20626 );
    xnor g36925 ( n29355 , n20056 , n20319 );
    not g36926 ( n10224 , n10113 );
    or g36927 ( n24139 , n42870 , n11105 );
    and g36928 ( n22983 , n15247 , n9034 );
    or g36929 ( n14409 , n38143 , n29299 );
    or g36930 ( n17748 , n39367 , n35403 );
    or g36931 ( n20084 , n15681 , n22853 );
    not g36932 ( n21654 , n35394 );
    not g36933 ( n18546 , n29461 );
    or g36934 ( n20965 , n40093 , n21938 );
    and g36935 ( n9518 , n38965 , n26356 );
    nor g36936 ( n28383 , n27593 , n823 );
    xnor g36937 ( n35611 , n5891 , n36536 );
    or g36938 ( n9052 , n32786 , n3670 );
    not g36939 ( n13009 , n38271 );
    or g36940 ( n2540 , n33675 , n10429 );
    xnor g36941 ( n11972 , n17049 , n37663 );
    or g36942 ( n2618 , n39439 , n15789 );
    or g36943 ( n33098 , n35528 , n14412 );
    or g36944 ( n21744 , n2630 , n38112 );
    not g36945 ( n21141 , n4822 );
    or g36946 ( n12027 , n10121 , n34949 );
    or g36947 ( n7600 , n40623 , n38151 );
    or g36948 ( n18513 , n10048 , n36687 );
    nor g36949 ( n2524 , n26636 , n9175 );
    nor g36950 ( n38600 , n9988 , n32751 );
    and g36951 ( n22615 , n35819 , n34729 );
    xnor g36952 ( n31847 , n708 , n3867 );
    nor g36953 ( n5869 , n19365 , n16210 );
    xnor g36954 ( n38243 , n18678 , n30028 );
    or g36955 ( n16935 , n20684 , n13498 );
    and g36956 ( n39753 , n40360 , n9606 );
    nor g36957 ( n34755 , n1507 , n4853 );
    or g36958 ( n2405 , n23449 , n27783 );
    or g36959 ( n36338 , n36378 , n8256 );
    or g36960 ( n9109 , n6558 , n31420 );
    nor g36961 ( n14874 , n30465 , n1962 );
    nor g36962 ( n33998 , n1356 , n2957 );
    or g36963 ( n32809 , n12173 , n2729 );
    or g36964 ( n31422 , n15187 , n34225 );
    and g36965 ( n36422 , n16055 , n7062 );
    nor g36966 ( n30159 , n20237 , n4794 );
    not g36967 ( n1441 , n34136 );
    and g36968 ( n14378 , n36854 , n24792 );
    or g36969 ( n36192 , n10284 , n2077 );
    or g36970 ( n38929 , n3147 , n34621 );
    not g36971 ( n36092 , n38361 );
    not g36972 ( n4501 , n8182 );
    and g36973 ( n10503 , n31895 , n33156 );
    nor g36974 ( n40283 , n15261 , n40071 );
    and g36975 ( n20895 , n22096 , n26297 );
    or g36976 ( n20809 , n9540 , n1061 );
    or g36977 ( n7672 , n15031 , n19904 );
    and g36978 ( n18101 , n20769 , n26128 );
    or g36979 ( n16070 , n64 , n28758 );
    and g36980 ( n2643 , n10773 , n2808 );
    not g36981 ( n12495 , n169 );
    or g36982 ( n6597 , n13820 , n9067 );
    and g36983 ( n22297 , n4980 , n15270 );
    or g36984 ( n39901 , n17473 , n31091 );
    not g36985 ( n23130 , n10100 );
    and g36986 ( n25434 , n3478 , n7494 );
    and g36987 ( n27817 , n28602 , n16480 );
    nor g36988 ( n1240 , n19862 , n26352 );
    not g36989 ( n26740 , n40686 );
    or g36990 ( n40977 , n8899 , n38581 );
    xnor g36991 ( n12310 , n41098 , n9713 );
    or g36992 ( n30597 , n21111 , n5471 );
    xnor g36993 ( n3125 , n25619 , n30266 );
    and g36994 ( n39357 , n5627 , n352 );
    or g36995 ( n26463 , n3939 , n41418 );
    and g36996 ( n15809 , n16219 , n15641 );
    or g36997 ( n39049 , n23354 , n40787 );
    nor g36998 ( n31983 , n15272 , n16630 );
    and g36999 ( n11305 , n6076 , n37203 );
    and g37000 ( n7360 , n14516 , n14421 );
    and g37001 ( n30517 , n35241 , n3579 );
    and g37002 ( n14602 , n2003 , n40105 );
    and g37003 ( n41661 , n8382 , n22329 );
    and g37004 ( n24035 , n19990 , n34884 );
    and g37005 ( n14294 , n17731 , n35121 );
    and g37006 ( n27105 , n19654 , n3195 );
    or g37007 ( n22498 , n41056 , n22282 );
    or g37008 ( n2629 , n33755 , n36061 );
    xnor g37009 ( n32625 , n13261 , n18501 );
    and g37010 ( n2601 , n34214 , n13827 );
    or g37011 ( n14183 , n38764 , n37262 );
    not g37012 ( n39954 , n17527 );
    or g37013 ( n22028 , n12794 , n28663 );
    or g37014 ( n9108 , n14481 , n24900 );
    not g37015 ( n7585 , n9519 );
    or g37016 ( n29335 , n6949 , n38191 );
    or g37017 ( n26748 , n35526 , n2813 );
    or g37018 ( n11195 , n35412 , n35758 );
    xnor g37019 ( n34791 , n20974 , n5896 );
    xnor g37020 ( n11366 , n36712 , n31907 );
    not g37021 ( n14531 , n11812 );
    or g37022 ( n19338 , n41382 , n34650 );
    or g37023 ( n9882 , n23319 , n23904 );
    or g37024 ( n5612 , n8896 , n27126 );
    or g37025 ( n29933 , n5658 , n35443 );
    or g37026 ( n20040 , n28041 , n38006 );
    or g37027 ( n1228 , n16216 , n13051 );
    not g37028 ( n8232 , n30438 );
    or g37029 ( n11508 , n31978 , n16001 );
    nor g37030 ( n28385 , n1765 , n30051 );
    xnor g37031 ( n32299 , n21941 , n10473 );
    and g37032 ( n41266 , n2002 , n627 );
    or g37033 ( n37975 , n17112 , n20454 );
    and g37034 ( n1546 , n5990 , n10656 );
    and g37035 ( n8151 , n27197 , n39918 );
    nor g37036 ( n32646 , n34292 , n3845 );
    or g37037 ( n41315 , n10472 , n31625 );
    xnor g37038 ( n26380 , n17158 , n3321 );
    and g37039 ( n24765 , n6324 , n6062 );
    xnor g37040 ( n25981 , n40717 , n18776 );
    xnor g37041 ( n35139 , n31385 , n2941 );
    or g37042 ( n2918 , n165 , n6296 );
    or g37043 ( n9755 , n22023 , n5261 );
    or g37044 ( n2772 , n14749 , n1740 );
    nor g37045 ( n41034 , n6745 , n7251 );
    not g37046 ( n35486 , n29292 );
    and g37047 ( n18063 , n19525 , n34725 );
    and g37048 ( n27464 , n41587 , n3191 );
    nor g37049 ( n10873 , n6525 , n29651 );
    xnor g37050 ( n6864 , n16266 , n4638 );
    or g37051 ( n34763 , n34793 , n3251 );
    or g37052 ( n17354 , n3550 , n41029 );
    not g37053 ( n7753 , n34 );
    and g37054 ( n33743 , n34835 , n2010 );
    nor g37055 ( n38927 , n13683 , n11994 );
    xnor g37056 ( n12281 , n27371 , n8593 );
    or g37057 ( n6482 , n6370 , n29773 );
    and g37058 ( n14664 , n39633 , n19289 );
    and g37059 ( n32877 , n10820 , n24059 );
    or g37060 ( n25386 , n18455 , n3312 );
    and g37061 ( n34998 , n11580 , n17113 );
    or g37062 ( n1603 , n23427 , n34456 );
    and g37063 ( n6078 , n10298 , n23217 );
    or g37064 ( n19287 , n19067 , n29338 );
    not g37065 ( n22220 , n40113 );
    and g37066 ( n6080 , n31689 , n4291 );
    nor g37067 ( n11210 , n10929 , n7019 );
    not g37068 ( n3115 , n12636 );
    and g37069 ( n11834 , n42085 , n39853 );
    or g37070 ( n11543 , n27693 , n15064 );
    and g37071 ( n3570 , n24629 , n14843 );
    not g37072 ( n21689 , n17332 );
    or g37073 ( n28799 , n2451 , n24679 );
    or g37074 ( n19250 , n36213 , n22443 );
    and g37075 ( n34710 , n898 , n36293 );
    xnor g37076 ( n8746 , n352 , n5627 );
    or g37077 ( n40829 , n35026 , n24746 );
    or g37078 ( n31041 , n39186 , n14094 );
    and g37079 ( n19081 , n12712 , n17437 );
    not g37080 ( n36697 , n25207 );
    or g37081 ( n17831 , n38693 , n41845 );
    or g37082 ( n36402 , n3962 , n629 );
    or g37083 ( n14318 , n19540 , n28044 );
    or g37084 ( n38739 , n9566 , n40517 );
    not g37085 ( n38912 , n8051 );
    and g37086 ( n42763 , n32081 , n38457 );
    or g37087 ( n19372 , n4991 , n37779 );
    not g37088 ( n2074 , n13374 );
    nor g37089 ( n4288 , n14217 , n40401 );
    or g37090 ( n22438 , n2878 , n39515 );
    or g37091 ( n20060 , n35251 , n1783 );
    or g37092 ( n3778 , n29477 , n41532 );
    nor g37093 ( n30055 , n37662 , n20218 );
    or g37094 ( n13817 , n22816 , n2242 );
    or g37095 ( n24464 , n30660 , n24371 );
    and g37096 ( n37332 , n28369 , n15380 );
    xnor g37097 ( n30272 , n32470 , n17849 );
    not g37098 ( n34548 , n21007 );
    xnor g37099 ( n5317 , n40130 , n38032 );
    or g37100 ( n42495 , n40785 , n12978 );
    or g37101 ( n16021 , n2255 , n9847 );
    or g37102 ( n3671 , n821 , n29099 );
    and g37103 ( n23973 , n35404 , n100 );
    xnor g37104 ( n25151 , n41013 , n29619 );
    or g37105 ( n36142 , n7973 , n23703 );
    and g37106 ( n2820 , n17372 , n18302 );
    and g37107 ( n8078 , n23200 , n8368 );
    xnor g37108 ( n15683 , n18755 , n21921 );
    or g37109 ( n17192 , n22619 , n16092 );
    or g37110 ( n25493 , n32277 , n33293 );
    or g37111 ( n20885 , n32217 , n14913 );
    or g37112 ( n42629 , n39253 , n19908 );
    or g37113 ( n21485 , n29547 , n425 );
    nor g37114 ( n1220 , n32793 , n11349 );
    nor g37115 ( n14625 , n37071 , n24252 );
    or g37116 ( n1005 , n10153 , n11872 );
    and g37117 ( n21581 , n40183 , n36827 );
    and g37118 ( n2112 , n38990 , n22496 );
    or g37119 ( n42880 , n11222 , n1006 );
    nor g37120 ( n30779 , n39386 , n15870 );
    or g37121 ( n21125 , n8035 , n13888 );
    and g37122 ( n21538 , n31167 , n30021 );
    or g37123 ( n10573 , n31801 , n38343 );
    or g37124 ( n28381 , n32155 , n40323 );
    not g37125 ( n5007 , n24257 );
    and g37126 ( n21205 , n14783 , n31502 );
    or g37127 ( n17242 , n25588 , n3994 );
    or g37128 ( n5176 , n8618 , n9016 );
    xnor g37129 ( n18987 , n2645 , n34080 );
    xnor g37130 ( n34042 , n33838 , n42610 );
    or g37131 ( n24962 , n120 , n4477 );
    or g37132 ( n34340 , n186 , n33232 );
    not g37133 ( n42896 , n37694 );
    or g37134 ( n7259 , n8494 , n23282 );
    xnor g37135 ( n10292 , n7567 , n15661 );
    xnor g37136 ( n28534 , n23510 , n1067 );
    or g37137 ( n38606 , n26442 , n5588 );
    and g37138 ( n40854 , n7741 , n28543 );
    or g37139 ( n6408 , n24613 , n26051 );
    nor g37140 ( n8340 , n36117 , n3642 );
    nor g37141 ( n32173 , n17744 , n315 );
    or g37142 ( n37475 , n18403 , n25831 );
    and g37143 ( n21997 , n8630 , n29628 );
    or g37144 ( n33446 , n405 , n326 );
    and g37145 ( n27536 , n19175 , n3440 );
    or g37146 ( n12267 , n35320 , n17959 );
    not g37147 ( n26032 , n4149 );
    or g37148 ( n26605 , n16996 , n39651 );
    xnor g37149 ( n34015 , n19071 , n32257 );
    or g37150 ( n14661 , n17654 , n20678 );
    and g37151 ( n20066 , n35975 , n21797 );
    or g37152 ( n15945 , n24787 , n17643 );
    or g37153 ( n16009 , n34433 , n2991 );
    and g37154 ( n4159 , n13666 , n15864 );
    and g37155 ( n27645 , n577 , n1019 );
    not g37156 ( n6370 , n14055 );
    and g37157 ( n25429 , n109 , n12911 );
    and g37158 ( n25798 , n23149 , n909 );
    not g37159 ( n562 , n39082 );
    and g37160 ( n2654 , n8303 , n18832 );
    or g37161 ( n11801 , n40035 , n37787 );
    not g37162 ( n31368 , n40301 );
    not g37163 ( n10090 , n42097 );
    nor g37164 ( n4755 , n915 , n19844 );
    or g37165 ( n21472 , n845 , n12153 );
    and g37166 ( n36578 , n15061 , n10744 );
    not g37167 ( n42064 , n2199 );
    nor g37168 ( n8339 , n29296 , n20763 );
    nor g37169 ( n34631 , n39390 , n11956 );
    and g37170 ( n30744 , n28414 , n35200 );
    not g37171 ( n1847 , n5915 );
    not g37172 ( n12397 , n27063 );
    and g37173 ( n9375 , n17964 , n1821 );
    not g37174 ( n17994 , n7655 );
    or g37175 ( n19388 , n27552 , n17875 );
    or g37176 ( n13011 , n42077 , n3203 );
    or g37177 ( n21288 , n41913 , n40516 );
    or g37178 ( n27324 , n31418 , n28141 );
    or g37179 ( n11915 , n24656 , n30814 );
    not g37180 ( n32103 , n27854 );
    or g37181 ( n40640 , n2284 , n21002 );
    and g37182 ( n39299 , n23312 , n29496 );
    or g37183 ( n29901 , n38879 , n36197 );
    or g37184 ( n32156 , n39000 , n23116 );
    and g37185 ( n15789 , n8846 , n39542 );
    or g37186 ( n21450 , n3047 , n33693 );
    or g37187 ( n18505 , n26003 , n29562 );
    not g37188 ( n18835 , n16865 );
    not g37189 ( n29144 , n25163 );
    or g37190 ( n5994 , n8686 , n8353 );
    or g37191 ( n39125 , n13120 , n28745 );
    or g37192 ( n36999 , n23344 , n21819 );
    and g37193 ( n26520 , n25048 , n26181 );
    nor g37194 ( n27164 , n6776 , n39421 );
    not g37195 ( n17371 , n178 );
    or g37196 ( n31974 , n31786 , n31400 );
    or g37197 ( n7284 , n38986 , n946 );
    nor g37198 ( n850 , n10924 , n1392 );
    not g37199 ( n5650 , n20980 );
    and g37200 ( n39057 , n30252 , n38878 );
    and g37201 ( n38919 , n33672 , n28890 );
    nor g37202 ( n38870 , n24948 , n39407 );
    not g37203 ( n28516 , n27893 );
    xnor g37204 ( n17936 , n33050 , n35079 );
    and g37205 ( n942 , n21810 , n20738 );
    not g37206 ( n17148 , n35118 );
    and g37207 ( n4559 , n39198 , n5155 );
    or g37208 ( n20842 , n8109 , n4099 );
    not g37209 ( n32069 , n5675 );
    and g37210 ( n38428 , n469 , n4465 );
    and g37211 ( n12803 , n11274 , n23765 );
    and g37212 ( n16957 , n16349 , n37170 );
    or g37213 ( n28536 , n14407 , n40236 );
    or g37214 ( n33587 , n12105 , n1266 );
    and g37215 ( n37299 , n25895 , n8371 );
    not g37216 ( n28458 , n19580 );
    xnor g37217 ( n879 , n41450 , n4000 );
    or g37218 ( n20240 , n10698 , n3564 );
    or g37219 ( n10243 , n15282 , n1160 );
    or g37220 ( n8263 , n22037 , n29695 );
    and g37221 ( n26764 , n13799 , n38289 );
    or g37222 ( n35116 , n6578 , n14292 );
    not g37223 ( n37247 , n21876 );
    not g37224 ( n19873 , n6475 );
    and g37225 ( n7141 , n13082 , n17490 );
    and g37226 ( n5364 , n15097 , n42262 );
    and g37227 ( n2856 , n39190 , n1854 );
    or g37228 ( n33172 , n30444 , n35549 );
    xnor g37229 ( n27206 , n31099 , n34643 );
    xnor g37230 ( n14919 , n15706 , n42073 );
    nor g37231 ( n2817 , n2118 , n1131 );
    or g37232 ( n727 , n16046 , n3744 );
    nor g37233 ( n19729 , n11380 , n32748 );
    or g37234 ( n33157 , n36308 , n9962 );
    or g37235 ( n22817 , n32873 , n23130 );
    nor g37236 ( n17071 , n15611 , n19975 );
    or g37237 ( n29350 , n12105 , n7765 );
    nor g37238 ( n28484 , n24507 , n36906 );
    or g37239 ( n34261 , n17563 , n39844 );
    not g37240 ( n2012 , n27756 );
    or g37241 ( n416 , n3868 , n21608 );
    not g37242 ( n24336 , n21077 );
    or g37243 ( n8620 , n550 , n9928 );
    not g37244 ( n24592 , n38444 );
    xnor g37245 ( n39615 , n30809 , n29926 );
    or g37246 ( n39181 , n2322 , n14944 );
    nor g37247 ( n32467 , n25588 , n5551 );
    xnor g37248 ( n33751 , n12057 , n3754 );
    nor g37249 ( n15875 , n28879 , n10038 );
    xnor g37250 ( n24947 , n30832 , n22275 );
    and g37251 ( n8115 , n8944 , n23635 );
    and g37252 ( n9813 , n25745 , n12333 );
    or g37253 ( n4125 , n21833 , n41007 );
    not g37254 ( n21666 , n25616 );
    nor g37255 ( n31490 , n4102 , n30672 );
    or g37256 ( n8477 , n28531 , n41903 );
    not g37257 ( n5509 , n31881 );
    or g37258 ( n28877 , n8026 , n40588 );
    xnor g37259 ( n33950 , n32049 , n3168 );
    or g37260 ( n22015 , n269 , n14734 );
    xnor g37261 ( n31239 , n41811 , n35761 );
    or g37262 ( n5706 , n26407 , n27642 );
    xnor g37263 ( n7503 , n30397 , n7623 );
    xnor g37264 ( n30320 , n27762 , n30909 );
    or g37265 ( n27063 , n40228 , n35432 );
    xnor g37266 ( n7029 , n28464 , n4255 );
    nor g37267 ( n42345 , n22176 , n40282 );
    xnor g37268 ( n25692 , n7489 , n30031 );
    not g37269 ( n3455 , n36939 );
    or g37270 ( n21780 , n25456 , n5653 );
    nor g37271 ( n13576 , n39917 , n30982 );
    and g37272 ( n27631 , n10104 , n35353 );
    or g37273 ( n6210 , n27388 , n27926 );
    and g37274 ( n9063 , n5028 , n31054 );
    xnor g37275 ( n399 , n27026 , n7050 );
    or g37276 ( n36353 , n609 , n1922 );
    or g37277 ( n33749 , n18719 , n27686 );
    xnor g37278 ( n2164 , n19599 , n16798 );
    not g37279 ( n1224 , n31665 );
    and g37280 ( n28171 , n23906 , n30367 );
    or g37281 ( n6998 , n40109 , n31809 );
    or g37282 ( n27986 , n36564 , n25233 );
    not g37283 ( n16161 , n32094 );
    and g37284 ( n41862 , n34416 , n27354 );
    not g37285 ( n10704 , n39642 );
    and g37286 ( n39237 , n32907 , n18217 );
    nor g37287 ( n13281 , n28712 , n38455 );
    or g37288 ( n9532 , n42747 , n36848 );
    and g37289 ( n20196 , n30565 , n42562 );
    or g37290 ( n1693 , n9718 , n8823 );
    or g37291 ( n8741 , n16892 , n22872 );
    or g37292 ( n23382 , n157 , n2175 );
    and g37293 ( n25928 , n32966 , n17419 );
    and g37294 ( n3660 , n37165 , n19063 );
    nor g37295 ( n35970 , n34565 , n2470 );
    or g37296 ( n30595 , n42115 , n9799 );
    not g37297 ( n9322 , n28282 );
    and g37298 ( n20207 , n5429 , n20598 );
    or g37299 ( n22720 , n4926 , n31732 );
    not g37300 ( n14475 , n5675 );
    not g37301 ( n23509 , n18915 );
    and g37302 ( n6086 , n24046 , n30063 );
    or g37303 ( n31604 , n34326 , n3314 );
    nor g37304 ( n25372 , n34565 , n13000 );
    or g37305 ( n19697 , n39828 , n12696 );
    or g37306 ( n16080 , n7979 , n31503 );
    or g37307 ( n7025 , n26935 , n13130 );
    or g37308 ( n4763 , n3224 , n16170 );
    not g37309 ( n22184 , n41030 );
    not g37310 ( n2184 , n29799 );
    or g37311 ( n38591 , n27281 , n40228 );
    or g37312 ( n24629 , n2815 , n16031 );
    and g37313 ( n34965 , n24522 , n39172 );
    or g37314 ( n9124 , n39373 , n37263 );
    xnor g37315 ( n6651 , n5001 , n30665 );
    nor g37316 ( n39578 , n24549 , n30086 );
    xnor g37317 ( n15266 , n36506 , n34565 );
    nor g37318 ( n16818 , n38485 , n29241 );
    or g37319 ( n20007 , n2053 , n42534 );
    nor g37320 ( n27690 , n17744 , n32411 );
    or g37321 ( n9445 , n36848 , n6582 );
    xnor g37322 ( n20724 , n22922 , n24347 );
    not g37323 ( n22306 , n32831 );
    or g37324 ( n12362 , n36646 , n15436 );
    or g37325 ( n36982 , n1309 , n19890 );
    not g37326 ( n22345 , n22629 );
    not g37327 ( n5661 , n31364 );
    or g37328 ( n9924 , n28735 , n36239 );
    or g37329 ( n7930 , n17833 , n41657 );
    not g37330 ( n22558 , n37760 );
    nor g37331 ( n25852 , n28276 , n8041 );
    nor g37332 ( n31317 , n30515 , n4917 );
    or g37333 ( n42201 , n4994 , n33556 );
    or g37334 ( n28063 , n7864 , n4160 );
    or g37335 ( n22986 , n28468 , n21783 );
    or g37336 ( n41749 , n9608 , n42364 );
    xnor g37337 ( n11988 , n8656 , n39515 );
    not g37338 ( n41847 , n34922 );
    not g37339 ( n12209 , n16655 );
    or g37340 ( n12908 , n5964 , n7683 );
    and g37341 ( n8581 , n3877 , n4224 );
    and g37342 ( n42462 , n28855 , n40503 );
    or g37343 ( n19710 , n9047 , n37787 );
    or g37344 ( n2690 , n17767 , n1846 );
    or g37345 ( n2691 , n22788 , n33489 );
    or g37346 ( n11954 , n6214 , n4016 );
    or g37347 ( n7382 , n158 , n701 );
    and g37348 ( n40202 , n13296 , n10252 );
    or g37349 ( n8046 , n1060 , n5220 );
    not g37350 ( n11409 , n2661 );
    and g37351 ( n8177 , n14725 , n38272 );
    or g37352 ( n32891 , n9417 , n20194 );
    or g37353 ( n6417 , n31901 , n7823 );
    and g37354 ( n12002 , n32391 , n38445 );
    nor g37355 ( n9721 , n17583 , n11863 );
    and g37356 ( n9217 , n20808 , n10176 );
    nor g37357 ( n7699 , n6132 , n31301 );
    or g37358 ( n24986 , n14481 , n30461 );
    and g37359 ( n32324 , n23571 , n31237 );
    nor g37360 ( n31883 , n14475 , n35337 );
    xnor g37361 ( n6714 , n38378 , n8341 );
    nor g37362 ( n32969 , n27258 , n21318 );
    xnor g37363 ( n35877 , n13444 , n3235 );
    and g37364 ( n5589 , n5598 , n35150 );
    or g37365 ( n7596 , n26599 , n2836 );
    and g37366 ( n28093 , n17155 , n38625 );
    and g37367 ( n31961 , n17781 , n10524 );
    and g37368 ( n31192 , n18657 , n35671 );
    nor g37369 ( n17923 , n18866 , n19664 );
    xnor g37370 ( n41036 , n23197 , n19315 );
    or g37371 ( n3836 , n11270 , n15882 );
    not g37372 ( n41293 , n39742 );
    xnor g37373 ( n15483 , n20272 , n26405 );
    xnor g37374 ( n24862 , n37210 , n42841 );
    xnor g37375 ( n1166 , n27644 , n24024 );
    or g37376 ( n2160 , n5845 , n2597 );
    or g37377 ( n14210 , n10832 , n28447 );
    or g37378 ( n32017 , n2608 , n22708 );
    or g37379 ( n6759 , n31707 , n9134 );
    not g37380 ( n17688 , n19254 );
    and g37381 ( n29546 , n18287 , n26117 );
    nor g37382 ( n2827 , n2214 , n22693 );
    and g37383 ( n40386 , n19586 , n29248 );
    nor g37384 ( n1677 , n30736 , n31561 );
    xnor g37385 ( n921 , n16742 , n19919 );
    or g37386 ( n21776 , n34225 , n28705 );
    not g37387 ( n18401 , n15435 );
    or g37388 ( n22231 , n9692 , n15342 );
    or g37389 ( n3849 , n32133 , n3856 );
    and g37390 ( n38569 , n21835 , n34380 );
    not g37391 ( n21942 , n24810 );
    nor g37392 ( n33804 , n35285 , n29986 );
    or g37393 ( n23615 , n1422 , n12153 );
    nor g37394 ( n4069 , n17792 , n30127 );
    nor g37395 ( n21783 , n39623 , n22356 );
    not g37396 ( n34627 , n32781 );
    nor g37397 ( n3160 , n35509 , n23726 );
    and g37398 ( n20194 , n22189 , n29747 );
    or g37399 ( n7392 , n27961 , n40157 );
    xnor g37400 ( n6980 , n12837 , n20098 );
    not g37401 ( n18202 , n40276 );
    or g37402 ( n13593 , n9474 , n41779 );
    or g37403 ( n35594 , n37882 , n32242 );
    or g37404 ( n14567 , n32100 , n39464 );
    and g37405 ( n24537 , n38830 , n4230 );
    xnor g37406 ( n40397 , n23371 , n16478 );
    nor g37407 ( n28292 , n25781 , n8581 );
    nor g37408 ( n33575 , n24625 , n32214 );
    nor g37409 ( n18319 , n8494 , n18486 );
    not g37410 ( n39852 , n4746 );
    xnor g37411 ( n31581 , n5759 , n5764 );
    nor g37412 ( n7756 , n16532 , n18166 );
    or g37413 ( n11474 , n29596 , n7964 );
    nor g37414 ( n34767 , n23398 , n33421 );
    or g37415 ( n9643 , n394 , n11392 );
    or g37416 ( n12486 , n5881 , n37363 );
    or g37417 ( n5732 , n4140 , n40380 );
    nor g37418 ( n5717 , n26168 , n7893 );
    xnor g37419 ( n33599 , n40513 , n32613 );
    or g37420 ( n40327 , n15064 , n8144 );
    nor g37421 ( n36869 , n35488 , n27896 );
    or g37422 ( n19096 , n8750 , n40612 );
    not g37423 ( n20141 , n20157 );
    or g37424 ( n922 , n31095 , n37250 );
    or g37425 ( n14542 , n28149 , n40317 );
    or g37426 ( n32615 , n12112 , n24902 );
    nor g37427 ( n21526 , n18866 , n36832 );
    not g37428 ( n19471 , n30877 );
    or g37429 ( n9963 , n11476 , n38731 );
    not g37430 ( n26916 , n24846 );
    or g37431 ( n39894 , n21334 , n1961 );
    or g37432 ( n31642 , n28594 , n25907 );
    or g37433 ( n32554 , n1416 , n1705 );
    nor g37434 ( n755 , n16969 , n6942 );
    xnor g37435 ( n37276 , n2862 , n42634 );
    and g37436 ( n13277 , n24082 , n34420 );
    and g37437 ( n33108 , n37070 , n42574 );
    or g37438 ( n3201 , n28444 , n15733 );
    or g37439 ( n28829 , n32245 , n3535 );
    and g37440 ( n11320 , n20257 , n25079 );
    and g37441 ( n42779 , n36068 , n17146 );
    nor g37442 ( n14167 , n17182 , n26479 );
    or g37443 ( n21908 , n19197 , n6359 );
    xnor g37444 ( n11153 , n35727 , n8479 );
    xnor g37445 ( n37026 , n174 , n871 );
    or g37446 ( n22338 , n11288 , n22681 );
    not g37447 ( n37662 , n25592 );
    nor g37448 ( n41094 , n20878 , n13307 );
    xnor g37449 ( n34098 , n25701 , n11984 );
    or g37450 ( n34825 , n33027 , n42001 );
    xnor g37451 ( n24654 , n38371 , n17218 );
    not g37452 ( n10392 , n35358 );
    or g37453 ( n19854 , n41040 , n33184 );
    xnor g37454 ( n7298 , n35727 , n10170 );
    and g37455 ( n42311 , n38705 , n34236 );
    or g37456 ( n5427 , n21044 , n37993 );
    and g37457 ( n11797 , n4832 , n27858 );
    and g37458 ( n34069 , n4939 , n41028 );
    or g37459 ( n7945 , n39612 , n40787 );
    not g37460 ( n5718 , n41321 );
    or g37461 ( n35396 , n12848 , n34793 );
    or g37462 ( n27729 , n15096 , n31368 );
    not g37463 ( n40740 , n38481 );
    and g37464 ( n30852 , n329 , n13125 );
    and g37465 ( n33530 , n18599 , n595 );
    or g37466 ( n36725 , n21201 , n10965 );
    or g37467 ( n28656 , n23444 , n19085 );
    nor g37468 ( n12688 , n32261 , n41670 );
    or g37469 ( n39771 , n6815 , n27738 );
    or g37470 ( n18160 , n17908 , n6328 );
    nor g37471 ( n32113 , n6303 , n39749 );
    or g37472 ( n38726 , n28954 , n360 );
    or g37473 ( n9094 , n3318 , n38519 );
    xnor g37474 ( n19085 , n10176 , n20808 );
    or g37475 ( n40007 , n9084 , n31095 );
    and g37476 ( n6006 , n36748 , n18094 );
    or g37477 ( n39099 , n36376 , n16844 );
    or g37478 ( n28399 , n24183 , n340 );
    xnor g37479 ( n41231 , n40698 , n21227 );
    or g37480 ( n28310 , n10460 , n38505 );
    and g37481 ( n23998 , n36329 , n34147 );
    not g37482 ( n34698 , n31775 );
    xnor g37483 ( n26049 , n42064 , n40676 );
    or g37484 ( n20779 , n38487 , n24986 );
    or g37485 ( n28406 , n32347 , n21856 );
    and g37486 ( n8361 , n784 , n24493 );
    xnor g37487 ( n25860 , n28443 , n42532 );
    not g37488 ( n7276 , n11011 );
    nor g37489 ( n40816 , n24640 , n21556 );
    and g37490 ( n32748 , n20692 , n11839 );
    not g37491 ( n26799 , n39585 );
    not g37492 ( n37031 , n20792 );
    or g37493 ( n5784 , n13483 , n28289 );
    not g37494 ( n22888 , n31764 );
    nor g37495 ( n11114 , n39198 , n5155 );
    or g37496 ( n10252 , n6025 , n25252 );
    or g37497 ( n30876 , n4670 , n33777 );
    or g37498 ( n40856 , n33972 , n41624 );
    not g37499 ( n24423 , n25610 );
    nor g37500 ( n21844 , n22109 , n40859 );
    not g37501 ( n1385 , n24381 );
    or g37502 ( n24458 , n37031 , n39616 );
    not g37503 ( n10192 , n30989 );
    or g37504 ( n29541 , n12383 , n10742 );
    xnor g37505 ( n30026 , n37829 , n9308 );
    or g37506 ( n37394 , n11800 , n36760 );
    xnor g37507 ( n38301 , n7922 , n6904 );
    and g37508 ( n1444 , n6261 , n42259 );
    nor g37509 ( n2708 , n33586 , n22503 );
    nor g37510 ( n16714 , n10598 , n37010 );
    or g37511 ( n7368 , n8841 , n1206 );
    or g37512 ( n36957 , n25343 , n42411 );
    and g37513 ( n12562 , n22672 , n13202 );
    and g37514 ( n2180 , n12391 , n36495 );
    xnor g37515 ( n12042 , n21381 , n26914 );
    not g37516 ( n34687 , n19651 );
    xnor g37517 ( n34174 , n3248 , n24416 );
    and g37518 ( n30974 , n34313 , n6918 );
    and g37519 ( n8945 , n30682 , n11462 );
    and g37520 ( n8712 , n27056 , n28460 );
    nor g37521 ( n31644 , n17578 , n21925 );
    not g37522 ( n16866 , n6260 );
    or g37523 ( n30586 , n25273 , n6299 );
    or g37524 ( n42764 , n39227 , n15292 );
    nor g37525 ( n15175 , n5964 , n41787 );
    nor g37526 ( n12765 , n33838 , n12847 );
    or g37527 ( n35527 , n33744 , n3676 );
    and g37528 ( n11941 , n20789 , n32857 );
    not g37529 ( n26363 , n35480 );
    and g37530 ( n25900 , n26460 , n23581 );
    or g37531 ( n20579 , n36117 , n18132 );
    xnor g37532 ( n20881 , n4185 , n42604 );
    or g37533 ( n41024 , n12186 , n8033 );
    not g37534 ( n16280 , n7845 );
    nor g37535 ( n857 , n38029 , n14939 );
    or g37536 ( n5954 , n17021 , n22379 );
    not g37537 ( n36222 , n10457 );
    not g37538 ( n29601 , n24832 );
    and g37539 ( n26946 , n41451 , n992 );
    and g37540 ( n441 , n15203 , n35380 );
    xnor g37541 ( n42142 , n25849 , n29288 );
    and g37542 ( n21562 , n32272 , n33110 );
    and g37543 ( n173 , n6081 , n2543 );
    and g37544 ( n37891 , n6317 , n16225 );
    or g37545 ( n1427 , n11708 , n35761 );
    or g37546 ( n10265 , n15681 , n11142 );
    not g37547 ( n16803 , n10442 );
    not g37548 ( n31069 , n4912 );
    and g37549 ( n28723 , n23731 , n41164 );
    or g37550 ( n8555 , n10873 , n26147 );
    or g37551 ( n5648 , n5358 , n15365 );
    or g37552 ( n9305 , n34292 , n31323 );
    or g37553 ( n5895 , n28643 , n19838 );
    not g37554 ( n38939 , n7963 );
    nor g37555 ( n13049 , n42272 , n20746 );
    not g37556 ( n15282 , n28843 );
    or g37557 ( n10870 , n2655 , n11970 );
    and g37558 ( n42603 , n8935 , n32004 );
    or g37559 ( n28198 , n20775 , n35695 );
    nor g37560 ( n6271 , n17272 , n29738 );
    nor g37561 ( n4262 , n32874 , n18300 );
    and g37562 ( n18068 , n20335 , n25773 );
    and g37563 ( n36051 , n27224 , n28655 );
    or g37564 ( n34272 , n24836 , n40848 );
    or g37565 ( n21940 , n19309 , n17015 );
    not g37566 ( n4218 , n6379 );
    or g37567 ( n18252 , n12841 , n37572 );
    or g37568 ( n10421 , n10269 , n31091 );
    xnor g37569 ( n14194 , n21534 , n14899 );
    nor g37570 ( n32316 , n35887 , n2286 );
    not g37571 ( n22432 , n21117 );
    not g37572 ( n21253 , n40671 );
    or g37573 ( n23128 , n22523 , n12439 );
    not g37574 ( n478 , n34922 );
    nor g37575 ( n4240 , n34065 , n15067 );
    xnor g37576 ( n15733 , n16441 , n34565 );
    and g37577 ( n31513 , n39960 , n27940 );
    or g37578 ( n39584 , n4303 , n7363 );
    or g37579 ( n21588 , n28947 , n37224 );
    or g37580 ( n5293 , n12765 , n5761 );
    xnor g37581 ( n16770 , n5441 , n30355 );
    or g37582 ( n27462 , n39506 , n3856 );
    nor g37583 ( n24852 , n30110 , n5989 );
    or g37584 ( n1671 , n3508 , n36393 );
    and g37585 ( n32149 , n4261 , n33598 );
    and g37586 ( n22513 , n26907 , n30986 );
    xnor g37587 ( n13306 , n4334 , n9750 );
    and g37588 ( n41957 , n8089 , n6206 );
    nor g37589 ( n39422 , n36181 , n40932 );
    or g37590 ( n41821 , n17780 , n12433 );
    not g37591 ( n25756 , n29711 );
    nor g37592 ( n9444 , n38762 , n6684 );
    not g37593 ( n2060 , n29271 );
    xnor g37594 ( n2459 , n549 , n23488 );
    not g37595 ( n25286 , n12362 );
    and g37596 ( n28056 , n16936 , n19587 );
    or g37597 ( n21916 , n21111 , n18377 );
    not g37598 ( n10183 , n1784 );
    or g37599 ( n34336 , n11295 , n27261 );
    or g37600 ( n24429 , n39815 , n36983 );
    or g37601 ( n19050 , n35224 , n42179 );
    not g37602 ( n16909 , n1450 );
    and g37603 ( n18170 , n7844 , n41347 );
    or g37604 ( n22256 , n23990 , n33494 );
    xnor g37605 ( n41271 , n15812 , n27894 );
    or g37606 ( n42869 , n38405 , n31263 );
    or g37607 ( n21932 , n17853 , n8977 );
    not g37608 ( n16124 , n36263 );
    or g37609 ( n34314 , n38119 , n22830 );
    or g37610 ( n40167 , n2012 , n10913 );
    or g37611 ( n39101 , n21695 , n35531 );
    or g37612 ( n19377 , n15075 , n25847 );
    and g37613 ( n17512 , n9828 , n3707 );
    or g37614 ( n21370 , n33725 , n32101 );
    or g37615 ( n30639 , n2316 , n17404 );
    nor g37616 ( n20315 , n17906 , n33008 );
    nor g37617 ( n31737 , n37732 , n23837 );
    nor g37618 ( n26698 , n34292 , n29533 );
    and g37619 ( n37010 , n30095 , n41012 );
    and g37620 ( n42367 , n8282 , n1140 );
    not g37621 ( n32371 , n41939 );
    or g37622 ( n16167 , n3396 , n42704 );
    nor g37623 ( n18222 , n1730 , n24984 );
    and g37624 ( n40303 , n30716 , n15723 );
    or g37625 ( n20139 , n5573 , n16686 );
    and g37626 ( n35273 , n25953 , n22277 );
    and g37627 ( n25298 , n12681 , n36237 );
    and g37628 ( n37984 , n39125 , n15159 );
    xnor g37629 ( n8135 , n21973 , n14448 );
    or g37630 ( n24 , n1353 , n29630 );
    or g37631 ( n29496 , n29437 , n29260 );
    xnor g37632 ( n11927 , n18530 , n18504 );
    or g37633 ( n4103 , n3466 , n27058 );
    nor g37634 ( n3851 , n26990 , n29383 );
    xnor g37635 ( n42656 , n2174 , n27401 );
    and g37636 ( n18140 , n2950 , n19732 );
    xnor g37637 ( n33299 , n34562 , n5198 );
    or g37638 ( n42676 , n18464 , n22218 );
    and g37639 ( n21098 , n23609 , n40789 );
    not g37640 ( n3524 , n33563 );
    or g37641 ( n21853 , n19728 , n3771 );
    or g37642 ( n22860 , n33105 , n9633 );
    or g37643 ( n20149 , n25537 , n14053 );
    or g37644 ( n17612 , n34485 , n22988 );
    nor g37645 ( n15455 , n32328 , n15457 );
    xnor g37646 ( n32996 , n26402 , n23293 );
    or g37647 ( n1384 , n40375 , n8578 );
    nor g37648 ( n9700 , n31861 , n3382 );
    nor g37649 ( n22598 , n19300 , n30028 );
    and g37650 ( n25367 , n8196 , n9086 );
    not g37651 ( n34404 , n24045 );
    or g37652 ( n9972 , n5927 , n16169 );
    and g37653 ( n37791 , n14698 , n17531 );
    not g37654 ( n31107 , n16253 );
    nor g37655 ( n20751 , n9902 , n9071 );
    xnor g37656 ( n30879 , n255 , n1751 );
    or g37657 ( n1285 , n16789 , n30848 );
    nor g37658 ( n22711 , n29568 , n35486 );
    or g37659 ( n12933 , n36131 , n31509 );
    or g37660 ( n9888 , n20810 , n23703 );
    not g37661 ( n2463 , n31640 );
    nor g37662 ( n3947 , n35301 , n19404 );
    or g37663 ( n11513 , n15528 , n25626 );
    xnor g37664 ( n2570 , n39556 , n40857 );
    not g37665 ( n21893 , n23847 );
    not g37666 ( n31043 , n7681 );
    or g37667 ( n15654 , n14945 , n41799 );
    and g37668 ( n18917 , n22571 , n33988 );
    or g37669 ( n17660 , n8859 , n35685 );
    nor g37670 ( n15581 , n19665 , n26914 );
    and g37671 ( n42280 , n36472 , n14880 );
    not g37672 ( n16676 , n25044 );
    nor g37673 ( n2045 , n37017 , n5901 );
    nor g37674 ( n17411 , n38563 , n29008 );
    or g37675 ( n41734 , n13488 , n36021 );
    and g37676 ( n10010 , n17715 , n1117 );
    nor g37677 ( n38698 , n19532 , n13681 );
    and g37678 ( n22639 , n42252 , n28693 );
    or g37679 ( n15174 , n39991 , n31057 );
    and g37680 ( n3648 , n12466 , n23474 );
    or g37681 ( n14599 , n36844 , n32510 );
    or g37682 ( n14011 , n4668 , n11709 );
    or g37683 ( n38079 , n35287 , n31102 );
    nor g37684 ( n27027 , n33190 , n13733 );
    and g37685 ( n29139 , n35687 , n28260 );
    xnor g37686 ( n31119 , n28673 , n28206 );
    and g37687 ( n2301 , n6184 , n3050 );
    or g37688 ( n25166 , n18421 , n14057 );
    or g37689 ( n16098 , n13820 , n22928 );
    xnor g37690 ( n20948 , n22263 , n1518 );
    or g37691 ( n16989 , n28996 , n41337 );
    and g37692 ( n21433 , n9593 , n4297 );
    nor g37693 ( n20452 , n139 , n8448 );
    or g37694 ( n25167 , n6240 , n7938 );
    nor g37695 ( n498 , n9989 , n28284 );
    or g37696 ( n10655 , n23462 , n21581 );
    not g37697 ( n32506 , n11879 );
    xnor g37698 ( n10416 , n36046 , n12670 );
    xnor g37699 ( n13936 , n41053 , n19909 );
    or g37700 ( n23573 , n8787 , n23547 );
    and g37701 ( n17998 , n19871 , n10797 );
    nor g37702 ( n5719 , n35086 , n4656 );
    not g37703 ( n40870 , n6473 );
    or g37704 ( n36016 , n991 , n5964 );
    or g37705 ( n2644 , n18314 , n7640 );
    not g37706 ( n41230 , n16119 );
    or g37707 ( n4291 , n15131 , n16372 );
    and g37708 ( n31530 , n19162 , n23643 );
    xnor g37709 ( n8836 , n898 , n36528 );
    or g37710 ( n32260 , n41705 , n26809 );
    and g37711 ( n6912 , n31310 , n19951 );
    xnor g37712 ( n36638 , n36998 , n28786 );
    or g37713 ( n9231 , n30455 , n42762 );
    xnor g37714 ( n38477 , n21534 , n30067 );
    or g37715 ( n22265 , n24588 , n36790 );
    xnor g37716 ( n8190 , n4495 , n29452 );
    not g37717 ( n37250 , n8734 );
    and g37718 ( n29970 , n6731 , n27716 );
    xnor g37719 ( n4844 , n39104 , n23127 );
    not g37720 ( n4869 , n21293 );
    or g37721 ( n24941 , n19229 , n10012 );
    not g37722 ( n16320 , n40299 );
    and g37723 ( n41021 , n39622 , n23316 );
    not g37724 ( n38636 , n7042 );
    not g37725 ( n14055 , n28843 );
    xnor g37726 ( n32953 , n2174 , n673 );
    xnor g37727 ( n12238 , n12281 , n34979 );
    or g37728 ( n29289 , n19380 , n16682 );
    xnor g37729 ( n15060 , n21534 , n196 );
    not g37730 ( n42447 , n17467 );
    or g37731 ( n5944 , n16462 , n36555 );
    and g37732 ( n38067 , n23436 , n6015 );
    or g37733 ( n34398 , n33398 , n11410 );
    nor g37734 ( n36441 , n31351 , n39474 );
    or g37735 ( n11975 , n29178 , n14154 );
    and g37736 ( n42157 , n6697 , n21453 );
    nor g37737 ( n31649 , n15437 , n23604 );
    not g37738 ( n30846 , n458 );
    or g37739 ( n3697 , n1995 , n10964 );
    or g37740 ( n8405 , n7829 , n41319 );
    xnor g37741 ( n5270 , n3068 , n13448 );
    not g37742 ( n347 , n21825 );
    and g37743 ( n20351 , n17285 , n38880 );
    and g37744 ( n4598 , n16347 , n25379 );
    xnor g37745 ( n5810 , n42064 , n15904 );
    or g37746 ( n7721 , n39970 , n41243 );
    or g37747 ( n31910 , n38142 , n5295 );
    xnor g37748 ( n19555 , n31099 , n38063 );
    or g37749 ( n30710 , n19795 , n10707 );
    and g37750 ( n37728 , n31863 , n19059 );
    xnor g37751 ( n11612 , n38128 , n31383 );
    nor g37752 ( n36877 , n30725 , n27842 );
    or g37753 ( n29 , n31721 , n4798 );
    or g37754 ( n5797 , n5543 , n14009 );
    or g37755 ( n2169 , n41139 , n13866 );
    or g37756 ( n17864 , n12752 , n39804 );
    and g37757 ( n15940 , n6506 , n10705 );
    not g37758 ( n13967 , n12087 );
    and g37759 ( n27132 , n19738 , n8557 );
    or g37760 ( n38055 , n8493 , n15065 );
    not g37761 ( n11178 , n15956 );
    xnor g37762 ( n28217 , n41358 , n3941 );
    nor g37763 ( n29574 , n23761 , n4803 );
    or g37764 ( n21883 , n33275 , n18167 );
    and g37765 ( n3945 , n24890 , n744 );
    not g37766 ( n33973 , n19178 );
    or g37767 ( n39527 , n1352 , n9054 );
    and g37768 ( n13170 , n8522 , n38610 );
    nor g37769 ( n31836 , n59 , n871 );
    not g37770 ( n3740 , n19236 );
    and g37771 ( n4747 , n13408 , n20011 );
    xnor g37772 ( n15145 , n105 , n29228 );
    or g37773 ( n22961 , n34552 , n36344 );
    and g37774 ( n17025 , n13001 , n34482 );
    or g37775 ( n35627 , n19784 , n15262 );
    xnor g37776 ( n18303 , n5144 , n2333 );
    nor g37777 ( n2310 , n23040 , n30400 );
    or g37778 ( n20703 , n7364 , n17576 );
    or g37779 ( n20129 , n26040 , n33445 );
    and g37780 ( n14373 , n34056 , n14525 );
    or g37781 ( n23269 , n1151 , n42452 );
    or g37782 ( n37079 , n30578 , n6633 );
    xnor g37783 ( n10652 , n16746 , n28598 );
    and g37784 ( n22517 , n6585 , n10431 );
    or g37785 ( n15924 , n5959 , n27967 );
    and g37786 ( n39193 , n31408 , n30954 );
    and g37787 ( n23206 , n14193 , n13020 );
    not g37788 ( n24687 , n30438 );
    or g37789 ( n16322 , n31991 , n28028 );
    or g37790 ( n36472 , n6769 , n13687 );
    or g37791 ( n13541 , n41297 , n10400 );
    or g37792 ( n1443 , n39659 , n35365 );
    and g37793 ( n5770 , n34111 , n24487 );
    and g37794 ( n27203 , n23305 , n7662 );
    or g37795 ( n12295 , n20717 , n560 );
    or g37796 ( n19597 , n24454 , n39173 );
    xnor g37797 ( n4864 , n20487 , n33619 );
    not g37798 ( n42558 , n7975 );
    nor g37799 ( n38019 , n17006 , n24954 );
    and g37800 ( n8420 , n41483 , n33326 );
    xnor g37801 ( n25450 , n18530 , n36485 );
    and g37802 ( n30386 , n13583 , n3452 );
    not g37803 ( n24843 , n24377 );
    and g37804 ( n16174 , n15575 , n3752 );
    xnor g37805 ( n5956 , n20831 , n14707 );
    or g37806 ( n38705 , n9504 , n34288 );
    and g37807 ( n33363 , n10276 , n19341 );
    or g37808 ( n16950 , n41294 , n31139 );
    nor g37809 ( n10147 , n18027 , n22506 );
    not g37810 ( n35553 , n5605 );
    or g37811 ( n19048 , n28213 , n26962 );
    nor g37812 ( n19487 , n39182 , n699 );
    not g37813 ( n34796 , n25649 );
    xnor g37814 ( n32917 , n105 , n30472 );
    not g37815 ( n12344 , n12907 );
    xnor g37816 ( n21887 , n11931 , n31988 );
    not g37817 ( n20209 , n37115 );
    nor g37818 ( n18911 , n23324 , n11355 );
    xnor g37819 ( n17115 , n302 , n24215 );
    and g37820 ( n31420 , n2560 , n2522 );
    nor g37821 ( n3149 , n14496 , n2843 );
    or g37822 ( n40731 , n35649 , n37185 );
    xnor g37823 ( n13798 , n15972 , n12122 );
    or g37824 ( n34207 , n35963 , n5631 );
    xnor g37825 ( n39136 , n37073 , n34565 );
    or g37826 ( n18195 , n2387 , n27616 );
    xnor g37827 ( n24499 , n21880 , n23299 );
    nor g37828 ( n32714 , n13175 , n12780 );
    nor g37829 ( n20606 , n18424 , n25238 );
    nor g37830 ( n40066 , n32548 , n14213 );
    not g37831 ( n24164 , n12240 );
    or g37832 ( n3963 , n19067 , n19548 );
    or g37833 ( n21127 , n4535 , n9541 );
    not g37834 ( n25607 , n25936 );
    or g37835 ( n4867 , n27311 , n24229 );
    not g37836 ( n11059 , n4508 );
    nor g37837 ( n38718 , n5964 , n41928 );
    nor g37838 ( n27875 , n38059 , n5999 );
    or g37839 ( n10817 , n11368 , n3399 );
    and g37840 ( n30114 , n39242 , n14845 );
    not g37841 ( n5254 , n8066 );
    not g37842 ( n36250 , n17625 );
    or g37843 ( n25867 , n23233 , n734 );
    or g37844 ( n39343 , n26992 , n9913 );
    or g37845 ( n34655 , n39539 , n32409 );
    or g37846 ( n1473 , n2110 , n41562 );
    or g37847 ( n4514 , n22175 , n30800 );
    and g37848 ( n23693 , n38879 , n39377 );
    or g37849 ( n979 , n15064 , n22729 );
    or g37850 ( n33925 , n18698 , n13113 );
    and g37851 ( n42857 , n32459 , n9018 );
    or g37852 ( n19408 , n27261 , n15780 );
    nor g37853 ( n1732 , n22473 , n4593 );
    and g37854 ( n42546 , n37135 , n278 );
    not g37855 ( n13683 , n19607 );
    xnor g37856 ( n10142 , n29423 , n20361 );
    xnor g37857 ( n3032 , n21559 , n12847 );
    or g37858 ( n8371 , n10608 , n33718 );
    not g37859 ( n39991 , n32716 );
    and g37860 ( n26604 , n17591 , n12445 );
    not g37861 ( n13422 , n62 );
    or g37862 ( n38680 , n29898 , n37890 );
    nor g37863 ( n15262 , n17120 , n41032 );
    not g37864 ( n28347 , n29948 );
    or g37865 ( n11137 , n19668 , n713 );
    and g37866 ( n8101 , n42822 , n24533 );
    or g37867 ( n22594 , n17241 , n42899 );
    and g37868 ( n38833 , n39555 , n2150 );
    and g37869 ( n22146 , n35237 , n26486 );
    or g37870 ( n36206 , n12112 , n38127 );
    not g37871 ( n25409 , n30569 );
    or g37872 ( n26900 , n13457 , n14487 );
    or g37873 ( n6737 , n5402 , n11237 );
    xnor g37874 ( n15626 , n38899 , n23466 );
    or g37875 ( n15557 , n33981 , n9936 );
    not g37876 ( n7016 , n144 );
    or g37877 ( n10340 , n22989 , n10591 );
    or g37878 ( n22810 , n28323 , n38140 );
    and g37879 ( n9858 , n13327 , n41619 );
    nor g37880 ( n1068 , n35009 , n1988 );
    not g37881 ( n2370 , n40375 );
    or g37882 ( n39682 , n24454 , n37395 );
    or g37883 ( n4792 , n39915 , n36235 );
    xnor g37884 ( n28394 , n24546 , n11196 );
    or g37885 ( n29482 , n36983 , n41855 );
    and g37886 ( n32472 , n4205 , n28907 );
    or g37887 ( n365 , n11008 , n27096 );
    or g37888 ( n35955 , n34485 , n9514 );
    or g37889 ( n15243 , n42052 , n31271 );
    xnor g37890 ( n4265 , n8591 , n35848 );
    not g37891 ( n19818 , n19113 );
    and g37892 ( n29914 , n5452 , n4232 );
    and g37893 ( n41438 , n1056 , n20182 );
    or g37894 ( n9104 , n41723 , n34796 );
    not g37895 ( n18563 , n15132 );
    and g37896 ( n27816 , n8385 , n17447 );
    or g37897 ( n1573 , n35321 , n29250 );
    and g37898 ( n27192 , n33157 , n15534 );
    and g37899 ( n34339 , n23890 , n10023 );
    nor g37900 ( n13101 , n5320 , n39616 );
    or g37901 ( n28704 , n10998 , n27092 );
    and g37902 ( n9464 , n23363 , n16070 );
    and g37903 ( n33878 , n18636 , n32561 );
    xnor g37904 ( n22356 , n13444 , n882 );
    or g37905 ( n4342 , n857 , n9967 );
    or g37906 ( n3489 , n11877 , n19796 );
    or g37907 ( n21743 , n32711 , n583 );
    xnor g37908 ( n24507 , n42064 , n41839 );
    or g37909 ( n24963 , n19464 , n29780 );
    and g37910 ( n37129 , n9083 , n21576 );
    not g37911 ( n31001 , n35288 );
    or g37912 ( n39285 , n19802 , n33775 );
    and g37913 ( n9184 , n11835 , n22690 );
    or g37914 ( n26373 , n40041 , n25610 );
    not g37915 ( n11932 , n14367 );
    or g37916 ( n10432 , n5220 , n12400 );
    nor g37917 ( n40850 , n1002 , n12296 );
    or g37918 ( n16972 , n39942 , n40323 );
    not g37919 ( n31671 , n33545 );
    and g37920 ( n8679 , n21724 , n36202 );
    xnor g37921 ( n34943 , n31989 , n33254 );
    not g37922 ( n3835 , n22426 );
    or g37923 ( n25229 , n40769 , n15063 );
    and g37924 ( n5409 , n3114 , n25883 );
    or g37925 ( n11776 , n313 , n23649 );
    and g37926 ( n27862 , n9681 , n20529 );
    not g37927 ( n1386 , n29537 );
    xnor g37928 ( n31931 , n27789 , n24537 );
    or g37929 ( n23281 , n8806 , n4612 );
    or g37930 ( n12964 , n19803 , n29210 );
    or g37931 ( n8513 , n38307 , n11082 );
    and g37932 ( n4941 , n6639 , n21162 );
    or g37933 ( n5619 , n27127 , n38910 );
    and g37934 ( n15479 , n18740 , n31757 );
    or g37935 ( n22058 , n35977 , n42471 );
    or g37936 ( n41510 , n7375 , n21555 );
    or g37937 ( n37999 , n31140 , n1534 );
    not g37938 ( n13735 , n15693 );
    or g37939 ( n31880 , n29187 , n10609 );
    or g37940 ( n25728 , n10496 , n2514 );
    or g37941 ( n38087 , n448 , n39213 );
    not g37942 ( n28373 , n25974 );
    xnor g37943 ( n21741 , n32253 , n980 );
    nor g37944 ( n8440 , n18391 , n37240 );
    nor g37945 ( n569 , n19260 , n7354 );
    not g37946 ( n6761 , n12687 );
    or g37947 ( n41372 , n5896 , n30090 );
    xnor g37948 ( n41867 , n6621 , n14216 );
    not g37949 ( n25700 , n22009 );
    nor g37950 ( n23007 , n15325 , n22727 );
    or g37951 ( n25758 , n24016 , n23414 );
    or g37952 ( n32084 , n19486 , n5250 );
    xnor g37953 ( n39070 , n25985 , n3508 );
    or g37954 ( n31833 , n11897 , n17899 );
    xnor g37955 ( n19501 , n38899 , n6990 );
    and g37956 ( n29965 , n5887 , n31365 );
    and g37957 ( n30101 , n32941 , n30747 );
    not g37958 ( n35876 , n41603 );
    or g37959 ( n37934 , n12129 , n42310 );
    xnor g37960 ( n15648 , n16746 , n33248 );
    and g37961 ( n22552 , n35684 , n20402 );
    or g37962 ( n75 , n34305 , n35171 );
    xnor g37963 ( n32193 , n14312 , n16364 );
    not g37964 ( n12285 , n12962 );
    not g37965 ( n2456 , n33788 );
    not g37966 ( n18702 , n1903 );
    or g37967 ( n38010 , n15687 , n36327 );
    or g37968 ( n23194 , n34017 , n41878 );
    and g37969 ( n2848 , n26472 , n40800 );
    or g37970 ( n21093 , n34643 , n13866 );
    and g37971 ( n13605 , n8524 , n32096 );
    and g37972 ( n28904 , n34435 , n10046 );
    and g37973 ( n17947 , n16517 , n13842 );
    and g37974 ( n6869 , n38265 , n31287 );
    and g37975 ( n34560 , n37196 , n1087 );
    not g37976 ( n4388 , n33313 );
    xnor g37977 ( n39051 , n13444 , n30867 );
    and g37978 ( n36378 , n17354 , n15991 );
    and g37979 ( n22701 , n26697 , n41138 );
    or g37980 ( n39370 , n41584 , n9303 );
    or g37981 ( n20465 , n41250 , n10230 );
    or g37982 ( n16986 , n15185 , n30655 );
    and g37983 ( n12924 , n17189 , n38616 );
    and g37984 ( n12243 , n5056 , n12458 );
    and g37985 ( n30479 , n17697 , n1282 );
    or g37986 ( n4203 , n41767 , n9710 );
    xnor g37987 ( n1809 , n18350 , n38734 );
    not g37988 ( n31986 , n19583 );
    not g37989 ( n29906 , n35121 );
    or g37990 ( n24028 , n8082 , n2515 );
    and g37991 ( n11695 , n25139 , n41801 );
    nor g37992 ( n20701 , n8634 , n29160 );
    xnor g37993 ( n11329 , n2005 , n33447 );
    not g37994 ( n29426 , n28826 );
    not g37995 ( n38826 , n42907 );
    not g37996 ( n4397 , n22916 );
    nor g37997 ( n28291 , n26680 , n6105 );
    or g37998 ( n34247 , n7475 , n8963 );
    nor g37999 ( n8245 , n34323 , n41416 );
    nor g38000 ( n10413 , n36636 , n34555 );
    or g38001 ( n4216 , n26225 , n2565 );
    or g38002 ( n35929 , n6905 , n20478 );
    nor g38003 ( n9998 , n14707 , n11734 );
    or g38004 ( n42889 , n37851 , n13634 );
    nor g38005 ( n26867 , n21846 , n10452 );
    or g38006 ( n31450 , n33951 , n2793 );
    or g38007 ( n39006 , n17725 , n36995 );
    nor g38008 ( n14049 , n2199 , n41839 );
    or g38009 ( n32861 , n37239 , n21440 );
    nor g38010 ( n3056 , n28617 , n25453 );
    or g38011 ( n24409 , n19864 , n569 );
    xnor g38012 ( n34245 , n18678 , n25228 );
    or g38013 ( n6356 , n17984 , n3254 );
    and g38014 ( n11306 , n1801 , n35282 );
    and g38015 ( n24295 , n40027 , n13264 );
    and g38016 ( n21142 , n29676 , n29670 );
    nor g38017 ( n2167 , n17051 , n16775 );
    and g38018 ( n5475 , n12208 , n35627 );
    nor g38019 ( n34201 , n31792 , n3031 );
    or g38020 ( n2473 , n12275 , n23511 );
    or g38021 ( n26464 , n9108 , n17679 );
    not g38022 ( n39778 , n4934 );
    or g38023 ( n11919 , n11917 , n27111 );
    nor g38024 ( n27169 , n13801 , n21055 );
    and g38025 ( n3552 , n31160 , n35865 );
    not g38026 ( n8618 , n38675 );
    or g38027 ( n5972 , n12959 , n13695 );
    not g38028 ( n11670 , n36076 );
    and g38029 ( n1389 , n4774 , n5321 );
    or g38030 ( n41251 , n7685 , n32061 );
    or g38031 ( n16296 , n7196 , n7747 );
    or g38032 ( n39943 , n2825 , n32744 );
    or g38033 ( n1691 , n18221 , n2204 );
    not g38034 ( n16073 , n27125 );
    not g38035 ( n41906 , n1269 );
    not g38036 ( n14472 , n30956 );
    and g38037 ( n33940 , n1161 , n10726 );
    xnor g38038 ( n19586 , n32624 , n5386 );
    xnor g38039 ( n30201 , n185 , n36766 );
    or g38040 ( n28899 , n16161 , n34171 );
    not g38041 ( n5422 , n22574 );
    and g38042 ( n23079 , n24937 , n25422 );
    not g38043 ( n11509 , n38793 );
    not g38044 ( n13848 , n33662 );
    and g38045 ( n26098 , n26612 , n39209 );
    or g38046 ( n34512 , n41995 , n2112 );
    or g38047 ( n10942 , n32529 , n28157 );
    nor g38048 ( n39569 , n26279 , n1126 );
    and g38049 ( n42408 , n4691 , n9102 );
    xnor g38050 ( n20847 , n17220 , n38864 );
    nor g38051 ( n10094 , n15672 , n24313 );
    or g38052 ( n13087 , n8155 , n40554 );
    or g38053 ( n11158 , n4305 , n3046 );
    or g38054 ( n22410 , n20521 , n23031 );
    and g38055 ( n2591 , n4811 , n7625 );
    xnor g38056 ( n22148 , n7001 , n14449 );
    not g38057 ( n38175 , n23430 );
    nor g38058 ( n6586 , n39412 , n18879 );
    nor g38059 ( n29325 , n22243 , n37901 );
    and g38060 ( n34824 , n14097 , n24034 );
    and g38061 ( n39799 , n28126 , n23281 );
    nor g38062 ( n24615 , n6865 , n26159 );
    nor g38063 ( n9024 , n4941 , n11576 );
    and g38064 ( n37008 , n29467 , n16732 );
    or g38065 ( n4793 , n40710 , n13964 );
    or g38066 ( n41735 , n5403 , n25303 );
    nor g38067 ( n29411 , n920 , n37138 );
    and g38068 ( n41121 , n7628 , n16344 );
    or g38069 ( n41506 , n20250 , n358 );
    and g38070 ( n18771 , n8810 , n42087 );
    or g38071 ( n32066 , n29686 , n17287 );
    not g38072 ( n6852 , n15195 );
    or g38073 ( n3693 , n9319 , n28518 );
    or g38074 ( n18980 , n26113 , n9055 );
    nor g38075 ( n34535 , n29052 , n19909 );
    or g38076 ( n30351 , n1138 , n36619 );
    or g38077 ( n26833 , n30082 , n21663 );
    xnor g38078 ( n17973 , n41766 , n20887 );
    nor g38079 ( n37798 , n23351 , n16956 );
    or g38080 ( n35312 , n12495 , n19354 );
    xnor g38081 ( n40247 , n566 , n25161 );
    nor g38082 ( n39008 , n41781 , n8513 );
    nor g38083 ( n10912 , n39456 , n34041 );
    xnor g38084 ( n39942 , n17854 , n28380 );
    or g38085 ( n26045 , n21929 , n10205 );
    xnor g38086 ( n32721 , n24505 , n8808 );
    xnor g38087 ( n5316 , n23011 , n5896 );
    or g38088 ( n41325 , n35534 , n6818 );
    and g38089 ( n29488 , n37764 , n30898 );
    and g38090 ( n12553 , n25483 , n22856 );
    or g38091 ( n22080 , n21206 , n39503 );
    or g38092 ( n18594 , n23047 , n14571 );
    or g38093 ( n8435 , n28647 , n6772 );
    nor g38094 ( n24147 , n11352 , n9389 );
    xnor g38095 ( n28992 , n38378 , n8040 );
    xnor g38096 ( n36384 , n27900 , n12898 );
    or g38097 ( n2211 , n19662 , n29911 );
    or g38098 ( n15725 , n29425 , n17381 );
    or g38099 ( n28137 , n7613 , n30155 );
    and g38100 ( n22031 , n9499 , n33498 );
    xnor g38101 ( n26800 , n19760 , n33829 );
    nor g38102 ( n7117 , n8790 , n10410 );
    or g38103 ( n16524 , n9752 , n4368 );
    or g38104 ( n16816 , n39948 , n19310 );
    or g38105 ( n3183 , n26514 , n37697 );
    and g38106 ( n11033 , n18967 , n23203 );
    and g38107 ( n33113 , n12214 , n20898 );
    or g38108 ( n23100 , n21977 , n34267 );
    nor g38109 ( n9466 , n23783 , n21796 );
    nor g38110 ( n36312 , n12516 , n33969 );
    not g38111 ( n29256 , n874 );
    and g38112 ( n2592 , n36409 , n6830 );
    not g38113 ( n24831 , n19907 );
    and g38114 ( n32040 , n17969 , n551 );
    and g38115 ( n29197 , n21149 , n19297 );
    nor g38116 ( n16840 , n7286 , n29115 );
    nor g38117 ( n35491 , n17525 , n29931 );
    xnor g38118 ( n39205 , n4636 , n39591 );
    or g38119 ( n37504 , n29980 , n14586 );
    xnor g38120 ( n22068 , n37558 , n8494 );
    or g38121 ( n18684 , n20250 , n24878 );
    xnor g38122 ( n31894 , n760 , n27583 );
    and g38123 ( n36327 , n23911 , n34086 );
    nor g38124 ( n29075 , n39449 , n15040 );
    or g38125 ( n40672 , n2460 , n19639 );
    and g38126 ( n19590 , n9436 , n38765 );
    or g38127 ( n9731 , n4492 , n20899 );
    or g38128 ( n15551 , n4717 , n22640 );
    nor g38129 ( n14770 , n16143 , n10940 );
    or g38130 ( n13288 , n10384 , n14769 );
    nor g38131 ( n39973 , n31633 , n9565 );
    not g38132 ( n42531 , n25093 );
    xnor g38133 ( n15530 , n31956 , n33569 );
    not g38134 ( n21421 , n30575 );
    xnor g38135 ( n2566 , n36009 , n26946 );
    and g38136 ( n33988 , n21534 , n40221 );
    or g38137 ( n13431 , n22714 , n25206 );
    or g38138 ( n12539 , n20503 , n12975 );
    nor g38139 ( n28575 , n22290 , n21140 );
    nor g38140 ( n11703 , n33787 , n11770 );
    and g38141 ( n36517 , n7618 , n12231 );
    nor g38142 ( n29194 , n25588 , n14745 );
    and g38143 ( n10266 , n19938 , n21271 );
    xnor g38144 ( n40604 , n32731 , n27831 );
    or g38145 ( n7633 , n9597 , n13568 );
    or g38146 ( n17039 , n14016 , n9042 );
    xnor g38147 ( n36857 , n39214 , n11748 );
    or g38148 ( n10321 , n38119 , n37487 );
    not g38149 ( n14930 , n32847 );
    or g38150 ( n25934 , n29251 , n5261 );
    or g38151 ( n27777 , n37916 , n36866 );
    or g38152 ( n25278 , n8494 , n36517 );
    or g38153 ( n20281 , n23965 , n36687 );
    and g38154 ( n17696 , n36046 , n5430 );
    or g38155 ( n21706 , n42405 , n32846 );
    or g38156 ( n22575 , n27225 , n22061 );
    xnor g38157 ( n15811 , n3735 , n19852 );
    and g38158 ( n17663 , n42089 , n19287 );
    or g38159 ( n1101 , n26553 , n11829 );
    xnor g38160 ( n5998 , n136 , n32830 );
    or g38161 ( n23719 , n4752 , n39839 );
    not g38162 ( n34061 , n41463 );
    and g38163 ( n26595 , n771 , n31169 );
    or g38164 ( n39586 , n21752 , n23 );
    and g38165 ( n40387 , n21746 , n42505 );
    or g38166 ( n725 , n26234 , n32602 );
    not g38167 ( n25122 , n34320 );
    and g38168 ( n6524 , n24413 , n26552 );
    not g38169 ( n878 , n18387 );
    or g38170 ( n39982 , n27232 , n882 );
    and g38171 ( n35230 , n33741 , n31955 );
    or g38172 ( n3007 , n42409 , n12077 );
    nor g38173 ( n16494 , n17427 , n18976 );
    nor g38174 ( n4020 , n5964 , n34169 );
    not g38175 ( n29457 , n27478 );
    xnor g38176 ( n25088 , n41013 , n12937 );
    not g38177 ( n9870 , n40484 );
    not g38178 ( n32191 , n23008 );
    not g38179 ( n4341 , n35759 );
    xnor g38180 ( n32423 , n6688 , n20350 );
    nor g38181 ( n29763 , n3857 , n7932 );
    nor g38182 ( n25062 , n3462 , n39936 );
    or g38183 ( n42292 , n13404 , n7116 );
    not g38184 ( n36249 , n9285 );
    or g38185 ( n23123 , n19099 , n34664 );
    or g38186 ( n23840 , n38507 , n27540 );
    or g38187 ( n14566 , n8000 , n8567 );
    or g38188 ( n27589 , n405 , n30970 );
    and g38189 ( n21038 , n36838 , n10452 );
    not g38190 ( n10363 , n10706 );
    nor g38191 ( n11598 , n32132 , n20926 );
    or g38192 ( n13358 , n40625 , n4454 );
    and g38193 ( n32487 , n12223 , n12903 );
    not g38194 ( n35866 , n25649 );
    nor g38195 ( n8740 , n4370 , n41014 );
    and g38196 ( n12987 , n4330 , n36990 );
    or g38197 ( n5251 , n1702 , n28206 );
    xnor g38198 ( n26912 , n6625 , n40948 );
    or g38199 ( n8948 , n3868 , n21252 );
    and g38200 ( n10557 , n23770 , n32843 );
    not g38201 ( n5813 , n28949 );
    or g38202 ( n19386 , n14312 , n16364 );
    nor g38203 ( n11672 , n39266 , n18504 );
    and g38204 ( n38282 , n5781 , n14215 );
    nor g38205 ( n21884 , n4795 , n30007 );
    or g38206 ( n12801 , n3919 , n12235 );
    not g38207 ( n23502 , n4873 );
    xnor g38208 ( n20582 , n26345 , n39998 );
    not g38209 ( n20615 , n4841 );
    not g38210 ( n20681 , n19050 );
    or g38211 ( n11276 , n36303 , n12699 );
    and g38212 ( n39786 , n18900 , n2177 );
    or g38213 ( n41180 , n36738 , n17383 );
    and g38214 ( n32735 , n29818 , n4313 );
    or g38215 ( n22508 , n41592 , n14569 );
    and g38216 ( n24121 , n32851 , n14439 );
    or g38217 ( n29446 , n10967 , n1934 );
    or g38218 ( n39577 , n39327 , n15661 );
    not g38219 ( n6316 , n263 );
    nor g38220 ( n14195 , n14471 , n10170 );
    xnor g38221 ( n24976 , n34235 , n40879 );
    not g38222 ( n28006 , n39527 );
    or g38223 ( n37251 , n35483 , n24484 );
    not g38224 ( n30071 , n4708 );
    nor g38225 ( n40844 , n39444 , n24568 );
    or g38226 ( n3012 , n6573 , n32247 );
    and g38227 ( n12045 , n14355 , n1475 );
    and g38228 ( n38924 , n8185 , n18437 );
    nor g38229 ( n15444 , n6132 , n13944 );
    not g38230 ( n17144 , n7182 );
    xnor g38231 ( n11758 , n6688 , n26931 );
    or g38232 ( n24789 , n22002 , n32385 );
    or g38233 ( n30753 , n8040 , n27540 );
    xnor g38234 ( n35398 , n25292 , n20918 );
    and g38235 ( n36168 , n36246 , n28295 );
    or g38236 ( n21027 , n36389 , n34806 );
    and g38237 ( n29536 , n29222 , n41251 );
    and g38238 ( n36233 , n37349 , n438 );
    or g38239 ( n36156 , n5140 , n22714 );
    not g38240 ( n4961 , n768 );
    not g38241 ( n41761 , n11353 );
    xnor g38242 ( n9041 , n39217 , n5774 );
    or g38243 ( n2474 , n2701 , n15795 );
    or g38244 ( n34492 , n888 , n442 );
    not g38245 ( n25207 , n23541 );
    and g38246 ( n30839 , n39321 , n21585 );
    or g38247 ( n8497 , n14861 , n31306 );
    and g38248 ( n35779 , n18384 , n5326 );
    xnor g38249 ( n42282 , n34731 , n17002 );
    and g38250 ( n20816 , n32286 , n27496 );
    or g38251 ( n23794 , n6446 , n28082 );
    xnor g38252 ( n41341 , n35938 , n2901 );
    and g38253 ( n42328 , n1305 , n40535 );
    xnor g38254 ( n34926 , n16473 , n9518 );
    or g38255 ( n4846 , n20978 , n7833 );
    nor g38256 ( n26179 , n27697 , n3499 );
    xnor g38257 ( n1250 , n39921 , n28044 );
    xnor g38258 ( n40682 , n21973 , n28607 );
    or g38259 ( n11953 , n19459 , n1975 );
    nor g38260 ( n37665 , n22915 , n19081 );
    not g38261 ( n26904 , n16987 );
    xnor g38262 ( n42570 , n14311 , n15161 );
    or g38263 ( n5202 , n5564 , n7526 );
    and g38264 ( n30938 , n33535 , n630 );
    not g38265 ( n17175 , n10114 );
    not g38266 ( n8876 , n29206 );
    not g38267 ( n39195 , n15778 );
    or g38268 ( n20603 , n7180 , n18836 );
    xnor g38269 ( n28084 , n784 , n15639 );
    or g38270 ( n34291 , n14407 , n63 );
    not g38271 ( n4043 , n2513 );
    xnor g38272 ( n25876 , n35687 , n28260 );
    or g38273 ( n14079 , n37850 , n2565 );
    and g38274 ( n31333 , n26733 , n41522 );
    and g38275 ( n20375 , n4314 , n1033 );
    and g38276 ( n23366 , n13863 , n31745 );
    or g38277 ( n24050 , n34153 , n15315 );
    nor g38278 ( n24234 , n17193 , n25669 );
    not g38279 ( n3829 , n13966 );
    or g38280 ( n32934 , n33423 , n34412 );
    or g38281 ( n1881 , n15282 , n14664 );
    nor g38282 ( n21088 , n5685 , n13711 );
    not g38283 ( n1452 , n36338 );
    or g38284 ( n501 , n38249 , n16622 );
    not g38285 ( n20411 , n32001 );
    and g38286 ( n5879 , n24338 , n40395 );
    xnor g38287 ( n11414 , n20804 , n1122 );
    and g38288 ( n6192 , n21937 , n11450 );
    not g38289 ( n16699 , n13784 );
    and g38290 ( n17566 , n12407 , n40466 );
    nor g38291 ( n42083 , n8857 , n8980 );
    or g38292 ( n16213 , n41008 , n3788 );
    and g38293 ( n33502 , n24641 , n19977 );
    or g38294 ( n15644 , n6560 , n39984 );
    or g38295 ( n42914 , n2149 , n16066 );
    not g38296 ( n7622 , n9719 );
    not g38297 ( n19196 , n13009 );
    not g38298 ( n25668 , n21034 );
    or g38299 ( n1944 , n18314 , n34166 );
    not g38300 ( n421 , n2163 );
    and g38301 ( n29612 , n33100 , n9386 );
    or g38302 ( n13614 , n1567 , n13692 );
    or g38303 ( n29929 , n17452 , n15578 );
    xnor g38304 ( n26909 , n39415 , n6721 );
    not g38305 ( n27358 , n12170 );
    or g38306 ( n24969 , n26298 , n35994 );
    not g38307 ( n2935 , n23147 );
    and g38308 ( n35809 , n6376 , n22575 );
    or g38309 ( n26420 , n24315 , n23949 );
    or g38310 ( n15798 , n31924 , n26731 );
    or g38311 ( n21506 , n28774 , n40270 );
    not g38312 ( n27127 , n30826 );
    and g38313 ( n33997 , n105 , n15977 );
    and g38314 ( n5424 , n10844 , n41683 );
    or g38315 ( n31500 , n13480 , n42706 );
    nor g38316 ( n25737 , n22385 , n31247 );
    xnor g38317 ( n7608 , n21448 , n33873 );
    not g38318 ( n455 , n8649 );
    nor g38319 ( n37858 , n3770 , n41619 );
    and g38320 ( n30936 , n33559 , n14866 );
    nor g38321 ( n2121 , n33981 , n9837 );
    and g38322 ( n8979 , n20398 , n32621 );
    or g38323 ( n18098 , n17759 , n37994 );
    or g38324 ( n20392 , n40070 , n7988 );
    or g38325 ( n14565 , n33134 , n26000 );
    and g38326 ( n12227 , n22820 , n6471 );
    or g38327 ( n40651 , n32499 , n2217 );
    and g38328 ( n31856 , n42430 , n33163 );
    or g38329 ( n25646 , n29068 , n29485 );
    or g38330 ( n42587 , n34461 , n23243 );
    nor g38331 ( n36416 , n38290 , n16353 );
    xnor g38332 ( n20377 , n22296 , n26971 );
    and g38333 ( n16768 , n12270 , n2736 );
    xnor g38334 ( n5957 , n36998 , n7009 );
    or g38335 ( n29665 , n4717 , n1281 );
    and g38336 ( n21207 , n23549 , n11912 );
    xnor g38337 ( n35428 , n4712 , n41139 );
    nor g38338 ( n13909 , n13621 , n5417 );
    not g38339 ( n20222 , n21915 );
    and g38340 ( n3919 , n6007 , n20281 );
    not g38341 ( n32476 , n18915 );
    not g38342 ( n14219 , n25067 );
    or g38343 ( n5958 , n11374 , n431 );
    not g38344 ( n19571 , n13234 );
    and g38345 ( n9912 , n7022 , n34556 );
    or g38346 ( n36339 , n38653 , n1354 );
    or g38347 ( n32380 , n36856 , n5613 );
    and g38348 ( n5386 , n28384 , n37023 );
    and g38349 ( n33029 , n41398 , n39492 );
    or g38350 ( n17366 , n23801 , n6004 );
    or g38351 ( n21587 , n11067 , n2612 );
    xnor g38352 ( n29971 , n20323 , n14853 );
    nor g38353 ( n28740 , n41534 , n30266 );
    and g38354 ( n15691 , n13908 , n19323 );
    not g38355 ( n19030 , n8121 );
    xnor g38356 ( n41056 , n29611 , n1918 );
    or g38357 ( n6579 , n15239 , n22532 );
    or g38358 ( n19732 , n37869 , n27912 );
    and g38359 ( n6811 , n37810 , n19373 );
    xnor g38360 ( n14476 , n8439 , n40077 );
    and g38361 ( n4449 , n11846 , n4320 );
    or g38362 ( n24672 , n40884 , n25285 );
    nor g38363 ( n40904 , n25588 , n42537 );
    or g38364 ( n29748 , n25273 , n9423 );
    not g38365 ( n14723 , n5915 );
    nor g38366 ( n8313 , n38879 , n23924 );
    xnor g38367 ( n25707 , n38785 , n6789 );
    nor g38368 ( n34542 , n26018 , n40267 );
    and g38369 ( n23065 , n20291 , n35107 );
    and g38370 ( n31605 , n12303 , n89 );
    and g38371 ( n3855 , n22283 , n42635 );
    not g38372 ( n31691 , n28192 );
    and g38373 ( n16995 , n13850 , n19713 );
    not g38374 ( n27861 , n38153 );
    and g38375 ( n32151 , n8607 , n8030 );
    or g38376 ( n34519 , n39483 , n39980 );
    or g38377 ( n17749 , n31382 , n27629 );
    and g38378 ( n254 , n19053 , n574 );
    xnor g38379 ( n6634 , n25619 , n36494 );
    not g38380 ( n6978 , n7999 );
    xnor g38381 ( n39652 , n24980 , n32441 );
    or g38382 ( n9363 , n3255 , n18319 );
    or g38383 ( n20951 , n28221 , n11960 );
    or g38384 ( n23108 , n23690 , n40132 );
    not g38385 ( n17903 , n12822 );
    and g38386 ( n22167 , n155 , n34966 );
    and g38387 ( n13713 , n28219 , n24145 );
    not g38388 ( n19052 , n38828 );
    or g38389 ( n11627 , n21774 , n19242 );
    not g38390 ( n32018 , n1123 );
    or g38391 ( n32122 , n11340 , n2813 );
    and g38392 ( n41401 , n37166 , n10389 );
    and g38393 ( n4689 , n32412 , n41232 );
    and g38394 ( n35719 , n27811 , n36594 );
    or g38395 ( n20769 , n6430 , n1090 );
    or g38396 ( n15464 , n41186 , n14395 );
    and g38397 ( n3630 , n4111 , n36085 );
    or g38398 ( n671 , n21683 , n21860 );
    or g38399 ( n35620 , n41462 , n3645 );
    or g38400 ( n34524 , n22821 , n19664 );
    xnor g38401 ( n41994 , n34731 , n35180 );
    or g38402 ( n40045 , n36381 , n21363 );
    not g38403 ( n23322 , n6984 );
    or g38404 ( n11030 , n40588 , n17556 );
    or g38405 ( n11096 , n5232 , n18992 );
    and g38406 ( n35736 , n17905 , n42727 );
    or g38407 ( n22347 , n14735 , n2847 );
    or g38408 ( n21113 , n23041 , n9479 );
    and g38409 ( n41449 , n36998 , n21057 );
    and g38410 ( n42394 , n41508 , n578 );
    not g38411 ( n41357 , n32119 );
    xnor g38412 ( n18350 , n13444 , n17410 );
    and g38413 ( n29217 , n4137 , n3297 );
    xnor g38414 ( n30514 , n26898 , n12462 );
    or g38415 ( n32621 , n15823 , n13642 );
    and g38416 ( n23047 , n875 , n29993 );
    not g38417 ( n40600 , n24716 );
    nor g38418 ( n27974 , n17712 , n33852 );
    nor g38419 ( n8470 , n25588 , n13384 );
    xnor g38420 ( n3861 , n566 , n32 );
    or g38421 ( n15634 , n4266 , n9357 );
    and g38422 ( n4564 , n8889 , n838 );
    or g38423 ( n22661 , n7058 , n6086 );
    not g38424 ( n37057 , n9678 );
    not g38425 ( n15752 , n19367 );
    nor g38426 ( n35726 , n18520 , n25579 );
    and g38427 ( n23183 , n8366 , n17465 );
    or g38428 ( n33816 , n32549 , n2034 );
    or g38429 ( n6449 , n3237 , n24836 );
    and g38430 ( n40878 , n31637 , n12085 );
    or g38431 ( n10085 , n29822 , n33828 );
    and g38432 ( n20367 , n37172 , n28826 );
    and g38433 ( n33724 , n23927 , n34364 );
    or g38434 ( n18109 , n12847 , n38266 );
    and g38435 ( n7012 , n19150 , n12451 );
    or g38436 ( n36170 , n40591 , n22007 );
    not g38437 ( n14185 , n16066 );
    and g38438 ( n13021 , n4888 , n35396 );
    and g38439 ( n23738 , n40813 , n3043 );
    or g38440 ( n9019 , n5116 , n24812 );
    and g38441 ( n4893 , n21497 , n16722 );
    and g38442 ( n25335 , n31187 , n18240 );
    or g38443 ( n31524 , n15264 , n29545 );
    or g38444 ( n12604 , n35625 , n1479 );
    and g38445 ( n16129 , n30927 , n33933 );
    xnor g38446 ( n35233 , n8836 , n22860 );
    nor g38447 ( n14612 , n18145 , n33299 );
    or g38448 ( n34302 , n28212 , n17474 );
    or g38449 ( n22655 , n40110 , n7285 );
    nor g38450 ( n18106 , n30590 , n38942 );
    or g38451 ( n21086 , n15070 , n33304 );
    or g38452 ( n14123 , n30881 , n1378 );
    nor g38453 ( n22976 , n9422 , n8423 );
    nor g38454 ( n38976 , n39330 , n14800 );
    nor g38455 ( n27312 , n14530 , n13730 );
    xnor g38456 ( n26525 , n22879 , n7483 );
    and g38457 ( n291 , n24620 , n30891 );
    not g38458 ( n39870 , n24956 );
    and g38459 ( n3402 , n9073 , n40727 );
    or g38460 ( n6847 , n6215 , n1510 );
    not g38461 ( n16746 , n7673 );
    or g38462 ( n2821 , n6632 , n1940 );
    or g38463 ( n20528 , n550 , n34638 );
    and g38464 ( n33535 , n18059 , n4944 );
    or g38465 ( n13463 , n37978 , n1387 );
    xnor g38466 ( n39246 , n105 , n27211 );
    and g38467 ( n32112 , n25744 , n18720 );
    or g38468 ( n29820 , n23102 , n19848 );
    and g38469 ( n35364 , n14329 , n33126 );
    not g38470 ( n40295 , n9005 );
    or g38471 ( n40734 , n13741 , n32146 );
    or g38472 ( n28099 , n19130 , n27526 );
    or g38473 ( n5338 , n19969 , n15999 );
    or g38474 ( n24201 , n25109 , n13368 );
    not g38475 ( n26572 , n2689 );
    and g38476 ( n9162 , n35008 , n10321 );
    or g38477 ( n32077 , n37177 , n34569 );
    xnor g38478 ( n29634 , n33511 , n2968 );
    or g38479 ( n10096 , n25583 , n946 );
    or g38480 ( n5394 , n26542 , n7635 );
    nor g38481 ( n5829 , n25588 , n21538 );
    or g38482 ( n40208 , n6526 , n5007 );
    nor g38483 ( n16178 , n31746 , n3671 );
    xnor g38484 ( n5981 , n40781 , n32156 );
    and g38485 ( n5291 , n41001 , n7868 );
    and g38486 ( n29111 , n9897 , n33668 );
    xnor g38487 ( n20220 , n15281 , n26731 );
    nor g38488 ( n40073 , n1617 , n8593 );
    and g38489 ( n8703 , n21892 , n26390 );
    or g38490 ( n5817 , n27439 , n4747 );
    and g38491 ( n11 , n24964 , n4714 );
    and g38492 ( n16563 , n199 , n22665 );
    not g38493 ( n3891 , n12076 );
    or g38494 ( n1561 , n6229 , n3246 );
    or g38495 ( n7089 , n9750 , n6842 );
    and g38496 ( n31070 , n37356 , n5231 );
    or g38497 ( n11540 , n40955 , n26215 );
    xnor g38498 ( n22642 , n27767 , n37642 );
    xnor g38499 ( n26891 , n41900 , n14444 );
    or g38500 ( n39734 , n6636 , n20581 );
    not g38501 ( n41564 , n33891 );
    or g38502 ( n31714 , n39050 , n28408 );
    and g38503 ( n30790 , n5909 , n7739 );
    or g38504 ( n38086 , n14455 , n29035 );
    not g38505 ( n38752 , n41117 );
    or g38506 ( n40162 , n748 , n42870 );
    or g38507 ( n3831 , n18387 , n23094 );
    xnor g38508 ( n34471 , n41013 , n26982 );
    or g38509 ( n21022 , n7670 , n13478 );
    or g38510 ( n12662 , n76 , n7021 );
    xnor g38511 ( n38577 , n2839 , n704 );
    or g38512 ( n3205 , n28430 , n4717 );
    or g38513 ( n37157 , n30118 , n33262 );
    or g38514 ( n7182 , n12705 , n12891 );
    or g38515 ( n5275 , n1370 , n42726 );
    and g38516 ( n10241 , n14183 , n28412 );
    not g38517 ( n19519 , n8759 );
    and g38518 ( n12967 , n15779 , n9366 );
    and g38519 ( n8009 , n3608 , n27391 );
    and g38520 ( n38815 , n8996 , n34937 );
    or g38521 ( n2168 , n33815 , n3874 );
    not g38522 ( n21738 , n31909 );
    and g38523 ( n26994 , n35827 , n2981 );
    nor g38524 ( n34316 , n33508 , n8780 );
    not g38525 ( n33160 , n32722 );
    not g38526 ( n18257 , n41959 );
    not g38527 ( n4558 , n23170 );
    nor g38528 ( n19438 , n41563 , n41791 );
    xnor g38529 ( n8850 , n23304 , n38729 );
    and g38530 ( n15387 , n35172 , n19981 );
    xnor g38531 ( n6933 , n9810 , n18307 );
    or g38532 ( n29133 , n30875 , n6316 );
    or g38533 ( n22798 , n24356 , n9162 );
    xnor g38534 ( n24175 , n28333 , n4436 );
    or g38535 ( n4945 , n2916 , n2689 );
    not g38536 ( n13084 , n4151 );
    or g38537 ( n20356 , n3893 , n34199 );
    or g38538 ( n28203 , n31691 , n17203 );
    or g38539 ( n27617 , n4305 , n40539 );
    and g38540 ( n10892 , n23231 , n41106 );
    or g38541 ( n25232 , n17001 , n21528 );
    xnor g38542 ( n19213 , n24159 , n22666 );
    and g38543 ( n863 , n1041 , n37746 );
    or g38544 ( n23532 , n31303 , n39536 );
    or g38545 ( n8705 , n27926 , n28065 );
    xnor g38546 ( n7661 , n4334 , n38120 );
    or g38547 ( n31788 , n6411 , n19497 );
    not g38548 ( n12318 , n7681 );
    or g38549 ( n34327 , n41961 , n39379 );
    xnor g38550 ( n34178 , n2659 , n7742 );
    xnor g38551 ( n13023 , n2632 , n25329 );
    xnor g38552 ( n7695 , n298 , n29602 );
    not g38553 ( n30826 , n42497 );
    nor g38554 ( n21292 , n3369 , n15108 );
    nor g38555 ( n28522 , n8660 , n28172 );
    xnor g38556 ( n11289 , n22263 , n27669 );
    or g38557 ( n16038 , n32939 , n28859 );
    not g38558 ( n5904 , n13668 );
    xnor g38559 ( n13386 , n39645 , n18279 );
    or g38560 ( n22364 , n15449 , n11828 );
    and g38561 ( n16941 , n6318 , n30353 );
    nor g38562 ( n1360 , n9674 , n36750 );
    not g38563 ( n21954 , n26268 );
    or g38564 ( n29581 , n20699 , n42882 );
    nor g38565 ( n9910 , n4949 , n13170 );
    not g38566 ( n8857 , n17234 );
    or g38567 ( n26612 , n991 , n13989 );
    or g38568 ( n31023 , n3311 , n33223 );
    nor g38569 ( n19167 , n37025 , n3344 );
    and g38570 ( n20722 , n18674 , n33065 );
    xnor g38571 ( n18926 , n19628 , n29870 );
    xnor g38572 ( n2651 , n29740 , n37843 );
    or g38573 ( n12793 , n5475 , n316 );
    or g38574 ( n37741 , n30479 , n37035 );
    or g38575 ( n32500 , n24264 , n38061 );
    nor g38576 ( n13923 , n9421 , n33425 );
    or g38577 ( n32765 , n37212 , n10087 );
    and g38578 ( n5434 , n42663 , n24494 );
    not g38579 ( n26786 , n15756 );
    xnor g38580 ( n41634 , n35727 , n30767 );
    nor g38581 ( n26384 , n31857 , n2542 );
    and g38582 ( n22548 , n2952 , n7249 );
    and g38583 ( n32518 , n6422 , n15901 );
    or g38584 ( n5405 , n1994 , n12679 );
    not g38585 ( n23411 , n21488 );
    and g38586 ( n805 , n5971 , n7791 );
    not g38587 ( n9142 , n20553 );
    not g38588 ( n30820 , n15439 );
    nor g38589 ( n39317 , n9568 , n1108 );
    or g38590 ( n20869 , n8707 , n5910 );
    and g38591 ( n16416 , n35906 , n35060 );
    not g38592 ( n28080 , n39226 );
    or g38593 ( n28893 , n4670 , n14814 );
    or g38594 ( n22228 , n8128 , n17763 );
    or g38595 ( n34101 , n5844 , n36848 );
    nor g38596 ( n7772 , n14471 , n12601 );
    or g38597 ( n40866 , n674 , n21662 );
    or g38598 ( n11937 , n8996 , n34937 );
    or g38599 ( n20692 , n24729 , n9790 );
    nor g38600 ( n12738 , n21652 , n2992 );
    or g38601 ( n2736 , n34960 , n33304 );
    nor g38602 ( n36887 , n14471 , n31049 );
    or g38603 ( n36588 , n24453 , n35304 );
    nor g38604 ( n21224 , n3343 , n23960 );
    or g38605 ( n33000 , n22294 , n34118 );
    or g38606 ( n6518 , n7996 , n23740 );
    or g38607 ( n3085 , n42327 , n11504 );
    or g38608 ( n38275 , n20324 , n26879 );
    or g38609 ( n6384 , n37886 , n24330 );
    or g38610 ( n4362 , n18895 , n2095 );
    or g38611 ( n38277 , n37152 , n29735 );
    not g38612 ( n6841 , n35759 );
    and g38613 ( n11775 , n11608 , n40410 );
    and g38614 ( n16001 , n7407 , n2257 );
    or g38615 ( n28429 , n1716 , n39839 );
    and g38616 ( n32332 , n21247 , n3173 );
    and g38617 ( n18879 , n2027 , n35885 );
    xnor g38618 ( n37418 , n7641 , n34823 );
    or g38619 ( n37696 , n20681 , n12525 );
    or g38620 ( n20195 , n33704 , n18087 );
    and g38621 ( n27510 , n7936 , n38737 );
    nor g38622 ( n30566 , n27762 , n27194 );
    or g38623 ( n33684 , n14252 , n22977 );
    xnor g38624 ( n16138 , n21592 , n20687 );
    xnor g38625 ( n18892 , n21141 , n29653 );
    or g38626 ( n24725 , n30371 , n15317 );
    nor g38627 ( n8199 , n1011 , n42874 );
    xnor g38628 ( n10797 , n17647 , n29234 );
    and g38629 ( n12718 , n39315 , n37537 );
    nor g38630 ( n16837 , n21347 , n20521 );
    not g38631 ( n20884 , n33451 );
    and g38632 ( n24910 , n27650 , n9374 );
    nor g38633 ( n19918 , n18754 , n32658 );
    or g38634 ( n324 , n17193 , n11821 );
    xnor g38635 ( n12521 , n11436 , n88 );
    nor g38636 ( n8691 , n35665 , n25412 );
    or g38637 ( n19633 , n33549 , n14487 );
    not g38638 ( n36104 , n28821 );
    or g38639 ( n22890 , n21836 , n28440 );
    and g38640 ( n26298 , n25153 , n30950 );
    or g38641 ( n42526 , n34549 , n36087 );
    or g38642 ( n10794 , n32786 , n16362 );
    and g38643 ( n9068 , n37372 , n15811 );
    xnor g38644 ( n39490 , n6884 , n24225 );
    or g38645 ( n22140 , n25047 , n17686 );
    nor g38646 ( n5577 , n16866 , n40732 );
    xnor g38647 ( n40875 , n25619 , n33946 );
    or g38648 ( n15297 , n7356 , n30031 );
    or g38649 ( n19851 , n16109 , n20594 );
    or g38650 ( n31673 , n37076 , n33307 );
    or g38651 ( n42149 , n34751 , n15735 );
    or g38652 ( n30209 , n11327 , n24075 );
    or g38653 ( n9811 , n31485 , n42812 );
    nor g38654 ( n19331 , n11531 , n24143 );
    or g38655 ( n32184 , n24824 , n34293 );
    not g38656 ( n26515 , n28949 );
    and g38657 ( n12306 , n16922 , n7353 );
    or g38658 ( n9598 , n6138 , n40080 );
    or g38659 ( n14727 , n34994 , n18485 );
    not g38660 ( n15220 , n20068 );
    and g38661 ( n4675 , n9768 , n14555 );
    nor g38662 ( n19565 , n38342 , n1836 );
    or g38663 ( n33999 , n33394 , n950 );
    and g38664 ( n15278 , n25629 , n4038 );
    or g38665 ( n5550 , n27128 , n16724 );
    or g38666 ( n41919 , n19873 , n2415 );
    nor g38667 ( n25352 , n34565 , n20825 );
    or g38668 ( n10931 , n10205 , n31769 );
    not g38669 ( n10707 , n9874 );
    and g38670 ( n31258 , n1779 , n20933 );
    and g38671 ( n12234 , n31328 , n28367 );
    xnor g38672 ( n2261 , n7489 , n42288 );
    or g38673 ( n20518 , n12890 , n21558 );
    and g38674 ( n30269 , n19285 , n10514 );
    not g38675 ( n11531 , n3539 );
    or g38676 ( n19018 , n9809 , n19773 );
    or g38677 ( n12165 , n31707 , n19560 );
    or g38678 ( n10046 , n16013 , n42533 );
    or g38679 ( n6096 , n16109 , n37484 );
    and g38680 ( n36659 , n38079 , n2860 );
    or g38681 ( n35535 , n15224 , n8586 );
    not g38682 ( n28407 , n27766 );
    and g38683 ( n28969 , n20605 , n3510 );
    not g38684 ( n317 , n30570 );
    or g38685 ( n40667 , n19976 , n21981 );
    or g38686 ( n9973 , n42638 , n10953 );
    and g38687 ( n21673 , n27852 , n27346 );
    and g38688 ( n37229 , n15549 , n29921 );
    not g38689 ( n7004 , n5940 );
    or g38690 ( n26013 , n35001 , n3954 );
    or g38691 ( n40003 , n24666 , n7070 );
    or g38692 ( n11562 , n28364 , n15421 );
    or g38693 ( n26055 , n37107 , n21019 );
    not g38694 ( n735 , n5873 );
    and g38695 ( n4929 , n28240 , n29617 );
    not g38696 ( n17229 , n14888 );
    and g38697 ( n37064 , n9493 , n10227 );
    nor g38698 ( n32315 , n29098 , n22884 );
    nor g38699 ( n27518 , n941 , n2724 );
    not g38700 ( n32261 , n3930 );
    nor g38701 ( n37440 , n23914 , n20290 );
    xnor g38702 ( n25259 , n30943 , n35119 );
    or g38703 ( n34656 , n41000 , n25221 );
    or g38704 ( n38148 , n11417 , n38786 );
    not g38705 ( n4266 , n38486 );
    or g38706 ( n19956 , n42683 , n25626 );
    or g38707 ( n37291 , n7174 , n26580 );
    and g38708 ( n32309 , n18633 , n19195 );
    xnor g38709 ( n17676 , n40191 , n22018 );
    and g38710 ( n22186 , n16518 , n40628 );
    and g38711 ( n26765 , n1691 , n18614 );
    or g38712 ( n3512 , n691 , n33621 );
    or g38713 ( n29877 , n19311 , n17502 );
    not g38714 ( n33434 , n24378 );
    or g38715 ( n1330 , n41548 , n4715 );
    not g38716 ( n27465 , n14563 );
    or g38717 ( n6038 , n18685 , n14177 );
    nor g38718 ( n9567 , n32916 , n36969 );
    and g38719 ( n8998 , n35709 , n2574 );
    and g38720 ( n14699 , n33882 , n42261 );
    not g38721 ( n31866 , n41148 );
    and g38722 ( n29707 , n25842 , n23939 );
    and g38723 ( n10208 , n19021 , n2874 );
    not g38724 ( n14668 , n40635 );
    or g38725 ( n1420 , n2947 , n715 );
    nor g38726 ( n3220 , n16475 , n11649 );
    xnor g38727 ( n8250 , n13683 , n36205 );
    or g38728 ( n40569 , n19446 , n19104 );
    not g38729 ( n24943 , n10962 );
    or g38730 ( n11994 , n5194 , n39772 );
    or g38731 ( n13295 , n14383 , n27165 );
    not g38732 ( n3531 , n5515 );
    and g38733 ( n42369 , n14058 , n31022 );
    nor g38734 ( n10648 , n34052 , n8042 );
    and g38735 ( n5057 , n21741 , n21262 );
    xnor g38736 ( n41248 , n35727 , n25969 );
    xnor g38737 ( n9778 , n7342 , n12975 );
    or g38738 ( n38838 , n8004 , n9704 );
    nor g38739 ( n42486 , n14821 , n34636 );
    not g38740 ( n23689 , n39158 );
    xnor g38741 ( n14469 , n28867 , n14138 );
    nor g38742 ( n22867 , n7554 , n7431 );
    or g38743 ( n18922 , n39708 , n36644 );
    or g38744 ( n23799 , n4460 , n29316 );
    or g38745 ( n17103 , n19850 , n17364 );
    nor g38746 ( n4451 , n40550 , n13333 );
    not g38747 ( n7299 , n40511 );
    or g38748 ( n6034 , n26689 , n23396 );
    and g38749 ( n37292 , n28285 , n37226 );
    or g38750 ( n35962 , n19126 , n36447 );
    xnor g38751 ( n30227 , n28541 , n34128 );
    not g38752 ( n41323 , n387 );
    or g38753 ( n16867 , n14030 , n17623 );
    or g38754 ( n20419 , n19110 , n14057 );
    and g38755 ( n6118 , n27853 , n8118 );
    or g38756 ( n11397 , n40375 , n8911 );
    and g38757 ( n5265 , n1547 , n459 );
    xnor g38758 ( n25800 , n23867 , n7765 );
    nor g38759 ( n42753 , n16640 , n34989 );
    not g38760 ( n10377 , n33707 );
    and g38761 ( n40669 , n21463 , n320 );
    or g38762 ( n351 , n19455 , n18072 );
    or g38763 ( n5418 , n31728 , n37711 );
    xnor g38764 ( n24700 , n35361 , n25298 );
    not g38765 ( n1631 , n26332 );
    not g38766 ( n39475 , n39537 );
    nor g38767 ( n6708 , n4140 , n31339 );
    and g38768 ( n37185 , n29855 , n38380 );
    nor g38769 ( n33411 , n16410 , n28416 );
    or g38770 ( n36990 , n5063 , n12788 );
    and g38771 ( n15719 , n17619 , n5972 );
    or g38772 ( n36766 , n13414 , n41160 );
    or g38773 ( n38005 , n40694 , n35094 );
    or g38774 ( n40190 , n24054 , n36473 );
    or g38775 ( n30267 , n40713 , n308 );
    or g38776 ( n14369 , n16761 , n22016 );
    nor g38777 ( n38855 , n14707 , n35160 );
    nor g38778 ( n41624 , n9448 , n29829 );
    nor g38779 ( n17700 , n1110 , n34194 );
    not g38780 ( n19485 , n35025 );
    not g38781 ( n492 , n39253 );
    nor g38782 ( n4405 , n38946 , n19921 );
    or g38783 ( n38775 , n7903 , n38418 );
    not g38784 ( n21652 , n32558 );
    or g38785 ( n1184 , n40899 , n3969 );
    or g38786 ( n23410 , n3544 , n4533 );
    or g38787 ( n10317 , n3583 , n11971 );
    or g38788 ( n31488 , n40339 , n5813 );
    xnor g38789 ( n33937 , n6625 , n27709 );
    or g38790 ( n39369 , n17626 , n6912 );
    not g38791 ( n3226 , n34306 );
    and g38792 ( n22078 , n28581 , n30246 );
    or g38793 ( n6100 , n4070 , n4841 );
    not g38794 ( n21025 , n5993 );
    xnor g38795 ( n13831 , n7836 , n9727 );
    or g38796 ( n29961 , n11707 , n21533 );
    or g38797 ( n5383 , n1183 , n8682 );
    xnor g38798 ( n42146 , n784 , n930 );
    or g38799 ( n40158 , n18166 , n36815 );
    or g38800 ( n33600 , n755 , n29803 );
    or g38801 ( n20541 , n31195 , n2565 );
    and g38802 ( n18156 , n27310 , n41643 );
    or g38803 ( n35229 , n1767 , n35970 );
    nor g38804 ( n1649 , n24636 , n31259 );
    and g38805 ( n1415 , n42563 , n17688 );
    not g38806 ( n6517 , n25977 );
    or g38807 ( n10227 , n11601 , n37279 );
    or g38808 ( n26751 , n36641 , n32975 );
    and g38809 ( n21275 , n20211 , n18369 );
    nor g38810 ( n35804 , n10617 , n7659 );
    or g38811 ( n3375 , n9084 , n33228 );
    and g38812 ( n2511 , n16653 , n20812 );
    and g38813 ( n26171 , n18991 , n30375 );
    not g38814 ( n29939 , n25670 );
    nor g38815 ( n35002 , n37539 , n10718 );
    or g38816 ( n15680 , n36585 , n39093 );
    not g38817 ( n20503 , n294 );
    or g38818 ( n5024 , n31542 , n19737 );
    and g38819 ( n38795 , n13091 , n8007 );
    nor g38820 ( n40973 , n96 , n12478 );
    or g38821 ( n28798 , n12656 , n42824 );
    or g38822 ( n38114 , n19169 , n28123 );
    xnor g38823 ( n8653 , n15522 , n3004 );
    or g38824 ( n31659 , n37365 , n31503 );
    or g38825 ( n38823 , n3217 , n16724 );
    or g38826 ( n24996 , n34081 , n10953 );
    nor g38827 ( n22069 , n5896 , n39612 );
    and g38828 ( n13421 , n3188 , n16689 );
    and g38829 ( n33709 , n37838 , n40217 );
    nor g38830 ( n3803 , n42792 , n27372 );
    not g38831 ( n33892 , n21997 );
    not g38832 ( n34891 , n23357 );
    not g38833 ( n2632 , n37873 );
    not g38834 ( n15556 , n354 );
    not g38835 ( n36071 , n35604 );
    or g38836 ( n3841 , n18438 , n28055 );
    or g38837 ( n4167 , n20030 , n39155 );
    and g38838 ( n16054 , n1517 , n38188 );
    or g38839 ( n34868 , n5348 , n30471 );
    or g38840 ( n16958 , n32256 , n2694 );
    nor g38841 ( n39779 , n24149 , n39319 );
    and g38842 ( n39037 , n12799 , n8792 );
    not g38843 ( n27137 , n15356 );
    or g38844 ( n34808 , n34569 , n12995 );
    not g38845 ( n13437 , n8655 );
    and g38846 ( n25814 , n34460 , n17349 );
    xnor g38847 ( n14347 , n21534 , n28547 );
    nor g38848 ( n34570 , n12837 , n6837 );
    or g38849 ( n5990 , n29169 , n12137 );
    not g38850 ( n22371 , n15778 );
    not g38851 ( n36161 , n35890 );
    xnor g38852 ( n24078 , n13313 , n2199 );
    or g38853 ( n16212 , n9673 , n27549 );
    or g38854 ( n23308 , n34082 , n7316 );
    or g38855 ( n31246 , n19584 , n26563 );
    or g38856 ( n37617 , n40302 , n41413 );
    or g38857 ( n14046 , n34760 , n40626 );
    xnor g38858 ( n28436 , n12389 , n30620 );
    nor g38859 ( n36396 , n13249 , n9043 );
    not g38860 ( n29799 , n3680 );
    or g38861 ( n16484 , n16272 , n8712 );
    or g38862 ( n37449 , n9915 , n39194 );
    or g38863 ( n23350 , n30235 , n25000 );
    xnor g38864 ( n41133 , n5457 , n13314 );
    not g38865 ( n19049 , n19620 );
    and g38866 ( n21852 , n18754 , n32658 );
    not g38867 ( n38975 , n40140 );
    and g38868 ( n32879 , n41195 , n19263 );
    or g38869 ( n13956 , n41961 , n5181 );
    or g38870 ( n6441 , n10633 , n41879 );
    not g38871 ( n36286 , n9599 );
    or g38872 ( n847 , n27091 , n39536 );
    and g38873 ( n30447 , n34846 , n36018 );
    or g38874 ( n9386 , n28846 , n27743 );
    not g38875 ( n18963 , n17821 );
    nor g38876 ( n19069 , n40163 , n35432 );
    or g38877 ( n24891 , n16158 , n36445 );
    or g38878 ( n17033 , n7900 , n22991 );
    xnor g38879 ( n34139 , n24067 , n34668 );
    xnor g38880 ( n1371 , n22128 , n17340 );
    or g38881 ( n6961 , n545 , n27392 );
    or g38882 ( n39076 , n41288 , n16678 );
    or g38883 ( n24320 , n12100 , n20684 );
    not g38884 ( n9800 , n41202 );
    not g38885 ( n42054 , n21871 );
    and g38886 ( n34797 , n10721 , n38003 );
    nor g38887 ( n37586 , n10881 , n27575 );
    nor g38888 ( n41160 , n27524 , n40304 );
    xnor g38889 ( n91 , n18530 , n14726 );
    and g38890 ( n5610 , n13073 , n34848 );
    or g38891 ( n30033 , n14854 , n7347 );
    and g38892 ( n25743 , n8310 , n32616 );
    not g38893 ( n41182 , n19897 );
    and g38894 ( n3480 , n9672 , n26544 );
    and g38895 ( n3029 , n35727 , n12746 );
    or g38896 ( n19530 , n9519 , n30278 );
    nor g38897 ( n8681 , n9020 , n15370 );
    xnor g38898 ( n3336 , n105 , n34133 );
    nor g38899 ( n15451 , n13593 , n17414 );
    and g38900 ( n36084 , n39591 , n4636 );
    or g38901 ( n15209 , n1971 , n34248 );
    or g38902 ( n8388 , n19922 , n9456 );
    and g38903 ( n12910 , n7817 , n2196 );
    or g38904 ( n15966 , n32302 , n1734 );
    and g38905 ( n18978 , n29398 , n14588 );
    and g38906 ( n11052 , n24529 , n38212 );
    nor g38907 ( n27202 , n23971 , n17134 );
    xnor g38908 ( n3634 , n4340 , n24635 );
    xnor g38909 ( n26103 , n2921 , n40126 );
    nor g38910 ( n14897 , n30237 , n35848 );
    nor g38911 ( n10670 , n17551 , n18008 );
    or g38912 ( n10957 , n36099 , n24061 );
    not g38913 ( n15006 , n15589 );
    xnor g38914 ( n19132 , n22670 , n39266 );
    not g38915 ( n24510 , n13054 );
    or g38916 ( n40060 , n27873 , n20632 );
    or g38917 ( n39504 , n41425 , n32180 );
    or g38918 ( n37766 , n38461 , n21942 );
    xnor g38919 ( n23470 , n31460 , n27480 );
    not g38920 ( n26147 , n28662 );
    and g38921 ( n21950 , n30161 , n3805 );
    xnor g38922 ( n41536 , n34602 , n22390 );
    and g38923 ( n30777 , n20339 , n3197 );
    and g38924 ( n2876 , n29465 , n568 );
    or g38925 ( n15326 , n22734 , n21510 );
    or g38926 ( n34713 , n23942 , n33955 );
    or g38927 ( n27695 , n37131 , n39973 );
    not g38928 ( n6415 , n2535 );
    or g38929 ( n5627 , n23777 , n14095 );
    or g38930 ( n35551 , n6503 , n29955 );
    nor g38931 ( n18663 , n24209 , n26833 );
    or g38932 ( n29463 , n31997 , n28539 );
    or g38933 ( n26195 , n20587 , n6042 );
    nor g38934 ( n5100 , n23431 , n37360 );
    xnor g38935 ( n32388 , n1917 , n35990 );
    or g38936 ( n12609 , n31030 , n30822 );
    and g38937 ( n19631 , n23477 , n35305 );
    not g38938 ( n39213 , n112 );
    or g38939 ( n20022 , n12286 , n29998 );
    and g38940 ( n25200 , n22245 , n13253 );
    nor g38941 ( n35697 , n33258 , n40034 );
    xnor g38942 ( n19718 , n25619 , n1993 );
    or g38943 ( n3944 , n14112 , n6212 );
    or g38944 ( n4770 , n34391 , n36875 );
    nor g38945 ( n14341 , n32461 , n10003 );
    or g38946 ( n17939 , n27357 , n28690 );
    and g38947 ( n40807 , n30604 , n305 );
    not g38948 ( n23893 , n40227 );
    and g38949 ( n9928 , n4252 , n1331 );
    xnor g38950 ( n16811 , n1762 , n29788 );
    or g38951 ( n41617 , n3506 , n24496 );
    or g38952 ( n34196 , n39233 , n22631 );
    and g38953 ( n13178 , n10114 , n31416 );
    or g38954 ( n20739 , n2146 , n25666 );
    nor g38955 ( n2044 , n8694 , n12449 );
    or g38956 ( n14719 , n19221 , n22543 );
    and g38957 ( n40930 , n18270 , n10615 );
    nor g38958 ( n32355 , n14707 , n25803 );
    or g38959 ( n41070 , n19673 , n17847 );
    xnor g38960 ( n38267 , n6625 , n6126 );
    xnor g38961 ( n6175 , n39531 , n21337 );
    or g38962 ( n25441 , n5085 , n904 );
    xnor g38963 ( n40424 , n38668 , n19761 );
    or g38964 ( n29889 , n6629 , n36647 );
    not g38965 ( n25958 , n14778 );
    and g38966 ( n38456 , n15887 , n35003 );
    nor g38967 ( n25824 , n6762 , n6859 );
    xnor g38968 ( n13484 , n12146 , n31101 );
    xnor g38969 ( n20648 , n1011 , n37862 );
    or g38970 ( n11017 , n22732 , n27631 );
    not g38971 ( n38650 , n18719 );
    not g38972 ( n22212 , n29394 );
    or g38973 ( n23961 , n22821 , n40504 );
    xnor g38974 ( n36759 , n31989 , n10515 );
    or g38975 ( n24970 , n9255 , n884 );
    and g38976 ( n5473 , n1157 , n16796 );
    or g38977 ( n664 , n34558 , n30131 );
    or g38978 ( n15538 , n5718 , n13923 );
    nor g38979 ( n1400 , n39191 , n27115 );
    nor g38980 ( n1322 , n38879 , n13199 );
    not g38981 ( n37819 , n6600 );
    or g38982 ( n23046 , n29849 , n28341 );
    and g38983 ( n30243 , n24166 , n25514 );
    not g38984 ( n33 , n33217 );
    nor g38985 ( n6208 , n32718 , n15071 );
    or g38986 ( n25171 , n9105 , n14902 );
    or g38987 ( n3612 , n94 , n15948 );
    xnor g38988 ( n15121 , n42071 , n20689 );
    xnor g38989 ( n42683 , n25075 , n17974 );
    or g38990 ( n20527 , n8674 , n2740 );
    nor g38991 ( n4606 , n5936 , n30787 );
    or g38992 ( n15741 , n40477 , n20921 );
    not g38993 ( n20167 , n38991 );
    or g38994 ( n26176 , n2419 , n4922 );
    xnor g38995 ( n24928 , n20310 , n18271 );
    not g38996 ( n15721 , n563 );
    or g38997 ( n31506 , n5893 , n521 );
    and g38998 ( n26197 , n17048 , n22930 );
    xnor g38999 ( n17668 , n42064 , n39502 );
    or g39000 ( n23215 , n24376 , n19845 );
    nor g39001 ( n11604 , n23275 , n27763 );
    and g39002 ( n33546 , n7563 , n31470 );
    and g39003 ( n39967 , n4663 , n17348 );
    or g39004 ( n37833 , n11356 , n19688 );
    or g39005 ( n42562 , n34997 , n1210 );
    not g39006 ( n21026 , n28042 );
    xnor g39007 ( n37239 , n31129 , n8494 );
    and g39008 ( n10857 , n41959 , n2189 );
    or g39009 ( n19155 , n25806 , n10002 );
    not g39010 ( n38806 , n6790 );
    xnor g39011 ( n24545 , n27644 , n36972 );
    not g39012 ( n1602 , n16357 );
    not g39013 ( n17494 , n1755 );
    not g39014 ( n6512 , n14233 );
    or g39015 ( n32413 , n32800 , n40853 );
    and g39016 ( n13294 , n35420 , n28936 );
    or g39017 ( n15 , n23457 , n14501 );
    or g39018 ( n38495 , n22548 , n20606 );
    nor g39019 ( n22287 , n23330 , n2303 );
    or g39020 ( n8321 , n29627 , n29884 );
    not g39021 ( n19984 , n9101 );
    or g39022 ( n23705 , n25356 , n19540 );
    not g39023 ( n23456 , n19118 );
    xnor g39024 ( n20397 , n15591 , n32133 );
    and g39025 ( n349 , n16601 , n12463 );
    not g39026 ( n6632 , n14224 );
    or g39027 ( n4993 , n36641 , n23314 );
    nor g39028 ( n920 , n9180 , n8892 );
    or g39029 ( n15465 , n40178 , n35131 );
    or g39030 ( n3187 , n14471 , n17398 );
    and g39031 ( n11253 , n31947 , n30632 );
    or g39032 ( n23469 , n12303 , n89 );
    not g39033 ( n27712 , n40954 );
    and g39034 ( n36101 , n12257 , n40198 );
    xnor g39035 ( n39349 , n5013 , n2410 );
    nor g39036 ( n37188 , n23162 , n11157 );
    or g39037 ( n20520 , n1952 , n34569 );
    xnor g39038 ( n13546 , n12146 , n27735 );
    or g39039 ( n13225 , n26227 , n26028 );
    and g39040 ( n34842 , n24346 , n2075 );
    nor g39041 ( n481 , n32475 , n19005 );
    or g39042 ( n14175 , n19990 , n36235 );
    or g39043 ( n18890 , n28774 , n42509 );
    or g39044 ( n20391 , n40845 , n16586 );
    xnor g39045 ( n9401 , n12024 , n35459 );
    and g39046 ( n9216 , n38742 , n16086 );
    xnor g39047 ( n2342 , n28185 , n9524 );
    nor g39048 ( n13686 , n14707 , n13980 );
    or g39049 ( n35763 , n35337 , n7901 );
    or g39050 ( n2122 , n40860 , n31940 );
    and g39051 ( n25779 , n20723 , n34607 );
    nor g39052 ( n10651 , n22170 , n15001 );
    or g39053 ( n39655 , n30072 , n1749 );
    not g39054 ( n19523 , n29987 );
    xnor g39055 ( n32201 , n1499 , n37043 );
    or g39056 ( n38206 , n1972 , n41207 );
    or g39057 ( n10238 , n26308 , n18075 );
    or g39058 ( n38682 , n18640 , n21725 );
    xnor g39059 ( n37765 , n6625 , n11734 );
    or g39060 ( n5306 , n29914 , n19434 );
    xnor g39061 ( n9777 , n22263 , n9920 );
    and g39062 ( n2418 , n195 , n12276 );
    and g39063 ( n10069 , n30330 , n41184 );
    and g39064 ( n659 , n6142 , n11479 );
    not g39065 ( n38695 , n10 );
    not g39066 ( n21301 , n31626 );
    and g39067 ( n13094 , n24428 , n36808 );
    not g39068 ( n21361 , n2604 );
    and g39069 ( n20796 , n14865 , n4997 );
    or g39070 ( n23912 , n10559 , n40983 );
    not g39071 ( n20383 , n20900 );
    or g39072 ( n10960 , n27208 , n7802 );
    and g39073 ( n33175 , n23608 , n16707 );
    xnor g39074 ( n42056 , n5891 , n28116 );
    or g39075 ( n29801 , n42340 , n41458 );
    or g39076 ( n1480 , n24780 , n41780 );
    and g39077 ( n20042 , n42010 , n18596 );
    or g39078 ( n38278 , n9809 , n26335 );
    xnor g39079 ( n33656 , n25118 , n8094 );
    xnor g39080 ( n21321 , n31099 , n42006 );
    nor g39081 ( n31221 , n14471 , n35192 );
    or g39082 ( n25293 , n25634 , n32112 );
    or g39083 ( n12237 , n6031 , n31055 );
    or g39084 ( n14189 , n30399 , n28273 );
    and g39085 ( n17681 , n33690 , n40992 );
    xnor g39086 ( n8812 , n5144 , n38213 );
    not g39087 ( n23239 , n9353 );
    not g39088 ( n29131 , n12578 );
    nor g39089 ( n4155 , n16598 , n38401 );
    or g39090 ( n17787 , n33239 , n37467 );
    or g39091 ( n14679 , n32741 , n16520 );
    nor g39092 ( n33924 , n10716 , n8864 );
    xnor g39093 ( n31620 , n20487 , n1870 );
    nor g39094 ( n37964 , n30862 , n5839 );
    not g39095 ( n23085 , n39226 );
    nor g39096 ( n41019 , n29640 , n1618 );
    or g39097 ( n34185 , n12907 , n30410 );
    or g39098 ( n21798 , n14411 , n8412 );
    nor g39099 ( n13880 , n22702 , n29171 );
    or g39100 ( n7533 , n8341 , n37247 );
    and g39101 ( n1865 , n41586 , n8249 );
    or g39102 ( n10089 , n28115 , n2148 );
    xnor g39103 ( n7502 , n2781 , n5896 );
    or g39104 ( n26246 , n18708 , n8722 );
    and g39105 ( n27545 , n27550 , n26143 );
    and g39106 ( n5532 , n41171 , n21468 );
    nor g39107 ( n32377 , n5826 , n14368 );
    xnor g39108 ( n6340 , n751 , n11661 );
    or g39109 ( n39863 , n36117 , n14557 );
    nor g39110 ( n40135 , n23123 , n11986 );
    or g39111 ( n14792 , n8442 , n16134 );
    not g39112 ( n40570 , n16781 );
    or g39113 ( n35392 , n35833 , n27102 );
    nor g39114 ( n38960 , n11130 , n15103 );
    or g39115 ( n3651 , n13885 , n2283 );
    or g39116 ( n21437 , n11374 , n35518 );
    or g39117 ( n11519 , n18741 , n15889 );
    or g39118 ( n7631 , n20071 , n31997 );
    not g39119 ( n2193 , n5696 );
    or g39120 ( n9925 , n141 , n19517 );
    and g39121 ( n24603 , n21637 , n27167 );
    or g39122 ( n11605 , n26342 , n19497 );
    and g39123 ( n8328 , n42353 , n19112 );
    xnor g39124 ( n23399 , n11846 , n4320 );
    or g39125 ( n30776 , n28718 , n20220 );
    nor g39126 ( n15553 , n17617 , n25342 );
    nor g39127 ( n36515 , n31394 , n36208 );
    or g39128 ( n40028 , n14622 , n17284 );
    or g39129 ( n9178 , n41006 , n13093 );
    or g39130 ( n38868 , n39213 , n5039 );
    not g39131 ( n7400 , n27638 );
    not g39132 ( n32226 , n31382 );
    and g39133 ( n16691 , n17255 , n19209 );
    nor g39134 ( n12194 , n40280 , n19949 );
    or g39135 ( n37242 , n7131 , n29932 );
    not g39136 ( n13820 , n30869 );
    not g39137 ( n20130 , n1420 );
    or g39138 ( n34894 , n16106 , n39825 );
    and g39139 ( n2836 , n32336 , n21008 );
    nor g39140 ( n37533 , n35301 , n4446 );
    xnor g39141 ( n1413 , n37709 , n3588 );
    or g39142 ( n30095 , n34499 , n8999 );
    and g39143 ( n30131 , n28110 , n39530 );
    not g39144 ( n29543 , n10617 );
    or g39145 ( n9529 , n11321 , n28434 );
    or g39146 ( n17497 , n41730 , n37740 );
    or g39147 ( n36018 , n18114 , n33289 );
    not g39148 ( n30896 , n35814 );
    and g39149 ( n16595 , n13444 , n40000 );
    and g39150 ( n35586 , n29917 , n10671 );
    or g39151 ( n1875 , n15776 , n41990 );
    and g39152 ( n30797 , n35727 , n25708 );
    or g39153 ( n12544 , n7628 , n10278 );
    and g39154 ( n39807 , n27141 , n12 );
    or g39155 ( n28011 , n6403 , n313 );
    not g39156 ( n31128 , n32056 );
    and g39157 ( n37353 , n15835 , n30106 );
    and g39158 ( n42207 , n40264 , n34771 );
    and g39159 ( n1256 , n2441 , n42474 );
    nor g39160 ( n39805 , n2263 , n27121 );
    and g39161 ( n37028 , n14979 , n29190 );
    not g39162 ( n39178 , n38828 );
    not g39163 ( n34569 , n3084 );
    nor g39164 ( n37053 , n15261 , n410 );
    xnor g39165 ( n17867 , n27596 , n19893 );
    nor g39166 ( n11653 , n41616 , n42746 );
    or g39167 ( n11889 , n33767 , n12715 );
    or g39168 ( n41929 , n9508 , n34430 );
    not g39169 ( n16510 , n42636 );
    not g39170 ( n18335 , n30902 );
    nor g39171 ( n26524 , n22049 , n7620 );
    nor g39172 ( n31501 , n25088 , n21790 );
    or g39173 ( n25558 , n1074 , n34225 );
    or g39174 ( n5739 , n26092 , n29504 );
    nor g39175 ( n30756 , n23619 , n39596 );
    or g39176 ( n26981 , n42852 , n28610 );
    and g39177 ( n6115 , n20961 , n22637 );
    nor g39178 ( n4310 , n27370 , n26827 );
    not g39179 ( n36132 , n20714 );
    or g39180 ( n9854 , n13536 , n14838 );
    not g39181 ( n20544 , n14810 );
    or g39182 ( n40692 , n32087 , n21050 );
    and g39183 ( n11707 , n33310 , n14116 );
    and g39184 ( n7216 , n6921 , n6928 );
    and g39185 ( n21603 , n23684 , n26299 );
    or g39186 ( n41646 , n40612 , n15320 );
    or g39187 ( n36160 , n39402 , n460 );
    and g39188 ( n7114 , n22117 , n306 );
    or g39189 ( n4113 , n25547 , n32770 );
    or g39190 ( n9223 , n16010 , n4452 );
    and g39191 ( n33566 , n32818 , n24445 );
    xnor g39192 ( n34864 , n7585 , n3702 );
    not g39193 ( n11525 , n34922 );
    and g39194 ( n35403 , n29478 , n2357 );
    or g39195 ( n22581 , n4824 , n26933 );
    not g39196 ( n24621 , n36731 );
    nor g39197 ( n28167 , n15217 , n18204 );
    and g39198 ( n41389 , n31353 , n10138 );
    and g39199 ( n16359 , n38209 , n40920 );
    or g39200 ( n23107 , n26298 , n24312 );
    or g39201 ( n15777 , n26915 , n9767 );
    or g39202 ( n25613 , n16598 , n21444 );
    xnor g39203 ( n21397 , n25641 , n15471 );
    and g39204 ( n8881 , n27227 , n10267 );
    or g39205 ( n20552 , n34569 , n191 );
    not g39206 ( n36154 , n20416 );
    nor g39207 ( n41496 , n8125 , n9120 );
    or g39208 ( n35601 , n40978 , n15452 );
    nor g39209 ( n8665 , n11393 , n41864 );
    not g39210 ( n15358 , n16756 );
    nor g39211 ( n18571 , n9180 , n9203 );
    not g39212 ( n17823 , n17567 );
    or g39213 ( n15817 , n32901 , n28827 );
    nor g39214 ( n14966 , n18907 , n11418 );
    nor g39215 ( n30741 , n30985 , n2990 );
    nor g39216 ( n12001 , n8494 , n10476 );
    and g39217 ( n10330 , n3596 , n2534 );
    or g39218 ( n37109 , n9064 , n40520 );
    nor g39219 ( n22828 , n1521 , n37448 );
    or g39220 ( n6897 , n38463 , n24973 );
    nor g39221 ( n40933 , n11526 , n7965 );
    not g39222 ( n34954 , n31246 );
    or g39223 ( n9516 , n34202 , n5343 );
    or g39224 ( n32631 , n36789 , n32315 );
    or g39225 ( n29881 , n18394 , n28500 );
    and g39226 ( n35256 , n23196 , n7942 );
    or g39227 ( n33046 , n5585 , n14360 );
    and g39228 ( n14716 , n31205 , n5080 );
    nor g39229 ( n4607 , n8494 , n3537 );
    and g39230 ( n2838 , n3340 , n30607 );
    or g39231 ( n12481 , n36962 , n35272 );
    not g39232 ( n23707 , n23654 );
    nor g39233 ( n36210 , n3769 , n32044 );
    not g39234 ( n3459 , n10061 );
    and g39235 ( n29619 , n13834 , n33388 );
    nor g39236 ( n7237 , n24536 , n6849 );
    or g39237 ( n11833 , n34791 , n37774 );
    or g39238 ( n12691 , n20932 , n4229 );
    not g39239 ( n22767 , n2253 );
    or g39240 ( n6360 , n16306 , n4376 );
    or g39241 ( n2622 , n8031 , n17991 );
    or g39242 ( n14337 , n22456 , n18644 );
    not g39243 ( n15708 , n22074 );
    and g39244 ( n20788 , n6780 , n37485 );
    nor g39245 ( n21072 , n41306 , n6197 );
    or g39246 ( n25992 , n24729 , n21275 );
    or g39247 ( n25256 , n12867 , n34669 );
    not g39248 ( n6560 , n8465 );
    or g39249 ( n33659 , n39108 , n18521 );
    nor g39250 ( n12859 , n36104 , n35708 );
    or g39251 ( n11717 , n41349 , n16440 );
    nor g39252 ( n41596 , n40108 , n2816 );
    or g39253 ( n28090 , n25721 , n21195 );
    xnor g39254 ( n28734 , n302 , n20071 );
    or g39255 ( n10449 , n37806 , n18751 );
    nor g39256 ( n6141 , n39189 , n19906 );
    or g39257 ( n15650 , n15572 , n42361 );
    nor g39258 ( n7726 , n40332 , n41396 );
    not g39259 ( n5607 , n39579 );
    not g39260 ( n34675 , n13319 );
    or g39261 ( n5019 , n35301 , n20722 );
    and g39262 ( n16724 , n15447 , n1807 );
    not g39263 ( n3148 , n11108 );
    not g39264 ( n35450 , n3198 );
    and g39265 ( n34461 , n21614 , n14674 );
    not g39266 ( n39407 , n9302 );
    xnor g39267 ( n7320 , n15972 , n38305 );
    or g39268 ( n38592 , n31782 , n3410 );
    xnor g39269 ( n9934 , n11046 , n4641 );
    and g39270 ( n26655 , n30997 , n22526 );
    not g39271 ( n23696 , n5084 );
    and g39272 ( n28732 , n27427 , n17127 );
    xnor g39273 ( n39952 , n34154 , n13363 );
    not g39274 ( n20596 , n27033 );
    or g39275 ( n40575 , n3720 , n14535 );
    and g39276 ( n35360 , n27713 , n42889 );
    and g39277 ( n40504 , n35860 , n22996 );
    and g39278 ( n40065 , n36429 , n35392 );
    xnor g39279 ( n28787 , n527 , n28492 );
    not g39280 ( n21498 , n26277 );
    nor g39281 ( n37562 , n26680 , n2924 );
    and g39282 ( n12244 , n39704 , n37518 );
    and g39283 ( n29368 , n20248 , n41064 );
    nor g39284 ( n37037 , n10379 , n25378 );
    xnor g39285 ( n8133 , n10024 , n17194 );
    xnor g39286 ( n36681 , n26689 , n4076 );
    or g39287 ( n21573 , n25184 , n9201 );
    and g39288 ( n39173 , n13221 , n17807 );
    nor g39289 ( n39169 , n5977 , n36584 );
    or g39290 ( n22573 , n40673 , n7790 );
    nor g39291 ( n22108 , n38157 , n26498 );
    and g39292 ( n16104 , n25585 , n18290 );
    or g39293 ( n3079 , n42361 , n39088 );
    and g39294 ( n37898 , n39727 , n31435 );
    nor g39295 ( n9392 , n28708 , n22616 );
    not g39296 ( n10950 , n3362 );
    not g39297 ( n16891 , n861 );
    and g39298 ( n38001 , n36737 , n4269 );
    or g39299 ( n27605 , n41957 , n8715 );
    or g39300 ( n37786 , n3292 , n21682 );
    xnor g39301 ( n3519 , n9307 , n33961 );
    or g39302 ( n19176 , n37894 , n3728 );
    and g39303 ( n17460 , n21070 , n21316 );
    xnor g39304 ( n32333 , n17299 , n25109 );
    not g39305 ( n24958 , n29890 );
    nor g39306 ( n31770 , n42390 , n14919 );
    xnor g39307 ( n33343 , n9155 , n41245 );
    or g39308 ( n17876 , n25233 , n17786 );
    nor g39309 ( n11074 , n15070 , n15080 );
    xnor g39310 ( n34121 , n41013 , n30666 );
    or g39311 ( n37965 , n21466 , n13028 );
    or g39312 ( n2706 , n36739 , n32827 );
    not g39313 ( n32160 , n21675 );
    and g39314 ( n37799 , n15083 , n28182 );
    and g39315 ( n40287 , n26458 , n29666 );
    not g39316 ( n35266 , n10142 );
    not g39317 ( n9748 , n22415 );
    or g39318 ( n33180 , n27552 , n27877 );
    nor g39319 ( n4158 , n2263 , n41136 );
    not g39320 ( n11867 , n10554 );
    or g39321 ( n23992 , n35324 , n32812 );
    and g39322 ( n28571 , n42897 , n19093 );
    or g39323 ( n37209 , n30775 , n22986 );
    xnor g39324 ( n36131 , n28867 , n28904 );
    or g39325 ( n35976 , n26354 , n21900 );
    not g39326 ( n16249 , n33844 );
    xnor g39327 ( n33331 , n39722 , n24431 );
    xnor g39328 ( n41511 , n6625 , n8772 );
    xnor g39329 ( n26187 , n15289 , n2939 );
    or g39330 ( n37815 , n20531 , n3398 );
    or g39331 ( n3707 , n26116 , n657 );
    and g39332 ( n40276 , n10428 , n31709 );
    or g39333 ( n1856 , n24216 , n23931 );
    and g39334 ( n25987 , n14413 , n32229 );
    and g39335 ( n3643 , n19417 , n39964 );
    xnor g39336 ( n8383 , n906 , n24798 );
    and g39337 ( n11093 , n15135 , n5158 );
    or g39338 ( n30565 , n42343 , n38523 );
    nor g39339 ( n15256 , n6573 , n22512 );
    xnor g39340 ( n13290 , n41358 , n7041 );
    nor g39341 ( n6662 , n20820 , n1759 );
    not g39342 ( n27593 , n32384 );
    or g39343 ( n5747 , n30147 , n9935 );
    and g39344 ( n16928 , n19343 , n23889 );
    xnor g39345 ( n15493 , n26123 , n21443 );
    xnor g39346 ( n1661 , n23360 , n13879 );
    or g39347 ( n4071 , n28786 , n3311 );
    xnor g39348 ( n16696 , n36667 , n11660 );
    or g39349 ( n34979 , n20205 , n42057 );
    and g39350 ( n34099 , n20275 , n35987 );
    not g39351 ( n27802 , n28681 );
    nor g39352 ( n21289 , n25334 , n3190 );
    or g39353 ( n27656 , n26397 , n27508 );
    and g39354 ( n37457 , n25547 , n5827 );
    and g39355 ( n41793 , n1312 , n40249 );
    or g39356 ( n23817 , n21882 , n16575 );
    xnor g39357 ( n13865 , n20555 , n30319 );
    and g39358 ( n40448 , n7992 , n34102 );
    or g39359 ( n39242 , n34041 , n3856 );
    xnor g39360 ( n20583 , n27243 , n24377 );
    xnor g39361 ( n14928 , n14979 , n29190 );
    nor g39362 ( n4947 , n14188 , n7504 );
    and g39363 ( n25705 , n30833 , n6133 );
    or g39364 ( n36803 , n22048 , n3323 );
    or g39365 ( n30475 , n24898 , n8216 );
    or g39366 ( n13356 , n31265 , n16421 );
    not g39367 ( n33884 , n19485 );
    and g39368 ( n30450 , n3793 , n23111 );
    xnor g39369 ( n24975 , n34617 , n13891 );
    and g39370 ( n26947 , n5616 , n28047 );
    xnor g39371 ( n9300 , n37539 , n17720 );
    or g39372 ( n26293 , n11254 , n26545 );
    nor g39373 ( n39151 , n11319 , n32681 );
    xnor g39374 ( n138 , n31989 , n14894 );
    and g39375 ( n38008 , n31338 , n38086 );
    and g39376 ( n1035 , n27747 , n11616 );
    or g39377 ( n2730 , n17346 , n28357 );
    or g39378 ( n1089 , n18424 , n40272 );
    or g39379 ( n24485 , n19221 , n31370 );
    or g39380 ( n8932 , n27721 , n28206 );
    xnor g39381 ( n37548 , n30778 , n22034 );
    nor g39382 ( n5329 , n25875 , n14877 );
    and g39383 ( n12762 , n26513 , n2371 );
    not g39384 ( n9241 , n5566 );
    not g39385 ( n8656 , n29474 );
    or g39386 ( n24128 , n1985 , n31860 );
    or g39387 ( n22304 , n4585 , n5467 );
    not g39388 ( n2564 , n28133 );
    xnor g39389 ( n13895 , n32470 , n12665 );
    or g39390 ( n26707 , n24147 , n27738 );
    or g39391 ( n7160 , n33946 , n244 );
    or g39392 ( n40096 , n1312 , n40249 );
    xnor g39393 ( n41697 , n784 , n870 );
    or g39394 ( n34799 , n27773 , n27127 );
    not g39395 ( n6541 , n26290 );
    and g39396 ( n38869 , n24700 , n25091 );
    or g39397 ( n42684 , n18563 , n7333 );
    and g39398 ( n3088 , n13110 , n39048 );
    or g39399 ( n11365 , n5292 , n13520 );
    or g39400 ( n3043 , n9384 , n16683 );
    xnor g39401 ( n24306 , n22103 , n1774 );
    or g39402 ( n9282 , n4473 , n1995 );
    xnor g39403 ( n26513 , n33416 , n31301 );
    nor g39404 ( n4337 , n23101 , n3036 );
    or g39405 ( n10522 , n1023 , n38560 );
    or g39406 ( n10695 , n5348 , n15294 );
    and g39407 ( n39625 , n37526 , n4163 );
    and g39408 ( n21833 , n33896 , n4348 );
    or g39409 ( n10882 , n13667 , n22313 );
    not g39410 ( n792 , n26515 );
    not g39411 ( n11288 , n18176 );
    xnor g39412 ( n5674 , n36628 , n41723 );
    nor g39413 ( n26632 , n39384 , n11483 );
    or g39414 ( n4958 , n33144 , n8338 );
    or g39415 ( n12584 , n30110 , n15082 );
    xnor g39416 ( n1907 , n15972 , n457 );
    not g39417 ( n7991 , n5843 );
    nor g39418 ( n26088 , n2199 , n33900 );
    nor g39419 ( n2401 , n9465 , n40715 );
    xnor g39420 ( n35199 , n25619 , n26281 );
    or g39421 ( n35106 , n35109 , n17785 );
    nor g39422 ( n28312 , n20904 , n33447 );
    or g39423 ( n1614 , n40814 , n1035 );
    or g39424 ( n2842 , n39983 , n28908 );
    and g39425 ( n30283 , n38895 , n38759 );
    xnor g39426 ( n443 , n12769 , n27933 );
    or g39427 ( n8583 , n23380 , n3543 );
    or g39428 ( n4120 , n5444 , n7294 );
    or g39429 ( n24225 , n4504 , n3229 );
    and g39430 ( n28633 , n40533 , n36054 );
    or g39431 ( n1766 , n21442 , n19497 );
    and g39432 ( n24300 , n39434 , n23752 );
    or g39433 ( n22689 , n22969 , n1425 );
    xnor g39434 ( n28070 , n11051 , n11305 );
    not g39435 ( n1116 , n15056 );
    or g39436 ( n40841 , n22389 , n10709 );
    and g39437 ( n37970 , n19609 , n42207 );
    or g39438 ( n32776 , n18542 , n41993 );
    or g39439 ( n37813 , n6282 , n38153 );
    not g39440 ( n22585 , n11403 );
    nor g39441 ( n28230 , n39829 , n3141 );
    nor g39442 ( n22707 , n33981 , n11306 );
    or g39443 ( n26821 , n15222 , n12317 );
    xnor g39444 ( n29087 , n31989 , n10691 );
    not g39445 ( n5850 , n2018 );
    nor g39446 ( n31543 , n6377 , n15790 );
    nor g39447 ( n28733 , n5964 , n35554 );
    and g39448 ( n42288 , n14715 , n32555 );
    or g39449 ( n36920 , n41063 , n38874 );
    xnor g39450 ( n35741 , n21826 , n30976 );
    not g39451 ( n28648 , n39200 );
    or g39452 ( n20247 , n28032 , n23747 );
    not g39453 ( n10720 , n25947 );
    or g39454 ( n41753 , n39439 , n33248 );
    nor g39455 ( n32929 , n2257 , n42246 );
    xnor g39456 ( n8400 , n25582 , n28025 );
    or g39457 ( n7494 , n2199 , n12887 );
    and g39458 ( n27036 , n26750 , n10376 );
    or g39459 ( n33011 , n39462 , n34646 );
    or g39460 ( n30147 , n8539 , n15653 );
    and g39461 ( n30393 , n5095 , n8554 );
    and g39462 ( n1701 , n16105 , n25455 );
    and g39463 ( n37996 , n7323 , n17582 );
    xnor g39464 ( n42162 , n4877 , n207 );
    or g39465 ( n17094 , n25336 , n10850 );
    or g39466 ( n37206 , n5701 , n18898 );
    not g39467 ( n13628 , n6441 );
    or g39468 ( n26532 , n12130 , n9000 );
    and g39469 ( n38998 , n13789 , n16428 );
    not g39470 ( n26650 , n39870 );
    nor g39471 ( n14694 , n35134 , n24135 );
    or g39472 ( n17866 , n23582 , n3311 );
    not g39473 ( n13881 , n34115 );
    and g39474 ( n23651 , n15992 , n21789 );
    xnor g39475 ( n23600 , n41013 , n34712 );
    xnor g39476 ( n16469 , n31051 , n5964 );
    xnor g39477 ( n19904 , n20436 , n35301 );
    and g39478 ( n41714 , n30962 , n23734 );
    nor g39479 ( n23126 , n40902 , n38867 );
    or g39480 ( n33347 , n29988 , n3112 );
    xnor g39481 ( n23490 , n12282 , n14651 );
    and g39482 ( n15302 , n35472 , n24669 );
    xnor g39483 ( n1435 , n34731 , n12698 );
    or g39484 ( n38023 , n42229 , n33537 );
    or g39485 ( n12067 , n31843 , n23879 );
    or g39486 ( n1781 , n41472 , n13348 );
    and g39487 ( n17656 , n37546 , n31599 );
    or g39488 ( n38637 , n36235 , n38698 );
    or g39489 ( n15978 , n20200 , n8989 );
    nor g39490 ( n38582 , n40728 , n15085 );
    and g39491 ( n33071 , n2604 , n20153 );
    not g39492 ( n28184 , n2366 );
    or g39493 ( n20475 , n23563 , n38078 );
    or g39494 ( n20857 , n37879 , n19244 );
    or g39495 ( n885 , n16417 , n30540 );
    and g39496 ( n832 , n36678 , n6801 );
    xnor g39497 ( n37423 , n21941 , n19809 );
    or g39498 ( n33791 , n20477 , n34374 );
    nor g39499 ( n29480 , n1141 , n27954 );
    xnor g39500 ( n27687 , n30326 , n2199 );
    or g39501 ( n28179 , n41534 , n30853 );
    and g39502 ( n6734 , n9249 , n42011 );
    and g39503 ( n28074 , n27281 , n12042 );
    or g39504 ( n25905 , n1507 , n32549 );
    or g39505 ( n22793 , n39905 , n26112 );
    or g39506 ( n12533 , n4034 , n4830 );
    or g39507 ( n37000 , n15064 , n13449 );
    not g39508 ( n31474 , n27419 );
    or g39509 ( n30457 , n23323 , n12714 );
    and g39510 ( n1263 , n18963 , n24805 );
    xnor g39511 ( n22736 , n27396 , n31614 );
    xnor g39512 ( n38856 , n203 , n34292 );
    and g39513 ( n31949 , n37536 , n20838 );
    and g39514 ( n1226 , n23532 , n5127 );
    and g39515 ( n38135 , n5700 , n16187 );
    or g39516 ( n9866 , n33268 , n26586 );
    or g39517 ( n22566 , n39699 , n19457 );
    or g39518 ( n37746 , n42816 , n21502 );
    and g39519 ( n37553 , n3232 , n13342 );
    or g39520 ( n11388 , n29135 , n9202 );
    or g39521 ( n17186 , n16116 , n21659 );
    or g39522 ( n9729 , n17253 , n20877 );
    xnor g39523 ( n12657 , n5808 , n35036 );
    or g39524 ( n39644 , n23795 , n12669 );
    xnor g39525 ( n25616 , n3855 , n8494 );
    and g39526 ( n29552 , n22629 , n33993 );
    or g39527 ( n6434 , n9821 , n7378 );
    or g39528 ( n23367 , n22742 , n5048 );
    xnor g39529 ( n17019 , n26210 , n36279 );
    not g39530 ( n2799 , n12224 );
    or g39531 ( n40691 , n33066 , n2012 );
    and g39532 ( n3367 , n3176 , n6532 );
    or g39533 ( n11462 , n2346 , n28837 );
    or g39534 ( n41701 , n30603 , n36641 );
    and g39535 ( n12789 , n21097 , n24842 );
    not g39536 ( n5147 , n25288 );
    or g39537 ( n36591 , n25573 , n13872 );
    nor g39538 ( n6915 , n5353 , n30837 );
    or g39539 ( n27117 , n1859 , n14211 );
    not g39540 ( n36235 , n499 );
    and g39541 ( n20473 , n24289 , n13579 );
    nor g39542 ( n15405 , n25588 , n11229 );
    xnor g39543 ( n13173 , n31460 , n39373 );
    xnor g39544 ( n31391 , n3501 , n14471 );
    or g39545 ( n23048 , n33795 , n23069 );
    xnor g39546 ( n20026 , n21415 , n4884 );
    and g39547 ( n7558 , n30327 , n26012 );
    or g39548 ( n24133 , n18968 , n27111 );
    or g39549 ( n26318 , n33981 , n8468 );
    and g39550 ( n10888 , n18656 , n37383 );
    nor g39551 ( n9467 , n7063 , n37841 );
    or g39552 ( n22497 , n10752 , n30225 );
    xnor g39553 ( n7774 , n5708 , n26411 );
    nor g39554 ( n35184 , n28710 , n3606 );
    nor g39555 ( n9021 , n12787 , n39368 );
    or g39556 ( n42037 , n26130 , n16163 );
    not g39557 ( n14758 , n9512 );
    and g39558 ( n12840 , n31799 , n16790 );
    xnor g39559 ( n28473 , n4872 , n27327 );
    not g39560 ( n23819 , n10388 );
    and g39561 ( n990 , n4529 , n7693 );
    or g39562 ( n24720 , n18798 , n3091 );
    not g39563 ( n33889 , n41430 );
    or g39564 ( n12466 , n34842 , n6560 );
    or g39565 ( n6498 , n18857 , n36580 );
    xnor g39566 ( n19584 , n41318 , n14707 );
    not g39567 ( n3106 , n2635 );
    xnor g39568 ( n42866 , n13444 , n39884 );
    or g39569 ( n40098 , n34565 , n3514 );
    xnor g39570 ( n42347 , n32297 , n29368 );
    and g39571 ( n24973 , n36888 , n27615 );
    or g39572 ( n36729 , n12392 , n24564 );
    and g39573 ( n38729 , n41792 , n32067 );
    nor g39574 ( n22375 , n38650 , n1616 );
    or g39575 ( n25658 , n137 , n6694 );
    or g39576 ( n25773 , n1696 , n19207 );
    xnor g39577 ( n7478 , n20539 , n14893 );
    and g39578 ( n21788 , n42413 , n10133 );
    or g39579 ( n42578 , n40703 , n18706 );
    or g39580 ( n25472 , n10249 , n18937 );
    xnor g39581 ( n26955 , n37210 , n38678 );
    or g39582 ( n12712 , n19294 , n2802 );
    not g39583 ( n38173 , n26575 );
    and g39584 ( n22448 , n4423 , n14518 );
    or g39585 ( n8424 , n1447 , n26854 );
    or g39586 ( n40417 , n6273 , n13744 );
    or g39587 ( n21350 , n5140 , n5602 );
    not g39588 ( n20462 , n22303 );
    or g39589 ( n4523 , n12354 , n4669 );
    or g39590 ( n20642 , n32277 , n31991 );
    or g39591 ( n1376 , n2284 , n9479 );
    and g39592 ( n38052 , n10909 , n16716 );
    not g39593 ( n25413 , n8357 );
    or g39594 ( n25593 , n30550 , n42797 );
    or g39595 ( n7128 , n41809 , n6316 );
    or g39596 ( n37158 , n25576 , n38239 );
    or g39597 ( n8247 , n24134 , n14825 );
    or g39598 ( n30915 , n10491 , n3330 );
    nor g39599 ( n29061 , n15289 , n16692 );
    or g39600 ( n4628 , n16904 , n11144 );
    not g39601 ( n17483 , n7914 );
    and g39602 ( n10402 , n28004 , n19051 );
    nor g39603 ( n31851 , n23511 , n29857 );
    not g39604 ( n27188 , n499 );
    or g39605 ( n39359 , n11417 , n39958 );
    xnor g39606 ( n12004 , n585 , n11626 );
    and g39607 ( n34060 , n22433 , n33001 );
    nor g39608 ( n38028 , n1891 , n41619 );
    or g39609 ( n11355 , n9910 , n36578 );
    or g39610 ( n6652 , n26904 , n36080 );
    or g39611 ( n25415 , n20797 , n17070 );
    and g39612 ( n5774 , n23704 , n17962 );
    not g39613 ( n32265 , n20311 );
    not g39614 ( n1069 , n3339 );
    or g39615 ( n28306 , n36052 , n30620 );
    not g39616 ( n41065 , n34933 );
    nor g39617 ( n30498 , n24115 , n26478 );
    not g39618 ( n190 , n36612 );
    nor g39619 ( n4220 , n24549 , n29320 );
    xnor g39620 ( n39886 , n12605 , n16556 );
    or g39621 ( n27067 , n18190 , n3386 );
    nor g39622 ( n2745 , n40086 , n42532 );
    and g39623 ( n22758 , n21534 , n37560 );
    or g39624 ( n2749 , n17526 , n37836 );
    or g39625 ( n2137 , n1980 , n15624 );
    xnor g39626 ( n15153 , n21877 , n11820 );
    or g39627 ( n35078 , n28390 , n32892 );
    xnor g39628 ( n19856 , n31099 , n23621 );
    or g39629 ( n5562 , n6712 , n17729 );
    or g39630 ( n28687 , n27952 , n29287 );
    nor g39631 ( n33529 , n212 , n40873 );
    not g39632 ( n37083 , n12634 );
    or g39633 ( n15105 , n16575 , n27606 );
    or g39634 ( n24959 , n38314 , n31911 );
    or g39635 ( n13114 , n11622 , n4355 );
    or g39636 ( n10300 , n25939 , n33537 );
    not g39637 ( n29138 , n26434 );
    or g39638 ( n22283 , n32772 , n15505 );
    nor g39639 ( n28204 , n39266 , n8891 );
    and g39640 ( n41382 , n5234 , n25816 );
    not g39641 ( n24718 , n21530 );
    nor g39642 ( n33993 , n9001 , n6292 );
    nor g39643 ( n13562 , n9792 , n31300 );
    or g39644 ( n42797 , n25130 , n31707 );
    or g39645 ( n9091 , n23472 , n23756 );
    or g39646 ( n21753 , n12980 , n34967 );
    and g39647 ( n26884 , n19837 , n11602 );
    and g39648 ( n9967 , n40982 , n36516 );
    nor g39649 ( n31139 , n6147 , n18149 );
    or g39650 ( n41672 , n41625 , n30233 );
    or g39651 ( n24360 , n22203 , n37671 );
    or g39652 ( n21009 , n4895 , n37904 );
    or g39653 ( n531 , n37072 , n22597 );
    xnor g39654 ( n9661 , n35347 , n22876 );
    or g39655 ( n26015 , n19701 , n33263 );
    or g39656 ( n28169 , n17120 , n912 );
    not g39657 ( n18475 , n32597 );
    and g39658 ( n38048 , n2098 , n40774 );
    or g39659 ( n13231 , n711 , n33858 );
    xnor g39660 ( n17387 , n3068 , n12914 );
    or g39661 ( n5903 , n12764 , n38142 );
    or g39662 ( n39622 , n8681 , n5083 );
    or g39663 ( n41711 , n28149 , n41581 );
    or g39664 ( n18431 , n25233 , n13004 );
    or g39665 ( n26562 , n29058 , n26594 );
    or g39666 ( n40818 , n27921 , n40483 );
    not g39667 ( n30605 , n19229 );
    or g39668 ( n30111 , n14481 , n14273 );
    not g39669 ( n8475 , n8215 );
    and g39670 ( n6792 , n44 , n36746 );
    or g39671 ( n20662 , n5962 , n3946 );
    xnor g39672 ( n39754 , n36009 , n18703 );
    or g39673 ( n9572 , n38208 , n42349 );
    and g39674 ( n8198 , n984 , n13591 );
    nor g39675 ( n777 , n17768 , n41688 );
    nor g39676 ( n34360 , n34565 , n36506 );
    nor g39677 ( n19695 , n5788 , n41204 );
    xnor g39678 ( n35984 , n35140 , n5896 );
    and g39679 ( n40300 , n8947 , n6879 );
    nor g39680 ( n11079 , n35874 , n18889 );
    or g39681 ( n29105 , n24979 , n27540 );
    or g39682 ( n19759 , n19969 , n39027 );
    and g39683 ( n7612 , n32981 , n15326 );
    nor g39684 ( n8082 , n38621 , n40139 );
    or g39685 ( n28047 , n34195 , n37724 );
    and g39686 ( n4023 , n42363 , n23409 );
    and g39687 ( n39521 , n42772 , n31507 );
    nor g39688 ( n36574 , n8494 , n17356 );
    or g39689 ( n40580 , n12840 , n26789 );
    and g39690 ( n37516 , n36338 , n14251 );
    xnor g39691 ( n28248 , n17220 , n38924 );
    xnor g39692 ( n3918 , n12145 , n5937 );
    nor g39693 ( n16680 , n17120 , n29344 );
    not g39694 ( n11050 , n26992 );
    or g39695 ( n34707 , n27685 , n37584 );
    and g39696 ( n1086 , n15495 , n2313 );
    not g39697 ( n2985 , n2825 );
    not g39698 ( n37800 , n17386 );
    or g39699 ( n19234 , n12698 , n11814 );
    xnor g39700 ( n1081 , n12146 , n10155 );
    or g39701 ( n8264 , n36365 , n15392 );
    or g39702 ( n5544 , n28867 , n36851 );
    or g39703 ( n26084 , n27878 , n34195 );
    or g39704 ( n35885 , n33560 , n5090 );
    or g39705 ( n20898 , n14851 , n30447 );
    or g39706 ( n38190 , n38781 , n24151 );
    or g39707 ( n3762 , n25053 , n38937 );
    or g39708 ( n1094 , n24626 , n26330 );
    xnor g39709 ( n31532 , n25619 , n35131 );
    and g39710 ( n19422 , n25111 , n9120 );
    xnor g39711 ( n25823 , n15524 , n17031 );
    or g39712 ( n13794 , n20993 , n20498 );
    not g39713 ( n1997 , n13144 );
    or g39714 ( n16165 , n2193 , n26891 );
    or g39715 ( n29235 , n9218 , n790 );
    not g39716 ( n23694 , n32727 );
    or g39717 ( n12838 , n20138 , n28485 );
    not g39718 ( n10791 , n19526 );
    and g39719 ( n29430 , n8785 , n42835 );
    not g39720 ( n28053 , n3172 );
    or g39721 ( n16460 , n20246 , n16891 );
    or g39722 ( n36599 , n7604 , n5779 );
    not g39723 ( n33780 , n53 );
    not g39724 ( n27744 , n56 );
    or g39725 ( n16435 , n37664 , n15255 );
    and g39726 ( n21094 , n30722 , n30836 );
    and g39727 ( n38958 , n34622 , n33458 );
    not g39728 ( n4669 , n24447 );
    or g39729 ( n5223 , n23971 , n2362 );
    not g39730 ( n41955 , n39158 );
    or g39731 ( n8158 , n24212 , n3504 );
    and g39732 ( n39048 , n13656 , n23654 );
    not g39733 ( n5445 , n26014 );
    or g39734 ( n2371 , n10518 , n8384 );
    or g39735 ( n37717 , n17042 , n39350 );
    or g39736 ( n5489 , n8014 , n28402 );
    nor g39737 ( n5624 , n38873 , n25796 );
    or g39738 ( n4581 , n10625 , n39949 );
    xnor g39739 ( n4343 , n42003 , n4374 );
    or g39740 ( n19207 , n23707 , n25064 );
    or g39741 ( n19976 , n25430 , n7616 );
    and g39742 ( n34726 , n2176 , n41988 );
    or g39743 ( n39956 , n6632 , n28596 );
    nor g39744 ( n1952 , n21727 , n19492 );
    or g39745 ( n5058 , n17948 , n4329 );
    xnor g39746 ( n11584 , n18530 , n34418 );
    or g39747 ( n41064 , n7864 , n33619 );
    or g39748 ( n2574 , n3444 , n17623 );
    and g39749 ( n9847 , n15732 , n21477 );
    or g39750 ( n13083 , n38659 , n34553 );
    or g39751 ( n38672 , n12867 , n24784 );
    and g39752 ( n35093 , n7562 , n2423 );
    nor g39753 ( n35437 , n30546 , n42848 );
    not g39754 ( n35588 , n7207 );
    or g39755 ( n42080 , n20932 , n1462 );
    xnor g39756 ( n40048 , n6164 , n27521 );
    not g39757 ( n23228 , n32057 );
    or g39758 ( n6729 , n9275 , n14618 );
    and g39759 ( n12756 , n27144 , n29594 );
    not g39760 ( n38211 , n20766 );
    or g39761 ( n28512 , n17427 , n4076 );
    or g39762 ( n13378 , n3781 , n41628 );
    and g39763 ( n30088 , n2682 , n27050 );
    not g39764 ( n36344 , n14900 );
    or g39765 ( n1359 , n39420 , n11753 );
    xnor g39766 ( n38902 , n3296 , n1686 );
    and g39767 ( n9328 , n38446 , n25977 );
    or g39768 ( n24377 , n20142 , n26203 );
    nor g39769 ( n26744 , n36271 , n28356 );
    or g39770 ( n39670 , n32800 , n7893 );
    or g39771 ( n29175 , n18424 , n22928 );
    or g39772 ( n25421 , n16016 , n17030 );
    and g39773 ( n30046 , n10257 , n12300 );
    xnor g39774 ( n25976 , n13984 , n11205 );
    or g39775 ( n35694 , n18334 , n4355 );
    nor g39776 ( n23446 , n42282 , n38728 );
    xnor g39777 ( n14920 , n22437 , n40074 );
    and g39778 ( n8530 , n6224 , n37407 );
    xnor g39779 ( n26114 , n38350 , n1266 );
    and g39780 ( n40543 , n4049 , n2866 );
    or g39781 ( n39985 , n40728 , n12315 );
    not g39782 ( n38807 , n27562 );
    xnor g39783 ( n20285 , n22998 , n25588 );
    or g39784 ( n26812 , n10199 , n33117 );
    or g39785 ( n31193 , n11806 , n13813 );
    or g39786 ( n12513 , n40664 , n2296 );
    or g39787 ( n25387 , n17410 , n14501 );
    and g39788 ( n20865 , n5451 , n3111 );
    and g39789 ( n25383 , n10273 , n7895 );
    or g39790 ( n25037 , n22509 , n41037 );
    and g39791 ( n26071 , n34099 , n42827 );
    and g39792 ( n32063 , n3153 , n42022 );
    xnor g39793 ( n31566 , n11304 , n4419 );
    nor g39794 ( n4778 , n21545 , n4483 );
    and g39795 ( n12796 , n34185 , n11083 );
    or g39796 ( n18443 , n26832 , n6359 );
    and g39797 ( n15762 , n23600 , n24090 );
    or g39798 ( n39698 , n31035 , n6098 );
    not g39799 ( n15457 , n41191 );
    or g39800 ( n18248 , n16496 , n5282 );
    not g39801 ( n17578 , n37248 );
    and g39802 ( n32326 , n38946 , n19921 );
    or g39803 ( n8396 , n26075 , n15421 );
    and g39804 ( n35432 , n6497 , n1832 );
    and g39805 ( n42841 , n31673 , n22565 );
    and g39806 ( n22858 , n35428 , n6795 );
    or g39807 ( n11227 , n30263 , n20189 );
    or g39808 ( n5436 , n14048 , n16002 );
    or g39809 ( n24543 , n22025 , n25626 );
    or g39810 ( n26462 , n25902 , n42254 );
    and g39811 ( n15943 , n26131 , n5709 );
    xnor g39812 ( n1594 , n34731 , n4751 );
    nor g39813 ( n7341 , n10522 , n6951 );
    or g39814 ( n36303 , n23750 , n2565 );
    or g39815 ( n4413 , n24264 , n12967 );
    nor g39816 ( n28832 , n18866 , n31751 );
    and g39817 ( n870 , n27935 , n38449 );
    xnor g39818 ( n4554 , n31896 , n28845 );
    or g39819 ( n14915 , n36585 , n35306 );
    or g39820 ( n17591 , n17828 , n5524 );
    or g39821 ( n32944 , n38423 , n31464 );
    nor g39822 ( n40945 , n28261 , n16877 );
    or g39823 ( n22403 , n32228 , n19352 );
    nor g39824 ( n10975 , n35611 , n9838 );
    or g39825 ( n30819 , n18976 , n33289 );
    nor g39826 ( n32288 , n36042 , n35821 );
    or g39827 ( n42116 , n11438 , n31421 );
    nor g39828 ( n9343 , n36625 , n18842 );
    xnor g39829 ( n5494 , n6621 , n11190 );
    and g39830 ( n38056 , n29145 , n19569 );
    or g39831 ( n499 , n37430 , n8105 );
    or g39832 ( n2981 , n19392 , n19171 );
    or g39833 ( n40552 , n20092 , n34956 );
    or g39834 ( n35228 , n38953 , n29507 );
    and g39835 ( n17124 , n4064 , n40205 );
    xnor g39836 ( n36552 , n42064 , n12887 );
    or g39837 ( n32821 , n34016 , n35772 );
    not g39838 ( n21789 , n28498 );
    or g39839 ( n23076 , n39913 , n16741 );
    xnor g39840 ( n25140 , n42131 , n34593 );
    or g39841 ( n8537 , n17193 , n8541 );
    nor g39842 ( n4461 , n36238 , n33359 );
    and g39843 ( n19783 , n17228 , n2620 );
    nor g39844 ( n32638 , n24182 , n17716 );
    and g39845 ( n387 , n7451 , n2520 );
    or g39846 ( n31197 , n12776 , n38379 );
    not g39847 ( n17527 , n11085 );
    or g39848 ( n26619 , n37415 , n41836 );
    xnor g39849 ( n937 , n9370 , n41809 );
    nor g39850 ( n21059 , n34402 , n35889 );
    or g39851 ( n13302 , n36789 , n36282 );
    or g39852 ( n6427 , n4207 , n34569 );
    xnor g39853 ( n26907 , n12146 , n20381 );
    xnor g39854 ( n8061 , n35876 , n25205 );
    nor g39855 ( n40716 , n6149 , n18802 );
    and g39856 ( n26295 , n23938 , n15408 );
    or g39857 ( n22042 , n23176 , n439 );
    or g39858 ( n15851 , n6930 , n38753 );
    and g39859 ( n35815 , n20651 , n20438 );
    and g39860 ( n19589 , n41031 , n10877 );
    and g39861 ( n32293 , n26221 , n28244 );
    and g39862 ( n26714 , n40029 , n33808 );
    xnor g39863 ( n23565 , n18235 , n15925 );
    or g39864 ( n32546 , n17874 , n27347 );
    or g39865 ( n32128 , n25830 , n5504 );
    nor g39866 ( n25813 , n28353 , n34264 );
    or g39867 ( n3688 , n19221 , n29531 );
    and g39868 ( n35321 , n31226 , n42014 );
    and g39869 ( n8384 , n26703 , n31329 );
    or g39870 ( n21452 , n31227 , n1509 );
    or g39871 ( n34176 , n17903 , n11641 );
    or g39872 ( n25462 , n42909 , n5110 );
    nor g39873 ( n32036 , n10939 , n6524 );
    not g39874 ( n39921 , n3425 );
    and g39875 ( n33398 , n17663 , n17902 );
    and g39876 ( n29752 , n20320 , n18396 );
    not g39877 ( n8390 , n32507 );
    and g39878 ( n10467 , n39029 , n40425 );
    or g39879 ( n33018 , n19645 , n16273 );
    xnor g39880 ( n38077 , n26864 , n36436 );
    or g39881 ( n19606 , n5365 , n1735 );
    or g39882 ( n27339 , n13777 , n42775 );
    or g39883 ( n25953 , n17037 , n3728 );
    and g39884 ( n2563 , n20380 , n15920 );
    not g39885 ( n24426 , n18110 );
    or g39886 ( n20059 , n2368 , n41271 );
    or g39887 ( n2757 , n14904 , n39123 );
    or g39888 ( n35824 , n23292 , n24383 );
    and g39889 ( n19484 , n26447 , n9739 );
    xnor g39890 ( n42036 , n8194 , n41799 );
    or g39891 ( n22518 , n29943 , n4043 );
    not g39892 ( n2135 , n40372 );
    and g39893 ( n37519 , n671 , n12743 );
    or g39894 ( n35038 , n38725 , n13804 );
    and g39895 ( n23842 , n156 , n17462 );
    or g39896 ( n16086 , n22723 , n16488 );
    or g39897 ( n9996 , n395 , n19422 );
    or g39898 ( n129 , n13640 , n3160 );
    or g39899 ( n42286 , n22143 , n26001 );
    xnor g39900 ( n25611 , n9180 , n38237 );
    or g39901 ( n29275 , n29520 , n6290 );
    not g39902 ( n39489 , n23184 );
    and g39903 ( n23071 , n27421 , n24981 );
    xnor g39904 ( n41631 , n3316 , n34565 );
    or g39905 ( n11156 , n11143 , n981 );
    and g39906 ( n363 , n37071 , n24252 );
    and g39907 ( n22065 , n40991 , n38398 );
    and g39908 ( n38525 , n14654 , n24337 );
    not g39909 ( n13398 , n18012 );
    nor g39910 ( n21864 , n38879 , n8111 );
    nor g39911 ( n7754 , n38829 , n3302 );
    and g39912 ( n22602 , n564 , n3626 );
    and g39913 ( n15714 , n7622 , n1700 );
    and g39914 ( n6335 , n30244 , n24710 );
    or g39915 ( n18411 , n38615 , n37633 );
    and g39916 ( n14980 , n2137 , n32692 );
    or g39917 ( n35335 , n16060 , n15564 );
    or g39918 ( n6656 , n14723 , n12850 );
    or g39919 ( n35592 , n33835 , n22282 );
    or g39920 ( n22613 , n34793 , n18084 );
    or g39921 ( n33664 , n20928 , n25626 );
    nor g39922 ( n29950 , n27875 , n37275 );
    or g39923 ( n12795 , n21235 , n23226 );
    or g39924 ( n39891 , n34190 , n39893 );
    or g39925 ( n1008 , n29372 , n1167 );
    not g39926 ( n41116 , n1477 );
    or g39927 ( n15660 , n698 , n34793 );
    xnor g39928 ( n40883 , n34352 , n8294 );
    not g39929 ( n27686 , n1616 );
    and g39930 ( n33139 , n38081 , n32998 );
    or g39931 ( n19423 , n19958 , n16595 );
    or g39932 ( n21644 , n295 , n11968 );
    or g39933 ( n15862 , n3427 , n37183 );
    or g39934 ( n41551 , n1426 , n735 );
    or g39935 ( n8357 , n11271 , n2073 );
    not g39936 ( n22728 , n34833 );
    and g39937 ( n36812 , n7119 , n34647 );
    and g39938 ( n41126 , n31229 , n6040 );
    or g39939 ( n21548 , n9549 , n20041 );
    or g39940 ( n17403 , n1980 , n19325 );
    xnor g39941 ( n6695 , n29740 , n4816 );
    or g39942 ( n4396 , n20141 , n5677 );
    not g39943 ( n39327 , n22128 );
    or g39944 ( n35169 , n7409 , n27037 );
    or g39945 ( n37405 , n4787 , n38751 );
    and g39946 ( n2204 , n8515 , n33415 );
    and g39947 ( n27804 , n8186 , n40308 );
    not g39948 ( n28837 , n35356 );
    or g39949 ( n23932 , n27311 , n18639 );
    not g39950 ( n2323 , n29625 );
    xnor g39951 ( n8025 , n39559 , n21805 );
    xnor g39952 ( n15887 , n32470 , n32167 );
    not g39953 ( n5759 , n42550 );
    and g39954 ( n39056 , n5516 , n25472 );
    and g39955 ( n29498 , n37897 , n34579 );
    and g39956 ( n11789 , n11360 , n6123 );
    not g39957 ( n7615 , n31668 );
    nor g39958 ( n11761 , n28684 , n14188 );
    and g39959 ( n34000 , n17800 , n17392 );
    not g39960 ( n32264 , n35315 );
    not g39961 ( n24317 , n25035 );
    or g39962 ( n30442 , n10986 , n42535 );
    not g39963 ( n17276 , n42811 );
    or g39964 ( n11334 , n31046 , n15165 );
    nor g39965 ( n29787 , n5964 , n939 );
    or g39966 ( n38043 , n36833 , n4522 );
    not g39967 ( n8938 , n14421 );
    or g39968 ( n23364 , n19911 , n37342 );
    not g39969 ( n4776 , n14439 );
    or g39970 ( n23471 , n22173 , n122 );
    or g39971 ( n28793 , n7752 , n8626 );
    and g39972 ( n33033 , n13502 , n15019 );
    nor g39973 ( n20862 , n155 , n34966 );
    or g39974 ( n25503 , n21521 , n12663 );
    not g39975 ( n24093 , n35455 );
    xnor g39976 ( n21599 , n13296 , n8581 );
    xnor g39977 ( n16102 , n5606 , n21200 );
    or g39978 ( n40789 , n22648 , n15707 );
    not g39979 ( n33289 , n17327 );
    xnor g39980 ( n31250 , n38334 , n37260 );
    nor g39981 ( n15513 , n34307 , n13484 );
    and g39982 ( n9163 , n8010 , n22068 );
    or g39983 ( n26837 , n40512 , n12056 );
    and g39984 ( n37916 , n7063 , n37841 );
    or g39985 ( n4939 , n41756 , n21007 );
    or g39986 ( n40378 , n5004 , n38006 );
    or g39987 ( n11750 , n16586 , n21160 );
    and g39988 ( n9840 , n40919 , n37206 );
    not g39989 ( n24356 , n21293 );
    and g39990 ( n40477 , n1945 , n10436 );
    or g39991 ( n33510 , n33344 , n4689 );
    and g39992 ( n15671 , n41816 , n21693 );
    or g39993 ( n9261 , n22091 , n42488 );
    or g39994 ( n10482 , n37898 , n15411 );
    not g39995 ( n366 , n6809 );
    and g39996 ( n37925 , n25662 , n15742 );
    not g39997 ( n30540 , n21518 );
    not g39998 ( n14224 , n8900 );
    not g39999 ( n9544 , n23369 );
    and g40000 ( n31886 , n25428 , n982 );
    or g40001 ( n7352 , n855 , n22715 );
    nor g40002 ( n11579 , n42580 , n10452 );
    and g40003 ( n39749 , n41005 , n23952 );
    or g40004 ( n919 , n12295 , n12236 );
    not g40005 ( n31924 , n5947 );
    not g40006 ( n246 , n13301 );
    not g40007 ( n39243 , n26558 );
    nor g40008 ( n22943 , n22057 , n967 );
    or g40009 ( n34368 , n4081 , n36235 );
    nor g40010 ( n15615 , n37771 , n8701 );
    or g40011 ( n17601 , n40751 , n17605 );
    and g40012 ( n19210 , n26154 , n39400 );
    xnor g40013 ( n3468 , n20904 , n13605 );
    and g40014 ( n3659 , n37276 , n40171 );
    or g40015 ( n41149 , n481 , n18296 );
    or g40016 ( n8179 , n4018 , n17599 );
    not g40017 ( n38947 , n13072 );
    or g40018 ( n5694 , n1162 , n11485 );
    nor g40019 ( n26626 , n36117 , n11637 );
    and g40020 ( n35997 , n36607 , n39834 );
    xnor g40021 ( n24420 , n21954 , n32719 );
    xnor g40022 ( n5948 , n6962 , n10406 );
    and g40023 ( n36479 , n34382 , n39156 );
    or g40024 ( n15489 , n32997 , n40114 );
    and g40025 ( n3356 , n24930 , n31262 );
    or g40026 ( n11104 , n2746 , n42370 );
    xnor g40027 ( n32155 , n9242 , n32249 );
    not g40028 ( n17196 , n26973 );
    or g40029 ( n34439 , n16378 , n9241 );
    or g40030 ( n5855 , n26561 , n28608 );
    not g40031 ( n19602 , n9637 );
    or g40032 ( n5135 , n39952 , n39804 );
    or g40033 ( n1033 , n19530 , n31578 );
    nor g40034 ( n14304 , n41534 , n37332 );
    not g40035 ( n6322 , n34384 );
    not g40036 ( n37835 , n18251 );
    or g40037 ( n24353 , n37928 , n17729 );
    nor g40038 ( n19482 , n10676 , n8844 );
    and g40039 ( n35831 , n6820 , n34958 );
    or g40040 ( n19315 , n26183 , n880 );
    xnor g40041 ( n34795 , n15617 , n1320 );
    or g40042 ( n1105 , n6415 , n34740 );
    or g40043 ( n40408 , n27321 , n27515 );
    nor g40044 ( n14986 , n9616 , n12379 );
    or g40045 ( n6070 , n37167 , n1645 );
    or g40046 ( n37802 , n3654 , n3031 );
    or g40047 ( n42731 , n12955 , n19585 );
    not g40048 ( n30510 , n17131 );
    not g40049 ( n35813 , n12098 );
    xnor g40050 ( n22207 , n31099 , n19151 );
    or g40051 ( n30991 , n37935 , n41182 );
    and g40052 ( n5256 , n25713 , n13137 );
    or g40053 ( n14254 , n21267 , n3729 );
    or g40054 ( n34859 , n40978 , n20337 );
    or g40055 ( n39300 , n22692 , n35461 );
    or g40056 ( n26466 , n19221 , n25448 );
    xnor g40057 ( n18141 , n12174 , n15378 );
    not g40058 ( n6402 , n31222 );
    nor g40059 ( n16706 , n6313 , n21645 );
    and g40060 ( n23452 , n34386 , n27560 );
    or g40061 ( n31103 , n17744 , n34204 );
    not g40062 ( n42121 , n22110 );
    not g40063 ( n8565 , n16664 );
    not g40064 ( n9525 , n2829 );
    and g40065 ( n15485 , n35924 , n41917 );
    nor g40066 ( n9284 , n4140 , n30354 );
    xnor g40067 ( n258 , n105 , n2155 );
    xnor g40068 ( n1042 , n14864 , n30389 );
    or g40069 ( n7064 , n38168 , n17194 );
    or g40070 ( n25632 , n30619 , n19057 );
    or g40071 ( n19390 , n32855 , n5984 );
    and g40072 ( n12839 , n30642 , n22774 );
    or g40073 ( n1834 , n14597 , n26094 );
    xnor g40074 ( n14466 , n41040 , n9766 );
    xnor g40075 ( n41908 , n480 , n7608 );
    or g40076 ( n31439 , n11882 , n42374 );
    not g40077 ( n8163 , n8209 );
    not g40078 ( n14268 , n38576 );
    xnor g40079 ( n39233 , n20770 , n18076 );
    xnor g40080 ( n11812 , n35727 , n16134 );
    or g40081 ( n40248 , n42871 , n5066 );
    or g40082 ( n20875 , n28149 , n7350 );
    or g40083 ( n40897 , n37600 , n21723 );
    not g40084 ( n3128 , n22506 );
    xnor g40085 ( n1461 , n894 , n36319 );
    or g40086 ( n8333 , n34411 , n11642 );
    xnor g40087 ( n6901 , n34731 , n40947 );
    nor g40088 ( n23828 , n4365 , n7251 );
    or g40089 ( n30694 , n13495 , n30719 );
    and g40090 ( n10549 , n8051 , n38368 );
    nor g40091 ( n24751 , n36823 , n35544 );
    or g40092 ( n42885 , n32200 , n25504 );
    nor g40093 ( n29222 , n20020 , n27115 );
    and g40094 ( n8762 , n42866 , n9587 );
    nor g40095 ( n24790 , n20852 , n21368 );
    nor g40096 ( n7361 , n19519 , n27047 );
    or g40097 ( n34146 , n15109 , n27241 );
    or g40098 ( n33500 , n16116 , n34755 );
    not g40099 ( n10306 , n7532 );
    or g40100 ( n8320 , n41221 , n479 );
    and g40101 ( n17714 , n1084 , n11922 );
    or g40102 ( n31906 , n3679 , n9903 );
    nor g40103 ( n36325 , n25697 , n26799 );
    or g40104 ( n13219 , n20882 , n13718 );
    or g40105 ( n41686 , n36815 , n23957 );
    or g40106 ( n7739 , n15836 , n10250 );
    or g40107 ( n7918 , n2685 , n41641 );
    or g40108 ( n8291 , n25451 , n9986 );
    and g40109 ( n40660 , n21996 , n30831 );
    xnor g40110 ( n17989 , n23867 , n30011 );
    not g40111 ( n5305 , n36853 );
    and g40112 ( n5567 , n21589 , n14710 );
    nor g40113 ( n9537 , n36265 , n26253 );
    and g40114 ( n22762 , n36231 , n26560 );
    xnor g40115 ( n29886 , n38685 , n314 );
    or g40116 ( n797 , n7404 , n42074 );
    or g40117 ( n27233 , n17405 , n14027 );
    xnor g40118 ( n3061 , n30513 , n20816 );
    or g40119 ( n8910 , n15484 , n16636 );
    xnor g40120 ( n32134 , n18840 , n1024 );
    and g40121 ( n1642 , n4244 , n34506 );
    not g40122 ( n31607 , n29475 );
    or g40123 ( n3956 , n26916 , n13012 );
    nor g40124 ( n13993 , n30754 , n24815 );
    or g40125 ( n14584 , n13651 , n38335 );
    not g40126 ( n5675 , n14656 );
    and g40127 ( n41030 , n6060 , n9223 );
    and g40128 ( n33039 , n215 , n29433 );
    and g40129 ( n42077 , n11201 , n24214 );
    or g40130 ( n3644 , n10106 , n24578 );
    not g40131 ( n2292 , n24023 );
    or g40132 ( n11408 , n32809 , n29986 );
    or g40133 ( n25791 , n18686 , n15555 );
    or g40134 ( n33736 , n14707 , n15743 );
    nor g40135 ( n2259 , n23535 , n8420 );
    not g40136 ( n24705 , n36640 );
    and g40137 ( n7687 , n20956 , n1446 );
    not g40138 ( n40487 , n5288 );
    not g40139 ( n29595 , n6372 );
    or g40140 ( n40196 , n35089 , n16100 );
    and g40141 ( n42538 , n9211 , n15694 );
    xnor g40142 ( n42499 , n6962 , n18879 );
    xnor g40143 ( n21845 , n32154 , n11863 );
    and g40144 ( n9824 , n37284 , n28756 );
    and g40145 ( n35859 , n22204 , n8248 );
    or g40146 ( n17885 , n19416 , n33497 );
    xnor g40147 ( n27157 , n11694 , n8664 );
    or g40148 ( n23021 , n15759 , n18236 );
    and g40149 ( n23503 , n5058 , n7298 );
    nor g40150 ( n13833 , n24734 , n12696 );
    or g40151 ( n35972 , n1780 , n5775 );
    or g40152 ( n32761 , n19043 , n22999 );
    xnor g40153 ( n36682 , n25519 , n16398 );
    or g40154 ( n42771 , n5140 , n14442 );
    and g40155 ( n14154 , n36805 , n30227 );
    not g40156 ( n4108 , n3416 );
    not g40157 ( n27552 , n11559 );
    or g40158 ( n24675 , n9329 , n14326 );
    and g40159 ( n41696 , n29723 , n37350 );
    or g40160 ( n25848 , n1105 , n4705 );
    xnor g40161 ( n7236 , n9900 , n37505 );
    xnor g40162 ( n27173 , n35727 , n33337 );
    and g40163 ( n4119 , n8112 , n32342 );
    and g40164 ( n10611 , n8290 , n21121 );
    or g40165 ( n31108 , n17180 , n22631 );
    nor g40166 ( n35677 , n18812 , n28525 );
    nor g40167 ( n20037 , n22117 , n306 );
    xnor g40168 ( n19001 , n566 , n10582 );
    xnor g40169 ( n1534 , n9607 , n36101 );
    xnor g40170 ( n19076 , n5144 , n33316 );
    or g40171 ( n11567 , n17576 , n14276 );
    not g40172 ( n16738 , n38721 );
    and g40173 ( n35673 , n33270 , n27309 );
    or g40174 ( n2162 , n18798 , n38994 );
    or g40175 ( n8124 , n39842 , n40421 );
    or g40176 ( n40307 , n8327 , n10622 );
    or g40177 ( n41802 , n20575 , n40323 );
    or g40178 ( n39784 , n22291 , n38701 );
    or g40179 ( n38568 , n27039 , n41754 );
    not g40180 ( n16841 , n32398 );
    or g40181 ( n19714 , n14432 , n5850 );
    not g40182 ( n34745 , n2239 );
    and g40183 ( n21278 , n23798 , n35967 );
    and g40184 ( n2155 , n11662 , n22959 );
    not g40185 ( n31523 , n36034 );
    nor g40186 ( n41645 , n2199 , n30886 );
    not g40187 ( n7421 , n34330 );
    and g40188 ( n1549 , n29694 , n39818 );
    nor g40189 ( n26252 , n4154 , n10269 );
    xnor g40190 ( n20467 , n105 , n17678 );
    not g40191 ( n22243 , n41847 );
    or g40192 ( n8482 , n5101 , n10496 );
    xnor g40193 ( n2487 , n11436 , n22186 );
    xnor g40194 ( n18297 , n34329 , n1217 );
    or g40195 ( n29360 , n14481 , n35746 );
    xnor g40196 ( n29174 , n10084 , n35843 );
    or g40197 ( n28795 , n32980 , n20256 );
    and g40198 ( n42704 , n38005 , n27436 );
    or g40199 ( n14628 , n9508 , n19445 );
    or g40200 ( n22822 , n13220 , n26520 );
    not g40201 ( n18178 , n34611 );
    nor g40202 ( n23249 , n10828 , n20964 );
    xnor g40203 ( n6313 , n38899 , n34390 );
    or g40204 ( n19059 , n28025 , n34184 );
    and g40205 ( n6041 , n12554 , n7630 );
    and g40206 ( n13313 , n28853 , n41214 );
    xnor g40207 ( n20093 , n21184 , n13012 );
    or g40208 ( n26327 , n10635 , n40379 );
    and g40209 ( n23669 , n16215 , n13906 );
    or g40210 ( n32211 , n12621 , n36476 );
    and g40211 ( n34289 , n20919 , n37781 );
    not g40212 ( n3868 , n42016 );
    xnor g40213 ( n14119 , n39900 , n34563 );
    xnor g40214 ( n34057 , n22161 , n1716 );
    not g40215 ( n4444 , n1319 );
    not g40216 ( n39118 , n17918 );
    or g40217 ( n27009 , n18866 , n19371 );
    not g40218 ( n7980 , n18285 );
    nor g40219 ( n41574 , n28749 , n4964 );
    xnor g40220 ( n21605 , n21534 , n2694 );
    or g40221 ( n22680 , n28526 , n8617 );
    or g40222 ( n12270 , n37771 , n41370 );
    nor g40223 ( n6627 , n34480 , n16901 );
    not g40224 ( n5413 , n32384 );
    or g40225 ( n9112 , n32180 , n39316 );
    or g40226 ( n34058 , n40088 , n18236 );
    not g40227 ( n10676 , n34173 );
    or g40228 ( n41876 , n9508 , n30011 );
    and g40229 ( n5931 , n36307 , n31224 );
    nor g40230 ( n24459 , n9869 , n23117 );
    and g40231 ( n15025 , n40603 , n28851 );
    xnor g40232 ( n24526 , n24991 , n16734 );
    xnor g40233 ( n16775 , n29129 , n20321 );
    or g40234 ( n9845 , n12515 , n12867 );
    or g40235 ( n42319 , n14945 , n27326 );
    or g40236 ( n6410 , n2506 , n31671 );
    xnor g40237 ( n2929 , n23846 , n19846 );
    nor g40238 ( n28494 , n32414 , n10469 );
    or g40239 ( n262 , n29580 , n18495 );
    not g40240 ( n30959 , n18800 );
    or g40241 ( n23527 , n27306 , n32068 );
    and g40242 ( n17187 , n34092 , n7258 );
    not g40243 ( n20566 , n24141 );
    not g40244 ( n5261 , n13979 );
    not g40245 ( n20707 , n31965 );
    and g40246 ( n8355 , n15725 , n2618 );
    or g40247 ( n17020 , n2549 , n30822 );
    not g40248 ( n13447 , n4826 );
    or g40249 ( n17324 , n39671 , n24185 );
    and g40250 ( n40529 , n26454 , n8484 );
    and g40251 ( n31776 , n11420 , n24977 );
    not g40252 ( n5055 , n31557 );
    nor g40253 ( n9218 , n36104 , n41689 );
    xnor g40254 ( n23494 , n3028 , n14707 );
    and g40255 ( n16593 , n35439 , n14789 );
    or g40256 ( n21944 , n14996 , n3021 );
    or g40257 ( n16824 , n8950 , n22398 );
    and g40258 ( n16856 , n37943 , n14424 );
    or g40259 ( n40491 , n4611 , n28256 );
    not g40260 ( n7242 , n14589 );
    and g40261 ( n31603 , n18312 , n6567 );
    or g40262 ( n35888 , n22731 , n41213 );
    and g40263 ( n32130 , n28279 , n6136 );
    not g40264 ( n23109 , n30874 );
    and g40265 ( n1281 , n34595 , n25687 );
    xnor g40266 ( n22659 , n28217 , n5517 );
    or g40267 ( n26127 , n28345 , n33330 );
    nor g40268 ( n26766 , n31518 , n27115 );
    not g40269 ( n34106 , n613 );
    and g40270 ( n36447 , n4334 , n22661 );
    xnor g40271 ( n12349 , n13415 , n40218 );
    and g40272 ( n33580 , n9685 , n17673 );
    xnor g40273 ( n7521 , n2130 , n12061 );
    xnor g40274 ( n35014 , n38955 , n32460 );
    nor g40275 ( n31593 , n18051 , n16081 );
    or g40276 ( n4547 , n32258 , n13701 );
    or g40277 ( n8937 , n34286 , n11709 );
    or g40278 ( n3534 , n1097 , n328 );
    not g40279 ( n35387 , n204 );
    not g40280 ( n24200 , n31775 );
    nor g40281 ( n25084 , n22820 , n38238 );
    nor g40282 ( n4277 , n28553 , n11549 );
    not g40283 ( n40655 , n24825 );
    not g40284 ( n29389 , n140 );
    or g40285 ( n35652 , n15721 , n15827 );
    not g40286 ( n14384 , n42759 );
    or g40287 ( n36554 , n18294 , n3133 );
    nor g40288 ( n7214 , n20707 , n25133 );
    and g40289 ( n8516 , n19299 , n38961 );
    and g40290 ( n32437 , n27717 , n9093 );
    or g40291 ( n23412 , n4959 , n11515 );
    or g40292 ( n32840 , n7525 , n2129 );
    or g40293 ( n39739 , n38317 , n2203 );
    not g40294 ( n12876 , n25105 );
    or g40295 ( n28663 , n21279 , n41684 );
    not g40296 ( n22452 , n30936 );
    not g40297 ( n27153 , n5275 );
    or g40298 ( n19877 , n41961 , n12546 );
    nor g40299 ( n39303 , n2770 , n29847 );
    or g40300 ( n38794 , n39441 , n15306 );
    or g40301 ( n24619 , n38082 , n25318 );
    and g40302 ( n37219 , n17167 , n21715 );
    or g40303 ( n26700 , n36574 , n30165 );
    not g40304 ( n28517 , n26673 );
    not g40305 ( n42393 , n23824 );
    and g40306 ( n41203 , n22763 , n19978 );
    or g40307 ( n37501 , n2469 , n20174 );
    or g40308 ( n12373 , n35276 , n525 );
    or g40309 ( n11173 , n31992 , n13861 );
    not g40310 ( n6294 , n18159 );
    or g40311 ( n39324 , n8415 , n15866 );
    and g40312 ( n38793 , n35872 , n24557 );
    xnor g40313 ( n23567 , n14315 , n18313 );
    nor g40314 ( n19440 , n35297 , n32446 );
    xnor g40315 ( n12773 , n36009 , n22599 );
    and g40316 ( n8659 , n34822 , n9497 );
    not g40317 ( n32711 , n23184 );
    or g40318 ( n39467 , n4033 , n27059 );
    and g40319 ( n2252 , n20487 , n11764 );
    not g40320 ( n27633 , n35841 );
    nor g40321 ( n3511 , n38314 , n26578 );
    not g40322 ( n34017 , n7986 );
    and g40323 ( n28044 , n5735 , n19696 );
    nor g40324 ( n18666 , n28328 , n1899 );
    or g40325 ( n36910 , n310 , n6720 );
    and g40326 ( n31860 , n18503 , n28267 );
    nor g40327 ( n4238 , n17193 , n8602 );
    not g40328 ( n2226 , n35496 );
    nor g40329 ( n16499 , n25657 , n19574 );
    or g40330 ( n26251 , n27884 , n5587 );
    not g40331 ( n12190 , n35759 );
    nor g40332 ( n12330 , n39473 , n1845 );
    or g40333 ( n25682 , n29766 , n16466 );
    not g40334 ( n38196 , n36298 );
    and g40335 ( n30007 , n35828 , n5477 );
    xnor g40336 ( n2165 , n31532 , n6360 );
    or g40337 ( n13133 , n567 , n8874 );
    and g40338 ( n1948 , n6696 , n20372 );
    or g40339 ( n11241 , n21919 , n24927 );
    xnor g40340 ( n21647 , n23058 , n27076 );
    or g40341 ( n5288 , n36813 , n6679 );
    nor g40342 ( n24882 , n42794 , n20628 );
    and g40343 ( n42793 , n20994 , n42303 );
    or g40344 ( n42678 , n15505 , n23787 );
    not g40345 ( n5013 , n15693 );
    not g40346 ( n21767 , n38934 );
    not g40347 ( n2850 , n31620 );
    xnor g40348 ( n17928 , n31099 , n15554 );
    and g40349 ( n13085 , n24404 , n38866 );
    nor g40350 ( n13823 , n23318 , n4847 );
    not g40351 ( n40978 , n16076 );
    not g40352 ( n40210 , n18090 );
    xnor g40353 ( n20019 , n21610 , n6515 );
    nor g40354 ( n25736 , n141 , n6501 );
    not g40355 ( n36153 , n6854 );
    or g40356 ( n26568 , n38621 , n38223 );
    or g40357 ( n10104 , n41516 , n26140 );
    not g40358 ( n21957 , n26358 );
    and g40359 ( n7996 , n33386 , n39440 );
    and g40360 ( n38748 , n24071 , n2934 );
    or g40361 ( n41055 , n19765 , n21697 );
    not g40362 ( n42850 , n18369 );
    xnor g40363 ( n15623 , n21141 , n26478 );
    or g40364 ( n23038 , n42068 , n30224 );
    not g40365 ( n18209 , n21451 );
    or g40366 ( n14334 , n4788 , n9824 );
    or g40367 ( n6860 , n42300 , n26606 );
    or g40368 ( n1103 , n18000 , n27007 );
    not g40369 ( n4908 , n25205 );
    and g40370 ( n35646 , n21406 , n16700 );
    not g40371 ( n23510 , n13523 );
    not g40372 ( n32747 , n38701 );
    xnor g40373 ( n1698 , n42064 , n18978 );
    or g40374 ( n31920 , n29358 , n10654 );
    and g40375 ( n42840 , n30310 , n41183 );
    xnor g40376 ( n15136 , n25552 , n11673 );
    and g40377 ( n22727 , n7455 , n20139 );
    or g40378 ( n12183 , n42798 , n11554 );
    not g40379 ( n38661 , n3140 );
    not g40380 ( n38828 , n39861 );
    and g40381 ( n16237 , n19611 , n35300 );
    and g40382 ( n40712 , n35242 , n6926 );
    or g40383 ( n35114 , n9732 , n12129 );
    nor g40384 ( n35921 , n383 , n2899 );
    not g40385 ( n27575 , n20630 );
    or g40386 ( n11160 , n38323 , n30824 );
    nor g40387 ( n35692 , n16039 , n32798 );
    and g40388 ( n29000 , n35053 , n39009 );
    or g40389 ( n5373 , n35151 , n32194 );
    not g40390 ( n33038 , n20882 );
    or g40391 ( n18371 , n10914 , n6478 );
    or g40392 ( n23062 , n16114 , n25486 );
    or g40393 ( n17737 , n30936 , n1485 );
    or g40394 ( n35957 , n12666 , n13021 );
    or g40395 ( n15805 , n2783 , n26334 );
    and g40396 ( n18927 , n3022 , n692 );
    or g40397 ( n13906 , n14788 , n9455 );
    and g40398 ( n41136 , n7875 , n16674 );
    and g40399 ( n22744 , n12060 , n4434 );
    not g40400 ( n17918 , n10010 );
    nor g40401 ( n15332 , n9035 , n41089 );
    or g40402 ( n29090 , n26996 , n20189 );
    or g40403 ( n34568 , n36240 , n6619 );
    and g40404 ( n15242 , n38989 , n12472 );
    and g40405 ( n24281 , n37089 , n39011 );
    xnor g40406 ( n41807 , n12836 , n15098 );
    nor g40407 ( n38611 , n12864 , n8263 );
    and g40408 ( n35728 , n30012 , n4475 );
    or g40409 ( n20833 , n29239 , n33234 );
    nor g40410 ( n28440 , n32069 , n4854 );
    xnor g40411 ( n35376 , n5041 , n12726 );
    or g40412 ( n5451 , n40331 , n2531 );
    and g40413 ( n12898 , n371 , n26661 );
    and g40414 ( n29673 , n7217 , n32022 );
    xnor g40415 ( n16565 , n38190 , n22382 );
    xnor g40416 ( n15593 , n26440 , n15334 );
    nor g40417 ( n7189 , n42740 , n20062 );
    or g40418 ( n8007 , n7174 , n27531 );
    or g40419 ( n35519 , n17808 , n12165 );
    and g40420 ( n2272 , n40438 , n922 );
    or g40421 ( n38848 , n17985 , n13866 );
    not g40422 ( n17967 , n5594 );
    not g40423 ( n30677 , n19855 );
    not g40424 ( n12266 , n10523 );
    not g40425 ( n26441 , n22303 );
    or g40426 ( n31008 , n38704 , n7660 );
    not g40427 ( n13379 , n30590 );
    xnor g40428 ( n12192 , n1469 , n26665 );
    or g40429 ( n7825 , n37780 , n13765 );
    not g40430 ( n10779 , n12367 );
    or g40431 ( n13271 , n14499 , n40957 );
    nor g40432 ( n39509 , n33981 , n17002 );
    nor g40433 ( n26389 , n33198 , n13262 );
    not g40434 ( n13597 , n8747 );
    not g40435 ( n14507 , n37325 );
    or g40436 ( n10301 , n9765 , n17445 );
    not g40437 ( n15425 , n19605 );
    and g40438 ( n10966 , n38863 , n8328 );
    and g40439 ( n18685 , n12405 , n29828 );
    or g40440 ( n12323 , n42532 , n3856 );
    or g40441 ( n23875 , n33924 , n25077 );
    or g40442 ( n35718 , n34997 , n35636 );
    not g40443 ( n10710 , n33714 );
    nor g40444 ( n34910 , n22473 , n19986 );
    or g40445 ( n19944 , n7092 , n28398 );
    and g40446 ( n13341 , n17660 , n19440 );
    not g40447 ( n18427 , n3428 );
    not g40448 ( n5625 , n1246 );
    and g40449 ( n24771 , n38917 , n5736 );
    or g40450 ( n31706 , n295 , n40494 );
    xnor g40451 ( n27927 , n29854 , n37292 );
    or g40452 ( n23536 , n34527 , n6521 );
    xnor g40453 ( n11236 , n15887 , n35003 );
    xnor g40454 ( n7520 , n31474 , n39304 );
    xnor g40455 ( n32047 , n105 , n33522 );
    xnor g40456 ( n15442 , n784 , n10665 );
    xnor g40457 ( n12752 , n33876 , n9381 );
    and g40458 ( n10378 , n28542 , n15126 );
    xnor g40459 ( n5746 , n34810 , n18893 );
    not g40460 ( n8794 , n26343 );
    and g40461 ( n32719 , n28668 , n42130 );
    or g40462 ( n35202 , n36283 , n279 );
    xnor g40463 ( n17396 , n588 , n31461 );
    and g40464 ( n29443 , n24333 , n35201 );
    and g40465 ( n25598 , n36998 , n31989 );
    and g40466 ( n36621 , n17519 , n42711 );
    and g40467 ( n10223 , n38147 , n12322 );
    or g40468 ( n31398 , n13505 , n24371 );
    or g40469 ( n15575 , n18140 , n10240 );
    nor g40470 ( n22654 , n18093 , n16362 );
    not g40471 ( n12666 , n8081 );
    and g40472 ( n6348 , n13864 , n21587 );
    and g40473 ( n867 , n10342 , n21605 );
    and g40474 ( n22044 , n14720 , n26745 );
    or g40475 ( n2236 , n24053 , n4441 );
    and g40476 ( n32503 , n15699 , n34257 );
    or g40477 ( n27528 , n24872 , n12228 );
    not g40478 ( n24696 , n4945 );
    or g40479 ( n964 , n37771 , n13970 );
    not g40480 ( n41278 , n7888 );
    xnor g40481 ( n25058 , n33253 , n28780 );
    and g40482 ( n35118 , n41583 , n18361 );
    not g40483 ( n35531 , n39581 );
    or g40484 ( n9270 , n31194 , n21807 );
    xnor g40485 ( n18344 , n15742 , n25662 );
    or g40486 ( n21704 , n20995 , n20083 );
    and g40487 ( n25903 , n36855 , n2461 );
    xnor g40488 ( n39143 , n37969 , n35728 );
    and g40489 ( n26549 , n4728 , n891 );
    nor g40490 ( n21569 , n12064 , n1552 );
    not g40491 ( n27385 , n32019 );
    or g40492 ( n36057 , n38463 , n23989 );
    or g40493 ( n38514 , n24018 , n7645 );
    or g40494 ( n8737 , n28097 , n7372 );
    or g40495 ( n4150 , n3745 , n11456 );
    nor g40496 ( n30719 , n23066 , n13541 );
    xnor g40497 ( n35799 , n29189 , n4817 );
    and g40498 ( n14868 , n23093 , n9875 );
    and g40499 ( n711 , n36478 , n7909 );
    xnor g40500 ( n19344 , n7023 , n12163 );
    or g40501 ( n11384 , n20350 , n14569 );
    and g40502 ( n32089 , n22392 , n18729 );
    and g40503 ( n30383 , n26598 , n10305 );
    xnor g40504 ( n26722 , n15706 , n441 );
    not g40505 ( n9627 , n20146 );
    xnor g40506 ( n33061 , n16745 , n33128 );
    nor g40507 ( n1225 , n35318 , n1672 );
    or g40508 ( n32577 , n38489 , n3781 );
    or g40509 ( n15985 , n3443 , n25018 );
    or g40510 ( n8251 , n9192 , n17681 );
    or g40511 ( n12446 , n3876 , n8087 );
    and g40512 ( n20622 , n39912 , n42843 );
    not g40513 ( n39559 , n19651 );
    not g40514 ( n27992 , n7477 );
    and g40515 ( n12252 , n39882 , n9463 );
    and g40516 ( n27783 , n31105 , n17508 );
    or g40517 ( n1230 , n10356 , n16908 );
    and g40518 ( n42119 , n16569 , n32380 );
    nor g40519 ( n22079 , n9168 , n29059 );
    or g40520 ( n22674 , n39709 , n19902 );
    and g40521 ( n29363 , n9092 , n20260 );
    or g40522 ( n3189 , n26523 , n11828 );
    nor g40523 ( n11793 , n28407 , n33479 );
    not g40524 ( n10251 , n30185 );
    nor g40525 ( n15908 , n13643 , n20870 );
    and g40526 ( n25782 , n40938 , n35916 );
    and g40527 ( n26782 , n17328 , n23720 );
    and g40528 ( n37011 , n38145 , n1346 );
    or g40529 ( n39497 , n18672 , n14630 );
    xnor g40530 ( n37816 , n7741 , n28543 );
    and g40531 ( n31336 , n4138 , n25999 );
    or g40532 ( n23093 , n21813 , n35729 );
    and g40533 ( n13536 , n3491 , n1431 );
    and g40534 ( n37939 , n39417 , n28008 );
    not g40535 ( n31122 , n40600 );
    not g40536 ( n37446 , n16552 );
    or g40537 ( n15323 , n11597 , n32256 );
    not g40538 ( n37163 , n40927 );
    and g40539 ( n8523 , n20046 , n13779 );
    xnor g40540 ( n3251 , n9449 , n22878 );
    and g40541 ( n21203 , n5233 , n7317 );
    or g40542 ( n4319 , n587 , n28165 );
    not g40543 ( n29135 , n2018 );
    xnor g40544 ( n1297 , n30830 , n21671 );
    xnor g40545 ( n31611 , n24278 , n22718 );
    and g40546 ( n11774 , n17274 , n6204 );
    xnor g40547 ( n8144 , n31615 , n14100 );
    and g40548 ( n28113 , n28964 , n25841 );
    not g40549 ( n26542 , n3490 );
    and g40550 ( n360 , n40099 , n13196 );
    nor g40551 ( n16464 , n186 , n32024 );
    and g40552 ( n20176 , n29692 , n7161 );
    or g40553 ( n12055 , n40785 , n11604 );
    or g40554 ( n7531 , n972 , n6691 );
    and g40555 ( n30173 , n39666 , n28627 );
    xnor g40556 ( n33324 , n11023 , n11643 );
    or g40557 ( n25227 , n16054 , n20065 );
    not g40558 ( n38556 , n40674 );
    and g40559 ( n6432 , n1394 , n25093 );
    or g40560 ( n7123 , n40229 , n21064 );
    or g40561 ( n12596 , n8563 , n10292 );
    xnor g40562 ( n40988 , n2714 , n8065 );
    and g40563 ( n39966 , n12934 , n32464 );
    and g40564 ( n27798 , n20894 , n9100 );
    and g40565 ( n29842 , n5885 , n12659 );
    and g40566 ( n3719 , n17132 , n5949 );
    and g40567 ( n24221 , n19226 , n10383 );
    or g40568 ( n25333 , n20133 , n3905 );
    or g40569 ( n14633 , n34609 , n9713 );
    or g40570 ( n11943 , n40611 , n1479 );
    and g40571 ( n27431 , n28052 , n24412 );
    nor g40572 ( n27725 , n12389 , n15440 );
    not g40573 ( n30358 , n3000 );
    not g40574 ( n35678 , n6054 );
    or g40575 ( n31133 , n16155 , n42850 );
    xnor g40576 ( n37691 , n25985 , n12802 );
    not g40577 ( n29577 , n7188 );
    xnor g40578 ( n42169 , n29740 , n18132 );
    xnor g40579 ( n30032 , n34585 , n5601 );
    and g40580 ( n34967 , n31726 , n22882 );
    xnor g40581 ( n32143 , n33416 , n19682 );
    xnor g40582 ( n42312 , n36998 , n33376 );
    and g40583 ( n15904 , n38948 , n2796 );
    and g40584 ( n40983 , n31904 , n13131 );
    or g40585 ( n36187 , n2742 , n30749 );
    or g40586 ( n39190 , n966 , n17090 );
    or g40587 ( n19967 , n26592 , n42448 );
    nor g40588 ( n304 , n27328 , n559 );
    nor g40589 ( n21676 , n2734 , n39477 );
    not g40590 ( n41538 , n26171 );
    and g40591 ( n20831 , n34689 , n15304 );
    or g40592 ( n7310 , n3548 , n4660 );
    and g40593 ( n13745 , n12779 , n16704 );
    xnor g40594 ( n7121 , n41697 , n95 );
    or g40595 ( n42597 , n39844 , n28143 );
    or g40596 ( n3650 , n39439 , n21583 );
    or g40597 ( n4139 , n3363 , n11177 );
    not g40598 ( n28125 , n26872 );
    or g40599 ( n40334 , n41074 , n36644 );
    xnor g40600 ( n8249 , n40086 , n20899 );
    and g40601 ( n30274 , n13697 , n20361 );
    or g40602 ( n31269 , n131 , n14373 );
    nor g40603 ( n23972 , n31078 , n34867 );
    and g40604 ( n123 , n10303 , n31868 );
    or g40605 ( n24492 , n12051 , n29865 );
    nor g40606 ( n18508 , n42146 , n424 );
    not g40607 ( n36397 , n23309 );
    and g40608 ( n41186 , n30033 , n29736 );
    or g40609 ( n23418 , n5680 , n6719 );
    or g40610 ( n12008 , n8494 , n5964 );
    nor g40611 ( n1189 , n24364 , n23461 );
    xnor g40612 ( n30073 , n30492 , n17326 );
    not g40613 ( n3759 , n29560 );
    or g40614 ( n17004 , n35674 , n17595 );
    xnor g40615 ( n31592 , n39532 , n32430 );
    or g40616 ( n31544 , n33691 , n22593 );
    not g40617 ( n19251 , n8317 );
    or g40618 ( n30524 , n24259 , n34728 );
    or g40619 ( n40843 , n23139 , n6588 );
    or g40620 ( n10154 , n1788 , n12298 );
    nor g40621 ( n17670 , n8922 , n14544 );
    and g40622 ( n34549 , n16754 , n9949 );
    not g40623 ( n10017 , n15831 );
    nor g40624 ( n17991 , n6995 , n41626 );
    or g40625 ( n27821 , n18022 , n42218 );
    nor g40626 ( n38164 , n13657 , n17959 );
    or g40627 ( n1951 , n36870 , n3072 );
    or g40628 ( n41512 , n34586 , n20312 );
    or g40629 ( n36278 , n7423 , n40151 );
    not g40630 ( n5795 , n22306 );
    xnor g40631 ( n22874 , n36444 , n23989 );
    and g40632 ( n38505 , n29409 , n12496 );
    or g40633 ( n34595 , n1407 , n21372 );
    or g40634 ( n13072 , n166 , n36214 );
    or g40635 ( n18325 , n15303 , n13560 );
    xnor g40636 ( n2468 , n12146 , n28130 );
    not g40637 ( n7492 , n4722 );
    xnor g40638 ( n17810 , n31962 , n39613 );
    or g40639 ( n35988 , n10103 , n40648 );
    xnor g40640 ( n9373 , n2227 , n10598 );
    or g40641 ( n19502 , n32550 , n5128 );
    and g40642 ( n13310 , n24325 , n41675 );
    or g40643 ( n29270 , n14875 , n36071 );
    and g40644 ( n24185 , n9242 , n32249 );
    nor g40645 ( n29339 , n29424 , n39305 );
    or g40646 ( n23155 , n7378 , n25312 );
    or g40647 ( n22295 , n15116 , n34296 );
    or g40648 ( n26997 , n18662 , n20621 );
    and g40649 ( n36067 , n18145 , n33299 );
    xnor g40650 ( n27972 , n22128 , n41097 );
    xnor g40651 ( n33225 , n25601 , n39338 );
    and g40652 ( n23881 , n29794 , n12118 );
    nor g40653 ( n19457 , n12225 , n30889 );
    and g40654 ( n19110 , n36591 , n36753 );
    and g40655 ( n32943 , n23639 , n26033 );
    xnor g40656 ( n14231 , n29740 , n15540 );
    not g40657 ( n6377 , n39095 );
    not g40658 ( n16872 , n17764 );
    and g40659 ( n9646 , n1886 , n37458 );
    nor g40660 ( n27919 , n34097 , n4248 );
    and g40661 ( n29240 , n35552 , n2307 );
    nor g40662 ( n14141 , n6574 , n23996 );
    nor g40663 ( n34486 , n22625 , n4495 );
    and g40664 ( n23314 , n24414 , n3200 );
    nor g40665 ( n6925 , n17698 , n12195 );
    or g40666 ( n12097 , n34993 , n17895 );
    xnor g40667 ( n22641 , n20647 , n38930 );
    or g40668 ( n27014 , n16598 , n36504 );
    not g40669 ( n36315 , n31336 );
    or g40670 ( n31639 , n7223 , n26554 );
    or g40671 ( n2059 , n30207 , n22239 );
    or g40672 ( n17837 , n18835 , n11118 );
    and g40673 ( n27567 , n34600 , n33645 );
    and g40674 ( n7493 , n9526 , n1744 );
    or g40675 ( n13935 , n15282 , n23335 );
    or g40676 ( n22189 , n12011 , n117 );
    and g40677 ( n32513 , n21356 , n33958 );
    or g40678 ( n3865 , n40110 , n2218 );
    nor g40679 ( n5524 , n32069 , n4839 );
    and g40680 ( n27374 , n26756 , n8001 );
    and g40681 ( n31218 , n39005 , n13578 );
    not g40682 ( n40391 , n2562 );
    and g40683 ( n23618 , n18423 , n33399 );
    and g40684 ( n7831 , n32507 , n4592 );
    or g40685 ( n17633 , n6929 , n37037 );
    and g40686 ( n32923 , n40108 , n2816 );
    xnor g40687 ( n10352 , n23322 , n34119 );
    not g40688 ( n42143 , n7518 );
    not g40689 ( n27682 , n9158 );
    not g40690 ( n24734 , n1419 );
    and g40691 ( n23542 , n36192 , n39325 );
    or g40692 ( n35380 , n734 , n41405 );
    or g40693 ( n39650 , n9145 , n29840 );
    or g40694 ( n36997 , n15053 , n40259 );
    xnor g40695 ( n38097 , n40861 , n38127 );
    not g40696 ( n25382 , n13540 );
    and g40697 ( n19376 , n27641 , n34776 );
    or g40698 ( n14100 , n805 , n19736 );
    xnor g40699 ( n3499 , n36009 , n37065 );
    and g40700 ( n21910 , n27066 , n5715 );
    xnor g40701 ( n34355 , n34562 , n38461 );
    or g40702 ( n9204 , n19084 , n3503 );
    or g40703 ( n34421 , n23192 , n19159 );
    or g40704 ( n109 , n36200 , n24501 );
    xnor g40705 ( n21639 , n21495 , n15984 );
    or g40706 ( n4204 , n15307 , n39536 );
    xnor g40707 ( n41917 , n5759 , n8324 );
    or g40708 ( n6382 , n31405 , n24110 );
    and g40709 ( n28117 , n13546 , n4134 );
    or g40710 ( n19751 , n28785 , n29431 );
    and g40711 ( n32174 , n19172 , n15679 );
    or g40712 ( n29004 , n22562 , n19140 );
    not g40713 ( n9511 , n27205 );
    xnor g40714 ( n36196 , n28221 , n33981 );
    nor g40715 ( n2040 , n32265 , n26810 );
    and g40716 ( n10603 , n25901 , n19204 );
    or g40717 ( n16041 , n8047 , n27702 );
    not g40718 ( n24800 , n40136 );
    or g40719 ( n33814 , n38879 , n711 );
    and g40720 ( n796 , n37673 , n29463 );
    or g40721 ( n10938 , n36972 , n28253 );
    not g40722 ( n24879 , n29715 );
    nor g40723 ( n37470 , n13476 , n40204 );
    nor g40724 ( n35096 , n25588 , n16684 );
    and g40725 ( n19446 , n29907 , n10951 );
    and g40726 ( n9451 , n6994 , n29428 );
    or g40727 ( n13617 , n641 , n644 );
    or g40728 ( n10144 , n36195 , n28239 );
    and g40729 ( n28809 , n6895 , n42579 );
    nor g40730 ( n42314 , n19008 , n15761 );
    and g40731 ( n19402 , n23351 , n16956 );
    xnor g40732 ( n18417 , n2317 , n20328 );
    not g40733 ( n39896 , n36490 );
    and g40734 ( n25453 , n30731 , n6100 );
    and g40735 ( n34505 , n10122 , n11959 );
    nor g40736 ( n40200 , n5953 , n18705 );
    xnor g40737 ( n3621 , n5144 , n32123 );
    nor g40738 ( n40044 , n4105 , n38784 );
    or g40739 ( n6089 , n37308 , n35635 );
    or g40740 ( n9625 , n3954 , n26023 );
    or g40741 ( n38930 , n17446 , n12846 );
    not g40742 ( n14379 , n354 );
    and g40743 ( n26234 , n22644 , n19640 );
    xnor g40744 ( n7358 , n30549 , n27616 );
    xnor g40745 ( n24774 , n1863 , n6672 );
    and g40746 ( n38603 , n42854 , n22265 );
    or g40747 ( n5936 , n35138 , n17059 );
    nor g40748 ( n20837 , n19033 , n41114 );
    and g40749 ( n22199 , n37066 , n10776 );
    nor g40750 ( n7202 , n18143 , n16677 );
    or g40751 ( n14757 , n24199 , n31671 );
    or g40752 ( n26830 , n2507 , n9700 );
    or g40753 ( n7440 , n1917 , n35149 );
    not g40754 ( n23211 , n26515 );
    or g40755 ( n37491 , n7375 , n16136 );
    and g40756 ( n2479 , n27173 , n10261 );
    or g40757 ( n29483 , n7839 , n11968 );
    xnor g40758 ( n25312 , n5043 , n42593 );
    nor g40759 ( n16443 , n24833 , n17095 );
    nor g40760 ( n35895 , n29408 , n2944 );
    or g40761 ( n4978 , n33031 , n19984 );
    or g40762 ( n41490 , n1320 , n16150 );
    or g40763 ( n32081 , n29970 , n34728 );
    or g40764 ( n73 , n34762 , n13865 );
    and g40765 ( n36179 , n10994 , n1277 );
    nor g40766 ( n7660 , n28792 , n25605 );
    or g40767 ( n14588 , n38450 , n2296 );
    and g40768 ( n34079 , n33880 , n36232 );
    xnor g40769 ( n20890 , n24505 , n27192 );
    not g40770 ( n32170 , n31815 );
    nor g40771 ( n38821 , n36441 , n11005 );
    or g40772 ( n17278 , n36945 , n40882 );
    nor g40773 ( n11090 , n22861 , n36676 );
    or g40774 ( n14593 , n3282 , n529 );
    and g40775 ( n20118 , n13109 , n40897 );
    and g40776 ( n31898 , n17939 , n142 );
    and g40777 ( n15374 , n7136 , n16385 );
    not g40778 ( n21309 , n39082 );
    xnor g40779 ( n12338 , n21192 , n10180 );
    not g40780 ( n26540 , n26463 );
    and g40781 ( n12559 , n33109 , n36229 );
    and g40782 ( n22733 , n17878 , n35421 );
    xnor g40783 ( n9906 , n28541 , n23496 );
    or g40784 ( n11121 , n22090 , n32180 );
    xnor g40785 ( n21507 , n35813 , n25851 );
    and g40786 ( n9265 , n20910 , n12916 );
    or g40787 ( n28277 , n36211 , n39250 );
    xnor g40788 ( n18755 , n18530 , n27507 );
    or g40789 ( n5448 , n13699 , n30259 );
    and g40790 ( n30875 , n13581 , n38501 );
    not g40791 ( n19119 , n25936 );
    xnor g40792 ( n6568 , n502 , n38859 );
    or g40793 ( n26923 , n1644 , n13554 );
    or g40794 ( n15496 , n15037 , n23206 );
    and g40795 ( n18847 , n31319 , n31282 );
    not g40796 ( n17563 , n23948 );
    or g40797 ( n28040 , n17568 , n28643 );
    nor g40798 ( n30612 , n22577 , n15907 );
    not g40799 ( n18142 , n22009 );
    or g40800 ( n19425 , n16530 , n9107 );
    or g40801 ( n28412 , n8284 , n34267 );
    not g40802 ( n23944 , n19952 );
    or g40803 ( n8330 , n13157 , n30274 );
    or g40804 ( n22653 , n20709 , n4462 );
    xnor g40805 ( n14273 , n42277 , n21228 );
    and g40806 ( n6765 , n3611 , n13434 );
    nor g40807 ( n23315 , n28636 , n34663 );
    and g40808 ( n33946 , n35806 , n33116 );
    not g40809 ( n485 , n2103 );
    and g40810 ( n26729 , n15330 , n30388 );
    or g40811 ( n9631 , n38213 , n10491 );
    xnor g40812 ( n21963 , n10226 , n12886 );
    or g40813 ( n38092 , n11964 , n36157 );
    or g40814 ( n12971 , n7118 , n10559 );
    not g40815 ( n13921 , n2135 );
    or g40816 ( n23248 , n23462 , n12025 );
    not g40817 ( n5608 , n4163 );
    not g40818 ( n27257 , n41427 );
    nor g40819 ( n9258 , n25709 , n21613 );
    not g40820 ( n23572 , n36154 );
    and g40821 ( n7783 , n2168 , n21758 );
    and g40822 ( n30578 , n28712 , n38455 );
    not g40823 ( n5124 , n19735 );
    nor g40824 ( n20757 , n14530 , n13115 );
    and g40825 ( n22945 , n18175 , n6344 );
    not g40826 ( n17511 , n18008 );
    or g40827 ( n32053 , n30473 , n17894 );
    or g40828 ( n3545 , n16530 , n15074 );
    or g40829 ( n35654 , n20286 , n35269 );
    and g40830 ( n35431 , n25532 , n6805 );
    and g40831 ( n467 , n29450 , n1553 );
    or g40832 ( n9227 , n1275 , n41215 );
    and g40833 ( n4853 , n39901 , n33150 );
    not g40834 ( n24778 , n33726 );
    or g40835 ( n19634 , n27661 , n1387 );
    or g40836 ( n20348 , n18885 , n9926 );
    and g40837 ( n33473 , n1298 , n27095 );
    or g40838 ( n19699 , n26172 , n6872 );
    not g40839 ( n26565 , n19248 );
    and g40840 ( n17362 , n2405 , n4498 );
    xnor g40841 ( n7388 , n22940 , n35716 );
    and g40842 ( n10878 , n10628 , n23208 );
    not g40843 ( n7617 , n31486 );
    nor g40844 ( n11613 , n30189 , n13598 );
    or g40845 ( n27717 , n35879 , n25161 );
    and g40846 ( n12084 , n23822 , n872 );
    and g40847 ( n32580 , n9104 , n2138 );
    xnor g40848 ( n28288 , n6760 , n21388 );
    and g40849 ( n15173 , n12088 , n5830 );
    xnor g40850 ( n7000 , n8194 , n40306 );
    nor g40851 ( n9679 , n16649 , n15351 );
    nor g40852 ( n9735 , n24819 , n37454 );
    and g40853 ( n19397 , n41617 , n15627 );
    nor g40854 ( n862 , n38789 , n16268 );
    xnor g40855 ( n1731 , n38749 , n25651 );
    and g40856 ( n17679 , n23252 , n17635 );
    nor g40857 ( n29155 , n33981 , n3562 );
    or g40858 ( n31921 , n11431 , n35374 );
    or g40859 ( n39130 , n12415 , n4625 );
    nor g40860 ( n641 , n39324 , n20061 );
    or g40861 ( n42279 , n2987 , n17173 );
    nor g40862 ( n12140 , n42436 , n17143 );
    not g40863 ( n27898 , n16010 );
    not g40864 ( n303 , n1868 );
    or g40865 ( n28470 , n16993 , n38175 );
    xnor g40866 ( n36056 , n29057 , n40746 );
    and g40867 ( n28206 , n15966 , n40569 );
    or g40868 ( n34417 , n26448 , n37625 );
    or g40869 ( n6870 , n32389 , n24436 );
    or g40870 ( n41640 , n24874 , n37045 );
    or g40871 ( n29487 , n14029 , n12456 );
    nor g40872 ( n11996 , n42441 , n34498 );
    and g40873 ( n22676 , n37658 , n5069 );
    or g40874 ( n35825 , n2193 , n2949 );
    and g40875 ( n13158 , n21130 , n27514 );
    xnor g40876 ( n21208 , n37436 , n12477 );
    or g40877 ( n12512 , n15095 , n33178 );
    or g40878 ( n26661 , n2563 , n15342 );
    or g40879 ( n3913 , n7073 , n39735 );
    not g40880 ( n36372 , n30851 );
    xnor g40881 ( n185 , n34735 , n1653 );
    and g40882 ( n22667 , n13344 , n35236 );
    and g40883 ( n18455 , n29386 , n42151 );
    not g40884 ( n34691 , n1743 );
    nor g40885 ( n27096 , n25547 , n39459 );
    not g40886 ( n6063 , n15916 );
    or g40887 ( n39842 , n42502 , n22409 );
    nor g40888 ( n21960 , n15409 , n16234 );
    not g40889 ( n21170 , n16702 );
    or g40890 ( n9907 , n9414 , n18602 );
    nor g40891 ( n28610 , n9235 , n29024 );
    and g40892 ( n15775 , n37078 , n37126 );
    or g40893 ( n13149 , n40419 , n6162 );
    not g40894 ( n33596 , n25836 );
    and g40895 ( n37232 , n22416 , n41141 );
    not g40896 ( n24898 , n26620 );
    or g40897 ( n18391 , n13536 , n33074 );
    xnor g40898 ( n28649 , n4060 , n41919 );
    and g40899 ( n23715 , n21941 , n13465 );
    xnor g40900 ( n38673 , n33189 , n11788 );
    xnor g40901 ( n25384 , n11436 , n17153 );
    or g40902 ( n22227 , n38107 , n15233 );
    xnor g40903 ( n42295 , n24997 , n34898 );
    and g40904 ( n32922 , n9271 , n11155 );
    nor g40905 ( n21363 , n39266 , n40303 );
    and g40906 ( n17021 , n11804 , n21464 );
    not g40907 ( n31321 , n18024 );
    xnor g40908 ( n35837 , n27734 , n7747 );
    or g40909 ( n32746 , n7356 , n21571 );
    not g40910 ( n12220 , n36521 );
    or g40911 ( n25083 , n13367 , n10755 );
    and g40912 ( n7534 , n3181 , n39485 );
    xnor g40913 ( n21412 , n36009 , n27851 );
    or g40914 ( n1748 , n27311 , n32488 );
    or g40915 ( n40394 , n33191 , n10136 );
    or g40916 ( n13272 , n8954 , n22489 );
    not g40917 ( n16586 , n499 );
    xnor g40918 ( n32422 , n784 , n13786 );
    or g40919 ( n37142 , n6510 , n40413 );
    not g40920 ( n19192 , n42452 );
    or g40921 ( n23036 , n22379 , n1857 );
    or g40922 ( n32343 , n32100 , n15903 );
    xnor g40923 ( n35563 , n13444 , n26301 );
    or g40924 ( n8509 , n39327 , n10976 );
    not g40925 ( n37705 , n15313 );
    or g40926 ( n4857 , n24595 , n24263 );
    not g40927 ( n13968 , n26383 );
    and g40928 ( n31234 , n18260 , n25919 );
    or g40929 ( n28845 , n3056 , n29583 );
    xnor g40930 ( n13204 , n3822 , n31330 );
    or g40931 ( n24100 , n26887 , n14944 );
    not g40932 ( n17932 , n23341 );
    nor g40933 ( n5840 , n28333 , n12803 );
    nor g40934 ( n20916 , n4174 , n18253 );
    or g40935 ( n38480 , n30896 , n11808 );
    nor g40936 ( n33612 , n17193 , n17506 );
    or g40937 ( n3025 , n40071 , n28253 );
    or g40938 ( n15515 , n30395 , n18207 );
    nor g40939 ( n42726 , n3795 , n33922 );
    or g40940 ( n34781 , n11640 , n16694 );
    not g40941 ( n22861 , n5552 );
    or g40942 ( n32099 , n28551 , n36812 );
    and g40943 ( n17585 , n17989 , n10552 );
    or g40944 ( n37887 , n9015 , n32203 );
    or g40945 ( n23050 , n49 , n4026 );
    and g40946 ( n13279 , n29001 , n1420 );
    nor g40947 ( n34533 , n17193 , n18428 );
    xnor g40948 ( n8391 , n9751 , n33381 );
    or g40949 ( n28324 , n35129 , n34594 );
    xnor g40950 ( n27422 , n23947 , n3736 );
    or g40951 ( n10201 , n41722 , n42586 );
    or g40952 ( n35560 , n24382 , n39408 );
    xnor g40953 ( n15579 , n40617 , n15409 );
    xnor g40954 ( n8934 , n39704 , n37518 );
    or g40955 ( n2049 , n41961 , n23224 );
    not g40956 ( n7568 , n31145 );
    nor g40957 ( n41052 , n28782 , n5879 );
    or g40958 ( n4980 , n22652 , n425 );
    or g40959 ( n15240 , n16941 , n36052 );
    and g40960 ( n21552 , n40866 , n14627 );
    and g40961 ( n6826 , n14041 , n20642 );
    not g40962 ( n40278 , n30244 );
    xnor g40963 ( n31547 , n40380 , n4140 );
    xnor g40964 ( n22787 , n19116 , n40480 );
    not g40965 ( n19848 , n21881 );
    nor g40966 ( n7653 , n31992 , n25804 );
    and g40967 ( n36095 , n5267 , n11584 );
    not g40968 ( n15753 , n17328 );
    not g40969 ( n3410 , n17301 );
    not g40970 ( n2561 , n24096 );
    or g40971 ( n37542 , n930 , n37263 );
    and g40972 ( n32147 , n7248 , n33844 );
    nor g40973 ( n29136 , n1507 , n8447 );
    nor g40974 ( n3370 , n35288 , n12162 );
    not g40975 ( n7839 , n3085 );
    nor g40976 ( n27228 , n13474 , n31773 );
    or g40977 ( n15739 , n5508 , n3681 );
    not g40978 ( n31134 , n21550 );
    or g40979 ( n13986 , n39056 , n36687 );
    not g40980 ( n8900 , n28755 );
    nor g40981 ( n36559 , n18526 , n26878 );
    or g40982 ( n12092 , n3764 , n33437 );
    not g40983 ( n16821 , n35487 );
    or g40984 ( n33255 , n21993 , n35840 );
    nor g40985 ( n35628 , n41793 , n18290 );
    xnor g40986 ( n2381 , n2342 , n4458 );
    or g40987 ( n10951 , n35234 , n31131 );
    and g40988 ( n3587 , n22094 , n12615 );
    xnor g40989 ( n30099 , n24136 , n30574 );
    or g40990 ( n21705 , n35534 , n31827 );
    and g40991 ( n13786 , n27571 , n4576 );
    not g40992 ( n17723 , n4971 );
    or g40993 ( n11861 , n5671 , n13466 );
    nor g40994 ( n3421 , n25976 , n16049 );
    and g40995 ( n4585 , n39979 , n42472 );
    not g40996 ( n27150 , n25355 );
    and g40997 ( n19724 , n16107 , n36039 );
    not g40998 ( n41758 , n25892 );
    not g40999 ( n30546 , n8523 );
    and g41000 ( n21243 , n30009 , n17653 );
    or g41001 ( n37844 , n26869 , n11321 );
    or g41002 ( n4030 , n21254 , n21234 );
    or g41003 ( n41477 , n27447 , n20461 );
    or g41004 ( n6253 , n39026 , n36213 );
    or g41005 ( n20181 , n20174 , n149 );
    and g41006 ( n16066 , n22720 , n30075 );
    or g41007 ( n8525 , n322 , n33941 );
    not g41008 ( n41703 , n36334 );
    or g41009 ( n36551 , n1715 , n40386 );
    or g41010 ( n42093 , n16490 , n37733 );
    or g41011 ( n37236 , n17442 , n37804 );
    or g41012 ( n16806 , n6315 , n12947 );
    not g41013 ( n1379 , n37032 );
    or g41014 ( n42647 , n26549 , n5813 );
    not g41015 ( n4386 , n15992 );
    not g41016 ( n36296 , n2932 );
    not g41017 ( n17381 , n33083 );
    not g41018 ( n3764 , n6557 );
    and g41019 ( n15689 , n13139 , n6336 );
    and g41020 ( n27372 , n27000 , n42720 );
    or g41021 ( n42278 , n25478 , n2304 );
    and g41022 ( n37720 , n22860 , n8836 );
    xnor g41023 ( n40687 , n12146 , n33113 );
    nor g41024 ( n29943 , n32084 , n26773 );
    or g41025 ( n16672 , n40409 , n9580 );
    or g41026 ( n22836 , n33256 , n12152 );
    and g41027 ( n7785 , n39917 , n30982 );
    xnor g41028 ( n12148 , n105 , n24322 );
    not g41029 ( n28228 , n8139 );
    xnor g41030 ( n36165 , n29740 , n39781 );
    nor g41031 ( n20657 , n7356 , n37154 );
    and g41032 ( n7833 , n40069 , n26284 );
    or g41033 ( n12076 , n20866 , n21165 );
    or g41034 ( n9861 , n27311 , n23530 );
    not g41035 ( n8696 , n40614 );
    or g41036 ( n23874 , n32356 , n35231 );
    or g41037 ( n33474 , n10345 , n256 );
    nor g41038 ( n39241 , n39035 , n1128 );
    not g41039 ( n39302 , n19019 );
    xnor g41040 ( n32590 , n23867 , n29254 );
    or g41041 ( n4246 , n34648 , n4564 );
    or g41042 ( n13132 , n25142 , n29874 );
    or g41043 ( n8520 , n36500 , n16843 );
    and g41044 ( n38817 , n14390 , n1142 );
    and g41045 ( n732 , n15941 , n8500 );
    and g41046 ( n11796 , n14285 , n13708 );
    not g41047 ( n7375 , n42710 );
    not g41048 ( n6754 , n42554 );
    and g41049 ( n16016 , n14331 , n31787 );
    or g41050 ( n7528 , n24588 , n6119 );
    or g41051 ( n42721 , n11562 , n14728 );
    not g41052 ( n22582 , n16750 );
    not g41053 ( n39764 , n22009 );
    or g41054 ( n12935 , n38389 , n23309 );
    and g41055 ( n40857 , n23227 , n30753 );
    nor g41056 ( n37496 , n23697 , n2541 );
    xnor g41057 ( n32414 , n24210 , n21857 );
    or g41058 ( n20919 , n18389 , n1630 );
    or g41059 ( n27474 , n33760 , n34010 );
    nor g41060 ( n31032 , n13736 , n19988 );
    or g41061 ( n41307 , n27848 , n40323 );
    or g41062 ( n3180 , n34390 , n33775 );
    or g41063 ( n12329 , n9370 , n29788 );
    or g41064 ( n613 , n34603 , n18057 );
    or g41065 ( n24086 , n32863 , n12351 );
    nor g41066 ( n42882 , n8842 , n40980 );
    or g41067 ( n19279 , n7575 , n41891 );
    and g41068 ( n6990 , n16542 , n40165 );
    nor g41069 ( n24032 , n35042 , n9120 );
    and g41070 ( n396 , n30144 , n14405 );
    or g41071 ( n682 , n24454 , n32437 );
    xnor g41072 ( n28839 , n141 , n19632 );
    or g41073 ( n35903 , n4744 , n12998 );
    and g41074 ( n15335 , n32128 , n24120 );
    or g41075 ( n29460 , n3531 , n22180 );
    or g41076 ( n16375 , n39826 , n28487 );
    not g41077 ( n37811 , n3898 );
    not g41078 ( n16236 , n30054 );
    and g41079 ( n20016 , n35323 , n40562 );
    or g41080 ( n24707 , n36437 , n36658 );
    or g41081 ( n17554 , n14308 , n21761 );
    xnor g41082 ( n7530 , n19514 , n10719 );
    xnor g41083 ( n11880 , n20382 , n4140 );
    and g41084 ( n22050 , n37966 , n29860 );
    nor g41085 ( n39430 , n32669 , n22368 );
    or g41086 ( n8576 , n12459 , n31156 );
    and g41087 ( n12416 , n40759 , n9373 );
    not g41088 ( n32852 , n38580 );
    or g41089 ( n40690 , n28407 , n6436 );
    and g41090 ( n12299 , n10218 , n27854 );
    not g41091 ( n20860 , n192 );
    or g41092 ( n4057 , n41329 , n8735 );
    not g41093 ( n26061 , n28214 );
    xnor g41094 ( n12536 , n9250 , n22988 );
    nor g41095 ( n34188 , n31088 , n4826 );
    or g41096 ( n25099 , n40271 , n29184 );
    and g41097 ( n22559 , n1621 , n38988 );
    or g41098 ( n7101 , n5081 , n11750 );
    and g41099 ( n16709 , n32836 , n22195 );
    or g41100 ( n38329 , n3555 , n33718 );
    not g41101 ( n2548 , n273 );
    or g41102 ( n12905 , n8345 , n6474 );
    not g41103 ( n1734 , n16506 );
    and g41104 ( n8019 , n6741 , n35446 );
    xnor g41105 ( n3663 , n784 , n10333 );
    nor g41106 ( n2107 , n19580 , n5042 );
    and g41107 ( n10754 , n2350 , n34122 );
    not g41108 ( n27555 , n27463 );
    or g41109 ( n15283 , n36203 , n35474 );
    not g41110 ( n22947 , n4855 );
    or g41111 ( n14570 , n11417 , n41448 );
    or g41112 ( n32882 , n8847 , n16995 );
    not g41113 ( n5123 , n7347 );
    or g41114 ( n30679 , n40663 , n38142 );
    or g41115 ( n26918 , n29831 , n9356 );
    and g41116 ( n12527 , n21735 , n5890 );
    or g41117 ( n35462 , n11052 , n39954 );
    not g41118 ( n37495 , n7672 );
    or g41119 ( n8885 , n19811 , n2617 );
    or g41120 ( n34144 , n15185 , n17614 );
    not g41121 ( n37020 , n9344 );
    or g41122 ( n5045 , n15244 , n27628 );
    or g41123 ( n17223 , n18866 , n33254 );
    or g41124 ( n11840 , n9970 , n21778 );
    not g41125 ( n328 , n25345 );
    not g41126 ( n39100 , n19007 );
    and g41127 ( n33217 , n21878 , n28798 );
    or g41128 ( n31481 , n31432 , n29558 );
    or g41129 ( n4583 , n41534 , n17559 );
    xnor g41130 ( n9465 , n22879 , n5839 );
    not g41131 ( n22797 , n12578 );
    and g41132 ( n1459 , n41261 , n39203 );
    nor g41133 ( n7575 , n36598 , n33426 );
    or g41134 ( n17219 , n12619 , n25451 );
    or g41135 ( n1278 , n20031 , n6109 );
    or g41136 ( n24919 , n12756 , n14501 );
    and g41137 ( n7295 , n17117 , n30804 );
    or g41138 ( n1284 , n17827 , n39814 );
    not g41139 ( n15396 , n31075 );
    xnor g41140 ( n31564 , n31989 , n19450 );
    or g41141 ( n31612 , n731 , n20198 );
    not g41142 ( n32814 , n40531 );
    and g41143 ( n2542 , n38831 , n16019 );
    not g41144 ( n23040 , n26575 );
    and g41145 ( n15791 , n35122 , n13410 );
    or g41146 ( n24342 , n38529 , n33858 );
    not g41147 ( n26964 , n13696 );
    nor g41148 ( n34161 , n22625 , n22014 );
    and g41149 ( n31068 , n36876 , n28719 );
    or g41150 ( n31494 , n25808 , n25504 );
    nor g41151 ( n11490 , n21824 , n16869 );
    or g41152 ( n14572 , n25588 , n42195 );
    or g41153 ( n29599 , n32137 , n27981 );
    nor g41154 ( n19655 , n16830 , n29720 );
    and g41155 ( n2704 , n28201 , n23464 );
    and g41156 ( n19151 , n27472 , n42126 );
    not g41157 ( n13491 , n19035 );
    or g41158 ( n29515 , n19041 , n10945 );
    xnor g41159 ( n37950 , n7417 , n17744 );
    not g41160 ( n28404 , n13784 );
    nor g41161 ( n13532 , n535 , n30637 );
    or g41162 ( n7955 , n40033 , n42220 );
    xnor g41163 ( n41467 , n453 , n12371 );
    and g41164 ( n7188 , n14660 , n31588 );
    or g41165 ( n31394 , n15707 , n17858 );
    or g41166 ( n2240 , n6960 , n2863 );
    and g41167 ( n16426 , n34271 , n38015 );
    or g41168 ( n32850 , n35500 , n9315 );
    or g41169 ( n23976 , n35223 , n8429 );
    not g41170 ( n25097 , n33585 );
    or g41171 ( n3904 , n3583 , n2554 );
    not g41172 ( n30768 , n40927 );
    and g41173 ( n11685 , n12944 , n34088 );
    or g41174 ( n7024 , n512 , n7129 );
    or g41175 ( n26398 , n31261 , n16673 );
    not g41176 ( n22454 , n26749 );
    nor g41177 ( n32141 , n24404 , n38866 );
    or g41178 ( n23401 , n30044 , n17726 );
    or g41179 ( n5443 , n33216 , n36167 );
    or g41180 ( n29975 , n17739 , n11216 );
    nor g41181 ( n6599 , n34354 , n28687 );
    or g41182 ( n23579 , n7839 , n22757 );
    or g41183 ( n22208 , n4333 , n35497 );
    or g41184 ( n7951 , n4099 , n34353 );
    not g41185 ( n4340 , n8232 );
    or g41186 ( n11027 , n34114 , n1972 );
    nor g41187 ( n11935 , n16396 , n8804 );
    or g41188 ( n14138 , n42067 , n25885 );
    nor g41189 ( n3016 , n32085 , n32838 );
    not g41190 ( n38058 , n41301 );
    xnor g41191 ( n22708 , n15347 , n18680 );
    or g41192 ( n41953 , n12706 , n41361 );
    and g41193 ( n37659 , n30755 , n42728 );
    and g41194 ( n1608 , n6470 , n19208 );
    and g41195 ( n30658 , n3772 , n934 );
    nor g41196 ( n11756 , n6762 , n23860 );
    not g41197 ( n6211 , n42116 );
    not g41198 ( n4707 , n39393 );
    or g41199 ( n2531 , n37952 , n5133 );
    not g41200 ( n39773 , n6367 );
    or g41201 ( n26694 , n9313 , n23152 );
    nor g41202 ( n23538 , n37163 , n14081 );
    or g41203 ( n16749 , n6249 , n39796 );
    and g41204 ( n38381 , n11980 , n12843 );
    or g41205 ( n16849 , n23447 , n32983 );
    or g41206 ( n35203 , n38463 , n28453 );
    nor g41207 ( n309 , n9336 , n9238 );
    or g41208 ( n33699 , n15113 , n41344 );
    and g41209 ( n41567 , n32190 , n15122 );
    or g41210 ( n31248 , n4018 , n18425 );
    not g41211 ( n7460 , n20593 );
    or g41212 ( n18413 , n28970 , n2597 );
    or g41213 ( n36493 , n40368 , n21884 );
    xnor g41214 ( n12328 , n28541 , n13854 );
    nor g41215 ( n8214 , n38879 , n21976 );
    nor g41216 ( n3467 , n18275 , n42751 );
    xnor g41217 ( n15321 , n34731 , n34315 );
    not g41218 ( n15443 , n15841 );
    or g41219 ( n38782 , n37964 , n15404 );
    and g41220 ( n12168 , n41805 , n38837 );
    nor g41221 ( n26865 , n34090 , n8094 );
    or g41222 ( n23526 , n1788 , n939 );
    not g41223 ( n19787 , n30126 );
    xnor g41224 ( n1474 , n12524 , n5142 );
    or g41225 ( n37281 , n9477 , n26305 );
    nor g41226 ( n4372 , n9371 , n1603 );
    nor g41227 ( n31978 , n9573 , n41619 );
    xnor g41228 ( n16539 , n21957 , n8355 );
    not g41229 ( n4385 , n7035 );
    not g41230 ( n21415 , n10943 );
    or g41231 ( n12912 , n14622 , n1293 );
    or g41232 ( n5304 , n28138 , n42416 );
    xnor g41233 ( n8862 , n23510 , n15484 );
    or g41234 ( n15369 , n20913 , n14776 );
    and g41235 ( n7798 , n31637 , n28630 );
    or g41236 ( n17852 , n15064 , n2208 );
    or g41237 ( n12360 , n25781 , n13594 );
    or g41238 ( n26715 , n26116 , n33502 );
    and g41239 ( n36030 , n26644 , n32054 );
    and g41240 ( n5289 , n14862 , n37757 );
    or g41241 ( n8248 , n1735 , n25200 );
    not g41242 ( n34664 , n31159 );
    not g41243 ( n36712 , n38898 );
    nor g41244 ( n31600 , n14279 , n12172 );
    or g41245 ( n31930 , n30263 , n38574 );
    or g41246 ( n32074 , n31309 , n30821 );
    nor g41247 ( n42754 , n784 , n27922 );
    nor g41248 ( n27454 , n27281 , n19180 );
    or g41249 ( n19162 , n24662 , n12210 );
    xnor g41250 ( n25539 , n105 , n40339 );
    nor g41251 ( n41474 , n39544 , n29752 );
    or g41252 ( n22937 , n23006 , n6655 );
    xnor g41253 ( n20876 , n6625 , n13980 );
    and g41254 ( n34215 , n26184 , n30261 );
    nor g41255 ( n13757 , n33292 , n3336 );
    or g41256 ( n40458 , n3634 , n35689 );
    nor g41257 ( n18686 , n41728 , n23280 );
    and g41258 ( n25389 , n29226 , n19874 );
    nor g41259 ( n30134 , n32069 , n35269 );
    not g41260 ( n30889 , n35737 );
    or g41261 ( n16446 , n37980 , n21872 );
    or g41262 ( n42900 , n36408 , n22670 );
    not g41263 ( n29147 , n14712 );
    and g41264 ( n4892 , n8348 , n26396 );
    or g41265 ( n40355 , n13273 , n5789 );
    or g41266 ( n24968 , n26272 , n18975 );
    nor g41267 ( n17279 , n22184 , n23624 );
    nor g41268 ( n23189 , n14471 , n15107 );
    not g41269 ( n6578 , n32887 );
    not g41270 ( n14837 , n11589 );
    or g41271 ( n23650 , n12285 , n10017 );
    not g41272 ( n20083 , n17163 );
    and g41273 ( n5779 , n34918 , n11379 );
    or g41274 ( n21967 , n3941 , n20446 );
    and g41275 ( n8914 , n30734 , n32176 );
    and g41276 ( n13664 , n40087 , n979 );
    nor g41277 ( n30882 , n32015 , n28552 );
    xnor g41278 ( n41818 , n27184 , n1168 );
    nor g41279 ( n37108 , n6565 , n40317 );
    or g41280 ( n10827 , n14956 , n12059 );
    or g41281 ( n14349 , n9523 , n5243 );
    and g41282 ( n11071 , n3986 , n5996 );
    or g41283 ( n18040 , n8576 , n1244 );
    not g41284 ( n37378 , n10435 );
    not g41285 ( n7433 , n7597 );
    nor g41286 ( n30670 , n39645 , n29521 );
    nor g41287 ( n33380 , n3447 , n38816 );
    and g41288 ( n26281 , n10566 , n15878 );
    and g41289 ( n37290 , n19481 , n22058 );
    and g41290 ( n6066 , n21320 , n14303 );
    or g41291 ( n17933 , n21071 , n17855 );
    and g41292 ( n41484 , n24914 , n6430 );
    and g41293 ( n2114 , n36784 , n42268 );
    and g41294 ( n37994 , n21999 , n4286 );
    nor g41295 ( n26860 , n20128 , n42687 );
    or g41296 ( n27040 , n39137 , n23320 );
    or g41297 ( n3458 , n10396 , n8311 );
    or g41298 ( n32005 , n33655 , n35848 );
    nor g41299 ( n17110 , n19424 , n34332 );
    or g41300 ( n36964 , n35483 , n17638 );
    xnor g41301 ( n28621 , n42725 , n34669 );
    nor g41302 ( n41011 , n22151 , n25016 );
    not g41303 ( n6660 , n37088 );
    and g41304 ( n8803 , n8800 , n985 );
    nor g41305 ( n28386 , n4920 , n16386 );
    or g41306 ( n16954 , n39283 , n29261 );
    and g41307 ( n21855 , n31429 , n35877 );
    or g41308 ( n34351 , n33134 , n88 );
    or g41309 ( n28585 , n39593 , n14063 );
    not g41310 ( n6756 , n25333 );
    xnor g41311 ( n32658 , n32154 , n6838 );
    xnor g41312 ( n4027 , n4511 , n8516 );
    or g41313 ( n37769 , n3781 , n2442 );
    and g41314 ( n36571 , n19146 , n38854 );
    or g41315 ( n35624 , n15681 , n11006 );
    and g41316 ( n13894 , n37975 , n41310 );
    or g41317 ( n28422 , n31677 , n17466 );
    xnor g41318 ( n5169 , n29740 , n3642 );
    or g41319 ( n14574 , n37712 , n6328 );
    xnor g41320 ( n12557 , n17476 , n35400 );
    or g41321 ( n16358 , n28080 , n4181 );
    nor g41322 ( n28246 , n31724 , n28425 );
    and g41323 ( n30062 , n24659 , n3428 );
    or g41324 ( n603 , n30263 , n11660 );
    not g41325 ( n21536 , n35535 );
    not g41326 ( n31007 , n16210 );
    or g41327 ( n2424 , n16101 , n39363 );
    not g41328 ( n7296 , n12041 );
    and g41329 ( n26908 , n26350 , n22194 );
    and g41330 ( n14643 , n17650 , n19395 );
    not g41331 ( n6087 , n23188 );
    not g41332 ( n14487 , n36723 );
    and g41333 ( n10856 , n40967 , n11769 );
    or g41334 ( n33759 , n32003 , n10655 );
    xnor g41335 ( n38984 , n37437 , n620 );
    or g41336 ( n3808 , n41539 , n14944 );
    not g41337 ( n439 , n13979 );
    and g41338 ( n6051 , n8494 , n34181 );
    or g41339 ( n23754 , n6507 , n18432 );
    and g41340 ( n13758 , n18386 , n31554 );
    not g41341 ( n15140 , n31945 );
    nor g41342 ( n10233 , n1301 , n28438 );
    xnor g41343 ( n27500 , n11692 , n14254 );
    not g41344 ( n27111 , n33438 );
    not g41345 ( n32346 , n7686 );
    xnor g41346 ( n21414 , n4491 , n33955 );
    or g41347 ( n28814 , n12061 , n19866 );
    xnor g41348 ( n28686 , n35074 , n14860 );
    not g41349 ( n41321 , n1842 );
    and g41350 ( n23933 , n30449 , n20774 );
    not g41351 ( n21709 , n3899 );
    or g41352 ( n23824 , n16521 , n17411 );
    or g41353 ( n30016 , n21072 , n26078 );
    nor g41354 ( n17073 , n20390 , n4483 );
    and g41355 ( n19015 , n19759 , n19877 );
    xnor g41356 ( n728 , n29740 , n33912 );
    nor g41357 ( n39334 , n1081 , n214 );
    or g41358 ( n12664 , n29373 , n21028 );
    not g41359 ( n865 , n21065 );
    and g41360 ( n10170 , n42178 , n29687 );
    not g41361 ( n36590 , n9028 );
    or g41362 ( n16241 , n12181 , n38022 );
    nor g41363 ( n39026 , n37302 , n7520 );
    not g41364 ( n38121 , n30713 );
    or g41365 ( n40466 , n39366 , n13721 );
    not g41366 ( n36413 , n27206 );
    or g41367 ( n38141 , n18236 , n22464 );
    xnor g41368 ( n5410 , n6625 , n30799 );
    not g41369 ( n15261 , n33220 );
    or g41370 ( n39468 , n40295 , n17505 );
    or g41371 ( n30734 , n12856 , n28234 );
    nor g41372 ( n26554 , n9616 , n35019 );
    or g41373 ( n22643 , n38387 , n17312 );
    or g41374 ( n7147 , n40913 , n6307 );
    and g41375 ( n37399 , n14839 , n38204 );
    and g41376 ( n15255 , n35017 , n25186 );
    or g41377 ( n21416 , n38463 , n35187 );
    nor g41378 ( n14794 , n39266 , n23757 );
    and g41379 ( n31675 , n9058 , n5825 );
    xnor g41380 ( n16030 , n23070 , n11150 );
    or g41381 ( n38934 , n17800 , n17392 );
    nor g41382 ( n33094 , n38511 , n41004 );
    nor g41383 ( n11028 , n5611 , n28905 );
    xnor g41384 ( n271 , n39848 , n2199 );
    and g41385 ( n4462 , n18218 , n2243 );
    not g41386 ( n11147 , n24687 );
    or g41387 ( n29269 , n42487 , n21772 );
    not g41388 ( n36001 , n13099 );
    nor g41389 ( n8972 , n7356 , n26317 );
    xnor g41390 ( n22153 , n17708 , n20892 );
    or g41391 ( n33147 , n28111 , n5778 );
    or g41392 ( n12989 , n23256 , n19753 );
    not g41393 ( n35391 , n5478 );
    xnor g41394 ( n39298 , n6625 , n40043 );
    or g41395 ( n23514 , n25286 , n1324 );
    or g41396 ( n357 , n12565 , n20249 );
    nor g41397 ( n15980 , n21595 , n39687 );
    or g41398 ( n33568 , n42115 , n33964 );
    nor g41399 ( n17758 , n1075 , n14873 );
    not g41400 ( n19768 , n20441 );
    not g41401 ( n12224 , n25025 );
    xnor g41402 ( n38908 , n29854 , n33223 );
    xnor g41403 ( n9776 , n5891 , n18080 );
    or g41404 ( n1920 , n39059 , n13944 );
    not g41405 ( n3223 , n19928 );
    or g41406 ( n33429 , n8697 , n41429 );
    xnor g41407 ( n17155 , n28319 , n26809 );
    and g41408 ( n3526 , n13621 , n5417 );
    and g41409 ( n4612 , n24410 , n36624 );
    and g41410 ( n40306 , n13271 , n18692 );
    xnor g41411 ( n17937 , n29057 , n11312 );
    and g41412 ( n34470 , n12147 , n27149 );
    not g41413 ( n42842 , n33702 );
    xnor g41414 ( n12070 , n36567 , n34375 );
    and g41415 ( n15718 , n32622 , n3059 );
    or g41416 ( n9088 , n20760 , n5422 );
    nor g41417 ( n14923 , n23868 , n32587 );
    and g41418 ( n38448 , n37033 , n10891 );
    xnor g41419 ( n9555 , n14801 , n4674 );
    and g41420 ( n6898 , n7697 , n3778 );
    or g41421 ( n1832 , n8656 , n29730 );
    or g41422 ( n12928 , n18914 , n24024 );
    or g41423 ( n1627 , n9471 , n808 );
    or g41424 ( n35278 , n904 , n13599 );
    nor g41425 ( n15560 , n2083 , n32634 );
    or g41426 ( n29062 , n35386 , n6311 );
    xnor g41427 ( n27395 , n37896 , n23335 );
    and g41428 ( n37435 , n20885 , n19646 );
    xnor g41429 ( n62 , n35378 , n8494 );
    and g41430 ( n26097 , n35727 , n10863 );
    not g41431 ( n2146 , n21370 );
    or g41432 ( n34045 , n9484 , n21584 );
    nor g41433 ( n30834 , n38777 , n4360 );
    xnor g41434 ( n30042 , n1316 , n14345 );
    or g41435 ( n484 , n27287 , n24327 );
    and g41436 ( n22018 , n34488 , n12141 );
    or g41437 ( n11278 , n11076 , n40323 );
    or g41438 ( n5866 , n11651 , n17084 );
    and g41439 ( n38143 , n15263 , n39561 );
    or g41440 ( n10458 , n22199 , n28500 );
    and g41441 ( n20901 , n23014 , n21194 );
    or g41442 ( n14890 , n26933 , n32214 );
    nor g41443 ( n27775 , n5540 , n17564 );
    xnor g41444 ( n21407 , n35553 , n30610 );
    xnor g41445 ( n14017 , n5041 , n37913 );
    or g41446 ( n31708 , n39372 , n1044 );
    or g41447 ( n19686 , n24656 , n13564 );
    not g41448 ( n16194 , n8267 );
    and g41449 ( n38305 , n25984 , n5902 );
    or g41450 ( n33801 , n36420 , n8253 );
    nor g41451 ( n31038 , n28749 , n17862 );
    or g41452 ( n40441 , n10329 , n35080 );
    and g41453 ( n20179 , n8608 , n37734 );
    or g41454 ( n33844 , n36754 , n32388 );
    or g41455 ( n18674 , n3764 , n26630 );
    not g41456 ( n751 , n28003 );
    xnor g41457 ( n21891 , n9133 , n12791 );
    not g41458 ( n36070 , n16101 );
    or g41459 ( n39482 , n5868 , n4582 );
    or g41460 ( n489 , n9354 , n8679 );
    xnor g41461 ( n15941 , n29970 , n10598 );
    not g41462 ( n4904 , n25544 );
    or g41463 ( n33726 , n14321 , n21992 );
    or g41464 ( n4918 , n40981 , n40169 );
    and g41465 ( n39585 , n27373 , n27822 );
    and g41466 ( n3622 , n8046 , n40589 );
    or g41467 ( n18216 , n19468 , n40065 );
    nor g41468 ( n6272 , n29461 , n41896 );
    not g41469 ( n22278 , n597 );
    or g41470 ( n1148 , n6654 , n5183 );
    or g41471 ( n15279 , n39850 , n12635 );
    nor g41472 ( n321 , n15325 , n9986 );
    or g41473 ( n28493 , n8788 , n36022 );
    and g41474 ( n12546 , n689 , n7224 );
    and g41475 ( n28361 , n3076 , n31833 );
    not g41476 ( n35982 , n22644 );
    or g41477 ( n27602 , n34436 , n9311 );
    or g41478 ( n33317 , n6423 , n27203 );
    and g41479 ( n18652 , n1460 , n10689 );
    not g41480 ( n8035 , n14589 );
    or g41481 ( n4466 , n22057 , n34985 );
    or g41482 ( n9374 , n26545 , n25011 );
    or g41483 ( n40131 , n25966 , n31497 );
    and g41484 ( n30186 , n10243 , n916 );
    or g41485 ( n14113 , n20413 , n34609 );
    or g41486 ( n2248 , n38590 , n12637 );
    nor g41487 ( n5806 , n11115 , n32677 );
    and g41488 ( n33607 , n7661 , n31463 );
    or g41489 ( n5425 , n24620 , n30891 );
    xnor g41490 ( n14523 , n14596 , n6027 );
    and g41491 ( n16660 , n7489 , n3194 );
    xnor g41492 ( n4590 , n7915 , n5410 );
    or g41493 ( n36674 , n17566 , n28432 );
    not g41494 ( n8439 , n2919 );
    or g41495 ( n2581 , n40094 , n6359 );
    and g41496 ( n9207 , n26557 , n42094 );
    or g41497 ( n6489 , n12425 , n24030 );
    xnor g41498 ( n36829 , n21415 , n36518 );
    not g41499 ( n20310 , n39200 );
    and g41500 ( n41997 , n1566 , n11826 );
    nor g41501 ( n38235 , n36117 , n21080 );
    nor g41502 ( n28032 , n6754 , n29231 );
    or g41503 ( n34122 , n21426 , n37414 );
    and g41504 ( n34552 , n17290 , n19013 );
    and g41505 ( n31869 , n12111 , n33888 );
    or g41506 ( n8315 , n40145 , n21552 );
    and g41507 ( n39379 , n17245 , n13901 );
    xnor g41508 ( n10771 , n23742 , n14471 );
    xnor g41509 ( n42612 , n23867 , n39634 );
    nor g41510 ( n15931 , n36484 , n34165 );
    or g41511 ( n26528 , n42010 , n18596 );
    and g41512 ( n37454 , n9143 , n5880 );
    and g41513 ( n6468 , n12467 , n33741 );
    and g41514 ( n1144 , n14857 , n32354 );
    or g41515 ( n26436 , n42243 , n37031 );
    and g41516 ( n17780 , n29435 , n3341 );
    and g41517 ( n394 , n39858 , n22536 );
    or g41518 ( n1860 , n14707 , n38658 );
    or g41519 ( n14824 , n32762 , n970 );
    or g41520 ( n7272 , n7637 , n33226 );
    nor g41521 ( n3892 , n41343 , n14160 );
    and g41522 ( n12515 , n19255 , n34900 );
    or g41523 ( n30636 , n42659 , n4039 );
    or g41524 ( n9476 , n32683 , n36439 );
    xnor g41525 ( n2685 , n20386 , n36402 );
    or g41526 ( n32444 , n36804 , n20895 );
    or g41527 ( n19309 , n122 , n558 );
    or g41528 ( n2138 , n9625 , n18578 );
    and g41529 ( n39988 , n16444 , n42495 );
    and g41530 ( n12345 , n6776 , n39421 );
    and g41531 ( n586 , n31261 , n21195 );
    or g41532 ( n40849 , n9725 , n31497 );
    xnor g41533 ( n20415 , n14613 , n2126 );
    or g41534 ( n13070 , n20301 , n42603 );
    or g41535 ( n40986 , n40862 , n17857 );
    or g41536 ( n8785 , n35422 , n34949 );
    or g41537 ( n24109 , n33981 , n9443 );
    nor g41538 ( n29178 , n27721 , n34128 );
    nor g41539 ( n34769 , n6860 , n10127 );
    nor g41540 ( n15382 , n38712 , n40088 );
    or g41541 ( n22116 , n28263 , n9396 );
    nor g41542 ( n42625 , n21199 , n27933 );
    xnor g41543 ( n29481 , n21534 , n15759 );
    not g41544 ( n14443 , n9065 );
    or g41545 ( n30425 , n12542 , n14917 );
    nor g41546 ( n39275 , n14707 , n27374 );
    buf g41547 ( n19009 , n8407 );
    or g41548 ( n24767 , n12059 , n4757 );
    or g41549 ( n8764 , n6742 , n33453 );
    or g41550 ( n24881 , n644 , n30921 );
    nor g41551 ( n12255 , n18866 , n12121 );
    or g41552 ( n32164 , n4713 , n20517 );
    and g41553 ( n24931 , n21606 , n38651 );
    or g41554 ( n41488 , n40540 , n38858 );
    not g41555 ( n19202 , n12337 );
    or g41556 ( n551 , n2120 , n30626 );
    and g41557 ( n41528 , n33606 , n38470 );
    or g41558 ( n39872 , n30801 , n39856 );
    or g41559 ( n7562 , n38879 , n34643 );
    and g41560 ( n37427 , n34207 , n40564 );
    xnor g41561 ( n8529 , n2501 , n40342 );
    not g41562 ( n41462 , n8008 );
    not g41563 ( n25631 , n40753 );
    xnor g41564 ( n23797 , n12946 , n41070 );
    and g41565 ( n33680 , n28587 , n26658 );
    not g41566 ( n15474 , n36838 );
    not g41567 ( n36788 , n5244 );
    xnor g41568 ( n21484 , n4334 , n17164 );
    not g41569 ( n25105 , n5337 );
    or g41570 ( n33207 , n7070 , n10766 );
    or g41571 ( n5547 , n18826 , n4808 );
    and g41572 ( n25787 , n5601 , n34585 );
    xnor g41573 ( n6203 , n38173 , n29607 );
    and g41574 ( n10272 , n41020 , n27634 );
    and g41575 ( n17052 , n36914 , n10179 );
    or g41576 ( n20143 , n5102 , n29916 );
    or g41577 ( n12587 , n28021 , n24277 );
    nor g41578 ( n8584 , n28917 , n11152 );
    xnor g41579 ( n26261 , n11436 , n42144 );
    or g41580 ( n16424 , n16994 , n12448 );
    not g41581 ( n26570 , n15676 );
    xnor g41582 ( n2843 , n13735 , n2538 );
    or g41583 ( n29940 , n17045 , n37787 );
    xnor g41584 ( n7685 , n27644 , n14473 );
    and g41585 ( n30155 , n4417 , n22438 );
    nor g41586 ( n19600 , n38879 , n38063 );
    or g41587 ( n32382 , n38879 , n28729 );
    or g41588 ( n30342 , n9362 , n24490 );
    and g41589 ( n17169 , n24258 , n12032 );
    or g41590 ( n30858 , n18475 , n19888 );
    or g41591 ( n24082 , n19762 , n12417 );
    or g41592 ( n26292 , n27033 , n37077 );
    or g41593 ( n24474 , n10592 , n40306 );
    not g41594 ( n31201 , n38367 );
    not g41595 ( n28596 , n19226 );
    or g41596 ( n1654 , n38247 , n27430 );
    not g41597 ( n10452 , n42738 );
    not g41598 ( n7555 , n28817 );
    or g41599 ( n40998 , n9877 , n27683 );
    not g41600 ( n27840 , n22306 );
    or g41601 ( n19105 , n30861 , n11650 );
    not g41602 ( n40702 , n3178 );
    or g41603 ( n30515 , n29913 , n13024 );
    and g41604 ( n34036 , n37261 , n34878 );
    not g41605 ( n30648 , n30303 );
    xnor g41606 ( n30697 , n35938 , n28646 );
    not g41607 ( n29751 , n24847 );
    and g41608 ( n19290 , n42910 , n10877 );
    and g41609 ( n10032 , n5253 , n42043 );
    not g41610 ( n11133 , n8663 );
    and g41611 ( n22714 , n22435 , n15104 );
    and g41612 ( n3362 , n36449 , n24478 );
    or g41613 ( n7787 , n25573 , n25776 );
    and g41614 ( n18827 , n19504 , n20806 );
    nor g41615 ( n40429 , n9150 , n35869 );
    or g41616 ( n1755 , n40735 , n42743 );
    or g41617 ( n7886 , n4949 , n15952 );
    xnor g41618 ( n36274 , n41013 , n28078 );
    xnor g41619 ( n618 , n32351 , n31030 );
    or g41620 ( n33905 , n12175 , n8061 );
    nor g41621 ( n39865 , n13023 , n32162 );
    nor g41622 ( n38082 , n38261 , n12811 );
    not g41623 ( n37041 , n22097 );
    not g41624 ( n5808 , n19667 );
    not g41625 ( n41247 , n30469 );
    xnor g41626 ( n6030 , n11436 , n15500 );
    or g41627 ( n5969 , n23491 , n26731 );
    or g41628 ( n10745 , n42227 , n41943 );
    not g41629 ( n42320 , n32431 );
    nor g41630 ( n11035 , n15537 , n7212 );
    nor g41631 ( n24883 , n17764 , n40075 );
    or g41632 ( n6763 , n29649 , n32918 );
    xnor g41633 ( n19369 , n42898 , n22199 );
    or g41634 ( n26306 , n39489 , n4964 );
    or g41635 ( n36593 , n35969 , n13938 );
    or g41636 ( n9119 , n40210 , n12046 );
    not g41637 ( n41519 , n5600 );
    xnor g41638 ( n35616 , n32955 , n10120 );
    and g41639 ( n1993 , n24983 , n14111 );
    or g41640 ( n26504 , n5048 , n24463 );
    not g41641 ( n1496 , n33496 );
    and g41642 ( n10918 , n33935 , n42451 );
    xnor g41643 ( n12891 , n37742 , n33981 );
    xnor g41644 ( n3158 , n15111 , n2671 );
    xnor g41645 ( n33809 , n10782 , n29506 );
    nor g41646 ( n24375 , n33981 , n17078 );
    and g41647 ( n31211 , n1955 , n38682 );
    and g41648 ( n8994 , n18993 , n11532 );
    or g41649 ( n41173 , n37579 , n27535 );
    and g41650 ( n11069 , n16747 , n23336 );
    or g41651 ( n24368 , n25152 , n9983 );
    and g41652 ( n30472 , n4103 , n30052 );
    or g41653 ( n26467 , n28597 , n35831 );
    nor g41654 ( n26516 , n12521 , n23364 );
    or g41655 ( n29705 , n7737 , n41158 );
    and g41656 ( n39755 , n33207 , n5344 );
    or g41657 ( n27272 , n14481 , n32189 );
    xnor g41658 ( n40993 , n2753 , n27567 );
    or g41659 ( n18765 , n21879 , n10888 );
    nor g41660 ( n12852 , n21184 , n12234 );
    or g41661 ( n28542 , n1066 , n42361 );
    nor g41662 ( n18621 , n26419 , n38364 );
    not g41663 ( n14338 , n10779 );
    and g41664 ( n12104 , n1364 , n1304 );
    xnor g41665 ( n35345 , n41013 , n21157 );
    or g41666 ( n21345 , n34095 , n31321 );
    xnor g41667 ( n2385 , n3549 , n13381 );
    or g41668 ( n35034 , n20102 , n16466 );
    and g41669 ( n40629 , n32337 , n17242 );
    or g41670 ( n1697 , n18011 , n29249 );
    or g41671 ( n10270 , n15662 , n41651 );
    nor g41672 ( n3924 , n15118 , n6886 );
    or g41673 ( n41051 , n41760 , n12252 );
    not g41674 ( n40808 , n24802 );
    xnor g41675 ( n8238 , n24745 , n23771 );
    xnor g41676 ( n19211 , n105 , n37752 );
    or g41677 ( n694 , n39351 , n25158 );
    or g41678 ( n24806 , n10530 , n4372 );
    nor g41679 ( n335 , n33266 , n8802 );
    or g41680 ( n40793 , n27783 , n40994 );
    nor g41681 ( n27147 , n14226 , n2316 );
    and g41682 ( n331 , n2329 , n26080 );
    not g41683 ( n41705 , n17918 );
    and g41684 ( n2104 , n34394 , n10171 );
    or g41685 ( n19746 , n35386 , n22677 );
    nor g41686 ( n24138 , n5964 , n7682 );
    or g41687 ( n32774 , n12383 , n17418 );
    not g41688 ( n17086 , n7106 );
    or g41689 ( n20696 , n27454 , n40679 );
    and g41690 ( n23744 , n38526 , n10015 );
    or g41691 ( n3792 , n19599 , n16798 );
    not g41692 ( n38630 , n2089 );
    or g41693 ( n5727 , n7177 , n9785 );
    xnor g41694 ( n35424 , n18736 , n2542 );
    or g41695 ( n19047 , n21721 , n15830 );
    and g41696 ( n5498 , n26199 , n10977 );
    or g41697 ( n15069 , n28586 , n19553 );
    nor g41698 ( n11780 , n25173 , n2198 );
    not g41699 ( n20086 , n32001 );
    nor g41700 ( n18474 , n18928 , n610 );
    and g41701 ( n2768 , n18754 , n26742 );
    or g41702 ( n8905 , n7293 , n9958 );
    xnor g41703 ( n20733 , n28126 , n23281 );
    or g41704 ( n29572 , n42105 , n25907 );
    not g41705 ( n14932 , n40173 );
    or g41706 ( n40280 , n22013 , n24330 );
    and g41707 ( n825 , n993 , n10840 );
    xnor g41708 ( n3551 , n19596 , n18496 );
    not g41709 ( n39766 , n24622 );
    nor g41710 ( n14673 , n6145 , n3230 );
    or g41711 ( n23481 , n16897 , n20359 );
    and g41712 ( n21232 , n11491 , n33444 );
    or g41713 ( n19779 , n36363 , n37633 );
    nor g41714 ( n6775 , n13899 , n15986 );
    not g41715 ( n15437 , n8949 );
    or g41716 ( n17931 , n24644 , n27503 );
    and g41717 ( n25543 , n21167 , n12563 );
    or g41718 ( n35119 , n23148 , n39509 );
    nor g41719 ( n20152 , n38156 , n2869 );
    not g41720 ( n32786 , n9161 );
    and g41721 ( n21761 , n19801 , n15213 );
    and g41722 ( n4446 , n42035 , n37773 );
    nor g41723 ( n9903 , n14471 , n5518 );
    or g41724 ( n1434 , n40151 , n15092 );
    nor g41725 ( n5322 , n12779 , n16704 );
    and g41726 ( n7869 , n18790 , n1595 );
    and g41727 ( n11146 , n15343 , n38889 );
    not g41728 ( n2136 , n34137 );
    nor g41729 ( n21483 , n8633 , n188 );
    and g41730 ( n7649 , n9856 , n7581 );
    or g41731 ( n5439 , n13282 , n23042 );
    and g41732 ( n24766 , n8208 , n8140 );
    and g41733 ( n3692 , n39916 , n21609 );
    xnor g41734 ( n12359 , n37860 , n21883 );
    or g41735 ( n27487 , n5318 , n25626 );
    nor g41736 ( n33463 , n24373 , n9599 );
    or g41737 ( n3048 , n21430 , n37590 );
    and g41738 ( n40443 , n34240 , n41491 );
    and g41739 ( n8823 , n39429 , n19544 );
    and g41740 ( n5343 , n12268 , n21523 );
    xnor g41741 ( n41741 , n22263 , n20373 );
    nor g41742 ( n29208 , n9892 , n39747 );
    or g41743 ( n13953 , n17169 , n1337 );
    or g41744 ( n15865 , n22174 , n10872 );
    not g41745 ( n41662 , n21710 );
    or g41746 ( n35853 , n26280 , n37788 );
    and g41747 ( n10125 , n25723 , n18783 );
    and g41748 ( n18557 , n26997 , n28567 );
    xnor g41749 ( n957 , n17299 , n9265 );
    and g41750 ( n7935 , n30108 , n38246 );
    and g41751 ( n3550 , n34894 , n23766 );
    and g41752 ( n32691 , n2453 , n10366 );
    or g41753 ( n14003 , n24203 , n22881 );
    not g41754 ( n15379 , n7834 );
    or g41755 ( n21630 , n11259 , n17383 );
    or g41756 ( n16868 , n11119 , n10198 );
    or g41757 ( n16626 , n24216 , n32332 );
    and g41758 ( n14825 , n36271 , n28356 );
    or g41759 ( n1172 , n42186 , n3303 );
    or g41760 ( n29220 , n17193 , n20242 );
    and g41761 ( n40057 , n3125 , n4041 );
    xnor g41762 ( n39566 , n34731 , n12545 );
    or g41763 ( n24393 , n15096 , n34788 );
    xnor g41764 ( n1828 , n32701 , n23589 );
    xnor g41765 ( n39680 , n6278 , n25963 );
    nor g41766 ( n28014 , n25588 , n3439 );
    and g41767 ( n13867 , n8177 , n14479 );
    not g41768 ( n14117 , n14718 );
    nor g41769 ( n5534 , n3836 , n2625 );
    and g41770 ( n7485 , n8193 , n18418 );
    and g41771 ( n27998 , n22786 , n13962 );
    not g41772 ( n30513 , n35394 );
    nor g41773 ( n11721 , n17120 , n6874 );
    and g41774 ( n38184 , n16099 , n29326 );
    xnor g41775 ( n17628 , n42064 , n22945 );
    or g41776 ( n33290 , n21359 , n541 );
    nor g41777 ( n25628 , n25386 , n20536 );
    xnor g41778 ( n19617 , n34875 , n28539 );
    and g41779 ( n31641 , n39017 , n32220 );
    or g41780 ( n28449 , n25319 , n19803 );
    or g41781 ( n6064 , n34793 , n879 );
    not g41782 ( n726 , n10587 );
    or g41783 ( n42632 , n19811 , n25038 );
    or g41784 ( n13676 , n26226 , n16635 );
    or g41785 ( n25843 , n2394 , n500 );
    nor g41786 ( n5545 , n545 , n8019 );
    or g41787 ( n29465 , n550 , n15238 );
    or g41788 ( n35648 , n35483 , n10790 );
    or g41789 ( n35954 , n27943 , n25250 );
    or g41790 ( n39524 , n33464 , n25881 );
    and g41791 ( n24177 , n29606 , n36156 );
    not g41792 ( n784 , n8494 );
    nor g41793 ( n28812 , n29411 , n29688 );
    nor g41794 ( n38715 , n39266 , n22701 );
    not g41795 ( n34434 , n1029 );
    or g41796 ( n38802 , n437 , n4810 );
    nor g41797 ( n35086 , n1965 , n17043 );
    and g41798 ( n7085 , n30272 , n415 );
    or g41799 ( n6795 , n21352 , n10450 );
    and g41800 ( n40876 , n33276 , n6523 );
    not g41801 ( n7156 , n39452 );
    and g41802 ( n27315 , n34045 , n19705 );
    or g41803 ( n21726 , n2055 , n22463 );
    and g41804 ( n5518 , n20743 , n39044 );
    xnor g41805 ( n25406 , n37685 , n19672 );
    or g41806 ( n2369 , n3922 , n19003 );
    nor g41807 ( n42903 , n21634 , n8823 );
    and g41808 ( n30340 , n4520 , n30213 );
    nor g41809 ( n34318 , n33880 , n36232 );
    or g41810 ( n7657 , n14503 , n21129 );
    or g41811 ( n3559 , n19469 , n18694 );
    nor g41812 ( n18447 , n20490 , n22736 );
    or g41813 ( n36496 , n30078 , n7378 );
    or g41814 ( n24029 , n24665 , n12455 );
    or g41815 ( n27845 , n1114 , n1631 );
    or g41816 ( n39546 , n14611 , n12170 );
    or g41817 ( n38026 , n24131 , n923 );
    nor g41818 ( n24925 , n13338 , n19318 );
    xnor g41819 ( n19771 , n23755 , n25542 );
    nor g41820 ( n12385 , n11057 , n2807 );
    or g41821 ( n18029 , n9452 , n734 );
    xnor g41822 ( n13699 , n7723 , n19828 );
    not g41823 ( n19436 , n6116 );
    and g41824 ( n967 , n4777 , n35169 );
    not g41825 ( n40753 , n3140 );
    xnor g41826 ( n39885 , n40964 , n11280 );
    not g41827 ( n32041 , n37456 );
    xnor g41828 ( n11599 , n21946 , n5045 );
    xnor g41829 ( n6198 , n784 , n42510 );
    not g41830 ( n34024 , n13165 );
    nor g41831 ( n9369 , n10297 , n11439 );
    or g41832 ( n13250 , n4648 , n3410 );
    nor g41833 ( n28919 , n41761 , n41238 );
    and g41834 ( n36550 , n31930 , n17521 );
    xnor g41835 ( n33163 , n31099 , n22762 );
    and g41836 ( n20076 , n33920 , n9247 );
    and g41837 ( n18805 , n2164 , n41885 );
    or g41838 ( n13312 , n20341 , n29388 );
    not g41839 ( n3093 , n28910 );
    or g41840 ( n3877 , n28900 , n13470 );
    or g41841 ( n18832 , n38321 , n29158 );
    xnor g41842 ( n11628 , n42698 , n20595 );
    xnor g41843 ( n9046 , n32794 , n38117 );
    or g41844 ( n28182 , n21754 , n20170 );
    xnor g41845 ( n12919 , n35553 , n10733 );
    or g41846 ( n14620 , n9807 , n36605 );
    or g41847 ( n29722 , n2436 , n21025 );
    and g41848 ( n3302 , n28187 , n23288 );
    or g41849 ( n29794 , n11452 , n31430 );
    xnor g41850 ( n32766 , n9597 , n35533 );
    or g41851 ( n20361 , n34463 , n28401 );
    not g41852 ( n24689 , n17726 );
    or g41853 ( n24511 , n35355 , n6429 );
    and g41854 ( n40447 , n6799 , n30534 );
    and g41855 ( n10755 , n17207 , n32871 );
    xnor g41856 ( n41572 , n38222 , n5964 );
    or g41857 ( n42767 , n14941 , n34849 );
    or g41858 ( n16905 , n32574 , n10063 );
    not g41859 ( n27505 , n35208 );
    and g41860 ( n27701 , n38724 , n12951 );
    xnor g41861 ( n34479 , n784 , n36091 );
    or g41862 ( n40357 , n24371 , n28875 );
    or g41863 ( n18633 , n34292 , n12787 );
    or g41864 ( n19191 , n24196 , n31580 );
    nor g41865 ( n38688 , n40128 , n42867 );
    not g41866 ( n17691 , n6724 );
    not g41867 ( n13 , n23550 );
    and g41868 ( n39831 , n41818 , n37442 );
    and g41869 ( n14222 , n26449 , n24444 );
    xnor g41870 ( n30346 , n21982 , n25293 );
    xnor g41871 ( n7817 , n29740 , n37972 );
    and g41872 ( n33337 , n30745 , n35686 );
    and g41873 ( n21235 , n2191 , n3979 );
    or g41874 ( n16463 , n31553 , n6850 );
    or g41875 ( n13934 , n32150 , n31551 );
    or g41876 ( n8273 , n5120 , n12083 );
    and g41877 ( n36929 , n21458 , n27152 );
    or g41878 ( n16640 , n38718 , n41632 );
    or g41879 ( n130 , n22102 , n26417 );
    xnor g41880 ( n3369 , n39104 , n1369 );
    xnor g41881 ( n22891 , n8425 , n15442 );
    and g41882 ( n38303 , n30904 , n9219 );
    or g41883 ( n417 , n13676 , n4008 );
    or g41884 ( n41842 , n11174 , n13081 );
    xnor g41885 ( n34397 , n35509 , n10846 );
    not g41886 ( n24273 , n12332 );
    or g41887 ( n914 , n31174 , n16703 );
    and g41888 ( n24695 , n36523 , n30372 );
    and g41889 ( n38409 , n8654 , n34259 );
    or g41890 ( n37636 , n9617 , n28997 );
    and g41891 ( n16260 , n31385 , n2941 );
    xnor g41892 ( n42236 , n29858 , n12883 );
    and g41893 ( n11361 , n40085 , n36692 );
    or g41894 ( n5918 , n35386 , n42820 );
    and g41895 ( n15127 , n40113 , n19568 );
    or g41896 ( n30942 , n32283 , n38447 );
    and g41897 ( n8346 , n6287 , n23339 );
    or g41898 ( n38624 , n25033 , n7921 );
    or g41899 ( n33221 , n14417 , n11755 );
    and g41900 ( n22688 , n10283 , n41770 );
    and g41901 ( n19733 , n1706 , n2289 );
    and g41902 ( n17736 , n18193 , n31909 );
    not g41903 ( n11464 , n7390 );
    not g41904 ( n11900 , n25288 );
    or g41905 ( n25514 , n35963 , n22900 );
    or g41906 ( n26717 , n23088 , n42918 );
    and g41907 ( n36917 , n28459 , n17237 );
    or g41908 ( n40289 , n38762 , n28596 );
    nor g41909 ( n39819 , n12054 , n314 );
    not g41910 ( n8837 , n5940 );
    not g41911 ( n6584 , n35935 );
    and g41912 ( n17005 , n27348 , n24942 );
    nor g41913 ( n18464 , n12885 , n21069 );
    or g41914 ( n22393 , n22631 , n26380 );
    or g41915 ( n20501 , n32313 , n14281 );
    nor g41916 ( n12423 , n29859 , n18898 );
    nor g41917 ( n5962 , n2091 , n31767 );
    xnor g41918 ( n31097 , n6547 , n39651 );
    nor g41919 ( n11500 , n14125 , n22911 );
    nor g41920 ( n12022 , n19519 , n39173 );
    xnor g41921 ( n41608 , n27762 , n5085 );
    or g41922 ( n32198 , n36517 , n9748 );
    not g41923 ( n23353 , n12578 );
    or g41924 ( n1941 , n1642 , n14304 );
    and g41925 ( n5377 , n3412 , n7225 );
    or g41926 ( n1209 , n12927 , n41021 );
    or g41927 ( n28098 , n14622 , n34000 );
    and g41928 ( n40445 , n12054 , n3869 );
    or g41929 ( n33181 , n38029 , n40894 );
    or g41930 ( n8995 , n23552 , n25132 );
    or g41931 ( n4450 , n33981 , n456 );
    not g41932 ( n11658 , n30088 );
    or g41933 ( n12932 , n31268 , n15538 );
    or g41934 ( n41364 , n31153 , n36548 );
    and g41935 ( n7854 , n26169 , n17128 );
    nor g41936 ( n28041 , n1379 , n11783 );
    or g41937 ( n16317 , n5854 , n14809 );
    and g41938 ( n23480 , n39438 , n41404 );
    and g41939 ( n16832 , n19462 , n2521 );
    or g41940 ( n39866 , n32800 , n14829 );
    or g41941 ( n41926 , n35019 , n20978 );
    and g41942 ( n29100 , n20212 , n20213 );
    or g41943 ( n2465 , n7590 , n440 );
    or g41944 ( n18281 , n3764 , n38420 );
    not g41945 ( n33080 , n34800 );
    not g41946 ( n23263 , n6679 );
    or g41947 ( n22277 , n7150 , n23182 );
    nor g41948 ( n1620 , n14467 , n7279 );
    or g41949 ( n33449 , n33464 , n21873 );
    and g41950 ( n33718 , n12349 , n17278 );
    not g41951 ( n31361 , n23365 );
    or g41952 ( n36784 , n38829 , n13824 );
    nor g41953 ( n16807 , n12888 , n21271 );
    not g41954 ( n27142 , n28530 );
    and g41955 ( n39730 , n695 , n6601 );
    nor g41956 ( n18748 , n17744 , n18273 );
    or g41957 ( n37190 , n14602 , n26031 );
    not g41958 ( n20393 , n16075 );
    or g41959 ( n34097 , n6156 , n19790 );
    and g41960 ( n28715 , n19876 , n19716 );
    or g41961 ( n9166 , n6423 , n6105 );
    or g41962 ( n38478 , n16308 , n3900 );
    nor g41963 ( n37086 , n42427 , n37188 );
    not g41964 ( n39556 , n40861 );
    nor g41965 ( n29291 , n3835 , n29770 );
    or g41966 ( n10591 , n38119 , n23805 );
    not g41967 ( n28999 , n25949 );
    or g41968 ( n40362 , n41420 , n15342 );
    and g41969 ( n14621 , n7769 , n29760 );
    nor g41970 ( n23122 , n12828 , n21666 );
    and g41971 ( n13814 , n26236 , n34935 );
    or g41972 ( n24518 , n981 , n5136 );
    or g41973 ( n39084 , n23292 , n21550 );
    and g41974 ( n24048 , n35035 , n29392 );
    or g41975 ( n30133 , n13529 , n40492 );
    and g41976 ( n12982 , n37327 , n28193 );
    and g41977 ( n27480 , n30654 , n23178 );
    or g41978 ( n19216 , n4848 , n40420 );
    or g41979 ( n17645 , n15282 , n41129 );
    or g41980 ( n13293 , n7139 , n18267 );
    nor g41981 ( n39619 , n4334 , n22856 );
    and g41982 ( n10517 , n13444 , n31036 );
    or g41983 ( n12132 , n40183 , n36827 );
    or g41984 ( n4572 , n1688 , n8363 );
    or g41985 ( n5592 , n36815 , n31315 );
    and g41986 ( n36169 , n40849 , n7437 );
    and g41987 ( n37648 , n3040 , n25408 );
    or g41988 ( n39077 , n20631 , n23286 );
    and g41989 ( n28275 , n6084 , n22029 );
    or g41990 ( n22555 , n36835 , n13968 );
    not g41991 ( n25246 , n24868 );
    or g41992 ( n469 , n2786 , n3501 );
    nor g41993 ( n21102 , n7047 , n32333 );
    or g41994 ( n40267 , n37123 , n19331 );
    and g41995 ( n17505 , n24401 , n319 );
    or g41996 ( n37515 , n47 , n2587 );
    or g41997 ( n24851 , n17927 , n4446 );
    nor g41998 ( n1491 , n26017 , n35634 );
    and g41999 ( n1733 , n37888 , n39637 );
    or g42000 ( n8947 , n4952 , n29150 );
    or g42001 ( n23597 , n35870 , n25423 );
    nor g42002 ( n13197 , n59 , n38763 );
    not g42003 ( n8081 , n25345 );
    and g42004 ( n34010 , n15506 , n5293 );
    or g42005 ( n41872 , n15282 , n16553 );
    and g42006 ( n3750 , n10729 , n40361 );
    or g42007 ( n25654 , n33866 , n18507 );
    not g42008 ( n23847 , n27506 );
    or g42009 ( n12460 , n32274 , n18102 );
    and g42010 ( n13783 , n25982 , n39522 );
    and g42011 ( n1202 , n36778 , n19940 );
    or g42012 ( n35393 , n11417 , n26769 );
    and g42013 ( n24905 , n7602 , n565 );
    and g42014 ( n10296 , n1241 , n5752 );
    and g42015 ( n5538 , n8851 , n40334 );
    or g42016 ( n38349 , n40911 , n19159 );
    xnor g42017 ( n33863 , n39852 , n42462 );
    and g42018 ( n36300 , n39862 , n2247 );
    or g42019 ( n11475 , n18179 , n12456 );
    xnor g42020 ( n8577 , n33851 , n15754 );
    xnor g42021 ( n1295 , n39183 , n41634 );
    not g42022 ( n4302 , n6161 );
    or g42023 ( n28307 , n41441 , n31716 );
    not g42024 ( n1395 , n32272 );
    or g42025 ( n17171 , n35866 , n5218 );
    not g42026 ( n745 , n13810 );
    or g42027 ( n11963 , n15529 , n25416 );
    not g42028 ( n19607 , n29089 );
    not g42029 ( n10748 , n26749 );
    or g42030 ( n16592 , n18339 , n6247 );
    and g42031 ( n16839 , n23605 , n42148 );
    or g42032 ( n30792 , n42669 , n18654 );
    or g42033 ( n14131 , n42386 , n1908 );
    or g42034 ( n31158 , n10955 , n41389 );
    xnor g42035 ( n9841 , n9142 , n17304 );
    or g42036 ( n13727 , n10460 , n37395 );
    not g42037 ( n31220 , n40629 );
    xnor g42038 ( n40025 , n6914 , n15248 );
    and g42039 ( n26932 , n12974 , n19712 );
    not g42040 ( n28911 , n19515 );
    or g42041 ( n40091 , n11849 , n29919 );
    not g42042 ( n16862 , n17179 );
    or g42043 ( n38641 , n3781 , n4387 );
    or g42044 ( n36686 , n14707 , n37705 );
    or g42045 ( n18289 , n6365 , n13942 );
    and g42046 ( n2793 , n24681 , n26083 );
    or g42047 ( n1736 , n14259 , n14668 );
    and g42048 ( n31571 , n20891 , n12935 );
    or g42049 ( n13998 , n991 , n19811 );
    or g42050 ( n28709 , n12484 , n21928 );
    nor g42051 ( n24637 , n13981 , n1785 );
    nor g42052 ( n23397 , n38621 , n18078 );
    nor g42053 ( n2995 , n35553 , n37019 );
    and g42054 ( n35042 , n6249 , n39796 );
    xnor g42055 ( n3774 , n784 , n26947 );
    or g42056 ( n2652 , n33775 , n37360 );
    not g42057 ( n18727 , n24266 );
    not g42058 ( n7532 , n33108 );
    not g42059 ( n17830 , n6468 );
    and g42060 ( n29165 , n5165 , n39706 );
    and g42061 ( n3337 , n32023 , n1480 );
    or g42062 ( n41214 , n6462 , n11167 );
    xnor g42063 ( n41016 , n23947 , n42540 );
    xnor g42064 ( n16869 , n32253 , n23406 );
    xnor g42065 ( n34585 , n29740 , n21080 );
    or g42066 ( n10887 , n33262 , n5075 );
    xnor g42067 ( n51 , n25631 , n31869 );
    and g42068 ( n2495 , n10700 , n41505 );
    or g42069 ( n19025 , n25902 , n25553 );
    nor g42070 ( n20277 , n40902 , n5440 );
    nor g42071 ( n15329 , n38879 , n3097 );
    not g42072 ( n2680 , n11733 );
    nor g42073 ( n23383 , n14014 , n22205 );
    or g42074 ( n29357 , n8494 , n30318 );
    not g42075 ( n30018 , n37721 );
    and g42076 ( n21900 , n4684 , n38757 );
    or g42077 ( n798 , n30496 , n28522 );
    and g42078 ( n1265 , n31899 , n1682 );
    or g42079 ( n17675 , n23445 , n18269 );
    not g42080 ( n3619 , n2661 );
    and g42081 ( n8219 , n35597 , n29861 );
    or g42082 ( n10164 , n36772 , n21068 );
    and g42083 ( n35524 , n22927 , n6 );
    nor g42084 ( n3522 , n19700 , n12388 );
    and g42085 ( n34082 , n40692 , n34 );
    nor g42086 ( n40209 , n37685 , n15776 );
    or g42087 ( n9765 , n10095 , n30301 );
    and g42088 ( n12690 , n42398 , n7310 );
    xnor g42089 ( n28581 , n19592 , n37360 );
    and g42090 ( n26417 , n12543 , n1858 );
    or g42091 ( n15574 , n40261 , n3561 );
    or g42092 ( n4497 , n7616 , n12573 );
    or g42093 ( n23852 , n2209 , n23126 );
    nor g42094 ( n1447 , n14707 , n10081 );
    or g42095 ( n13834 , n22122 , n27768 );
    or g42096 ( n6920 , n23615 , n35456 );
    nor g42097 ( n41442 , n42413 , n10133 );
    not g42098 ( n26213 , n14299 );
    and g42099 ( n27367 , n23961 , n41454 );
    or g42100 ( n517 , n30358 , n40675 );
    nor g42101 ( n11520 , n40369 , n11828 );
    or g42102 ( n24669 , n5665 , n15848 );
    or g42103 ( n30466 , n39057 , n3873 );
    and g42104 ( n28359 , n33949 , n29257 );
    xnor g42105 ( n20908 , n27874 , n25179 );
    or g42106 ( n941 , n2224 , n8863 );
    or g42107 ( n22500 , n22121 , n23722 );
    or g42108 ( n2993 , n21046 , n39919 );
    and g42109 ( n12705 , n33959 , n15518 );
    or g42110 ( n11138 , n26900 , n11789 );
    or g42111 ( n23731 , n40730 , n5476 );
    and g42112 ( n18788 , n34196 , n4513 );
    and g42113 ( n13670 , n29181 , n34388 );
    and g42114 ( n12618 , n4175 , n42612 );
    and g42115 ( n1567 , n22049 , n7620 );
    not g42116 ( n40281 , n27905 );
    not g42117 ( n38805 , n34422 );
    and g42118 ( n23771 , n26913 , n19537 );
    or g42119 ( n36174 , n39292 , n20422 );
    or g42120 ( n6361 , n35471 , n23957 );
    not g42121 ( n8157 , n27545 );
    or g42122 ( n10019 , n5048 , n26096 );
    not g42123 ( n21372 , n22310 );
    not g42124 ( n9180 , n32277 );
    xnor g42125 ( n41541 , n24411 , n4365 );
    or g42126 ( n18977 , n41699 , n2835 );
    and g42127 ( n12540 , n36340 , n13142 );
    or g42128 ( n28272 , n22098 , n20694 );
    and g42129 ( n8074 , n26402 , n23293 );
    or g42130 ( n24694 , n3837 , n799 );
    or g42131 ( n6638 , n25136 , n20519 );
    not g42132 ( n30378 , n14514 );
    not g42133 ( n36762 , n7109 );
    or g42134 ( n22429 , n17888 , n6199 );
    or g42135 ( n7589 , n9475 , n6359 );
    or g42136 ( n15413 , n7838 , n19138 );
    nor g42137 ( n38075 , n34292 , n17005 );
    or g42138 ( n31903 , n19803 , n36172 );
    or g42139 ( n18410 , n33515 , n1100 );
    nor g42140 ( n39806 , n17906 , n40741 );
    or g42141 ( n41120 , n4339 , n17173 );
    or g42142 ( n24604 , n41667 , n33531 );
    and g42143 ( n1729 , n4525 , n31269 );
    and g42144 ( n35149 , n26926 , n29093 );
    or g42145 ( n2176 , n13810 , n904 );
    not g42146 ( n31261 , n877 );
    or g42147 ( n18318 , n34918 , n23145 );
    nor g42148 ( n30678 , n13604 , n31806 );
    and g42149 ( n42734 , n31084 , n7497 );
    or g42150 ( n18437 , n12220 , n21180 );
    or g42151 ( n22300 , n37682 , n8988 );
    or g42152 ( n11741 , n16899 , n38162 );
    or g42153 ( n42527 , n13282 , n10727 );
    or g42154 ( n19100 , n1789 , n17703 );
    not g42155 ( n20338 , n25325 );
    and g42156 ( n18315 , n7491 , n28738 );
    or g42157 ( n37174 , n26820 , n10646 );
    not g42158 ( n41947 , n1743 );
    or g42159 ( n6909 , n7603 , n30652 );
    not g42160 ( n9174 , n41277 );
    xnor g42161 ( n12151 , n16693 , n11683 );
    nor g42162 ( n30941 , n35262 , n9439 );
    or g42163 ( n39005 , n4655 , n17173 );
    nor g42164 ( n29026 , n31286 , n33432 );
    and g42165 ( n5199 , n24688 , n42038 );
    not g42166 ( n40679 , n7920 );
    and g42167 ( n39636 , n29243 , n863 );
    nor g42168 ( n32819 , n22710 , n24208 );
    nor g42169 ( n20880 , n16618 , n27623 );
    not g42170 ( n34114 , n5522 );
    or g42171 ( n29374 , n1549 , n34163 );
    not g42172 ( n7598 , n35224 );
    xnor g42173 ( n13564 , n30673 , n13829 );
    and g42174 ( n319 , n11382 , n7930 );
    and g42175 ( n9953 , n28761 , n20481 );
    and g42176 ( n11230 , n35146 , n38432 );
    not g42177 ( n17313 , n29094 );
    not g42178 ( n31265 , n22863 );
    xnor g42179 ( n28254 , n25283 , n5245 );
    or g42180 ( n16026 , n27781 , n17401 );
    or g42181 ( n32993 , n4951 , n10572 );
    or g42182 ( n27685 , n11346 , n9038 );
    not g42183 ( n28821 , n19120 );
    xnor g42184 ( n13274 , n17159 , n5989 );
    nor g42185 ( n37669 , n32721 , n14323 );
    nor g42186 ( n37430 , n6890 , n11488 );
    and g42187 ( n11925 , n5494 , n2019 );
    not g42188 ( n23097 , n3236 );
    nor g42189 ( n28015 , n15153 , n40394 );
    not g42190 ( n41569 , n16263 );
    not g42191 ( n3094 , n40486 );
    not g42192 ( n31958 , n42016 );
    not g42193 ( n5701 , n8081 );
    or g42194 ( n6940 , n3006 , n9183 );
    or g42195 ( n26418 , n38066 , n3055 );
    xnor g42196 ( n24388 , n26210 , n27105 );
    xnor g42197 ( n10635 , n25706 , n1507 );
    or g42198 ( n42005 , n15116 , n34864 );
    or g42199 ( n2826 , n17466 , n19104 );
    xnor g42200 ( n36576 , n33919 , n1937 );
    and g42201 ( n39507 , n26705 , n37946 );
    or g42202 ( n9333 , n29493 , n4237 );
    not g42203 ( n2232 , n21561 );
    or g42204 ( n19343 , n21296 , n12983 );
    and g42205 ( n2829 , n15148 , n15180 );
    and g42206 ( n29451 , n41343 , n14160 );
    and g42207 ( n4478 , n19075 , n15034 );
    not g42208 ( n23867 , n1743 );
    nor g42209 ( n33842 , n10676 , n10242 );
    or g42210 ( n16392 , n29214 , n21433 );
    and g42211 ( n36277 , n39450 , n24960 );
    and g42212 ( n39097 , n6697 , n193 );
    nor g42213 ( n36265 , n23678 , n20857 );
    or g42214 ( n34510 , n35735 , n14622 );
    and g42215 ( n19340 , n20713 , n27222 );
    or g42216 ( n10102 , n30376 , n34051 );
    or g42217 ( n14207 , n28163 , n35027 );
    or g42218 ( n36033 , n2401 , n10530 );
    xnor g42219 ( n34986 , n7922 , n14983 );
    nor g42220 ( n29073 , n35374 , n7251 );
    and g42221 ( n28067 , n18392 , n32396 );
    or g42222 ( n8298 , n29382 , n7490 );
    xnor g42223 ( n11348 , n32470 , n2732 );
    xnor g42224 ( n33821 , n21973 , n31027 );
    not g42225 ( n13248 , n33305 );
    or g42226 ( n16871 , n16598 , n20939 );
    nor g42227 ( n27637 , n27137 , n32274 );
    xnor g42228 ( n33365 , n39182 , n42894 );
    and g42229 ( n6839 , n20028 , n26527 );
    or g42230 ( n20923 , n32100 , n6169 );
    xnor g42231 ( n18942 , n105 , n19989 );
    or g42232 ( n12572 , n16910 , n14860 );
    xnor g42233 ( n39438 , n16418 , n34638 );
    xnor g42234 ( n7724 , n15611 , n23410 );
    and g42235 ( n20818 , n38583 , n36894 );
    or g42236 ( n40803 , n40563 , n19848 );
    or g42237 ( n27559 , n18782 , n12040 );
    or g42238 ( n22311 , n16903 , n12612 );
    xnor g42239 ( n10921 , n18530 , n36612 );
    or g42240 ( n13395 , n34191 , n3603 );
    and g42241 ( n36535 , n34872 , n30240 );
    and g42242 ( n17606 , n16035 , n10767 );
    and g42243 ( n33235 , n39333 , n21543 );
    or g42244 ( n42167 , n20742 , n40325 );
    or g42245 ( n18568 , n20817 , n4365 );
    not g42246 ( n42460 , n40925 );
    nor g42247 ( n20710 , n17510 , n24940 );
    nor g42248 ( n16916 , n1507 , n9798 );
    or g42249 ( n38308 , n18252 , n19423 );
    or g42250 ( n26474 , n42896 , n39001 );
    xnor g42251 ( n15331 , n7489 , n14985 );
    not g42252 ( n38721 , n15354 );
    nor g42253 ( n6720 , n37639 , n39939 );
    or g42254 ( n4744 , n32980 , n1065 );
    xnor g42255 ( n2243 , n12161 , n26667 );
    xnor g42256 ( n16059 , n37899 , n38374 );
    and g42257 ( n13553 , n9326 , n7438 );
    and g42258 ( n32263 , n32900 , n34304 );
    xnor g42259 ( n2363 , n28909 , n29971 );
    xnor g42260 ( n8813 , n21784 , n11166 );
    not g42261 ( n30044 , n12394 );
    and g42262 ( n15015 , n35205 , n28600 );
    and g42263 ( n30732 , n26880 , n11700 );
    and g42264 ( n32247 , n682 , n41017 );
    nor g42265 ( n40316 , n23330 , n21205 );
    or g42266 ( n28659 , n16541 , n17468 );
    or g42267 ( n2251 , n16109 , n1217 );
    and g42268 ( n17172 , n26253 , n23038 );
    or g42269 ( n18929 , n34686 , n19580 );
    or g42270 ( n35206 , n20726 , n13209 );
    and g42271 ( n41443 , n30248 , n12091 );
    or g42272 ( n7523 , n36522 , n38556 );
    or g42273 ( n11224 , n32082 , n23194 );
    and g42274 ( n40505 , n2070 , n8799 );
    or g42275 ( n8141 , n84 , n16899 );
    or g42276 ( n30699 , n33216 , n14928 );
    or g42277 ( n31383 , n33461 , n19327 );
    or g42278 ( n1864 , n253 , n18328 );
    not g42279 ( n3934 , n42338 );
    nor g42280 ( n3288 , n8904 , n3541 );
    nor g42281 ( n11470 , n29056 , n39814 );
    and g42282 ( n20567 , n12304 , n33429 );
    or g42283 ( n5600 , n35487 , n5271 );
    nor g42284 ( n36050 , n15070 , n38904 );
    and g42285 ( n32644 , n33231 , n42592 );
    or g42286 ( n41454 , n22823 , n11590 );
    or g42287 ( n32284 , n14508 , n7853 );
    nor g42288 ( n38969 , n1490 , n11477 );
    not g42289 ( n4896 , n30684 );
    or g42290 ( n38050 , n24639 , n40702 );
    xnor g42291 ( n14807 , n33053 , n30114 );
    or g42292 ( n21434 , n23694 , n27771 );
    or g42293 ( n4317 , n10898 , n38181 );
    not g42294 ( n36813 , n3098 );
    and g42295 ( n6669 , n24085 , n25952 );
    not g42296 ( n30132 , n5548 );
    and g42297 ( n1425 , n7608 , n480 );
    nor g42298 ( n22130 , n9711 , n21787 );
    nor g42299 ( n40052 , n17120 , n38743 );
    not g42300 ( n9607 , n38991 );
    nor g42301 ( n17075 , n29821 , n37561 );
    xnor g42302 ( n3286 , n38886 , n7227 );
    or g42303 ( n1237 , n27536 , n34083 );
    not g42304 ( n15678 , n10396 );
    not g42305 ( n25461 , n18884 );
    xnor g42306 ( n23781 , n24651 , n3825 );
    or g42307 ( n35186 , n25398 , n4221 );
    and g42308 ( n5584 , n2571 , n20304 );
    or g42309 ( n9433 , n31428 , n22379 );
    and g42310 ( n42675 , n29272 , n15321 );
    xnor g42311 ( n25861 , n35727 , n22499 );
    or g42312 ( n5618 , n14612 , n25924 );
    and g42313 ( n19659 , n40211 , n18036 );
    not g42314 ( n6957 , n25607 );
    nor g42315 ( n41857 , n24896 , n17163 );
    not g42316 ( n40180 , n30880 );
    or g42317 ( n17793 , n24384 , n16593 );
    or g42318 ( n22583 , n5546 , n1307 );
    or g42319 ( n31933 , n26028 , n37050 );
    and g42320 ( n40966 , n21733 , n6757 );
    and g42321 ( n10333 , n27959 , n36180 );
    and g42322 ( n15610 , n24184 , n15656 );
    or g42323 ( n20490 , n41333 , n7083 );
    xnor g42324 ( n42825 , n21301 , n30547 );
    or g42325 ( n28943 , n26915 , n8309 );
    or g42326 ( n24871 , n39954 , n3514 );
    xnor g42327 ( n23539 , n20487 , n28337 );
    nor g42328 ( n28713 , n2274 , n11587 );
    and g42329 ( n18421 , n22380 , n20006 );
    xnor g42330 ( n31830 , n17762 , n21061 );
    nor g42331 ( n15087 , n8787 , n7094 );
    or g42332 ( n42432 , n9544 , n27192 );
    or g42333 ( n2067 , n22456 , n24918 );
    or g42334 ( n438 , n14964 , n33173 );
    nor g42335 ( n41571 , n9318 , n26594 );
    not g42336 ( n37733 , n30287 );
    and g42337 ( n1488 , n3928 , n27343 );
    or g42338 ( n32541 , n14289 , n42066 );
    not g42339 ( n20296 , n30929 );
    and g42340 ( n21046 , n19638 , n7155 );
    not g42341 ( n35759 , n26749 );
    xnor g42342 ( n5234 , n19282 , n12733 );
    xnor g42343 ( n40474 , n16320 , n39749 );
    or g42344 ( n14092 , n414 , n17827 );
    xnor g42345 ( n36034 , n9460 , n23254 );
    not g42346 ( n31707 , n14055 );
    and g42347 ( n14014 , n16804 , n27833 );
    and g42348 ( n27936 , n1796 , n38491 );
    or g42349 ( n39387 , n28143 , n9867 );
    nor g42350 ( n34515 , n17697 , n1282 );
    or g42351 ( n4622 , n18798 , n38510 );
    nor g42352 ( n28714 , n41278 , n13630 );
    or g42353 ( n5132 , n19009 , n17540 );
    or g42354 ( n9500 , n42454 , n39690 );
    or g42355 ( n40630 , n4425 , n32735 );
    not g42356 ( n39508 , n38666 );
    not g42357 ( n29047 , n3280 );
    and g42358 ( n19627 , n10390 , n27291 );
    not g42359 ( n5279 , n15567 );
    and g42360 ( n37385 , n32158 , n21823 );
    not g42361 ( n8414 , n13383 );
    not g42362 ( n26862 , n38474 );
    or g42363 ( n4827 , n2745 , n27526 );
    or g42364 ( n24985 , n10720 , n931 );
    and g42365 ( n8941 , n18839 , n31230 );
    nor g42366 ( n19424 , n19353 , n12662 );
    nor g42367 ( n22703 , n42455 , n20055 );
    nor g42368 ( n18082 , n2923 , n35229 );
    nor g42369 ( n11467 , n35874 , n40116 );
    nor g42370 ( n26787 , n785 , n41717 );
    or g42371 ( n10556 , n24268 , n3811 );
    and g42372 ( n21359 , n27994 , n24213 );
    not g42373 ( n34522 , n35389 );
    or g42374 ( n9527 , n38905 , n39804 );
    or g42375 ( n4882 , n8539 , n15183 );
    nor g42376 ( n3591 , n18550 , n18706 );
    xnor g42377 ( n9499 , n10834 , n38977 );
    and g42378 ( n1417 , n16574 , n38635 );
    nor g42379 ( n32409 , n4983 , n32505 );
    xnor g42380 ( n6307 , n6625 , n23219 );
    xnor g42381 ( n26761 , n25198 , n12531 );
    nor g42382 ( n10766 , n38879 , n39621 );
    and g42383 ( n31818 , n40913 , n6307 );
    xnor g42384 ( n13863 , n784 , n27878 );
    nor g42385 ( n24245 , n31368 , n41346 );
    or g42386 ( n15204 , n9456 , n26982 );
    not g42387 ( n25067 , n40496 );
    or g42388 ( n18064 , n33141 , n8659 );
    not g42389 ( n18127 , n32241 );
    and g42390 ( n39282 , n34798 , n17584 );
    nor g42391 ( n33553 , n39456 , n39550 );
    not g42392 ( n28749 , n31138 );
    xnor g42393 ( n26555 , n31554 , n18386 );
    nor g42394 ( n38103 , n22168 , n33821 );
    xnor g42395 ( n3695 , n6625 , n25121 );
    and g42396 ( n32370 , n28534 , n26590 );
    not g42397 ( n30549 , n37306 );
    and g42398 ( n8899 , n32297 , n3860 );
    or g42399 ( n21903 , n23085 , n28171 );
    and g42400 ( n32745 , n34815 , n36878 );
    or g42401 ( n29530 , n10747 , n5867 );
    or g42402 ( n40864 , n32087 , n20406 );
    not g42403 ( n27789 , n18285 );
    and g42404 ( n1399 , n23360 , n13879 );
    nor g42405 ( n13917 , n26377 , n16067 );
    or g42406 ( n31943 , n28883 , n39563 );
    nor g42407 ( n7675 , n1927 , n38214 );
    or g42408 ( n11662 , n26915 , n34906 );
    or g42409 ( n2177 , n22202 , n40447 );
    or g42410 ( n25374 , n12075 , n29930 );
    nor g42411 ( n22239 , n36996 , n41887 );
    or g42412 ( n23074 , n24621 , n41962 );
    nor g42413 ( n29116 , n17393 , n11632 );
    or g42414 ( n39401 , n11890 , n15282 );
    nor g42415 ( n29447 , n1507 , n15255 );
    nor g42416 ( n11006 , n25337 , n26890 );
    or g42417 ( n41000 , n14503 , n22422 );
    or g42418 ( n23569 , n2628 , n39526 );
    xnor g42419 ( n34364 , n105 , n39694 );
    or g42420 ( n18237 , n16565 , n10898 );
    or g42421 ( n12094 , n31186 , n40178 );
    and g42422 ( n26482 , n15383 , n30940 );
    or g42423 ( n37874 , n12385 , n39063 );
    or g42424 ( n4459 , n33433 , n42610 );
    or g42425 ( n38134 , n41998 , n23183 );
    or g42426 ( n37324 , n28087 , n22997 );
    or g42427 ( n32281 , n41332 , n24894 );
    and g42428 ( n19774 , n443 , n31082 );
    nor g42429 ( n5785 , n4334 , n4971 );
    or g42430 ( n30211 , n5850 , n28388 );
    and g42431 ( n13804 , n13443 , n26685 );
    and g42432 ( n32827 , n11886 , n42836 );
    or g42433 ( n658 , n1025 , n35829 );
    not g42434 ( n453 , n26268 );
    and g42435 ( n42307 , n32897 , n12005 );
    nor g42436 ( n37580 , n465 , n18844 );
    xnor g42437 ( n2362 , n29692 , n7161 );
    nor g42438 ( n2237 , n13 , n16511 );
    not g42439 ( n9250 , n24876 );
    xnor g42440 ( n4655 , n20858 , n12798 );
    not g42441 ( n14840 , n10279 );
    not g42442 ( n22660 , n34654 );
    xnor g42443 ( n35399 , n6625 , n12923 );
    nor g42444 ( n26470 , n58 , n17351 );
    nor g42445 ( n3237 , n22057 , n7048 );
    or g42446 ( n40002 , n36377 , n11901 );
    xnor g42447 ( n21646 , n5174 , n11269 );
    and g42448 ( n34854 , n9788 , n7627 );
    or g42449 ( n6698 , n36411 , n8498 );
    and g42450 ( n16081 , n5060 , n28001 );
    and g42451 ( n6467 , n38672 , n11519 );
    or g42452 ( n14335 , n32683 , n8408 );
    nor g42453 ( n27412 , n9951 , n25202 );
    or g42454 ( n8287 , n20897 , n28487 );
    xnor g42455 ( n37762 , n12954 , n21691 );
    and g42456 ( n32239 , n27961 , n31546 );
    or g42457 ( n6994 , n15382 , n42077 );
    and g42458 ( n3629 , n3044 , n40522 );
    or g42459 ( n5801 , n33624 , n13860 );
    or g42460 ( n30621 , n5310 , n5284 );
    xnor g42461 ( n23994 , n31099 , n20934 );
    not g42462 ( n25191 , n19720 );
    or g42463 ( n9728 , n19090 , n8214 );
    and g42464 ( n8967 , n42884 , n11555 );
    xnor g42465 ( n8098 , n7870 , n28400 );
    xnor g42466 ( n11719 , n24862 , n20981 );
    not g42467 ( n27965 , n40953 );
    not g42468 ( n42572 , n101 );
    or g42469 ( n7273 , n14898 , n17532 );
    or g42470 ( n19124 , n18182 , n17321 );
    or g42471 ( n27281 , n991 , n20949 );
    not g42472 ( n7143 , n37801 );
    or g42473 ( n9600 , n2454 , n26922 );
    nor g42474 ( n30647 , n29592 , n33769 );
    or g42475 ( n9348 , n37664 , n22249 );
    xnor g42476 ( n31505 , n35727 , n42308 );
    and g42477 ( n9470 , n23780 , n26163 );
    and g42478 ( n20660 , n8364 , n27689 );
    nor g42479 ( n19905 , n11245 , n23437 );
    and g42480 ( n23006 , n12163 , n7023 );
    or g42481 ( n23340 , n17393 , n32714 );
    or g42482 ( n74 , n18121 , n11814 );
    nor g42483 ( n29282 , n36117 , n33912 );
    and g42484 ( n24187 , n42572 , n18991 );
    or g42485 ( n19573 , n25136 , n39411 );
    not g42486 ( n18424 , n8641 );
    nor g42487 ( n28783 , n12873 , n19433 );
    or g42488 ( n28773 , n38702 , n24077 );
    or g42489 ( n5502 , n781 , n19496 );
    and g42490 ( n39501 , n27281 , n19180 );
    not g42491 ( n17768 , n31142 );
    and g42492 ( n23002 , n35470 , n2635 );
    not g42493 ( n7116 , n4426 );
    xnor g42494 ( n16822 , n14758 , n32125 );
    not g42495 ( n9150 , n31781 );
    or g42496 ( n36318 , n5849 , n21772 );
    or g42497 ( n23232 , n39358 , n23703 );
    and g42498 ( n27619 , n18266 , n22596 );
    or g42499 ( n5652 , n2935 , n3952 );
    nor g42500 ( n28984 , n11636 , n39278 );
    and g42501 ( n18593 , n14701 , n34032 );
    xnor g42502 ( n25063 , n10408 , n16243 );
    xnor g42503 ( n40941 , n34731 , n576 );
    xnor g42504 ( n30379 , n38326 , n3807 );
    nor g42505 ( n42520 , n16780 , n11510 );
    or g42506 ( n19749 , n609 , n22108 );
    or g42507 ( n30039 , n9642 , n5941 );
    and g42508 ( n36029 , n21880 , n23299 );
    not g42509 ( n23445 , n9492 );
    not g42510 ( n35656 , n26610 );
    nor g42511 ( n25615 , n29973 , n11711 );
    nor g42512 ( n16470 , n38577 , n30000 );
    not g42513 ( n13002 , n36526 );
    or g42514 ( n24025 , n35730 , n30652 );
    and g42515 ( n24322 , n17618 , n35893 );
    or g42516 ( n4629 , n41526 , n37606 );
    or g42517 ( n17209 , n25033 , n5741 );
    and g42518 ( n40140 , n7153 , n34302 );
    not g42519 ( n25780 , n36404 );
    or g42520 ( n18824 , n23991 , n15387 );
    or g42521 ( n22124 , n11126 , n7616 );
    not g42522 ( n39348 , n14222 );
    not g42523 ( n20795 , n22704 );
    nor g42524 ( n16078 , n1779 , n20933 );
    and g42525 ( n8699 , n5448 , n26259 );
    not g42526 ( n34075 , n13262 );
    xnor g42527 ( n21991 , n28225 , n14368 );
    or g42528 ( n37450 , n2696 , n28837 );
    not g42529 ( n16717 , n30463 );
    not g42530 ( n13207 , n34472 );
    and g42531 ( n9255 , n22787 , n13672 );
    xnor g42532 ( n23937 , n11633 , n13021 );
    or g42533 ( n29486 , n38570 , n23926 );
    or g42534 ( n33234 , n42405 , n40448 );
    nor g42535 ( n14177 , n17744 , n31809 );
    or g42536 ( n6822 , n16255 , n26888 );
    xnor g42537 ( n19019 , n25299 , n5529 );
    and g42538 ( n14626 , n30156 , n11927 );
    nor g42539 ( n8242 , n9945 , n5214 );
    or g42540 ( n11089 , n42457 , n14967 );
    not g42541 ( n35174 , n14799 );
    or g42542 ( n27200 , n39524 , n25077 );
    or g42543 ( n8071 , n2668 , n3568 );
    not g42544 ( n6358 , n8734 );
    or g42545 ( n7369 , n2564 , n5714 );
    nor g42546 ( n10349 , n42111 , n34782 );
    or g42547 ( n27099 , n4669 , n35736 );
    or g42548 ( n15076 , n10674 , n19354 );
    or g42549 ( n22857 , n7839 , n8963 );
    and g42550 ( n27527 , n18400 , n41747 );
    not g42551 ( n36352 , n6496 );
    or g42552 ( n5143 , n15781 , n12053 );
    and g42553 ( n15799 , n34868 , n1121 );
    and g42554 ( n31301 , n24827 , n14802 );
    not g42555 ( n22473 , n10779 );
    nor g42556 ( n42026 , n38462 , n42388 );
    or g42557 ( n23213 , n11976 , n7157 );
    and g42558 ( n17297 , n1242 , n19023 );
    or g42559 ( n4734 , n20754 , n23928 );
    xnor g42560 ( n33850 , n2005 , n33813 );
    and g42561 ( n24776 , n12406 , n33176 );
    or g42562 ( n21467 , n40210 , n24857 );
    not g42563 ( n38081 , n40499 );
    or g42564 ( n33395 , n28607 , n24114 );
    nor g42565 ( n14085 , n2149 , n21046 );
    nor g42566 ( n40970 , n10903 , n12840 );
    xnor g42567 ( n17273 , n25050 , n22481 );
    and g42568 ( n12206 , n40454 , n42037 );
    or g42569 ( n13286 , n41580 , n6178 );
    and g42570 ( n23701 , n31658 , n26501 );
    and g42571 ( n15674 , n30790 , n38856 );
    not g42572 ( n37847 , n13627 );
    nor g42573 ( n11480 , n17097 , n18148 );
    nor g42574 ( n40497 , n38494 , n12171 );
    or g42575 ( n7072 , n14407 , n30040 );
    xnor g42576 ( n11473 , n22773 , n10878 );
    and g42577 ( n11504 , n15259 , n13748 );
    or g42578 ( n1007 , n22274 , n40481 );
    and g42579 ( n11706 , n37743 , n41311 );
    or g42580 ( n35770 , n32335 , n17104 );
    xnor g42581 ( n35842 , n35727 , n20985 );
    or g42582 ( n7803 , n24215 , n41649 );
    or g42583 ( n22527 , n17654 , n17884 );
    or g42584 ( n7852 , n12049 , n42786 );
    or g42585 ( n38877 , n38919 , n6290 );
    or g42586 ( n6451 , n5115 , n11026 );
    xnor g42587 ( n33342 , n37922 , n41216 );
    or g42588 ( n3810 , n24609 , n3916 );
    or g42589 ( n11242 , n39699 , n32370 );
    and g42590 ( n1043 , n8748 , n23128 );
    or g42591 ( n9434 , n7410 , n41353 );
    and g42592 ( n27912 , n36469 , n19319 );
    and g42593 ( n1696 , n9789 , n12470 );
    xnor g42594 ( n17099 , n26579 , n3506 );
    nor g42595 ( n25711 , n2199 , n23426 );
    not g42596 ( n33068 , n28665 );
    and g42597 ( n18412 , n3998 , n835 );
    nor g42598 ( n3618 , n16780 , n16081 );
    or g42599 ( n23105 , n20234 , n26927 );
    not g42600 ( n40773 , n20111 );
    and g42601 ( n12558 , n35390 , n34839 );
    or g42602 ( n4211 , n8611 , n13232 );
    xnor g42603 ( n8466 , n21648 , n10712 );
    not g42604 ( n94 , n15396 );
    not g42605 ( n31783 , n20220 );
    or g42606 ( n23084 , n17031 , n14944 );
    or g42607 ( n23362 , n27712 , n18808 );
    nor g42608 ( n7329 , n26294 , n21353 );
    not g42609 ( n40010 , n30706 );
    nor g42610 ( n41527 , n6908 , n4010 );
    or g42611 ( n39834 , n41009 , n40239 );
    or g42612 ( n32227 , n19828 , n32068 );
    and g42613 ( n2762 , n17053 , n32604 );
    or g42614 ( n19947 , n20935 , n26895 );
    xnor g42615 ( n1803 , n24979 , n14471 );
    and g42616 ( n29406 , n2806 , n35953 );
    not g42617 ( n38163 , n21387 );
    nor g42618 ( n25089 , n6687 , n23403 );
    nor g42619 ( n389 , n15567 , n29084 );
    nor g42620 ( n30255 , n10509 , n15598 );
    or g42621 ( n22232 , n10035 , n7839 );
    and g42622 ( n28471 , n38599 , n8295 );
    or g42623 ( n3666 , n39828 , n35270 );
    and g42624 ( n10222 , n700 , n21575 );
    nor g42625 ( n25144 , n18866 , n5365 );
    and g42626 ( n12915 , n15235 , n33992 );
    or g42627 ( n28199 , n16109 , n13172 );
    not g42628 ( n7281 , n19392 );
    and g42629 ( n22681 , n10409 , n11720 );
    or g42630 ( n14445 , n9145 , n24893 );
    and g42631 ( n35755 , n11657 , n10715 );
    nor g42632 ( n30228 , n38879 , n34477 );
    and g42633 ( n27303 , n34919 , n18661 );
    or g42634 ( n19286 , n29947 , n4623 );
    or g42635 ( n18516 , n18916 , n26228 );
    or g42636 ( n11037 , n9795 , n17035 );
    xnor g42637 ( n28237 , n35867 , n24905 );
    or g42638 ( n4417 , n6009 , n10957 );
    not g42639 ( n22608 , n19369 );
    nor g42640 ( n20442 , n20974 , n9883 );
    not g42641 ( n13697 , n2060 );
    or g42642 ( n19529 , n29882 , n17104 );
    not g42643 ( n15800 , n12098 );
    or g42644 ( n12949 , n9564 , n265 );
    and g42645 ( n13374 , n5098 , n37421 );
    or g42646 ( n5006 , n24972 , n30590 );
    or g42647 ( n18864 , n29276 , n24642 );
    and g42648 ( n31442 , n24556 , n30478 );
    and g42649 ( n20594 , n6017 , n11738 );
    xnor g42650 ( n20602 , n35727 , n36838 );
    and g42651 ( n17605 , n18049 , n12597 );
    and g42652 ( n27660 , n22810 , n1897 );
    or g42653 ( n25856 , n8004 , n35805 );
    or g42654 ( n2895 , n26924 , n30263 );
    not g42655 ( n31559 , n9740 );
    or g42656 ( n9156 , n34310 , n27037 );
    and g42657 ( n34905 , n20060 , n37082 );
    and g42658 ( n16887 , n3036 , n26048 );
    not g42659 ( n24165 , n12651 );
    nor g42660 ( n880 , n24750 , n10272 );
    xnor g42661 ( n8911 , n31857 , n466 );
    nor g42662 ( n27796 , n4546 , n38727 );
    nor g42663 ( n296 , n25815 , n30494 );
    not g42664 ( n28188 , n11592 );
    xnor g42665 ( n4014 , n38188 , n1517 );
    or g42666 ( n11926 , n19610 , n39924 );
    and g42667 ( n31516 , n34208 , n1551 );
    or g42668 ( n33110 , n19602 , n6080 );
    not g42669 ( n7936 , n17058 );
    not g42670 ( n15982 , n16302 );
    xnor g42671 ( n14478 , n26680 , n24857 );
    xnor g42672 ( n918 , n10623 , n23565 );
    or g42673 ( n9320 , n27018 , n20176 );
    or g42674 ( n6974 , n9831 , n25216 );
    xnor g42675 ( n8616 , n12954 , n37648 );
    or g42676 ( n20463 , n19260 , n9122 );
    and g42677 ( n17410 , n27099 , n21656 );
    or g42678 ( n12483 , n4065 , n40505 );
    xnor g42679 ( n33226 , n40279 , n9169 );
    and g42680 ( n25833 , n9643 , n34333 );
    or g42681 ( n6743 , n29215 , n30652 );
    not g42682 ( n31362 , n32397 );
    not g42683 ( n21306 , n28411 );
    and g42684 ( n8162 , n12386 , n3152 );
    nor g42685 ( n24418 , n29751 , n6160 );
    not g42686 ( n4085 , n4491 );
    not g42687 ( n24156 , n41847 );
    and g42688 ( n10846 , n26893 , n8925 );
    not g42689 ( n16552 , n25835 );
    or g42690 ( n15645 , n24621 , n30269 );
    or g42691 ( n22717 , n39539 , n184 );
    xnor g42692 ( n19609 , n27572 , n10378 );
    nor g42693 ( n37481 , n5763 , n36267 );
    xnor g42694 ( n11407 , n40 , n3254 );
    nor g42695 ( n2078 , n18866 , n9710 );
    or g42696 ( n4555 , n34171 , n27092 );
    and g42697 ( n34534 , n15463 , n28679 );
    nor g42698 ( n28374 , n32446 , n15172 );
    or g42699 ( n13311 , n28468 , n35233 );
    not g42700 ( n13366 , n42441 );
    or g42701 ( n27795 , n6446 , n41890 );
    or g42702 ( n10607 , n28443 , n37270 );
    not g42703 ( n40070 , n15901 );
    not g42704 ( n4483 , n38197 );
    and g42705 ( n24724 , n10583 , n14082 );
    or g42706 ( n42011 , n41705 , n35859 );
    and g42707 ( n15751 , n16392 , n14059 );
    not g42708 ( n31052 , n761 );
    nor g42709 ( n23562 , n32804 , n37040 );
    and g42710 ( n3874 , n23187 , n16813 );
    not g42711 ( n33321 , n263 );
    or g42712 ( n33208 , n13298 , n34391 );
    xnor g42713 ( n26046 , n5073 , n28363 );
    nor g42714 ( n22901 , n33981 , n20650 );
    not g42715 ( n12867 , n25978 );
    or g42716 ( n15770 , n28674 , n26740 );
    or g42717 ( n21755 , n42340 , n34669 );
    xnor g42718 ( n5821 , n10806 , n12288 );
    not g42719 ( n40455 , n3178 );
    and g42720 ( n14700 , n28397 , n1118 );
    or g42721 ( n21343 , n16910 , n39521 );
    or g42722 ( n16132 , n18504 , n3801 );
    nor g42723 ( n12988 , n27599 , n42501 );
    or g42724 ( n21488 , n25131 , n42138 );
    and g42725 ( n39311 , n21027 , n13932 );
    or g42726 ( n38380 , n32472 , n14937 );
    xnor g42727 ( n4556 , n30513 , n36128 );
    nor g42728 ( n31335 , n15623 , n24616 );
    xnor g42729 ( n2964 , n38609 , n1170 );
    xnor g42730 ( n13445 , n16693 , n4797 );
    or g42731 ( n37604 , n38771 , n7616 );
    or g42732 ( n33030 , n10358 , n42535 );
    xnor g42733 ( n19107 , n5759 , n17394 );
    and g42734 ( n39426 , n9666 , n27901 );
    not g42735 ( n27082 , n35812 );
    or g42736 ( n5836 , n25907 , n6027 );
    or g42737 ( n24290 , n42163 , n26663 );
    and g42738 ( n27787 , n16112 , n37095 );
    not g42739 ( n8651 , n32563 );
    and g42740 ( n4363 , n5519 , n2294 );
    not g42741 ( n42535 , n30794 );
    xnor g42742 ( n22525 , n7342 , n5997 );
    or g42743 ( n34157 , n24407 , n13273 );
    nor g42744 ( n20935 , n22519 , n3750 );
    or g42745 ( n31672 , n4717 , n32027 );
    and g42746 ( n32599 , n30299 , n33714 );
    and g42747 ( n22442 , n29663 , n12707 );
    or g42748 ( n10429 , n32933 , n4099 );
    xnor g42749 ( n10814 , n11633 , n3503 );
    or g42750 ( n6913 , n42577 , n13339 );
    or g42751 ( n14225 , n22409 , n30167 );
    nor g42752 ( n34809 , n1507 , n3927 );
    or g42753 ( n37469 , n40946 , n5868 );
    xnor g42754 ( n19966 , n17583 , n2549 );
    or g42755 ( n20327 , n19084 , n26654 );
    or g42756 ( n35017 , n40627 , n21886 );
    or g42757 ( n20336 , n2193 , n14327 );
    nor g42758 ( n23295 , n23478 , n26887 );
    xnor g42759 ( n5257 , n22637 , n20961 );
    or g42760 ( n40721 , n23273 , n14524 );
    or g42761 ( n31862 , n19335 , n4052 );
    xnor g42762 ( n40501 , n7585 , n13154 );
    and g42763 ( n30523 , n29369 , n26110 );
    not g42764 ( n37077 , n11852 );
    and g42765 ( n30671 , n2413 , n27115 );
    and g42766 ( n3668 , n42688 , n4844 );
    nor g42767 ( n25243 , n11147 , n4866 );
    xnor g42768 ( n36145 , n42725 , n117 );
    not g42769 ( n34648 , n7604 );
    or g42770 ( n40890 , n24183 , n26077 );
    or g42771 ( n9844 , n17961 , n5578 );
    or g42772 ( n7855 , n550 , n12505 );
    nor g42773 ( n27191 , n34565 , n38038 );
    or g42774 ( n21615 , n21111 , n24421 );
    or g42775 ( n14097 , n5109 , n39018 );
    or g42776 ( n27854 , n26401 , n29121 );
    or g42777 ( n15284 , n27092 , n36733 );
    and g42778 ( n31699 , n32461 , n32706 );
    and g42779 ( n29526 , n30492 , n17326 );
    or g42780 ( n30934 , n7925 , n27234 );
    or g42781 ( n21756 , n12529 , n5379 );
    xnor g42782 ( n25354 , n40 , n27865 );
    or g42783 ( n39255 , n40028 , n6277 );
    or g42784 ( n611 , n15470 , n20874 );
    or g42785 ( n14616 , n12570 , n23123 );
    or g42786 ( n3961 , n37513 , n22651 );
    or g42787 ( n29237 , n22381 , n13885 );
    nor g42788 ( n35550 , n6477 , n24922 );
    and g42789 ( n38594 , n1080 , n41289 );
    nor g42790 ( n28623 , n20193 , n19322 );
endmodule
