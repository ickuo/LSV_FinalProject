// Benchmark "top" written by ABC on Sun Dec 21 18:07:49 2025

module top ( 
    n7, n9, n12, n19, n33, n38, n39, n60, n64, n77, n84, n92, n119, n128,
    n132, n157, n179, n186, n187, n190, n228, n236, n238, n239, n257, n261,
    n270, n288, n297, n307, n319, n321, n326, n335, n342, n371, n377, n378,
    n380, n384, n386, n387, n389, n403, n448, n457, n482, n488, n495, n504,
    n516, n520, n530, n541, n544, n560, n564, n565, n566, n579, n591, n600,
    n601, n606, n617, n627, n636, n643, n668, n676, n697, n708, n714, n715,
    n721, n754, n758, n760, n779, n801, n807, n813, n830, n841, n850, n887,
    n894, n912, n917, n918, n937, n946, n955, n961, n962, n966, n971, n984,
    n999, n1016, n1033, n1039, n1043, n1058, n1088, n1095, n1097, n1100,
    n1119, n1125, n1135, n1150, n1172, n1175, n1177, n1180, n1181, n1182,
    n1205, n1207, n1219, n1227, n1238, n1279, n1281, n1288, n1299, n1338,
    n1353, n1357, n1361, n1362, n1363, n1366, n1391, n1396, n1402, n1406,
    n1408, n1426, n1427, n1435, n1436, n1454, n1463, n1471, n1485, n1498,
    n1503, n1515, n1518, n1519, n1534, n1540, n1553, n1568, n1575, n1598,
    n1613, n1632, n1633, n1649, n1655, n1660, n1663, n1674, n1675, n1700,
    n1707, n1729, n1740, n1743, n1753, n1755, n1756, n1768, n1788, n1790,
    n18, n56, n61, n66, n67, n75, n83, n101, n107, n112, n117, n123, n129,
    n130, n158, n165, n168, n173, n193, n211, n222, n235, n245, n249, n259,
    n262, n264, n315, n320, n337, n357, n361, n370, n375, n379, n381, n413,
    n417, n454, n456, n476, n487, n542, n547, n567, n574, n596, n611, n623,
    n635, n649, n661, n673, n722, n765, n776, n786, n793, n824, n840, n845,
    n849, n860, n878, n882, n889, n944, n951, n964, n967, n974, n1027,
    n1044, n1047, n1050, n1065, n1087, n1096, n1110, n1140, n1163, n1186,
    n1224, n1233, n1269, n1270, n1297, n1314, n1322, n1346, n1355, n1370,
    n1377, n1378, n1390, n1409, n1414, n1425, n1462, n1464, n1491, n1495,
    n1510, n1511, n1543, n1584, n1587, n1631, n1654, n1657, n1676, n1682,
    n1697, n1698, n1708, n1710, n1721, n1733, n1761, n1780, n1784, n1793,
    n1794  );
  input  n7, n9, n12, n19, n33, n38, n39, n60, n64, n77, n84, n92, n119,
    n128, n132, n157, n179, n186, n187, n190, n228, n236, n238, n239, n257,
    n261, n270, n288, n297, n307, n319, n321, n326, n335, n342, n371, n377,
    n378, n380, n384, n386, n387, n389, n403, n448, n457, n482, n488, n495,
    n504, n516, n520, n530, n541, n544, n560, n564, n565, n566, n579, n591,
    n600, n601, n606, n617, n627, n636, n643, n668, n676, n697, n708, n714,
    n715, n721, n754, n758, n760, n779, n801, n807, n813, n830, n841, n850,
    n887, n894, n912, n917, n918, n937, n946, n955, n961, n962, n966, n971,
    n984, n999, n1016, n1033, n1039, n1043, n1058, n1088, n1095, n1097,
    n1100, n1119, n1125, n1135, n1150, n1172, n1175, n1177, n1180, n1181,
    n1182, n1205, n1207, n1219, n1227, n1238, n1279, n1281, n1288, n1299,
    n1338, n1353, n1357, n1361, n1362, n1363, n1366, n1391, n1396, n1402,
    n1406, n1408, n1426, n1427, n1435, n1436, n1454, n1463, n1471, n1485,
    n1498, n1503, n1515, n1518, n1519, n1534, n1540, n1553, n1568, n1575,
    n1598, n1613, n1632, n1633, n1649, n1655, n1660, n1663, n1674, n1675,
    n1700, n1707, n1729, n1740, n1743, n1753, n1755, n1756, n1768, n1788,
    n1790;
  output n18, n56, n61, n66, n67, n75, n83, n101, n107, n112, n117, n123,
    n129, n130, n158, n165, n168, n173, n193, n211, n222, n235, n245, n249,
    n259, n262, n264, n315, n320, n337, n357, n361, n370, n375, n379, n381,
    n413, n417, n454, n456, n476, n487, n542, n547, n567, n574, n596, n611,
    n623, n635, n649, n661, n673, n722, n765, n776, n786, n793, n824, n840,
    n845, n849, n860, n878, n882, n889, n944, n951, n964, n967, n974,
    n1027, n1044, n1047, n1050, n1065, n1087, n1096, n1110, n1140, n1163,
    n1186, n1224, n1233, n1269, n1270, n1297, n1314, n1322, n1346, n1355,
    n1370, n1377, n1378, n1390, n1409, n1414, n1425, n1462, n1464, n1491,
    n1495, n1510, n1511, n1543, n1584, n1587, n1631, n1654, n1657, n1676,
    n1682, n1697, n1698, n1708, n1710, n1721, n1733, n1761, n1780, n1784,
    n1793, n1794;
  wire new_n302, new_n303, new_n304, new_n305, new_n306, new_n307_1,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315_1, new_n316, new_n317, new_n318, new_n319_1, new_n320_1,
    new_n321_1, new_n322, new_n323, new_n324, new_n325, new_n326_1,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335_1, new_n336, new_n337_1, new_n338, new_n339,
    new_n340, new_n341, new_n342_1, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n356, new_n357_1, new_n358, new_n359, new_n360,
    new_n361_1, new_n362, new_n363, new_n364, new_n365, new_n366, new_n367,
    new_n368, new_n369, new_n370_1, new_n371_1, new_n372, new_n374,
    new_n375_1, new_n376, new_n377_1, new_n378_1, new_n379_1, new_n380_1,
    new_n381_1, new_n382, new_n383, new_n384_1, new_n385, new_n386_1,
    new_n387_1, new_n388, new_n389_1, new_n390, new_n391, new_n392,
    new_n393, new_n394, new_n395, new_n396, new_n397, new_n398, new_n399,
    new_n400, new_n401, new_n402, new_n403_1, new_n404, new_n405, new_n406,
    new_n407, new_n408, new_n409, new_n410, new_n411, new_n412, new_n413_1,
    new_n414, new_n415, new_n416, new_n417_1, new_n418, new_n419, new_n420,
    new_n421, new_n422, new_n423, new_n424, new_n425, new_n426, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n432, new_n433, new_n434,
    new_n435, new_n436, new_n437, new_n438, new_n439, new_n441, new_n442,
    new_n443, new_n445, new_n446, new_n447, new_n448_1, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454_1, new_n455, new_n456_1,
    new_n457_1, new_n458, new_n459, new_n460, new_n461, new_n462, new_n463,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476_1, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482_1, new_n483, new_n484, new_n485,
    new_n486, new_n487_1, new_n488_1, new_n490, new_n491, new_n492,
    new_n493, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504_1, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516_1, new_n517, new_n518, new_n519, new_n520_1, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530_1, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n542_1, new_n543,
    new_n544_1, new_n545, new_n546, new_n547_1, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n560_1, new_n561, new_n563, new_n564_1,
    new_n565_1, new_n566_1, new_n567_1, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574_1, new_n575, new_n576, new_n577,
    new_n578, new_n579_1, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591_1,
    new_n592, new_n593, new_n594, new_n595, new_n596_1, new_n597, new_n598,
    new_n599, new_n600_1, new_n601_1, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611_1, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617_1, new_n619, new_n620,
    new_n621, new_n622, new_n623_1, new_n624, new_n625, new_n627_1,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635_1,
    new_n636_1, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643_1, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649_1, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661_1, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668_1, new_n669,
    new_n670, new_n671, new_n672, new_n673_1, new_n674, new_n675,
    new_n676_1, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697_1, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708_1, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714_1, new_n715_1, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722_1, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754_1, new_n756, new_n757, new_n758_1, new_n759,
    new_n760_1, new_n761, new_n762, new_n763, new_n765_1, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776_1, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801_1, new_n802, new_n803, new_n805,
    new_n806, new_n807_1, new_n808, new_n811, new_n812, new_n813_1,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824_1, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830_1, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n838, new_n839, new_n840_1, new_n841_1,
    new_n842, new_n843, new_n844, new_n845_1, new_n846, new_n847, new_n848,
    new_n849_1, new_n850_1, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860_1, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878_1, new_n879, new_n880, new_n881, new_n882_1,
    new_n883, new_n884, new_n885, new_n886, new_n887_1, new_n888,
    new_n889_1, new_n890, new_n891, new_n892, new_n893, new_n894_1,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912_1, new_n913, new_n914, new_n915, new_n916,
    new_n917_1, new_n918_1, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937_1, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944_1, new_n945, new_n946_1,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955_1, new_n956, new_n957, new_n959, new_n960, new_n961_1,
    new_n962_1, new_n963, new_n964_1, new_n965, new_n967_1, new_n968,
    new_n969, new_n970, new_n971_1, new_n972, new_n973, new_n974_1,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984_1, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999_1, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016_1, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027_1, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033_1, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039_1, new_n1040, new_n1041, new_n1042, new_n1043_1,
    new_n1044_1, new_n1045, new_n1046, new_n1047_1, new_n1048, new_n1049,
    new_n1050_1, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058_1, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065_1, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087_1, new_n1088_1, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095_1, new_n1096_1, new_n1097_1,
    new_n1098, new_n1099, new_n1100_1, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110_1, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119_1, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125_1, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135_1, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140_1, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150_1, new_n1151,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163_1, new_n1164, new_n1165,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172_1,
    new_n1173, new_n1174, new_n1175_1, new_n1176, new_n1177_1, new_n1178,
    new_n1179, new_n1180_1, new_n1182_1, new_n1183, new_n1184, new_n1185,
    new_n1186_1, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1206,
    new_n1207_1, new_n1208, new_n1209, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224_1, new_n1225, new_n1227_1, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233_1, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238_1, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269_1, new_n1270_1, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279_1, new_n1280, new_n1281_1, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288_1, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297_1, new_n1298, new_n1299_1, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314_1, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322_1, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338_1, new_n1339, new_n1340, new_n1341, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346_1, new_n1347, new_n1348, new_n1349,
    new_n1350, new_n1351, new_n1352, new_n1353_1, new_n1354, new_n1355_1,
    new_n1356, new_n1357_1, new_n1358, new_n1359, new_n1360, new_n1361_1,
    new_n1362_1, new_n1363_1, new_n1364, new_n1365, new_n1366_1, new_n1367,
    new_n1368, new_n1369, new_n1370_1, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1377_1, new_n1378_1, new_n1379, new_n1380, new_n1381,
    new_n1382, new_n1384, new_n1386, new_n1387, new_n1388, new_n1389,
    new_n1390_1, new_n1391_1, new_n1393, new_n1394, new_n1395, new_n1396_1,
    new_n1397, new_n1398, new_n1399, new_n1401, new_n1402_1, new_n1403,
    new_n1404, new_n1405, new_n1406_1, new_n1408_1, new_n1409_1, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1415, new_n1416, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1423, new_n1424,
    new_n1426_1, new_n1427_1, new_n1428, new_n1430, new_n1432, new_n1433,
    new_n1434, new_n1435_1, new_n1436_1, new_n1437, new_n1438, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1448, new_n1449, new_n1450, new_n1451, new_n1452, new_n1453,
    new_n1456, new_n1457, new_n1458, new_n1459, new_n1460, new_n1461,
    new_n1462_1, new_n1464_1, new_n1465, new_n1466, new_n1467, new_n1468,
    new_n1469, new_n1470, new_n1472, new_n1473, new_n1474, new_n1475,
    new_n1476, new_n1477, new_n1478, new_n1479, new_n1480, new_n1481,
    new_n1482, new_n1483, new_n1484, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491_1, new_n1492, new_n1494, new_n1495_1,
    new_n1496, new_n1497, new_n1498_1, new_n1499, new_n1501, new_n1502,
    new_n1503_1, new_n1504, new_n1505, new_n1506, new_n1507, new_n1509,
    new_n1510_1, new_n1511_1, new_n1512, new_n1513, new_n1514, new_n1516,
    new_n1517, new_n1518_1, new_n1519_1, new_n1520, new_n1521, new_n1524,
    new_n1525, new_n1526, new_n1528, new_n1529, new_n1530, new_n1531,
    new_n1532, new_n1533, new_n1534_1, new_n1536, new_n1537, new_n1538,
    new_n1539, new_n1540_1, new_n1541, new_n1543_1, new_n1544, new_n1545,
    new_n1546, new_n1547, new_n1548, new_n1551, new_n1552, new_n1553_1,
    new_n1554, new_n1555, new_n1556, new_n1557, new_n1559, new_n1560,
    new_n1561, new_n1562, new_n1563, new_n1565, new_n1566, new_n1567,
    new_n1568_1, new_n1569, new_n1570, new_n1571, new_n1573, new_n1574,
    new_n1575_1, new_n1576, new_n1577, new_n1578, new_n1581, new_n1582,
    new_n1583, new_n1584_1, new_n1585, new_n1586, new_n1587_1, new_n1589,
    new_n1590, new_n1591, new_n1592, new_n1593, new_n1594, new_n1595;
  assign new_n302 = ~n186 & n560;
  assign new_n303 = ~n261 & n579;
  assign new_n304 = n504 & n917;
  assign new_n305 = ~n504 & n1553;
  assign new_n306 = ~new_n304 & ~new_n305;
  assign new_n307_1 = n1755 & ~new_n306;
  assign new_n308 = ~n1755 & new_n306;
  assign new_n309 = ~new_n307_1 & ~new_n308;
  assign new_n310 = n504 & n887;
  assign new_n311 = ~n504 & n1729;
  assign new_n312 = ~new_n310 & ~new_n311;
  assign new_n313 = n1135 & ~new_n312;
  assign new_n314 = ~n1135 & new_n312;
  assign new_n315_1 = ~new_n313 & ~new_n314;
  assign new_n316 = n504 & n1436;
  assign new_n317 = n319 & ~n504;
  assign new_n318 = ~new_n316 & ~new_n317;
  assign new_n319_1 = n1402 & ~new_n318;
  assign new_n320_1 = ~n1402 & new_n318;
  assign new_n321_1 = ~new_n319_1 & ~new_n320_1;
  assign new_n322 = n504 & n961;
  assign new_n323 = ~n504 & n1238;
  assign new_n324 = ~new_n322 & ~new_n323;
  assign new_n325 = ~n1100 & new_n324;
  assign new_n326_1 = n1100 & ~new_n324;
  assign new_n327 = ~new_n325 & ~new_n326_1;
  assign new_n328 = n504 & n1632;
  assign new_n329 = ~n504 & n1498;
  assign new_n330 = ~new_n328 & ~new_n329;
  assign new_n331 = n1039 & ~new_n330;
  assign new_n332 = ~n1039 & new_n330;
  assign new_n333 = ~new_n331 & ~new_n332;
  assign new_n334 = n504 & n1396;
  assign new_n335_1 = ~n504 & n617;
  assign new_n336 = ~new_n334 & ~new_n335_1;
  assign new_n337_1 = n39 & ~new_n336;
  assign new_n338 = ~n39 & new_n336;
  assign new_n339 = ~new_n337_1 & ~new_n338;
  assign new_n340 = new_n333 & new_n339;
  assign new_n341 = new_n327 & new_n340;
  assign new_n342_1 = new_n321_1 & new_n341;
  assign new_n343 = new_n315_1 & new_n342_1;
  assign new_n344 = new_n333 & new_n337_1;
  assign new_n345 = ~new_n326_1 & ~new_n331;
  assign new_n346 = ~new_n344 & new_n345;
  assign new_n347 = ~new_n325 & ~new_n346;
  assign new_n348 = ~new_n319_1 & ~new_n347;
  assign new_n349 = ~new_n320_1 & ~new_n348;
  assign new_n350 = ~new_n313 & ~new_n349;
  assign new_n351 = ~new_n314 & ~new_n350;
  assign new_n352 = ~new_n343 & ~new_n351;
  assign new_n353 = ~n1279 & ~new_n351;
  assign new_n354 = ~new_n352 & ~new_n353;
  assign new_n355 = new_n309 & new_n354;
  assign new_n356 = ~new_n309 & ~new_n354;
  assign new_n357_1 = ~new_n355 & ~new_n356;
  assign new_n358 = new_n303 & new_n357_1;
  assign new_n359 = ~n261 & ~n579;
  assign new_n360 = n1288 & n1553;
  assign new_n361_1 = n721 & ~n1553;
  assign new_n362 = n1755 & ~new_n361_1;
  assign new_n363 = ~new_n360 & new_n362;
  assign new_n364 = ~n1519 & ~n1553;
  assign new_n365 = ~n77 & n1553;
  assign new_n366 = ~new_n364 & ~new_n365;
  assign new_n367 = ~n1755 & new_n366;
  assign new_n368 = ~new_n363 & ~new_n367;
  assign new_n369 = new_n359 & new_n368;
  assign new_n370_1 = n261 & ~n579;
  assign new_n371_1 = n984 & new_n370_1;
  assign new_n372 = ~new_n369 & ~new_n371_1;
  assign n370 = ~new_n358 & new_n372;
  assign new_n374 = new_n302 & ~n370;
  assign new_n375_1 = n186 & n560;
  assign new_n376 = n19 & new_n375_1;
  assign new_n377_1 = n186 & ~n560;
  assign new_n378_1 = n955 & new_n377_1;
  assign new_n379_1 = ~n186 & ~n560;
  assign new_n380_1 = n600 & n894;
  assign new_n381_1 = ~n600 & n946;
  assign new_n382 = ~new_n380_1 & ~new_n381_1;
  assign new_n383 = n1406 & ~new_n382;
  assign new_n384_1 = ~n1406 & new_n382;
  assign new_n385 = ~new_n383 & ~new_n384_1;
  assign new_n386_1 = n600 & ~n1568;
  assign new_n387_1 = n238 & ~new_n386_1;
  assign new_n388 = ~n238 & new_n386_1;
  assign new_n389_1 = ~new_n387_1 & ~new_n388;
  assign new_n390 = n600 & n1707;
  assign new_n391 = n380 & ~n600;
  assign new_n392 = ~new_n390 & ~new_n391;
  assign new_n393 = n1391 & ~new_n392;
  assign new_n394 = ~n1391 & new_n392;
  assign new_n395 = ~new_n393 & ~new_n394;
  assign new_n396 = new_n389_1 & new_n395;
  assign new_n397 = n600 & n937;
  assign new_n398 = ~n600 & n1435;
  assign new_n399 = ~new_n397 & ~new_n398;
  assign new_n400 = n1016 & ~new_n399;
  assign new_n401 = ~n1016 & new_n399;
  assign new_n402 = ~new_n400 & ~new_n401;
  assign new_n403_1 = n448 & n600;
  assign new_n404 = ~n600 & n1043;
  assign new_n405 = ~new_n403_1 & ~new_n404;
  assign new_n406 = ~n1125 & new_n405;
  assign new_n407 = n1125 & ~new_n405;
  assign new_n408 = n600 & n1338;
  assign new_n409 = ~n600 & n1515;
  assign new_n410 = ~new_n408 & ~new_n409;
  assign new_n411 = ~new_n407 & new_n410;
  assign new_n412 = ~new_n406 & new_n411;
  assign new_n413_1 = new_n402 & new_n412;
  assign new_n414 = new_n396 & new_n413_1;
  assign new_n415 = n1788 & new_n414;
  assign new_n416 = ~new_n406 & ~new_n411;
  assign new_n417_1 = ~new_n400 & ~new_n416;
  assign new_n418 = ~new_n401 & ~new_n417_1;
  assign new_n419 = ~new_n387_1 & ~new_n418;
  assign new_n420 = ~new_n388 & ~new_n419;
  assign new_n421 = ~new_n393 & ~new_n420;
  assign new_n422 = ~new_n394 & ~new_n421;
  assign new_n423 = ~new_n415 & ~new_n422;
  assign new_n424 = ~new_n385 & ~new_n423;
  assign new_n425 = new_n385 & new_n423;
  assign new_n426 = ~new_n424 & ~new_n425;
  assign new_n427 = new_n303 & ~new_n426;
  assign new_n428 = ~n946 & ~n1227;
  assign new_n429 = ~n591 & n946;
  assign new_n430 = n1406 & ~new_n429;
  assign new_n431 = ~new_n428 & new_n430;
  assign new_n432 = n807 & n946;
  assign new_n433 = n714 & ~n946;
  assign new_n434 = ~new_n432 & ~new_n433;
  assign new_n435 = ~n1406 & new_n434;
  assign new_n436 = ~new_n431 & ~new_n435;
  assign new_n437 = new_n359 & new_n436;
  assign new_n438 = n1097 & new_n370_1;
  assign new_n439 = ~new_n437 & ~new_n438;
  assign n964 = ~new_n427 & new_n439;
  assign new_n441 = new_n379_1 & ~n964;
  assign new_n442 = ~new_n378_1 & ~new_n441;
  assign new_n443 = ~new_n376 & new_n442;
  assign n18 = new_n374 | ~new_n443;
  assign new_n445 = n228 & ~n1205;
  assign new_n446 = n1279 & new_n339;
  assign new_n447 = ~new_n337_1 & ~new_n446;
  assign new_n448_1 = new_n333 & ~new_n447;
  assign new_n449 = ~new_n333 & new_n447;
  assign new_n450 = ~new_n448_1 & ~new_n449;
  assign new_n451 = new_n303 & new_n450;
  assign new_n452 = n1288 & n1498;
  assign new_n453 = n721 & ~n1498;
  assign new_n454_1 = n1039 & ~new_n453;
  assign new_n455 = ~new_n452 & new_n454_1;
  assign new_n456_1 = ~n1498 & ~n1519;
  assign new_n457_1 = ~n77 & n1498;
  assign new_n458 = ~new_n456_1 & ~new_n457_1;
  assign new_n459 = ~n1039 & new_n458;
  assign new_n460 = ~new_n455 & ~new_n459;
  assign new_n461 = new_n359 & new_n460;
  assign new_n462 = n1633 & new_n370_1;
  assign new_n463 = ~new_n461 & ~new_n462;
  assign n1346 = ~new_n451 & new_n463;
  assign new_n465 = new_n445 & ~n1346;
  assign new_n466 = ~n228 & n1205;
  assign new_n467 = n1180 & new_n466;
  assign new_n468 = n228 & n1205;
  assign new_n469 = n7 & new_n468;
  assign new_n470 = ~n228 & ~n1205;
  assign new_n471 = ~new_n406 & ~new_n407;
  assign new_n472 = ~n1788 & new_n410;
  assign new_n473 = ~new_n471 & new_n472;
  assign new_n474 = new_n471 & ~new_n472;
  assign new_n475 = new_n303 & ~new_n474;
  assign new_n476_1 = ~new_n473 & new_n475;
  assign new_n477 = n668 & new_n370_1;
  assign new_n478 = n1043 & n1288;
  assign new_n479 = n721 & ~n1043;
  assign new_n480 = n1125 & ~new_n479;
  assign new_n481 = ~new_n478 & new_n480;
  assign new_n482_1 = ~n1043 & ~n1519;
  assign new_n483 = ~n77 & n1043;
  assign new_n484 = ~new_n482_1 & ~new_n483;
  assign new_n485 = ~n1125 & new_n484;
  assign new_n486 = ~new_n481 & ~new_n485;
  assign new_n487_1 = new_n359 & new_n486;
  assign new_n488_1 = ~new_n477 & ~new_n487_1;
  assign n168 = ~new_n476_1 & new_n488_1;
  assign new_n490 = new_n470 & ~n168;
  assign new_n491 = ~new_n469 & ~new_n490;
  assign new_n492 = ~new_n467 & new_n491;
  assign new_n493 = ~new_n465 & new_n492;
  assign n56 = n1534 & ~new_n493;
  assign n67 = ~n544 & n1471;
  assign new_n496 = n600 & n1426;
  assign new_n497 = ~n600 & n966;
  assign new_n498 = ~new_n496 & ~new_n497;
  assign new_n499 = n326 & ~new_n498;
  assign new_n500 = ~n326 & new_n498;
  assign new_n501 = ~new_n499 & ~new_n500;
  assign new_n502 = new_n383 & new_n501;
  assign new_n503 = ~new_n499 & ~new_n502;
  assign new_n504_1 = new_n385 & new_n501;
  assign new_n505 = ~new_n423 & new_n504_1;
  assign new_n506 = new_n503 & ~new_n505;
  assign new_n507 = n600 & n971;
  assign new_n508 = ~n600 & n1518;
  assign new_n509 = ~new_n507 & ~new_n508;
  assign new_n510 = ~new_n506 & ~new_n509;
  assign new_n511 = new_n503 & new_n509;
  assign new_n512 = ~new_n505 & new_n511;
  assign new_n513 = ~new_n510 & ~new_n512;
  assign new_n514 = new_n303 & ~new_n513;
  assign new_n515 = n591 & n1518;
  assign new_n516_1 = n1227 & ~n1518;
  assign new_n517 = ~new_n515 & ~new_n516_1;
  assign new_n518 = new_n359 & new_n517;
  assign new_n519 = n813 & new_n370_1;
  assign new_n520_1 = ~new_n518 & ~new_n519;
  assign n75 = ~new_n514 & new_n520_1;
  assign new_n522 = ~new_n341 & ~new_n347;
  assign new_n523 = ~n1279 & ~new_n347;
  assign new_n524 = ~new_n522 & ~new_n523;
  assign new_n525 = new_n321_1 & new_n524;
  assign new_n526 = ~new_n321_1 & ~new_n524;
  assign new_n527 = ~new_n525 & ~new_n526;
  assign new_n528 = new_n303 & new_n527;
  assign new_n529 = n319 & n1288;
  assign new_n530_1 = ~n319 & n721;
  assign new_n531 = n1402 & ~new_n530_1;
  assign new_n532 = ~new_n529 & new_n531;
  assign new_n533 = ~n319 & ~n1519;
  assign new_n534 = ~n77 & n319;
  assign new_n535 = ~new_n533 & ~new_n534;
  assign new_n536 = ~n1402 & new_n535;
  assign new_n537 = ~new_n532 & ~new_n536;
  assign new_n538 = new_n359 & new_n537;
  assign new_n539 = n999 & new_n370_1;
  assign new_n540 = ~new_n538 & ~new_n539;
  assign n1710 = ~new_n528 & new_n540;
  assign new_n542_1 = new_n302 & ~n1710;
  assign new_n543 = n1540 & new_n377_1;
  assign new_n544_1 = n565 & new_n375_1;
  assign new_n545 = ~new_n407 & ~new_n474;
  assign new_n546 = new_n402 & ~new_n545;
  assign new_n547_1 = ~new_n400 & ~new_n546;
  assign new_n548 = ~new_n389_1 & new_n547_1;
  assign new_n549 = new_n389_1 & ~new_n547_1;
  assign new_n550 = ~new_n548 & ~new_n549;
  assign new_n551 = new_n303 & new_n550;
  assign new_n552 = n238 & n1288;
  assign new_n553 = ~n77 & ~n238;
  assign new_n554 = ~new_n552 & ~new_n553;
  assign new_n555 = new_n359 & ~new_n554;
  assign new_n556 = n1361 & new_n370_1;
  assign new_n557 = ~new_n555 & ~new_n556;
  assign n487 = ~new_n551 & new_n557;
  assign new_n559 = new_n379_1 & ~n487;
  assign new_n560_1 = ~new_n544_1 & ~new_n559;
  assign new_n561 = ~new_n543 & new_n560_1;
  assign n83 = new_n542_1 | ~new_n561;
  assign new_n563 = n504 & n1408;
  assign new_n564_1 = ~n504 & n708;
  assign new_n565_1 = ~new_n563 & ~new_n564_1;
  assign new_n566_1 = n60 & ~new_n565_1;
  assign new_n567_1 = ~n60 & new_n565_1;
  assign new_n568 = ~new_n566_1 & ~new_n567_1;
  assign new_n569 = n504 & n801;
  assign new_n570 = ~n504 & n1660;
  assign new_n571 = ~new_n569 & ~new_n570;
  assign new_n572 = ~n1575 & new_n571;
  assign new_n573 = n1575 & ~new_n571;
  assign new_n574_1 = ~new_n572 & ~new_n573;
  assign new_n575 = n504 & n1485;
  assign new_n576 = ~n504 & n1172;
  assign new_n577 = ~new_n575 & ~new_n576;
  assign new_n578 = n697 & ~new_n577;
  assign new_n579_1 = ~n697 & new_n577;
  assign new_n580 = ~new_n578 & ~new_n579_1;
  assign new_n581 = new_n309 & new_n580;
  assign new_n582 = new_n574_1 & new_n581;
  assign new_n583 = new_n307_1 & new_n580;
  assign new_n584 = ~new_n578 & ~new_n583;
  assign new_n585 = ~new_n572 & ~new_n584;
  assign new_n586 = ~new_n573 & ~new_n585;
  assign new_n587 = ~new_n582 & new_n586;
  assign new_n588 = ~new_n354 & new_n586;
  assign new_n589 = ~new_n587 & ~new_n588;
  assign new_n590 = ~new_n568 & new_n589;
  assign new_n591_1 = new_n568 & ~new_n589;
  assign new_n592 = ~new_n590 & ~new_n591_1;
  assign new_n593 = new_n303 & ~new_n592;
  assign new_n594 = ~n708 & ~n1227;
  assign new_n595 = ~n591 & n708;
  assign new_n596_1 = n60 & ~new_n595;
  assign new_n597 = ~new_n594 & new_n596_1;
  assign new_n598 = n708 & n807;
  assign new_n599 = ~n708 & n714;
  assign new_n600_1 = ~new_n598 & ~new_n599;
  assign new_n601_1 = ~n60 & new_n600_1;
  assign new_n602 = ~new_n597 & ~new_n601_1;
  assign new_n603 = new_n359 & new_n602;
  assign new_n604 = n850 & new_n370_1;
  assign new_n605 = ~new_n603 & ~new_n604;
  assign n123 = ~new_n593 & new_n605;
  assign new_n607 = new_n302 & ~n123;
  assign new_n608 = n1177 & new_n377_1;
  assign new_n609 = n754 & new_n375_1;
  assign new_n610 = n389 & n600;
  assign new_n611_1 = n288 & ~n600;
  assign new_n612 = ~new_n610 & ~new_n611_1;
  assign new_n613 = new_n509 & new_n612;
  assign new_n614 = ~new_n509 & ~new_n612;
  assign new_n615 = ~new_n613 & ~new_n614;
  assign new_n616 = new_n506 & ~new_n615;
  assign new_n617_1 = ~new_n506 & ~new_n612;
  assign n1793 = ~new_n616 & ~new_n617_1;
  assign new_n619 = new_n303 & ~n1793;
  assign new_n620 = n482 & new_n370_1;
  assign new_n621 = n288 & n807;
  assign new_n622 = ~n288 & n714;
  assign new_n623_1 = ~new_n621 & ~new_n622;
  assign new_n624 = new_n359 & ~new_n623_1;
  assign new_n625 = ~new_n620 & ~new_n624;
  assign n1027 = ~new_n619 & new_n625;
  assign new_n627_1 = new_n379_1 & ~n1027;
  assign new_n628 = ~new_n609 & ~new_n627_1;
  assign new_n629 = ~new_n608 & new_n628;
  assign n101 = new_n607 | ~new_n629;
  assign new_n631 = n1172 & n1288;
  assign new_n632 = n721 & ~n1172;
  assign new_n633 = n697 & ~new_n632;
  assign new_n634 = ~new_n631 & new_n633;
  assign new_n635_1 = ~n1172 & ~n1519;
  assign new_n636_1 = ~n77 & n1172;
  assign new_n637 = ~new_n635_1 & ~new_n636_1;
  assign new_n638 = ~n697 & new_n637;
  assign new_n639 = ~new_n634 & ~new_n638;
  assign new_n640 = n1288 & n1729;
  assign new_n641 = n721 & ~n1729;
  assign new_n642 = n1135 & ~new_n641;
  assign new_n643_1 = ~new_n640 & new_n642;
  assign new_n644 = ~n1519 & ~n1729;
  assign new_n645 = ~n77 & n1729;
  assign new_n646 = ~new_n644 & ~new_n645;
  assign new_n647 = ~n1135 & new_n646;
  assign new_n648 = ~new_n643_1 & ~new_n647;
  assign new_n649_1 = ~new_n639 & ~new_n648;
  assign new_n650 = n1238 & n1288;
  assign new_n651 = n721 & ~n1238;
  assign new_n652 = n1100 & ~new_n651;
  assign new_n653 = ~new_n650 & new_n652;
  assign new_n654 = ~n1238 & ~n1519;
  assign new_n655 = ~n77 & n1238;
  assign new_n656 = ~new_n654 & ~new_n655;
  assign new_n657 = ~n1100 & new_n656;
  assign new_n658 = ~new_n653 & ~new_n657;
  assign new_n659 = n1288 & n1660;
  assign new_n660 = n721 & ~n1660;
  assign new_n661_1 = n1575 & ~new_n660;
  assign new_n662 = ~new_n659 & new_n661_1;
  assign new_n663 = ~n1519 & ~n1660;
  assign new_n664 = ~n77 & n1660;
  assign new_n665 = ~new_n663 & ~new_n664;
  assign new_n666 = ~n1575 & new_n665;
  assign new_n667 = ~new_n662 & ~new_n666;
  assign new_n668_1 = ~new_n658 & ~new_n667;
  assign new_n669 = ~new_n460 & ~new_n602;
  assign new_n670 = new_n668_1 & new_n669;
  assign new_n671 = ~new_n368 & ~new_n537;
  assign new_n672 = n617 & n1288;
  assign new_n673_1 = ~n617 & n721;
  assign new_n674 = n39 & ~new_n673_1;
  assign new_n675 = ~new_n672 & new_n674;
  assign new_n676_1 = ~n617 & ~n1519;
  assign new_n677 = ~n77 & n617;
  assign new_n678 = ~new_n676_1 & ~new_n677;
  assign new_n679 = ~n39 & new_n678;
  assign new_n680 = ~new_n675 & ~new_n679;
  assign new_n681 = new_n671 & ~new_n680;
  assign new_n682 = new_n670 & new_n681;
  assign n107 = new_n649_1 & new_n682;
  assign n117 = ~n601 | ~n841;
  assign new_n685 = new_n504_1 & new_n509;
  assign new_n686 = new_n422 & new_n685;
  assign new_n687 = new_n511 & new_n612;
  assign n130 = new_n686 | ~new_n687;
  assign new_n689 = n378 & ~n627;
  assign new_n690 = ~n123 & new_n689;
  assign new_n691 = ~n378 & ~n627;
  assign new_n692 = ~n1027 & new_n691;
  assign new_n693 = n378 & n627;
  assign new_n694 = n830 & new_n693;
  assign new_n695 = ~n378 & n627;
  assign new_n696 = n1033 & new_n695;
  assign new_n697_1 = ~new_n694 & ~new_n696;
  assign new_n698 = ~new_n692 & new_n697_1;
  assign new_n699 = ~new_n690 & new_n698;
  assign n158 = n1534 & ~new_n699;
  assign new_n701 = n1788 & ~new_n410;
  assign new_n702 = ~new_n472 & ~new_n701;
  assign new_n703 = ~new_n402 & new_n545;
  assign new_n704 = ~new_n546 & ~new_n703;
  assign new_n705 = new_n471 & ~new_n704;
  assign new_n706 = new_n702 & new_n705;
  assign new_n707 = ~new_n383 & new_n423;
  assign new_n708_1 = ~new_n384_1 & ~new_n707;
  assign new_n709 = ~new_n501 & new_n708_1;
  assign new_n710 = new_n501 & ~new_n708_1;
  assign new_n711 = ~new_n709 & ~new_n710;
  assign new_n712 = ~new_n550 & new_n711;
  assign new_n713 = new_n706 & new_n712;
  assign new_n714_1 = ~new_n387_1 & ~new_n549;
  assign new_n715_1 = ~new_n395 & new_n714_1;
  assign new_n716 = new_n395 & ~new_n714_1;
  assign new_n717 = ~new_n715_1 & ~new_n716;
  assign new_n718 = new_n426 & ~new_n717;
  assign new_n719 = n1793 & new_n718;
  assign new_n720 = new_n513 & new_n719;
  assign n165 = new_n713 & new_n720;
  assign new_n722_1 = ~new_n308 & new_n580;
  assign new_n723 = ~new_n578 & ~new_n722_1;
  assign new_n724 = ~new_n354 & new_n584;
  assign new_n725 = ~new_n723 & ~new_n724;
  assign new_n726 = ~new_n574_1 & new_n725;
  assign new_n727 = new_n574_1 & ~new_n725;
  assign new_n728 = ~new_n726 & ~new_n727;
  assign new_n729 = new_n303 & ~new_n728;
  assign new_n730 = new_n359 & new_n667;
  assign new_n731 = n386 & new_n370_1;
  assign new_n732 = ~new_n730 & ~new_n731;
  assign n1087 = ~new_n729 & new_n732;
  assign new_n734 = new_n302 & ~n1087;
  assign new_n735 = n384 & new_n377_1;
  assign new_n736 = n297 & new_n375_1;
  assign new_n737 = new_n379_1 & ~n75;
  assign new_n738 = ~new_n736 & ~new_n737;
  assign new_n739 = ~new_n735 & new_n738;
  assign n211 = new_n734 | ~new_n739;
  assign new_n741 = ~n370 & new_n689;
  assign new_n742 = ~n964 & new_n691;
  assign new_n743 = n715 & new_n693;
  assign new_n744 = n128 & new_n695;
  assign new_n745 = ~new_n743 & ~new_n744;
  assign new_n746 = ~new_n742 & new_n745;
  assign new_n747 = ~new_n741 & new_n746;
  assign n222 = n1534 & ~new_n747;
  assign new_n749 = new_n504_1 & new_n613;
  assign n235 = new_n414 & new_n749;
  assign new_n751 = n1219 & ~n1281;
  assign new_n752 = n1088 & n1281;
  assign new_n753 = ~n117 & ~new_n752;
  assign new_n754_1 = ~new_n751 & new_n753;
  assign n245 = n1613 & ~new_n754_1;
  assign new_n756 = ~new_n319_1 & ~new_n525;
  assign new_n757 = ~new_n315_1 & new_n756;
  assign new_n758_1 = new_n315_1 & ~new_n756;
  assign new_n759 = ~new_n757 & ~new_n758_1;
  assign new_n760_1 = new_n303 & new_n759;
  assign new_n761 = new_n359 & new_n648;
  assign new_n762 = n157 & new_n370_1;
  assign new_n763 = ~new_n761 & ~new_n762;
  assign n1631 = ~new_n760_1 & new_n763;
  assign new_n765_1 = new_n689 & ~n1631;
  assign new_n766 = new_n303 & new_n717;
  assign new_n767 = n380 & n1288;
  assign new_n768 = ~n380 & n721;
  assign new_n769 = n1391 & ~new_n768;
  assign new_n770 = ~new_n767 & new_n769;
  assign new_n771 = ~n380 & ~n1519;
  assign new_n772 = ~n77 & n380;
  assign new_n773 = ~new_n771 & ~new_n772;
  assign new_n774 = ~n1391 & new_n773;
  assign new_n775 = ~new_n770 & ~new_n774;
  assign new_n776_1 = new_n359 & new_n775;
  assign new_n777 = n1095 & new_n370_1;
  assign new_n778 = ~new_n776_1 & ~new_n777;
  assign n1495 = ~new_n766 & new_n778;
  assign new_n780 = new_n691 & ~n1495;
  assign new_n781 = n236 & new_n693;
  assign new_n782 = n1743 & new_n695;
  assign new_n783 = ~new_n781 & ~new_n782;
  assign new_n784 = ~new_n780 & new_n783;
  assign new_n785 = ~new_n765_1 & new_n784;
  assign n249 = n1534 & ~new_n785;
  assign new_n787 = ~n1279 & ~new_n339;
  assign new_n788 = ~new_n446 & ~new_n787;
  assign new_n789 = new_n303 & new_n788;
  assign new_n790 = new_n359 & new_n680;
  assign new_n791 = n190 & new_n370_1;
  assign new_n792 = ~new_n790 & ~new_n791;
  assign n259 = ~new_n789 & new_n792;
  assign new_n794 = n758 & new_n693;
  assign new_n795 = new_n689 & ~n259;
  assign new_n796 = n1675 & new_n695;
  assign new_n797 = new_n303 & ~new_n702;
  assign new_n798 = n591 & n1515;
  assign new_n799 = n1227 & ~n1515;
  assign new_n800 = ~new_n798 & ~new_n799;
  assign new_n801_1 = new_n359 & new_n800;
  assign new_n802 = n1753 & new_n370_1;
  assign new_n803 = ~new_n801_1 & ~new_n802;
  assign n454 = ~new_n797 & new_n803;
  assign new_n805 = new_n691 & ~n454;
  assign new_n806 = ~new_n796 & ~new_n805;
  assign new_n807_1 = ~new_n795 & new_n806;
  assign new_n808 = ~new_n794 & new_n807_1;
  assign n262 = n1534 & ~new_n808;
  assign n1491 = ~n119 | ~n1768;
  assign new_n811 = ~new_n382 & new_n498;
  assign new_n812 = new_n382 & ~new_n498;
  assign new_n813_1 = ~new_n811 & ~new_n812;
  assign new_n814 = new_n615 & ~new_n813_1;
  assign new_n815 = ~new_n615 & new_n813_1;
  assign new_n816 = ~new_n814 & ~new_n815;
  assign new_n817 = new_n399 & new_n816;
  assign new_n818 = ~new_n399 & ~new_n816;
  assign new_n819 = ~new_n817 & ~new_n818;
  assign new_n820 = ~n600 & ~n643;
  assign new_n821 = ~n541 & n600;
  assign new_n822 = ~new_n820 & ~new_n821;
  assign new_n823 = ~new_n410 & new_n822;
  assign new_n824_1 = new_n410 & ~new_n822;
  assign new_n825 = ~new_n823 & ~new_n824_1;
  assign new_n826 = ~new_n386_1 & new_n392;
  assign new_n827 = n1707 & new_n386_1;
  assign new_n828 = ~new_n826 & ~new_n827;
  assign new_n829 = new_n405 & new_n828;
  assign new_n830_1 = ~new_n405 & ~new_n828;
  assign new_n831 = ~new_n829 & ~new_n830_1;
  assign new_n832 = ~new_n825 & new_n831;
  assign new_n833 = new_n825 & ~new_n831;
  assign new_n834 = ~new_n832 & ~new_n833;
  assign new_n835 = new_n819 & ~new_n834;
  assign new_n836 = ~new_n819 & new_n834;
  assign n320 = new_n835 | new_n836;
  assign new_n838 = ~n1491 & ~n320;
  assign new_n839 = ~n504 & ~n1674;
  assign new_n840_1 = ~n64 & n504;
  assign new_n841_1 = ~new_n839 & ~new_n840_1;
  assign new_n842 = ~new_n565_1 & new_n841_1;
  assign new_n843 = new_n565_1 & ~new_n841_1;
  assign new_n844 = ~new_n842 & ~new_n843;
  assign new_n845_1 = new_n306 & new_n312;
  assign new_n846 = ~new_n306 & ~new_n312;
  assign new_n847 = ~new_n845_1 & ~new_n846;
  assign new_n848 = new_n844 & new_n847;
  assign new_n849_1 = ~new_n844 & ~new_n847;
  assign new_n850_1 = ~new_n848 & ~new_n849_1;
  assign new_n851 = new_n318 & new_n324;
  assign new_n852 = ~new_n318 & ~new_n324;
  assign new_n853 = ~new_n851 & ~new_n852;
  assign new_n854 = ~new_n571 & new_n577;
  assign new_n855 = new_n571 & ~new_n577;
  assign new_n856 = ~new_n854 & ~new_n855;
  assign new_n857 = ~new_n853 & new_n856;
  assign new_n858 = new_n853 & ~new_n856;
  assign new_n859 = ~new_n857 & ~new_n858;
  assign new_n860_1 = new_n330 & new_n336;
  assign new_n861 = ~new_n330 & ~new_n336;
  assign new_n862 = ~new_n860_1 & ~new_n861;
  assign new_n863 = new_n859 & ~new_n862;
  assign new_n864 = ~new_n859 & new_n862;
  assign new_n865 = ~new_n863 & ~new_n864;
  assign new_n866 = ~new_n850_1 & ~new_n865;
  assign new_n867 = new_n850_1 & new_n865;
  assign n547 = new_n866 | new_n867;
  assign new_n869 = ~n1660 & n1729;
  assign new_n870 = n1660 & ~n1729;
  assign new_n871 = ~new_n869 & ~new_n870;
  assign new_n872 = n708 & n1553;
  assign new_n873 = ~n708 & ~n1553;
  assign new_n874 = ~new_n872 & ~new_n873;
  assign new_n875 = ~new_n871 & new_n874;
  assign new_n876 = new_n871 & ~new_n874;
  assign new_n877 = ~new_n875 & ~new_n876;
  assign new_n878_1 = ~n1498 & n1674;
  assign new_n879 = n1498 & ~n1674;
  assign new_n880 = ~new_n878_1 & ~new_n879;
  assign new_n881 = n617 & n1238;
  assign new_n882_1 = ~n617 & ~n1238;
  assign new_n883 = ~new_n881 & ~new_n882_1;
  assign new_n884 = new_n880 & new_n883;
  assign new_n885 = ~new_n880 & ~new_n883;
  assign new_n886 = ~new_n884 & ~new_n885;
  assign new_n887_1 = n319 & n1172;
  assign new_n888 = ~n319 & ~n1172;
  assign new_n889_1 = ~new_n887_1 & ~new_n888;
  assign new_n890 = new_n886 & ~new_n889_1;
  assign new_n891 = ~new_n886 & new_n889_1;
  assign new_n892 = ~new_n890 & ~new_n891;
  assign new_n893 = ~new_n877 & ~new_n892;
  assign new_n894_1 = new_n877 & new_n892;
  assign n878 = ~new_n893 & ~new_n894_1;
  assign new_n896 = ~n1435 & n1518;
  assign new_n897 = n1435 & ~n1518;
  assign new_n898 = ~new_n896 & ~new_n897;
  assign new_n899 = n288 & n1043;
  assign new_n900 = ~n288 & ~n1043;
  assign new_n901 = ~new_n899 & ~new_n900;
  assign new_n902 = new_n898 & new_n901;
  assign new_n903 = ~new_n898 & ~new_n901;
  assign new_n904 = ~new_n902 & ~new_n903;
  assign new_n905 = n380 & n643;
  assign new_n906 = ~n380 & ~n643;
  assign new_n907 = ~new_n905 & ~new_n906;
  assign new_n908 = n1515 & ~new_n907;
  assign new_n909 = ~n1515 & new_n907;
  assign new_n910 = ~new_n908 & ~new_n909;
  assign new_n911 = n946 & n966;
  assign new_n912_1 = ~n946 & ~n966;
  assign new_n913 = ~new_n911 & ~new_n912_1;
  assign new_n914 = new_n910 & ~new_n913;
  assign new_n915 = ~new_n910 & new_n913;
  assign new_n916 = ~new_n914 & ~new_n915;
  assign new_n917_1 = ~new_n904 & ~new_n916;
  assign new_n918_1 = new_n904 & new_n916;
  assign n1511 = ~new_n917_1 & ~new_n918_1;
  assign n1047 = n92 & n457;
  assign new_n921 = n516 & n1047;
  assign new_n922 = n1503 & new_n921;
  assign new_n923 = ~n1511 & new_n922;
  assign new_n924 = ~n878 & new_n923;
  assign new_n925 = ~n547 & new_n924;
  assign n264 = new_n838 & new_n925;
  assign new_n927 = ~new_n307_1 & ~new_n354;
  assign new_n928 = ~new_n308 & ~new_n927;
  assign new_n929 = ~new_n580 & ~new_n928;
  assign new_n930 = new_n580 & new_n928;
  assign new_n931 = ~new_n929 & ~new_n930;
  assign new_n932 = new_n303 & new_n931;
  assign new_n933 = new_n359 & new_n639;
  assign new_n934 = n779 & new_n370_1;
  assign new_n935 = ~new_n933 & ~new_n934;
  assign n456 = ~new_n932 & new_n935;
  assign new_n937_1 = new_n445 & ~n456;
  assign new_n938 = new_n303 & ~new_n711;
  assign new_n939 = ~n966 & ~n1227;
  assign new_n940 = ~n591 & n966;
  assign new_n941 = n326 & ~new_n940;
  assign new_n942 = ~new_n939 & new_n941;
  assign new_n943 = n807 & n966;
  assign new_n944_1 = n714 & ~n966;
  assign new_n945 = ~new_n943 & ~new_n944_1;
  assign new_n946_1 = ~n326 & new_n945;
  assign new_n947 = ~new_n942 & ~new_n946_1;
  assign new_n948 = new_n359 & new_n947;
  assign new_n949 = n1182 & new_n370_1;
  assign new_n950 = ~new_n948 & ~new_n949;
  assign n882 = ~new_n938 & new_n950;
  assign new_n952 = new_n470 & ~n882;
  assign new_n953 = n270 & new_n466;
  assign new_n954 = n335 & new_n468;
  assign new_n955_1 = ~new_n953 & ~new_n954;
  assign new_n956 = ~new_n952 & new_n955_1;
  assign new_n957 = ~new_n937_1 & new_n956;
  assign n315 = n1534 & ~new_n957;
  assign new_n959 = n1675 & new_n466;
  assign new_n960 = new_n445 & ~n259;
  assign new_n961_1 = n758 & new_n468;
  assign new_n962_1 = new_n470 & ~n454;
  assign new_n963 = ~new_n961_1 & ~new_n962_1;
  assign new_n964_1 = ~new_n960 & new_n963;
  assign new_n965 = ~new_n959 & new_n964_1;
  assign n337 = n1534 & ~new_n965;
  assign new_n967_1 = new_n339 & new_n349;
  assign new_n968 = ~new_n339 & ~new_n349;
  assign new_n969 = ~new_n967_1 & ~new_n968;
  assign new_n970 = ~new_n327 & new_n969;
  assign new_n971_1 = new_n327 & ~new_n969;
  assign new_n972 = ~new_n970 & ~new_n971_1;
  assign new_n973 = ~new_n325 & ~new_n337_1;
  assign new_n974_1 = ~new_n345 & new_n973;
  assign new_n975 = new_n337_1 & ~new_n347;
  assign new_n976 = ~new_n974_1 & ~new_n975;
  assign new_n977 = ~new_n331 & ~new_n344;
  assign new_n978 = new_n315_1 & new_n977;
  assign new_n979 = ~new_n315_1 & ~new_n977;
  assign new_n980 = ~new_n978 & ~new_n979;
  assign new_n981 = new_n321_1 & new_n333;
  assign new_n982 = ~new_n321_1 & ~new_n333;
  assign new_n983 = ~new_n981 & ~new_n982;
  assign new_n984_1 = new_n980 & ~new_n983;
  assign new_n985 = ~new_n980 & new_n983;
  assign new_n986 = ~new_n984_1 & ~new_n985;
  assign new_n987 = new_n976 & ~new_n986;
  assign new_n988 = ~new_n976 & new_n986;
  assign new_n989 = ~new_n987 & ~new_n988;
  assign new_n990 = ~new_n972 & new_n989;
  assign new_n991 = new_n972 & ~new_n989;
  assign new_n992 = ~n1175 & ~new_n991;
  assign new_n993 = ~new_n990 & new_n992;
  assign new_n994 = ~new_n332 & ~new_n338;
  assign new_n995 = ~new_n331 & new_n338;
  assign new_n996 = ~new_n994 & ~new_n995;
  assign new_n997 = ~new_n315_1 & new_n327;
  assign new_n998 = new_n315_1 & ~new_n327;
  assign new_n999_1 = ~new_n997 & ~new_n998;
  assign new_n1000 = new_n996 & new_n999_1;
  assign new_n1001 = ~new_n996 & ~new_n999_1;
  assign new_n1002 = ~new_n1000 & ~new_n1001;
  assign new_n1003 = new_n522 & ~new_n1002;
  assign new_n1004 = ~new_n522 & new_n1002;
  assign new_n1005 = ~new_n1003 & ~new_n1004;
  assign new_n1006 = ~new_n969 & new_n983;
  assign new_n1007 = ~new_n342_1 & ~new_n983;
  assign new_n1008 = new_n969 & new_n1007;
  assign new_n1009 = ~new_n1006 & ~new_n1008;
  assign new_n1010 = ~new_n1005 & new_n1009;
  assign new_n1011 = new_n1005 & ~new_n1009;
  assign new_n1012 = n1175 & ~new_n1011;
  assign new_n1013 = ~new_n1010 & new_n1012;
  assign new_n1014 = ~new_n993 & ~new_n1013;
  assign new_n1015 = new_n308 & ~new_n580;
  assign new_n1016_1 = ~new_n722_1 & ~new_n1015;
  assign new_n1017 = new_n568 & new_n574_1;
  assign new_n1018 = ~new_n568 & ~new_n574_1;
  assign new_n1019 = ~new_n1017 & ~new_n1018;
  assign new_n1020 = ~new_n573 & new_n584;
  assign new_n1021 = ~new_n585 & ~new_n1020;
  assign new_n1022 = ~new_n1019 & new_n1021;
  assign new_n1023 = new_n1019 & ~new_n1021;
  assign new_n1024 = ~new_n1022 & ~new_n1023;
  assign new_n1025 = new_n1016_1 & new_n1024;
  assign new_n1026 = ~new_n1016_1 & ~new_n1024;
  assign new_n1027_1 = ~new_n1025 & ~new_n1026;
  assign new_n1028 = ~new_n351 & new_n1027_1;
  assign new_n1029 = ~new_n343 & new_n1028;
  assign new_n1030 = ~new_n307_1 & ~new_n580;
  assign new_n1031 = ~new_n583 & ~new_n1030;
  assign new_n1032 = ~new_n1019 & new_n1031;
  assign new_n1033_1 = new_n1019 & ~new_n1031;
  assign new_n1034 = ~new_n1032 & ~new_n1033_1;
  assign new_n1035 = ~new_n723 & new_n1034;
  assign new_n1036 = new_n723 & ~new_n1034;
  assign new_n1037 = ~new_n1035 & ~new_n1036;
  assign new_n1038 = new_n587 & new_n1037;
  assign new_n1039_1 = ~new_n587 & ~new_n1037;
  assign new_n1040 = ~new_n1038 & ~new_n1039_1;
  assign new_n1041 = new_n351 & new_n1040;
  assign new_n1042 = ~n1175 & ~new_n1041;
  assign new_n1043_1 = ~new_n1028 & new_n1042;
  assign new_n1044_1 = ~new_n352 & new_n1040;
  assign new_n1045 = n1175 & ~new_n1044_1;
  assign new_n1046 = ~new_n1043_1 & ~new_n1045;
  assign new_n1047_1 = ~new_n1029 & ~new_n1046;
  assign new_n1048 = new_n1014 & ~new_n1047_1;
  assign new_n1049 = ~new_n1014 & new_n1047_1;
  assign new_n1050_1 = n579 & ~new_n1049;
  assign new_n1051 = ~new_n1048 & new_n1050_1;
  assign new_n1052 = ~n617 & ~n1227;
  assign new_n1053 = ~n591 & n617;
  assign new_n1054 = n39 & ~new_n1053;
  assign new_n1055 = ~new_n1052 & new_n1054;
  assign new_n1056 = n617 & n807;
  assign new_n1057 = ~n617 & n714;
  assign new_n1058_1 = ~new_n1056 & ~new_n1057;
  assign new_n1059 = ~n39 & new_n1058_1;
  assign new_n1060 = ~new_n1055 & ~new_n1059;
  assign new_n1061 = ~n1227 & ~n1498;
  assign new_n1062 = ~n591 & n1498;
  assign new_n1063 = n1039 & ~new_n1062;
  assign new_n1064 = ~new_n1061 & new_n1063;
  assign new_n1065_1 = n807 & n1498;
  assign new_n1066 = n714 & ~n1498;
  assign new_n1067 = ~new_n1065_1 & ~new_n1066;
  assign new_n1068 = ~n1039 & new_n1067;
  assign new_n1069 = ~new_n1064 & ~new_n1068;
  assign new_n1070 = ~n319 & ~n1227;
  assign new_n1071 = n319 & ~n591;
  assign new_n1072 = n1402 & ~new_n1071;
  assign new_n1073 = ~new_n1070 & new_n1072;
  assign new_n1074 = n319 & n807;
  assign new_n1075 = ~n319 & n714;
  assign new_n1076 = ~new_n1074 & ~new_n1075;
  assign new_n1077 = ~n1402 & new_n1076;
  assign new_n1078 = ~new_n1073 & ~new_n1077;
  assign new_n1079 = new_n1069 & new_n1078;
  assign new_n1080 = ~new_n1069 & ~new_n1078;
  assign new_n1081 = ~new_n1079 & ~new_n1080;
  assign new_n1082 = new_n1060 & ~new_n1081;
  assign new_n1083 = ~new_n1060 & new_n1081;
  assign new_n1084 = ~new_n1082 & ~new_n1083;
  assign new_n1085 = ~n1172 & ~n1227;
  assign new_n1086 = ~n591 & n1172;
  assign new_n1087_1 = n697 & ~new_n1086;
  assign new_n1088_1 = ~new_n1085 & new_n1087_1;
  assign new_n1089 = n807 & n1172;
  assign new_n1090 = n714 & ~n1172;
  assign new_n1091 = ~new_n1089 & ~new_n1090;
  assign new_n1092 = ~n697 & new_n1091;
  assign new_n1093 = ~new_n1088_1 & ~new_n1092;
  assign new_n1094 = ~n1227 & ~n1660;
  assign new_n1095_1 = ~n591 & n1660;
  assign new_n1096_1 = n1575 & ~new_n1095_1;
  assign new_n1097_1 = ~new_n1094 & new_n1096_1;
  assign new_n1098 = n807 & n1660;
  assign new_n1099 = n714 & ~n1660;
  assign new_n1100_1 = ~new_n1098 & ~new_n1099;
  assign new_n1101 = ~n1575 & new_n1100_1;
  assign new_n1102 = ~new_n1097_1 & ~new_n1101;
  assign new_n1103 = ~new_n1093 & new_n1102;
  assign new_n1104 = new_n1093 & ~new_n1102;
  assign new_n1105 = ~new_n1103 & ~new_n1104;
  assign new_n1106 = ~n1227 & ~n1553;
  assign new_n1107 = ~n591 & n1553;
  assign new_n1108 = n1755 & ~new_n1107;
  assign new_n1109 = ~new_n1106 & new_n1108;
  assign new_n1110_1 = n807 & n1553;
  assign new_n1111 = n714 & ~n1553;
  assign new_n1112 = ~new_n1110_1 & ~new_n1111;
  assign new_n1113 = ~n1755 & new_n1112;
  assign new_n1114 = ~new_n1109 & ~new_n1113;
  assign new_n1115 = new_n602 & new_n1114;
  assign new_n1116 = ~new_n602 & ~new_n1114;
  assign new_n1117 = ~new_n1115 & ~new_n1116;
  assign new_n1118 = new_n1105 & new_n1117;
  assign new_n1119_1 = ~new_n1105 & ~new_n1117;
  assign new_n1120 = ~new_n1118 & ~new_n1119_1;
  assign new_n1121 = ~n1227 & ~n1729;
  assign new_n1122 = ~n591 & n1729;
  assign new_n1123 = n1135 & ~new_n1122;
  assign new_n1124 = ~new_n1121 & new_n1123;
  assign new_n1125_1 = n807 & n1729;
  assign new_n1126 = n714 & ~n1729;
  assign new_n1127 = ~new_n1125_1 & ~new_n1126;
  assign new_n1128 = ~n1135 & new_n1127;
  assign new_n1129 = ~new_n1124 & ~new_n1128;
  assign new_n1130 = ~n1227 & ~n1238;
  assign new_n1131 = ~n591 & n1238;
  assign new_n1132 = n1100 & ~new_n1131;
  assign new_n1133 = ~new_n1130 & new_n1132;
  assign new_n1134 = n807 & n1238;
  assign new_n1135_1 = n714 & ~n1238;
  assign new_n1136 = ~new_n1134 & ~new_n1135_1;
  assign new_n1137 = ~n1100 & new_n1136;
  assign new_n1138 = ~new_n1133 & ~new_n1137;
  assign new_n1139 = ~new_n1129 & new_n1138;
  assign new_n1140_1 = new_n1129 & ~new_n1138;
  assign new_n1141 = ~new_n1139 & ~new_n1140_1;
  assign new_n1142 = ~new_n1120 & new_n1141;
  assign new_n1143 = new_n1120 & ~new_n1141;
  assign new_n1144 = ~new_n1142 & ~new_n1143;
  assign new_n1145 = new_n1084 & ~new_n1144;
  assign new_n1146 = ~new_n1084 & new_n1144;
  assign new_n1147 = ~n261 & ~new_n1146;
  assign new_n1148 = ~new_n1145 & new_n1147;
  assign new_n1149 = ~new_n303 & ~new_n1148;
  assign new_n1150_1 = ~new_n1051 & ~new_n1149;
  assign new_n1151 = ~n132 & new_n370_1;
  assign n361 = ~new_n1150_1 & ~new_n1151;
  assign new_n1153 = n371 & ~n1281;
  assign new_n1154 = n636 & n1281;
  assign new_n1155 = ~n117 & ~new_n1154;
  assign new_n1156 = ~new_n1153 & new_n1155;
  assign n379 = n1613 & ~new_n1156;
  assign new_n1158 = ~new_n331 & ~new_n448_1;
  assign new_n1159 = ~new_n327 & new_n1158;
  assign new_n1160 = new_n327 & ~new_n1158;
  assign new_n1161 = ~new_n1159 & ~new_n1160;
  assign new_n1162 = new_n303 & new_n1161;
  assign new_n1163_1 = new_n359 & new_n658;
  assign new_n1164 = n9 & new_n370_1;
  assign new_n1165 = ~new_n1163_1 & ~new_n1164;
  assign n1110 = ~new_n1162 & new_n1165;
  assign new_n1167 = new_n302 & ~n1110;
  assign new_n1168 = new_n303 & new_n704;
  assign new_n1169 = n1288 & n1435;
  assign new_n1170 = n721 & ~n1435;
  assign new_n1171 = n1016 & ~new_n1170;
  assign new_n1172_1 = ~new_n1169 & new_n1171;
  assign new_n1173 = ~n1435 & ~n1519;
  assign new_n1174 = ~n77 & n1435;
  assign new_n1175_1 = ~new_n1173 & ~new_n1174;
  assign new_n1176 = ~n1016 & new_n1175_1;
  assign new_n1177_1 = ~new_n1172_1 & ~new_n1176;
  assign new_n1178 = new_n359 & new_n1177_1;
  assign new_n1179 = n1740 & new_n370_1;
  assign new_n1180_1 = ~new_n1178 & ~new_n1179;
  assign n1314 = ~new_n1168 & new_n1180_1;
  assign new_n1182_1 = new_n379_1 & ~n1314;
  assign new_n1183 = n564 & new_n375_1;
  assign new_n1184 = n1655 & new_n377_1;
  assign new_n1185 = ~new_n1183 & ~new_n1184;
  assign new_n1186_1 = ~new_n1182_1 & new_n1185;
  assign n381 = new_n1167 | ~new_n1186_1;
  assign new_n1188 = ~n307 & n377;
  assign new_n1189 = ~n456 & new_n1188;
  assign new_n1190 = n307 & ~n377;
  assign new_n1191 = n488 & new_n1190;
  assign new_n1192 = n307 & n377;
  assign new_n1193 = n1150 & new_n1192;
  assign new_n1194 = ~n307 & ~n377;
  assign new_n1195 = ~n882 & new_n1194;
  assign new_n1196 = ~new_n1193 & ~new_n1195;
  assign new_n1197 = ~new_n1191 & new_n1196;
  assign n413 = new_n1189 | ~new_n1197;
  assign new_n1199 = ~n123 & new_n1188;
  assign new_n1200 = n1177 & new_n1190;
  assign new_n1201 = n754 & new_n1192;
  assign new_n1202 = ~n1027 & new_n1194;
  assign new_n1203 = ~new_n1201 & ~new_n1202;
  assign new_n1204 = ~new_n1200 & new_n1203;
  assign n417 = new_n1199 | ~new_n1204;
  assign new_n1206 = n1181 & ~n1281;
  assign new_n1207_1 = n12 & n1281;
  assign new_n1208 = ~n117 & ~new_n1207_1;
  assign new_n1209 = ~new_n1206 & new_n1208;
  assign n476 = n1613 & ~new_n1209;
  assign new_n1211 = ~n487 & new_n691;
  assign new_n1212 = ~n1710 & new_n689;
  assign new_n1213 = n1362 & new_n693;
  assign new_n1214 = n1598 & new_n695;
  assign new_n1215 = ~new_n1213 & ~new_n1214;
  assign new_n1216 = ~new_n1212 & new_n1215;
  assign new_n1217 = ~new_n1211 & new_n1216;
  assign n567 = n1534 & ~new_n1217;
  assign n574 = ~n1454 | n117;
  assign new_n1220 = new_n302 & ~n456;
  assign new_n1221 = n488 & new_n377_1;
  assign new_n1222 = n1150 & new_n375_1;
  assign new_n1223 = new_n379_1 & ~n882;
  assign new_n1224_1 = ~new_n1222 & ~new_n1223;
  assign new_n1225 = ~new_n1221 & new_n1224_1;
  assign n596 = new_n1220 | ~new_n1225;
  assign new_n1227_1 = ~n257 & ~n1281;
  assign new_n1228 = n1281 & ~n1363;
  assign new_n1229 = ~n117 & ~new_n1228;
  assign n623 = new_n1227_1 | ~new_n1229;
  assign new_n1231 = n261 & n520;
  assign new_n1232 = ~new_n1150_1 & ~new_n1231;
  assign new_n1233_1 = new_n1188 & ~new_n1232;
  assign new_n1234 = n261 & n321;
  assign new_n1235 = new_n384_1 & ~new_n499;
  assign new_n1236 = ~new_n384_1 & ~new_n503;
  assign new_n1237 = ~new_n1235 & ~new_n1236;
  assign new_n1238_1 = ~new_n615 & new_n1237;
  assign new_n1239 = new_n615 & ~new_n1237;
  assign new_n1240 = ~new_n1238_1 & ~new_n1239;
  assign new_n1241 = new_n500 & new_n509;
  assign new_n1242 = new_n501 & ~new_n511;
  assign new_n1243 = ~new_n1241 & ~new_n1242;
  assign new_n1244 = ~new_n1240 & ~new_n1243;
  assign new_n1245 = new_n1240 & new_n1243;
  assign new_n1246 = ~new_n1244 & ~new_n1245;
  assign new_n1247 = ~new_n422 & new_n1246;
  assign new_n1248 = ~new_n414 & new_n1247;
  assign new_n1249 = ~new_n383 & ~new_n501;
  assign new_n1250 = ~new_n502 & ~new_n1249;
  assign new_n1251 = ~new_n615 & new_n1250;
  assign new_n1252 = new_n615 & ~new_n1250;
  assign new_n1253 = ~new_n1251 & ~new_n1252;
  assign new_n1254 = new_n503 & ~new_n509;
  assign new_n1255 = ~new_n504_1 & new_n1254;
  assign new_n1256 = new_n1253 & new_n1255;
  assign new_n1257 = ~new_n1253 & ~new_n1255;
  assign new_n1258 = ~new_n1256 & ~new_n1257;
  assign new_n1259 = new_n414 & ~new_n1258;
  assign new_n1260 = n1366 & ~new_n1259;
  assign new_n1261 = new_n422 & ~new_n1258;
  assign new_n1262 = new_n1260 & ~new_n1261;
  assign new_n1263 = ~new_n1248 & new_n1262;
  assign new_n1264 = ~new_n1247 & ~new_n1261;
  assign new_n1265 = ~n1366 & new_n1264;
  assign new_n1266 = ~new_n1263 & ~new_n1265;
  assign new_n1267 = ~new_n401 & new_n416;
  assign new_n1268 = ~new_n417_1 & ~new_n1267;
  assign new_n1269_1 = ~new_n389_1 & ~new_n395;
  assign new_n1270_1 = ~new_n396 & ~new_n1269_1;
  assign new_n1271 = new_n402 & new_n471;
  assign new_n1272 = ~new_n402 & ~new_n471;
  assign new_n1273 = ~new_n1271 & ~new_n1272;
  assign new_n1274 = new_n1270_1 & ~new_n1273;
  assign new_n1275 = ~new_n1270_1 & new_n1273;
  assign new_n1276 = ~new_n1274 & ~new_n1275;
  assign new_n1277 = ~new_n1268 & new_n1276;
  assign new_n1278 = new_n1268 & ~new_n1276;
  assign new_n1279_1 = ~new_n1277 & ~new_n1278;
  assign new_n1280 = new_n420 & new_n1279_1;
  assign new_n1281_1 = ~new_n420 & ~new_n1279_1;
  assign new_n1282 = ~n1366 & ~new_n1281_1;
  assign new_n1283 = ~new_n1280 & new_n1282;
  assign new_n1284 = ~new_n413_1 & ~new_n418;
  assign new_n1285 = ~new_n387_1 & new_n1284;
  assign new_n1286 = ~new_n388 & ~new_n1284;
  assign new_n1287 = ~new_n1285 & ~new_n1286;
  assign new_n1288_1 = ~new_n410 & ~new_n471;
  assign new_n1289 = ~new_n412 & ~new_n1288_1;
  assign new_n1290 = ~new_n402 & new_n406;
  assign new_n1291 = new_n402 & ~new_n406;
  assign new_n1292 = ~new_n1290 & ~new_n1291;
  assign new_n1293 = new_n1270_1 & ~new_n1292;
  assign new_n1294 = ~new_n1270_1 & new_n1292;
  assign new_n1295 = ~new_n1293 & ~new_n1294;
  assign new_n1296 = new_n1289 & new_n1295;
  assign new_n1297_1 = ~new_n1289 & ~new_n1295;
  assign new_n1298 = ~new_n1296 & ~new_n1297_1;
  assign new_n1299_1 = new_n1287 & new_n1298;
  assign new_n1300 = ~new_n1287 & ~new_n1298;
  assign new_n1301 = ~new_n1299_1 & ~new_n1300;
  assign new_n1302 = n1366 & new_n1301;
  assign new_n1303 = ~new_n1283 & ~new_n1302;
  assign new_n1304 = ~new_n1266 & new_n1303;
  assign new_n1305 = new_n1266 & ~new_n1303;
  assign new_n1306 = n579 & ~new_n1305;
  assign new_n1307 = ~new_n1304 & new_n1306;
  assign new_n1308 = ~n1227 & ~n1435;
  assign new_n1309 = ~n591 & n1435;
  assign new_n1310 = n1016 & ~new_n1309;
  assign new_n1311 = ~new_n1308 & new_n1310;
  assign new_n1312 = n807 & n1435;
  assign new_n1313 = n714 & ~n1435;
  assign new_n1314_1 = ~new_n1312 & ~new_n1313;
  assign new_n1315 = ~n1016 & new_n1314_1;
  assign new_n1316 = ~new_n1311 & ~new_n1315;
  assign new_n1317 = n238 & n591;
  assign new_n1318 = ~n238 & ~n807;
  assign new_n1319 = ~new_n1317 & ~new_n1318;
  assign new_n1320 = ~new_n800 & new_n1319;
  assign new_n1321 = new_n800 & ~new_n1319;
  assign new_n1322_1 = ~new_n1320 & ~new_n1321;
  assign new_n1323 = ~new_n1316 & new_n1322_1;
  assign new_n1324 = new_n1316 & ~new_n1322_1;
  assign new_n1325 = ~new_n1323 & ~new_n1324;
  assign new_n1326 = ~n380 & ~n1227;
  assign new_n1327 = n380 & ~n591;
  assign new_n1328 = n1391 & ~new_n1327;
  assign new_n1329 = ~new_n1326 & new_n1328;
  assign new_n1330 = n380 & n807;
  assign new_n1331 = ~n380 & n714;
  assign new_n1332 = ~new_n1330 & ~new_n1331;
  assign new_n1333 = ~n1391 & new_n1332;
  assign new_n1334 = ~new_n1329 & ~new_n1333;
  assign new_n1335 = ~n1043 & ~n1227;
  assign new_n1336 = ~n591 & n1043;
  assign new_n1337 = n1125 & ~new_n1336;
  assign new_n1338_1 = ~new_n1335 & new_n1337;
  assign new_n1339 = n807 & n1043;
  assign new_n1340 = n714 & ~n1043;
  assign new_n1341 = ~new_n1339 & ~new_n1340;
  assign new_n1342 = ~n1125 & new_n1341;
  assign new_n1343 = ~new_n1338_1 & ~new_n1342;
  assign new_n1344 = new_n1334 & new_n1343;
  assign new_n1345 = ~new_n1334 & ~new_n1343;
  assign new_n1346_1 = ~new_n1344 & ~new_n1345;
  assign new_n1347 = ~new_n1325 & new_n1346_1;
  assign new_n1348 = new_n1325 & ~new_n1346_1;
  assign new_n1349 = ~new_n1347 & ~new_n1348;
  assign new_n1350 = ~new_n623_1 & new_n947;
  assign new_n1351 = new_n623_1 & ~new_n947;
  assign new_n1352 = ~new_n1350 & ~new_n1351;
  assign new_n1353_1 = new_n436 & new_n517;
  assign new_n1354 = ~new_n436 & ~new_n517;
  assign new_n1355_1 = ~new_n1353_1 & ~new_n1354;
  assign new_n1356 = new_n1352 & new_n1355_1;
  assign new_n1357_1 = ~new_n1352 & ~new_n1355_1;
  assign new_n1358 = ~new_n1356 & ~new_n1357_1;
  assign new_n1359 = ~new_n1349 & new_n1358;
  assign new_n1360 = new_n1349 & ~new_n1358;
  assign new_n1361_1 = ~new_n1359 & ~new_n1360;
  assign new_n1362_1 = ~n579 & new_n1361_1;
  assign new_n1363_1 = ~n261 & ~new_n1362_1;
  assign new_n1364 = ~new_n1307 & new_n1363_1;
  assign new_n1365 = ~new_n1234 & ~new_n1364;
  assign new_n1366_1 = new_n1194 & ~new_n1365;
  assign new_n1367 = n1756 & new_n1190;
  assign new_n1368 = n187 & new_n1192;
  assign new_n1369 = ~new_n1367 & ~new_n1368;
  assign new_n1370_1 = ~new_n1366_1 & new_n1369;
  assign n635 = new_n1233_1 | ~new_n1370_1;
  assign new_n1372 = ~n1281 & n1299;
  assign new_n1373 = n403 & n1281;
  assign new_n1374 = ~n117 & ~new_n1373;
  assign new_n1375 = ~new_n1372 & new_n1374;
  assign n649 = n1613 & ~new_n1375;
  assign new_n1377_1 = new_n302 & ~new_n1232;
  assign new_n1378_1 = new_n379_1 & ~new_n1365;
  assign new_n1379 = n187 & new_n375_1;
  assign new_n1380 = n1756 & new_n377_1;
  assign new_n1381 = ~new_n1379 & ~new_n1380;
  assign new_n1382 = ~new_n1378_1 & new_n1381;
  assign n661 = new_n1377_1 | ~new_n1382;
  assign new_n1384 = new_n581 & new_n1017;
  assign n673 = new_n343 & new_n1384;
  assign new_n1386 = ~n1087 & new_n1188;
  assign new_n1387 = n297 & new_n1192;
  assign new_n1388 = n384 & new_n1190;
  assign new_n1389 = ~n75 & new_n1194;
  assign new_n1390_1 = ~new_n1388 & ~new_n1389;
  assign new_n1391_1 = ~new_n1387 & new_n1390_1;
  assign n722 = new_n1386 | ~new_n1391_1;
  assign new_n1393 = ~n964 & new_n470;
  assign new_n1394 = ~n370 & new_n445;
  assign new_n1395 = n715 & new_n468;
  assign new_n1396_1 = n128 & new_n466;
  assign new_n1397 = ~new_n1395 & ~new_n1396_1;
  assign new_n1398 = ~new_n1394 & new_n1397;
  assign new_n1399 = ~new_n1393 & new_n1398;
  assign n786 = n1534 & ~new_n1399;
  assign new_n1401 = ~n1110 & new_n1188;
  assign new_n1402_1 = ~n1314 & new_n1194;
  assign new_n1403 = n564 & new_n1192;
  assign new_n1404 = n1655 & new_n1190;
  assign new_n1405 = ~new_n1403 & ~new_n1404;
  assign new_n1406_1 = ~new_n1402_1 & new_n1405;
  assign n824 = new_n1401 | ~new_n1406_1;
  assign new_n1408_1 = ~n1346 & new_n1188;
  assign new_n1409_1 = ~n168 & new_n1194;
  assign new_n1410 = n760 & new_n1190;
  assign new_n1411 = n179 & new_n1192;
  assign new_n1412 = ~new_n1410 & ~new_n1411;
  assign new_n1413 = ~new_n1409_1 & new_n1412;
  assign n840 = new_n1408_1 | ~new_n1413;
  assign new_n1415 = ~n1790 & ~new_n512;
  assign new_n1416 = n1790 & new_n512;
  assign n889 = new_n1415 | new_n1416;
  assign new_n1418 = ~n75 & new_n691;
  assign new_n1419 = new_n689 & ~n1087;
  assign new_n1420 = n1353 & new_n693;
  assign new_n1421 = n530 & new_n695;
  assign new_n1422 = ~new_n1420 & ~new_n1421;
  assign new_n1423 = ~new_n1419 & new_n1422;
  assign new_n1424 = ~new_n1418 & new_n1423;
  assign n944 = n1534 & ~new_n1424;
  assign new_n1426_1 = ~n1281 & ~n1700;
  assign new_n1427_1 = ~n38 & n1281;
  assign new_n1428 = ~n117 & ~new_n1427_1;
  assign n951 = new_n1426_1 | ~new_n1428;
  assign new_n1430 = ~n33 & new_n370_1;
  assign n974 = ~new_n1364 & ~new_n1430;
  assign new_n1432 = n1180 & new_n695;
  assign new_n1433 = ~n1346 & new_n689;
  assign new_n1434 = n7 & new_n693;
  assign new_n1435_1 = ~n168 & new_n691;
  assign new_n1436_1 = ~new_n1434 & ~new_n1435_1;
  assign new_n1437 = ~new_n1433 & new_n1436_1;
  assign new_n1438 = ~new_n1432 & new_n1437;
  assign n1050 = n1534 & ~new_n1438;
  assign new_n1440 = n1663 & new_n466;
  assign new_n1441 = new_n445 & ~new_n1232;
  assign new_n1442 = n962 & new_n468;
  assign new_n1443 = new_n470 & ~new_n1365;
  assign new_n1444 = ~new_n1442 & ~new_n1443;
  assign new_n1445 = ~new_n1441 & new_n1444;
  assign new_n1446 = ~new_n1440 & new_n1445;
  assign n1065 = ~n1534 | new_n1446;
  assign new_n1448 = ~n1710 & new_n1188;
  assign new_n1449 = n1540 & new_n1190;
  assign new_n1450 = n565 & new_n1192;
  assign new_n1451 = ~n487 & new_n1194;
  assign new_n1452 = ~new_n1450 & ~new_n1451;
  assign new_n1453 = ~new_n1449 & new_n1452;
  assign n1096 = new_n1448 | ~new_n1453;
  assign n1163 = ~n1463 | n117;
  assign new_n1456 = new_n689 & ~n456;
  assign new_n1457 = new_n691 & ~n882;
  assign new_n1458 = n270 & new_n695;
  assign new_n1459 = n335 & new_n693;
  assign new_n1460 = ~new_n1458 & ~new_n1459;
  assign new_n1461 = ~new_n1457 & new_n1460;
  assign new_n1462_1 = ~new_n1456 & new_n1461;
  assign n1186 = n1534 & ~new_n1462_1;
  assign new_n1464_1 = ~new_n788 & ~new_n931;
  assign new_n1465 = ~new_n357_1 & new_n728;
  assign new_n1466 = new_n1464_1 & new_n1465;
  assign new_n1467 = ~new_n450 & ~new_n527;
  assign new_n1468 = ~new_n759 & new_n1467;
  assign new_n1469 = new_n592 & ~new_n1161;
  assign new_n1470 = new_n1468 & new_n1469;
  assign n1224 = new_n1466 & new_n1470;
  assign new_n1472 = n1357 & n1649;
  assign new_n1473 = n1790 & new_n612;
  assign new_n1474 = ~n1790 & ~new_n612;
  assign new_n1475 = ~new_n1473 & ~new_n1474;
  assign new_n1476 = ~n342 & new_n1475;
  assign new_n1477 = n342 & ~n1793;
  assign new_n1478 = n495 & ~new_n1477;
  assign new_n1479 = ~new_n1476 & new_n1478;
  assign new_n1480 = ~n342 & ~new_n623_1;
  assign new_n1481 = n342 & n482;
  assign new_n1482 = ~n495 & ~new_n1481;
  assign new_n1483 = ~new_n1480 & new_n1482;
  assign new_n1484 = ~new_n1479 & ~new_n1483;
  assign n1269 = ~new_n1472 & new_n1484;
  assign new_n1486 = new_n445 & ~n1110;
  assign new_n1487 = n387 & new_n466;
  assign new_n1488 = n606 & new_n468;
  assign new_n1489 = new_n470 & ~n1314;
  assign new_n1490 = ~new_n1488 & ~new_n1489;
  assign new_n1491_1 = ~new_n1487 & new_n1490;
  assign new_n1492 = ~new_n1486 & new_n1491_1;
  assign n1270 = n1534 & ~new_n1492;
  assign new_n1494 = new_n302 & ~n259;
  assign new_n1495_1 = new_n379_1 & ~n454;
  assign new_n1496 = n676 & new_n375_1;
  assign new_n1497 = n1207 & new_n377_1;
  assign new_n1498_1 = ~new_n1496 & ~new_n1497;
  assign new_n1499 = ~new_n1495_1 & new_n1498_1;
  assign n1297 = new_n1494 | ~new_n1499;
  assign new_n1501 = new_n689 & ~new_n1232;
  assign new_n1502 = n962 & new_n693;
  assign new_n1503_1 = n1663 & new_n695;
  assign new_n1504 = new_n691 & ~new_n1365;
  assign new_n1505 = ~new_n1503_1 & ~new_n1504;
  assign new_n1506 = ~new_n1502 & new_n1505;
  assign new_n1507 = ~new_n1501 & new_n1506;
  assign n1322 = ~n1534 | new_n1507;
  assign new_n1509 = ~n1631 & new_n1188;
  assign new_n1510_1 = n239 & new_n1190;
  assign new_n1511_1 = n1119 & new_n1192;
  assign new_n1512 = ~n1495 & new_n1194;
  assign new_n1513 = ~new_n1511_1 & ~new_n1512;
  assign new_n1514 = ~new_n1510_1 & new_n1513;
  assign n1377 = new_n1509 | ~new_n1514;
  assign new_n1516 = ~n259 & new_n1188;
  assign new_n1517 = ~n454 & new_n1194;
  assign new_n1518_1 = n676 & new_n1192;
  assign new_n1519_1 = n1207 & new_n1190;
  assign new_n1520 = ~new_n1518_1 & ~new_n1519_1;
  assign new_n1521 = ~new_n1517 & new_n1520;
  assign n1390 = new_n1516 | ~new_n1521;
  assign n1409 = ~n841 | n1427;
  assign new_n1524 = new_n351 & new_n582;
  assign new_n1525 = new_n586 & ~new_n1524;
  assign new_n1526 = ~new_n566_1 & new_n1525;
  assign n1414 = ~new_n567_1 & ~new_n1526;
  assign new_n1528 = new_n470 & ~n1027;
  assign new_n1529 = new_n445 & ~n123;
  assign new_n1530 = n1033 & new_n466;
  assign new_n1531 = n830 & new_n468;
  assign new_n1532 = ~new_n1530 & ~new_n1531;
  assign new_n1533 = ~new_n1529 & new_n1532;
  assign new_n1534_1 = ~new_n1528 & new_n1533;
  assign n1462 = n1534 & ~new_n1534_1;
  assign new_n1536 = new_n302 & ~n1631;
  assign new_n1537 = n239 & new_n377_1;
  assign new_n1538 = n1119 & new_n375_1;
  assign new_n1539 = new_n379_1 & ~n1495;
  assign new_n1540_1 = ~new_n1538 & ~new_n1539;
  assign new_n1541 = ~new_n1537 & new_n1540_1;
  assign n1510 = new_n1536 | ~new_n1541;
  assign new_n1543_1 = ~n370 & new_n1188;
  assign new_n1544 = n19 & new_n1192;
  assign new_n1545 = n955 & new_n1190;
  assign new_n1546 = ~n964 & new_n1194;
  assign new_n1547 = ~new_n1545 & ~new_n1546;
  assign new_n1548 = ~new_n1544 & new_n1547;
  assign n1543 = new_n1543_1 | ~new_n1548;
  assign n1584 = n912 & n1613;
  assign new_n1551 = new_n470 & ~n75;
  assign new_n1552 = new_n445 & ~n1087;
  assign new_n1553_1 = n1353 & new_n468;
  assign new_n1554 = n530 & new_n466;
  assign new_n1555 = ~new_n1553_1 & ~new_n1554;
  assign new_n1556 = ~new_n1552 & new_n1555;
  assign new_n1557 = ~new_n1551 & new_n1556;
  assign n1587 = n1534 & ~new_n1557;
  assign new_n1559 = new_n554 & ~new_n800;
  assign new_n1560 = new_n1351 & new_n1559;
  assign new_n1561 = ~new_n486 & ~new_n775;
  assign new_n1562 = ~new_n1177_1 & new_n1561;
  assign new_n1563 = new_n1354 & new_n1562;
  assign n1708 = new_n1560 & new_n1563;
  assign new_n1565 = new_n689 & ~n1110;
  assign new_n1566 = n606 & new_n693;
  assign new_n1567 = n387 & new_n695;
  assign new_n1568_1 = new_n691 & ~n1314;
  assign new_n1569 = ~new_n1567 & ~new_n1568_1;
  assign new_n1570 = ~new_n1566 & new_n1569;
  assign new_n1571 = ~new_n1565 & new_n1570;
  assign n1733 = n1534 & ~new_n1571;
  assign new_n1573 = new_n302 & ~n1346;
  assign new_n1574 = new_n379_1 & ~n168;
  assign new_n1575_1 = n760 & new_n377_1;
  assign new_n1576 = n179 & new_n375_1;
  assign new_n1577 = ~new_n1575_1 & ~new_n1576;
  assign new_n1578 = ~new_n1574 & new_n1577;
  assign n1761 = new_n1573 | ~new_n1578;
  assign n1780 = n84 & n1058;
  assign new_n1581 = new_n470 & ~n1495;
  assign new_n1582 = new_n445 & ~n1631;
  assign new_n1583 = n236 & new_n468;
  assign new_n1584_1 = n1743 & new_n466;
  assign new_n1585 = ~new_n1583 & ~new_n1584_1;
  assign new_n1586 = ~new_n1582 & new_n1585;
  assign new_n1587_1 = ~new_n1581 & new_n1586;
  assign n1784 = n1534 & ~new_n1587_1;
  assign new_n1589 = new_n445 & ~n1710;
  assign new_n1590 = new_n470 & ~n487;
  assign new_n1591 = n1362 & new_n468;
  assign new_n1592 = n1598 & new_n466;
  assign new_n1593 = ~new_n1591 & ~new_n1592;
  assign new_n1594 = ~new_n1590 & new_n1593;
  assign new_n1595 = ~new_n1589 & new_n1594;
  assign n1794 = n1534 & ~new_n1595;
  assign n61 = ~n1503;
  assign n112 = ~n448;
  assign n193 = ~n937;
  assign n357 = ~n566;
  assign n765 = ~n918;
  assign n849 = ~n516;
  assign n1140 = ~n1568;
  assign n1370 = ~n92;
  assign n1464 = ~n389;
  assign n1654 = ~n457;
  assign n1676 = ~n1338;
  assign n66 = n389;
  assign n129 = n566;
  assign n173 = n84;
  assign n375 = n84;
  assign n542 = n84;
  assign n611 = n84;
  assign n776 = n1613;
  assign n793 = n544;
  assign n845 = n1613;
  assign n860 = n623;
  assign n967 = n357;
  assign n1044 = n765;
  assign n1233 = n765;
  assign n1355 = n288;
  assign n1378 = n84;
  assign n1425 = n1534;
  assign n1657 = n389;
  assign n1682 = n130;
  assign n1697 = n1414;
  assign n1698 = n673;
  assign n1721 = n235;
endmodule


