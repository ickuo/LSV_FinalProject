module top( n8 , n46 , n74 , n91 , n126 , n203 , n271 , n278 , n389 , 
n394 , n411 , n427 , n451 , n462 , n490 , n498 , n543 , n650 , n656 , 
n666 , n674 , n682 , n702 , n730 , n737 , n760 , n844 , n884 , n948 , 
n977 , n1027 , n1093 , n1094 , n1122 , n1124 , n1222 , n1265 , n1268 , n1329 , 
n1347 , n1545 , n1568 , n1637 , n1702 , n1739 , n1763 , n1776 , n1827 , n1900 , 
n1927 , n1951 , n2027 , n2048 , n2061 , n2126 , n2164 , n2166 , n2175 , n2201 , 
n2223 , n2311 , n2334 , n2407 , n2454 , n2556 , n2559 , n2572 , n2573 , n2615 , 
n2672 , n2674 , n2699 , n2734 , n2895 , n3090 , n3130 , n3166 , n3242 , n3263 , 
n3340 , n3367 , n3388 , n3506 , n3532 , n3603 , n3652 , n3655 , n3673 , n3775 , 
n3799 , n3804 , n3833 , n3854 , n3893 , n3901 , n3910 , n3972 , n4000 , n4022 , 
n4039 , n4117 , n4125 , n4131 , n4147 , n4154 , n4172 , n4175 , n4225 , n4279 , 
n4282 , n4292 , n4305 , n4345 , n4437 , n4541 , n4604 , n4615 , n4659 , n4672 , 
n4755 , n4774 , n4785 , n4858 , n4895 , n4907 , n4971 , n5009 , n5014 , n5023 , 
n5033 , n5046 , n5077 , n5184 , n5185 , n5225 , n5430 , n5449 , n5467 , n5479 , 
n5502 , n5550 , n5586 , n5601 , n5725 , n5786 , n5806 , n5851 , n5943 , n5950 , 
n5960 , n5987 , n6007 , n6012 , n6054 , n6114 , n6147 , n6198 , n6251 , n6258 , 
n6270 , n6275 , n6314 , n6362 , n6436 , n6460 , n6480 , n6517 , n6555 , n6586 , 
n6680 , n6682 , n6693 , n6696 , n6703 , n6758 , n6786 , n6791 , n6810 , n6853 , 
n6873 , n6946 , n6952 , n6979 , n6999 , n7071 , n7073 , n7104 , n7132 , n7152 , 
n7246 , n7265 , n7272 , n7282 , n7354 , n7382 , n7450 , n7652 , n7655 , n7667 , 
n7748 , n7771 , n7825 , n7832 , n7941 , n7972 , n7988 , n8002 , n8044 , n8068 , 
n8073 , n8085 , n8124 , n8144 , n8204 , n8215 , n8262 , n8302 , n8306 , n8315 , 
n8397 , n8439 , n8463 , n8471 , n8486 , n8550 , n8552 , n8598 , n8604 , n8635 , 
n8649 , n8737 , n8746 , n8780 , n8799 , n8800 , n8873 , n8892 , n8909 , n8926 , 
n8997 , n9026 , n9096 , n9110 , n9154 , n9186 , n9252 , n9314 , n9342 , n9437 , 
n9447 , n9543 , n9544 , n9555 , n9570 , n9589 , n9665 , n9717 , n9830 , n9893 , 
n9921 , n9936 , n9977 , n10050 , n10051 , n10061 , n10080 , n10112 , n10147 , n10255 , 
n10278 , n10283 , n10378 , n10407 , n10426 , n10446 , n10466 , n10470 , n10515 , n10573 , 
n10591 , n10615 , n10630 , n10736 , n10750 , n10765 , n10791 , n10802 , n10862 , n10912 , 
n10915 , n10945 , n11122 , n11143 , n11158 , n11269 , n11345 , n11393 , n11404 , n11463 , 
n11529 , n11534 , n11590 , n11605 , n11627 , n11664 , n11666 , n11756 , n11776 , n11822 , 
n11842 , n11847 , n11854 , n11875 , n11902 , n11930 , n11933 , n11961 , n12009 , n12012 , 
n12025 , n12032 , n12142 , n12166 , n12218 , n12232 , n12270 , n12321 , n12336 , n12355 , 
n12535 , n12573 , n12614 , n12782 , n12829 , n12885 , n12927 , n12976 , n12989 , n13000 , 
n13010 , n13045 , n13093 , n13102 , n13109 , n13114 , n13141 , n13186 , n13224 , n13231 , 
n13295 , n13316 , n13363 , n13364 , n13509 , n13511 , n13561 , n13577 , n13625 , n13636 , 
n13639 , n13658 , n13693 , n13760 , n13814 , n13853 , n13870 , n13882 , n13890 , n13944 , 
n13953 , n13959 , n13992 , n14072 , n14163 , n14289 , n14293 , n14303 , n14307 , n14330 , 
n14399 , n14408 , n14463 , n14464 , n14475 , n14483 );
    input n74 , n203 , n271 , n394 , n411 , n427 , n462 , n498 , n650 , 
n656 , n666 , n674 , n702 , n730 , n737 , n760 , n844 , n977 , n1027 , 
n1093 , n1222 , n1265 , n1268 , n1347 , n1568 , n1637 , n1702 , n1763 , n1776 , 
n2048 , n2061 , n2164 , n2166 , n2201 , n2334 , n2454 , n2573 , n2615 , n2674 , 
n2699 , n2895 , n3130 , n3166 , n3263 , n3367 , n3388 , n3506 , n3532 , n3652 , 
n3655 , n3673 , n3775 , n3799 , n3804 , n3833 , n3893 , n3910 , n3972 , n4000 , 
n4022 , n4039 , n4117 , n4131 , n4147 , n4154 , n4172 , n4175 , n4225 , n4282 , 
n4292 , n4615 , n4659 , n4755 , n4774 , n4785 , n4895 , n4907 , n5009 , n5014 , 
n5023 , n5033 , n5046 , n5077 , n5184 , n5185 , n5225 , n5430 , n5449 , n5467 , 
n5502 , n5601 , n5725 , n5786 , n5943 , n5950 , n5960 , n6007 , n6054 , n6114 , 
n6147 , n6251 , n6258 , n6270 , n6362 , n6436 , n6460 , n6480 , n6517 , n6555 , 
n6586 , n6680 , n6693 , n6703 , n6758 , n6791 , n6810 , n6873 , n6946 , n6999 , 
n7104 , n7272 , n7282 , n7354 , n7450 , n7652 , n7667 , n7748 , n7832 , n7941 , 
n7972 , n7988 , n8002 , n8044 , n8073 , n8204 , n8262 , n8302 , n8315 , n8397 , 
n8439 , n8463 , n8486 , n8550 , n8552 , n8598 , n8635 , n8649 , n8737 , n8746 , 
n8780 , n8799 , n8800 , n8873 , n8892 , n8926 , n8997 , n9026 , n9110 , n9154 , 
n9186 , n9252 , n9314 , n9543 , n9544 , n9555 , n9589 , n9830 , n9893 , n9921 , 
n9936 , n9977 , n10050 , n10051 , n10061 , n10080 , n10112 , n10147 , n10255 , n10278 , 
n10283 , n10378 , n10407 , n10426 , n10446 , n10466 , n10470 , n10573 , n10615 , n10630 , 
n10736 , n10750 , n10765 , n10862 , n10912 , n10945 , n11143 , n11158 , n11269 , n11345 , 
n11404 , n11529 , n11590 , n11605 , n11666 , n11756 , n11776 , n11842 , n11854 , n11875 , 
n11902 , n11930 , n11933 , n11961 , n12009 , n12012 , n12025 , n12142 , n12218 , n12270 , 
n12321 , n12336 , n12573 , n12614 , n12782 , n12829 , n12885 , n12927 , n12976 , n13000 , 
n13093 , n13102 , n13109 , n13186 , n13224 , n13231 , n13295 , n13363 , n13364 , n13509 , 
n13511 , n13561 , n13625 , n13636 , n13814 , n13882 , n13890 , n13944 , n13992 , n14072 , 
n14163 , n14293 , n14303 , n14408 , n14464 , n14475 , n14483 ;
    output n8 , n46 , n91 , n126 , n278 , n389 , n451 , n490 , n543 , 
n682 , n884 , n948 , n1094 , n1122 , n1124 , n1329 , n1545 , n1739 , n1827 , 
n1900 , n1927 , n1951 , n2027 , n2126 , n2175 , n2223 , n2311 , n2407 , n2556 , 
n2559 , n2572 , n2672 , n2734 , n3090 , n3242 , n3340 , n3603 , n3854 , n3901 , 
n4125 , n4279 , n4305 , n4345 , n4437 , n4541 , n4604 , n4672 , n4858 , n4971 , 
n5479 , n5550 , n5586 , n5806 , n5851 , n5987 , n6012 , n6198 , n6275 , n6314 , 
n6682 , n6696 , n6786 , n6853 , n6952 , n6979 , n7071 , n7073 , n7132 , n7152 , 
n7246 , n7265 , n7382 , n7655 , n7771 , n7825 , n8068 , n8085 , n8124 , n8144 , 
n8215 , n8306 , n8471 , n8604 , n8909 , n9096 , n9342 , n9437 , n9447 , n9570 , 
n9665 , n9717 , n10515 , n10591 , n10791 , n10802 , n10915 , n11122 , n11393 , n11463 , 
n11534 , n11627 , n11664 , n11822 , n11847 , n12032 , n12166 , n12232 , n12355 , n12535 , 
n12989 , n13010 , n13045 , n13114 , n13141 , n13316 , n13577 , n13639 , n13658 , n13693 , 
n13760 , n13853 , n13870 , n13953 , n13959 , n14289 , n14307 , n14330 , n14399 , n14463 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n9 , 
n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
n40 , n41 , n42 , n43 , n44 , n45 , n47 , n48 , n49 , n50 , 
n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
n71 , n72 , n73 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , 
n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n92 , 
n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , 
n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , 
n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , 
n123 , n124 , n125 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , 
n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , 
n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , 
n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , 
n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , 
n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , 
n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , 
n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n204 , 
n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , 
n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , 
n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , 
n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , 
n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , 
n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , 
n265 , n266 , n267 , n268 , n269 , n270 , n272 , n273 , n274 , n275 , 
n276 , n277 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , 
n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , 
n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , 
n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , 
n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , 
n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , 
n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , 
n387 , n388 , n390 , n391 , n392 , n393 , n395 , n396 , n397 , n398 , 
n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , 
n409 , n410 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
n420 , n421 , n422 , n423 , n424 , n425 , n426 , n428 , n429 , n430 , 
n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , 
n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , 
n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , 
n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , 
n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , 
n483 , n484 , n485 , n486 , n487 , n488 , n489 , n491 , n492 , n493 , 
n494 , n495 , n496 , n497 , n499 , n500 , n501 , n502 , n503 , n504 , 
n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , 
n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , 
n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , 
n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n544 , n545 , 
n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , 
n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , 
n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , 
n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , 
n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , 
n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , 
n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , 
n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , 
n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , 
n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , 
n646 , n647 , n648 , n649 , n651 , n652 , n653 , n654 , n655 , n657 , 
n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n667 , n668 , 
n669 , n670 , n671 , n672 , n673 , n675 , n676 , n677 , n678 , n679 , 
n680 , n681 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , 
n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , 
n701 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , 
n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , 
n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n731 , n732 , 
n733 , n734 , n735 , n736 , n738 , n739 , n740 , n741 , n742 , n743 , 
n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , 
n754 , n755 , n756 , n757 , n758 , n759 , n761 , n762 , n763 , n764 , 
n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , 
n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , 
n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , 
n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , 
n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , 
n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , 
n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , 
n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n845 , 
n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , 
n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , 
n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , 
n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n885 , n886 , 
n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , 
n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , 
n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , 
n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , 
n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , 
n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , 
n947 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , 
n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , 
n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n978 , 
n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , 
n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , 
n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , 
n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , 
n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1028 , n1029 , 
n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
n1090 , n1091 , n1092 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , 
n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , 
n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , 
n1123 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , 
n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , 
n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , 
n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , 
n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , 
n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , 
n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , 
n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , 
n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , 
n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1223 , n1224 , 
n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , 
n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , 
n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , 
n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , 
n1266 , n1267 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , 
n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , 
n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , 
n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , 
n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , 
n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , 
n1327 , n1328 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , 
n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1348 , 
n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , 
n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , 
n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , 
n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , 
n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , 
n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , 
n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , 
n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , 
n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , 
n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , 
n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , 
n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , 
n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , 
n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , 
n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , 
n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , 
n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , 
n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , 
n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , 
n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1546 , n1547 , n1548 , n1549 , 
n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1569 , n1570 , 
n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , 
n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , 
n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , 
n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , 
n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , 
n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , 
n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1638 , n1639 , n1640 , n1641 , 
n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , 
n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , 
n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , 
n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , 
n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , 
n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , 
n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , 
n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , 
n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , 
n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1740 , n1741 , n1742 , n1743 , 
n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , 
n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1764 , 
n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , 
n1775 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , 
n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , 
n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , 
n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , 
n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , 
n1826 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , 
n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , 
n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , 
n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , 
n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , 
n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , 
n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , 
n1897 , n1898 , n1899 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , 
n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , 
n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1928 , 
n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , 
n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , 
n1949 , n1950 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2028 , n2029 , n2030 , 
n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , 
n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2049 , n2050 , n2051 , 
n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2062 , 
n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , 
n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , 
n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , 
n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , 
n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , 
n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , 
n2123 , n2124 , n2125 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , 
n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , 
n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , 
n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , 
n2165 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2176 , 
n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , 
n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , 
n2197 , n2198 , n2199 , n2200 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , 
n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , 
n2218 , n2219 , n2220 , n2221 , n2222 , n2224 , n2225 , n2226 , n2227 , n2228 , 
n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , 
n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , 
n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , 
n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , 
n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , 
n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , 
n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , 
n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , 
n2309 , n2310 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
n2330 , n2331 , n2332 , n2333 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , 
n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , 
n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , 
n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , 
n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , 
n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , 
n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2408 , n2409 , n2410 , n2411 , 
n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , 
n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , 
n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , 
n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , 
n2452 , n2453 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , 
n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , 
n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , 
n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , 
n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , 
n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , 
n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , 
n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , 
n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , 
n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , 
n2553 , n2554 , n2555 , n2557 , n2558 , n2560 , n2561 , n2562 , n2563 , n2564 , 
n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2574 , n2575 , n2576 , 
n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , 
n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , 
n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , 
n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2616 , n2617 , 
n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , 
n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , 
n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , 
n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , 
n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , 
n2668 , n2669 , n2670 , n2671 , n2673 , n2675 , n2676 , n2677 , n2678 , n2679 , 
n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2700 , 
n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , 
n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , 
n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , 
n2731 , n2732 , n2733 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , 
n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , 
n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , 
n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , 
n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , 
n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , 
n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , 
n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , 
n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , 
n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , 
n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , 
n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , 
n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , 
n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , 
n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , 
n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , 
n2892 , n2893 , n2894 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , 
n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , 
n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , 
n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , 
n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , 
n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , 
n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , 
n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , 
n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , 
n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , 
n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , 
n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , 
n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , 
n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , 
n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , 
n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , 
n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , 
n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , 
n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , 
n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3091 , n3092 , n3093 , 
n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , 
n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , 
n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , 
n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3131 , n3132 , n3133 , n3134 , 
n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , 
n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , 
n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , 
n3165 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , 
n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , 
n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , 
n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , 
n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , 
n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , 
n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , 
n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3243 , n3244 , n3245 , n3246 , 
n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , 
n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3264 , n3265 , n3266 , n3267 , 
n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , 
n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , 
n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , 
n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , 
n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , 
n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , 
n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , 
n3338 , n3339 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , 
n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , 
n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3368 , n3369 , 
n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3389 , n3390 , 
n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , 
n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , 
n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , 
n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , 
n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , 
n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , 
n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , 
n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , 
n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , 
n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
n3501 , n3502 , n3503 , n3504 , n3505 , n3507 , n3508 , n3509 , n3510 , n3511 , 
n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , 
n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , 
n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , 
n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , 
n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , 
n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , 
n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , 
n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , 
n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , 
n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , 
n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , 
n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , 
n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , 
n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3653 , n3654 , 
n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , 
n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3674 , n3675 , n3676 , 
n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , 
n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , 
n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , 
n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , 
n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , 
n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , 
n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , 
n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , 
n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , 
n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3776 , n3777 , 
n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , 
n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , 
n3798 , n3800 , n3801 , n3802 , n3803 , n3805 , n3806 , n3807 , n3808 , n3809 , 
n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , 
n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , 
n3830 , n3831 , n3832 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , 
n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , 
n3851 , n3852 , n3853 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , 
n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , 
n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , 
n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , 
n3892 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3902 , n3903 , 
n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3911 , n3912 , n3913 , n3914 , 
n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , 
n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , 
n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , 
n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , 
n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , 
n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3973 , n3974 , n3975 , 
n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , 
n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , 
n3996 , n3997 , n3998 , n3999 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , 
n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , 
n4017 , n4018 , n4019 , n4020 , n4021 , n4023 , n4024 , n4025 , n4026 , n4027 , 
n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , 
n4038 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , 
n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , 
n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , 
n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , 
n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , 
n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , 
n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , 
n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4118 , n4119 , 
n4120 , n4121 , n4122 , n4123 , n4124 , n4126 , n4127 , n4128 , n4129 , n4130 , 
n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , 
n4142 , n4143 , n4144 , n4145 , n4146 , n4148 , n4149 , n4150 , n4151 , n4152 , 
n4153 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , 
n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4173 , n4174 , 
n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , 
n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , 
n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , 
n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , 
n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4226 , 
n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , 
n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , 
n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , 
n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , 
n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , 
n4277 , n4278 , n4280 , n4281 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , 
n4289 , n4290 , n4291 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , 
n4300 , n4301 , n4302 , n4303 , n4304 , n4306 , n4307 , n4308 , n4309 , n4310 , 
n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , 
n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
n4341 , n4342 , n4343 , n4344 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , 
n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , 
n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , 
n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , 
n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , 
n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , 
n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , 
n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , 
n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , 
n4432 , n4433 , n4434 , n4435 , n4436 , n4438 , n4439 , n4440 , n4441 , n4442 , 
n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , 
n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , 
n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , 
n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , 
n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , 
n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , 
n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , 
n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , 
n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , 
n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4542 , n4543 , 
n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , 
n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , 
n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , 
n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , 
n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , 
n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , 
n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , 
n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , 
n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , 
n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , 
n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , 
n4656 , n4657 , n4658 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , 
n4667 , n4668 , n4669 , n4670 , n4671 , n4673 , n4674 , n4675 , n4676 , n4677 , 
n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , 
n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , 
n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , 
n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , 
n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , 
n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , 
n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , 
n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4756 , n4757 , n4758 , 
n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , 
n4769 , n4770 , n4771 , n4772 , n4773 , n4775 , n4776 , n4777 , n4778 , n4779 , 
n4780 , n4781 , n4782 , n4783 , n4784 , n4786 , n4787 , n4788 , n4789 , n4790 , 
n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4859 , n4860 , n4861 , 
n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , 
n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , 
n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , 
n4892 , n4893 , n4894 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , 
n4903 , n4904 , n4905 , n4906 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , 
n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , 
n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , 
n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , 
n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , 
n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , 
n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4972 , n4973 , n4974 , 
n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , 
n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , 
n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , 
n5005 , n5006 , n5007 , n5008 , n5010 , n5011 , n5012 , n5013 , n5015 , n5016 , 
n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5024 , n5025 , n5026 , n5027 , 
n5028 , n5029 , n5030 , n5031 , n5032 , n5034 , n5035 , n5036 , n5037 , n5038 , 
n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5047 , n5048 , n5049 , 
n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , 
n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , 
n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5078 , n5079 , n5080 , 
n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
n5181 , n5182 , n5183 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , 
n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , 
n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , 
n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , 
n5223 , n5224 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , 
n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , 
n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , 
n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , 
n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , 
n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , 
n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , 
n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , 
n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , 
n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , 
n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , 
n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , 
n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , 
n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , 
n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , 
n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , 
n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , 
n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , 
n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , 
n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , 
n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5431 , n5432 , n5433 , n5434 , 
n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , 
n5445 , n5446 , n5447 , n5448 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , 
n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , 
n5466 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , 
n5477 , n5478 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , 
n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , 
n5498 , n5499 , n5500 , n5501 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , 
n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , 
n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , 
n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , 
n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , 
n5549 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , 
n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , 
n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , 
n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5587 , n5588 , n5589 , n5590 , 
n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , 
n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , 
n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , 
n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , 
n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , 
n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , 
n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , 
n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , 
n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , 
n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , 
n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , 
n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , 
n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , 
n5722 , n5723 , n5724 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , 
n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , 
n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , 
n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , 
n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , 
n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , 
n5783 , n5784 , n5785 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , 
n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , 
n5804 , n5805 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , 
n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , 
n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , 
n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , 
n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5852 , n5853 , n5854 , n5855 , 
n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , 
n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , 
n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , 
n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , 
n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , 
n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , 
n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , 
n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , 
n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5944 , n5945 , n5946 , 
n5947 , n5948 , n5949 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , 
n5958 , n5959 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , 
n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , 
n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5988 , n5989 , 
n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , 
n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6008 , n6009 , n6010 , 
n6011 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , 
n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , 
n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , 
n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , 
n6052 , n6053 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , 
n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , 
n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , 
n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , 
n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , 
n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , 
n6113 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , 
n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , 
n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , 
n6144 , n6145 , n6146 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , 
n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , 
n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , 
n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , 
n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , 
n6195 , n6196 , n6197 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , 
n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , 
n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , 
n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , 
n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , 
n6246 , n6247 , n6248 , n6249 , n6250 , n6252 , n6253 , n6254 , n6255 , n6256 , 
n6257 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , 
n6268 , n6269 , n6271 , n6272 , n6273 , n6274 , n6276 , n6277 , n6278 , n6279 , 
n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , 
n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , 
n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , 
n6310 , n6311 , n6312 , n6313 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , 
n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , 
n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , 
n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , 
n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , 
n6361 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , 
n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , 
n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , 
n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , 
n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , 
n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , 
n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , 
n6432 , n6433 , n6434 , n6435 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , 
n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , 
n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6461 , n6462 , n6463 , 
n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , 
n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6481 , n6482 , n6483 , n6484 , 
n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , 
n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , 
n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , 
n6515 , n6516 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , 
n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , 
n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , 
n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6556 , 
n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , 
n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , 
n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6587 , 
n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , 
n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , 
n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , 
n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , 
n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , 
n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , 
n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , 
n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , 
n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , 
n6678 , n6679 , n6681 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , 
n6690 , n6691 , n6692 , n6694 , n6695 , n6697 , n6698 , n6699 , n6700 , n6701 , 
n6702 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , 
n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , 
n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , 
n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , 
n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , 
n6753 , n6754 , n6755 , n6756 , n6757 , n6759 , n6760 , n6761 , n6762 , n6763 , 
n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , 
n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , 
n6784 , n6785 , n6787 , n6788 , n6789 , n6790 , n6792 , n6793 , n6794 , n6795 , 
n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , 
n6806 , n6807 , n6808 , n6809 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , 
n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , 
n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , 
n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , 
n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6854 , n6855 , n6856 , n6857 , 
n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , 
n6868 , n6869 , n6870 , n6871 , n6872 , n6874 , n6875 , n6876 , n6877 , n6878 , 
n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , 
n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , 
n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , 
n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , 
n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , 
n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , 
n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6947 , n6948 , n6949 , 
n6950 , n6951 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , 
n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , 
n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6980 , n6981 , 
n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , 
n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n7000 , n7001 , n7002 , 
n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , 
n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , 
n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , 
n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , 
n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , 
n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , 
n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7072 , n7074 , 
n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , 
n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , 
n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7105 , 
n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , 
n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , 
n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7133 , n7134 , n7135 , n7136 , 
n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , 
n7147 , n7148 , n7149 , n7150 , n7151 , n7153 , n7154 , n7155 , n7156 , n7157 , 
n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , 
n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , 
n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , 
n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , 
n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , 
n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , 
n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , 
n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , 
n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7247 , n7248 , 
n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , 
n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7266 , n7267 , n7268 , n7269 , 
n7270 , n7271 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , 
n7281 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , 
n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , 
n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , 
n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , 
n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , 
n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , 
n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , 
n7352 , n7353 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , 
n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , 
n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7383 , 
n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , 
n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , 
n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , 
n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , 
n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , 
n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , 
n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7451 , n7452 , n7453 , n7454 , 
n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , 
n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , 
n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , 
n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , 
n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , 
n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , 
n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , 
n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , 
n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , 
n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , 
n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , 
n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , 
n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , 
n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , 
n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , 
n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , 
n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , 
n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , 
n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , 
n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7653 , n7654 , n7656 , 
n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , 
n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , 
n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , 
n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , 
n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , 
n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , 
n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , 
n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , 
n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , 
n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , 
n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , 
n7769 , n7770 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , 
n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , 
n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , 
n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , 
n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , 
n7820 , n7821 , n7822 , n7823 , n7824 , n7826 , n7827 , n7828 , n7829 , n7830 , 
n7831 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , 
n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , 
n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , 
n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , 
n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , 
n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , 
n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , 
n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , 
n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , 
n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , 
n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7942 , 
n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , 
n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , 
n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7973 , 
n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , 
n7984 , n7985 , n7986 , n7987 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , 
n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8003 , n8004 , n8005 , 
n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , 
n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , 
n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , 
n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8045 , n8046 , 
n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , 
n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , 
n8067 , n8069 , n8070 , n8071 , n8072 , n8074 , n8075 , n8076 , n8077 , n8078 , 
n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8086 , n8087 , n8088 , n8089 , 
n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , 
n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , 
n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , 
n8120 , n8121 , n8122 , n8123 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , 
n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , 
n8141 , n8142 , n8143 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , 
n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , 
n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , 
n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , 
n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , 
n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , 
n8202 , n8203 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , 
n8213 , n8214 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , 
n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , 
n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , 
n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , 
n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8263 , n8264 , 
n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , 
n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , 
n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , 
n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8303 , n8304 , n8305 , 
n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8316 , n8317 , 
n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , 
n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , 
n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , 
n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , 
n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , 
n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , 
n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , 
n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8398 , 
n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , 
n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , 
n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , 
n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , 
n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , 
n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , 
n8460 , n8461 , n8462 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , 
n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , 
n8482 , n8483 , n8484 , n8485 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , 
n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , 
n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , 
n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , 
n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , 
n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , 
n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8551 , n8553 , n8554 , 
n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , 
n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , 
n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , 
n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , 
n8595 , n8596 , n8597 , n8599 , n8600 , n8601 , n8602 , n8603 , n8605 , n8606 , 
n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , 
n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , 
n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8636 , n8637 , 
n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , 
n8648 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , 
n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , 
n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , 
n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , 
n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , 
n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , 
n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , 
n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , 
n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8738 , n8739 , 
n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8747 , n8748 , n8749 , n8750 , 
n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , 
n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , 
n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8781 , 
n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , 
n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8801 , n8802 , n8803 , 
n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , 
n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , 
n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , 
n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , 
n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , 
n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , 
n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8874 , 
n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , 
n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8893 , n8894 , n8895 , 
n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , 
n8906 , n8907 , n8908 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , 
n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8927 , 
n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , 
n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , 
n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , 
n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , 
n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , 
n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , 
n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8998 , 
n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , 
n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , 
n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9027 , n9028 , n9029 , 
n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , 
n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , 
n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , 
n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , 
n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , 
n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , 
n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9097 , n9098 , n9099 , n9100 , 
n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9111 , 
n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , 
n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , 
n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , 
n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , 
n9152 , n9153 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , 
n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , 
n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , 
n9183 , n9184 , n9185 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , 
n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , 
n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , 
n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , 
n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , 
n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , 
n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9253 , n9254 , 
n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , 
n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , 
n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , 
n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , 
n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , 
n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9315 , 
n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , 
n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , 
n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9343 , n9344 , n9345 , n9346 , 
n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , 
n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , 
n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , 
n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , 
n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , 
n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , 
n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , 
n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , 
n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , 
n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9448 , 
n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , 
n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , 
n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , 
n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , 
n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , 
n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , 
n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , 
n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , 
n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , 
n9539 , n9540 , n9541 , n9542 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , 
n9551 , n9552 , n9553 , n9554 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , 
n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9571 , n9572 , 
n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , 
n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9590 , n9591 , n9592 , n9593 , 
n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , 
n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , 
n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , 
n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , 
n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , 
n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , 
n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , 
n9664 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , 
n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , 
n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , 
n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , 
n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , 
n9715 , n9716 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , 
n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , 
n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , 
n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , 
n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , 
n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , 
n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , 
n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , 
n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , 
n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , 
n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , 
n9826 , n9827 , n9828 , n9829 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , 
n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , 
n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , 
n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , 
n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , 
n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , 
n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9894 , n9895 , n9896 , n9897 , 
n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , 
n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , 
n9918 , n9919 , n9920 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , 
n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9937 , n9938 , n9939 , 
n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , 
n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , 
n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , 
n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9978 , n9979 , n9980 , 
n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , 
n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , 
n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , 
n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , 
n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , 
n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , 
n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10052 , 
n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10062 , n10063 , 
n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , 
n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10081 , n10082 , n10083 , n10084 , 
n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , 
n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , 
n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10113 , n10114 , n10115 , 
n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , 
n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , 
n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , 
n10146 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , 
n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , 
n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , 
n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , 
n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , 
n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , 
n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , 
n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , 
n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , 
n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , 
n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10256 , n10257 , 
n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , 
n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , 
n10279 , n10280 , n10281 , n10282 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , 
n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , 
n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , 
n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , 
n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , 
n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , 
n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , 
n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , 
n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , 
n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10379 , n10380 , 
n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , 
n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , 
n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10408 , n10409 , n10410 , n10411 , 
n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , 
n10422 , n10423 , n10424 , n10425 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , 
n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , 
n10443 , n10444 , n10445 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , 
n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , 
n10464 , n10465 , n10467 , n10468 , n10469 , n10471 , n10472 , n10473 , n10474 , n10475 , 
n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , 
n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , 
n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , 
n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10516 , 
n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , 
n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , 
n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , 
n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , 
n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , 
n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10574 , n10575 , n10576 , n10577 , 
n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , 
n10588 , n10589 , n10590 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , 
n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , 
n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10616 , n10617 , n10618 , n10619 , 
n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , 
n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , 
n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , 
n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , 
n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , 
n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , 
n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , 
n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , 
n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , 
n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , 
n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , 
n10731 , n10732 , n10733 , n10734 , n10735 , n10737 , n10738 , n10739 , n10740 , n10741 , 
n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10751 , n10752 , 
n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , 
n10763 , n10764 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , 
n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , 
n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10792 , n10793 , n10794 , 
n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10803 , n10804 , n10805 , 
n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , 
n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , 
n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , 
n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , 
n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , 
n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10863 , n10864 , n10865 , n10866 , 
n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , 
n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , 
n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , 
n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , 
n10907 , n10908 , n10909 , n10910 , n10911 , n10913 , n10914 , n10916 , n10917 , n10918 , 
n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , 
n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , 
n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10946 , n10947 , n10948 , n10949 , 
n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , 
n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , 
n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , 
n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , 
n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , 
n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , 
n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , 
n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , 
n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , 
n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , 
n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , 
n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , 
n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , 
n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , 
n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , 
n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , 
n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , 
n11120 , n11121 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , 
n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , 
n11141 , n11142 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , 
n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11159 , n11160 , n11161 , n11162 , 
n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , 
n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , 
n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , 
n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , 
n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , 
n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , 
n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , 
n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , 
n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , 
n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , 
n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11270 , n11271 , n11272 , n11273 , 
n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , 
n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , 
n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , 
n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , 
n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , 
n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , 
n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , 
n11344 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , 
n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , 
n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , 
n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , 
n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11394 , n11395 , 
n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11405 , n11406 , 
n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , 
n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , 
n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , 
n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , 
n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , 
n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11464 , n11465 , n11466 , n11467 , 
n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , 
n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , 
n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , 
n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , 
n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , 
n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , 
n11528 , n11530 , n11531 , n11532 , n11533 , n11535 , n11536 , n11537 , n11538 , n11539 , 
n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , 
n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , 
n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , 
n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , 
n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , 
n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , 
n11601 , n11602 , n11603 , n11604 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , 
n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , 
n11622 , n11623 , n11624 , n11625 , n11626 , n11628 , n11629 , n11630 , n11631 , n11632 , 
n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , 
n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , 
n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , 
n11663 , n11665 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , 
n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , 
n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , 
n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , 
n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , 
n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , 
n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , 
n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , 
n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , 
n11755 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , 
n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , 
n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , 
n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , 
n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , 
n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , 
n11817 , n11818 , n11819 , n11820 , n11821 , n11823 , n11824 , n11825 , n11826 , n11827 , 
n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , 
n11838 , n11839 , n11840 , n11841 , n11843 , n11844 , n11845 , n11846 , n11848 , n11849 , 
n11850 , n11851 , n11852 , n11853 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , 
n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , 
n11871 , n11872 , n11873 , n11874 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , 
n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , 
n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , 
n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , 
n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , 
n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11931 , n11932 , n11934 , 
n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , 
n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , 
n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11962 , n11963 , n11964 , n11965 , 
n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , 
n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , 
n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , 
n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , 
n12006 , n12007 , n12008 , n12010 , n12011 , n12013 , n12014 , n12015 , n12016 , n12017 , 
n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12026 , n12027 , n12028 , 
n12029 , n12030 , n12031 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , 
n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , 
n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , 
n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , 
n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , 
n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , 
n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , 
n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , 
n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , 
n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , 
n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , 
n12140 , n12141 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , 
n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , 
n12161 , n12162 , n12163 , n12164 , n12165 , n12167 , n12168 , n12169 , n12170 , n12171 , 
n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , 
n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , 
n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , 
n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , 
n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12219 , n12220 , n12221 , n12222 , 
n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12233 , 
n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , 
n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , 
n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , 
n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12271 , n12272 , n12273 , n12274 , 
n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , 
n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , 
n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , 
n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , 
n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12322 , n12323 , n12324 , n12325 , 
n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , 
n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , 
n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12356 , n12357 , 
n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , 
n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , 
n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , 
n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , 
n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , 
n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , 
n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , 
n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , 
n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , 
n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , 
n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , 
n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , 
n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , 
n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , 
n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , 
n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , 
n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , 
n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12536 , n12537 , n12538 , 
n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , 
n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , 
n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , 
n12569 , n12570 , n12571 , n12572 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , 
n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , 
n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , 
n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , 
n12610 , n12611 , n12612 , n12613 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , 
n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , 
n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , 
n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , 
n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , 
n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , 
n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , 
n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , 
n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , 
n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , 
n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , 
n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , 
n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , 
n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , 
n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , 
n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , 
n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , 
n12781 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , 
n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , 
n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , 
n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , 
n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12830 , n12831 , n12832 , 
n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , 
n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , 
n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , 
n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , 
n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , 
n12883 , n12884 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , 
n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , 
n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , 
n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , 
n12924 , n12925 , n12926 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , 
n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , 
n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , 
n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , 
n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , 
n12975 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , 
n12986 , n12987 , n12988 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , 
n12997 , n12998 , n12999 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , 
n13008 , n13009 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , 
n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , 
n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , 
n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13046 , n13047 , n13048 , n13049 , 
n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , 
n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , 
n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , 
n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , 
n13090 , n13091 , n13092 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , 
n13101 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13110 , n13111 , n13112 , 
n13113 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , 
n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , 
n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13142 , n13143 , n13144 , 
n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , 
n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , 
n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , 
n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , 
n13185 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , 
n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , 
n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , 
n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13225 , n13226 , 
n13227 , n13228 , n13229 , n13230 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , 
n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , 
n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , 
n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , 
n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , 
n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , 
n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13296 , n13297 , n13298 , 
n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , 
n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13317 , n13318 , n13319 , 
n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , 
n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , 
n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , 
n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , 
n13360 , n13361 , n13362 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , 
n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , 
n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , 
n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , 
n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , 
n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , 
n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , 
n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , 
n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , 
n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , 
n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , 
n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , 
n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , 
n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , 
n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13510 , n13512 , n13513 , 
n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , 
n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , 
n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , 
n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , 
n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13562 , n13563 , n13564 , 
n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , 
n13575 , n13576 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , 
n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , 
n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , 
n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , 
n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13626 , 
n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13637 , 
n13638 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , 
n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13659 , 
n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , 
n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , 
n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , 
n13690 , n13691 , n13692 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , 
n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , 
n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , 
n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , 
n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , 
n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , 
n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13761 , 
n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , 
n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , 
n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , 
n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , 
n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , 
n13812 , n13813 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , 
n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , 
n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , 
n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , 
n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , 
n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13871 , n13872 , n13873 , n13874 , 
n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13883 , n13884 , n13885 , 
n13886 , n13887 , n13888 , n13889 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , 
n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , 
n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , 
n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , 
n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , 
n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13945 , n13946 , n13947 , 
n13948 , n13949 , n13950 , n13951 , n13952 , n13954 , n13955 , n13956 , n13957 , n13958 , 
n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , 
n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , 
n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , 
n13990 , n13991 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , 
n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , 
n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , 
n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , 
n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , 
n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , 
n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , 
n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , 
n14071 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , 
n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , 
n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , 
n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , 
n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , 
n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , 
n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , 
n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , 
n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , 
n14162 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , 
n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , 
n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , 
n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , 
n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , 
n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , 
n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , 
n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , 
n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , 
n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , 
n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , 
n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , 
n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14290 , n14291 , n14292 , n14294 , 
n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14304 , n14305 , 
n14306 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , 
n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , 
n14327 , n14328 , n14329 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , 
n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , 
n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , 
n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , 
n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , 
n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , 
n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , 
n14398 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14409 , 
n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , 
n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , 
n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , 
n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , 
n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , 
n14460 , n14461 , n14462 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , 
n14472 , n14473 , n14474 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , 
n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , 
n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , 
n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , 
n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , 
n14524 , n14525 , n14526 ;
    or g0 ( n6289 , n9151 , n3294 );
    nor g1 ( n7757 , n12807 , n10319 );
    not g2 ( n2651 , n13041 );
    or g3 ( n10364 , n12601 , n9558 );
    not g4 ( n1362 , n7322 );
    or g5 ( n6140 , n4052 , n8064 );
    not g6 ( n8630 , n13734 );
    and g7 ( n14021 , n4289 , n6390 );
    and g8 ( n6317 , n5240 , n5350 );
    or g9 ( n13791 , n4871 , n5786 );
    and g10 ( n178 , n11607 , n9635 );
    or g11 ( n1013 , n12528 , n7972 );
    and g12 ( n5244 , n406 , n40 );
    or g13 ( n2507 , n14188 , n14051 );
    nor g14 ( n10110 , n4544 , n11112 );
    and g15 ( n12465 , n13676 , n4145 );
    not g16 ( n2021 , n5795 );
    and g17 ( n180 , n4102 , n11811 );
    and g18 ( n5358 , n3986 , n2419 );
    nor g19 ( n2530 , n2597 , n7614 );
    and g20 ( n7263 , n7529 , n8354 );
    and g21 ( n9031 , n11687 , n5664 );
    nor g22 ( n12876 , n1944 , n5100 );
    not g23 ( n12900 , n5725 );
    and g24 ( n13931 , n4300 , n5032 );
    not g25 ( n9422 , n1894 );
    or g26 ( n10151 , n4967 , n8596 );
    and g27 ( n10115 , n3271 , n3260 );
    or g28 ( n2332 , n4022 , n11875 );
    or g29 ( n13604 , n5715 , n13570 );
    or g30 ( n10494 , n7116 , n7870 );
    and g31 ( n12899 , n11142 , n12366 );
    and g32 ( n12249 , n10994 , n9776 );
    and g33 ( n1389 , n12918 , n5537 );
    not g34 ( n1944 , n11302 );
    not g35 ( n14312 , n3287 );
    or g36 ( n11237 , n12870 , n9767 );
    nor g37 ( n5724 , n11180 , n2128 );
    not g38 ( n5129 , n1243 );
    or g39 ( n7303 , n12020 , n6027 );
    or g40 ( n7754 , n3804 , n7652 );
    and g41 ( n667 , n14373 , n3634 );
    nor g42 ( n1675 , n10233 , n7403 );
    and g43 ( n4909 , n4354 , n3671 );
    not g44 ( n3977 , n10824 );
    and g45 ( n1030 , n5229 , n8184 );
    nor g46 ( n1263 , n9806 , n9496 );
    and g47 ( n10882 , n14042 , n2697 );
    or g48 ( n10974 , n10871 , n12320 );
    or g49 ( n13428 , n11558 , n7538 );
    and g50 ( n7180 , n13103 , n12346 );
    or g51 ( n10950 , n976 , n437 );
    not g52 ( n2889 , n13425 );
    and g53 ( n5592 , n4098 , n3065 );
    or g54 ( n10914 , n10808 , n13594 );
    and g55 ( n9665 , n13511 , n9733 );
    and g56 ( n4403 , n8801 , n10549 );
    or g57 ( n13412 , n13083 , n942 );
    and g58 ( n7567 , n14286 , n7644 );
    not g59 ( n781 , n7339 );
    or g60 ( n2362 , n3093 , n3943 );
    not g61 ( n6672 , n6357 );
    or g62 ( n14005 , n5236 , n11954 );
    and g63 ( n7129 , n13297 , n187 );
    or g64 ( n5481 , n2949 , n9091 );
    nor g65 ( n32 , n4913 , n8126 );
    and g66 ( n4943 , n3212 , n4990 );
    nor g67 ( n9606 , n1473 , n6423 );
    and g68 ( n6879 , n2177 , n2552 );
    not g69 ( n8081 , n4036 );
    or g70 ( n13550 , n10960 , n5342 );
    or g71 ( n3660 , n1137 , n11790 );
    and g72 ( n7712 , n14093 , n5157 );
    not g73 ( n1612 , n3572 );
    or g74 ( n8287 , n9229 , n7331 );
    or g75 ( n10768 , n11647 , n1547 );
    not g76 ( n1571 , n8357 );
    or g77 ( n10012 , n6383 , n10051 );
    not g78 ( n8432 , n8524 );
    or g79 ( n3531 , n8376 , n9589 );
    and g80 ( n114 , n4851 , n14280 );
    or g81 ( n13990 , n13507 , n6436 );
    or g82 ( n1358 , n12401 , n5643 );
    nor g83 ( n13163 , n4924 , n5324 );
    and g84 ( n4951 , n4856 , n6884 );
    or g85 ( n4953 , n666 , n13511 );
    and g86 ( n13989 , n4433 , n12947 );
    and g87 ( n6927 , n4422 , n7485 );
    or g88 ( n12632 , n13220 , n7191 );
    and g89 ( n1237 , n10763 , n14040 );
    nor g90 ( n11299 , n7011 , n12162 );
    not g91 ( n6595 , n5627 );
    not g92 ( n8048 , n12014 );
    or g93 ( n1817 , n9375 , n5095 );
    not g94 ( n3861 , n2958 );
    and g95 ( n10345 , n5092 , n5407 );
    and g96 ( n10477 , n7421 , n3669 );
    or g97 ( n6283 , n9353 , n11650 );
    or g98 ( n8753 , n13087 , n4518 );
    not g99 ( n7689 , n7056 );
    not g100 ( n11411 , n4266 );
    or g101 ( n8957 , n14282 , n12902 );
    or g102 ( n3822 , n11345 , n5786 );
    or g103 ( n10518 , n14450 , n10147 );
    not g104 ( n5897 , n13967 );
    nor g105 ( n2125 , n12904 , n10607 );
    nor g106 ( n9733 , n5237 , n8944 );
    and g107 ( n3022 , n6822 , n9199 );
    or g108 ( n13113 , n11710 , n7021 );
    not g109 ( n230 , n5178 );
    or g110 ( n2015 , n9140 , n13351 );
    or g111 ( n5150 , n10019 , n6737 );
    nor g112 ( n10329 , n13356 , n9372 );
    or g113 ( n14316 , n7219 , n6307 );
    or g114 ( n2931 , n5064 , n4181 );
    not g115 ( n14134 , n7940 );
    and g116 ( n3978 , n8950 , n7597 );
    or g117 ( n10926 , n5807 , n12141 );
    or g118 ( n2400 , n8908 , n11465 );
    or g119 ( n3379 , n5064 , n4227 );
    and g120 ( n3473 , n14260 , n4003 );
    and g121 ( n4506 , n1876 , n13713 );
    or g122 ( n1570 , n2878 , n2225 );
    not g123 ( n7120 , n9193 );
    and g124 ( n4303 , n14321 , n515 );
    nor g125 ( n7496 , n8189 , n12030 );
    nor g126 ( n13881 , n906 , n11277 );
    not g127 ( n8378 , n409 );
    and g128 ( n10354 , n55 , n876 );
    or g129 ( n671 , n6242 , n10752 );
    or g130 ( n10988 , n14419 , n7643 );
    not g131 ( n9461 , n10395 );
    and g132 ( n1521 , n13555 , n5463 );
    nor g133 ( n9282 , n4195 , n5747 );
    and g134 ( n923 , n2533 , n872 );
    or g135 ( n475 , n14366 , n43 );
    or g136 ( n10159 , n10461 , n11364 );
    not g137 ( n742 , n241 );
    or g138 ( n2487 , n8582 , n4719 );
    and g139 ( n6976 , n2224 , n13663 );
    and g140 ( n11242 , n7957 , n7138 );
    or g141 ( n13973 , n3394 , n13859 );
    and g142 ( n10150 , n14313 , n8116 );
    nor g143 ( n6327 , n6672 , n12268 );
    or g144 ( n8613 , n5450 , n6229 );
    or g145 ( n13372 , n12353 , n12385 );
    and g146 ( n4979 , n14213 , n13576 );
    or g147 ( n5403 , n3886 , n13790 );
    or g148 ( n10140 , n10560 , n3600 );
    and g149 ( n7473 , n13297 , n6951 );
    or g150 ( n1260 , n12768 , n8737 );
    or g151 ( n12910 , n2888 , n3360 );
    nor g152 ( n11192 , n9795 , n14259 );
    and g153 ( n2440 , n286 , n6562 );
    or g154 ( n9122 , n12100 , n3017 );
    or g155 ( n6330 , n5234 , n9338 );
    and g156 ( n577 , n8412 , n9010 );
    and g157 ( n5991 , n1539 , n8103 );
    not g158 ( n13206 , n1813 );
    or g159 ( n3358 , n13698 , n12441 );
    not g160 ( n11824 , n730 );
    and g161 ( n8532 , n1431 , n9764 );
    or g162 ( n1239 , n3667 , n7380 );
    or g163 ( n5700 , n6350 , n11949 );
    and g164 ( n9728 , n10589 , n7148 );
    or g165 ( n8319 , n3419 , n13363 );
    not g166 ( n234 , n12489 );
    or g167 ( n12215 , n9806 , n3147 );
    not g168 ( n1210 , n427 );
    or g169 ( n13229 , n2949 , n12427 );
    and g170 ( n5227 , n13367 , n13687 );
    and g171 ( n5884 , n6016 , n4531 );
    not g172 ( n13142 , n3455 );
    not g173 ( n10751 , n6989 );
    or g174 ( n4124 , n3025 , n13332 );
    or g175 ( n6783 , n14107 , n1670 );
    and g176 ( n10728 , n3766 , n10226 );
    not g177 ( n12046 , n2503 );
    or g178 ( n14459 , n12047 , n3153 );
    nor g179 ( n10148 , n13977 , n12002 );
    not g180 ( n225 , n13734 );
    or g181 ( n10452 , n5570 , n2786 );
    and g182 ( n4081 , n646 , n12722 );
    or g183 ( n14045 , n1821 , n1663 );
    and g184 ( n6055 , n6937 , n5756 );
    or g185 ( n5661 , n14449 , n13228 );
    or g186 ( n2053 , n390 , n3250 );
    nor g187 ( n1666 , n12453 , n1611 );
    nor g188 ( n5425 , n5209 , n3973 );
    and g189 ( n7269 , n9297 , n3135 );
    not g190 ( n1247 , n4535 );
    nor g191 ( n11078 , n12087 , n266 );
    not g192 ( n9429 , n11541 );
    or g193 ( n13292 , n163 , n7679 );
    not g194 ( n11582 , n9046 );
    or g195 ( n119 , n5139 , n112 );
    not g196 ( n7886 , n316 );
    not g197 ( n14368 , n9679 );
    and g198 ( n9468 , n12039 , n4393 );
    and g199 ( n10145 , n1520 , n12538 );
    and g200 ( n8413 , n1254 , n176 );
    and g201 ( n7977 , n7391 , n10720 );
    not g202 ( n2850 , n1706 );
    and g203 ( n13895 , n3715 , n13290 );
    or g204 ( n5453 , n2901 , n11010 );
    nor g205 ( n5577 , n900 , n1159 );
    nor g206 ( n3528 , n7551 , n4673 );
    and g207 ( n5191 , n1489 , n3415 );
    nor g208 ( n7459 , n13707 , n12055 );
    nor g209 ( n4201 , n14058 , n7577 );
    not g210 ( n5876 , n14135 );
    or g211 ( n132 , n12820 , n12260 );
    nor g212 ( n6384 , n13361 , n1887 );
    or g213 ( n12909 , n2608 , n6270 );
    and g214 ( n4115 , n6649 , n1186 );
    or g215 ( n6694 , n1051 , n13427 );
    and g216 ( n7923 , n12335 , n566 );
    and g217 ( n9196 , n3424 , n13690 );
    and g218 ( n9257 , n7961 , n14348 );
    and g219 ( n3378 , n14063 , n1429 );
    not g220 ( n904 , n5675 );
    or g221 ( n7591 , n12994 , n4852 );
    nor g222 ( n3557 , n2417 , n5339 );
    and g223 ( n3007 , n9041 , n53 );
    or g224 ( n13692 , n9375 , n292 );
    or g225 ( n11829 , n9218 , n1730 );
    or g226 ( n9459 , n747 , n14064 );
    nor g227 ( n12492 , n14216 , n11505 );
    not g228 ( n7739 , n12846 );
    or g229 ( n2077 , n10089 , n4450 );
    or g230 ( n599 , n2055 , n3975 );
    or g231 ( n621 , n3134 , n11268 );
    or g232 ( n6340 , n12759 , n14415 );
    not g233 ( n2958 , n744 );
    or g234 ( n9993 , n13718 , n2296 );
    and g235 ( n8041 , n1662 , n9420 );
    or g236 ( n13836 , n1480 , n8774 );
    and g237 ( n9379 , n12721 , n6215 );
    and g238 ( n10898 , n6649 , n7074 );
    not g239 ( n2692 , n2520 );
    or g240 ( n5328 , n28 , n1759 );
    and g241 ( n7005 , n1071 , n8665 );
    nor g242 ( n2054 , n10535 , n11034 );
    and g243 ( n5117 , n2067 , n6643 );
    and g244 ( n5794 , n1140 , n4191 );
    or g245 ( n5551 , n839 , n3185 );
    and g246 ( n3416 , n9920 , n11878 );
    and g247 ( n11617 , n2608 , n12132 );
    not g248 ( n5873 , n4022 );
    nor g249 ( n14485 , n4092 , n5385 );
    and g250 ( n14203 , n14227 , n13897 );
    and g251 ( n8222 , n392 , n11789 );
    not g252 ( n2784 , n7086 );
    or g253 ( n7805 , n3047 , n5590 );
    not g254 ( n8401 , n7275 );
    and g255 ( n9719 , n9564 , n1104 );
    not g256 ( n10930 , n14075 );
    and g257 ( n7762 , n8025 , n12129 );
    or g258 ( n4832 , n5800 , n9845 );
    not g259 ( n10338 , n3577 );
    or g260 ( n4103 , n6891 , n12575 );
    and g261 ( n13822 , n3952 , n10487 );
    and g262 ( n4028 , n12460 , n5859 );
    and g263 ( n4453 , n1339 , n7868 );
    and g264 ( n8514 , n13103 , n7290 );
    or g265 ( n12004 , n850 , n12983 );
    not g266 ( n3182 , n14164 );
    and g267 ( n11464 , n13952 , n12180 );
    or g268 ( n12070 , n2597 , n2062 );
    nor g269 ( n6184 , n3034 , n6131 );
    and g270 ( n9658 , n13650 , n1748 );
    not g271 ( n10730 , n13158 );
    and g272 ( n11610 , n8431 , n11351 );
    and g273 ( n14151 , n4844 , n2140 );
    or g274 ( n9814 , n13675 , n13972 );
    or g275 ( n1947 , n5084 , n8260 );
    not g276 ( n13399 , n2409 );
    and g277 ( n11778 , n12808 , n11452 );
    not g278 ( n5800 , n5242 );
    or g279 ( n12124 , n11048 , n9473 );
    not g280 ( n5432 , n13752 );
    and g281 ( n356 , n679 , n11927 );
    nor g282 ( n10349 , n9810 , n1469 );
    not g283 ( n6119 , n7533 );
    and g284 ( n6187 , n2985 , n11919 );
    and g285 ( n12032 , n8550 , n11192 );
    or g286 ( n8367 , n6109 , n2070 );
    not g287 ( n7808 , n10603 );
    nor g288 ( n3524 , n9124 , n1323 );
    or g289 ( n10771 , n12023 , n9312 );
    or g290 ( n7945 , n5587 , n4516 );
    or g291 ( n4219 , n8638 , n829 );
    or g292 ( n6543 , n7250 , n9003 );
    and g293 ( n3081 , n11411 , n3788 );
    or g294 ( n3507 , n11048 , n14513 );
    and g295 ( n5701 , n13535 , n1630 );
    and g296 ( n11650 , n406 , n2019 );
    or g297 ( n10677 , n7011 , n8863 );
    not g298 ( n11094 , n11415 );
    or g299 ( n1128 , n2897 , n12487 );
    or g300 ( n1493 , n1051 , n13543 );
    not g301 ( n4856 , n2744 );
    and g302 ( n5692 , n3607 , n10293 );
    not g303 ( n12075 , n11152 );
    nor g304 ( n6194 , n12087 , n3436 );
    not g305 ( n2761 , n1676 );
    or g306 ( n807 , n1844 , n14232 );
    or g307 ( n11565 , n10300 , n5433 );
    and g308 ( n3945 , n6822 , n2377 );
    and g309 ( n4966 , n8252 , n12430 );
    or g310 ( n12554 , n283 , n7190 );
    or g311 ( n7001 , n12353 , n1384 );
    and g312 ( n9647 , n2985 , n3283 );
    or g313 ( n563 , n2857 , n7982 );
    and g314 ( n7089 , n406 , n13 );
    or g315 ( n9258 , n10331 , n8968 );
    not g316 ( n1697 , n1220 );
    and g317 ( n10039 , n11028 , n7268 );
    not g318 ( n7919 , n13437 );
    or g319 ( n2773 , n11011 , n3246 );
    or g320 ( n12803 , n2790 , n11480 );
    not g321 ( n11048 , n11152 );
    not g322 ( n14245 , n12336 );
    and g323 ( n13564 , n889 , n2585 );
    or g324 ( n11789 , n6730 , n3299 );
    nor g325 ( n6081 , n12693 , n1782 );
    or g326 ( n13036 , n10351 , n7918 );
    and g327 ( n693 , n6854 , n13957 );
    and g328 ( n13901 , n1161 , n13128 );
    and g329 ( n5877 , n10134 , n4955 );
    or g330 ( n3982 , n4978 , n7155 );
    or g331 ( n6574 , n7122 , n6722 );
    or g332 ( n6648 , n11036 , n11273 );
    not g333 ( n6849 , n10466 );
    and g334 ( n8064 , n13236 , n13216 );
    not g335 ( n7519 , n11792 );
    or g336 ( n3555 , n7862 , n10379 );
    or g337 ( n4229 , n2510 , n3878 );
    and g338 ( n9680 , n4880 , n10324 );
    or g339 ( n3836 , n13446 , n7487 );
    and g340 ( n2578 , n13952 , n9827 );
    and g341 ( n13748 , n10072 , n11126 );
    and g342 ( n11639 , n2682 , n9993 );
    not g343 ( n4865 , n3542 );
    or g344 ( n2712 , n7003 , n1270 );
    not g345 ( n2643 , n11715 );
    or g346 ( n4834 , n13806 , n10935 );
    and g347 ( n3433 , n13656 , n9333 );
    and g348 ( n8535 , n3635 , n1216 );
    and g349 ( n5541 , n13877 , n10725 );
    and g350 ( n13660 , n11569 , n9112 );
    and g351 ( n1528 , n13555 , n9034 );
    or g352 ( n6880 , n8908 , n2496 );
    and g353 ( n1930 , n13433 , n11344 );
    not g354 ( n6822 , n6559 );
    or g355 ( n5349 , n3193 , n3142 );
    or g356 ( n8956 , n11360 , n12596 );
    and g357 ( n6526 , n10710 , n5965 );
    not g358 ( n766 , n4317 );
    and g359 ( n3026 , n1339 , n8846 );
    not g360 ( n7575 , n8565 );
    not g361 ( n6109 , n4606 );
    and g362 ( n12245 , n2983 , n8614 );
    and g363 ( n5293 , n11867 , n2411 );
    or g364 ( n2093 , n3800 , n8935 );
    not g365 ( n7238 , n11071 );
    and g366 ( n10169 , n10032 , n3656 );
    nor g367 ( n3716 , n12934 , n3464 );
    or g368 ( n5013 , n14404 , n9774 );
    or g369 ( n3422 , n6781 , n13546 );
    and g370 ( n1624 , n13069 , n8837 );
    nor g371 ( n9847 , n1697 , n8720 );
    or g372 ( n13517 , n6288 , n14169 );
    or g373 ( n12662 , n4407 , n10223 );
    nor g374 ( n164 , n8378 , n3964 );
    and g375 ( n7866 , n2099 , n14226 );
    and g376 ( n7440 , n8630 , n140 );
    and g377 ( n4434 , n12013 , n8017 );
    or g378 ( n4669 , n511 , n6553 );
    and g379 ( n3190 , n8066 , n1913 );
    or g380 ( n5256 , n7612 , n12573 );
    and g381 ( n97 , n1876 , n14338 );
    or g382 ( n469 , n10224 , n12365 );
    and g383 ( n10299 , n80 , n11237 );
    and g384 ( n8893 , n8427 , n3178 );
    and g385 ( n2447 , n5999 , n13452 );
    or g386 ( n2106 , n12278 , n7466 );
    or g387 ( n464 , n838 , n9489 );
    or g388 ( n11193 , n10960 , n12073 );
    and g389 ( n2723 , n4573 , n11068 );
    or g390 ( n11344 , n4180 , n9316 );
    not g391 ( n4244 , n7681 );
    nor g392 ( n4477 , n10323 , n2988 );
    or g393 ( n8706 , n10846 , n14408 );
    or g394 ( n7036 , n7354 , n13363 );
    or g395 ( n11846 , n1147 , n5771 );
    and g396 ( n1824 , n1489 , n863 );
    not g397 ( n4554 , n4135 );
    and g398 ( n3256 , n2724 , n11973 );
    and g399 ( n14179 , n7627 , n6188 );
    or g400 ( n7260 , n5603 , n3385 );
    and g401 ( n6220 , n10072 , n12861 );
    and g402 ( n7201 , n6389 , n10895 );
    or g403 ( n10990 , n4468 , n13479 );
    not g404 ( n2608 , n9830 );
    not g405 ( n8897 , n8148 );
    or g406 ( n4074 , n12428 , n14142 );
    or g407 ( n11295 , n4033 , n12341 );
    or g408 ( n8394 , n8045 , n9419 );
    and g409 ( n1025 , n1047 , n1208 );
    and g410 ( n3373 , n2587 , n7554 );
    and g411 ( n5161 , n5279 , n267 );
    and g412 ( n9966 , n3491 , n4649 );
    not g413 ( n12998 , n5268 );
    or g414 ( n9487 , n2098 , n1314 );
    and g415 ( n2385 , n3268 , n1503 );
    or g416 ( n2683 , n3559 , n4351 );
    and g417 ( n10172 , n14286 , n10157 );
    or g418 ( n2944 , n10035 , n5555 );
    or g419 ( n8826 , n769 , n7520 );
    or g420 ( n11318 , n69 , n4870 );
    nor g421 ( n1403 , n2889 , n606 );
    and g422 ( n1719 , n405 , n6165 );
    and g423 ( n12980 , n776 , n3930 );
    or g424 ( n8924 , n3320 , n14340 );
    and g425 ( n12466 , n5459 , n7869 );
    and g426 ( n4603 , n12092 , n14361 );
    not g427 ( n1478 , n10047 );
    not g428 ( n873 , n5153 );
    not g429 ( n1193 , n13003 );
    or g430 ( n9554 , n10834 , n941 );
    and g431 ( n14229 , n14450 , n13415 );
    and g432 ( n3295 , n12460 , n13188 );
    nor g433 ( n8617 , n9601 , n1954 );
    or g434 ( n14226 , n10019 , n10727 );
    and g435 ( n6709 , n405 , n4701 );
    not g436 ( n1914 , n13901 );
    and g437 ( n12916 , n5825 , n8525 );
    or g438 ( n4875 , n11048 , n13872 );
    or g439 ( n9166 , n10136 , n4505 );
    and g440 ( n10531 , n5252 , n9116 );
    and g441 ( n10629 , n752 , n9465 );
    or g442 ( n12777 , n12820 , n13918 );
    and g443 ( n8934 , n2587 , n7878 );
    and g444 ( n12734 , n9972 , n764 );
    not g445 ( n412 , n3357 );
    or g446 ( n6291 , n5472 , n756 );
    nor g447 ( n3421 , n4877 , n3997 );
    and g448 ( n2640 , n5458 , n9397 );
    nor g449 ( n527 , n7886 , n8388 );
    and g450 ( n8554 , n1924 , n13923 );
    or g451 ( n12658 , n848 , n9936 );
    and g452 ( n13493 , n5317 , n6890 );
    or g453 ( n11181 , n8332 , n72 );
    or g454 ( n11082 , n28 , n7947 );
    and g455 ( n9757 , n350 , n8365 );
    or g456 ( n7119 , n12543 , n4040 );
    not g457 ( n6981 , n977 );
    or g458 ( n1279 , n4923 , n13750 );
    or g459 ( n12954 , n8747 , n6571 );
    nor g460 ( n6841 , n9305 , n13053 );
    or g461 ( n6115 , n6350 , n1968 );
    or g462 ( n11399 , n5236 , n11899 );
    or g463 ( n8526 , n1137 , n10910 );
    not g464 ( n6288 , n9959 );
    and g465 ( n2909 , n7768 , n3127 );
    nor g466 ( n9318 , n11697 , n4975 );
    and g467 ( n1395 , n7171 , n2627 );
    nor g468 ( n5958 , n4978 , n2189 );
    and g469 ( n14037 , n4790 , n3993 );
    and g470 ( n145 , n904 , n14224 );
    and g471 ( n12196 , n2783 , n9599 );
    nor g472 ( n5376 , n1127 , n725 );
    not g473 ( n9613 , n2816 );
    nor g474 ( n6048 , n1771 , n4696 );
    or g475 ( n10667 , n11176 , n2551 );
    and g476 ( n10802 , n13186 , n6448 );
    or g477 ( n1499 , n4128 , n10292 );
    or g478 ( n5924 , n5450 , n14448 );
    and g479 ( n12188 , n6649 , n3300 );
    nor g480 ( n4694 , n13875 , n7606 );
    and g481 ( n6928 , n400 , n10231 );
    or g482 ( n3086 , n14319 , n11596 );
    and g483 ( n7404 , n11654 , n6742 );
    and g484 ( n7811 , n10660 , n8706 );
    or g485 ( n11502 , n1660 , n167 );
    or g486 ( n3392 , n6206 , n5604 );
    and g487 ( n13934 , n7717 , n7218 );
    and g488 ( n6701 , n5048 , n9957 );
    nor g489 ( n9444 , n13283 , n2522 );
    or g490 ( n12115 , n5493 , n2632 );
    and g491 ( n13161 , n12039 , n4141 );
    and g492 ( n5043 , n8247 , n4964 );
    or g493 ( n3729 , n14430 , n13320 );
    not g494 ( n6434 , n10529 );
    and g495 ( n12313 , n13404 , n9528 );
    or g496 ( n14182 , n11576 , n10594 );
    and g497 ( n8745 , n432 , n10504 );
    not g498 ( n1489 , n5525 );
    and g499 ( n13479 , n7691 , n7504 );
    or g500 ( n12168 , n9206 , n5449 );
    nor g501 ( n13337 , n12922 , n5654 );
    nor g502 ( n13009 , n4144 , n12878 );
    and g503 ( n8794 , n3419 , n6144 );
    not g504 ( n7745 , n3926 );
    not g505 ( n13317 , n12909 );
    and g506 ( n1618 , n10408 , n5903 );
    and g507 ( n12128 , n9232 , n6621 );
    or g508 ( n12713 , n7898 , n8776 );
    and g509 ( n5423 , n7392 , n8292 );
    and g510 ( n10167 , n13700 , n12108 );
    and g511 ( n2516 , n7208 , n10836 );
    nor g512 ( n3726 , n6266 , n2854 );
    not g513 ( n8786 , n230 );
    and g514 ( n4312 , n2904 , n5506 );
    or g515 ( n11146 , n7708 , n8302 );
    or g516 ( n8570 , n13854 , n8954 );
    nor g517 ( n5597 , n1713 , n10604 );
    and g518 ( n12043 , n4788 , n1923 );
    and g519 ( n13601 , n12620 , n6983 );
    and g520 ( n2728 , n10458 , n7110 );
    and g521 ( n7283 , n5948 , n10778 );
    nor g522 ( n7841 , n12403 , n11898 );
    not g523 ( n11676 , n8598 );
    and g524 ( n2223 , n4175 , n6721 );
    and g525 ( n3571 , n2461 , n2526 );
    and g526 ( n382 , n2788 , n12304 );
    or g527 ( n104 , n13074 , n7797 );
    not g528 ( n11861 , n11195 );
    or g529 ( n8652 , n7887 , n4387 );
    nor g530 ( n1492 , n5762 , n7582 );
    not g531 ( n9984 , n1267 );
    nor g532 ( n1910 , n3768 , n13378 );
    or g533 ( n324 , n4195 , n1732 );
    and g534 ( n11500 , n10855 , n4680 );
    nor g535 ( n10373 , n12075 , n8143 );
    and g536 ( n7205 , n8358 , n14184 );
    and g537 ( n404 , n12057 , n13773 );
    nor g538 ( n8943 , n4877 , n11260 );
    or g539 ( n3668 , n8816 , n4916 );
    and g540 ( n11187 , n3370 , n5682 );
    and g541 ( n7543 , n965 , n2105 );
    or g542 ( n2836 , n747 , n12867 );
    nor g543 ( n14526 , n4829 , n13632 );
    and g544 ( n4737 , n2224 , n10514 );
    or g545 ( n2009 , n8799 , n12614 );
    not g546 ( n9795 , n2772 );
    not g547 ( n1813 , n2371 );
    or g548 ( n11691 , n8581 , n11461 );
    or g549 ( n10794 , n12292 , n6440 );
    or g550 ( n13689 , n6205 , n9237 );
    or g551 ( n11061 , n6046 , n9434 );
    nor g552 ( n2844 , n8301 , n7105 );
    not g553 ( n5266 , n5901 );
    and g554 ( n10835 , n2330 , n6599 );
    or g555 ( n5464 , n1061 , n8585 );
    or g556 ( n10117 , n11303 , n2078 );
    and g557 ( n9961 , n6192 , n269 );
    and g558 ( n5173 , n4098 , n12914 );
    or g559 ( n4495 , n8986 , n4768 );
    nor g560 ( n7013 , n11094 , n8982 );
    or g561 ( n10777 , n2149 , n3295 );
    and g562 ( n4613 , n6016 , n8254 );
    and g563 ( n5629 , n3405 , n9298 );
    nor g564 ( n10739 , n12705 , n10235 );
    and g565 ( n1132 , n286 , n4190 );
    or g566 ( n1698 , n4908 , n6550 );
    and g567 ( n8030 , n8393 , n5346 );
    or g568 ( n2565 , n4407 , n6591 );
    and g569 ( n17 , n11679 , n7635 );
    and g570 ( n3314 , n1266 , n4411 );
    and g571 ( n1673 , n4394 , n11528 );
    nor g572 ( n3937 , n8663 , n10952 );
    not g573 ( n5409 , n1833 );
    or g574 ( n1191 , n228 , n10137 );
    or g575 ( n6861 , n9819 , n1093 );
    or g576 ( n5270 , n4435 , n11855 );
    and g577 ( n3240 , n11157 , n3690 );
    and g578 ( n6921 , n10338 , n8915 );
    or g579 ( n3711 , n11724 , n136 );
    and g580 ( n7592 , n687 , n3379 );
    and g581 ( n10979 , n14351 , n12137 );
    and g582 ( n13577 , n9110 , n467 );
    and g583 ( n4332 , n8702 , n10389 );
    and g584 ( n2472 , n3233 , n11617 );
    and g585 ( n4505 , n4095 , n10545 );
    nor g586 ( n4079 , n7904 , n12430 );
    and g587 ( n3855 , n12335 , n9676 );
    and g588 ( n7836 , n2942 , n5452 );
    or g589 ( n12547 , n976 , n6924 );
    or g590 ( n10698 , n14404 , n9222 );
    and g591 ( n3714 , n8250 , n9777 );
    or g592 ( n10702 , n13847 , n9860 );
    and g593 ( n2120 , n4574 , n14185 );
    or g594 ( n896 , n2179 , n4587 );
    and g595 ( n115 , n14210 , n10000 );
    or g596 ( n8297 , n7462 , n5215 );
    and g597 ( n12516 , n12015 , n2392 );
    not g598 ( n3361 , n13983 );
    or g599 ( n661 , n13991 , n14444 );
    not g600 ( n3640 , n8899 );
    nor g601 ( n14019 , n3822 , n11763 );
    not g602 ( n6975 , n2011 );
    and g603 ( n14493 , n10855 , n12796 );
    or g604 ( n11750 , n9807 , n7713 );
    not g605 ( n8582 , n2918 );
    not g606 ( n4871 , n3532 );
    or g607 ( n10850 , n2229 , n8077 );
    and g608 ( n4011 , n12226 , n1510 );
    or g609 ( n7341 , n11722 , n10826 );
    and g610 ( n13559 , n8043 , n13280 );
    and g611 ( n3514 , n1854 , n2839 );
    and g612 ( n12177 , n501 , n4192 );
    and g613 ( n2169 , n2064 , n13292 );
    not g614 ( n5172 , n521 );
    and g615 ( n9895 , n2587 , n1067 );
    and g616 ( n4387 , n406 , n10926 );
    nor g617 ( n14390 , n882 , n11671 );
    and g618 ( n5663 , n4382 , n7758 );
    or g619 ( n6100 , n7914 , n1146 );
    not g620 ( n5468 , n3007 );
    or g621 ( n12578 , n6373 , n8588 );
    not g622 ( n7418 , n11456 );
    or g623 ( n9810 , n4147 , n10378 );
    or g624 ( n5121 , n5570 , n6800 );
    nor g625 ( n4 , n6797 , n8449 );
    nor g626 ( n11709 , n5365 , n4645 );
    nor g627 ( n11796 , n1480 , n6646 );
    and g628 ( n2777 , n1354 , n14105 );
    nor g629 ( n10554 , n13201 , n10900 );
    and g630 ( n260 , n4422 , n7330 );
    not g631 ( n12092 , n13383 );
    and g632 ( n12444 , n6536 , n510 );
    nor g633 ( n6094 , n14370 , n6918 );
    not g634 ( n320 , n5950 );
    nor g635 ( n6502 , n8592 , n13214 );
    and g636 ( n10738 , n12092 , n8725 );
    not g637 ( n4498 , n12249 );
    or g638 ( n3108 , n2747 , n9173 );
    or g639 ( n2205 , n172 , n1704 );
    and g640 ( n5272 , n2330 , n9857 );
    nor g641 ( n3380 , n11998 , n10655 );
    or g642 ( n3218 , n6271 , n6748 );
    not g643 ( n7678 , n238 );
    not g644 ( n12918 , n13219 );
    and g645 ( n5167 , n6128 , n9161 );
    not g646 ( n4233 , n4465 );
    and g647 ( n1087 , n9724 , n1516 );
    or g648 ( n3860 , n9442 , n12550 );
    and g649 ( n11390 , n13107 , n677 );
    not g650 ( n3099 , n5974 );
    and g651 ( n12309 , n12229 , n5988 );
    or g652 ( n4707 , n5507 , n12775 );
    or g653 ( n149 , n7003 , n5746 );
    and g654 ( n12386 , n7779 , n372 );
    and g655 ( n4198 , n7203 , n14445 );
    and g656 ( n12383 , n6135 , n12788 );
    not g657 ( n6754 , n11975 );
    nor g658 ( n3848 , n11325 , n11999 );
    or g659 ( n12816 , n11576 , n5367 );
    nor g660 ( n1954 , n9035 , n7143 );
    not g661 ( n8115 , n6074 );
    and g662 ( n5872 , n348 , n13207 );
    and g663 ( n6071 , n1427 , n6005 );
    and g664 ( n842 , n7826 , n12497 );
    or g665 ( n9884 , n11951 , n5136 );
    or g666 ( n8411 , n5936 , n485 );
    and g667 ( n2210 , n4757 , n13143 );
    nor g668 ( n4396 , n5780 , n14243 );
    and g669 ( n721 , n4581 , n1008 );
    or g670 ( n4441 , n11804 , n4436 );
    and g671 ( n3597 , n2643 , n9761 );
    and g672 ( n2273 , n7826 , n9538 );
    or g673 ( n12792 , n6109 , n10060 );
    or g674 ( n1785 , n12549 , n13614 );
    not g675 ( n12933 , n12321 );
    not g676 ( n1588 , n8656 );
    nor g677 ( n13273 , n5468 , n4063 );
    or g678 ( n4370 , n3161 , n531 );
    or g679 ( n214 , n5800 , n1877 );
    and g680 ( n3055 , n8300 , n3570 );
    and g681 ( n10463 , n3405 , n2013 );
    not g682 ( n2808 , n4510 );
    and g683 ( n2502 , n1117 , n3617 );
    nor g684 ( n13159 , n3546 , n2345 );
    or g685 ( n12991 , n2315 , n2196 );
    or g686 ( n10037 , n7898 , n2388 );
    and g687 ( n5882 , n1904 , n9221 );
    not g688 ( n7419 , n1478 );
    not g689 ( n12304 , n13714 );
    or g690 ( n9271 , n12759 , n7730 );
    and g691 ( n2364 , n4347 , n14462 );
    or g692 ( n9120 , n4340 , n3391 );
    or g693 ( n190 , n1362 , n13031 );
    and g694 ( n9867 , n14351 , n10891 );
    and g695 ( n12272 , n6848 , n1165 );
    not g696 ( n7026 , n6559 );
    nor g697 ( n11371 , n11259 , n5199 );
    and g698 ( n3220 , n14465 , n6775 );
    or g699 ( n1422 , n13155 , n10526 );
    not g700 ( n7809 , n9231 );
    and g701 ( n3312 , n10595 , n4616 );
    or g702 ( n12432 , n8096 , n8955 );
    or g703 ( n7044 , n116 , n8634 );
    not g704 ( n7430 , n11331 );
    or g705 ( n1835 , n8396 , n1078 );
    not g706 ( n13823 , n4928 );
    or g707 ( n9264 , n7430 , n12418 );
    or g708 ( n5021 , n900 , n7746 );
    not g709 ( n14110 , n12687 );
    or g710 ( n2732 , n3826 , n12234 );
    or g711 ( n12602 , n1261 , n3448 );
    and g712 ( n3297 , n904 , n6876 );
    or g713 ( n8150 , n5406 , n1931 );
    or g714 ( n4026 , n850 , n7964 );
    not g715 ( n6848 , n4292 );
    or g716 ( n4817 , n5493 , n10948 );
    and g717 ( n3481 , n12013 , n8788 );
    and g718 ( n13315 , n10357 , n14140 );
    or g719 ( n4676 , n12625 , n1963 );
    and g720 ( n471 , n6753 , n7119 );
    and g721 ( n6557 , n3405 , n4420 );
    or g722 ( n14138 , n7358 , n8281 );
    or g723 ( n6107 , n2315 , n8808 );
    and g724 ( n877 , n3942 , n9346 );
    and g725 ( n4830 , n11676 , n6408 );
    not g726 ( n14377 , n9721 );
    and g727 ( n6262 , n12185 , n6717 );
    and g728 ( n5723 , n3169 , n5211 );
    and g729 ( n12026 , n13362 , n12597 );
    or g730 ( n12285 , n4908 , n471 );
    nor g731 ( n8874 , n11580 , n6191 );
    not g732 ( n7391 , n11369 );
    not g733 ( n5088 , n1639 );
    or g734 ( n9143 , n10933 , n9823 );
    and g735 ( n13929 , n3672 , n8842 );
    nor g736 ( n9033 , n4092 , n13984 );
    or g737 ( n8173 , n1821 , n9663 );
    or g738 ( n1846 , n7156 , n1113 );
    not g739 ( n11171 , n2970 );
    or g740 ( n5834 , n1348 , n1706 );
    or g741 ( n4888 , n4544 , n3378 );
    or g742 ( n8847 , n13867 , n10061 );
    or g743 ( n8891 , n9211 , n8832 );
    not g744 ( n10280 , n5738 );
    and g745 ( n12434 , n1729 , n4087 );
    not g746 ( n5137 , n6657 );
    or g747 ( n7744 , n6344 , n12819 );
    not g748 ( n4698 , n6362 );
    or g749 ( n13079 , n10523 , n5681 );
    or g750 ( n10928 , n3047 , n8024 );
    or g751 ( n10868 , n817 , n577 );
    and g752 ( n575 , n5553 , n2968 );
    and g753 ( n3828 , n6343 , n6901 );
    not g754 ( n10276 , n2428 );
    and g755 ( n3767 , n3986 , n7260 );
    and g756 ( n8604 , n5786 , n2183 );
    nor g757 ( n12119 , n8277 , n5676 );
    and g758 ( n2095 , n12858 , n9098 );
    or g759 ( n8491 , n820 , n13302 );
    and g760 ( n285 , n4690 , n11663 );
    and g761 ( n2018 , n6625 , n3599 );
    or g762 ( n697 , n781 , n10546 );
    nor g763 ( n1432 , n1844 , n10823 );
    and g764 ( n3203 , n678 , n6453 );
    and g765 ( n5549 , n7433 , n13132 );
    nor g766 ( n6121 , n7754 , n6948 );
    or g767 ( n10829 , n1623 , n7763 );
    or g768 ( n13883 , n7122 , n8264 );
    nor g769 ( n4337 , n1628 , n13070 );
    and g770 ( n7147 , n1708 , n14323 );
    and g771 ( n4161 , n1937 , n13293 );
    and g772 ( n9949 , n10247 , n6286 );
    and g773 ( n3981 , n6486 , n798 );
    and g774 ( n6491 , n5062 , n520 );
    and g775 ( n5101 , n11803 , n14308 );
    nor g776 ( n2947 , n5986 , n1762 );
    nor g777 ( n4363 , n10179 , n11964 );
    and g778 ( n2078 , n4244 , n10404 );
    nor g779 ( n1194 , n919 , n11685 );
    and g780 ( n8698 , n1788 , n9077 );
    or g781 ( n9195 , n9541 , n7080 );
    or g782 ( n11703 , n8897 , n2083 );
    and g783 ( n326 , n55 , n11256 );
    or g784 ( n13120 , n13978 , n468 );
    or g785 ( n11742 , n12633 , n8678 );
    or g786 ( n13115 , n3219 , n8625 );
    and g787 ( n3407 , n8950 , n2954 );
    and g788 ( n4678 , n2527 , n3329 );
    or g789 ( n4072 , n14376 , n13364 );
    or g790 ( n10010 , n12023 , n2771 );
    not g791 ( n10929 , n8131 );
    and g792 ( n8165 , n14091 , n5087 );
    not g793 ( n4491 , n2470 );
    not g794 ( n7359 , n8272 );
    and g795 ( n5178 , n4871 , n11763 );
    or g796 ( n8898 , n9289 , n2825 );
    or g797 ( n2810 , n10781 , n2247 );
    and g798 ( n36 , n748 , n7950 );
    or g799 ( n3044 , n12820 , n2321 );
    or g800 ( n13764 , n12994 , n8931 );
    and g801 ( n4779 , n225 , n3205 );
    and g802 ( n9093 , n2378 , n8491 );
    or g803 ( n12090 , n12149 , n7836 );
    not g804 ( n8172 , n565 );
    and g805 ( n11555 , n13676 , n2842 );
    and g806 ( n4148 , n7970 , n4689 );
    and g807 ( n7533 , n10660 , n7087 );
    nor g808 ( n8481 , n1425 , n13400 );
    not g809 ( n11176 , n1060 );
    or g810 ( n996 , n10024 , n9421 );
    nor g811 ( n6028 , n2086 , n9785 );
    or g812 ( n8191 , n11580 , n6736 );
    and g813 ( n9568 , n3932 , n5707 );
    not g814 ( n10383 , n12687 );
    or g815 ( n3953 , n10960 , n10113 );
    nor g816 ( n2807 , n14238 , n8201 );
    and g817 ( n8054 , n6343 , n8387 );
    and g818 ( n2716 , n8692 , n12291 );
    and g819 ( n10880 , n2067 , n8472 );
    and g820 ( n6212 , n5188 , n11778 );
    or g821 ( n9168 , n791 , n9870 );
    and g822 ( n2085 , n2177 , n4459 );
    or g823 ( n9412 , n14282 , n4909 );
    and g824 ( n9741 , n14150 , n853 );
    and g825 ( n13683 , n4581 , n8731 );
    or g826 ( n7780 , n647 , n6846 );
    and g827 ( n8546 , n222 , n174 );
    and g828 ( n10684 , n14260 , n5911 );
    and g829 ( n39 , n9232 , n12134 );
    or g830 ( n6453 , n3527 , n5272 );
    and g831 ( n10421 , n5335 , n8344 );
    or g832 ( n4319 , n11379 , n1155 );
    or g833 ( n11734 , n2857 , n6526 );
    or g834 ( n3350 , n1660 , n2299 );
    nor g835 ( n11332 , n9216 , n4469 );
    and g836 ( n5578 , n432 , n464 );
    and g837 ( n13116 , n13209 , n6569 );
    and g838 ( n8708 , n8300 , n899 );
    and g839 ( n596 , n3365 , n9621 );
    or g840 ( n9906 , n10534 , n5953 );
    or g841 ( n8445 , n6781 , n9919 );
    and g842 ( n2476 , n2998 , n6973 );
    not g843 ( n4239 , n9354 );
    not g844 ( n7677 , n8168 );
    not g845 ( n11702 , n3313 );
    nor g846 ( n7439 , n10309 , n11755 );
    not g847 ( n14435 , n4939 );
    or g848 ( n10131 , n10383 , n0 );
    and g849 ( n4016 , n8232 , n6880 );
    or g850 ( n11337 , n10637 , n12356 );
    or g851 ( n8797 , n555 , n1743 );
    or g852 ( n291 , n172 , n12502 );
    and g853 ( n45 , n6609 , n9598 );
    not g854 ( n10651 , n5905 );
    and g855 ( n11042 , n10566 , n3253 );
    and g856 ( n5203 , n8801 , n5284 );
    or g857 ( n11785 , n9422 , n6465 );
    or g858 ( n1609 , n13112 , n5656 );
    nor g859 ( n13839 , n13190 , n12467 );
    or g860 ( n7483 , n14198 , n5530 );
    not g861 ( n4447 , n6586 );
    nor g862 ( n7431 , n9546 , n9203 );
    and g863 ( n14375 , n10197 , n1336 );
    and g864 ( n497 , n13745 , n2366 );
    nor g865 ( n12626 , n12311 , n491 );
    or g866 ( n8521 , n12992 , n656 );
    and g867 ( n4489 , n13342 , n6523 );
    and g868 ( n8049 , n2804 , n6640 );
    nor g869 ( n9094 , n2218 , n4664 );
    and g870 ( n5242 , n4047 , n10236 );
    or g871 ( n692 , n4123 , n10862 );
    nor g872 ( n47 , n4608 , n4507 );
    not g873 ( n251 , n14354 );
    or g874 ( n7505 , n8980 , n1942 );
    and g875 ( n1726 , n11406 , n4780 );
    not g876 ( n10650 , n8345 );
    and g877 ( n4425 , n9972 , n11029 );
    and g878 ( n6380 , n536 , n9085 );
    not g879 ( n12404 , n11547 );
    and g880 ( n10947 , n4655 , n4339 );
    not g881 ( n9745 , n3356 );
    or g882 ( n87 , n3076 , n12608 );
    nor g883 ( n8139 , n11094 , n9498 );
    or g884 ( n5766 , n9806 , n9457 );
    nor g885 ( n9519 , n11580 , n2350 );
    or g886 ( n4428 , n6891 , n943 );
    and g887 ( n9426 , n1788 , n14014 );
    or g888 ( n6681 , n12651 , n11984 );
    and g889 ( n4334 , n14465 , n3684 );
    and g890 ( n7064 , n5980 , n7077 );
    or g891 ( n3184 , n4602 , n7316 );
    and g892 ( n3189 , n2961 , n11522 );
    nor g893 ( n9675 , n13248 , n5714 );
    and g894 ( n1164 , n13421 , n10227 );
    not g895 ( n400 , n7652 );
    and g896 ( n1782 , n2758 , n10442 );
    or g897 ( n8782 , n1628 , n11242 );
    and g898 ( n11407 , n1857 , n9828 );
    and g899 ( n2475 , n3762 , n4067 );
    not g900 ( n9245 , n13231 );
    or g901 ( n11072 , n10871 , n7854 );
    or g902 ( n10404 , n10449 , n10365 );
    or g903 ( n9175 , n1840 , n1721 );
    not g904 ( n9403 , n7064 );
    or g905 ( n6623 , n12968 , n9256 );
    nor g906 ( n11432 , n10977 , n11802 );
    not g907 ( n6933 , n9377 );
    nor g908 ( n5883 , n13981 , n2122 );
    or g909 ( n2404 , n4562 , n4032 );
    and g910 ( n1497 , n7768 , n12908 );
    nor g911 ( n1486 , n6039 , n11926 );
    and g912 ( n8936 , n9191 , n12350 );
    and g913 ( n10144 , n10197 , n2993 );
    or g914 ( n8273 , n12494 , n4122 );
    nor g915 ( n7170 , n329 , n6172 );
    nor g916 ( n6403 , n1617 , n2879 );
    or g917 ( n1276 , n12934 , n1467 );
    not g918 ( n8692 , n4824 );
    or g919 ( n8255 , n1535 , n3240 );
    not g920 ( n7662 , n4835 );
    or g921 ( n10293 , n227 , n3081 );
    nor g922 ( n7985 , n300 , n11246 );
    and g923 ( n10833 , n12147 , n2840 );
    not g924 ( n11838 , n8451 );
    and g925 ( n2618 , n10458 , n13245 );
    or g926 ( n12707 , n4340 , n14131 );
    or g927 ( n4168 , n7888 , n8514 );
    or g928 ( n4474 , n3093 , n2144 );
    or g929 ( n6961 , n11953 , n12125 );
    or g930 ( n2662 , n6544 , n2808 );
    or g931 ( n10670 , n12414 , n5877 );
    nor g932 ( n1682 , n4877 , n701 );
    or g933 ( n9833 , n8986 , n9240 );
    and g934 ( n11207 , n706 , n277 );
    or g935 ( n13014 , n1711 , n8010 );
    or g936 ( n12083 , n1602 , n13504 );
    not g937 ( n11620 , n4465 );
    nor g938 ( n9192 , n7720 , n5982 );
    and g939 ( n4815 , n7068 , n10983 );
    and g940 ( n10787 , n5975 , n987 );
    or g941 ( n10639 , n619 , n5051 );
    not g942 ( n1708 , n7052 );
    nor g943 ( n8534 , n8015 , n11434 );
    or g944 ( n13838 , n13706 , n4025 );
    or g945 ( n10954 , n769 , n27 );
    or g946 ( n6678 , n4092 , n699 );
    nor g947 ( n14080 , n10715 , n5075 );
    and g948 ( n8933 , n6157 , n6468 );
    or g949 ( n1438 , n4822 , n683 );
    and g950 ( n14340 , n13676 , n12686 );
    not g951 ( n5450 , n630 );
    and g952 ( n12634 , n13367 , n12223 );
    not g953 ( n8216 , n8750 );
    or g954 ( n715 , n1391 , n1408 );
    and g955 ( n7256 , n13227 , n1590 );
    and g956 ( n11423 , n14227 , n10771 );
    not g957 ( n10617 , n1178 );
    not g958 ( n6971 , n2918 );
    or g959 ( n7055 , n5406 , n9370 );
    not g960 ( n3309 , n6308 );
    and g961 ( n8077 , n6051 , n3399 );
    and g962 ( n1314 , n5279 , n13077 );
    or g963 ( n13198 , n3667 , n8265 );
    not g964 ( n3034 , n1161 );
    and g965 ( n5679 , n12521 , n3938 );
    and g966 ( n6626 , n7060 , n4031 );
    or g967 ( n7478 , n6654 , n10252 );
    and g968 ( n13752 , n11852 , n9142 );
    or g969 ( n6503 , n1198 , n758 );
    and g970 ( n3803 , n13626 , n6104 );
    nor g971 ( n9408 , n8825 , n9901 );
    or g972 ( n2560 , n2055 , n6882 );
    and g973 ( n7563 , n3813 , n12744 );
    nor g974 ( n4944 , n10189 , n1777 );
    not g975 ( n9952 , n14011 );
    or g976 ( n6862 , n5493 , n2722 );
    or g977 ( n6338 , n7971 , n14423 );
    or g978 ( n9221 , n1538 , n6769 );
    or g979 ( n7932 , n10731 , n7361 );
    and g980 ( n767 , n12404 , n13157 );
    and g981 ( n4381 , n8147 , n9682 );
    and g982 ( n2538 , n1489 , n444 );
    and g983 ( n7414 , n6754 , n1244 );
    or g984 ( n10563 , n3445 , n4997 );
    and g985 ( n3223 , n4932 , n1052 );
    and g986 ( n12883 , n5948 , n7213 );
    or g987 ( n3023 , n10245 , n2634 );
    or g988 ( n2211 , n1821 , n6976 );
    nor g989 ( n12891 , n4270 , n1790 );
    and g990 ( n13613 , n6507 , n3425 );
    and g991 ( n12895 , n4102 , n11604 );
    and g992 ( n3522 , n5940 , n10429 );
    or g993 ( n13789 , n8980 , n9883 );
    or g994 ( n1005 , n5715 , n2777 );
    nor g995 ( n8643 , n31 , n9253 );
    and g996 ( n5799 , n11674 , n1296 );
    or g997 ( n10053 , n11620 , n6204 );
    or g998 ( n5393 , n1728 , n8587 );
    and g999 ( n7460 , n2820 , n5900 );
    or g1000 ( n8887 , n9589 , n11404 );
    nor g1001 ( n8466 , n7919 , n9150 );
    or g1002 ( n915 , n1202 , n8919 );
    and g1003 ( n6545 , n6316 , n4116 );
    not g1004 ( n14006 , n4615 );
    or g1005 ( n3995 , n12764 , n127 );
    and g1006 ( n11733 , n4102 , n13019 );
    and g1007 ( n12512 , n10457 , n10964 );
    or g1008 ( n6959 , n7700 , n11053 );
    or g1009 ( n13059 , n8714 , n11586 );
    or g1010 ( n8042 , n6706 , n11370 );
    nor g1011 ( n3145 , n3443 , n3581 );
    or g1012 ( n9165 , n954 , n9515 );
    and g1013 ( n3498 , n7779 , n3793 );
    or g1014 ( n4044 , n13142 , n10616 );
    and g1015 ( n7469 , n6486 , n5274 );
    or g1016 ( n3832 , n1613 , n10027 );
    and g1017 ( n9930 , n4690 , n14082 );
    not g1018 ( n13003 , n11120 );
    and g1019 ( n5733 , n10822 , n9561 );
    and g1020 ( n3242 , n6147 , n685 );
    and g1021 ( n4850 , n12741 , n13731 );
    and g1022 ( n10194 , n286 , n2439 );
    nor g1023 ( n6419 , n7375 , n5611 );
    not g1024 ( n3405 , n1911 );
    and g1025 ( n2654 , n6744 , n10474 );
    nor g1026 ( n10344 , n11285 , n7555 );
    or g1027 ( n6169 , n14466 , n8089 );
    and g1028 ( n3854 , n3799 , n10776 );
    not g1029 ( n390 , n10204 );
    not g1030 ( n10089 , n6123 );
    not g1031 ( n8969 , n1894 );
    and g1032 ( n388 , n3586 , n4170 );
    not g1033 ( n1728 , n2484 );
    and g1034 ( n4948 , n4276 , n14148 );
    and g1035 ( n3829 , n13367 , n9540 );
    and g1036 ( n10008 , n6354 , n6814 );
    nor g1037 ( n3677 , n12288 , n731 );
    and g1038 ( n13606 , n3536 , n13928 );
    or g1039 ( n4894 , n12391 , n8550 );
    and g1040 ( n10075 , n12461 , n2737 );
    or g1041 ( n7565 , n2878 , n6355 );
    or g1042 ( n12384 , n4913 , n6231 );
    and g1043 ( n1399 , n8386 , n8194 );
    and g1044 ( n4256 , n4614 , n8039 );
    nor g1045 ( n13353 , n1417 , n4730 );
    and g1046 ( n885 , n5634 , n2524 );
    or g1047 ( n5111 , n13083 , n13478 );
    or g1048 ( n10445 , n11935 , n6152 );
    or g1049 ( n11786 , n5732 , n8845 );
    and g1050 ( n4364 , n2322 , n8772 );
    and g1051 ( n12822 , n8372 , n13692 );
    and g1052 ( n1745 , n8386 , n275 );
    and g1053 ( n7107 , n5229 , n1134 );
    and g1054 ( n9171 , n11329 , n2348 );
    or g1055 ( n13396 , n13978 , n9649 );
    or g1056 ( n8713 , n8747 , n5968 );
    nor g1057 ( n4086 , n12568 , n5323 );
    and g1058 ( n12385 , n8238 , n1396 );
    or g1059 ( n8690 , n10857 , n9693 );
    or g1060 ( n2872 , n1051 , n4706 );
    and g1061 ( n1952 , n13535 , n8340 );
    or g1062 ( n689 , n1031 , n8785 );
    or g1063 ( n8574 , n8209 , n13688 );
    not g1064 ( n9824 , n4050 );
    nor g1065 ( n4916 , n8543 , n2483 );
    nor g1066 ( n6736 , n9176 , n244 );
    and g1067 ( n1369 , n8855 , n12094 );
    nor g1068 ( n13387 , n8223 , n3413 );
    not g1069 ( n1354 , n442 );
    nor g1070 ( n4917 , n11584 , n4763 );
    or g1071 ( n8998 , n5891 , n8128 );
    and g1072 ( n9886 , n7057 , n7498 );
    not g1073 ( n5429 , n13765 );
    and g1074 ( n1866 , n3332 , n5776 );
    and g1075 ( n2668 , n2445 , n13348 );
    not g1076 ( n4639 , n7518 );
    or g1077 ( n13897 , n8748 , n2376 );
    and g1078 ( n1551 , n2465 , n35 );
    not g1079 ( n5483 , n12249 );
    not g1080 ( n13240 , n2744 );
    not g1081 ( n1255 , n13154 );
    or g1082 ( n9217 , n7481 , n1896 );
    not g1083 ( n820 , n13901 );
    and g1084 ( n12720 , n13078 , n353 );
    nor g1085 ( n6070 , n8378 , n13377 );
    and g1086 ( n8761 , n2961 , n11389 );
    or g1087 ( n12556 , n4925 , n6056 );
    or g1088 ( n12767 , n172 , n2059 );
    or g1089 ( n953 , n9422 , n11081 );
    not g1090 ( n9035 , n8595 );
    and g1091 ( n1505 , n1414 , n12484 );
    or g1092 ( n6950 , n14449 , n11649 );
    and g1093 ( n1545 , n4117 , n9840 );
    not g1094 ( n3211 , n4533 );
    or g1095 ( n12239 , n12211 , n8522 );
    or g1096 ( n3669 , n13016 , n6825 );
    or g1097 ( n2513 , n12112 , n8621 );
    and g1098 ( n8067 , n5088 , n10411 );
    or g1099 ( n5881 , n9353 , n12845 );
    or g1100 ( n1892 , n12712 , n3750 );
    or g1101 ( n13610 , n7971 , n11560 );
    or g1102 ( n12108 , n194 , n4552 );
    and g1103 ( n5386 , n7670 , n1504 );
    and g1104 ( n13802 , n7429 , n1523 );
    or g1105 ( n12213 , n9140 , n13741 );
    and g1106 ( n3519 , n5825 , n4762 );
    nor g1107 ( n8467 , n9035 , n1869 );
    or g1108 ( n422 , n791 , n12817 );
    or g1109 ( n1557 , n6556 , n10736 );
    or g1110 ( n1590 , n100 , n869 );
    and g1111 ( n5602 , n5279 , n10860 );
    and g1112 ( n12276 , n11142 , n8062 );
    or g1113 ( n13510 , n838 , n10194 );
    or g1114 ( n3650 , n3076 , n12359 );
    and g1115 ( n8379 , n10134 , n2754 );
    nor g1116 ( n7555 , n1218 , n3302 );
    not g1117 ( n11129 , n2094 );
    or g1118 ( n7268 , n13978 , n3695 );
    or g1119 ( n12981 , n3120 , n4288 );
    nor g1120 ( n3225 , n13310 , n6513 );
    not g1121 ( n772 , n12323 );
    or g1122 ( n2964 , n6607 , n6985 );
    nor g1123 ( n8880 , n4195 , n12275 );
    nor g1124 ( n1234 , n4988 , n6403 );
    or g1125 ( n1038 , n3125 , n138 );
    and g1126 ( n8455 , n1414 , n5740 );
    and g1127 ( n2353 , n10084 , n6398 );
    or g1128 ( n9343 , n13847 , n9279 );
    not g1129 ( n2417 , n6451 );
    and g1130 ( n10222 , n13626 , n8946 );
    and g1131 ( n8909 , n9589 , n1196 );
    and g1132 ( n1861 , n7997 , n7925 );
    or g1133 ( n2955 , n7364 , n9283 );
    or g1134 ( n4232 , n791 , n10116 );
    nor g1135 ( n14352 , n10803 , n14019 );
    and g1136 ( n10437 , n3942 , n6958 );
    or g1137 ( n866 , n234 , n1439 );
    not g1138 ( n3290 , n1312 );
    or g1139 ( n13685 , n2089 , n11471 );
    or g1140 ( n3074 , n11542 , n2285 );
    not g1141 ( n8701 , n2484 );
    or g1142 ( n8837 , n8881 , n7544 );
    and g1143 ( n6786 , n11875 , n4247 );
    nor g1144 ( n3890 , n12294 , n10002 );
    nor g1145 ( n2768 , n8462 , n12454 );
    and g1146 ( n6247 , n4104 , n3687 );
    and g1147 ( n5927 , n12953 , n14189 );
    or g1148 ( n2896 , n7011 , n8418 );
    and g1149 ( n4336 , n6016 , n8675 );
    or g1150 ( n6552 , n8983 , n5205 );
    or g1151 ( n12972 , n412 , n10132 );
    or g1152 ( n13291 , n12019 , n2582 );
    nor g1153 ( n2122 , n4561 , n7879 );
    nor g1154 ( n11044 , n13276 , n12539 );
    or g1155 ( n12476 , n7812 , n10430 );
    or g1156 ( n14424 , n7530 , n10986 );
    nor g1157 ( n12681 , n11047 , n10390 );
    nor g1158 ( n6325 , n9414 , n14236 );
    and g1159 ( n5433 , n1804 , n3149 );
    nor g1160 ( n3638 , n425 , n4301 );
    and g1161 ( n1754 , n5825 , n4021 );
    and g1162 ( n7155 , n2021 , n1211 );
    and g1163 ( n8735 , n14016 , n4963 );
    and g1164 ( n2220 , n1610 , n8973 );
    and g1165 ( n13788 , n2445 , n4878 );
    and g1166 ( n10944 , n11950 , n1856 );
    or g1167 ( n8723 , n5695 , n6033 );
    and g1168 ( n12619 , n5062 , n11386 );
    and g1169 ( n9916 , n7284 , n1566 );
    or g1170 ( n2124 , n3088 , n12381 );
    or g1171 ( n11720 , n11097 , n4401 );
    or g1172 ( n6547 , n492 , n12374 );
    or g1173 ( n13767 , n4052 , n12059 );
    or g1174 ( n13506 , n7803 , n3328 );
    or g1175 ( n12967 , n12292 , n9030 );
    and g1176 ( n274 , n12018 , n2553 );
    or g1177 ( n5910 , n3099 , n743 );
    or g1178 ( n9261 , n12428 , n9013 );
    and g1179 ( n8813 , n692 , n8349 );
    or g1180 ( n14386 , n5409 , n589 );
    nor g1181 ( n1953 , n14370 , n11767 );
    not g1182 ( n11569 , n11547 );
    nor g1183 ( n3906 , n7364 , n14052 );
    and g1184 ( n3513 , n13362 , n1828 );
    and g1185 ( n5205 , n11142 , n10669 );
    not g1186 ( n13937 , n11574 );
    nor g1187 ( n9432 , n8197 , n6864 );
    not g1188 ( n9280 , n10765 );
    nor g1189 ( n330 , n10402 , n14070 );
    and g1190 ( n8227 , n9972 , n3636 );
    or g1191 ( n4796 , n11171 , n5422 );
    or g1192 ( n4310 , n11621 , n8317 );
    or g1193 ( n2687 , n2790 , n7093 );
    nor g1194 ( n9634 , n9550 , n12111 );
    not g1195 ( n1701 , n10775 );
    or g1196 ( n12137 , n12023 , n3563 );
    nor g1197 ( n4575 , n6672 , n12988 );
    or g1198 ( n5052 , n13806 , n4513 );
    and g1199 ( n4329 , n200 , n14509 );
    or g1200 ( n4940 , n2272 , n13534 );
    nor g1201 ( n7094 , n13050 , n10959 );
    and g1202 ( n3624 , n8047 , n479 );
    or g1203 ( n12462 , n10781 , n1456 );
    and g1204 ( n3326 , n11422 , n3555 );
    or g1205 ( n13250 , n5362 , n11349 );
    and g1206 ( n12053 , n2783 , n8889 );
    or g1207 ( n6692 , n4498 , n11645 );
    and g1208 ( n13541 , n14260 , n3001 );
    or g1209 ( n4459 , n5064 , n2167 );
    or g1210 ( n5029 , n14200 , n9026 );
    not g1211 ( n7211 , n2432 );
    and g1212 ( n10633 , n7187 , n1737 );
    and g1213 ( n3360 , n12449 , n6347 );
    or g1214 ( n3679 , n9541 , n3407 );
    and g1215 ( n13567 , n7419 , n8764 );
    or g1216 ( n6685 , n7914 , n6597 );
    or g1217 ( n2815 , n100 , n14441 );
    or g1218 ( n2342 , n11572 , n12574 );
    or g1219 ( n3974 , n8983 , n1288 );
    or g1220 ( n8383 , n8452 , n4712 );
    and g1221 ( n7324 , n13147 , n4625 );
    nor g1222 ( n13753 , n9806 , n14297 );
    or g1223 ( n11527 , n4205 , n12916 );
    and g1224 ( n8626 , n10516 , n110 );
    or g1225 ( n9449 , n4205 , n3291 );
    nor g1226 ( n11928 , n8209 , n7160 );
    and g1227 ( n13047 , n7618 , n1959 );
    and g1228 ( n14518 , n9509 , n6662 );
    not g1229 ( n2422 , n13447 );
    or g1230 ( n7497 , n1189 , n7821 );
    or g1231 ( n3091 , n5936 , n4569 );
    or g1232 ( n12896 , n4033 , n9310 );
    and g1233 ( n1751 , n776 , n12392 );
    and g1234 ( n52 , n14038 , n2379 );
    not g1235 ( n6090 , n12394 );
    or g1236 ( n7384 , n10637 , n14344 );
    not g1237 ( n264 , n9388 );
    and g1238 ( n4169 , n6537 , n13858 );
    or g1239 ( n9937 , n6206 , n13647 );
    and g1240 ( n13795 , n14213 , n13256 );
    or g1241 ( n256 , n6323 , n5027 );
    and g1242 ( n1151 , n1431 , n3122 );
    and g1243 ( n13719 , n3286 , n10049 );
    nor g1244 ( n1858 , n13941 , n9820 );
    not g1245 ( n12018 , n7621 );
    and g1246 ( n7761 , n13464 , n14451 );
    or g1247 ( n2963 , n7963 , n4147 );
    or g1248 ( n11592 , n6654 , n13161 );
    or g1249 ( n12470 , n2412 , n9259 );
    not g1250 ( n13338 , n9865 );
    nor g1251 ( n1019 , n1685 , n10065 );
    and g1252 ( n11416 , n8630 , n8362 );
    and g1253 ( n544 , n3097 , n13666 );
    not g1254 ( n2548 , n3822 );
    or g1255 ( n4432 , n7122 , n12514 );
    and g1256 ( n11211 , n13359 , n12742 );
    or g1257 ( n10412 , n3667 , n693 );
    not g1258 ( n11392 , n13186 );
    and g1259 ( n7040 , n14351 , n11907 );
    and g1260 ( n6029 , n10854 , n3574 );
    and g1261 ( n5074 , n11213 , n8314 );
    or g1262 ( n7671 , n12020 , n11825 );
    and g1263 ( n9348 , n7079 , n12080 );
    not g1264 ( n6062 , n10897 );
    or g1265 ( n9556 , n1202 , n5767 );
    or g1266 ( n5451 , n194 , n6269 );
    or g1267 ( n4626 , n2098 , n7164 );
    or g1268 ( n6962 , n11839 , n1072 );
    or g1269 ( n6770 , n4128 , n13493 );
    and g1270 ( n10986 , n12521 , n8987 );
    and g1271 ( n7951 , n2985 , n1135 );
    nor g1272 ( n2443 , n6424 , n1055 );
    not g1273 ( n2465 , n6905 );
    and g1274 ( n5166 , n8721 , n6984 );
    or g1275 ( n13392 , n5625 , n7374 );
    nor g1276 ( n2610 , n13875 , n206 );
    not g1277 ( n5460 , n834 );
    and g1278 ( n2616 , n7852 , n1236 );
    and g1279 ( n5755 , n8786 , n12221 );
    and g1280 ( n13820 , n9571 , n9603 );
    and g1281 ( n1674 , n6157 , n11521 );
    and g1282 ( n11185 , n6013 , n5667 );
    and g1283 ( n7039 , n5459 , n9438 );
    and g1284 ( n7680 , n6830 , n3698 );
    or g1285 ( n2984 , n12601 , n4943 );
    or g1286 ( n4776 , n12821 , n8627 );
    not g1287 ( n2012 , n12976 );
    not g1288 ( n3161 , n9959 );
    and g1289 ( n12067 , n11867 , n13618 );
    and g1290 ( n13565 , n3401 , n12488 );
    or g1291 ( n11754 , n10713 , n10145 );
    or g1292 ( n11249 , n480 , n4198 );
    nor g1293 ( n11929 , n4092 , n9207 );
    and g1294 ( n6265 , n11093 , n7332 );
    or g1295 ( n7672 , n10449 , n10553 );
    and g1296 ( n5818 , n2367 , n9391 );
    and g1297 ( n10643 , n6525 , n10435 );
    not g1298 ( n8112 , n13109 );
    or g1299 ( n2174 , n4741 , n10114 );
    and g1300 ( n1461 , n8605 , n6815 );
    and g1301 ( n7417 , n5240 , n7189 );
    or g1302 ( n6011 , n3799 , n8746 );
    nor g1303 ( n6889 , n600 , n2646 );
    or g1304 ( n14205 , n9174 , n8988 );
    or g1305 ( n7839 , n8304 , n2151 );
    or g1306 ( n9621 , n12149 , n5060 );
    and g1307 ( n3919 , n13755 , n5372 );
    and g1308 ( n9074 , n11484 , n5993 );
    and g1309 ( n935 , n12147 , n9247 );
    or g1310 ( n7706 , n14366 , n9715 );
    and g1311 ( n8124 , n9154 , n8991 );
    and g1312 ( n11144 , n5434 , n9146 );
    not g1313 ( n11548 , n11324 );
    and g1314 ( n7539 , n8020 , n7303 );
    not g1315 ( n6211 , n12086 );
    or g1316 ( n4075 , n9269 , n2372 );
    not g1317 ( n3709 , n6054 );
    or g1318 ( n342 , n3546 , n10071 );
    not g1319 ( n14388 , n11474 );
    or g1320 ( n4571 , n1044 , n447 );
    and g1321 ( n4809 , n11240 , n12237 );
    or g1322 ( n1525 , n5587 , n232 );
    and g1323 ( n6902 , n1678 , n3392 );
    not g1324 ( n4898 , n10985 );
    and g1325 ( n2007 , n687 , n7286 );
    not g1326 ( n931 , n2355 );
    nor g1327 ( n14017 , n5429 , n4409 );
    and g1328 ( n9355 , n6957 , n7975 );
    and g1329 ( n2771 , n12592 , n12554 );
    and g1330 ( n7992 , n2564 , n2931 );
    and g1331 ( n7864 , n12265 , n125 );
    not g1332 ( n4091 , n8288 );
    and g1333 ( n8410 , n986 , n5295 );
    and g1334 ( n1951 , n10050 , n11088 );
    nor g1335 ( n6278 , n10136 , n10041 );
    nor g1336 ( n11757 , n4518 , n220 );
    or g1337 ( n2307 , n9856 , n3522 );
    or g1338 ( n10795 , n9403 , n2905 );
    and g1339 ( n12649 , n10710 , n2793 );
    nor g1340 ( n3990 , n8458 , n2990 );
    or g1341 ( n11887 , n6629 , n8839 );
    and g1342 ( n668 , n13362 , n4488 );
    and g1343 ( n5851 , n13944 , n4183 );
    nor g1344 ( n11050 , n9423 , n2010 );
    or g1345 ( n4452 , n3394 , n6608 );
    and g1346 ( n14089 , n7221 , n161 );
    and g1347 ( n982 , n4619 , n12723 );
    and g1348 ( n7623 , n11336 , n4073 );
    or g1349 ( n3665 , n11510 , n10251 );
    and g1350 ( n13558 , n13860 , n4452 );
    nor g1351 ( n9590 , n10036 , n9309 );
    not g1352 ( n9953 , n8650 );
    or g1353 ( n13191 , n2784 , n2701 );
    or g1354 ( n7845 , n9864 , n1237 );
    nor g1355 ( n2115 , n4284 , n11916 );
    nor g1356 ( n8929 , n1760 , n5208 );
    nor g1357 ( n11562 , n48 , n3894 );
    or g1358 ( n13091 , n815 , n10615 );
    or g1359 ( n10487 , n8452 , n10070 );
    or g1360 ( n7137 , n12149 , n1994 );
    and g1361 ( n3556 , n6898 , n8687 );
    and g1362 ( n3810 , n9191 , n4229 );
    not g1363 ( n3365 , n1571 );
    nor g1364 ( n13829 , n900 , n12706 );
    not g1365 ( n235 , n11901 );
    not g1366 ( n8242 , n7339 );
    or g1367 ( n10939 , n2387 , n9958 );
    and g1368 ( n4078 , n9297 , n8659 );
    not g1369 ( n12449 , n8524 );
    and g1370 ( n5342 , n1904 , n10146 );
    and g1371 ( n9717 , n6873 , n1241 );
    nor g1372 ( n8720 , n13327 , n9799 );
    and g1373 ( n4521 , n428 , n1038 );
    and g1374 ( n654 , n2533 , n9165 );
    or g1375 ( n2785 , n11121 , n4920 );
    nor g1376 ( n5100 , n163 , n8590 );
    not g1377 ( n1850 , n4175 );
    and g1378 ( n13647 , n7203 , n10543 );
    and g1379 ( n5307 , n12445 , n2124 );
    not g1380 ( n6544 , n2609 );
    not g1381 ( n13806 , n7086 );
    and g1382 ( n11374 , n4581 , n2887 );
    or g1383 ( n6901 , n11909 , n7103 );
    and g1384 ( n12731 , n12986 , n7449 );
    not g1385 ( n12592 , n1724 );
    and g1386 ( n13314 , n11300 , n12289 );
    nor g1387 ( n11000 , n2780 , n12654 );
    or g1388 ( n3122 , n648 , n4628 );
    not g1389 ( n4803 , n9416 );
    and g1390 ( n13574 , n8111 , n4460 );
    not g1391 ( n1023 , n3054 );
    not g1392 ( n10619 , n9543 );
    and g1393 ( n7854 , n11636 , n5829 );
    or g1394 ( n1131 , n766 , n2464 );
    not g1395 ( n5229 , n9450 );
    and g1396 ( n9891 , n8630 , n1570 );
    not g1397 ( n4634 , n7200 );
    or g1398 ( n92 , n4239 , n5802 );
    and g1399 ( n5801 , n3724 , n5931 );
    and g1400 ( n557 , n986 , n7078 );
    not g1401 ( n2983 , n13734 );
    and g1402 ( n7317 , n4244 , n1750 );
    or g1403 ( n9975 , n7358 , n13649 );
    and g1404 ( n13812 , n3923 , n9424 );
    or g1405 ( n6468 , n11951 , n7385 );
    and g1406 ( n13693 , n74 , n7669 );
    and g1407 ( n13234 , n11066 , n4510 );
    or g1408 ( n994 , n12324 , n1918 );
    or g1409 ( n2532 , n4898 , n10437 );
    or g1410 ( n8710 , n14110 , n7482 );
    and g1411 ( n8648 , n7057 , n13886 );
    or g1412 ( n12830 , n10781 , n13262 );
    or g1413 ( n8764 , n77 , n2476 );
    or g1414 ( n11222 , n8527 , n13322 );
    or g1415 ( n3398 , n4045 , n1369 );
    or g1416 ( n3013 , n13016 , n7199 );
    or g1417 ( n1208 , n13806 , n4833 );
    and g1418 ( n4053 , n7208 , n13150 );
    or g1419 ( n1424 , n13875 , n12067 );
    and g1420 ( n8705 , n6527 , n7396 );
    and g1421 ( n5588 , n8965 , n4220 );
    or g1422 ( n8348 , n5575 , n13782 );
    and g1423 ( n4662 , n5053 , n8803 );
    or g1424 ( n6294 , n5315 , n12778 );
    or g1425 ( n11716 , n12019 , n7369 );
    or g1426 ( n7110 , n1538 , n6626 );
    or g1427 ( n13452 , n555 , n10744 );
    and g1428 ( n8303 , n9297 , n4872 );
    not g1429 ( n6389 , n5990 );
    and g1430 ( n14129 , n1937 , n12393 );
    or g1431 ( n12818 , n11420 , n2633 );
    nor g1432 ( n12508 , n3944 , n2052 );
    and g1433 ( n3605 , n200 , n11298 );
    or g1434 ( n3664 , n820 , n4660 );
    and g1435 ( n3456 , n11220 , n10126 );
    and g1436 ( n2325 , n13781 , n2260 );
    or g1437 ( n4537 , n2843 , n1364 );
    not g1438 ( n1538 , n777 );
    not g1439 ( n6537 , n3775 );
    or g1440 ( n9912 , n387 , n9517 );
    and g1441 ( n11783 , n6822 , n11229 );
    and g1442 ( n11532 , n12858 , n7694 );
    or g1443 ( n5212 , n2098 , n2749 );
    or g1444 ( n4116 , n9429 , n14359 );
    or g1445 ( n1387 , n12601 , n3157 );
    and g1446 ( n5235 , n3536 , n13335 );
    and g1447 ( n6483 , n5275 , n10993 );
    and g1448 ( n11645 , n8025 , n11890 );
    not g1449 ( n2564 , n12503 );
    nor g1450 ( n12761 , n3165 , n4912 );
    or g1451 ( n10703 , n6595 , n14482 );
    and g1452 ( n14396 , n10072 , n7051 );
    nor g1453 ( n2917 , n1914 , n2113 );
    or g1454 ( n1597 , n2025 , n1624 );
    not g1455 ( n5839 , n10837 );
    nor g1456 ( n6972 , n7227 , n10938 );
    or g1457 ( n8012 , n3011 , n11064 );
    and g1458 ( n2922 , n7419 , n13691 );
    not g1459 ( n4065 , n2934 );
    and g1460 ( n255 , n1117 , n9072 );
    not g1461 ( n7768 , n1955 );
    and g1462 ( n8322 , n13252 , n1181 );
    not g1463 ( n7624 , n13476 );
    not g1464 ( n4572 , n11582 );
    or g1465 ( n5124 , n6857 , n3883 );
    not g1466 ( n12159 , n448 );
    not g1467 ( n6781 , n3681 );
    or g1468 ( n2428 , n12025 , n3673 );
    and g1469 ( n7471 , n13404 , n847 );
    and g1470 ( n5524 , n10357 , n9195 );
    or g1471 ( n10267 , n8332 , n7960 );
    or g1472 ( n11849 , n317 , n9576 );
    and g1473 ( n2083 , n11093 , n10163 );
    and g1474 ( n10252 , n1489 , n11137 );
    not g1475 ( n11558 , n8813 );
    and g1476 ( n2736 , n13860 , n8779 );
    and g1477 ( n1388 , n6556 , n8795 );
    or g1478 ( n4421 , n5762 , n12882 );
    not g1479 ( n7963 , n6251 );
    and g1480 ( n12365 , n2942 , n3903 );
    or g1481 ( n6414 , n5997 , n12638 );
    or g1482 ( n5309 , n7678 , n12570 );
    not g1483 ( n6519 , n7086 );
    and g1484 ( n12665 , n12802 , n9906 );
    or g1485 ( n12289 , n3168 , n721 );
    and g1486 ( n2939 , n225 , n9356 );
    or g1487 ( n11284 , n2181 , n8308 );
    not g1488 ( n5999 , n3361 );
    and g1489 ( n617 , n8697 , n14094 );
    not g1490 ( n4589 , n6855 );
    or g1491 ( n2252 , n2908 , n2391 );
    and g1492 ( n4720 , n7710 , n12886 );
    or g1493 ( n9915 , n4357 , n2447 );
    or g1494 ( n10385 , n4739 , n14469 );
    not g1495 ( n11251 , n1932 );
    nor g1496 ( n1042 , n11714 , n2611 );
    and g1497 ( n4160 , n10302 , n9374 );
    or g1498 ( n10213 , n9174 , n4643 );
    not g1499 ( n3210 , n10314 );
    not g1500 ( n9792 , n11158 );
    not g1501 ( n13516 , n5242 );
    not g1502 ( n13525 , n6787 );
    or g1503 ( n3138 , n9289 , n13620 );
    or g1504 ( n8505 , n11440 , n14265 );
    nor g1505 ( n592 , n3132 , n2703 );
    nor g1506 ( n2199 , n12968 , n8276 );
    not g1507 ( n9718 , n13429 );
    and g1508 ( n5186 , n5857 , n672 );
    not g1509 ( n7116 , n2970 );
    and g1510 ( n4513 , n3724 , n11957 );
    and g1511 ( n1603 , n327 , n3152 );
    and g1512 ( n5213 , n12542 , n13329 );
    nor g1513 ( n11755 , n13324 , n10308 );
    and g1514 ( n6063 , n4790 , n2966 );
    or g1515 ( n7488 , n4233 , n9178 );
    or g1516 ( n8915 , n5562 , n5474 );
    and g1517 ( n10676 , n8769 , n8509 );
    and g1518 ( n9386 , n12953 , n193 );
    nor g1519 ( n11945 , n473 , n933 );
    not g1520 ( n13720 , n6460 );
    and g1521 ( n6738 , n2583 , n1491 );
    nor g1522 ( n8999 , n1820 , n14352 );
    and g1523 ( n2622 , n11470 , n5652 );
    nor g1524 ( n5916 , n5919 , n9787 );
    or g1525 ( n947 , n8877 , n3654 );
    not g1526 ( n3400 , n13084 );
    or g1527 ( n7074 , n2694 , n13152 );
    nor g1528 ( n11184 , n1681 , n9205 );
    or g1529 ( n571 , n1028 , n5970 );
    or g1530 ( n503 , n4925 , n10366 );
    or g1531 ( n9055 , n10351 , n10598 );
    and g1532 ( n3323 , n4880 , n4640 );
    or g1533 ( n8331 , n7678 , n1592 );
    not g1534 ( n11584 , n12358 );
    not g1535 ( n11262 , n9252 );
    or g1536 ( n6779 , n1198 , n10007 );
    or g1537 ( n4290 , n9226 , n9712 );
    not g1538 ( n12079 , n513 );
    not g1539 ( n12335 , n12970 );
    not g1540 ( n584 , n11788 );
    not g1541 ( n11572 , n7064 );
    or g1542 ( n4941 , n7229 , n3721 );
    and g1543 ( n14259 , n225 , n12690 );
    and g1544 ( n6978 , n10384 , n5905 );
    or g1545 ( n6892 , n10062 , n10093 );
    nor g1546 ( n3963 , n9046 , n7714 );
    not g1547 ( n3530 , n10012 );
    and g1548 ( n3544 , n8376 , n2854 );
    and g1549 ( n9135 , n7221 , n11974 );
    or g1550 ( n12524 , n13854 , n8054 );
    and g1551 ( n14427 , n5926 , n6633 );
    not g1552 ( n882 , n3054 );
    or g1553 ( n5829 , n4807 , n12150 );
    not g1554 ( n3097 , n5613 );
    and g1555 ( n9062 , n12445 , n12297 );
    or g1556 ( n1410 , n10019 , n96 );
    not g1557 ( n12712 , n7600 );
    not g1558 ( n12622 , n11541 );
    or g1559 ( n6528 , n1189 , n7733 );
    and g1560 ( n5381 , n222 , n757 );
    or g1561 ( n10983 , n12622 , n14037 );
    or g1562 ( n5721 , n5409 , n6539 );
    and g1563 ( n2228 , n7429 , n9001 );
    or g1564 ( n14439 , n1711 , n4138 );
    or g1565 ( n9331 , n6090 , n11758 );
    or g1566 ( n2977 , n10019 , n11517 );
    or g1567 ( n5416 , n5855 , n4907 );
    not g1568 ( n12167 , n3833 );
    or g1569 ( n6796 , n3093 , n8239 );
    or g1570 ( n2711 , n329 , n7991 );
    and g1571 ( n7760 , n5489 , n8886 );
    not g1572 ( n1152 , n4769 );
    or g1573 ( n4141 , n3569 , n19 );
    nor g1574 ( n10271 , n6765 , n2323 );
    not g1575 ( n11121 , n14412 );
    and g1576 ( n107 , n6311 , n280 );
    and g1577 ( n5843 , n9345 , n135 );
    or g1578 ( n3005 , n4207 , n10869 );
    and g1579 ( n279 , n10815 , n4038 );
    not g1580 ( n3942 , n3440 );
    or g1581 ( n8187 , n13016 , n10371 );
    and g1582 ( n5708 , n12858 , n7114 );
    or g1583 ( n790 , n2318 , n10941 );
    or g1584 ( n4667 , n8034 , n10477 );
    or g1585 ( n4578 , n11105 , n7232 );
    or g1586 ( n5639 , n6288 , n1993 );
    nor g1587 ( n7024 , n5919 , n3749 );
    or g1588 ( n10981 , n1480 , n13494 );
    and g1589 ( n13076 , n1962 , n7270 );
    nor g1590 ( n2113 , n8856 , n3769 );
    and g1591 ( n315 , n12475 , n11782 );
    not g1592 ( n4790 , n9450 );
    or g1593 ( n11108 , n1223 , n14440 );
    not g1594 ( n10134 , n6139 );
    or g1595 ( n3490 , n8015 , n12655 );
    and g1596 ( n9401 , n231 , n12532 );
    not g1597 ( n11090 , n10629 );
    and g1598 ( n12001 , n11679 , n11725 );
    and g1599 ( n9632 , n5434 , n4993 );
    or g1600 ( n10559 , n10154 , n5515 );
    and g1601 ( n10204 , n4533 , n2848 );
    or g1602 ( n8803 , n1189 , n3962 );
    or g1603 ( n10612 , n4435 , n8615 );
    and g1604 ( n683 , n4394 , n10640 );
    not g1605 ( n4822 , n9580 );
    or g1606 ( n3281 , n2750 , n12656 );
    or g1607 ( n13590 , n317 , n11074 );
    or g1608 ( n13612 , n11935 , n12875 );
    not g1609 ( n1074 , n1639 );
    not g1610 ( n2177 , n12503 );
    and g1611 ( n5538 , n14093 , n13254 );
    nor g1612 ( n9701 , n11305 , n66 );
    nor g1613 ( n8751 , n4233 , n7244 );
    or g1614 ( n13803 , n5977 , n10013 );
    not g1615 ( n4722 , n8451 );
    or g1616 ( n11914 , n3320 , n5499 );
    nor g1617 ( n10263 , n5986 , n6047 );
    and g1618 ( n10171 , n14093 , n4635 );
    or g1619 ( n4087 , n8209 , n2498 );
    or g1620 ( n11356 , n2750 , n11639 );
    or g1621 ( n14323 , n4180 , n14431 );
    and g1622 ( n3486 , n9705 , n324 );
    or g1623 ( n9184 , n12576 , n156 );
    or g1624 ( n10621 , n10331 , n4053 );
    not g1625 ( n4439 , n2069 );
    or g1626 ( n2740 , n4033 , n12523 );
    not g1627 ( n5975 , n5449 );
    or g1628 ( n2466 , n11405 , n9999 );
    and g1629 ( n12716 , n627 , n8408 );
    and g1630 ( n1607 , n8412 , n13215 );
    or g1631 ( n13797 , n234 , n9667 );
    and g1632 ( n3274 , n4546 , n7425 );
    or g1633 ( n10202 , n8986 , n4732 );
    nor g1634 ( n13265 , n11765 , n11054 );
    and g1635 ( n707 , n6130 , n7366 );
    nor g1636 ( n9380 , n10312 , n6284 );
    and g1637 ( n8770 , n14091 , n3358 );
    not g1638 ( n2669 , n6829 );
    not g1639 ( n2566 , n13983 );
    nor g1640 ( n11732 , n13324 , n8072 );
    or g1641 ( n243 , n1660 , n7102 );
    or g1642 ( n13935 , n11360 , n9624 );
    or g1643 ( n6576 , n390 , n8356 );
    or g1644 ( n4778 , n14088 , n10361 );
    or g1645 ( n3288 , n1258 , n10605 );
    not g1646 ( n7898 , n13696 );
    or g1647 ( n1981 , n11303 , n601 );
    and g1648 ( n7276 , n12250 , n14159 );
    or g1649 ( n1284 , n14282 , n2751 );
    and g1650 ( n12520 , n11838 , n6934 );
    or g1651 ( n2685 , n6288 , n5609 );
    nor g1652 ( n5339 , n11285 , n10109 );
    nor g1653 ( n6279 , n2017 , n14017 );
    nor g1654 ( n5714 , n194 , n11184 );
    or g1655 ( n6632 , n8172 , n12734 );
    not g1656 ( n10512 , n10912 );
    or g1657 ( n7586 , n7736 , n579 );
    or g1658 ( n13177 , n1669 , n9699 );
    and g1659 ( n12027 , n9275 , n6970 );
    or g1660 ( n7649 , n4741 , n8110 );
    or g1661 ( n13195 , n7997 , n6517 );
    and g1662 ( n10521 , n10015 , n8187 );
    nor g1663 ( n9652 , n329 , n8902 );
    and g1664 ( n12892 , n541 , n12173 );
    or g1665 ( n11952 , n13675 , n3488 );
    and g1666 ( n10405 , n11867 , n13736 );
    and g1667 ( n1464 , n13252 , n9691 );
    and g1668 ( n12607 , n6527 , n2767 );
    or g1669 ( n8230 , n1535 , n13251 );
    nor g1670 ( n6 , n6953 , n12456 );
    not g1671 ( n9557 , n13784 );
    and g1672 ( n12326 , n4790 , n3238 );
    not g1673 ( n7188 , n12397 );
    or g1674 ( n3346 , n9211 , n916 );
    or g1675 ( n2355 , n3910 , n5467 );
    nor g1676 ( n2150 , n14466 , n8186 );
    or g1677 ( n4140 , n11459 , n1305 );
    or g1678 ( n11937 , n13718 , n12333 );
    not g1679 ( n2111 , n7441 );
    not g1680 ( n5288 , n13593 );
    not g1681 ( n1724 , n4595 );
    or g1682 ( n2991 , n1261 , n3426 );
    or g1683 ( n346 , n4468 , n4381 );
    and g1684 ( n3195 , n2564 , n6575 );
    or g1685 ( n6951 , n12712 , n12140 );
    and g1686 ( n8161 , n2669 , n6594 );
    or g1687 ( n8661 , n930 , n13583 );
    not g1688 ( n14074 , n10446 );
    or g1689 ( n1826 , n11542 , n12648 );
    and g1690 ( n9373 , n9819 , n8309 );
    or g1691 ( n7545 , n10136 , n13768 );
    and g1692 ( n8559 , n13484 , n12372 );
    and g1693 ( n7844 , n9952 , n11391 );
    not g1694 ( n5488 , n10282 );
    nor g1695 ( n10462 , n11680 , n1399 );
    or g1696 ( n3984 , n12400 , n10074 );
    or g1697 ( n9194 , n14401 , n6068 );
    or g1698 ( n11253 , n7736 , n7864 );
    not g1699 ( n14157 , n9197 );
    or g1700 ( n11836 , n839 , n3496 );
    and g1701 ( n4291 , n13078 , n861 );
    and g1702 ( n14487 , n14042 , n7083 );
    or g1703 ( n615 , n5315 , n13909 );
    or g1704 ( n14164 , n2080 , n10278 );
    or g1705 ( n8886 , n820 , n8705 );
    and g1706 ( n2860 , n13520 , n6757 );
    not g1707 ( n14249 , n14303 );
    and g1708 ( n4094 , n12412 , n5984 );
    not g1709 ( n568 , n3007 );
    or g1710 ( n12558 , n14337 , n11905 );
    or g1711 ( n4649 , n6711 , n3297 );
    and g1712 ( n1287 , n12542 , n922 );
    and g1713 ( n8596 , n13641 , n1394 );
    and g1714 ( n11833 , n9564 , n2410 );
    not g1715 ( n638 , n1843 );
    nor g1716 ( n12396 , n163 , n8612 );
    not g1717 ( n28 , n4203 );
    not g1718 ( n10310 , n3655 );
    or g1719 ( n1067 , n2229 , n2101 );
    and g1720 ( n1558 , n6318 , n14242 );
    and g1721 ( n1267 , n8500 , n13752 );
    and g1722 ( n9123 , n9191 , n13483 );
    and g1723 ( n11081 , n873 , n10158 );
    or g1724 ( n5452 , n9218 , n8494 );
    or g1725 ( n12738 , n13017 , n5185 );
    or g1726 ( n13926 , n12633 , n2517 );
    or g1727 ( n7904 , n8800 , n203 );
    and g1728 ( n9189 , n3485 , n7274 );
    and g1729 ( n14393 , n4095 , n6956 );
    or g1730 ( n825 , n2694 , n2351 );
    and g1731 ( n6151 , n13464 , n243 );
    and g1732 ( n655 , n3097 , n10246 );
    and g1733 ( n6126 , n4018 , n6912 );
    or g1734 ( n2489 , n4544 , n3198 );
    not g1735 ( n3587 , n2405 );
    not g1736 ( n7612 , n4131 );
    or g1737 ( n7498 , n10834 , n5146 );
    or g1738 ( n6890 , n8881 , n9636 );
    and g1739 ( n12367 , n12229 , n3869 );
    and g1740 ( n1994 , n2422 , n5397 );
    and g1741 ( n6656 , n12038 , n2602 );
    or g1742 ( n7822 , n12303 , n8262 );
    or g1743 ( n71 , n5483 , n11934 );
    or g1744 ( n12247 , n14466 , n6395 );
    nor g1745 ( n3924 , n7683 , n12451 );
    not g1746 ( n900 , n426 );
    nor g1747 ( n12612 , n3255 , n7386 );
    or g1748 ( n8788 , n12428 , n9426 );
    and g1749 ( n14064 , n2158 , n10667 );
    and g1750 ( n14468 , n12986 , n4956 );
    nor g1751 ( n2695 , n12292 , n7709 );
    or g1752 ( n5889 , n13516 , n12577 );
    not g1753 ( n13017 , n7988 );
    nor g1754 ( n8473 , n11492 , n3771 );
    not g1755 ( n7481 , n9453 );
    and g1756 ( n4345 , n2615 , n5893 );
    not g1757 ( n1535 , n9580 );
    and g1758 ( n2250 , n1136 , n6298 );
    or g1759 ( n559 , n3093 , n13133 );
    or g1760 ( n1934 , n1728 , n1310 );
    and g1761 ( n12925 , n673 , n13371 );
    or g1762 ( n13012 , n1332 , n11269 );
    or g1763 ( n5552 , n13485 , n4511 );
    or g1764 ( n9970 , n7418 , n10370 );
    not g1765 ( n10312 , n2451 );
    and g1766 ( n6931 , n11503 , n3955 );
    or g1767 ( n4625 , n10637 , n9133 );
    or g1768 ( n9849 , n1576 , n4427 );
    and g1769 ( n13503 , n4095 , n5979 );
    nor g1770 ( n1174 , n13522 , n6094 );
    and g1771 ( n8342 , n5279 , n9638 );
    and g1772 ( n5612 , n5048 , n2282 );
    nor g1773 ( n14385 , n10620 , n6416 );
    and g1774 ( n13782 , n11484 , n6510 );
    nor g1775 ( n6512 , n13759 , n4096 );
    or g1776 ( n3949 , n14481 , n5281 );
    and g1777 ( n8906 , n12445 , n1230 );
    or g1778 ( n1706 , n13102 , n7354 );
    or g1779 ( n5295 , n14188 , n8436 );
    or g1780 ( n3508 , n4913 , n11191 );
    nor g1781 ( n1798 , n5848 , n10737 );
    not g1782 ( n2845 , n12614 );
    and g1783 ( n4585 , n6486 , n1598 );
    and g1784 ( n10272 , n13823 , n3137 );
    and g1785 ( n4555 , n6957 , n307 );
    and g1786 ( n12293 , n4614 , n10237 );
    not g1787 ( n791 , n10985 );
    or g1788 ( n508 , n85 , n9469 );
    not g1789 ( n2742 , n316 );
    and g1790 ( n8113 , n7779 , n9597 );
    or g1791 ( n3270 , n13155 , n1511 );
    or g1792 ( n11545 , n8582 , n1123 );
    and g1793 ( n12699 , n3424 , n13039 );
    or g1794 ( n9698 , n5834 , n2106 );
    or g1795 ( n2992 , n6471 , n7186 );
    nor g1796 ( n2314 , n7052 , n2795 );
    not g1797 ( n1840 , n1041 );
    nor g1798 ( n13249 , n584 , n4663 );
    and g1799 ( n2190 , n7673 , n2274 );
    or g1800 ( n11509 , n13501 , n6795 );
    and g1801 ( n9578 , n12412 , n5473 );
    and g1802 ( n11675 , n7767 , n9713 );
    or g1803 ( n12227 , n5132 , n686 );
    not g1804 ( n6788 , n6254 );
    or g1805 ( n9603 , n4357 , n1907 );
    not g1806 ( n8656 , n11195 );
    nor g1807 ( n11147 , n8529 , n6966 );
    or g1808 ( n12366 , n6629 , n4982 );
    or g1809 ( n2366 , n8480 , n5031 );
    or g1810 ( n3765 , n10238 , n10750 );
    or g1811 ( n5954 , n10383 , n6336 );
    and g1812 ( n4088 , n13952 , n10748 );
    or g1813 ( n7318 , n1136 , n3799 );
    not g1814 ( n12179 , n5416 );
    not g1815 ( n5780 , n2369 );
    not g1816 ( n13835 , n12096 );
    not g1817 ( n1662 , n14525 );
    nor g1818 ( n2856 , n12040 , n8677 );
    not g1819 ( n7704 , n11870 );
    and g1820 ( n3154 , n12015 , n4816 );
    and g1821 ( n5292 , n9509 , n13917 );
    or g1822 ( n4388 , n2908 , n5588 );
    and g1823 ( n215 , n13359 , n715 );
    not g1824 ( n4655 , n14525 );
    not g1825 ( n1117 , n9450 );
    or g1826 ( n3626 , n5236 , n4853 );
    and g1827 ( n10107 , n2669 , n10761 );
    not g1828 ( n13597 , n1769 );
    and g1829 ( n4870 , n13421 , n2818 );
    or g1830 ( n13204 , n10461 , n2675 );
    or g1831 ( n8038 , n11620 , n10230 );
    not g1832 ( n9716 , n13668 );
    or g1833 ( n1186 , n7438 , n10882 );
    not g1834 ( n7938 , n8892 );
    and g1835 ( n155 , n2669 , n7166 );
    nor g1836 ( n13145 , n6041 , n6246 );
    and g1837 ( n11388 , n3435 , n5673 );
    not g1838 ( n12147 , n9950 );
    or g1839 ( n8675 , n5472 , n7062 );
    and g1840 ( n1318 , n13575 , n5320 );
    and g1841 ( n1941 , n7043 , n12884 );
    or g1842 ( n8567 , n9931 , n2361 );
    not g1843 ( n13236 , n8122 );
    nor g1844 ( n12451 , n1127 , n13753 );
    and g1845 ( n13760 , n9921 , n2443 );
    or g1846 ( n420 , n13485 , n3547 );
    or g1847 ( n11818 , n11901 , n6011 );
    or g1848 ( n7115 , n12336 , n12782 );
    or g1849 ( n9957 , n2843 , n2693 );
    and g1850 ( n8750 , n1210 , n13912 );
    not g1851 ( n13779 , n10368 );
    or g1852 ( n13239 , n10781 , n495 );
    not g1853 ( n7862 , n13901 );
    and g1854 ( n9418 , n2527 , n3045 );
    and g1855 ( n5880 , n14091 , n11059 );
    and g1856 ( n3143 , n8692 , n8470 );
    not g1857 ( n7609 , n8349 );
    not g1858 ( n11479 , n8800 );
    and g1859 ( n5730 , n1520 , n5135 );
    or g1860 ( n9360 , n14401 , n12784 );
    or g1861 ( n11643 , n28 , n8328 );
    or g1862 ( n11321 , n4684 , n11648 );
    or g1863 ( n10130 , n11704 , n4658 );
    and g1864 ( n9644 , n1339 , n6925 );
    and g1865 ( n13891 , n3607 , n14291 );
    not g1866 ( n2181 , n1220 );
    not g1867 ( n11428 , n5257 );
    not g1868 ( n10015 , n10975 );
    and g1869 ( n10800 , n5823 , n1175 );
    or g1870 ( n9044 , n9442 , n5850 );
    and g1871 ( n3284 , n11793 , n6638 );
    and g1872 ( n14215 , n10969 , n9392 );
    nor g1873 ( n5513 , n13365 , n8407 );
    and g1874 ( n1307 , n3675 , n11146 );
    or g1875 ( n7846 , n9654 , n8204 );
    and g1876 ( n10319 , n5779 , n4969 );
    and g1877 ( n9596 , n8814 , n9718 );
    or g1878 ( n8171 , n13142 , n4235 );
    not g1879 ( n14188 , n7404 );
    nor g1880 ( n964 , n5897 , n13505 );
    or g1881 ( n1504 , n13698 , n10463 );
    and g1882 ( n10124 , n965 , n338 );
    or g1883 ( n4787 , n9140 , n14087 );
    and g1884 ( n8622 , n4614 , n3216 );
    or g1885 ( n1000 , n13518 , n12511 );
    not g1886 ( n11867 , n9613 );
    and g1887 ( n11677 , n9972 , n11787 );
    nor g1888 ( n9482 , n13835 , n13569 );
    not g1889 ( n10815 , n14501 );
    nor g1890 ( n9901 , n7575 , n2881 );
    or g1891 ( n2155 , n3800 , n3459 );
    not g1892 ( n4637 , n2470 );
    not g1893 ( n11621 , n7289 );
    or g1894 ( n12652 , n1356 , n9139 );
    or g1895 ( n6064 , n4791 , n10867 );
    not g1896 ( n10562 , n9592 );
    nor g1897 ( n123 , n5486 , n11798 );
    and g1898 ( n9873 , n6486 , n697 );
    and g1899 ( n9760 , n5459 , n9549 );
    or g1900 ( n11570 , n2401 , n5874 );
    not g1901 ( n13433 , n11425 );
    nor g1902 ( n7444 , n6428 , n7801 );
    or g1903 ( n13136 , n13885 , n197 );
    not g1904 ( n9743 , n11511 );
    and g1905 ( n3116 , n8768 , n9833 );
    and g1906 ( n5251 , n1071 , n14383 );
    and g1907 ( n241 , n10760 , n14057 );
    and g1908 ( n4467 , n4657 , n7096 );
    or g1909 ( n410 , n5234 , n1600 );
    or g1910 ( n6956 , n11094 , n3323 );
    and g1911 ( n9600 , n2709 , n8949 );
    or g1912 ( n5673 , n5266 , n11865 );
    or g1913 ( n2335 , n11121 , n13331 );
    or g1914 ( n11549 , n7700 , n11266 );
    not g1915 ( n5253 , n3007 );
    or g1916 ( n11186 , n4684 , n1459 );
    and g1917 ( n8108 , n12531 , n10445 );
    and g1918 ( n11219 , n5092 , n2453 );
    or g1919 ( n479 , n10394 , n5235 );
    and g1920 ( n1765 , n3709 , n8319 );
    or g1921 ( n7446 , n10731 , n8739 );
    and g1922 ( n2556 , n8799 , n7638 );
    or g1923 ( n10250 , n2510 , n12621 );
    or g1924 ( n10058 , n11739 , n5884 );
    not g1925 ( n12412 , n12403 );
    or g1926 ( n761 , n3871 , n6738 );
    or g1927 ( n9012 , n1223 , n2716 );
    or g1928 ( n12199 , n13718 , n2860 );
    and g1929 ( n13946 , n1125 , n5923 );
    or g1930 ( n7428 , n4840 , n6577 );
    or g1931 ( n270 , n4828 , n3470 );
    and g1932 ( n7837 , n1729 , n12205 );
    or g1933 ( n6337 , n14430 , n3048 );
    and g1934 ( n3029 , n8630 , n217 );
    and g1935 ( n12378 , n10032 , n12081 );
    not g1936 ( n5180 , n8813 );
    or g1937 ( n12178 , n478 , n3556 );
    and g1938 ( n7339 , n5218 , n7689 );
    and g1939 ( n5152 , n8605 , n546 );
    or g1940 ( n6005 , n8277 , n11986 );
    not g1941 ( n1699 , n4824 );
    nor g1942 ( n6715 , n2822 , n6217 );
    nor g1943 ( n4960 , n8209 , n2811 );
    or g1944 ( n4786 , n6640 , n5601 );
    not g1945 ( n3165 , n5734 );
    or g1946 ( n1974 , n1834 , n7926 );
    nor g1947 ( n8730 , n13327 , n11046 );
    and g1948 ( n2914 , n10622 , n3060 );
    or g1949 ( n8651 , n3777 , n4069 );
    and g1950 ( n158 , n873 , n4749 );
    and g1951 ( n9133 , n2527 , n1420 );
    or g1952 ( n13312 , n8527 , n265 );
    and g1953 ( n3121 , n7187 , n8339 );
    or g1954 ( n12680 , n12821 , n11858 );
    and g1955 ( n10047 , n320 , n115 );
    or g1956 ( n7113 , n14449 , n8606 );
    and g1957 ( n3267 , n5335 , n14195 );
    not g1958 ( n93 , n12872 );
    not g1959 ( n11405 , n4606 );
    or g1960 ( n5198 , n10089 , n2452 );
    not g1961 ( n13383 , n4835 );
    or g1962 ( n6884 , n13718 , n13480 );
    and g1963 ( n8444 , n10516 , n14514 );
    and g1964 ( n9845 , n12445 , n3659 );
    not g1965 ( n4123 , n6999 );
    and g1966 ( n881 , n6527 , n10364 );
    not g1967 ( n14450 , n11930 );
    not g1968 ( n3485 , n7275 );
    and g1969 ( n5174 , n6753 , n7001 );
    not g1970 ( n11510 , n8595 );
    or g1971 ( n13280 , n13413 , n3438 );
    or g1972 ( n5232 , n8210 , n3981 );
    or g1973 ( n12944 , n5315 , n1087 );
    and g1974 ( n2972 , n12445 , n6026 );
    not g1975 ( n12808 , n1347 );
    and g1976 ( n11552 , n5434 , n11399 );
    or g1977 ( n6179 , n4498 , n13099 );
    and g1978 ( n8979 , n103 , n7585 );
    and g1979 ( n4413 , n9953 , n5677 );
    and g1980 ( n8716 , n4156 , n4071 );
    or g1981 ( n13742 , n1356 , n4551 );
    not g1982 ( n2897 , n11456 );
    and g1983 ( n5750 , n11607 , n4710 );
    or g1984 ( n4561 , n10615 , n9830 );
    and g1985 ( n1642 , n1138 , n5379 );
    not g1986 ( n4690 , n13447 );
    and g1987 ( n758 , n9232 , n9814 );
    or g1988 ( n8842 , n10083 , n713 );
    and g1989 ( n5119 , n2521 , n6059 );
    or g1990 ( n6934 , n8034 , n4478 );
    or g1991 ( n7776 , n791 , n5190 );
    and g1992 ( n8275 , n6013 , n1829 );
    or g1993 ( n5093 , n9375 , n9772 );
    and g1994 ( n2045 , n12521 , n8026 );
    and g1995 ( n11258 , n10516 , n6259 );
    or g1996 ( n10955 , n116 , n1352 );
    nor g1997 ( n618 , n3394 , n9092 );
    and g1998 ( n604 , n5275 , n1803 );
    not g1999 ( n7433 , n13890 );
    or g2000 ( n12325 , n2897 , n2927 );
    not g2001 ( n3526 , n1784 );
    not g2002 ( n769 , n1966 );
    or g2003 ( n11084 , n9375 , n13929 );
    or g2004 ( n4012 , n13080 , n10405 );
    or g2005 ( n11391 , n5007 , n5213 );
    not g2006 ( n13458 , n14406 );
    nor g2007 ( n11054 , n5271 , n11190 );
    nor g2008 ( n2255 , n955 , n7514 );
    not g2009 ( n679 , n9314 );
    and g2010 ( n8615 , n10668 , n7468 );
    and g2011 ( n53 , n4887 , n2505 );
    or g2012 ( n6676 , n5493 , n5448 );
    not g2013 ( n10449 , n1214 );
    or g2014 ( n11904 , n13083 , n6991 );
    and g2015 ( n451 , n11842 , n8518 );
    or g2016 ( n9083 , n11935 , n3035 );
    and g2017 ( n4843 , n5475 , n2279 );
    nor g2018 ( n606 , n11581 , n5015 );
    or g2019 ( n6827 , n480 , n13271 );
    and g2020 ( n7306 , n6606 , n3106 );
    and g2021 ( n7487 , n3923 , n3095 );
    and g2022 ( n6320 , n3766 , n4254 );
    or g2023 ( n7758 , n673 , n11875 );
    and g2024 ( n13054 , n9102 , n12384 );
    and g2025 ( n7622 , n5825 , n12552 );
    nor g2026 ( n12826 , n7662 , n1337 );
    or g2027 ( n5804 , n13112 , n4263 );
    and g2028 ( n7061 , n6192 , n12519 );
    and g2029 ( n11539 , n9571 , n10954 );
    and g2030 ( n3179 , n1662 , n9607 );
    nor g2031 ( n5599 , n2405 , n4471 );
    and g2032 ( n9608 , n14521 , n13989 );
    not g2033 ( n7146 , n3493 );
    or g2034 ( n1096 , n1821 , n2796 );
    or g2035 ( n3411 , n5507 , n3511 );
    and g2036 ( n8728 , n3286 , n10955 );
    not g2037 ( n4913 , n13165 );
    or g2038 ( n6536 , n2505 , n12009 );
    or g2039 ( n6077 , n12428 , n3520 );
    not g2040 ( n329 , n5974 );
    and g2041 ( n5638 , n12421 , n6080 );
    and g2042 ( n3518 , n12147 , n11913 );
    not g2043 ( n9563 , n4169 );
    and g2044 ( n4450 , n14358 , n6892 );
    and g2045 ( n6851 , n15 , n4083 );
    not g2046 ( n9285 , n1833 );
    nor g2047 ( n532 , n4210 , n6723 );
    or g2048 ( n8285 , n4233 , n3831 );
    or g2049 ( n13491 , n12353 , n5845 );
    not g2050 ( n4200 , n3094 );
    and g2051 ( n9565 , n1117 , n7839 );
    or g2052 ( n12429 , n14088 , n10531 );
    or g2053 ( n262 , n9780 , n10103 );
    or g2054 ( n10505 , n9806 , n10022 );
    or g2055 ( n2805 , n4739 , n7299 );
    and g2056 ( n8268 , n2758 , n6968 );
    and g2057 ( n1842 , n13367 , n10572 );
    and g2058 ( n2762 , n8047 , n6718 );
    and g2059 ( n2650 , n1854 , n13686 );
    and g2060 ( n9822 , n2521 , n9061 );
    nor g2061 ( n3032 , n12292 , n9590 );
    and g2062 ( n719 , n8432 , n7037 );
    or g2063 ( n9731 , n12695 , n5610 );
    and g2064 ( n11442 , n12857 , n3646 );
    or g2065 ( n1471 , n6607 , n793 );
    or g2066 ( n3688 , n2272 , n2239 );
    and g2067 ( n5772 , n5825 , n13071 );
    not g2068 ( n2527 , n9583 );
    or g2069 ( n4341 , n177 , n13295 );
    and g2070 ( n1083 , n8432 , n10621 );
    not g2071 ( n12334 , n9329 );
    or g2072 ( n13082 , n3888 , n5500 );
    and g2073 ( n9406 , n13682 , n2002 );
    or g2074 ( n8492 , n412 , n10176 );
    and g2075 ( n12260 , n1937 , n12342 );
    nor g2076 ( n3934 , n1425 , n1283 );
    or g2077 ( n3404 , n6867 , n5772 );
    and g2078 ( n445 , n2527 , n3005 );
    and g2079 ( n8947 , n3724 , n925 );
    or g2080 ( n8940 , n13531 , n8579 );
    nor g2081 ( n12269 , n8592 , n2234 );
    nor g2082 ( n11469 , n1628 , n4756 );
    not g2083 ( n4711 , n355 );
    not g2084 ( n8592 , n81 );
    and g2085 ( n3631 , n638 , n8681 );
    and g2086 ( n6296 , n12953 , n11318 );
    or g2087 ( n1999 , n14337 , n10762 );
    or g2088 ( n10054 , n13547 , n1764 );
    nor g2089 ( n580 , n14377 , n6158 );
    or g2090 ( n1230 , n11223 , n12600 );
    or g2091 ( n13954 , n2111 , n7248 );
    nor g2092 ( n12028 , n619 , n2195 );
    not g2093 ( n3907 , n9778 );
    and g2094 ( n1291 , n1074 , n6481 );
    or g2095 ( n5836 , n7438 , n4111 );
    or g2096 ( n1917 , n9422 , n7508 );
    and g2097 ( n11685 , n9853 , n12763 );
    and g2098 ( n14437 , n11329 , n8609 );
    nor g2099 ( n12790 , n11455 , n10222 );
    or g2100 ( n9836 , n4876 , n2397 );
    and g2101 ( n12902 , n4354 , n519 );
    and g2102 ( n2075 , n12592 , n12206 );
    and g2103 ( n14406 , n13728 , n6482 );
    and g2104 ( n10610 , n6609 , n12510 );
    not g2105 ( n5603 , n12106 );
    or g2106 ( n2286 , n6263 , n13568 );
    not g2107 ( n7063 , n6807 );
    not g2108 ( n12990 , n14501 );
    not g2109 ( n11546 , n7455 );
    and g2110 ( n4661 , n9323 , n7489 );
    nor g2111 ( n8586 , n4978 , n5635 );
    and g2112 ( n7296 , n13860 , n8059 );
    or g2113 ( n9978 , n2843 , n12634 );
    or g2114 ( n5298 , n163 , n1642 );
    and g2115 ( n3754 , n2486 , n6908 );
    and g2116 ( n10726 , n8247 , n11234 );
    and g2117 ( n13351 , n11422 , n3892 );
    or g2118 ( n12532 , n7481 , n3416 );
    and g2119 ( n9881 , n1857 , n12222 );
    or g2120 ( n10671 , n4468 , n7647 );
    and g2121 ( n11178 , n8401 , n4905 );
    and g2122 ( n5631 , n7171 , n9017 );
    or g2123 ( n7694 , n5562 , n9401 );
    not g2124 ( n5558 , n1985 );
    and g2125 ( n7771 , n1763 , n2488 );
    or g2126 ( n2606 , n8452 , n13001 );
    not g2127 ( n2529 , n6873 );
    not g2128 ( n4284 , n8027 );
    and g2129 ( n9330 , n10367 , n10076 );
    or g2130 ( n561 , n555 , n2353 );
    and g2131 ( n4753 , n79 , n2471 );
    and g2132 ( n3551 , n2006 , n12469 );
    or g2133 ( n4801 , n2089 , n4584 );
    or g2134 ( n5769 , n747 , n972 );
    or g2135 ( n6750 , n9111 , n9951 );
    not g2136 ( n2783 , n10303 );
    or g2137 ( n3001 , n1006 , n8293 );
    and g2138 ( n10196 , n15 , n5793 );
    not g2139 ( n4007 , n12765 );
    nor g2140 ( n5611 , n5762 , n11791 );
    or g2141 ( n14067 , n116 , n4812 );
    not g2142 ( n5427 , n4169 );
    and g2143 ( n6755 , n10922 , n5706 );
    not g2144 ( n8747 , n2320 );
    and g2145 ( n2930 , n7826 , n8658 );
    or g2146 ( n7861 , n4065 , n6627 );
    and g2147 ( n3173 , n7768 , n11394 );
    or g2148 ( n14197 , n7481 , n9386 );
    nor g2149 ( n8058 , n700 , n1793 );
    nor g2150 ( n13924 , n1929 , n8459 );
    and g2151 ( n7581 , n8692 , n3342 );
    and g2152 ( n5790 , n11020 , n9934 );
    not g2153 ( n11360 , n13668 );
    or g2154 ( n1085 , n13978 , n10138 );
    and g2155 ( n14 , n1904 , n2200 );
    and g2156 ( n7659 , n5857 , n11128 );
    and g2157 ( n3723 , n13656 , n1131 );
    not g2158 ( n10820 , n11548 );
    not g2159 ( n627 , n5182 );
    and g2160 ( n1517 , n4574 , n13403 );
    and g2161 ( n12489 , n9156 , n3583 );
    or g2162 ( n2788 , n11328 , n3532 );
    or g2163 ( n14092 , n49 , n664 );
    and g2164 ( n12405 , n3365 , n2974 );
    or g2165 ( n11128 , n283 , n3447 );
    and g2166 ( n13514 , n7063 , n12070 );
    not g2167 ( n9008 , n13509 );
    or g2168 ( n12962 , n1741 , n7470 );
    or g2169 ( n12579 , n553 , n439 );
    and g2170 ( n11606 , n4123 , n848 );
    or g2171 ( n10574 , n12131 , n11960 );
    or g2172 ( n12379 , n3569 , n13029 );
    and g2173 ( n14000 , n808 , n5680 );
    not g2174 ( n1299 , n5595 );
    not g2175 ( n10400 , n12925 );
    not g2176 ( n3076 , n13234 );
    and g2177 ( n2913 , n14327 , n13935 );
    and g2178 ( n9686 , n9329 , n14312 );
    nor g2179 ( n12315 , n1086 , n10565 );
    or g2180 ( n8100 , n6603 , n11714 );
    and g2181 ( n6665 , n6389 , n5554 );
    and g2182 ( n2612 , n8801 , n12415 );
    and g2183 ( n8024 , n9321 , n2800 );
    not g2184 ( n11384 , n2166 );
    and g2185 ( n14270 , n12057 , n8914 );
    and g2186 ( n11109 , n1339 , n10946 );
    and g2187 ( n11074 , n11240 , n3194 );
    nor g2188 ( n1241 , n13467 , n4237 );
    nor g2189 ( n5635 , n4135 , n1321 );
    and g2190 ( n12751 , n7068 , n8385 );
    or g2191 ( n12266 , n11438 , n2852 );
    and g2192 ( n5531 , n12226 , n8142 );
    and g2193 ( n10105 , n12265 , n6337 );
    nor g2194 ( n3971 , n13811 , n9170 );
    and g2195 ( n14502 , n7957 , n5068 );
    and g2196 ( n8418 , n4018 , n12213 );
    nor g2197 ( n1012 , n4050 , n11418 );
    or g2198 ( n14152 , n769 , n2770 );
    and g2199 ( n5146 , n4095 , n418 );
    or g2200 ( n1135 , n2179 , n9706 );
    or g2201 ( n3693 , n10933 , n8716 );
    or g2202 ( n2046 , n8582 , n11613 );
    and g2203 ( n11400 , n1339 , n8338 );
    or g2204 ( n13094 , n10383 , n5152 );
    and g2205 ( n2852 , n3635 , n11594 );
    and g2206 ( n9193 , n12808 , n5183 );
    not g2207 ( n5764 , n304 );
    and g2208 ( n10502 , n5038 , n6425 );
    or g2209 ( n8489 , n14370 , n7844 );
    or g2210 ( n11149 , n782 , n10654 );
    and g2211 ( n5532 , n6838 , n12642 );
    not g2212 ( n6128 , n261 );
    and g2213 ( n13591 , n6192 , n10261 );
    not g2214 ( n6768 , n2503 );
    nor g2215 ( n6358 , n1697 , n964 );
    not g2216 ( n9819 , n10862 );
    or g2217 ( n13415 , n12636 , n7667 );
    and g2218 ( n9939 , n7081 , n11777 );
    or g2219 ( n2096 , n7530 , n5231 );
    or g2220 ( n5716 , n1391 , n564 );
    not g2221 ( n9509 , n2906 );
    or g2222 ( n2441 , n14481 , n10753 );
    nor g2223 ( n11678 , n4741 , n4109 );
    not g2224 ( n4771 , n2370 );
    or g2225 ( n4746 , n5362 , n10582 );
    and g2226 ( n3946 , n12933 , n13466 );
    or g2227 ( n10841 , n11171 , n14003 );
    or g2228 ( n4949 , n5591 , n13186 );
    or g2229 ( n2161 , n13516 , n1324 );
    or g2230 ( n9262 , n7462 , n12815 );
    or g2231 ( n11319 , n9442 , n5194 );
    and g2232 ( n14269 , n1125 , n5967 );
    nor g2233 ( n9203 , n7036 , n11 );
    and g2234 ( n6033 , n13246 , n4483 );
    and g2235 ( n11523 , n1100 , n402 );
    nor g2236 ( n2690 , n4865 , n13416 );
    or g2237 ( n13321 , n11123 , n4361 );
    or g2238 ( n8685 , n11739 , n12795 );
    not g2239 ( n11738 , n9936 );
    or g2240 ( n12051 , n12131 , n12058 );
    or g2241 ( n5025 , n13220 , n9101 );
    or g2242 ( n1360 , n9111 , n4577 );
    and g2243 ( n12711 , n5628 , n1974 );
    or g2244 ( n12668 , n4180 , n7319 );
    and g2245 ( n869 , n12953 , n11241 );
    or g2246 ( n9575 , n1258 , n10918 );
    or g2247 ( n11625 , n4807 , n5711 );
    and g2248 ( n9947 , n7081 , n8553 );
    and g2249 ( n12789 , n13103 , n12485 );
    and g2250 ( n505 , n2983 , n248 );
    and g2251 ( n318 , n5071 , n14147 );
    and g2252 ( n4080 , n13107 , n5662 );
    or g2253 ( n12499 , n10396 , n12871 );
    and g2254 ( n10830 , n673 , n63 );
    or g2255 ( n6575 , n4205 , n8113 );
    or g2256 ( n10761 , n2318 , n770 );
    and g2257 ( n13999 , n3608 , n14076 );
    not g2258 ( n888 , n12573 );
    and g2259 ( n2460 , n10556 , n9393 );
    and g2260 ( n13221 , n6389 , n9202 );
    or g2261 ( n6252 , n13446 , n7630 );
    not g2262 ( n5574 , n462 );
    and g2263 ( n12621 , n2564 , n13902 );
    nor g2264 ( n2795 , n3230 , n5166 );
    and g2265 ( n4243 , n541 , n13263 );
    and g2266 ( n5622 , n10678 , n13120 );
    or g2267 ( n12109 , n8983 , n8715 );
    and g2268 ( n11631 , n14213 , n2487 );
    or g2269 ( n4802 , n11303 , n5783 );
    and g2270 ( n5340 , n1678 , n6338 );
    or g2271 ( n7067 , n8969 , n10799 );
    or g2272 ( n5321 , n1409 , n271 );
    nor g2273 ( n9352 , n1417 , n2030 );
    or g2274 ( n1205 , n89 , n4996 );
    or g2275 ( n1986 , n4357 , n1842 );
    or g2276 ( n5230 , n6090 , n5880 );
    and g2277 ( n11393 , n7748 , n9595 );
    or g2278 ( n11932 , n11090 , n802 );
    or g2279 ( n8384 , n3134 , n11361 );
    and g2280 ( n4014 , n13555 , n3057 );
    and g2281 ( n6748 , n10084 , n170 );
    or g2282 ( n5066 , n9211 , n9501 );
    nor g2283 ( n1501 , n8337 , n4687 );
    nor g2284 ( n1338 , n5504 , n6199 );
    and g2285 ( n3159 , n13781 , n12481 );
    not g2286 ( n5823 , n3926 );
    and g2287 ( n6850 , n7208 , n465 );
    and g2288 ( n1636 , n2330 , n8313 );
    or g2289 ( n9339 , n7245 , n4854 );
    nor g2290 ( n2118 , n6888 , n13406 );
    or g2291 ( n358 , n5587 , n14214 );
    or g2292 ( n9934 , n11097 , n796 );
    and g2293 ( n2313 , n5053 , n2976 );
    not g2294 ( n361 , n4606 );
    nor g2295 ( n3139 , n5621 , n4797 );
    nor g2296 ( n4795 , n600 , n2554 );
    or g2297 ( n143 , n13875 , n13513 );
    or g2298 ( n1457 , n5936 , n5733 );
    and g2299 ( n9024 , n9952 , n2155 );
    or g2300 ( n9163 , n1202 , n13600 );
    not g2301 ( n8223 , n8224 );
    and g2302 ( n6152 , n3710 , n1239 );
    and g2303 ( n14490 , n11814 , n4733 );
    nor g2304 ( n2554 , n7887 , n4718 );
    not g2305 ( n8950 , n13908 );
    nor g2306 ( n8420 , n1577 , n4196 );
    nor g2307 ( n10588 , n4333 , n13709 );
    and g2308 ( n14172 , n13877 , n14113 );
    or g2309 ( n2462 , n2615 , n8737 );
    not g2310 ( n9525 , n6928 );
    or g2311 ( n4367 , n3273 , n1183 );
    and g2312 ( n7162 , n1125 , n6484 );
    or g2313 ( n5875 , n6672 , n6145 );
    or g2314 ( n7873 , n1494 , n4115 );
    nor g2315 ( n1509 , n4091 , n4458 );
    not g2316 ( n12112 , n11331 );
    and g2317 ( n1540 , n428 , n2047 );
    not g2318 ( n1428 , n5153 );
    and g2319 ( n2743 , n7670 , n10773 );
    or g2320 ( n4965 , n1112 , n11235 );
    and g2321 ( n10468 , n13745 , n2542 );
    nor g2322 ( n5626 , n12651 , n4383 );
    or g2323 ( n10790 , n10871 , n9109 );
    not g2324 ( n9345 , n10469 );
    and g2325 ( n11005 , n14145 , n5533 );
    not g2326 ( n9377 , n2468 );
    or g2327 ( n8059 , n11097 , n12011 );
    nor g2328 ( n5879 , n13050 , n10878 );
    not g2329 ( n8008 , n12675 );
    and g2330 ( n14165 , n3536 , n3585 );
    and g2331 ( n4136 , n1772 , n10701 );
    or g2332 ( n4058 , n8301 , n11764 );
    or g2333 ( n6104 , n14166 , n3408 );
    or g2334 ( n7490 , n1623 , n8395 );
    not g2335 ( n4174 , n10714 );
    and g2336 ( n6546 , n14376 , n2537 );
    or g2337 ( n7504 , n1061 , n3834 );
    and g2338 ( n10949 , n10815 , n10866 );
    and g2339 ( n11900 , n5137 , n14115 );
    or g2340 ( n2051 , n8980 , n4403 );
    nor g2341 ( n7617 , n478 , n9862 );
    and g2342 ( n9748 , n9885 , n2304 );
    and g2343 ( n4469 , n11814 , n10188 );
    or g2344 ( n2980 , n6711 , n8535 );
    or g2345 ( n9072 , n5234 , n6472 );
    nor g2346 ( n7244 , n10368 , n9586 );
    and g2347 ( n4277 , n10408 , n13510 );
    or g2348 ( n10350 , n9429 , n2414 );
    not g2349 ( n425 , n692 );
    and g2350 ( n11559 , n1904 , n13940 );
    nor g2351 ( n681 , n2241 , n3171 );
    or g2352 ( n11173 , n3120 , n6900 );
    and g2353 ( n6019 , n9571 , n9002 );
    or g2354 ( n13962 , n6373 , n1291 );
    or g2355 ( n1596 , n5977 , n3612 );
    and g2356 ( n5520 , n627 , n9759 );
    or g2357 ( n12616 , n5625 , n4641 );
    or g2358 ( n8498 , n2474 , n11158 );
    or g2359 ( n5380 , n6206 , n6015 );
    and g2360 ( n13697 , n1588 , n11378 );
    not g2361 ( n3785 , n10368 );
    and g2362 ( n10826 , n9113 , n1691 );
    or g2363 ( n10011 , n1356 , n1731 );
    or g2364 ( n12066 , n8378 , n1106 );
    or g2365 ( n10816 , n9078 , n12987 );
    and g2366 ( n4691 , n9650 , n7633 );
    or g2367 ( n9392 , n10035 , n9071 );
    or g2368 ( n484 , n10062 , n9641 );
    or g2369 ( n752 , n7433 , n6258 );
    or g2370 ( n4476 , n11572 , n14504 );
    and g2371 ( n276 , n7826 , n6688 );
    or g2372 ( n3838 , n13074 , n4184 );
    and g2373 ( n11060 , n7391 , n5273 );
    and g2374 ( n10797 , n13078 , n420 );
    nor g2375 ( n7340 , n9525 , n9138 );
    or g2376 ( n169 , n6891 , n4410 );
    and g2377 ( n108 , n4156 , n11836 );
    or g2378 ( n10163 , n5468 , n1162 );
    and g2379 ( n1601 , n1804 , n3042 );
    and g2380 ( n13046 , n11702 , n13705 );
    and g2381 ( n328 , n6316 , n7416 );
    and g2382 ( n8682 , n9654 , n11479 );
    nor g2383 ( n12879 , n1575 , n454 );
    nor g2384 ( n5216 , n2087 , n6444 );
    or g2385 ( n1631 , n8726 , n12417 );
    and g2386 ( n7729 , n6525 , n9441 );
    not g2387 ( n10523 , n7289 );
    and g2388 ( n7994 , n627 , n2691 );
    nor g2389 ( n11993 , n1914 , n14044 );
    and g2390 ( n11370 , n13641 , n7228 );
    or g2391 ( n1187 , n12543 , n12219 );
    nor g2392 ( n3779 , n1742 , n11929 );
    not g2393 ( n9853 , n8650 );
    nor g2394 ( n344 , n13981 , n5041 );
    and g2395 ( n1943 , n13877 , n4860 );
    and g2396 ( n8009 , n5918 , n9574 );
    and g2397 ( n3880 , n8789 , n13386 );
    or g2398 ( n9861 , n4562 , n13495 );
    and g2399 ( n8497 , n4346 , n12893 );
    nor g2400 ( n14362 , n3333 , n4524 );
    or g2401 ( n14409 , n8747 , n10661 );
    and g2402 ( n13961 , n2422 , n7410 );
    and g2403 ( n12113 , n5926 , n562 );
    or g2404 ( n672 , n5815 , n13225 );
    or g2405 ( n8807 , n2531 , n2705 );
    nor g2406 ( n12268 , n14524 , n3225 );
    and g2407 ( n13262 , n8358 , n8741 );
    and g2408 ( n12882 , n10134 , n4372 );
    nor g2409 ( n6395 , n13081 , n3702 );
    or g2410 ( n1926 , n8726 , n8166 );
    and g2411 ( n1716 , n14321 , n11742 );
    and g2412 ( n11106 , n13676 , n10991 );
    or g2413 ( n1116 , n13220 , n10478 );
    and g2414 ( n6659 , n7079 , n9428 );
    or g2415 ( n10508 , n8580 , n12823 );
    nor g2416 ( n13640 , n1638 , n11993 );
    or g2417 ( n1212 , n5454 , n3961 );
    not g2418 ( n12169 , n11055 );
    and g2419 ( n2641 , n11614 , n10951 );
    or g2420 ( n11782 , n1838 , n3859 );
    or g2421 ( n6904 , n4967 , n11466 );
    and g2422 ( n8974 , n11008 , n1271 );
    or g2423 ( n12486 , n13991 , n13533 );
    not g2424 ( n12611 , n6807 );
    or g2425 ( n12350 , n5450 , n11635 );
    and g2426 ( n3654 , n11702 , n3727 );
    and g2427 ( n12715 , n10247 , n8489 );
    or g2428 ( n3596 , n11953 , n9145 );
    and g2429 ( n9767 , n6838 , n6112 );
    and g2430 ( n7486 , n9953 , n14363 );
    and g2431 ( n14309 , n2378 , n10559 );
    or g2432 ( n3463 , n8638 , n13609 );
    and g2433 ( n4565 , n12229 , n3615 );
    or g2434 ( n917 , n28 , n7642 );
    and g2435 ( n12181 , n889 , n12562 );
    or g2436 ( n8553 , n12400 , n5085 );
    or g2437 ( n5740 , n13083 , n9642 );
    not g2438 ( n6242 , n10346 );
    and g2439 ( n84 , n7673 , n11431 );
    nor g2440 ( n8214 , n727 , n5116 );
    and g2441 ( n5744 , n7957 , n3228 );
    and g2442 ( n2240 , n678 , n12898 );
    not g2443 ( n11761 , n14118 );
    and g2444 ( n7835 , n865 , n14217 );
    not g2445 ( n11157 , n8963 );
    and g2446 ( n196 , n14120 , n10291 );
    not g2447 ( n11183 , n12331 );
    and g2448 ( n11689 , n9198 , n5808 );
    nor g2449 ( n1111 , n7091 , n7954 );
    or g2450 ( n2399 , n12821 , n5708 );
    or g2451 ( n5202 , n5139 , n2588 );
    nor g2452 ( n2948 , n2016 , n10441 );
    or g2453 ( n161 , n13547 , n2492 );
    or g2454 ( n10301 , n12351 , n11537 );
    nor g2455 ( n3101 , n4589 , n4079 );
    or g2456 ( n3956 , n4498 , n6138 );
    and g2457 ( n5010 , n9811 , n10100 );
    not g2458 ( n3028 , n13365 );
    and g2459 ( n9351 , n7267 , n12717 );
    and g2460 ( n9240 , n13489 , n755 );
    and g2461 ( n8850 , n2177 , n8055 );
    or g2462 ( n14241 , n1805 , n4568 );
    or g2463 ( n6437 , n10960 , n9645 );
    or g2464 ( n10824 , n8737 , n4615 );
    not g2465 ( n9592 , n7931 );
    or g2466 ( n160 , n13310 , n3908 );
    and g2467 ( n8968 , n3268 , n2297 );
    or g2468 ( n7332 , n568 , n9508 );
    or g2469 ( n4576 , n12414 , n12635 );
    not g2470 ( n496 , n2932 );
    and g2471 ( n7685 , n6311 , n10988 );
    or g2472 ( n12114 , n2246 , n11783 );
    or g2473 ( n10961 , n5570 , n624 );
    and g2474 ( n4675 , n13520 , n6552 );
    or g2475 ( n2056 , n3120 , n6863 );
    or g2476 ( n1430 , n3168 , n13261 );
    or g2477 ( n7261 , n12821 , n1687 );
    not g2478 ( n2724 , n13181 );
    nor g2479 ( n2276 , n13875 , n1149 );
    not g2480 ( n12904 , n4379 );
    and g2481 ( n1833 , n11511 , n12243 );
    and g2482 ( n12855 , n2021 , n12579 );
    and g2483 ( n11613 , n6609 , n2570 );
    or g2484 ( n7816 , n9941 , n10765 );
    and g2485 ( n5672 , n12425 , n8723 );
    and g2486 ( n2539 , n5092 , n12262 );
    nor g2487 ( n2851 , n8404 , n6324 );
    nor g2488 ( n12005 , n9078 , n7890 );
    and g2489 ( n7991 , n12611 , n6427 );
    and g2490 ( n4867 , n13246 , n2902 );
    nor g2491 ( n10625 , n14166 , n13124 );
    nor g2492 ( n1185 , n11765 , n11125 );
    or g2493 ( n2627 , n11688 , n10050 );
    not g2494 ( n10238 , n9589 );
    nor g2495 ( n1321 , n13875 , n11131 );
    and g2496 ( n4725 , n5825 , n2719 );
    and g2497 ( n3289 , n9571 , n13095 );
    and g2498 ( n3066 , n4844 , n11397 );
    nor g2499 ( n8199 , n11870 , n10287 );
    and g2500 ( n4709 , n3212 , n2885 );
    and g2501 ( n1629 , n13781 , n4802 );
    and g2502 ( n4510 , n9792 , n6383 );
    and g2503 ( n4896 , n1431 , n7108 );
    not g2504 ( n8247 , n5108 );
    and g2505 ( n5987 , n4659 , n12912 );
    and g2506 ( n11268 , n13407 , n9166 );
    or g2507 ( n9054 , n5139 , n7989 );
    or g2508 ( n13218 , n5641 , n6034 );
    or g2509 ( n8961 , n1031 , n5163 );
    or g2510 ( n8795 , n2067 , n6555 );
    not g2511 ( n309 , n5118 );
    or g2512 ( n332 , n5236 , n7613 );
    and g2513 ( n8888 , n14358 , n6267 );
    or g2514 ( n8488 , n5483 , n12501 );
    and g2515 ( n2283 , n2587 , n7055 );
    not g2516 ( n9776 , n6520 );
    and g2517 ( n1938 , n679 , n7397 );
    not g2518 ( n6614 , n99 );
    and g2519 ( n6310 , n11422 , n14049 );
    or g2520 ( n3993 , n13142 , n6309 );
    and g2521 ( n2816 , n5591 , n5645 );
    or g2522 ( n14105 , n2179 , n1195 );
    and g2523 ( n319 , n6957 , n11585 );
    or g2524 ( n12676 , n2908 , n7610 );
    not g2525 ( n5779 , n1495 );
    or g2526 ( n10227 , n2089 , n477 );
    and g2527 ( n166 , n2422 , n7038 );
    and g2528 ( n7289 , n461 , n6614 );
    and g2529 ( n11649 , n5071 , n11879 );
    or g2530 ( n88 , n838 , n9407 );
    not g2531 ( n2179 , n238 );
    not g2532 ( n13327 , n13967 );
    not g2533 ( n12288 , n3742 );
    nor g2534 ( n5542 , n8816 , n10082 );
    and g2535 ( n13222 , n687 , n4304 );
    and g2536 ( n1978 , n10408 , n528 );
    or g2537 ( n2698 , n11909 , n5692 );
    and g2538 ( n7764 , n10332 , n1967 );
    not g2539 ( n5226 , n7832 );
    and g2540 ( n7928 , n446 , n11603 );
    not g2541 ( n8043 , n6119 );
    or g2542 ( n6238 , n4988 , n4622 );
    and g2543 ( n4970 , n1047 , n2960 );
    and g2544 ( n587 , n3755 , n13824 );
    nor g2545 ( n6172 , n5852 , n8370 );
    and g2546 ( n13799 , n12998 , n9532 );
    not g2547 ( n8527 , n9686 );
    and g2548 ( n6268 , n320 , n3549 );
    and g2549 ( n10708 , n7768 , n7181 );
    and g2550 ( n13463 , n6016 , n5498 );
    or g2551 ( n13451 , n4684 , n6009 );
    and g2552 ( n9504 , n7691 , n8087 );
    or g2553 ( n14159 , n2229 , n12665 );
    and g2554 ( n13871 , n12335 , n11989 );
    not g2555 ( n8769 , n5427 );
    or g2556 ( n4972 , n10534 , n8379 );
    and g2557 ( n6025 , n13103 , n5828 );
    and g2558 ( n13918 , n8025 , n12375 );
    not g2559 ( n10638 , n7518 );
    nor g2560 ( n14096 , n799 , n5043 );
    and g2561 ( n6487 , n965 , n12138 );
    and g2562 ( n94 , n7427 , n14497 );
    and g2563 ( n13371 , n5975 , n11385 );
    and g2564 ( n7329 , n5857 , n10450 );
    and g2565 ( n6031 , n12802 , n12669 );
    and g2566 ( n282 , n9015 , n629 );
    nor g2567 ( n8086 , n2017 , n8939 );
    and g2568 ( n2861 , n7768 , n41 );
    and g2569 ( n13028 , n1140 , n905 );
    or g2570 ( n9117 , n14472 , n10156 );
    or g2571 ( n8921 , n1844 , n8178 );
    or g2572 ( n8510 , n6672 , n3061 );
    nor g2573 ( n10387 , n13675 , n10719 );
    not g2574 ( n5195 , n5852 );
    or g2575 ( n10288 , n1147 , n3784 );
    or g2576 ( n10474 , n14107 , n8523 );
    or g2577 ( n10184 , n8969 , n5566 );
    and g2578 ( n4706 , n4104 , n1410 );
    or g2579 ( n1992 , n13537 , n1928 );
    and g2580 ( n5500 , n4358 , n5233 );
    not g2581 ( n7245 , n9596 );
    or g2582 ( n6464 , n7683 , n9246 );
    and g2583 ( n741 , n4156 , n5551 );
    and g2584 ( n2092 , n7970 , n10670 );
    or g2585 ( n12631 , n5732 , n4904 );
    or g2586 ( n12796 , n4255 , n509 );
    not g2587 ( n7075 , n13408 );
    not g2588 ( n12265 , n9197 );
    nor g2589 ( n4782 , n13458 , n5649 );
    or g2590 ( n3264 , n8726 , n8182 );
    and g2591 ( n8128 , n13227 , n11095 );
    or g2592 ( n11348 , n1362 , n8602 );
    or g2593 ( n2386 , n7212 , n3163 );
    or g2594 ( n9635 , n10825 , n9605 );
    or g2595 ( n11359 , n2149 , n6237 );
    nor g2596 ( n5497 , n13310 , n2807 );
    or g2597 ( n5537 , n4807 , n14103 );
    or g2598 ( n6533 , n9864 , n6780 );
    or g2599 ( n9991 , n12870 , n5532 );
    and g2600 ( n11076 , n9315 , n13082 );
    and g2601 ( n9049 , n9724 , n2965 );
    not g2602 ( n11909 , n14354 );
    and g2603 ( n11456 , n9679 , n5959 );
    or g2604 ( n4217 , n12712 , n9755 );
    and g2605 ( n7140 , n12229 , n4062 );
    and g2606 ( n13205 , n7221 , n7135 );
    or g2607 ( n13602 , n10784 , n10262 );
    and g2608 ( n7383 , n8247 , n3839 );
    not g2609 ( n3815 , n5901 );
    or g2610 ( n5337 , n9111 , n2280 );
    or g2611 ( n11811 , n11123 , n6573 );
    and g2612 ( n13972 , n11614 , n978 );
    or g2613 ( n1684 , n4562 , n4674 );
    nor g2614 ( n1791 , n6768 , n5006 );
    or g2615 ( n13245 , n1538 , n1242 );
    or g2616 ( n10778 , n2645 , n14468 );
    or g2617 ( n11863 , n12601 , n11252 );
    not g2618 ( n8168 , n14181 );
    or g2619 ( n7604 , n5491 , n11753 );
    not g2620 ( n9191 , n5460 );
    not g2621 ( n11938 , n4342 );
    or g2622 ( n5145 , n11935 , n9472 );
    nor g2623 ( n5051 , n11481 , n11073 );
    and g2624 ( n4001 , n5940 , n8811 );
    not g2625 ( n14433 , n6743 );
    or g2626 ( n8949 , n11704 , n11939 );
    not g2627 ( n920 , n4715 );
    or g2628 ( n5734 , n2090 , n9314 );
    and g2629 ( n10067 , n6898 , n4395 );
    nor g2630 ( n6474 , n3003 , n6729 );
    and g2631 ( n13963 , n678 , n13762 );
    and g2632 ( n10334 , n9297 , n6962 );
    and g2633 ( n535 , n55 , n7150 );
    or g2634 ( n4879 , n10731 , n4994 );
    and g2635 ( n10578 , n8512 , n10623 );
    not g2636 ( n7050 , n4518 );
    and g2637 ( n9489 , n10367 , n4594 );
    nor g2638 ( n8577 , n14196 , n5210 );
    or g2639 ( n811 , n1031 , n1874 );
    not g2640 ( n11220 , n3356 );
    or g2641 ( n5508 , n3777 , n864 );
    not g2642 ( n1071 , n11715 );
    or g2643 ( n2023 , n2901 , n11686 );
    or g2644 ( n10931 , n747 , n7347 );
    or g2645 ( n590 , n9507 , n4166 );
    not g2646 ( n986 , n5951 );
    and g2647 ( n14225 , n12015 , n5766 );
    or g2648 ( n4596 , n13854 , n9385 );
    or g2649 ( n9791 , n8096 , n5016 );
    and g2650 ( n1439 , n11033 , n8297 );
    and g2651 ( n4057 , n13626 , n8790 );
    nor g2652 ( n8389 , n450 , n5542 );
    or g2653 ( n13736 , n9541 , n3978 );
    and g2654 ( n4609 , n4146 , n5131 );
    and g2655 ( n5627 , n7846 , n2738 );
    or g2656 ( n2329 , n14472 , n2569 );
    or g2657 ( n7399 , n4923 , n404 );
    or g2658 ( n3827 , n7462 , n5019 );
    or g2659 ( n6707 , n7683 , n5376 );
    and g2660 ( n4326 , n10367 , n14515 );
    not g2661 ( n11325 , n2202 );
    or g2662 ( n4499 , n4923 , n4413 );
    and g2663 ( n1663 , n4354 , n8981 );
    nor g2664 ( n8374 , n10609 , n11178 );
    nor g2665 ( n13996 , n5833 , n5669 );
    and g2666 ( n4740 , n3813 , n6812 );
    and g2667 ( n8083 , n1904 , n4495 );
    not g2668 ( n1955 , n6305 );
    or g2669 ( n6986 , n6781 , n13046 );
    not g2670 ( n9793 , n7036 );
    not g2671 ( n12858 , n6113 );
    and g2672 ( n7320 , n6697 , n13123 );
    nor g2673 ( n11609 , n9807 , n12920 );
    and g2674 ( n12152 , n10458 , n7300 );
    or g2675 ( n7114 , n5891 , n13127 );
    or g2676 ( n5996 , n1061 , n4621 );
    and g2677 ( n10711 , n103 , n7572 );
    and g2678 ( n9965 , n2904 , n6064 );
    or g2679 ( n5443 , n9716 , n1978 );
    not g2680 ( n2575 , n3233 );
    nor g2681 ( n4064 , n6520 , n6482 );
    and g2682 ( n7936 , n14093 , n660 );
    or g2683 ( n277 , n9716 , n3227 );
    and g2684 ( n4492 , n14157 , n11592 );
    and g2685 ( n188 , n7187 , n2869 );
    nor g2686 ( n1463 , n6883 , n13244 );
    or g2687 ( n14263 , n11094 , n4014 );
    not g2688 ( n4468 , n3616 );
    not g2689 ( n9562 , n3673 );
    nor g2690 ( n13471 , n7245 , n13573 );
    or g2691 ( n3697 , n12568 , n4330 );
    and g2692 ( n9852 , n5553 , n8637 );
    or g2693 ( n2858 , n8980 , n7254 );
    or g2694 ( n14371 , n5997 , n5008 );
    or g2695 ( n11346 , n2597 , n8698 );
    and g2696 ( n5442 , n12542 , n8771 );
    or g2697 ( n13532 , n12169 , n1176 );
    and g2698 ( n10486 , n11803 , n8905 );
    or g2699 ( n10258 , n2016 , n8289 );
    nor g2700 ( n9047 , n8081 , n2085 );
    not g2701 ( n162 , n13900 );
    or g2702 ( n2102 , n11704 , n13961 );
    and g2703 ( n7915 , n13650 , n10002 );
    not g2704 ( n11105 , n14154 );
    or g2705 ( n4145 , n5936 , n6148 );
    or g2706 ( n8237 , n8881 , n11063 );
    and g2707 ( n7853 , n3536 , n3261 );
    and g2708 ( n8221 , n12615 , n475 );
    not g2709 ( n7057 , n8555 );
    and g2710 ( n14012 , n2724 , n11963 );
    nor g2711 ( n13586 , n3210 , n1682 );
    and g2712 ( n11053 , n13863 , n1774 );
    not g2713 ( n6000 , n12691 );
    and g2714 ( n7926 , n7391 , n6003 );
    and g2715 ( n3612 , n7767 , n13043 );
    nor g2716 ( n6790 , n12548 , n10475 );
    or g2717 ( n9394 , n13706 , n810 );
    and g2718 ( n5901 , n1506 , n3704 );
    or g2719 ( n13390 , n8507 , n9154 );
    and g2720 ( n3020 , n3169 , n3665 );
    or g2721 ( n11468 , n1051 , n4789 );
    and g2722 ( n4257 , n12042 , n10081 );
    and g2723 ( n2522 , n2521 , n11941 );
    or g2724 ( n11794 , n14088 , n5624 );
    not g2725 ( n4928 , n12975 );
    not g2726 ( n11071 , n2241 );
    not g2727 ( n4627 , n6113 );
    not g2728 ( n11739 , n10108 );
    or g2729 ( n12190 , n3062 , n5340 );
    nor g2730 ( n3645 , n3428 , n3927 );
    and g2731 ( n7322 , n8884 , n11882 );
    or g2732 ( n6214 , n13537 , n5332 );
    or g2733 ( n8738 , n13112 , n9946 );
    or g2734 ( n11835 , n9856 , n1301 );
    or g2735 ( n14308 , n13108 , n816 );
    and g2736 ( n6307 , n5011 , n1885 );
    and g2737 ( n11250 , n4851 , n13766 );
    and g2738 ( n2786 , n9944 , n6084 );
    and g2739 ( n6831 , n2942 , n11982 );
    not g2740 ( n3168 , n777 );
    or g2741 ( n10168 , n12844 , n3292 );
    and g2742 ( n12501 , n10930 , n14262 );
    and g2743 ( n7544 , n11838 , n7974 );
    and g2744 ( n1766 , n4486 , n4864 );
    or g2745 ( n12703 , n13941 , n13646 );
    not g2746 ( n12500 , n11152 );
    and g2747 ( n2536 , n13362 , n6473 );
    or g2748 ( n7323 , n6781 , n13558 );
    or g2749 ( n10840 , n10539 , n42 );
    nor g2750 ( n6117 , n4637 , n6089 );
    or g2751 ( n4947 , n1137 , n1830 );
    nor g2752 ( n12198 , n7245 , n7658 );
    nor g2753 ( n1519 , n3132 , n6048 );
    nor g2754 ( n5860 , n588 , n575 );
    not g2755 ( n8427 , n9197 );
    and g2756 ( n11912 , n12042 , n8722 );
    and g2757 ( n14258 , n3268 , n10452 );
    or g2758 ( n170 , n9403 , n8622 );
    or g2759 ( n11594 , n11710 , n7276 );
    and g2760 ( n9720 , n5275 , n5887 );
    and g2761 ( n11905 , n5252 , n11228 );
    or g2762 ( n13178 , n8332 , n4843 );
    or g2763 ( n12406 , n8513 , n8410 );
    and g2764 ( n6601 , n1489 , n9209 );
    and g2765 ( n14015 , n3755 , n14281 );
    or g2766 ( n7435 , n7436 , n4238 );
    and g2767 ( n11968 , n457 , n6871 );
    or g2768 ( n6452 , n10154 , n4935 );
    not g2769 ( n14039 , n6480 );
    not g2770 ( n12800 , n6554 );
    and g2771 ( n12387 , n2082 , n13930 );
    nor g2772 ( n10924 , n2790 , n12530 );
    or g2773 ( n14102 , n361 , n1646 );
    nor g2774 ( n9614 , n12522 , n7500 );
    or g2775 ( n2074 , n781 , n1783 );
    and g2776 ( n12074 , n10767 , n1325 );
    nor g2777 ( n5343 , n6313 , n13422 );
    not g2778 ( n298 , n13356 );
    or g2779 ( n8938 , n3125 , n3431 );
    or g2780 ( n13052 , n1356 , n13042 );
    and g2781 ( n1979 , n3492 , n11190 );
    not g2782 ( n13130 , n3046 );
    and g2783 ( n11507 , n12105 , n12830 );
    and g2784 ( n2827 , n392 , n3429 );
    or g2785 ( n13469 , n7914 , n141 );
    and g2786 ( n122 , n3491 , n8941 );
    or g2787 ( n14108 , n11459 , n6372 );
    not g2788 ( n4261 , n8555 );
    and g2789 ( n9129 , n4856 , n9940 );
    and g2790 ( n9419 , n1427 , n2785 );
    or g2791 ( n13817 , n14198 , n13440 );
    and g2792 ( n9254 , n8238 , n4076 );
    not g2793 ( n14065 , n6946 );
    not g2794 ( n14120 , n1120 );
    or g2795 ( n12416 , n13706 , n2097 );
    or g2796 ( n13687 , n1044 , n14328 );
    and g2797 ( n11032 , n12389 , n11716 );
    or g2798 ( n8684 , n838 , n11800 );
    or g2799 ( n10672 , n1802 , n10080 );
    not g2800 ( n8638 , n8813 );
    or g2801 ( n5667 , n5144 , n1213 );
    not g2802 ( n2686 , n11788 );
    or g2803 ( n367 , n3445 , n10421 );
    or g2804 ( n418 , n8480 , n11553 );
    and g2805 ( n13294 , n8923 , n924 );
    or g2806 ( n14195 , n14058 , n4016 );
    not g2807 ( n8529 , n1997 );
    not g2808 ( n7934 , n13625 );
    nor g2809 ( n9378 , n4544 , n2398 );
    nor g2810 ( n1744 , n3444 , n6447 );
    and g2811 ( n3201 , n7779 , n13843 );
    or g2812 ( n8026 , n2055 , n4268 );
    not g2813 ( n12757 , n10965 );
    and g2814 ( n1841 , n8965 , n9114 );
    and g2815 ( n1062 , n4698 , n10198 );
    and g2816 ( n6058 , n11687 , n220 );
    or g2817 ( n7882 , n14029 , n2926 );
    and g2818 ( n4781 , n12259 , n728 );
    and g2819 ( n9656 , n5628 , n1565 );
    nor g2820 ( n8762 , n8877 , n13063 );
    or g2821 ( n3935 , n13155 , n10879 );
    or g2822 ( n8561 , n7364 , n13603 );
    and g2823 ( n6522 , n7419 , n8129 );
    and g2824 ( n9383 , n3 , n1292 );
    and g2825 ( n11415 , n11218 , n5782 );
    nor g2826 ( n8548 , n7359 , n8389 );
    or g2827 ( n7773 , n361 , n124 );
    or g2828 ( n2455 , n49 , n2648 );
    or g2829 ( n5831 , n11704 , n2278 );
    nor g2830 ( n9396 , n5391 , n5585 );
    and g2831 ( n4982 , n9811 , n1950 );
    and g2832 ( n9897 , n9617 , n11140 );
    or g2833 ( n10343 , n5406 , n10686 );
    or g2834 ( n10895 , n9229 , n6126 );
    and g2835 ( n7499 , n4300 , n14470 );
    or g2836 ( n6438 , n6654 , n10424 );
    not g2837 ( n5665 , n11347 );
    and g2838 ( n4859 , n1203 , n9008 );
    and g2839 ( n9322 , n1339 , n10003 );
    and g2840 ( n9421 , n10408 , n383 );
    or g2841 ( n9411 , n11121 , n12398 );
    and g2842 ( n4025 , n11674 , n3763 );
    not g2843 ( n6679 , n2996 );
    or g2844 ( n2357 , n13209 , n3910 );
    not g2845 ( n11474 , n6212 );
    and g2846 ( n2581 , n13535 , n3956 );
    not g2847 ( n2229 , n4609 );
    or g2848 ( n7924 , n6730 , n6216 );
    or g2849 ( n6469 , n1669 , n13423 );
    or g2850 ( n12781 , n9984 , n7195 );
    and g2851 ( n1935 , n5104 , n2898 );
    and g2852 ( n6359 , n10589 , n12261 );
    or g2853 ( n8501 , n7530 , n11419 );
    or g2854 ( n13275 , n6607 , n1345 );
    or g2855 ( n1415 , n480 , n13922 );
    or g2856 ( n7342 , n13155 , n8400 );
    not g2857 ( n12192 , n2332 );
    nor g2858 ( n7695 , n5480 , n1092 );
    nor g2859 ( n11280 , n8361 , n3582 );
    and g2860 ( n11467 , n1588 , n538 );
    or g2861 ( n236 , n3512 , n8283 );
    or g2862 ( n3979 , n13718 , n2490 );
    and g2863 ( n3423 , n13379 , n4012 );
    and g2864 ( n6935 , n14145 , n7085 );
    or g2865 ( n11462 , n4876 , n8967 );
    and g2866 ( n3246 , n5628 , n3036 );
    nor g2867 ( n2892 , n3802 , n6150 );
    and g2868 ( n3511 , n13952 , n6032 );
    or g2869 ( n8686 , n11048 , n4408 );
    nor g2870 ( n6729 , n10136 , n8481 );
    not g2871 ( n2752 , n10861 );
    not g2872 ( n1356 , n7819 );
    or g2873 ( n4593 , n5800 , n2373 );
    and g2874 ( n11039 , n6311 , n10875 );
    nor g2875 ( n483 , n13435 , n13939 );
    or g2876 ( n14069 , n1840 , n7185 );
    not g2877 ( n392 , n14525 );
    or g2878 ( n3856 , n5064 , n3519 );
    and g2879 ( n7239 , n12721 , n9262 );
    nor g2880 ( n13193 , n11706 , n5196 );
    and g2881 ( n6433 , n2158 , n8530 );
    or g2882 ( n5572 , n4052 , n11013 );
    or g2883 ( n5254 , n14481 , n12387 );
    not g2884 ( n12038 , n5153 );
    or g2885 ( n3348 , n10331 , n4813 );
    and g2886 ( n10799 , n12038 , n1884 );
    and g2887 ( n2426 , n9920 , n6045 );
    or g2888 ( n798 , n8242 , n10313 );
    or g2889 ( n6633 , n2843 , n14022 );
    not g2890 ( n8424 , n5761 );
    nor g2891 ( n4756 , n6326 , n11911 );
    or g2892 ( n5830 , n11440 , n13552 );
    and g2893 ( n7167 , n11220 , n8510 );
    or g2894 ( n3955 , n14404 , n2715 );
    and g2895 ( n7610 , n8965 , n8448 );
    or g2896 ( n3793 , n6607 , n13232 );
    or g2897 ( n10104 , n9423 , n4570 );
    and g2898 ( n8005 , n446 , n14237 );
    and g2899 ( n9106 , n12990 , n547 );
    and g2900 ( n6006 , n898 , n10950 );
    and g2901 ( n3567 , n11411 , n1286 );
    or g2902 ( n7576 , n12622 , n2502 );
    and g2903 ( n5961 , n8789 , n518 );
    not g2904 ( n13408 , n12069 );
    or g2905 ( n9844 , n11953 , n10711 );
    and g2906 ( n13593 , n12852 , n5398 );
    or g2907 ( n6446 , n4913 , n12376 );
    and g2908 ( n11893 , n11702 , n7360 );
    and g2909 ( n1122 , n12270 , n6384 );
    nor g2910 ( n6723 , n4082 , n356 );
    and g2911 ( n10433 , n3276 , n5249 );
    and g2912 ( n6922 , n11737 , n1785 );
    nor g2913 ( n3894 , n13213 , n14183 );
    or g2914 ( n9628 , n1660 , n205 );
    and g2915 ( n4374 , n5553 , n5456 );
    and g2916 ( n2320 , n5678 , n6099 );
    nor g2917 ( n3355 , n10637 , n13776 );
    not g2918 ( n5621 , n11350 );
    not g2919 ( n482 , n2462 );
    or g2920 ( n219 , n13991 , n4492 );
    and g2921 ( n4265 , n9238 , n5204 );
    nor g2922 ( n8154 , n12888 , n11566 );
    not g2923 ( n10197 , n9583 );
    or g2924 ( n12506 , n10360 , n7272 );
    or g2925 ( n1161 , n2924 , n6362 );
    and g2926 ( n9649 , n13863 , n13336 );
    and g2927 ( n2770 , n12421 , n3218 );
    or g2928 ( n1516 , n5406 , n4148 );
    not g2929 ( n116 , n14412 );
    or g2930 ( n10532 , n1261 , n10256 );
    or g2931 ( n9346 , n6706 , n6001 );
    nor g2932 ( n5243 , n5505 , n5497 );
    and g2933 ( n11823 , n4973 , n13619 );
    nor g2934 ( n5982 , n2057 , n3487 );
    nor g2935 ( n6125 , n10649 , n386 );
    or g2936 ( n11239 , n10289 , n13492 );
    or g2937 ( n7899 , n12651 , n2929 );
    not g2938 ( n222 , n1639 );
    or g2939 ( n9877 , n14282 , n7765 );
    not g2940 ( n10854 , n12450 );
    and g2941 ( n5436 , n5926 , n9915 );
    not g2942 ( n10781 , n5627 );
    and g2943 ( n11342 , n7911 , n5327 );
    and g2944 ( n9866 , n7970 , n4576 );
    or g2945 ( n14140 , n9541 , n4466 );
    and g2946 ( n5028 , n12521 , n357 );
    and g2947 ( n11224 , n3715 , n12212 );
    or g2948 ( n12221 , n6111 , n12184 );
    not g2949 ( n13967 , n7091 );
    nor g2950 ( n7197 , n2098 , n5938 );
    or g2951 ( n6098 , n9211 , n24 );
    and g2952 ( n7823 , n12105 , n11098 );
    or g2953 ( n2629 , n7898 , n13571 );
    and g2954 ( n11414 , n103 , n5670 );
    or g2955 ( n7637 , n2888 , n10870 );
    and g2956 ( n13257 , n12779 , n1210 );
    or g2957 ( n6236 , n4821 , n3707 );
    and g2958 ( n14382 , n2330 , n3335 );
    nor g2959 ( n2544 , n7359 , n7692 );
    and g2960 ( n10230 , n3785 , n694 );
    and g2961 ( n1215 , n9617 , n7198 );
    and g2962 ( n11986 , n10374 , n7607 );
    and g2963 ( n12166 , n7354 , n3734 );
    or g2964 ( n12080 , n3667 , n6604 );
    or g2965 ( n980 , n12139 , n812 );
    and g2966 ( n12331 , n8446 , n8131 );
    or g2967 ( n10992 , n900 , n11038 );
    or g2968 ( n14462 , n12131 , n12118 );
    not g2969 ( n6023 , n1568 );
    and g2970 ( n3784 , n2961 , n9522 );
    or g2971 ( n1690 , n584 , n5074 );
    and g2972 ( n5419 , n12953 , n9851 );
    nor g2973 ( n4093 , n8701 , n2515 );
    or g2974 ( n2959 , n9742 , n4005 );
    and g2975 ( n9481 , n3536 , n371 );
    not g2976 ( n3320 , n8148 );
    or g2977 ( n1058 , n11542 , n4543 );
    and g2978 ( n5168 , n2461 , n12854 );
    not g2979 ( n12200 , n5678 );
    and g2980 ( n7131 , n8849 , n11022 );
    and g2981 ( n1450 , n9080 , n7648 );
    not g2982 ( n1218 , n2577 );
    or g2983 ( n11660 , n7938 , n1268 );
    nor g2984 ( n10746 , n8015 , n14104 );
    and g2985 ( n12441 , n3405 , n8406 );
    and g2986 ( n4449 , n11737 , n652 );
    and g2987 ( n11375 , n13867 , n5663 );
    or g2988 ( n13774 , n6163 , n8753 );
    or g2989 ( n7910 , n5007 , n5442 );
    not g2990 ( n12057 , n8650 );
    or g2991 ( n5461 , n5815 , n2590 );
    and g2992 ( n3186 , n2422 , n2300 );
    not g2993 ( n11953 , n4317 );
    and g2994 ( n7865 , n13484 , n11202 );
    or g2995 ( n8149 , n9422 , n10207 );
    and g2996 ( n959 , n1804 , n671 );
    not g2997 ( n13572 , n3870 );
    not g2998 ( n3959 , n13476 );
    or g2999 ( n12337 , n5406 , n2092 );
    not g3000 ( n1526 , n13213 );
    not g3001 ( n12999 , n14320 );
    not g3002 ( n10374 , n8451 );
    or g3003 ( n6548 , n11620 , n13606 );
    or g3004 ( n9278 , n9742 , n6522 );
    or g3005 ( n4106 , n2086 , n5822 );
    not g3006 ( n3536 , n5460 );
    and g3007 ( n13397 , n8183 , n7807 );
    not g3008 ( n11472 , n3616 );
    and g3009 ( n1799 , n3424 , n1998 );
    or g3010 ( n11840 , n9353 , n2823 );
    and g3011 ( n5313 , n8393 , n11972 );
    or g3012 ( n4286 , n13518 , n3012 );
    or g3013 ( n8500 , n1850 , n10446 );
    nor g3014 ( n7008 , n6765 , n13313 );
    or g3015 ( n5466 , n766 , n2576 );
    and g3016 ( n5992 , n405 , n10143 );
    nor g3017 ( n701 , n11975 , n2424 );
    not g3018 ( n13447 , n6714 );
    and g3019 ( n2987 , n1452 , n499 );
    and g3020 ( n10526 , n8412 , n14069 );
    and g3021 ( n10242 , n2983 , n12476 );
    and g3022 ( n6668 , n8453 , n5863 );
    or g3023 ( n1199 , n11839 , n7040 );
    and g3024 ( n8948 , n11153 , n11750 );
    or g3025 ( n9327 , n11558 , n14264 );
    not g3026 ( n457 , n12450 );
    and g3027 ( n7062 , n2904 , n2836 );
    nor g3028 ( n4307 , n9529 , n7371 );
    or g3029 ( n6720 , n7530 , n1320 );
    and g3030 ( n10251 , n8630 , n1683 );
    not g3031 ( n13209 , n8873 );
    nor g3032 ( n237 , n2799 , n9039 );
    or g3033 ( n5793 , n10784 , n7977 );
    or g3034 ( n13733 , n9490 , n4700 );
    and g3035 ( n9283 , n7053 , n10839 );
    nor g3036 ( n13208 , n3248 , n13858 );
    and g3037 ( n7112 , n3286 , n11217 );
    and g3038 ( n11127 , n7370 , n13932 );
    or g3039 ( n12642 , n2761 , n5983 );
    not g3040 ( n6711 , n10346 );
    nor g3041 ( n14070 , n1112 , n4848 );
    and g3042 ( n13907 , n13641 , n10805 );
    or g3043 ( n768 , n3815 , n11311 );
    not g3044 ( n6130 , n5606 );
    or g3045 ( n14281 , n4033 , n12892 );
    or g3046 ( n4483 , n10523 , n11230 );
    or g3047 ( n11159 , n5807 , n10129 );
    or g3048 ( n9689 , n6039 , n1372 );
    nor g3049 ( n1777 , n8877 , n13670 );
    or g3050 ( n13737 , n3768 , n5826 );
    not g3051 ( n2069 , n1760 );
    or g3052 ( n4171 , n13226 , n9696 );
    nor g3053 ( n11805 , n5605 , n36 );
    nor g3054 ( n6817 , n584 , n6590 );
    and g3055 ( n5019 , n8183 , n5036 );
    nor g3056 ( n3702 , n7011 , n5410 );
    not g3057 ( n13421 , n6657 );
    or g3058 ( n6334 , n10624 , n617 );
    or g3059 ( n2837 , n4898 , n6110 );
    not g3060 ( n13298 , n3230 );
    and g3061 ( n1329 , n1268 , n2255 );
    and g3062 ( n13308 , n5471 , n11693 );
    and g3063 ( n13513 , n4619 , n11600 );
    and g3064 ( n12948 , n8692 , n7668 );
    not g3065 ( n13050 , n13158 );
    and g3066 ( n10605 , n1610 , n10123 );
    and g3067 ( n10484 , n7267 , n8256 );
    and g3068 ( n7461 , n5317 , n8237 );
    or g3069 ( n5994 , n5997 , n4223 );
    or g3070 ( n11236 , n8513 , n753 );
    and g3071 ( n9813 , n5926 , n13933 );
    or g3072 ( n4857 , n8969 , n6429 );
    or g3073 ( n12869 , n9111 , n8094 );
    nor g3074 ( n7981 , n448 , n3726 );
    nor g3075 ( n7946 , n3577 , n1063 );
    nor g3076 ( n11641 , n10241 , n2612 );
    and g3077 ( n10153 , n8697 , n7944 );
    nor g3078 ( n1712 , n10312 , n13148 );
    and g3079 ( n5479 , n14072 , n5728 );
    or g3080 ( n9438 , n14107 , n595 );
    or g3081 ( n763 , n4065 , n14015 );
    or g3082 ( n7111 , n8476 , n6411 );
    and g3083 ( n9979 , n11569 , n2436 );
    and g3084 ( n10490 , n4261 , n13305 );
    or g3085 ( n14167 , n2518 , n1867 );
    and g3086 ( n14171 , n13535 , n14345 );
    or g3087 ( n11873 , n2878 , n7042 );
    or g3088 ( n1351 , n1044 , n6919 );
    not g3089 ( n4407 , n1833 );
    not g3090 ( n500 , n4634 );
    and g3091 ( n6719 , n6724 , n8589 );
    or g3092 ( n259 , n7862 , n13732 );
    and g3093 ( n8588 , n222 , n14494 );
    or g3094 ( n6917 , n3545 , n8100 );
    or g3095 ( n10978 , n11123 , n5630 );
    and g3096 ( n2956 , n5071 , n6452 );
    and g3097 ( n5140 , n12460 , n7796 );
    or g3098 ( n2094 , n10050 , n5046 );
    nor g3099 ( n5893 , n7755 , n4662 );
    or g3100 ( n10023 , n1172 , n805 );
    and g3101 ( n12588 , n13756 , n3037 );
    not g3102 ( n13535 , n10322 );
    nor g3103 ( n13498 , n11428 , n8727 );
    and g3104 ( n8791 , n14327 , n5329 );
    nor g3105 ( n3909 , n2094 , n9017 );
    and g3106 ( n1600 , n11329 , n7517 );
    and g3107 ( n2192 , n14446 , n12682 );
    not g3108 ( n2055 , n4777 );
    or g3109 ( n2430 , n5647 , n6262 );
    not g3110 ( n10595 , n14332 );
    or g3111 ( n1630 , n5483 , n8342 );
    nor g3112 ( n9765 , n11667 , n6877 );
    and g3113 ( n12778 , n2587 , n2657 );
    or g3114 ( n6375 , n3168 , n12373 );
    nor g3115 ( n6567 , n2923 , n8134 );
    or g3116 ( n1035 , n1258 , n7531 );
    and g3117 ( n1482 , n13863 , n10831 );
    or g3118 ( n4327 , n1189 , n8343 );
    and g3119 ( n5246 , n2998 , n6464 );
    nor g3120 ( n12380 , n8752 , n10326 );
    and g3121 ( n11306 , n5458 , n10939 );
    and g3122 ( n3830 , n11411 , n14045 );
    and g3123 ( n2635 , n3724 , n4697 );
    or g3124 ( n6911 , n7116 , n7417 );
    not g3125 ( n5553 , n2619 );
    not g3126 ( n8376 , n1637 );
    or g3127 ( n14506 , n13675 , n12883 );
    not g3128 ( n11303 , n11456 );
    not g3129 ( n5035 , n56 );
    nor g3130 ( n2128 , n5833 , n11376 );
    and g3131 ( n7711 , n6609 , n6548 );
    nor g3132 ( n11812 , n7227 , n1675 );
    not g3133 ( n2180 , n9546 );
    or g3134 ( n14094 , n12633 , n9196 );
    or g3135 ( n9204 , n9269 , n1696 );
    or g3136 ( n2248 , n5800 , n2972 );
    and g3137 ( n6451 , n14210 , n12964 );
    nor g3138 ( n8072 , n1914 , n5912 );
    nor g3139 ( n10308 , n1914 , n13637 );
    and g3140 ( n6550 , n6753 , n7903 );
    or g3141 ( n3758 , n14058 , n6644 );
    and g3142 ( n10742 , n10072 , n1232 );
    and g3143 ( n7321 , n873 , n1015 );
    and g3144 ( n3000 , n4394 , n3050 );
    or g3145 ( n13356 , n5467 , n7282 );
    or g3146 ( n8037 , n9151 , n11494 );
    and g3147 ( n9474 , n13780 , n586 );
    or g3148 ( n3071 , n13847 , n8119 );
    and g3149 ( n5264 , n7053 , n10794 );
    and g3150 ( n7159 , n10909 , n6802 );
    not g3151 ( n7429 , n8168 );
    and g3152 ( n12014 , n8450 , n1469 );
    nor g3153 ( n1337 , n3427 , n10697 );
    or g3154 ( n611 , n3009 , n3609 );
    and g3155 ( n339 , n5948 , n13898 );
    and g3156 ( n11583 , n2367 , n13783 );
    and g3157 ( n2184 , n13236 , n14095 );
    not g3158 ( n4424 , n12189 );
    or g3159 ( n9089 , n11097 , n2325 );
    and g3160 ( n10027 , n4546 , n12729 );
    or g3161 ( n11669 , n14400 , n10684 );
    and g3162 ( n7154 , n6609 , n10053 );
    not g3163 ( n3271 , n4774 );
    nor g3164 ( n10823 , n10186 , n6476 );
    or g3165 ( n2821 , n1728 , n5179 );
    or g3166 ( n12029 , n7358 , n14278 );
    not g3167 ( n2562 , n14354 );
    or g3168 ( n9335 , n12500 , n2909 );
    not g3169 ( n12821 , n8272 );
    or g3170 ( n3213 , n14472 , n9464 );
    or g3171 ( n7174 , n3219 , n7283 );
    or g3172 ( n3282 , n2750 , n11958 );
    nor g3173 ( n13406 , n12568 , n12170 );
    and g3174 ( n10791 , n10378 , n2014 );
    and g3175 ( n608 , n9190 , n3783 );
    and g3176 ( n7031 , n8932 , n6619 );
    or g3177 ( n10701 , n2086 , n2647 );
    and g3178 ( n10704 , n5899 , n6136 );
    or g3179 ( n13813 , n10300 , n5796 );
    or g3180 ( n8509 , n1834 , n331 );
    or g3181 ( n5969 , n2761 , n5462 );
    or g3182 ( n1053 , n7476 , n5943 );
    and g3183 ( n11844 , n10562 , n12 );
    and g3184 ( n1878 , n898 , n3275 );
    not g3185 ( n512 , n8162 );
    not g3186 ( n2906 , n6855 );
    and g3187 ( n10113 , n8768 , n10409 );
    and g3188 ( n10755 , n9232 , n13115 );
    not g3189 ( n5606 , n8927 );
    not g3190 ( n11020 , n3313 );
    or g3191 ( n8170 , n5507 , n11464 );
    and g3192 ( n3563 , n6525 , n8373 );
    and g3193 ( n2221 , n9705 , n5200 );
    not g3194 ( n5548 , n630 );
    and g3195 ( n11021 , n11867 , n12639 );
    not g3196 ( n13875 , n4325 );
    or g3197 ( n12783 , n7678 , n596 );
    or g3198 ( n14428 , n251 , n12448 );
    and g3199 ( n6368 , n4484 , n7318 );
    or g3200 ( n10161 , n7898 , n12584 );
    or g3201 ( n5659 , n7250 , n8601 );
    and g3202 ( n3948 , n14120 , n2748 );
    not g3203 ( n4619 , n3922 );
    or g3204 ( n2506 , n9403 , n5991 );
    and g3205 ( n2725 , n13107 , n1658 );
    or g3206 ( n7337 , n553 , n13315 );
    or g3207 ( n11293 , n7684 , n8918 );
    and g3208 ( n10503 , n3635 , n14277 );
    and g3209 ( n6432 , n10589 , n859 );
    or g3210 ( n11139 , n1741 , n3409 );
    not g3211 ( n7589 , n2354 );
    not g3212 ( n12197 , n13084 );
    or g3213 ( n11450 , n781 , n2215 );
    and g3214 ( n8119 , n9069 , n4314 );
    and g3215 ( n10673 , n1266 , n11626 );
    and g3216 ( n9755 , n11748 , n12344 );
    and g3217 ( n12296 , n12013 , n11845 );
    nor g3218 ( n731 , n12968 , n4118 );
    or g3219 ( n8766 , n77 , n4902 );
    and g3220 ( n3720 , n8431 , n7560 );
    and g3221 ( n4805 , n4095 , n7833 );
    or g3222 ( n1653 , n10224 , n13729 );
    and g3223 ( n7784 , n2998 , n5878 );
    and g3224 ( n10900 , n3736 , n13195 );
    not g3225 ( n10314 , n1769 );
    or g3226 ( n3318 , n1623 , n535 );
    or g3227 ( n8905 , n13155 , n1607 );
    and g3228 ( n12945 , n4657 , n1597 );
    and g3229 ( n13382 , n14358 , n5443 );
    or g3230 ( n8446 , n6256 , n6946 );
    not g3231 ( n8714 , n7322 );
    or g3232 ( n10325 , n8015 , n7020 );
    and g3233 ( n12454 , n7852 , n13889 );
    or g3234 ( n4515 , n4382 , n4117 );
    or g3235 ( n10127 , n10539 , n7338 );
    and g3236 ( n1544 , n11384 , n12310 );
    nor g3237 ( n602 , n1838 , n12513 );
    not g3238 ( n4415 , n8223 );
    and g3239 ( n13649 , n231 , n12770 );
    and g3240 ( n2667 , n1193 , n4494 );
    and g3241 ( n11557 , n9188 , n4487 );
    nor g3242 ( n10355 , n8487 , n6368 );
    and g3243 ( n14278 , n13227 , n2591 );
    and g3244 ( n148 , n12229 , n13532 );
    nor g3245 ( n12008 , n7227 , n9137 );
    or g3246 ( n2253 , n11105 , n14299 );
    or g3247 ( n1654 , n3569 , n6101 );
    or g3248 ( n130 , n1031 , n9074 );
    nor g3249 ( n8464 , n2875 , n7617 );
    and g3250 ( n14394 , n8393 , n9382 );
    nor g3251 ( n10347 , n6888 , n3863 );
    and g3252 ( n7616 , n8412 , n4947 );
    not g3253 ( n1147 , n2934 );
    not g3254 ( n541 , n8650 );
    and g3255 ( n5530 , n10622 , n3013 );
    not g3256 ( n11495 , n14525 );
    not g3257 ( n6157 , n5427 );
    nor g3258 ( n8360 , n8209 , n9875 );
    not g3259 ( n10241 , n5788 );
    or g3260 ( n6611 , n4065 , n587 );
    not g3261 ( n12992 , n2615 );
    or g3262 ( n12360 , n14481 , n8664 );
    and g3263 ( n884 , n13224 , n5860 );
    and g3264 ( n13402 , n8401 , n6283 );
    not g3265 ( n5018 , n5921 );
    or g3266 ( n11719 , n10913 , n11250 );
    and g3267 ( n9774 , n4574 , n1667 );
    nor g3268 ( n6440 , n4046 , n6028 );
    or g3269 ( n12329 , n5180 , n12442 );
    and g3270 ( n2403 , n8950 , n13610 );
    and g3271 ( n13179 , n13850 , n8844 );
    not g3272 ( n2919 , n381 );
    and g3273 ( n8841 , n12611 , n3627 );
    or g3274 ( n10450 , n283 , n5930 );
    nor g3275 ( n5361 , n1838 , n6512 );
    or g3276 ( n5284 , n2790 , n2148 );
    and g3277 ( n12561 , n4300 , n11869 );
    not g3278 ( n12131 , n6332 );
    and g3279 ( n6204 , n3370 , n10240 );
    or g3280 ( n2416 , n12401 , n1256 );
    not g3281 ( n3443 , n3812 );
    and g3282 ( n11099 , n3766 , n6214 );
    nor g3283 ( n5400 , n619 , n9066 );
    or g3284 ( n8403 , n6690 , n11127 );
    nor g3285 ( n2999 , n2742 , n7170 );
    or g3286 ( n246 , n7122 , n6885 );
    and g3287 ( n10697 , n7618 , n13819 );
    or g3288 ( n10544 , n8513 , n4612 );
    not g3289 ( n6700 , n13756 );
    or g3290 ( n1560 , n14449 , n7760 );
    or g3291 ( n3682 , n11123 , n6739 );
    nor g3292 ( n3899 , n2086 , n5724 );
    or g3293 ( n8731 , n10383 , n8974 );
    and g3294 ( n7184 , n8450 , n2963 );
    not g3295 ( n4908 , n7064 );
    and g3296 ( n1466 , n11406 , n3860 );
    and g3297 ( n3231 , n783 , n1695 );
    not g3298 ( n9740 , n1417 );
    and g3299 ( n567 , n13433 , n8928 );
    or g3300 ( n7058 , n6109 , n8711 );
    and g3301 ( n1397 , n12425 , n5201 );
    or g3302 ( n6535 , n14029 , n12945 );
    not g3303 ( n6765 , n1984 );
    or g3304 ( n992 , n5315 , n7348 );
    and g3305 ( n2609 , n4320 , n13682 );
    or g3306 ( n5547 , n10834 , n4805 );
    not g3307 ( n2149 , n3284 );
    and g3308 ( n3483 , n4803 , n1541 );
    or g3309 ( n11901 , n271 , n3367 );
    and g3310 ( n3648 , n9345 , n3968 );
    not g3311 ( n13435 , n4415 );
    and g3312 ( n6367 , n1354 , n12547 );
    or g3313 ( n10100 , n194 , n12661 );
    nor g3314 ( n6751 , n1812 , n13585 );
    or g3315 ( n11907 , n11183 , n11552 );
    not g3316 ( n448 , n7258 );
    not g3317 ( n85 , n1894 );
    and g3318 ( n9605 , n9188 , n10683 );
    not g3319 ( n9705 , n10376 );
    and g3320 ( n13828 , n4880 , n9708 );
    not g3321 ( n3169 , n9592 );
    and g3322 ( n11124 , n8232 , n8125 );
    and g3323 ( n5922 , n10909 , n10832 );
    and g3324 ( n3573 , n1937 , n6801 );
    and g3325 ( n10906 , n10909 , n3108 );
    or g3326 ( n5445 , n11231 , n12856 );
    and g3327 ( n6445 , n2682 , n11091 );
    and g3328 ( n1739 , n12336 , n9432 );
    and g3329 ( n4262 , n9705 , n10795 );
    and g3330 ( n5709 , n6724 , n8435 );
    and g3331 ( n13725 , n5640 , n3760 );
    not g3332 ( n3212 , n1478 );
    nor g3333 ( n6404 , n10136 , n3934 );
    or g3334 ( n13431 , n6471 , n14473 );
    and g3335 ( n1123 , n6609 , n966 );
    and g3336 ( n10718 , n6649 , n825 );
    and g3337 ( n14431 , n10562 , n4945 );
    not g3338 ( n13723 , n1938 );
    and g3339 ( n3412 , n13626 , n8240 );
    not g3340 ( n5715 , n6332 );
    and g3341 ( n12277 , n11240 , n8962 );
    nor g3342 ( n491 , n573 , n8688 );
    or g3343 ( n12799 , n185 , n6987 );
    and g3344 ( n13732 , n6527 , n10098 );
    or g3345 ( n476 , n3427 , n4248 );
    and g3346 ( n6642 , n6854 , n10914 );
    and g3347 ( n91 , n3833 , n12664 );
    or g3348 ( n8234 , n2761 , n10724 );
    and g3349 ( n2568 , n14063 , n8053 );
    not g3350 ( n8490 , n10204 );
    and g3351 ( n4440 , n9345 , n3550 );
    nor g3352 ( n7072 , n6743 , n6228 );
    or g3353 ( n13635 , n12047 , n813 );
    or g3354 ( n9983 , n1061 , n9128 );
    or g3355 ( n7828 , n13108 , n3117 );
    nor g3356 ( n7955 , n4742 , n12028 );
    and g3357 ( n9919 , n13860 , n13689 );
    and g3358 ( n1167 , n13555 , n2306 );
    or g3359 ( n11057 , n4899 , n255 );
    or g3360 ( n9182 , n13968 , n11605 );
    nor g3361 ( n2541 , n11980 , n2118 );
    or g3362 ( n375 , n10449 , n5985 );
    or g3363 ( n44 , n12047 , n9943 );
    or g3364 ( n2501 , n8172 , n6061 );
    or g3365 ( n13043 , n9507 , n1098 );
    and g3366 ( n6450 , n7421 , n8014 );
    and g3367 ( n12733 , n13755 , n9892 );
    or g3368 ( n13117 , n2149 , n10796 );
    and g3369 ( n2718 , n4692 , n1295 );
    and g3370 ( n13025 , n7943 , n4155 );
    not g3371 ( n405 , n5613 );
    nor g3372 ( n10938 , n5278 , n4307 );
    or g3373 ( n11834 , n11710 , n9773 );
    and g3374 ( n7699 , n776 , n14304 );
    and g3375 ( n2710 , n2367 , n14459 );
    not g3376 ( n7004 , n8163 );
    and g3377 ( n11976 , n13484 , n4767 );
    or g3378 ( n14471 , n7684 , n13796 );
    and g3379 ( n3850 , n14213 , n9945 );
    and g3380 ( n11357 , n98 , n2386 );
    and g3381 ( n3548 , n7961 , n5636 );
    not g3382 ( n9546 , n8903 );
    and g3383 ( n1010 , n3442 , n11129 );
    and g3384 ( n4752 , n9198 , n3307 );
    or g3385 ( n13659 , n10824 , n3822 );
    and g3386 ( n1320 , n12521 , n3258 );
    nor g3387 ( n10321 , n1844 , n12923 );
    and g3388 ( n13695 , n1414 , n8200 );
    and g3389 ( n9017 , n11688 , n4311 );
    and g3390 ( n1898 , n13656 , n12368 );
    not g3391 ( n2005 , n4906 );
    or g3392 ( n2088 , n2901 , n12958 );
    not g3393 ( n13087 , n1045 );
    and g3394 ( n10686 , n12741 , n4861 );
    or g3395 ( n8391 , n7803 , n5090 );
    or g3396 ( n3819 , n3871 , n6049 );
    and g3397 ( n6429 , n1428 , n13281 );
    or g3398 ( n12479 , n12759 , n7456 );
    and g3399 ( n9910 , n7392 , n1048 );
    and g3400 ( n9105 , n12521 , n3053 );
    or g3401 ( n1923 , n3219 , n1794 );
    and g3402 ( n9131 , n1427 , n5322 );
    nor g3403 ( n9630 , n10593 , n6132 );
    and g3404 ( n1573 , n1662 , n7924 );
    or g3405 ( n10962 , n5450 , n1943 );
    or g3406 ( n5320 , n77 , n5246 );
    not g3407 ( n3093 , n6804 );
    not g3408 ( n2744 , n5151 );
    or g3409 ( n6379 , n511 , n6617 );
    not g3410 ( n9229 , n7289 );
    nor g3411 ( n12766 , n4464 , n3278 );
    and g3412 ( n13319 , n4098 , n4232 );
    and g3413 ( n2336 , n9052 , n801 );
    and g3414 ( n9063 , n13525 , n7753 );
    or g3415 ( n6756 , n13847 , n8282 );
    and g3416 ( n13966 , n4901 , n2448 );
    or g3417 ( n12382 , n12414 , n4555 );
    or g3418 ( n870 , n5362 , n688 );
    or g3419 ( n8781 , n14430 , n13166 );
    not g3420 ( n10620 , n7007 );
    nor g3421 ( n12627 , n12727 , n14123 );
    or g3422 ( n5526 , n13518 , n5674 );
    and g3423 ( n7134 , n8849 , n4857 );
    and g3424 ( n8177 , n12592 , n3626 );
    not g3425 ( n2089 , n6332 );
    and g3426 ( n7336 , n957 , n8975 );
    not g3427 ( n3125 , n11308 );
    or g3428 ( n4043 , n10035 , n11556 );
    and g3429 ( n184 , n14321 , n5846 );
    not g3430 ( n4033 , n9596 );
    and g3431 ( n5539 , n11495 , n822 );
    not g3432 ( n14481 , n11456 );
    not g3433 ( n2025 , n3046 );
    and g3434 ( n14289 , n14303 , n6630 );
    and g3435 ( n3961 , n79 , n4428 );
    and g3436 ( n2855 , n7911 , n7723 );
    or g3437 ( n1077 , n850 , n940 );
    or g3438 ( n1380 , n568 , n14171 );
    and g3439 ( n13264 , n3401 , n11640 );
    not g3440 ( n9297 , n12450 );
    not g3441 ( n727 , n11793 );
    nor g3442 ( n2420 , n10568 , n1765 );
    and g3443 ( n623 , n5312 , n3596 );
    nor g3444 ( n9907 , n2566 , n9065 );
    or g3445 ( n11879 , n13118 , n9748 );
    or g3446 ( n4860 , n5064 , n8035 );
    and g3447 ( n13135 , n1361 , n9138 );
    and g3448 ( n6865 , n2006 , n10881 );
    and g3449 ( n12230 , n9824 , n11297 );
    and g3450 ( n9627 , n11300 , n1248 );
    not g3451 ( n8964 , n12444 );
    and g3452 ( n4789 , n1857 , n934 );
    nor g3453 ( n13526 , n14455 , n5058 );
    or g3454 ( n4151 , n4821 , n5344 );
    nor g3455 ( n14254 , n6603 , n9611 );
    or g3456 ( n10118 , n2694 , n4679 );
    and g3457 ( n14132 , n13676 , n824 );
    not g3458 ( n3444 , n11052 );
    and g3459 ( n8046 , n10166 , n13014 );
    and g3460 ( n6991 , n5899 , n14499 );
    and g3461 ( n10758 , n12721 , n10352 );
    and g3462 ( n5845 , n8238 , n996 );
    and g3463 ( n9908 , n6899 , n1679 );
    or g3464 ( n11065 , n2790 , n12220 );
    and g3465 ( n9237 , n12335 , n1981 );
    and g3466 ( n12123 , n11220 , n9311 );
    and g3467 ( n6234 , n7208 , n12524 );
    not g3468 ( n7902 , n8903 );
    and g3469 ( n13913 , n5926 , n8858 );
    not g3470 ( n5569 , n1060 );
    and g3471 ( n8763 , n5062 , n10707 );
    not g3472 ( n3895 , n3799 );
    nor g3473 ( n9390 , n5762 , n558 );
    not g3474 ( n3333 , n14512 );
    or g3475 ( n11843 , n2901 , n13375 );
    or g3476 ( n7489 , n11223 , n3764 );
    or g3477 ( n8779 , n11097 , n11043 );
    or g3478 ( n6834 , n2750 , n11908 );
    and g3479 ( n14463 , n11776 , n3450 );
    or g3480 ( n9311 , n7436 , n13904 );
    not g3481 ( n9236 , n3428 );
    or g3482 ( n9532 , n12112 , n9910 );
    and g3483 ( n3807 , n12960 , n12201 );
    and g3484 ( n8 , n13509 , n1714 );
    not g3485 ( n2583 , n12930 );
    and g3486 ( n12183 , n12858 , n690 );
    and g3487 ( n5968 , n12404 , n13605 );
    nor g3488 ( n6365 , n8404 , n11116 );
    and g3489 ( n981 , n3370 , n571 );
    and g3490 ( n6579 , n12147 , n2605 );
    or g3491 ( n10757 , n8714 , n12459 );
    not g3492 ( n1425 , n12846 );
    or g3493 ( n6409 , n5084 , n10628 );
    and g3494 ( n72 , n8393 , n1700 );
    and g3495 ( n9064 , n5279 , n8469 );
    and g3496 ( n11 , n10760 , n7309 );
    and g3497 ( n5455 , n11403 , n7048 );
    and g3498 ( n6015 , n4655 , n3953 );
    or g3499 ( n548 , n5548 , n6879 );
    and g3500 ( n13020 , n7677 , n376 );
    and g3501 ( n8564 , n6625 , n5477 );
    and g3502 ( n9152 , n98 , n5658 );
    not g3503 ( n10936 , n3284 );
    and g3504 ( n9104 , n533 , n12452 );
    not g3505 ( n5252 , n5606 );
    not g3506 ( n8655 , n6436 );
    or g3507 ( n9486 , n7156 , n10657 );
    and g3508 ( n10972 , n7529 , n5713 );
    or g3509 ( n861 , n12576 , n1521 );
    or g3510 ( n10517 , n5807 , n11200 );
    or g3511 ( n11247 , n5833 , n3644 );
    or g3512 ( n11775 , n5234 , n2667 );
    and g3513 ( n1689 , n14120 , n13662 );
    and g3514 ( n12398 , n7443 , n11348 );
    not g3515 ( n12023 , n12331 );
    or g3516 ( n8870 , n185 , n3368 );
    or g3517 ( n13044 , n2888 , n6177 );
    nor g3518 ( n8143 , n7200 , n13551 );
    or g3519 ( n12305 , n283 , n10780 );
    or g3520 ( n2649 , n8748 , n12959 );
    and g3521 ( n6980 , n541 , n14349 );
    not g3522 ( n3845 , n7822 );
    or g3523 ( n11297 , n504 , n3029 );
    not g3524 ( n9176 , n10358 );
    nor g3525 ( n1527 , n9563 , n12390 );
    or g3526 ( n1644 , n10713 , n2141 );
    not g3527 ( n10234 , n7875 );
    nor g3528 ( n1180 , n12673 , n9737 );
    and g3529 ( n3408 , n7327 , n4153 );
    not g3530 ( n3986 , n5618 );
    and g3531 ( n9040 , n10458 , n13411 );
    and g3532 ( n4628 , n12592 , n12371 );
    not g3533 ( n7759 , n12924 );
    not g3534 ( n10566 , n355 );
    nor g3535 ( n9090 , n4213 , n12966 );
    or g3536 ( n12599 , n14400 , n3293 );
    nor g3537 ( n5728 , n12827 , n4256 );
    or g3538 ( n2 , n9230 , n2519 );
    and g3539 ( n14146 , n12542 , n13549 );
    not g3540 ( n1031 , n11308 );
    or g3541 ( n3960 , n251 , n988 );
    and g3542 ( n7896 , n6606 , n11815 );
    or g3543 ( n8916 , n12500 , n1497 );
    and g3544 ( n3704 , n7216 , n9654 );
    and g3545 ( n8310 , n2177 , n7829 );
    or g3546 ( n9887 , n12414 , n5531 );
    or g3547 ( n3102 , n11621 , n12931 );
    nor g3548 ( n8359 , n8529 , n8633 );
    and g3549 ( n2294 , n10922 , n11891 );
    or g3550 ( n10911 , n12131 , n7237 );
    nor g3551 ( n13842 , n8576 , n5183 );
    or g3552 ( n7522 , n3126 , n6201 );
    and g3553 ( n9457 , n5876 , n11652 );
    or g3554 ( n1932 , n10248 , n13561 );
    or g3555 ( n5896 , n11839 , n10979 );
    not g3556 ( n13979 , n11350 );
    or g3557 ( n11860 , n5800 , n5307 );
    and g3558 ( n4769 , n8975 , n1640 );
    and g3559 ( n6377 , n6318 , n4922 );
    or g3560 ( n7406 , n2111 , n11920 );
    nor g3561 ( n13238 , n2218 , n3101 );
    and g3562 ( n3539 , n10668 , n9843 );
    not g3563 ( n2080 , n7748 );
    not g3564 ( n12191 , n10406 );
    not g3565 ( n14321 , n9583 );
    nor g3566 ( n7638 , n9743 , n6057 );
    and g3567 ( n2940 , n12185 , n10618 );
    not g3568 ( n10461 , n4203 );
    or g3569 ( n13346 , n12968 , n14285 );
    or g3570 ( n7468 , n12047 , n7550 );
    and g3571 ( n7800 , n14358 , n13925 );
    or g3572 ( n5350 , n3164 , n1182 );
    and g3573 ( n3983 , n533 , n9692 );
    or g3574 ( n3545 , n8607 , n3457 );
    not g3575 ( n6397 , n12675 );
    nor g3576 ( n4463 , n3445 , n13085 );
    nor g3577 ( n13519 , n6020 , n6972 );
    not g3578 ( n7221 , n2932 );
    and g3579 ( n10485 , n9803 , n7879 );
    or g3580 ( n1507 , n3527 , n11225 );
    and g3581 ( n10048 , n2783 , n1870 );
    and g3582 ( n6859 , n873 , n6261 );
    or g3583 ( n1556 , n13706 , n10107 );
    or g3584 ( n11974 , n14366 , n6585 );
    or g3585 ( n56 , n10953 , n11961 );
    or g3586 ( n6490 , n4180 , n8945 );
    or g3587 ( n4038 , n8877 , n7296 );
    and g3588 ( n12490 , n1481 , n8093 );
    not g3589 ( n12421 , n3361 );
    or g3590 ( n11815 , n4340 , n5360 );
    and g3591 ( n10219 , n636 , n723 );
    and g3592 ( n486 , n6753 , n12082 );
    or g3593 ( n2595 , n5409 , n2654 );
    and g3594 ( n6207 , n1708 , n616 );
    nor g3595 ( n13011 , n5042 , n2395 );
    or g3596 ( n37 , n5454 , n11132 );
    or g3597 ( n3382 , n5507 , n785 );
    and g3598 ( n13106 , n706 , n2994 );
    or g3599 ( n7037 , n10539 , n7511 );
    nor g3600 ( n11505 , n3871 , n9690 );
    not g3601 ( n5732 , n9354 );
    or g3602 ( n4750 , n14404 , n12797 );
    and g3603 ( n4478 , n10229 , n7873 );
    and g3604 ( n11991 , n14446 , n132 );
    or g3605 ( n3579 , n13413 , n2555 );
    or g3606 ( n8416 , n10191 , n14287 );
    and g3607 ( n10603 , n9673 , n379 );
    and g3608 ( n11194 , n9885 , n729 );
    nor g3609 ( n7962 , n10254 , n1615 );
    and g3610 ( n4841 , n4790 , n11775 );
    and g3611 ( n2576 , n986 , n1883 );
    or g3612 ( n5248 , n2017 , n7315 );
    nor g3613 ( n5112 , n9107 , n9658 );
    and g3614 ( n5384 , n10822 , n3044 );
    and g3615 ( n2962 , n2682 , n13192 );
    not g3616 ( n2571 , n12102 );
    and g3617 ( n14234 , n13525 , n4286 );
    nor g3618 ( n2312 , n14370 , n2024 );
    not g3619 ( n6044 , n359 );
    not g3620 ( n9404 , n10714 );
    and g3621 ( n991 , n4445 , n12602 );
    and g3622 ( n3409 , n8769 , n1306 );
    and g3623 ( n9943 , n13656 , n10267 );
    nor g3624 ( n3413 , n4988 , n4808 );
    and g3625 ( n11563 , n11702 , n8958 );
    not g3626 ( n1582 , n6357 );
    or g3627 ( n12031 , n6471 , n9568 );
    not g3628 ( n10248 , n8737 );
    and g3629 ( n714 , n10589 , n3808 );
    and g3630 ( n8029 , n14465 , n9800 );
    or g3631 ( n4191 , n3164 , n9664 );
    or g3632 ( n10146 , n3168 , n13233 );
    and g3633 ( n12875 , n7079 , n13196 );
    and g3634 ( n12318 , n5999 , n10919 );
    not g3635 ( n5412 , n8647 );
    and g3636 ( n10093 , n8401 , n7493 );
    not g3637 ( n12149 , n8735 );
    or g3638 ( n8200 , n2686 , n16 );
    or g3639 ( n11869 , n11438 , n13173 );
    not g3640 ( n8572 , n13458 );
    and g3641 ( n8960 , n12475 , n1653 );
    and g3642 ( n13171 , n12953 , n2817 );
    or g3643 ( n11600 , n10933 , n13189 );
    and g3644 ( n9060 , n11838 , n13817 );
    or g3645 ( n2279 , n11011 , n10196 );
    nor g3646 ( n1869 , n13979 , n7035 );
    or g3647 ( n9674 , n8476 , n14375 );
    or g3648 ( n13199 , n12400 , n10135 );
    or g3649 ( n3515 , n2784 , n9826 );
    and g3650 ( n2637 , n12542 , n8445 );
    or g3651 ( n5078 , n1202 , n13223 );
    or g3652 ( n11982 , n9218 , n13020 );
    or g3653 ( n118 , n850 , n9530 );
    not g3654 ( n183 , n8179 );
    nor g3655 ( n10719 , n12957 , n13829 );
    or g3656 ( n13754 , n13774 , n10339 );
    and g3657 ( n6571 , n6899 , n13887 );
    and g3658 ( n9157 , n10969 , n4522 );
    nor g3659 ( n206 , n9291 , n1806 );
    and g3660 ( n6479 , n7081 , n13199 );
    or g3661 ( n6299 , n10191 , n6029 );
    or g3662 ( n11497 , n4913 , n6302 );
    and g3663 ( n10592 , n11950 , n8830 );
    not g3664 ( n4682 , n8341 );
    or g3665 ( n223 , n11576 , n2962 );
    or g3666 ( n5510 , n7219 , n1956 );
    or g3667 ( n6175 , n8964 , n2394 );
    and g3668 ( n2038 , n13952 , n12726 );
    or g3669 ( n8251 , n7898 , n3353 );
    or g3670 ( n11918 , n8452 , n8520 );
    or g3671 ( n12 , n11510 , n12349 );
    not g3672 ( n10072 , n9950 );
    nor g3673 ( n2014 , n5488 , n2418 );
    nor g3674 ( n7669 , n12079 , n843 );
    and g3675 ( n744 , n1855 , n9317 );
    or g3676 ( n4697 , n13537 , n11015 );
    and g3677 ( n11141 , n7768 , n5285 );
    and g3678 ( n3681 , n1365 , n9214 );
    and g3679 ( n6441 , n10357 , n2238 );
    and g3680 ( n8995 , n4394 , n3832 );
    and g3681 ( n12477 , n4806 , n14054 );
    and g3682 ( n12940 , n13850 , n1961 );
    not g3683 ( n13707 , n3616 );
    nor g3684 ( n6416 , n12292 , n6194 );
    nor g3685 ( n11439 , n6074 , n2475 );
    or g3686 ( n10052 , n11123 , n14522 );
    or g3687 ( n10333 , n10245 , n12833 );
    or g3688 ( n4872 , n492 , n14203 );
    or g3689 ( n9775 , n9742 , n6002 );
    and g3690 ( n11465 , n1140 , n1912 );
    and g3691 ( n6396 , n10015 , n11239 );
    or g3692 ( n10839 , n5603 , n9816 );
    or g3693 ( n10149 , n12870 , n211 );
    not g3694 ( n1576 , n11541 );
    and g3695 ( n6631 , n7081 , n3984 );
    and g3696 ( n1204 , n7392 , n6497 );
    or g3697 ( n13936 , n1613 , n14407 );
    and g3698 ( n5091 , n457 , n1532 );
    and g3699 ( n10879 , n1074 , n11871 );
    or g3700 ( n13653 , n2387 , n4977 );
    or g3701 ( n13691 , n5625 , n8778 );
    and g3702 ( n7967 , n10374 , n13349 );
    not g3703 ( n5188 , n6258 );
    or g3704 ( n12201 , n3320 , n6713 );
    and g3705 ( n1300 , n2669 , n11985 );
    or g3706 ( n8309 , n3736 , n6999 );
    or g3707 ( n8542 , n9806 , n6239 );
    not g3708 ( n2677 , n11066 );
    or g3709 ( n13927 , n2236 , n281 );
    or g3710 ( n875 , n12633 , n1650 );
    or g3711 ( n11963 , n6263 , n3543 );
    or g3712 ( n6344 , n10508 , n10201 );
    and g3713 ( n948 , n2674 , n10462 );
    or g3714 ( n10086 , n4791 , n5629 );
    or g3715 ( n4356 , n1805 , n7916 );
    or g3716 ( n8125 , n11171 , n337 );
    not g3717 ( n647 , n12331 );
    not g3718 ( n7203 , n7940 );
    and g3719 ( n13228 , n5489 , n1366 );
    or g3720 ( n13335 , n1875 , n12332 );
    or g3721 ( n221 , n11094 , n13487 );
    and g3722 ( n2826 , n9265 , n11287 );
    or g3723 ( n11110 , n5409 , n12466 );
    and g3724 ( n6222 , n3586 , n12707 );
    or g3725 ( n6080 , n9211 , n9809 );
    and g3726 ( n349 , n10922 , n4331 );
    or g3727 ( n11626 , n8332 , n11080 );
    and g3728 ( n12279 , n1401 , n957 );
    not g3729 ( n6016 , n4618 );
    and g3730 ( n3616 , n1109 , n2343 );
    or g3731 ( n1500 , n11438 , n8246 );
    not g3732 ( n6874 , n7023 );
    not g3733 ( n3521 , n9377 );
    nor g3734 ( n3170 , n5762 , n1426 );
    or g3735 ( n4995 , n4821 , n6378 );
    nor g3736 ( n11624 , n5432 , n12932 );
    or g3737 ( n7976 , n2897 , n6086 );
    or g3738 ( n13619 , n11472 , n1823 );
    and g3739 ( n9707 , n7068 , n13671 );
    not g3740 ( n10376 , n746 );
    nor g3741 ( n8939 , n5429 , n14136 );
    or g3742 ( n13884 , n5234 , n6940 );
    not g3743 ( n6020 , n7455 );
    or g3744 ( n2379 , n2878 , n11224 );
    or g3745 ( n3741 , n8517 , n70 );
    and g3746 ( n3384 , n7909 , n2501 );
    and g3747 ( n5586 , n8552 , n8547 );
    and g3748 ( n8224 , n10846 , n11291 );
    or g3749 ( n10467 , n7358 , n6818 );
    or g3750 ( n9041 , n7255 , n2573 );
    not g3751 ( n9742 , n13165 );
    and g3752 ( n8917 , n12092 , n13813 );
    or g3753 ( n9925 , n9422 , n14402 );
    and g3754 ( n9009 , n2486 , n3091 );
    nor g3755 ( n5536 , n6211 , n1319 );
    or g3756 ( n9082 , n5695 , n9084 );
    nor g3757 ( n1090 , n1383 , n14416 );
    or g3758 ( n9333 , n766 , n7640 );
    or g3759 ( n12540 , n8638 , n3383 );
    or g3760 ( n6775 , n11405 , n2812 );
    or g3761 ( n528 , n838 , n9330 );
    or g3762 ( n11693 , n817 , n967 );
    and g3763 ( n9624 , n3485 , n8684 );
    not g3764 ( n4618 , n11343 );
    or g3765 ( n3042 , n6711 , n534 );
    and g3766 ( n8167 , n4546 , n7899 );
    and g3767 ( n1373 , n8923 , n6811 );
    and g3768 ( n10937 , n10032 , n13355 );
    or g3769 ( n4158 , n6323 , n8181 );
    and g3770 ( n10135 , n8043 , n3390 );
    and g3771 ( n9826 , n12259 , n11754 );
    and g3772 ( n13303 , n5999 , n2326 );
    nor g3773 ( n10459 , n8065 , n13958 );
    and g3774 ( n9835 , n4486 , n5694 );
    or g3775 ( n10188 , n13485 , n3480 );
    or g3776 ( n7578 , n695 , n10541 );
    and g3777 ( n11740 , n1804 , n563 );
    or g3778 ( n3678 , n7812 , n1455 );
    and g3779 ( n2590 , n4554 , n9986 );
    or g3780 ( n846 , n11176 , n13397 );
    or g3781 ( n9973 , n5144 , n1930 );
    or g3782 ( n6923 , n3815 , n14012 );
    and g3783 ( n11322 , n10408 , n2732 );
    and g3784 ( n14218 , n3435 , n4024 );
    nor g3785 ( n1280 , n6062 , n2880 );
    nor g3786 ( n4542 , n10936 , n1839 );
    and g3787 ( n1756 , n428 , n8961 );
    and g3788 ( n6224 , n9345 , n5063 );
    or g3789 ( n9112 , n5575 , n3406 );
    or g3790 ( n13598 , n7212 , n4355 );
    and g3791 ( n5619 , n4156 , n4810 );
    and g3792 ( n4704 , n7798 , n10497 );
    or g3793 ( n2986 , n781 , n7157 );
    not g3794 ( n2597 , n8148 );
    and g3795 ( n7752 , n12475 , n6213 );
    and g3796 ( n10138 , n11020 , n9089 );
    not g3797 ( n4692 , n3443 );
    not g3798 ( n2709 , n1571 );
    and g3799 ( n11920 , n10134 , n640 );
    and g3800 ( n4885 , n5764 , n1815 );
    not g3801 ( n11951 , n3070 );
    or g3802 ( n5589 , n900 , n12868 );
    and g3803 ( n13309 , n13525 , n3778 );
    or g3804 ( n12484 , n584 , n10704 );
    and g3805 ( n1055 , n8769 , n12362 );
    and g3806 ( n429 , n9275 , n2056 );
    or g3807 ( n3135 , n492 , n8532 );
    and g3808 ( n12836 , n11636 , n2867 );
    and g3809 ( n13533 , n8427 , n4085 );
    or g3810 ( n11913 , n2645 , n9294 );
    and g3811 ( n7415 , n14120 , n2074 );
    or g3812 ( n4798 , n766 , n9267 );
    not g3813 ( n3559 , n1214 );
    and g3814 ( n1451 , n13359 , n2286 );
    or g3815 ( n7390 , n4447 , n5023 );
    not g3816 ( n11814 , n13038 );
    or g3817 ( n9843 , n12047 , n4548 );
    and g3818 ( n3499 , n8213 , n13635 );
    or g3819 ( n3689 , n10523 , n9938 );
    not g3820 ( n12673 , n7814 );
    nor g3821 ( n3226 , n478 , n453 );
    or g3822 ( n12510 , n10394 , n4271 );
    or g3823 ( n13611 , n2025 , n11102 );
    not g3824 ( n5486 , n3776 );
    nor g3825 ( n334 , n6085 , n5916 );
    and g3826 ( n4884 , n11313 , n11659 );
    not g3827 ( n10529 , n3344 );
    and g3828 ( n11463 , n13364 , n3217 );
    or g3829 ( n14233 , n12130 , n276 );
    and g3830 ( n4642 , n9564 , n10213 );
    and g3831 ( n5165 , n12101 , n11247 );
    and g3832 ( n12000 , n6130 , n9753 );
    and g3833 ( n1872 , n1662 , n5615 );
    and g3834 ( n6919 , n865 , n2342 );
    and g3835 ( n10682 , n6744 , n7897 );
    and g3836 ( n3695 , n13860 , n8562 );
    or g3837 ( n1039 , n234 , n10148 );
    and g3838 ( n7891 , n501 , n6533 );
    or g3839 ( n3307 , n5570 , n3339 );
    nor g3840 ( n352 , n5132 , n10709 );
    nor g3841 ( n651 , n1028 , n6715 );
    not g3842 ( n14178 , n11404 );
    or g3843 ( n4323 , n6857 , n7645 );
    and g3844 ( n13496 , n5628 , n3072 );
    or g3845 ( n9638 , n6596 , n6665 );
    not g3846 ( n9944 , n12930 );
    and g3847 ( n1753 , n6854 , n8924 );
    or g3848 ( n12645 , n9285 , n5245 );
    nor g3849 ( n12860 , n10323 , n1865 );
    and g3850 ( n7863 , n5335 , n13936 );
    nor g3851 ( n399 , n573 , n12492 );
    and g3852 ( n4902 , n13342 , n12479 );
    or g3853 ( n1643 , n11724 , n3451 );
    and g3854 ( n11541 , n7676 , n8341 );
    and g3855 ( n5604 , n7203 , n9358 );
    and g3856 ( n5447 , n7211 , n6950 );
    nor g3857 ( n4507 , n8527 , n8420 );
    and g3858 ( n5905 , n3222 , n13968 );
    and g3859 ( n204 , n1775 , n8570 );
    not g3860 ( n12324 , n4550 );
    or g3861 ( n9162 , n10191 , n635 );
    or g3862 ( n7029 , n9716 , n3140 );
    not g3863 ( n6730 , n81 );
    or g3864 ( n629 , n504 , n11416 );
    and g3865 ( n9381 , n8213 , n9048 );
    and g3866 ( n4328 , n11336 , n4936 );
    or g3867 ( n1512 , n839 , n11995 );
    and g3868 ( n11152 , n3976 , n8220 );
    or g3869 ( n1444 , n9230 , n6954 );
    and g3870 ( n874 , n13227 , n594 );
    or g3871 ( n5123 , n6288 , n5519 );
    and g3872 ( n6303 , n457 , n6547 );
    and g3873 ( n4004 , n9191 , n548 );
    nor g3874 ( n3372 , n5065 , n8180 );
    or g3875 ( n12017 , n9620 , n4893 );
    or g3876 ( n5683 , n11392 , n11854 );
    nor g3877 ( n68 , n11232 , n8762 );
    or g3878 ( n11746 , n4052 , n13876 );
    and g3879 ( n11381 , n13656 , n7872 );
    or g3880 ( n13756 , n3958 , n1265 );
    and g3881 ( n6666 , n12832 , n10315 );
    not g3882 ( n10973 , n637 );
    and g3883 ( n10268 , n808 , n6156 );
    and g3884 ( n1002 , n4614 , n11326 );
    and g3885 ( n5281 , n333 , n7408 );
    nor g3886 ( n9309 , n2086 , n7431 );
    not g3887 ( n2846 , n5435 );
    and g3888 ( n11064 , n10516 , n2977 );
    or g3889 ( n14349 , n13516 , n4389 );
    not g3890 ( n838 , n9169 );
    or g3891 ( n3782 , n6519 , n8156 );
    or g3892 ( n3599 , n4877 , n7414 );
    nor g3893 ( n12654 , n10309 , n11732 );
    or g3894 ( n2029 , n3222 , n8315 );
    nor g3895 ( n11427 , n1378 , n2390 );
    not g3896 ( n8337 , n3155 );
    or g3897 ( n13976 , n9747 , n1886 );
    or g3898 ( n9771 , n3886 , n2228 );
    or g3899 ( n5817 , n5472 , n9965 );
    not g3900 ( n10465 , n7660 );
    and g3901 ( n10410 , n4932 , n4683 );
    or g3902 ( n13581 , n2761 , n7751 );
    or g3903 ( n711 , n8575 , n12720 );
    not g3904 ( n9080 , n7662 );
    nor g3905 ( n4607 , n11047 , n708 );
    or g3906 ( n1433 , n9035 , n52 );
    not g3907 ( n14150 , n2417 );
    or g3908 ( n8055 , n6867 , n12386 );
    and g3909 ( n8293 , n8692 , n11149 );
    or g3910 ( n4934 , n8582 , n9460 );
    or g3911 ( n6967 , n8517 , n879 );
    or g3912 ( n4083 , n2877 , n11060 );
    or g3913 ( n14355 , n13501 , n6538 );
    or g3914 ( n3657 , n8490 , n4392 );
    not g3915 ( n7905 , n8631 );
    not g3916 ( n13860 , n3313 );
    and g3917 ( n9018 , n13755 , n10729 );
    or g3918 ( n12572 , n11362 , n5725 );
    and g3919 ( n9591 , n12013 , n59 );
    or g3920 ( n9746 , n10913 , n6540 );
    and g3921 ( n9317 , n8376 , n3113 );
    and g3922 ( n3299 , n11300 , n9341 );
    nor g3923 ( n5827 , n5715 , n5289 );
    and g3924 ( n336 , n13096 , n6334 );
    not g3925 ( n10784 , n3070 );
    or g3926 ( n6168 , n4898 , n8457 );
    nor g3927 ( n3621 , n7365 , n6345 );
    nor g3928 ( n4652 , n2932 , n665 );
    not g3929 ( n7187 , n11861 );
    and g3930 ( n4167 , n7026 , n1593 );
    nor g3931 ( n13637 , n9657 , n12911 );
    not g3932 ( n13002 , n4082 );
    not g3933 ( n3608 , n13000 );
    not g3934 ( n12019 , n12444 );
    or g3935 ( n1565 , n1834 , n14427 );
    and g3936 ( n8109 , n8605 , n12560 );
    and g3937 ( n10942 , n3743 , n13845 );
    or g3938 ( n2890 , n5647 , n11408 );
    or g3939 ( n3790 , n1006 , n2294 );
    or g3940 ( n2754 , n1147 , n8005 );
    and g3941 ( n1227 , n5764 , n12164 );
    and g3942 ( n9997 , n8043 , n7399 );
    not g3943 ( n2533 , n8122 );
    and g3944 ( n1655 , n6013 , n9973 );
    or g3945 ( n12544 , n11183 , n8632 );
    not g3946 ( n7249 , n10889 );
    nor g3947 ( n5676 , n4491 , n792 );
    not g3948 ( n7818 , n11590 );
    and g3949 ( n7877 , n9944 , n1574 );
    and g3950 ( n6012 , n5225 , n11987 );
    and g3951 ( n10727 , n12998 , n10740 );
    not g3952 ( n11722 , n12776 );
    or g3953 ( n572 , n100 , n2975 );
    and g3954 ( n942 , n9898 , n10491 );
    or g3955 ( n9954 , n9078 , n10228 );
    or g3956 ( n8299 , n7700 , n5790 );
    and g3957 ( n7144 , n13464 , n6297 );
    and g3958 ( n4712 , n1588 , n6543 );
    or g3959 ( n2772 , n6498 , n5430 );
    nor g3960 ( n5735 , n11047 , n5915 );
    and g3961 ( n12704 , n4803 , n6535 );
    or g3962 ( n13943 , n8969 , n8646 );
    nor g3963 ( n13939 , n4988 , n1822 );
    and g3964 ( n4586 , n4574 , n8285 );
    not g3965 ( n3635 , n5675 );
    or g3966 ( n305 , n5548 , n6361 );
    or g3967 ( n669 , n5710 , n5308 );
    not g3968 ( n11302 , n13981 );
    or g3969 ( n14326 , n2091 , n11590 );
    not g3970 ( n4464 , n1076 );
    or g3971 ( n2938 , n8209 , n4613 );
    or g3972 ( n9424 , n695 , n4440 );
    and g3973 ( n5290 , n6157 , n8202 );
    and g3974 ( n12841 , n13246 , n10677 );
    not g3975 ( n7670 , n1495 );
    not g3976 ( n14512 , n6765 );
    not g3977 ( n9456 , n4324 );
    or g3978 ( n7294 , n13518 , n9334 );
    and g3979 ( n10175 , n9015 , n10451 );
    and g3980 ( n4228 , n13078 , n13623 );
    and g3981 ( n6281 , n706 , n8956 );
    nor g3982 ( n10495 , n4105 , n857 );
    not g3983 ( n6196 , n1771 );
    not g3984 ( n9780 , n7875 );
    not g3985 ( n5365 , n670 );
    and g3986 ( n6645 , n7767 , n6789 );
    or g3987 ( n4714 , n2686 , n2528 );
    or g3988 ( n6530 , n5236 , n9016 );
    not g3989 ( n12531 , n6559 );
    or g3990 ( n13705 , n3394 , n13871 );
    and g3991 ( n6686 , n2082 , n621 );
    and g3992 ( n5561 , n889 , n8636 );
    or g3993 ( n8340 , n4498 , n14207 );
    or g3994 ( n13801 , n11315 , n8948 );
    not g3995 ( n4134 , n7754 );
    or g3996 ( n2147 , n4233 , n8591 );
    not g3997 ( n4923 , n9596 );
    and g3998 ( n5560 , n6531 , n12556 );
    or g3999 ( n4155 , n10781 , n11160 );
    and g4000 ( n11426 , n9941 , n459 );
    and g4001 ( n836 , n5553 , n5189 );
    nor g4002 ( n13709 , n4233 , n1627 );
    or g4003 ( n6508 , n9269 , n1549 );
    not g4004 ( n8620 , n5601 );
    or g4005 ( n3788 , n11739 , n1353 );
    and g4006 ( n354 , n12461 , n3102 );
    and g4007 ( n8326 , n11495 , n6437 );
    not g4008 ( n6111 , n2320 );
    and g4009 ( n12848 , n4347 , n10286 );
    and g4010 ( n2347 , n3097 , n7515 );
    not g4011 ( n7229 , n628 );
    and g4012 ( n2011 , n10025 , n2611 );
    or g4013 ( n8562 , n6205 , n7923 );
    nor g4014 ( n7403 , n9529 , n6075 );
    or g4015 ( n11059 , n3273 , n13073 );
    or g4016 ( n487 , n7912 , n1980 );
    not g4017 ( n673 , n10255 );
    or g4018 ( n5678 , n1447 , n10283 );
    or g4019 ( n1746 , n8151 , n388 );
    or g4020 ( n9802 , n2412 , n10759 );
    not g4021 ( n1838 , n8735 );
    not g4022 ( n5475 , n5951 );
    nor g4023 ( n199 , n7448 , n8794 );
    not g4024 ( n14351 , n11668 );
    nor g4025 ( n3027 , n2009 , n3760 );
    or g4026 ( n632 , n9226 , n1533 );
    or g4027 ( n8243 , n4821 , n14218 );
    and g4028 ( n13010 , n10061 , n489 );
    and g4029 ( n9545 , n12445 , n3150 );
    nor g4030 ( n8551 , n4092 , n6790 );
    or g4031 ( n8699 , n6046 , n7583 );
    and g4032 ( n13008 , n13597 , n7173 );
    not g4033 ( n4199 , n13696 );
    and g4034 ( n5280 , n9069 , n12424 );
    and g4035 ( n12667 , n13781 , n3949 );
    and g4036 ( n10413 , n4554 , n4041 );
    not g4037 ( n12400 , n2934 );
    or g4038 ( n11170 , n12759 , n12516 );
    or g4039 ( n14322 , n11980 , n13778 );
    nor g4040 ( n7999 , n7519 , n7458 );
    or g4041 ( n1774 , n6205 , n14325 );
    or g4042 ( n7628 , n10351 , n8229 );
    or g4043 ( n14345 , n12820 , n14143 );
    and g4044 ( n12369 , n4844 , n1116 );
    and g4045 ( n11553 , n4880 , n13475 );
    not g4046 ( n636 , n4000 );
    not g4047 ( n2016 , n12746 );
    or g4048 ( n9199 , n13083 , n13798 );
    and g4049 ( n597 , n13433 , n10011 );
    not g4050 ( n1821 , n10108 );
    and g4051 ( n289 , n4546 , n4796 );
    or g4052 ( n963 , n11223 , n13309 );
    not g4053 ( n11804 , n5242 );
    not g4054 ( n3628 , n498 );
    nor g4055 ( n5747 , n1342 , n4917 );
    and g4056 ( n2557 , n533 , n973 );
    not g4057 ( n4932 , n1784 );
    or g4058 ( n4616 , n2089 , n6006 );
    or g4059 ( n1908 , n12779 , n977 );
    or g4060 ( n6485 , n1875 , n12610 );
    or g4061 ( n8225 , n9804 , n3514 );
    not g4062 ( n10469 , n10965 );
    not g4063 ( n2241 , n1311 );
    or g4064 ( n3525 , n7250 , n6915 );
    or g4065 ( n5835 , n1613 , n8167 );
    or g4066 ( n12134 , n89 , n9455 );
    or g4067 ( n1750 , n10449 , n13488 );
    not g4068 ( n3736 , n12218 );
    or g4069 ( n308 , n2531 , n13587 );
    and g4070 ( n8662 , n3435 , n4723 );
    and g4071 ( n13497 , n1354 , n5962 );
    and g4072 ( n7893 , n6649 , n9788 );
    and g4073 ( n8003 , n14074 , n11283 );
    and g4074 ( n4308 , n2724 , n7271 );
    and g4075 ( n14380 , n9323 , n9782 );
    and g4076 ( n11209 , n2527 , n1163 );
    or g4077 ( n3098 , n10784 , n5436 );
    nor g4078 ( n7725 , n8701 , n9436 );
    or g4079 ( n11166 , n8969 , n9904 );
    or g4080 ( n3558 , n6090 , n5386 );
    or g4081 ( n7434 , n5468 , n1952 );
    and g4082 ( n9932 , n11329 , n3589 );
    and g4083 ( n2319 , n4614 , n13388 );
    or g4084 ( n4331 , n11440 , n4316 );
    and g4085 ( n12623 , n3169 , n851 );
    or g4086 ( n1211 , n6891 , n11741 );
    or g4087 ( n9363 , n4508 , n8852 );
    not g4088 ( n12401 , n628 );
    and g4089 ( n11476 , n1610 , n2489 );
    nor g4090 ( n2574 , n10342 , n4259 );
    and g4091 ( n10366 , n1266 , n12406 );
    or g4092 ( n5263 , n11315 , n8559 );
    and g4093 ( n9530 , n10229 , n2253 );
    nor g4094 ( n3146 , n5715 , n4610 );
    and g4095 ( n9214 , n888 , n1401 );
    and g4096 ( n6761 , n9898 , n434 );
    not g4097 ( n9151 , n14154 );
    or g4098 ( n444 , n2387 , n10807 );
    nor g4099 ( n8269 , n12248 , n12348 );
    or g4100 ( n10884 , n7862 , n4350 );
    or g4101 ( n8469 , n6596 , n12841 );
    and g4102 ( n395 , n3715 , n10863 );
    and g4103 ( n4893 , n8007 , n5889 );
    and g4104 ( n6060 , n10229 , n8037 );
    or g4105 ( n2282 , n769 , n7454 );
    and g4106 ( n10600 , n5335 , n6219 );
    and g4107 ( n11763 , n494 , n12995 );
    not g4108 ( n5354 , n9967 );
    and g4109 ( n6101 , n13297 , n10467 );
    or g4110 ( n1810 , n1582 , n12181 );
    nor g4111 ( n6239 , n6679 , n6421 );
    and g4112 ( n10596 , n14109 , n6518 );
    nor g4113 ( n9088 , n13153 , n12347 );
    and g4114 ( n7906 , n392 , n6142 );
    or g4115 ( n11366 , n11036 , n1982 );
    or g4116 ( n3110 , n9151 , n12383 );
    or g4117 ( n3068 , n10929 , n12097 );
    not g4118 ( n2086 , n12444 );
    and g4119 ( n14328 , n10084 , n4017 );
    not g4120 ( n9657 , n10617 );
    not g4121 ( n6609 , n920 );
    or g4122 ( n10432 , n1391 , n39 );
    and g4123 ( n4991 , n7612 , n4704 );
    or g4124 ( n8639 , n11420 , n1488 );
    nor g4125 ( n903 , n9984 , n5718 );
    and g4126 ( n6954 , n9617 , n7910 );
    or g4127 ( n5707 , n2111 , n6913 );
    and g4128 ( n9938 , n8923 , n4914 );
    nor g4129 ( n7701 , n6905 , n3027 );
    not g4130 ( n3696 , n5221 );
    or g4131 ( n13915 , n10960 , n7312 );
    and g4132 ( n6393 , n11569 , n811 );
    not g4133 ( n12351 , n9878 );
    or g4134 ( n7085 , n10024 , n1618 );
    not g4135 ( n10358 , n4633 );
    nor g4136 ( n4705 , n1028 , n6613 );
    and g4137 ( n3504 , n14063 , n4707 );
    nor g4138 ( n6133 , n6971 , n11578 );
    nor g4139 ( n1257 , n194 , n7008 );
    or g4140 ( n6003 , n13276 , n13878 );
    or g4141 ( n8344 , n1613 , n10587 );
    and g4142 ( n4954 , n2904 , n1039 );
    or g4143 ( n1020 , n4602 , n6079 );
    and g4144 ( n13543 , n4104 , n13449 );
    and g4145 ( n11245 , n1254 , n13879 );
    nor g4146 ( n10528 , n14238 , n3906 );
    or g4147 ( n14231 , n5587 , n13674 );
    or g4148 ( n1386 , n7803 , n14493 );
    or g4149 ( n12157 , n12295 , n2832 );
    not g4150 ( n10767 , n12522 );
    not g4151 ( n2194 , n8631 );
    and g4152 ( n7077 , n7484 , n7502 );
    or g4153 ( n11884 , n4435 , n3499 );
    or g4154 ( n10081 , n8480 , n1528 );
    and g4155 ( n1749 , n9811 , n1102 );
    not g4156 ( n1202 , n7289 );
    or g4157 ( n8654 , n6373 , n10038 );
    and g4158 ( n1368 , n6051 , n3184 );
    nor g4159 ( n8504 , n5848 , n399 );
    or g4160 ( n3115 , n5480 , n9251 );
    or g4161 ( n800 , n1711 , n3983 );
    or g4162 ( n3881 , n1728 , n12928 );
    nor g4163 ( n299 , n5504 , n7340 );
    or g4164 ( n2316 , n5188 , n2334 );
    or g4165 ( n7096 , n8045 , n6273 );
    and g4166 ( n12795 , n9321 , n6469 );
    or g4167 ( n4999 , n4791 , n7831 );
    or g4168 ( n10585 , n3047 , n13463 );
    not g4169 ( n3492 , n2164 );
    and g4170 ( n2995 , n6697 , n1975 );
    not g4171 ( n5505 , n10099 );
    or g4172 ( n12426 , n10857 , n1157 );
    and g4173 ( n3975 , n11313 , n8075 );
    and g4174 ( n13710 , n9345 , n1499 );
    not g4175 ( n7888 , n11331 );
    and g4176 ( n9250 , n7693 , n12302 );
    or g4177 ( n1022 , n11584 , n9871 );
    or g4178 ( n1789 , n10784 , n9813 );
    or g4179 ( n4866 , n10808 , n10872 );
    and g4180 ( n6647 , n3435 , n4961 );
    or g4181 ( n9808 , n8964 , n5568 );
    and g4182 ( n6145 , n12202 , n983 );
    and g4183 ( n4874 , n13107 , n10316 );
    not g4184 ( n4300 , n10372 );
    and g4185 ( n4577 , n14313 , n10887 );
    or g4186 ( n1498 , n11804 , n7895 );
    or g4187 ( n7046 , n4562 , n5961 );
    nor g4188 ( n5915 , n3428 , n8086 );
    and g4189 ( n10665 , n3986 , n12157 );
    and g4190 ( n5375 , n4790 , n8171 );
    or g4191 ( n7083 , n13941 , n8709 );
    and g4192 ( n6563 , n13227 , n7666 );
    nor g4193 ( n12672 , n10289 , n5879 );
    or g4194 ( n8174 , n13142 , n6174 );
    and g4195 ( n834 , n12037 , n3879 );
    or g4196 ( n7554 , n11542 , n1169 );
    or g4197 ( n7753 , n13518 , n5399 );
    and g4198 ( n13859 , n1247 , n8355 );
    or g4199 ( n7682 , n11384 , n6147 );
    not g4200 ( n15 , n9563 );
    and g4201 ( n2214 , n13338 , n780 );
    or g4202 ( n11431 , n49 , n6220 );
    nor g4203 ( n244 , n9807 , n12330 );
    nor g4204 ( n3487 , n9567 , n5005 );
    nor g4205 ( n13894 , n5172 , n4651 );
    or g4206 ( n13468 , n3527 , n9897 );
    and g4207 ( n2492 , n12683 , n7099 );
    and g4208 ( n4177 , n12015 , n12215 );
    and g4209 ( n8218 , n10197 , n8501 );
    not g4210 ( n2644 , n2723 );
    nor g4211 ( n12637 , n9423 , n9506 );
    nor g4212 ( n3642 , n7920 , n4477 );
    and g4213 ( n9955 , n14157 , n7478 );
    or g4214 ( n3024 , n8458 , n12689 );
    and g4215 ( n2126 , n4895 , n3798 );
    or g4216 ( n3442 , n1705 , n11529 );
    nor g4217 ( n5527 , n3344 , n2769 );
    and g4218 ( n1282 , n13575 , n1177 );
    nor g4219 ( n6477 , n3871 , n2813 );
    or g4220 ( n14221 , n7245 , n6282 );
    or g4221 ( n10056 , n10781 , n4598 );
    and g4222 ( n1620 , n8232 , n9551 );
    or g4223 ( n1811 , n1697 , n5325 );
    and g4224 ( n11712 , n13407 , n1144 );
    and g4225 ( n8377 , n9321 , n5373 );
    not g4226 ( n1677 , n8884 );
    or g4227 ( n3641 , n6672 , n1017 );
    or g4228 ( n2231 , n9285 , n8599 );
    or g4229 ( n8623 , n648 , n6776 );
    nor g4230 ( n11946 , n13941 , n14300 );
    and g4231 ( n12332 , n11950 , n8757 );
    and g4232 ( n9971 , n12768 , n8868 );
    nor g4233 ( n4196 , n13675 , n5722 );
    and g4234 ( n8919 , n5012 , n11082 );
    not g4235 ( n12189 , n5288 );
    or g4236 ( n2755 , n3877 , n12074 );
    and g4237 ( n4385 , n12768 , n8537 );
    or g4238 ( n449 , n5575 , n3468 );
    not g4239 ( n10975 , n2202 );
    and g4240 ( n11009 , n6128 , n12426 );
    or g4241 ( n13119 , n2750 , n5405 );
    or g4242 ( n14211 , n12764 , n7059 );
    not g4243 ( n3344 , n5886 );
    and g4244 ( n1245 , n14313 , n7494 );
    and g4245 ( n4520 , n13404 , n2003 );
    or g4246 ( n12613 , n89 , n14396 );
    or g4247 ( n12411 , n13130 , n13391 );
    and g4248 ( n13673 , n12998 , n14288 );
    nor g4249 ( n8863 , n2780 , n7439 );
    or g4250 ( n14397 , n3569 , n11278 );
    or g4251 ( n13576 , n14404 , n3077 );
    or g4252 ( n4849 , n4435 , n9619 );
    not g4253 ( n12960 , n5852 );
    nor g4254 ( n7030 , n3870 , n8190 );
    or g4255 ( n1752 , n13226 , n626 );
    not g4256 ( n3370 , n5460 );
    not g4257 ( n5084 , n777 );
    nor g4258 ( n14476 , n2790 , n13839 );
    or g4259 ( n6843 , n12633 , n6542 );
    not g4260 ( n3268 , n3402 );
    and g4261 ( n11899 , n79 , n2704 );
    nor g4262 ( n12700 , n11558 , n7557 );
    and g4263 ( n4166 , n98 , n14027 );
    or g4264 ( n11130 , n7389 , n8997 );
    nor g4265 ( n14318 , n8189 , n2798 );
    or g4266 ( n340 , n69 , n9180 );
    not g4267 ( n14009 , n6147 );
    or g4268 ( n6989 , n9154 , n3833 );
    or g4269 ( n13092 , n11951 , n11539 );
    and g4270 ( n7237 , n898 , n5508 );
    and g4271 ( n6076 , n4803 , n13938 );
    or g4272 ( n13125 , n8983 , n14114 );
    or g4273 ( n1632 , n974 , n5729 );
    or g4274 ( n9789 , n13485 , n9625 );
    and g4275 ( n4590 , n2783 , n1738 );
    or g4276 ( n6568 , n6596 , n11317 );
    or g4277 ( n12659 , n2236 , n14436 );
    and g4278 ( n13594 , n13676 , n11821 );
    and g4279 ( n12160 , n4690 , n2375 );
    or g4280 ( n3476 , n6971 , n11723 );
    nor g4281 ( n8840 , n7551 , n2163 );
    and g4282 ( n4222 , n5823 , n252 );
    and g4283 ( n6617 , n8432 , n10127 );
    and g4284 ( n12750 , n1247 , n11138 );
    not g4285 ( n4267 , n13992 );
    or g4286 ( n3933 , n8986 , n11374 );
    and g4287 ( n726 , n3401 , n6435 );
    nor g4288 ( n430 , n10342 , n4086 );
    and g4289 ( n8931 , n5823 , n14420 );
    and g4290 ( n5821 , n5926 , n14491 );
    or g4291 ( n12343 , n8242 , n8644 );
    or g4292 ( n3989 , n2845 , n12142 );
    and g4293 ( n11013 , n9315 , n11177 );
    or g4294 ( n13786 , n10224 , n313 );
    not g4295 ( n4270 , n12409 );
    nor g4296 ( n5540 , n6426 , n2133 );
    or g4297 ( n3258 , n14366 , n4884 );
    or g4298 ( n6619 , n3569 , n2138 );
    and g4299 ( n4197 , n7627 , n11970 );
    not g4300 ( n14216 , n14365 );
    not g4301 ( n1051 , n918 );
    or g4302 ( n10066 , n13074 , n6043 );
    not g4303 ( n1638 , n5333 );
    nor g4304 ( n5824 , n13310 , n9732 );
    and g4305 ( n1352 , n11838 , n13384 );
    and g4306 ( n7117 , n12741 , n12382 );
    not g4307 ( n9804 , n8813 );
    and g4308 ( n11349 , n12542 , n6959 );
    nor g4309 ( n6141 , n2212 , n4766 );
    or g4310 ( n9725 , n12695 , n12071 );
    and g4311 ( n7931 , n8721 , n2193 );
    nor g4312 ( n4383 , n13522 , n2312 );
    and g4313 ( n7959 , n9265 , n6230 );
    or g4314 ( n641 , n5454 , n8859 );
    and g4315 ( n7348 , n12250 , n3074 );
    and g4316 ( n3543 , n7043 , n150 );
    and g4317 ( n5047 , n222 , n12724 );
    or g4318 ( n10756 , n9742 , n6065 );
    and g4319 ( n5367 , n776 , n2231 );
    nor g4320 ( n14117 , n4200 , n11910 );
    nor g4321 ( n5649 , n8277 , n9841 );
    or g4322 ( n13143 , n1494 , n7893 );
    or g4323 ( n12951 , n14481 , n7958 );
    or g4324 ( n5677 , n9226 , n14380 );
    or g4325 ( n1939 , n2055 , n6993 );
    and g4326 ( n2141 , n1772 , n4931 );
    or g4327 ( n7517 , n1261 , n4845 );
    nor g4328 ( n1319 , n8527 , n4836 );
    not g4329 ( n6744 , n10828 );
    not g4330 ( n8752 , n11617 );
    not g4331 ( n2953 , n6067 );
    and g4332 ( n7707 , n7060 , n9394 );
    nor g4333 ( n11056 , n7418 , n4396 );
    and g4334 ( n11940 , n9617 , n13250 );
    or g4335 ( n7501 , n1356 , n5723 );
    or g4336 ( n1250 , n13130 , n6071 );
    or g4337 ( n13393 , n1669 , n6988 );
    and g4338 ( n1418 , n8238 , n5797 );
    and g4339 ( n12983 , n10229 , n14062 );
    and g4340 ( n13638 , n13078 , n9789 );
    not g4341 ( n7052 , n13135 );
    or g4342 ( n12233 , n14088 , n12000 );
    nor g4343 ( n9727 , n3107 , n8534 );
    not g4344 ( n12844 , n4777 );
    or g4345 ( n11271 , n6471 , n7566 );
    not g4346 ( n9950 , n13725 );
    and g4347 ( n2824 , n1254 , n12377 );
    or g4348 ( n6749 , n8828 , n2156 );
    and g4349 ( n6684 , n1071 , n10645 );
    and g4350 ( n8098 , n10408 , n13589 );
    and g4351 ( n7158 , n10506 , n2416 );
    and g4352 ( n2676 , n5048 , n4537 );
    or g4353 ( n3649 , n2686 , n1625 );
    and g4354 ( n4930 , n808 , n10488 );
    and g4355 ( n8157 , n11142 , n10777 );
    and g4356 ( n1155 , n9972 , n14453 );
    or g4357 ( n11227 , n6703 , n3893 );
    or g4358 ( n8323 , n12023 , n8531 );
    not g4359 ( n9871 , n13257 );
    and g4360 ( n1459 , n10302 , n7735 );
    or g4361 ( n12064 , n14188 , n9656 );
    and g4362 ( n12791 , n9297 , n14256 );
    not g4363 ( n7455 , n1378 );
    and g4364 ( n7686 , n10516 , n9535 );
    or g4365 ( n13633 , n787 , n462 );
    not g4366 ( n10084 , n10376 );
    and g4367 ( n14454 , n1452 , n7373 );
    not g4368 ( n4382 , n8262 );
    or g4369 ( n4968 , n8242 , n3713 );
    and g4370 ( n1879 , n14446 , n5114 );
    and g4371 ( n5031 , n3435 , n8862 );
    or g4372 ( n7051 , n10294 , n11161 );
    or g4373 ( n2730 , n9151 , n6166 );
    not g4374 ( n14370 , n2472 );
    or g4375 ( n2916 , n1582 , n5516 );
    or g4376 ( n6253 , n7229 , n3666 );
    or g4377 ( n9882 , n11379 , n14253 );
    or g4378 ( n4826 , n4807 , n2157 );
    nor g4379 ( n4283 , n5391 , n4523 );
    or g4380 ( n11661 , n7212 , n11514 );
    nor g4381 ( n2703 , n3019 , n11496 );
    nor g4382 ( n4183 , n7130 , n2075 );
    or g4383 ( n9020 , n695 , n13710 );
    or g4384 ( n10838 , n11576 , n1289 );
    and g4385 ( n1308 , n12013 , n13852 );
    not g4386 ( n14093 , n442 );
    or g4387 ( n3233 , n7590 , n7450 );
    or g4388 ( n7526 , n1362 , n12961 );
    or g4389 ( n3542 , n6600 , n14475 );
    not g4390 ( n10289 , n14154 );
    and g4391 ( n9523 , n2783 , n11366 );
    or g4392 ( n2954 , n480 , n5539 );
    not g4393 ( n3054 , n1462 );
    or g4394 ( n7735 , n8242 , n5411 );
    not g4395 ( n5738 , n12107 );
    and g4396 ( n5727 , n3932 , n9043 );
    nor g4397 ( n12740 , n2016 , n2344 );
    and g4398 ( n13527 , n1775 , n3819 );
    or g4399 ( n6230 , n10191 , n12791 );
    nor g4400 ( n1976 , n11309 , n1091 );
    or g4401 ( n13794 , n9507 , n9979 );
    not g4402 ( n13759 , n7027 );
    or g4403 ( n11323 , n2149 , n10813 );
    not g4404 ( n600 , n10046 );
    and g4405 ( n8131 , n2925 , n1946 );
    or g4406 ( n5249 , n11183 , n12151 );
    not g4407 ( n5904 , n5149 );
    nor g4408 ( n9213 , n5197 , n13893 );
    not g4409 ( n12107 , n11426 );
    or g4410 ( n1066 , n10834 , n4291 );
    or g4411 ( n11383 , n1189 , n11368 );
    or g4412 ( n4130 , n5084 , n11487 );
    nor g4413 ( n14517 , n3132 , n4287 );
    and g4414 ( n6280 , n8007 , n762 );
    not g4415 ( n11679 , n10376 );
    or g4416 ( n10875 , n1834 , n6701 );
    and g4417 ( n13122 , n11033 , n6767 );
    and g4418 ( n6417 , n3212 , n994 );
    nor g4419 ( n6195 , n13677 , n1263 );
    and g4420 ( n9155 , n2064 , n7253 );
    and g4421 ( n3377 , n6753 , n11921 );
    and g4422 ( n10766 , n11157 , n3758 );
    or g4423 ( n1651 , n6781 , n2736 );
    and g4424 ( n19 , n12858 , n8773 );
    nor g4425 ( n6374 , n13707 , n6407 );
    or g4426 ( n8941 , n6242 , n7952 );
    or g4427 ( n2003 , n11285 , n2426 );
    or g4428 ( n13256 , n14404 , n11996 );
    and g4429 ( n403 , n1431 , n12674 );
    or g4430 ( n4482 , n5710 , n1573 );
    and g4431 ( n1584 , n4261 , n1105 );
    and g4432 ( n11010 , n9898 , n3259 );
    and g4433 ( n4975 , n5414 , n7141 );
    and g4434 ( n14230 , n6192 , n8042 );
    and g4435 ( n1407 , n10015 , n6704 );
    nor g4436 ( n10029 , n7920 , n12133 );
    nor g4437 ( n2350 , n11988 , n6893 );
    or g4438 ( n3016 , n3826 , n11826 );
    not g4439 ( n10571 , n6536 );
    nor g4440 ( n949 , n183 , n9744 );
    or g4441 ( n7133 , n3076 , n8597 );
    and g4442 ( n9370 , n12741 , n804 );
    and g4443 ( n9371 , n12345 , n3946 );
    not g4444 ( n13484 , n9994 );
    and g4445 ( n6049 , n8801 , n7378 );
    and g4446 ( n7569 , n14120 , n11458 );
    or g4447 ( n8475 , n8378 , n1550 );
    nor g4448 ( n2186 , n8301 , n12780 );
    not g4449 ( n670 , n5118 );
    and g4450 ( n12071 , n14157 , n14342 );
    or g4451 ( n6740 , n2272 , n3950 );
    or g4452 ( n9730 , n12500 , n7855 );
    or g4453 ( n5841 , n1701 , n6881 );
    not g4454 ( n6088 , n9971 );
    and g4455 ( n937 , n10360 , n2080 );
    and g4456 ( n7630 , n8300 , n12306 );
    and g4457 ( n6492 , n12265 , n8781 );
    or g4458 ( n2031 , n8034 , n8028 );
    not g4459 ( n776 , n2744 );
    not g4460 ( n5454 , n8695 );
    or g4461 ( n8541 , n8476 , n9573 );
    nor g4462 ( n928 , n10136 , n6949 );
    and g4463 ( n6762 , n3401 , n8350 );
    nor g4464 ( n10030 , n234 , n14126 );
    not g4465 ( n14360 , n4895 );
    or g4466 ( n14445 , n6730 , n12152 );
    or g4467 ( n11409 , n7803 , n6306 );
    and g4468 ( n7480 , n4359 , n8505 );
    and g4469 ( n3477 , n904 , n13287 );
    nor g4470 ( n5410 , n3876 , n8895 );
    or g4471 ( n2331 , n2562 , n4734 );
    or g4472 ( n3137 , n5084 , n3412 );
    or g4473 ( n7607 , n1362 , n6385 );
    not g4474 ( n8543 , n9172 );
    and g4475 ( n3931 , n10197 , n1416 );
    nor g4476 ( n14300 , n3395 , n4792 );
    or g4477 ( n9313 , n2597 , n4094 );
    not g4478 ( n7015 , n7146 );
    and g4479 ( n4983 , n10556 , n5124 );
    nor g4480 ( n11915 , n7334 , n2434 );
    and g4481 ( n2382 , n533 , n13770 );
    and g4482 ( n8641 , n10332 , n11340 );
    nor g4483 ( n740 , n4534 , n4694 );
    and g4484 ( n2665 , n13863 , n1634 );
    and g4485 ( n9744 , n10458 , n7824 );
    and g4486 ( n6306 , n12935 , n8804 );
    not g4487 ( n5871 , n6451 );
    not g4488 ( n2246 , n2484 );
    and g4489 ( n11365 , n2367 , n8273 );
    or g4490 ( n11871 , n2750 , n7699 );
    and g4491 ( n9905 , n12990 , n947 );
    or g4492 ( n7271 , n1198 , n202 );
    and g4493 ( n7374 , n12092 , n10217 );
    and g4494 ( n1720 , n4098 , n422 );
    and g4495 ( n8868 , n11738 , n6861 );
    or g4496 ( n1114 , n5625 , n1450 );
    nor g4497 ( n2561 , n5986 , n7422 );
    not g4498 ( n2875 , n11493 );
    not g4499 ( n1481 , n11259 );
    or g4500 ( n7732 , n13080 , n4837 );
    or g4501 ( n11199 , n251 , n13891 );
    and g4502 ( n5985 , n1876 , n1066 );
    or g4503 ( n11784 , n2089 , n7712 );
    or g4504 ( n22 , n12808 , n13890 );
    or g4505 ( n4724 , n9716 , n9189 );
    and g4506 ( n6752 , n3028 , n2172 );
    or g4507 ( n4942 , n2857 , n2026 );
    and g4508 ( n10522 , n6130 , n5995 );
    and g4509 ( n11622 , n11142 , n4735 );
    not g4510 ( n7887 , n9169 );
    and g4511 ( n531 , n9650 , n2810 );
    and g4512 ( n13138 , n7957 , n9839 );
    and g4513 ( n7381 , n7810 , n3697 );
    or g4514 ( n1950 , n412 , n2797 );
    and g4515 ( n812 , n9944 , n11199 );
    or g4516 ( n8831 , n1834 , n3082 );
    and g4517 ( n13667 , n11748 , n4293 );
    or g4518 ( n4743 , n10062 , n997 );
    and g4519 ( n8660 , n904 , n4754 );
    or g4520 ( n4066 , n10626 , n10601 );
    not g4521 ( n1640 , n7972 );
    and g4522 ( n3357 , n14219 , n4765 );
    or g4523 ( n5908 , n10650 , n6074 );
    and g4524 ( n10273 , n4806 , n11829 );
    nor g4525 ( n3670 , n4913 , n9088 );
    or g4526 ( n11279 , n11621 , n4846 );
    and g4527 ( n10471 , n3332 , n2427 );
    and g4528 ( n11934 , n12425 , n6169 );
    or g4529 ( n8093 , n8638 , n3452 );
    or g4530 ( n7494 , n11231 , n13582 );
    not g4531 ( n5237 , n4146 );
    or g4532 ( n10064 , n954 , n6929 );
    or g4533 ( n3095 , n14029 , n2863 );
    and g4534 ( n6866 , n13246 , n1485 );
    or g4535 ( n5632 , n14366 , n1049 );
    or g4536 ( n1608 , n2784 , n5264 );
    not g4537 ( n4502 , n8002 );
    not g4538 ( n12852 , n6791 );
    or g4539 ( n7378 , n4045 , n13395 );
    nor g4540 ( n11587 , n12136 , n3260 );
    and g4541 ( n11225 , n6167 , n13808 );
    not g4542 ( n12872 , n3918 );
    or g4543 ( n4532 , n5647 , n2301 );
    or g4544 ( n12770 , n100 , n2987 );
    and g4545 ( n2970 , n6554 , n5595 );
    not g4546 ( n3923 , n9416 );
    or g4547 ( n14364 , n5450 , n12810 );
    and g4548 ( n13233 , n7060 , n9602 );
    or g4549 ( n8296 , n6690 , n5378 );
    not g4550 ( n7826 , n6113 );
    not g4551 ( n5062 , n2692 );
    not g4552 ( n7389 , n3263 );
    or g4553 ( n8261 , n12401 , n1043 );
    or g4554 ( n9164 , n7527 , n11631 );
    and g4555 ( n1896 , n1452 , n340 );
    not g4556 ( n13037 , n11842 );
    and g4557 ( n6979 , n8635 , n7999 );
    and g4558 ( n4768 , n4581 , n891 );
    and g4559 ( n12771 , n12935 , n139 );
    or g4560 ( n13110 , n100 , n13398 );
    not g4561 ( n13850 , n13181 );
    not g4562 ( n10046 , n5429 );
    and g4563 ( n10675 , n10457 , n9695 );
    nor g4564 ( n12936 , n512 , n14336 );
    and g4565 ( n10434 , n7673 , n14506 );
    and g4566 ( n2414 , n7957 , n2478 );
    not g4567 ( n9414 , n10341 );
    and g4568 ( n1009 , n10367 , n12676 );
    or g4569 ( n10982 , n12494 , n5421 );
    or g4570 ( n10211 , n8513 , n11414 );
    nor g4571 ( n12708 , n788 , n676 );
    and g4572 ( n6661 , n5764 , n4226 );
    and g4573 ( n11310 , n11313 , n3786 );
    and g4574 ( n12785 , n8252 , n10998 );
    and g4575 ( n14173 , n5012 , n2117 );
    or g4576 ( n9497 , n10857 , n13296 );
    and g4577 ( n10190 , n2158 , n5336 );
    and g4578 ( n3566 , n12986 , n3085 );
    not g4579 ( n1431 , n11668 );
    or g4580 ( n10369 , n7156 , n13264 );
    nor g4581 ( n2034 , n7179 , n9526 );
    nor g4582 ( n2431 , n11285 , n818 );
    nor g4583 ( n8573 , n8701 , n3991 );
    and g4584 ( n735 , n1071 , n11708 );
    nor g4585 ( n9948 , n10400 , n13238 );
    or g4586 ( n12240 , n3914 , n97 );
    or g4587 ( n5828 , n7697 , n10925 );
    and g4588 ( n3936 , n5553 , n2921 );
    or g4589 ( n2427 , n7530 , n3478 );
    and g4590 ( n11421 , n10767 , n2567 );
    and g4591 ( n8471 , n9544 , n7799 );
    and g4592 ( n468 , n13863 , n605 );
    not g4593 ( n2868 , n6053 );
    or g4594 ( n10520 , n7914 , n958 );
    nor g4595 ( n9612 , n11488 , n1910 );
    and g4596 ( n10418 , n2322 , n6651 );
    or g4597 ( n6347 , n573 , n204 );
    and g4598 ( n5448 , n9015 , n5495 );
    or g4599 ( n2793 , n13847 , n4566 );
    and g4600 ( n10060 , n8232 , n1443 );
    or g4601 ( n1479 , n930 , n11942 );
    or g4602 ( n1394 , n12764 , n1949 );
    not g4603 ( n11713 , n9721 );
    and g4604 ( n6741 , n200 , n6911 );
    or g4605 ( n9770 , n11710 , n8934 );
    or g4606 ( n814 , n523 , n6808 );
    or g4607 ( n12485 , n11551 , n2525 );
    and g4608 ( n8155 , n9275 , n6238 );
    or g4609 ( n9828 , n10019 , n10596 );
    and g4610 ( n13090 , n1729 , n10928 );
    or g4611 ( n9448 , n2412 , n7990 );
    or g4612 ( n14438 , n2531 , n8152 );
    or g4613 ( n10891 , n11183 , n9286 );
    or g4614 ( n3167 , n5641 , n9895 );
    not g4615 ( n3120 , n9354 );
    or g4616 ( n8438 , n5007 , n1287 );
    and g4617 ( n2176 , n8512 , n945 );
    or g4618 ( n7253 , n14337 , n2539 );
    or g4619 ( n5297 , n3826 , n8236 );
    and g4620 ( n3069 , n8025 , n2053 );
    or g4621 ( n11890 , n8490 , n3223 );
    or g4622 ( n11760 , n8701 , n8455 );
    and g4623 ( n3387 , n3672 , n7182 );
    nor g4624 ( n9520 , n7683 , n13648 );
    nor g4625 ( n10001 , n7588 , n12740 );
    and g4626 ( n9878 , n9350 , n9640 );
    not g4627 ( n3873 , n2409 );
    not g4628 ( n8524 , n10787 );
    not g4629 ( n6905 , n5151 );
    and g4630 ( n14344 , n3332 , n875 );
    or g4631 ( n11452 , n350 , n9977 );
    or g4632 ( n11307 , n3888 , n8756 );
    or g4633 ( n9452 , n4481 , n14061 );
    and g4634 ( n4912 , n1772 , n3393 );
    or g4635 ( n11518 , n11440 , n58 );
    or g4636 ( n5967 , n2874 , n5437 );
    nor g4637 ( n10041 , n3309 , n7013 );
    and g4638 ( n11996 , n8047 , n696 );
    and g4639 ( n951 , n4929 , n9014 );
    or g4640 ( n6860 , n8638 , n5726 );
    and g4641 ( n10734 , n9238 , n3243 );
    and g4642 ( n7012 , n7779 , n10021 );
    not g4643 ( n8096 , n1060 );
    and g4644 ( n4933 , n3986 , n5286 );
    or g4645 ( n4178 , n12351 , n8930 );
    nor g4646 ( n13585 , n7971 , n3439 );
    and g4647 ( n7791 , n3766 , n1412 );
    and g4648 ( n7937 , n14446 , n14511 );
    or g4649 ( n5336 , n11176 , n4862 );
    nor g4650 ( n9879 , n13477 , n13586 );
    and g4651 ( n9007 , n9232 , n2455 );
    nor g4652 ( n8276 , n4296 , n8231 );
    or g4653 ( n111 , n1391 , n10755 );
    or g4654 ( n6257 , n12844 , n11417 );
    and g4655 ( n8280 , n5553 , n4879 );
    and g4656 ( n3583 , n12900 , n7476 );
    not g4657 ( n3366 , n2048 );
    not g4658 ( n7696 , n4047 );
    or g4659 ( n13019 , n10234 , n1406 );
    or g4660 ( n9929 , n4923 , n8082 );
    or g4661 ( n8835 , n1741 , n5600 );
    and g4662 ( n5347 , n2758 , n5998 );
    and g4663 ( n12409 , n11837 , n7567 );
    or g4664 ( n10707 , n9780 , n6200 );
    and g4665 ( n7235 , n3710 , n11874 );
    or g4666 ( n1574 , n2562 , n12702 );
    not g4667 ( n2998 , n13383 );
    not g4668 ( n12968 , n2383 );
    and g4669 ( n7103 , n11406 , n8016 );
    and g4670 ( n826 , n2643 , n13809 );
    not g4671 ( n1929 , n6670 );
    or g4672 ( n13671 , n9429 , n12326 );
    nor g4673 ( n12664 , n14368 , n6686 );
    and g4674 ( n7002 , n6316 , n9849 );
    and g4675 ( n2193 , n3492 , n12572 );
    or g4676 ( n376 , n14472 , n10894 );
    not g4677 ( n12414 , n7441 );
    or g4678 ( n7766 , n6206 , n1154 );
    or g4679 ( n7243 , n11621 , n8563 );
    or g4680 ( n542 , n1821 , n4336 );
    nor g4681 ( n6284 , n13941 , n13353 );
    and g4682 ( n7295 , n7443 , n11611 );
    nor g4683 ( n7614 , n7334 , n613 );
    or g4684 ( n13563 , n8701 , n8482 );
    and g4685 ( n5276 , n12057 , n11860 );
    or g4686 ( n11725 , n4908 , n7603 );
    nor g4687 ( n1382 , n7940 , n12269 );
    or g4688 ( n6727 , n2897 , n12941 );
    and g4689 ( n14143 , n8025 , n5620 );
    or g4690 ( n7038 , n185 , n2425 );
    nor g4691 ( n7663 , n2790 , n5404 );
    and g4692 ( n897 , n3952 , n8383 );
    not g4693 ( n12522 , n6055 );
    or g4694 ( n10809 , n511 , n9045 );
    and g4695 ( n7087 , n10846 , n7390 );
    or g4696 ( n8820 , n9856 , n7061 );
    and g4697 ( n11254 , n446 , n3579 );
    and g4698 ( n1440 , n1071 , n8740 );
    and g4699 ( n3064 , n10516 , n5150 );
    not g4700 ( n6640 , n12270 );
    or g4701 ( n2802 , n4527 , n3652 );
    or g4702 ( n5073 , n11839 , n10214 );
    and g4703 ( n894 , n2587 , n8150 );
    or g4704 ( n929 , n7934 , n1776 );
    or g4705 ( n7568 , n9375 , n4489 );
    and g4706 ( n10002 , n11837 , n7266 );
    and g4707 ( n4751 , n14042 , n12093 );
    not g4708 ( n5279 , n9456 );
    and g4709 ( n9409 , n5823 , n12786 );
    and g4710 ( n3185 , n4655 , n1355 );
    or g4711 ( n9146 , n5815 , n7144 );
    and g4712 ( n3078 , n2064 , n12558 );
    not g4713 ( n8300 , n9416 );
    and g4714 ( n1435 , n6128 , n306 );
    and g4715 ( n2138 , n7826 , n9975 );
    not g4716 ( n12897 , n1742 );
    nor g4717 ( n1626 , n14419 , n10519 );
    not g4718 ( n14366 , n4777 );
    and g4719 ( n9434 , n783 , n1917 );
    nor g4720 ( n14186 , n12705 , n12956 );
    not g4721 ( n11488 , n8027 );
    and g4722 ( n3452 , n4163 , n13026 );
    or g4723 ( n11386 , n9780 , n9369 );
    or g4724 ( n13605 , n3768 , n8080 );
    and g4725 ( n12376 , n536 , n7568 );
    or g4726 ( n2893 , n13806 , n2635 );
    or g4727 ( n12505 , n13005 , n7388 );
    or g4728 ( n13862 , n8252 , n203 );
    and g4729 ( n8967 , n12620 , n13642 );
    or g4730 ( n8087 , n1061 , n6008 );
    and g4731 ( n4475 , n12092 , n11565 );
    or g4732 ( n1581 , n10289 , n1304 );
    or g4733 ( n3728 , n8828 , n11436 );
    nor g4734 ( n10782 , n3768 , n1050 );
    and g4735 ( n5869 , n12832 , n3136 );
    or g4736 ( n10658 , n5570 , n3315 );
    and g4737 ( n5930 , n2021 , n960 );
    and g4738 ( n12752 , n6311 , n3376 );
    and g4739 ( n9572 , n231 , n3866 );
    not g4740 ( n11316 , n7681 );
    and g4741 ( n13751 , n7627 , n60 );
    or g4742 ( n9415 , n10825 , n14255 );
    or g4743 ( n3038 , n7971 , n14122 );
    not g4744 ( n14252 , n5033 );
    or g4745 ( n3698 , n2888 , n1204 );
    or g4746 ( n13805 , n390 , n7201 );
    or g4747 ( n1281 , n12821 , n11532 );
    not g4748 ( n9069 , n3967 );
    and g4749 ( n5535 , n9952 , n5445 );
    nor g4750 ( n13340 , n6039 , n13265 );
    nor g4751 ( n3217 , n12179 , n8222 );
    and g4752 ( n14033 , n8401 , n6493 );
    and g4753 ( n4920 , n7443 , n7629 );
    or g4754 ( n13515 , n11472 , n8318 );
    or g4755 ( n10438 , n8452 , n11467 );
    nor g4756 ( n6501 , n5840 , n10733 );
    or g4757 ( n1792 , n3047 , n644 );
    and g4758 ( n7070 , n7627 , n7830 );
    and g4759 ( n8865 , n1876 , n2368 );
    or g4760 ( n2448 , n13083 , n152 );
    and g4761 ( n8674 , n5275 , n293 );
    or g4762 ( n1001 , n6471 , n5727 );
    and g4763 ( n7916 , n4525 , n5920 );
    and g4764 ( n7993 , n12531 , n7559 );
    or g4765 ( n2493 , n10936 , n6349 );
    and g4766 ( n13983 , n3736 , n609 );
    nor g4767 ( n8000 , n3400 , n4542 );
    or g4768 ( n2117 , n9140 , n12586 );
    or g4769 ( n5155 , n4498 , n11520 );
    not g4770 ( n9211 , n409 );
    or g4771 ( n2172 , n7116 , n9980 );
    and g4772 ( n1197 , n14213 , n4306 );
    not g4773 ( n428 , n11547 );
    or g4774 ( n1441 , n5715 , n10679 );
    or g4775 ( n12122 , n5800 , n9545 );
    and g4776 ( n10968 , n7267 , n2206 );
    or g4777 ( n10297 , n12169 , n7128 );
    not g4778 ( n13103 , n8524 );
    and g4779 ( n4911 , n4359 , n11956 );
    or g4780 ( n3516 , n3219 , n12812 );
    or g4781 ( n7723 , n7697 , n6974 );
    or g4782 ( n966 , n13074 , n2774 );
    or g4783 ( n11354 , n5139 , n6092 );
    or g4784 ( n12728 , n12601 , n12822 );
    not g4785 ( n393 , n7336 );
    and g4786 ( n8988 , n1354 , n7656 );
    and g4787 ( n1709 , n7043 , n691 );
    and g4788 ( n8719 , n1772 , n11669 );
    nor g4789 ( n6782 , n827 , n2235 );
    or g4790 ( n13714 , n5786 , n8552 );
    and g4791 ( n6589 , n14157 , n7571 );
    or g4792 ( n8460 , n7862 , n3369 );
    not g4793 ( n2961 , n6119 );
    and g4794 ( n13065 , n501 , n5717 );
    and g4795 ( n11736 , n11300 , n10455 );
    nor g4796 ( n5076 , n8647 , n1395 );
    and g4797 ( n9784 , n1125 , n11779 );
    and g4798 ( n11395 , n12265 , n14209 );
    and g4799 ( n11822 , n8746 , n1976 );
    or g4800 ( n8425 , n4620 , n3465 );
    not g4801 ( n14376 , n4907 );
    and g4802 ( n5356 , n11093 , n10018 );
    and g4803 ( n11367 , n8238 , n11653 );
    or g4804 ( n5706 , n782 , n12216 );
    or g4805 ( n13960 , n6090 , n2830 );
    and g4806 ( n8265 , n12611 , n4866 );
    nor g4807 ( n5255 , n3196 , n10924 );
    or g4808 ( n2110 , n8581 , n3592 );
    and g4809 ( n3718 , n8789 , n1916 );
    nor g4810 ( n3927 , n7759 , n9022 );
    not g4811 ( n13941 , n1010 );
    not g4812 ( n11748 , n5871 );
    nor g4813 ( n2757 , n12934 , n10460 );
    or g4814 ( n9454 , n10523 , n1373 );
    and g4815 ( n6273 , n1427 , n5693 );
    and g4816 ( n509 , n3766 , n13004 );
    or g4817 ( n5218 , n8528 , n2166 );
    and g4818 ( n9059 , n12998 , n10989 );
    not g4819 ( n12970 , n10423 );
    and g4820 ( n11595 , n3268 , n11087 );
    and g4821 ( n13481 , n8386 , n5867 );
    not g4822 ( n11313 , n9865 );
    and g4823 ( n8872 , n4657 , n14523 );
    or g4824 ( n14066 , n8908 , n3987 );
    and g4825 ( n8668 , n4973 , n2991 );
    or g4826 ( n5032 , n6711 , n145 );
    not g4827 ( n494 , n8997 );
    not g4828 ( n13061 , n5702 );
    or g4829 ( n109 , n6706 , n7891 );
    and g4830 ( n11461 , n11411 , n3251 );
    and g4831 ( n13169 , n5053 , n5202 );
    and g4832 ( n7199 , n9265 , n14421 );
    or g4833 ( n10964 , n5180 , n10599 );
    or g4834 ( n5223 , n4840 , n62 );
    or g4835 ( n859 , n11171 , n12565 );
    and g4836 ( n970 , n5999 , n8703 );
    nor g4837 ( n11711 , n4589 , n8257 );
    or g4838 ( n5346 , n1844 , n4137 );
    and g4839 ( n5338 , n5628 , n9962 );
    or g4840 ( n6494 , n2901 , n13880 );
    not g4841 ( n5825 , n2619 );
    not g4842 ( n5990 , n12175 );
    or g4843 ( n712 , n9856 , n10182 );
    or g4844 ( n6594 , n9984 , n9470 );
    and g4845 ( n2452 , n14327 , n6352 );
    not g4846 ( n14038 , n5665 );
    or g4847 ( n12246 , n5800 , n4661 );
    not g4848 ( n8899 , n14075 );
    or g4849 ( n5175 , n10331 , n11595 );
    or g4850 ( n10284 , n48 , n9790 );
    and g4851 ( n10042 , n14157 , n11276 );
    or g4852 ( n6481 , n1137 , n4539 );
    and g4853 ( n631 , n5348 , n4211 );
    and g4854 ( n11701 , n6822 , n1690 );
    or g4855 ( n14361 , n10300 , n14392 );
    and g4856 ( n12565 , n678 , n1507 );
    not g4857 ( n13547 , n4777 );
    or g4858 ( n3152 , n9422 , n10743 );
    nor g4859 ( n5396 , n4491 , n8861 );
    not g4860 ( n11607 , n11861 );
    and g4861 ( n13146 , n13780 , n6574 );
    and g4862 ( n759 , n12620 , n11857 );
    and g4863 ( n12457 , n6051 , n5837 );
    or g4864 ( n1286 , n14282 , n9609 );
    or g4865 ( n4423 , n2401 , n9468 );
    or g4866 ( n4640 , n2949 , n10966 );
    and g4867 ( n5515 , n9102 , n8864 );
    and g4868 ( n11741 , n10357 , n10187 );
    or g4869 ( n14077 , n1701 , n1895 );
    or g4870 ( n10414 , n8304 , n991 );
    nor g4871 ( n5521 , n7075 , n3874 );
    and g4872 ( n6216 , n8768 , n6375 );
    and g4873 ( n12725 , n103 , n8076 );
    and g4874 ( n4157 , n11484 , n3891 );
    not g4875 ( n2369 , n11771 );
    nor g4876 ( n1040 , n4544 , n6137 );
    nor g4877 ( n12780 , n12280 , n1375 );
    or g4878 ( n7595 , n2645 , n9697 );
    and g4879 ( n385 , n9885 , n11526 );
    and g4880 ( n972 , n2158 , n5572 );
    and g4881 ( n11506 , n9705 , n12463 );
    and g4882 ( n4622 , n4102 , n12553 );
    or g4883 ( n1958 , n4650 , n4615 );
    or g4884 ( n1365 , n5512 , n4131 );
    or g4885 ( n8415 , n12020 , n1151 );
    or g4886 ( n421 , n394 , n1268 );
    or g4887 ( n8971 , n13885 , n1449 );
    nor g4888 ( n8370 , n2597 , n9968 );
    and g4889 ( n9663 , n2224 , n3558 );
    not g4890 ( n1112 , n2934 );
    and g4891 ( n1201 , n6135 , n2457 );
    or g4892 ( n13410 , n5603 , n6820 );
    or g4893 ( n12415 , n251 , n13237 );
    not g4894 ( n11484 , n7802 );
    or g4895 ( n11731 , n6242 , n13624 );
    nor g4896 ( n4503 , n10186 , n1626 );
    or g4897 ( n12210 , n5139 , n732 );
    or g4898 ( n4910 , n8897 , n335 );
    nor g4899 ( n4109 , n9601 , n8467 );
    not g4900 ( n8798 , n11343 );
    not g4901 ( n10166 , n2958 );
    and g4902 ( n8854 , n2724 , n3396 );
    not g4903 ( n5952 , n4258 );
    and g4904 ( n2384 , n13236 , n1303 );
    and g4905 ( n12915 , n4627 , n12271 );
    or g4906 ( n14494 , n1840 , n4159 );
    and g4907 ( n12809 , n13745 , n1474 );
    and g4908 ( n1242 , n13489 , n10510 );
    or g4909 ( n6431 , n4468 , n9255 );
    and g4910 ( n4295 , n6311 , n12104 );
    and g4911 ( n2863 , n4657 , n13611 );
    not g4912 ( n4901 , n9967 );
    nor g4913 ( n1902 , n12569 , n10110 );
    not g4914 ( n10479 , n2791 );
    or g4915 ( n6165 , n7898 , n9646 );
    not g4916 ( n12254 , n2069 );
    and g4917 ( n7242 , n10855 , n8561 );
    or g4918 ( n11780 , n9742 , n1282 );
    or g4919 ( n640 , n12400 , n12072 );
    and g4920 ( n14276 , n4422 , n8996 );
    or g4921 ( n5477 , n7249 , n288 );
    not g4922 ( n4045 , n14354 );
    or g4923 ( n8017 , n8897 , n5311 );
    or g4924 ( n4485 , n4239 , n6491 );
    nor g4925 ( n6401 , n4091 , n5392 );
    or g4926 ( n876 , n8476 , n4303 );
    or g4927 ( n2885 , n77 , n642 );
    and g4928 ( n11872 , n13096 , n5841 );
    not g4929 ( n327 , n1458 );
    and g4930 ( n10379 , n10820 , n11497 );
    and g4931 ( n12828 , n4394 , n1264 );
    not g4932 ( n12015 , n10372 );
    and g4933 ( n2588 , n1231 , n250 );
    not g4934 ( n3037 , n11151 );
    or g4935 ( n9243 , n11980 , n3936 );
    or g4936 ( n7558 , n1051 , n245 );
    and g4937 ( n5141 , n12683 , n9249 );
    and g4938 ( n3533 , n6606 , n2872 );
    and g4939 ( n8084 , n10647 , n12753 );
    or g4940 ( n7217 , n5450 , n7592 );
    nor g4941 ( n12706 , n7052 , n9328 );
    not g4942 ( n13575 , n12765 );
    or g4943 ( n11828 , n1044 , n13311 );
    and g4944 ( n1294 , n12042 , n14097 );
    or g4945 ( n14523 , n2025 , n8728 );
    or g4946 ( n1778 , n3777 , n5616 );
    not g4947 ( n7683 , n9878 );
    and g4948 ( n10264 , n14038 , n14503 );
    not g4949 ( n8812 , n14464 );
    and g4950 ( n3315 , n6343 , n13357 );
    or g4951 ( n7650 , n11621 , n734 );
    or g4952 ( n6312 , n4199 , n9466 );
    not g4953 ( n9197 , n2778 );
    and g4954 ( n13727 , n8386 , n4926 );
    and g4955 ( n5511 , n405 , n9655 );
    and g4956 ( n10101 , n1354 , n7510 );
    and g4957 ( n5973 , n12226 , n4965 );
    or g4958 ( n3930 , n5409 , n12813 );
    and g4959 ( n1183 , n11033 , n12432 );
    and g4960 ( n10807 , n13297 , n6176 );
    or g4961 ( n2946 , n6436 , n11590 );
    or g4962 ( n1996 , n4481 , n13176 );
    or g4963 ( n13210 , n11097 , n12378 );
    not g4964 ( n1729 , n4266 );
    not g4965 ( n4156 , n13908 );
    and g4966 ( n9029 , n7852 , n11413 );
    or g4967 ( n3811 , n1006 , n11196 );
    or g4968 ( n4519 , n5861 , n3105 );
    not g4969 ( n9216 , n4716 );
    or g4970 ( n3341 , n10383 , n2626 );
    not g4971 ( n8768 , n12697 );
    and g4972 ( n5617 , n12057 , n4593 );
    not g4973 ( n553 , n4325 );
    or g4974 ( n7593 , n5253 , n952 );
    or g4975 ( n9688 , n12651 , n5794 );
    not g4976 ( n12721 , n1911 );
    and g4977 ( n165 , n10562 , n13739 );
    nor g4978 ( n14416 , n13835 , n4547 );
    and g4979 ( n6301 , n1047 , n4349 );
    nor g4980 ( n10785 , n8825 , n5784 );
    or g4981 ( n10956 , n8045 , n2978 );
    or g4982 ( n13258 , n7912 , n12446 );
    not g4983 ( n4887 , n13363 );
    or g4984 ( n7856 , n69 , n5981 );
    or g4985 ( n7639 , n1820 , n8900 );
    not g4986 ( n12846 , n3309 );
    and g4987 ( n6877 , n6822 , n3649 );
    and g4988 ( n4410 , n1339 , n4234 );
    not g4989 ( n783 , n8168 );
    nor g4990 ( n4101 , n10824 , n4385 );
    nor g4991 ( n10203 , n421 , n1062 );
    not g4992 ( n11737 , n82 );
    nor g4993 ( n10709 , n911 , n1341 );
    not g4994 ( n8629 , n521 );
    or g4995 ( n1303 , n12075 , n10734 );
    and g4996 ( n5595 , n13466 , n7484 );
    and g4997 ( n5886 , n13035 , n857 );
    not g4998 ( n1876 , n8555 );
    nor g4999 ( n7548 , n6122 , n1604 );
    or g5000 ( n6878 , n2878 , n9858 );
    or g5001 ( n5395 , n9429 , n9565 );
    not g5002 ( n1172 , n6274 );
    and g5003 ( n7168 , n13850 , n11222 );
    or g5004 ( n11604 , n11123 , n6509 );
    or g5005 ( n7290 , n10539 , n14258 );
    and g5006 ( n4353 , n5825 , n6725 );
    and g5007 ( n10096 , n10556 , n11615 );
    and g5008 ( n1823 , n627 , n5639 );
    or g5009 ( n2945 , n511 , n9817 );
    nor g5010 ( n11376 , n742 , n4278 );
    or g5011 ( n6045 , n4508 , n11978 );
    and g5012 ( n11544 , n12998 , n4702 );
    or g5013 ( n12639 , n6857 , n1935 );
    nor g5014 ( n7634 , n1462 , n9021 );
    and g5015 ( n7995 , n11495 , n38 );
    not g5016 ( n11492 , n6196 );
    and g5017 ( n14154 , n7376 , n1868 );
    and g5018 ( n16 , n3710 , n7357 );
    not g5019 ( n7081 , n6139 );
    and g5020 ( n7884 , n9113 , n13044 );
    and g5021 ( n13608 , n3277 , n10931 );
    or g5022 ( n4592 , n7912 , n11009 );
    not g5023 ( n5570 , n4891 );
    and g5024 ( n11853 , n4619 , n12190 );
    or g5025 ( n1141 , n1602 , n5187 );
    not g5026 ( n12295 , n12106 );
    or g5027 ( n733 , n4180 , n9288 );
    and g5028 ( n7202 , n10815 , n6986 );
    and g5029 ( n8259 , n10767 , n2252 );
    or g5030 ( n12395 , n11315 , n6664 );
    and g5031 ( n7516 , n9617 , n7867 );
    not g5032 ( n13698 , n12489 );
    nor g5033 ( n6584 , n6039 , n13740 );
    or g5034 ( n2593 , n4239 , n153 );
    or g5035 ( n9144 , n10731 , n8320 );
    and g5036 ( n7587 , n3942 , n12352 );
    and g5037 ( n12058 , n14093 , n7722 );
    or g5038 ( n7420 , n6109 , n314 );
    or g5039 ( n2920 , n14319 , n14002 );
    not g5040 ( n4829 , n2996 );
    and g5041 ( n201 , n5226 , n6600 );
    not g5042 ( n11047 , n6123 );
    or g5043 ( n7869 , n8983 , n12276 );
    or g5044 ( n2146 , n10083 , n6182 );
    nor g5045 ( n2133 , n329 , n11154 );
    and g5046 ( n10207 , n1428 , n13873 );
    or g5047 ( n216 , n8592 , n12172 );
    or g5048 ( n12097 , n1268 , n4895 );
    and g5049 ( n8732 , n13572 , n9486 );
    and g5050 ( n4647 , n2367 , n4054 );
    nor g5051 ( n1149 , n9291 , n7109 );
    and g5052 ( n11068 , n12357 , n3008 );
    nor g5053 ( n1851 , n13557 , n5805 );
    and g5054 ( n5563 , n4156 , n2714 );
    and g5055 ( n1455 , n11220 , n12083 );
    and g5056 ( n5796 , n4300 , n13903 );
    and g5057 ( n4545 , n10084 , n7535 );
    nor g5058 ( n2769 , n619 , n12591 );
    and g5059 ( n6050 , n3952 , n1160 );
    nor g5060 ( n12743 , n5288 , n13208 );
    and g5061 ( n10555 , n8372 , n3024 );
    and g5062 ( n8482 , n4901 , n9479 );
    not g5063 ( n12096 , n448 );
    or g5064 ( n6778 , n10624 , n12422 );
    and g5065 ( n11960 , n14093 , n4173 );
    not g5066 ( n9107 , n8682 );
    and g5067 ( n8970 , n1855 , n3531 );
    or g5068 ( n5965 , n11710 , n5030 );
    and g5069 ( n8777 , n11470 , n9398 );
    and g5070 ( n7313 , n3366 , n7682 );
    or g5071 ( n11743 , n14249 , n13636 );
    and g5072 ( n13434 , n13017 , n1003 );
    not g5073 ( n4924 , n14320 );
    or g5074 ( n51 , n11420 , n12771 );
    or g5075 ( n7949 , n4828 , n11610 );
    and g5076 ( n10865 , n6754 , n3900 );
    and g5077 ( n7715 , n10338 , n13761 );
    and g5078 ( n5803 , n10678 , n1085 );
    and g5079 ( n10753 , n12857 , n6454 );
    or g5080 ( n9477 , n4239 , n3066 );
    and g5081 ( n9101 , n8111 , n2495 );
    and g5082 ( n3500 , n7810 , n11959 );
    or g5083 ( n7840 , n7481 , n7140 );
    or g5084 ( n13792 , n4239 , n11733 );
    and g5085 ( n6198 , n3673 , n1194 );
    and g5086 ( n9816 , n80 , n9763 );
    nor g5087 ( n4430 , n8277 , n6117 );
    nor g5088 ( n6963 , n9461 , n7087 );
    and g5089 ( n5711 , n4574 , n2147 );
    and g5090 ( n3035 , n9898 , n1118 );
    or g5091 ( n9827 , n8747 , n12587 );
    not g5092 ( n706 , n7507 );
    nor g5093 ( n11154 , n5852 , n11587 );
    nor g5094 ( n11260 , n9703 , n10006 );
    and g5095 ( n2598 , n4929 , n11204 );
    and g5096 ( n3772 , n965 , n961 );
    not g5097 ( n5815 , n8695 );
    or g5098 ( n3036 , n2877 , n750 );
    or g5099 ( n10398 , n11510 , n3720 );
    and g5100 ( n10601 , n12335 , n11728 );
    not g5101 ( n7627 , n7023 );
    or g5102 ( n1973 , n13885 , n5291 );
    nor g5103 ( n7834 , n6466 , n6546 );
    and g5104 ( n12252 , n5011 , n13506 );
    or g5105 ( n11718 , n3161 , n6943 );
    and g5106 ( n4552 , n11503 , n11545 );
    or g5107 ( n4399 , n13074 , n9029 );
    and g5108 ( n5760 , n4655 , n3683 );
    or g5109 ( n1232 , n10294 , n10942 );
    or g5110 ( n5514 , n8969 , n6656 );
    nor g5111 ( n7127 , n506 , n6400 );
    and g5112 ( n13868 , n2709 , n2102 );
    or g5113 ( n7859 , n3320 , n12640 );
    and g5114 ( n6924 , n13107 , n10130 );
    and g5115 ( n5767 , n5012 , n13204 );
    or g5116 ( n912 , n14404 , n2762 );
    or g5117 ( n8325 , n7212 , n3613 );
    nor g5118 ( n7740 , n8920 , n13816 );
    or g5119 ( n1057 , n8747 , n6393 );
    and g5120 ( n4672 , n12976 , n949 );
    nor g5121 ( n6191 , n9176 , n11609 );
    or g5122 ( n8088 , n14357 , n7748 );
    and g5123 ( n4384 , n6354 , n6098 );
    or g5124 ( n5935 , n12695 , n13301 );
    not g5125 ( n77 , n4550 );
    or g5126 ( n9678 , n251 , n9248 );
    or g5127 ( n5533 , n11360 , n13402 );
    not g5128 ( n2682 , n2744 );
    or g5129 ( n9837 , n1225 , n6480 );
    or g5130 ( n11868 , n10224 , n7782 );
    or g5131 ( n7727 , n12934 , n10663 );
    or g5132 ( n2471 , n6891 , n6441 );
    and g5133 ( n3383 , n5764 , n11135 );
    or g5134 ( n4518 , n9186 , n12336 );
    and g5135 ( n3611 , n6525 , n9786 );
    or g5136 ( n12363 , n5315 , n8305 );
    nor g5137 ( n6300 , n12278 , n8365 );
    not g5138 ( n7212 , n11308 );
    or g5139 ( n13856 , n3011 , n11477 );
    or g5140 ( n4600 , n6271 , n11506 );
    and g5141 ( n1301 , n5940 , n7428 );
    not g5142 ( n13376 , n11100 );
    or g5143 ( n10077 , n11420 , n6960 );
    or g5144 ( n6506 , n8748 , n13086 );
    not g5145 ( n6209 , n13426 );
    not g5146 ( n4708 , n9305 );
    not g5147 ( n10969 , n7902 );
    not g5148 ( n7588 , n9778 );
    or g5149 ( n11948 , n11472 , n10448 );
    or g5150 ( n1856 , n5064 , n8280 );
    nor g5151 ( n2323 , n12823 , n13434 );
    and g5152 ( n7939 , n7745 , n5395 );
    nor g5153 ( n12440 , n13317 , n6521 );
    and g5154 ( n12847 , n1117 , n10496 );
    and g5155 ( n14078 , n2783 , n11468 );
    nor g5156 ( n11101 , n12292 , n7788 );
    nor g5157 ( n12116 , n4313 , n13442 );
    not g5158 ( n5071 , n13360 );
    or g5159 ( n5620 , n8490 , n5287 );
    not g5160 ( n13446 , n9846 );
    not g5161 ( n4333 , n9604 );
    nor g5162 ( n3568 , n48 , n3940 );
    and g5163 ( n11758 , n14091 , n7014 );
    and g5164 ( n3750 , n13227 , n7840 );
    not g5165 ( n3826 , n9169 );
    or g5166 ( n649 , n8490 , n10920 );
    or g5167 ( n7173 , n7249 , n14018 );
    and g5168 ( n1968 , n6854 , n6982 );
    or g5169 ( n6096 , n1210 , n9893 );
    or g5170 ( n3852 , n3667 , n11577 );
    and g5171 ( n2157 , n11816 , n7488 );
    and g5172 ( n11908 , n4856 , n189 );
    not g5173 ( n103 , n5951 );
    and g5174 ( n10440 , n11679 , n4476 );
    and g5175 ( n12939 , n5458 , n3058 );
    and g5176 ( n14214 , n5092 , n6285 );
    not g5177 ( n3222 , n5225 );
    and g5178 ( n9712 , n9323 , n2178 );
    and g5179 ( n7385 , n13755 , n3717 );
    and g5180 ( n5644 , n533 , n11162 );
    nor g5181 ( n11533 , n12046 , n5364 );
    and g5182 ( n6673 , n2474 , n14326 );
    or g5183 ( n8406 , n11176 , n923 );
    or g5184 ( n11654 , n11824 , n3775 );
    or g5185 ( n5660 , n4544 , n5142 );
    or g5186 ( n14082 , n3886 , n9103 );
    not g5187 ( n12697 , n12975 );
    not g5188 ( n4180 , n7819 );
    or g5189 ( n1572 , n3877 , n13419 );
    and g5190 ( n7986 , n225 , n233 );
    not g5191 ( n13035 , n9026 );
    or g5192 ( n8013 , n4162 , n10498 );
    or g5193 ( n4082 , n13109 , n9110 );
    not g5194 ( n9015 , n9592 );
    nor g5195 ( n12388 , n8458 , n12826 );
    or g5196 ( n14503 , n7812 , n5476 );
    and g5197 ( n7010 , n8372 , n10281 );
    and g5198 ( n14169 , n1254 , n4124 );
    and g5199 ( n1213 , n7693 , n2174 );
    or g5200 ( n5885 , n7678 , n2349 );
    or g5201 ( n8039 , n4162 , n10812 );
    or g5202 ( n9471 , n9035 , n10525 );
    or g5203 ( n9 , n9226 , n9062 );
    and g5204 ( n5476 , n9745 , n7534 );
    or g5205 ( n10989 , n2888 , n4412 );
    and g5206 ( n8556 , n12461 , n2256 );
    not g5207 ( n695 , n565 );
    not g5208 ( n10909 , n7200 );
    or g5209 ( n9374 , n7156 , n13565 );
    or g5210 ( n1667 , n13074 , n9481 );
    and g5211 ( n4587 , n3365 , n5382 );
    and g5212 ( n10918 , n11336 , n4888 );
    and g5213 ( n10654 , n6486 , n2986 );
    or g5214 ( n2602 , n5732 , n8763 );
    not g5215 ( n11803 , n10177 );
    nor g5216 ( n2380 , n2098 , n7452 );
    or g5217 ( n9005 , n2315 , n13339 );
    or g5218 ( n8549 , n3047 , n6399 );
    or g5219 ( n8637 , n12568 , n5082 );
    not g5220 ( n11668 , n3324 );
    and g5221 ( n6040 , n12802 , n6218 );
    nor g5222 ( n3089 , n3871 , n5255 );
    and g5223 ( n2979 , n7810 , n1996 );
    nor g5224 ( n12530 , n13190 , n11165 );
    not g5225 ( n6122 , n4634 );
    or g5226 ( n6459 , n1006 , n11619 );
    and g5227 ( n3369 , n9885 , n4055 );
    not g5228 ( n2497 , n739 );
    or g5229 ( n11752 , n9807 , n2700 );
    or g5230 ( n12093 , n12020 , n11423 );
    nor g5231 ( n12312 , n9924 , n2834 );
    and g5232 ( n999 , n12858 , n7998 );
    not g5233 ( n5435 , n744 );
    or g5234 ( n3900 , n9864 , n8056 );
    or g5235 ( n7571 , n2401 , n1110 );
    or g5236 ( n14304 , n9285 , n7262 );
    or g5237 ( n7405 , n7122 , n5283 );
    nor g5238 ( n12677 , n228 , n9922 );
    not g5239 ( n573 , n4847 );
    or g5240 ( n9441 , n5236 , n12855 );
    not g5241 ( n12353 , n6123 );
    and g5242 ( n7021 , n1924 , n3653 );
    and g5243 ( n14020 , n2180 , n11108 );
    nor g5244 ( n9615 , n9078 , n11147 );
    or g5245 ( n6188 , n12149 , n12160 );
    not g5246 ( n11710 , n3021 );
    not g5247 ( n12303 , n11875 );
    or g5248 ( n14348 , n10089 , n8888 );
    or g5249 ( n10295 , n12428 , n12208 );
    and g5250 ( n4215 , n7909 , n4352 );
    nor g5251 ( n8388 , n329 , n3325 );
    nor g5252 ( n6407 , n14377 , n14208 );
    not g5253 ( n8027 , n2919 );
    and g5254 ( n14460 , n13342 , n2146 );
    not g5255 ( n10713 , n12106 );
    and g5256 ( n6166 , n6135 , n8261 );
    and g5257 ( n202 , n7043 , n12613 );
    and g5258 ( n6171 , n11406 , n12158 );
    not g5259 ( n7798 , n10051 );
    or g5260 ( n2829 , n5454 , n3245 );
    and g5261 ( n2741 , n7745 , n6376 );
    and g5262 ( n4804 , n1708 , n6862 );
    or g5263 ( n3275 , n3777 , n5614 );
    not g5264 ( n11882 , n1348 );
    nor g5265 ( n7035 , n1685 , n4889 );
    or g5266 ( n13263 , n9226 , n11025 );
    and g5267 ( n3021 , n5029 , n7050 );
    or g5268 ( n12671 , n9174 , n9484 );
    or g5269 ( n11341 , n10294 , n567 );
    and g5270 ( n4316 , n4486 , n8191 );
    and g5271 ( n12358 , n12132 , n12933 );
    not g5272 ( n2510 , n630 );
    and g5273 ( n12153 , n11406 , n6773 );
    not g5274 ( n13520 , n10828 );
    or g5275 ( n465 , n13854 , n4517 );
    or g5276 ( n10886 , n5641 , n11856 );
    not g5277 ( n7852 , n5460 );
    or g5278 ( n13058 , n13941 , n4 );
    or g5279 ( n2537 , n4573 , n13511 );
    not g5280 ( n865 , n12483 );
    or g5281 ( n3176 , n3219 , n8454 );
    and g5282 ( n4784 , n13379 , n9628 );
    not g5283 ( n3905 , n10099 );
    or g5284 ( n7950 , n227 , n10972 );
    or g5285 ( n12148 , n1685 , n3456 );
    and g5286 ( n466 , n12918 , n830 );
    or g5287 ( n10499 , n12324 , n7573 );
    or g5288 ( n3183 , n6654 , n13988 );
    or g5289 ( n1787 , n7076 , n7006 );
    not g5290 ( n5618 , n8809 );
    and g5291 ( n9514 , n8401 , n5297 );
    not g5292 ( n13074 , n4465 );
    or g5293 ( n13578 , n12625 , n1718 );
    and g5294 ( n14301 , n222 , n1965 );
    and g5295 ( n9081 , n627 , n11827 );
    and g5296 ( n9762 , n4973 , n5220 );
    or g5297 ( n3178 , n10560 , n10806 );
    and g5298 ( n3075 , n2310 , n8207 );
    nor g5299 ( n10128 , n458 , n3633 );
    nor g5300 ( n5247 , n4213 , n4430 );
    nor g5301 ( n12853 , n7588 , n2948 );
    and g5302 ( n6653 , n4657 , n342 );
    or g5303 ( n4019 , n13226 , n5818 );
    and g5304 ( n447 , n11679 , n14156 );
    or g5305 ( n41 , n2246 , n1567 );
    not g5306 ( n2236 , n1214 );
    nor g5307 ( n6430 , n3497 , n7850 );
    and g5308 ( n10935 , n3986 , n12774 );
    or g5309 ( n2402 , n4128 , n13719 );
    nor g5310 ( n11206 , n7188 , n1007 );
    or g5311 ( n12553 , n13220 , n8977 );
    or g5312 ( n6331 , n3559 , n1584 );
    and g5313 ( n10337 , n55 , n11337 );
    or g5314 ( n10253 , n7122 , n1709 );
    and g5315 ( n14378 , n2820 , n11248 );
    and g5316 ( n939 , n638 , n7703 );
    and g5317 ( n11682 , n10855 , n2955 );
    and g5318 ( n6745 , n10457 , n5768 );
    or g5319 ( n9413 , n185 , n8474 );
    or g5320 ( n3968 , n8045 , n13775 );
    and g5321 ( n7018 , n5779 , n2549 );
    not g5322 ( n10019 , n12776 );
    and g5323 ( n5608 , n4525 , n2307 );
    not g5324 ( n10922 , n4824 );
    not g5325 ( n5919 , n8925 );
    or g5326 ( n10454 , n11379 , n3648 );
    or g5327 ( n7974 , n1362 , n2914 );
    or g5328 ( n1491 , n11909 , n7506 );
    or g5329 ( n4411 , n5132 , n2467 );
    or g5330 ( n9057 , n647 , n7657 );
    or g5331 ( n2495 , n5507 , n12963 );
    nor g5332 ( n57 , n12630 , n9995 );
    and g5333 ( n9501 , n9705 , n2506 );
    not g5334 ( n8291 , n5197 );
    or g5335 ( n5972 , n10154 , n9805 );
    nor g5336 ( n9303 , n163 , n5521 );
    or g5337 ( n6876 , n6428 , n9687 );
    or g5338 ( n1236 , n1028 , n8850 );
    and g5339 ( n6521 , n706 , n4743 );
    or g5340 ( n12016 , n5483 , n5602 );
    and g5341 ( n10996 , n13535 , n5212 );
    and g5342 ( n10769 , n10969 , n8994 );
    and g5343 ( n5739 , n10705 , n7930 );
    or g5344 ( n9492 , n8172 , n11677 );
    or g5345 ( n7228 , n7003 , n5167 );
    or g5346 ( n7901 , n4407 , n6969 );
    and g5347 ( n14255 , n12460 , n4799 );
    and g5348 ( n5 , n12611 , n10335 );
    and g5349 ( n9710 , n10209 , n12016 );
    or g5350 ( n11588 , n4407 , n13822 );
    and g5351 ( n9446 , n9726 , n1490 );
    or g5352 ( n2139 , n11438 , n5408 );
    or g5353 ( n14511 , n4498 , n12943 );
    or g5354 ( n4318 , n7684 , n4088 );
    and g5355 ( n6913 , n12226 , n525 );
    or g5356 ( n7019 , n6711 , n11226 );
    and g5357 ( n13455 , n11163 , n3881 );
    and g5358 ( n12903 , n13338 , n2661 );
    not g5359 ( n2171 , n3345 );
    or g5360 ( n7149 , n251 , n10817 );
    nor g5361 ( n7124 , n5952 , n1084 );
    and g5362 ( n3746 , n80 , n12599 );
    or g5363 ( n6363 , n6519 , n4933 );
    and g5364 ( n1072 , n14227 , n5120 );
    or g5365 ( n7408 , n2236 , n5125 );
    and g5366 ( n3647 , n4806 , n12799 );
    and g5367 ( n3237 , n5918 , n10722 );
    or g5368 ( n6353 , n8821 , n11457 );
    not g5369 ( n13811 , n11435 );
    and g5370 ( n6322 , n9323 , n10120 );
    not g5371 ( n1125 , n168 );
    and g5372 ( n11992 , n8432 , n4915 );
    not g5373 ( n7697 , n4847 );
    not g5374 ( n954 , n11152 );
    or g5375 ( n13843 , n10731 , n12704 );
    not g5376 ( n11036 , n918 );
    or g5377 ( n4119 , n1914 , n7363 );
    or g5378 ( n9535 , n11722 , n759 );
    and g5379 ( n12685 , n4244 , n9234 );
    not g5380 ( n10506 , n10973 );
    and g5381 ( n3980 , n7909 , n5492 );
    not g5382 ( n4877 , n10889 );
    and g5383 ( n7312 , n8768 , n1947 );
    and g5384 ( n13114 , n10470 , n8269 );
    or g5385 ( n14496 , n12295 , n9004 );
    not g5386 ( n2874 , n10629 );
    not g5387 ( n718 , n5525 );
    and g5388 ( n9071 , n8692 , n9880 );
    nor g5389 ( n7143 , n5665 , n1019 );
    or g5390 ( n6637 , n7227 , n14301 );
    or g5391 ( n11866 , n695 , n3534 );
    nor g5392 ( n10921 , n2953 , n7202 );
    not g5393 ( n5575 , n11308 );
    and g5394 ( n8018 , n12265 , n443 );
    not g5395 ( n8511 , n3946 );
    and g5396 ( n9042 , n4394 , n7058 );
    nor g5397 ( n3769 , n4913 , n7740 );
    and g5398 ( n4566 , n9069 , n1001 );
    and g5399 ( n9537 , n4267 , n6673 );
    not g5400 ( n906 , n6053 );
    and g5401 ( n4952 , n13525 , n7294 );
    and g5402 ( n9739 , n3715 , n10208 );
    and g5403 ( n1465 , n4657 , n2042 );
    and g5404 ( n785 , n8786 , n11593 );
    and g5405 ( n6138 , n12425 , n8694 );
    and g5406 ( n13763 , n13484 , n11752 );
    and g5407 ( n6532 , n4509 , n2271 );
    not g5408 ( n6638 , n1548 );
    and g5409 ( n2600 , n6316 , n13757 );
    nor g5410 ( n9595 , n9266 , n3477 );
    or g5411 ( n293 , n11572 , n4703 );
    not g5412 ( n151 , n2354 );
    not g5413 ( n3777 , n238 );
    nor g5414 ( n11198 , n4741 , n8617 );
    and g5415 ( n1848 , n7677 , n2329 );
    and g5416 ( n4238 , n10332 , n2068 );
    and g5417 ( n8867 , n9853 , n1498 );
    and g5418 ( n11848 , n4445 , n14155 );
    or g5419 ( n14115 , n12131 , n3941 );
    nor g5420 ( n4212 , n14133 , n12380 );
    or g5421 ( n13724 , n11510 , n784 );
    or g5422 ( n11070 , n5266 , n5303 );
    or g5423 ( n7817 , n4233 , n13445 );
    and g5424 ( n13373 , n13484 , n11261 );
    or g5425 ( n7619 , n3888 , n4265 );
    or g5426 ( n5099 , n13220 , n8241 );
    and g5427 ( n6226 , n14358 , n634 );
    and g5428 ( n3534 , n9345 , n2402 );
    nor g5429 ( n6290 , n6085 , n68 );
    and g5430 ( n3105 , n8372 , n10068 );
    or g5431 ( n9061 , n8825 , n2313 );
    nor g5432 ( n14336 , n12934 , n13235 );
    not g5433 ( n1802 , n4282 );
    or g5434 ( n9329 , n263 , n4000 );
    or g5435 ( n2263 , n11105 , n14339 );
    or g5436 ( n7360 , n10626 , n1272 );
    and g5437 ( n10262 , n9571 , n8826 );
    nor g5438 ( n10460 , n7238 , n9177 );
    nor g5439 ( n12911 , n4913 , n14170 );
    or g5440 ( n2974 , n12149 , n6831 );
    and g5441 ( n10893 , n5317 , n9296 );
    nor g5442 ( n2660 , n6428 , n5527 );
    and g5443 ( n8696 , n2465 , n9225 );
    or g5444 ( n3304 , n12324 , n1142 );
    not g5445 ( n11724 , n3357 );
    and g5446 ( n1095 , n11484 , n6321 );
    or g5447 ( n7033 , n3099 , n9591 );
    and g5448 ( n13995 , n1854 , n14295 );
    and g5449 ( n6056 , n13656 , n13068 );
    and g5450 ( n12762 , n13656 , n11236 );
    nor g5451 ( n4090 , n7245 , n2044 );
    nor g5452 ( n14208 , n2218 , n11711 );
    or g5453 ( n7356 , n13016 , n102 );
    not g5454 ( n8452 , n2545 );
    nor g5455 ( n2666 , n1383 , n9482 );
    or g5456 ( n13418 , n7426 , n8933 );
    or g5457 ( n11134 , n13707 , n3703 );
    or g5458 ( n2628 , n7438 , n2242 );
    nor g5459 ( n13584 , n2428 , n13999 );
    or g5460 ( n1888 , n8517 , n2600 );
    and g5461 ( n11664 , n13814 , n11332 );
    and g5462 ( n7719 , n1047 , n1862 );
    and g5463 ( n8802 , n13227 , n14197 );
    and g5464 ( n6355 , n3715 , n5040 );
    or g5465 ( n6593 , n11722 , n11499 );
    and g5466 ( n10696 , n8250 , n4512 );
    not g5467 ( n13466 , n9544 );
    and g5468 ( n13259 , n12209 , n8233 );
    nor g5469 ( n10244 , n12651 , n13596 );
    or g5470 ( n6994 , n4255 , n962 );
    and g5471 ( n6785 , n2461 , n6528 );
    and g5472 ( n6832 , n2904 , n3824 );
    not g5473 ( n6670 , n7662 );
    not g5474 ( n12620 , n5268 );
    or g5475 ( n5680 , n9218 , n2763 );
    not g5476 ( n13255 , n8106 );
    and g5477 ( n8499 , n5088 , n3660 );
    and g5478 ( n6237 , n12772 , n7594 );
    nor g5479 ( n4570 , n8023 , n4960 );
    and g5480 ( n7642 , n5071 , n5972 );
    or g5481 ( n12129 , n5695 , n7794 );
    or g5482 ( n6297 , n1660 , n9644 );
    and g5483 ( n8264 , n7673 , n2894 );
    and g5484 ( n2884 , n11814 , n221 );
    or g5485 ( n9293 , n2518 , n14490 );
    or g5486 ( n4728 , n10331 , n4752 );
    not g5487 ( n511 , n11331 );
    and g5488 ( n7338 , n7208 , n12062 );
    or g5489 ( n8428 , n8301 , n4582 );
    and g5490 ( n7090 , n10820 , n6446 );
    and g5491 ( n6847 , n11636 , n11625 );
    and g5492 ( n8306 , n1093 , n3638 );
    and g5493 ( n6856 , n4445 , n8624 );
    and g5494 ( n849 , n865 , n3129 );
    and g5495 ( n3851 , n14388 , n6292 );
    or g5496 ( n12898 , n9230 , n1245 );
    and g5497 ( n14513 , n9238 , n10580 );
    or g5498 ( n9025 , n1172 , n680 );
    or g5499 ( n9301 , n3120 , n1989 );
    and g5500 ( n2219 , n14327 , n13486 );
    and g5501 ( n4297 , n9188 , n8492 );
    and g5502 ( n7280 , n9944 , n862 );
    or g5503 ( n11806 , n12500 , n5922 );
    or g5504 ( n10143 , n4199 , n10354 );
    not g5505 ( n5038 , n9305 );
    and g5506 ( n11361 , n1876 , n14167 );
    nor g5507 ( n11762 , n5480 , n8000 );
    and g5508 ( n6868 , n718 , n4695 );
    and g5509 ( n9201 , n10822 , n8971 );
    and g5510 ( n7952 , n10710 , n9770 );
    and g5511 ( n6808 , n12620 , n6379 );
    and g5512 ( n9004 , n12389 , n9808 );
    or g5513 ( n4819 , n14088 , n2853 );
    nor g5514 ( n9848 , n234 , n6325 );
    nor g5515 ( n4766 , n11047 , n10723 );
    nor g5516 ( n13140 , n4534 , n13168 );
    or g5517 ( n8129 , n12324 , n5906 );
    or g5518 ( n11729 , n10560 , n7031 );
    or g5519 ( n5770 , n6596 , n4493 );
    nor g5520 ( n7069 , n6085 , n14248 );
    and g5521 ( n1288 , n11142 , n26 );
    and g5522 ( n14469 , n14373 , n11007 );
    and g5523 ( n4764 , n7852 , n6485 );
    and g5524 ( n9646 , n55 , n1988 );
    and g5525 ( n967 , n12455 , n364 );
    or g5526 ( n6566 , n5406 , n902 );
    or g5527 ( n13524 , n6109 , n9299 );
    and g5528 ( n7797 , n7852 , n5924 );
    nor g5529 ( n12982 , n13675 , n3560 );
    and g5530 ( n11768 , n12460 , n3322 );
    not g5531 ( n3134 , n1214 );
    and g5532 ( n10546 , n2547 , n8107 );
    or g5533 ( n12420 , n14449 , n8423 );
    and g5534 ( n13045 , n12321 , n3410 );
    or g5535 ( n13384 , n1362 , n8717 );
    nor g5536 ( n5199 , n11558 , n8929 );
    nor g5537 ( n12467 , n7889 , n6185 );
    or g5538 ( n1336 , n4207 , n2045 );
    or g5539 ( n1008 , n14110 , n5759 );
    and g5540 ( n10311 , n3286 , n14059 );
    or g5541 ( n13933 , n2843 , n5638 );
    or g5542 ( n14118 , n2529 , n7988 );
    nor g5543 ( n8417 , n12254 , n9879 );
    and g5544 ( n7344 , n965 , n14144 );
    and g5545 ( n12417 , n646 , n13117 );
    and g5546 ( n12459 , n10015 , n7743 );
    or g5547 ( n3079 , n7076 , n2580 );
    not g5548 ( n14198 , n7322 );
    or g5549 ( n9127 , n1614 , n3068 );
    not g5550 ( n9571 , n11369 );
    nor g5551 ( n7164 , n1713 , n9019 );
    not g5552 ( n3932 , n7278 );
    or g5553 ( n3747 , n619 , n6040 );
    and g5554 ( n3853 , n4722 , n11014 );
    or g5555 ( n11135 , n13477 , n877 );
    nor g5556 ( n10885 , n8424 , n4575 );
    nor g5557 ( n9552 , n7971 , n2584 );
    or g5558 ( n10984 , n4407 , n897 );
    and g5559 ( n8565 , n11738 , n9373 );
    nor g5560 ( n9126 , n3309 , n809 );
    not g5561 ( n10285 , n3191 );
    not g5562 ( n2503 , n12904 );
    nor g5563 ( n886 , n7192 , n3479 );
    or g5564 ( n14027 , n5575 , n1095 );
    or g5565 ( n3609 , n9127 , n9698 );
    and g5566 ( n5428 , n12159 , n12713 );
    or g5567 ( n605 , n3076 , n1518 );
    nor g5568 ( n9458 , n2868 , n12677 );
    and g5569 ( n12974 , n4394 , n11683 );
    and g5570 ( n14473 , n6051 , n9887 );
    or g5571 ( n12328 , n12576 , n8662 );
    or g5572 ( n11217 , n116 , n13704 );
    and g5573 ( n2659 , n8431 , n11849 );
    and g5574 ( n8289 , n4486 , n4968 );
    not g5575 ( n7079 , n871 );
    nor g5576 ( n7643 , n3602 , n9704 );
    or g5577 ( n6518 , n12112 , n6342 );
    or g5578 ( n10327 , n8151 , n11255 );
    not g5579 ( n14042 , n12450 );
    or g5580 ( n8811 , n4840 , n4298 );
    and g5581 ( n7400 , n7909 , n14516 );
    or g5582 ( n5583 , n5359 , n2187 );
    or g5583 ( n8075 , n4822 , n9923 );
    and g5584 ( n8944 , n12802 , n5543 );
    not g5585 ( n14337 , n12874 );
    not g5586 ( n1028 , n630 );
    and g5587 ( n1289 , n2682 , n11937 );
    not g5588 ( n228 , n5901 );
    and g5589 ( n3752 , n6854 , n5089 );
    not g5590 ( n9604 , n12888 );
    or g5591 ( n13542 , n9136 , n6422 );
    and g5592 ( n9996 , n6625 , n9874 );
    nor g5593 ( n9785 , n11180 , n7783 );
    not g5594 ( n300 , n10787 );
    not g5595 ( n7980 , n1377 );
    or g5596 ( n12688 , n4407 , n13855 );
    and g5597 ( n7620 , n12389 , n9991 );
    nor g5598 ( n5938 , n3640 , n5966 );
    not g5599 ( n6797 , n9740 );
    not g5600 ( n11232 , n2257 );
    or g5601 ( n10049 , n11121 , n3853 );
    or g5602 ( n7014 , n13698 , n7106 );
    not g5603 ( n2799 , n10046 );
    nor g5604 ( n13670 , n5840 , n618 );
    not g5605 ( n5926 , n11369 );
    and g5606 ( n10899 , n1962 , n8211 );
    and g5607 ( n5555 , n4359 , n5830 );
    and g5608 ( n14365 , n8817 , n12785 );
    or g5609 ( n7118 , n766 , n892 );
    or g5610 ( n12424 , n2229 , n6031 );
    or g5611 ( n2326 , n1044 , n7835 );
    and g5612 ( n7185 , n776 , n11110 );
    or g5613 ( n5920 , n9856 , n3780 );
    and g5614 ( n3103 , n2461 , n7922 );
    and g5615 ( n3041 , n10374 , n7483 );
    not g5616 ( n3 , n14216 );
    and g5617 ( n10892 , n8849 , n10184 );
    or g5618 ( n5642 , n4468 , n4034 );
    and g5619 ( n2145 , n13407 , n5302 );
    or g5620 ( n9433 , n11620 , n10507 );
    and g5621 ( n13905 , n9898 , n1957 );
    or g5622 ( n10073 , n5234 , n7978 );
    not g5623 ( n4358 , n1955 );
    or g5624 ( n4915 , n11551 , n13607 );
    and g5625 ( n3033 , n7391 , n1 );
    and g5626 ( n3999 , n5088 , n13119 );
    not g5627 ( n10032 , n12970 );
    not g5628 ( n10714 , n6905 );
    or g5629 ( n3009 , n11749 , n2073 );
    or g5630 ( n13711 , n9529 , n2971 );
    not g5631 ( n6039 , n12394 );
    and g5632 ( n7206 , n4554 , n12840 );
    not g5633 ( n9898 , n871 );
    not g5634 ( n11113 , n8887 );
    or g5635 ( n12375 , n5695 , n9357 );
    or g5636 ( n6304 , n11621 , n12747 );
    and g5637 ( n12801 , n6157 , n11168 );
    and g5638 ( n9495 , n8768 , n6409 );
    or g5639 ( n10178 , n9620 , n773 );
    and g5640 ( n2498 , n9321 , n13960 );
    not g5641 ( n10233 , n7704 );
    and g5642 ( n5405 , n776 , n5865 );
    nor g5643 ( n7536 , n5558 , n1959 );
    and g5644 ( n5895 , n2846 , n419 );
    or g5645 ( n13536 , n9375 , n1036 );
    not g5646 ( n3164 , n2472 );
    and g5647 ( n1687 , n4627 , n6620 );
    or g5648 ( n9695 , n9804 , n4962 );
    or g5649 ( n11288 , n48 , n7127 );
    and g5650 ( n4813 , n9198 , n12242 );
    or g5651 ( n1537 , n5253 , n4114 );
    or g5652 ( n3552 , n8151 , n8433 );
    nor g5653 ( n9276 , n703 , n9647 );
    or g5654 ( n1264 , n11405 , n6432 );
    nor g5655 ( n13810 , n4544 , n3351 );
    not g5656 ( n12693 , n8500 );
    and g5657 ( n10070 , n646 , n2493 );
    and g5658 ( n10313 , n11153 , n11253 );
    or g5659 ( n11979 , n5548 , n5541 );
    and g5660 ( n2458 , n8605 , n10111 );
    or g5661 ( n13287 , n11710 , n3279 );
    and g5662 ( n3227 , n3204 , n5881 );
    not g5663 ( n12127 , n10236 );
    not g5664 ( n55 , n6787 );
    or g5665 ( n10572 , n6271 , n8734 );
    or g5666 ( n12371 , n283 , n3423 );
    and g5667 ( n5792 , n10763 , n8911 );
    and g5668 ( n2337 , n6957 , n10520 );
    and g5669 ( n14086 , n3607 , n10104 );
    and g5670 ( n12993 , n11702 , n12842 );
    nor g5671 ( n14324 , n4207 , n14318 );
    and g5672 ( n13152 , n8020 , n4075 );
    and g5673 ( n10896 , n12018 , n10845 );
    or g5674 ( n2162 , n553 , n4983 );
    and g5675 ( n9299 , n8232 , n2400 );
    or g5676 ( n4480 , n1613 , n8538 );
    or g5677 ( n1102 , n11724 , n2333 );
    nor g5678 ( n14520 , n584 , n13030 );
    or g5679 ( n11749 , n12581 , n1022 );
    and g5680 ( n12745 , n3672 , n6707 );
    and g5681 ( n153 , n5062 , n6500 );
    not g5682 ( n2619 , n3812 );
    and g5683 ( n2832 , n12389 , n10997 );
    or g5684 ( n13940 , n8986 , n1273 );
    and g5685 ( n743 , n12013 , n4827 );
    or g5686 ( n993 , n10234 , n7553 );
    not g5687 ( n7803 , n10629 );
    and g5688 ( n7382 , n844 , n2892 );
    or g5689 ( n7177 , n12480 , n3655 );
    and g5690 ( n363 , n9944 , n76 );
    not g5691 ( n4562 , n7064 );
    not g5692 ( n14060 , n12278 );
    and g5693 ( n6478 , n4655 , n14108 );
    and g5694 ( n5791 , n1775 , n13789 );
    and g5695 ( n7224 , n5229 , n10414 );
    nor g5696 ( n11747 , n2468 , n14112 );
    and g5697 ( n8365 , n10059 , n7395 );
    or g5698 ( n1922 , n11804 , n8906 );
    not g5699 ( n13677 , n5294 );
    or g5700 ( n9582 , n10154 , n3215 );
    or g5701 ( n4931 , n8964 , n14020 );
    or g5702 ( n9077 , n568 , n2192 );
    or g5703 ( n8327 , n3800 , n279 );
    or g5704 ( n960 , n13080 , n11021 );
    and g5705 ( n9918 , n12620 , n9264 );
    or g5706 ( n10789 , n13718 , n14160 );
    not g5707 ( n10649 , n4708 );
    nor g5708 ( n5978 , n4207 , n7496 );
    or g5709 ( n10328 , n4807 , n3994 );
    and g5710 ( n4703 , n8789 , n8160 );
    not g5711 ( n13108 , n6264 );
    or g5712 ( n13430 , n3025 , n7205 );
    or g5713 ( n7653 , n10560 , n12754 );
    not g5714 ( n12503 , n9193 );
    or g5715 ( n12317 , n13698 , n7239 );
    and g5716 ( n220 , n13035 , n6022 );
    and g5717 ( n7319 , n10562 , n10398 );
    or g5718 ( n1836 , n9174 , n8244 );
    and g5719 ( n3004 , n706 , n12443 );
    and g5720 ( n373 , n9890 , n10558 );
    not g5721 ( n11998 , n11071 );
    or g5722 ( n1853 , n11285 , n3631 );
    nor g5723 ( n4164 , n9913 , n12848 );
    or g5724 ( n757 , n1137 , n9129 );
    or g5725 ( n1961 , n1391 , n10434 );
    and g5726 ( n2642 , n1117 , n410 );
    and g5727 ( n3898 , n5275 , n12285 );
    and g5728 ( n102 , n6135 , n6420 );
    not g5729 ( n7122 , n9686 );
    and g5730 ( n6091 , n7421 , n2213 );
    or g5731 ( n5357 , n6242 , n4236 );
    and g5732 ( n13170 , n11950 , n9729 );
    or g5733 ( n4194 , n5762 , n1666 );
    not g5734 ( n3345 , n4589 );
    or g5735 ( n10611 , n7530 , n8221 );
    or g5736 ( n7449 , n5493 , n6240 );
    and g5737 ( n4209 , n4806 , n9771 );
    or g5738 ( n9839 , n13142 , n6856 );
    not g5739 ( n12727 , n14016 );
    or g5740 ( n11241 , n12169 , n9402 );
    or g5741 ( n14458 , n85 , n5773 );
    nor g5742 ( n11449 , n7229 , n4738 );
    and g5743 ( n46 , n10080 , n7474 );
    or g5744 ( n9220 , n3062 , n1502 );
    nor g5745 ( n12347 , n8458 , n3651 );
    or g5746 ( n3202 , n12351 , n7987 );
    and g5747 ( n7982 , n2322 , n12363 );
    and g5748 ( n1549 , n3276 , n4514 );
    or g5749 ( n3630 , n11459 , n14 );
    and g5750 ( n10804 , n14388 , n2207 );
    and g5751 ( n8134 , n9245 , n416 );
    or g5752 ( n8846 , n3062 , n10564 );
    not g5753 ( n2866 , n6965 );
    not g5754 ( n889 , n168 );
    nor g5755 ( n3582 , n1243 , n14229 );
    and g5756 ( n9086 , n9726 , n2139 );
    not g5757 ( n14455 , n9172 );
    and g5758 ( n9917 , n9015 , n11286 );
    and g5759 ( n12407 , n5011 , n13949 );
    nor g5760 ( n8127 , n13477 , n9521 );
    and g5761 ( n13251 , n11157 , n14102 );
    and g5762 ( n9569 , n13745 , n5552 );
    or g5763 ( n593 , n850 , n6091 );
    not g5764 ( n7023 , n8357 );
    and g5765 ( n6186 , n536 , n13180 );
    or g5766 ( n9550 , n3263 , n11345 );
    and g5767 ( n5826 , n1481 , n10821 );
    and g5768 ( n11694 , n6311 , n13092 );
    or g5769 ( n10420 , n1711 , n11675 );
    or g5770 ( n12237 , n1602 , n4873 );
    nor g5771 ( n11926 , n151 , n10030 );
    and g5772 ( n9664 , n14313 , n7194 );
    and g5773 ( n11278 , n4627 , n10788 );
    and g5774 ( n5421 , n5312 , n971 );
    or g5775 ( n8422 , n2089 , n10171 );
    and g5776 ( n12702 , n11406 , n9044 );
    or g5777 ( n7466 , n74 , n13109 );
    or g5778 ( n6223 , n5362 , n10039 );
    or g5779 ( n10549 , n4045 , n2509 );
    or g5780 ( n3335 , n5007 , n3913 );
    not g5781 ( n12357 , n6810 );
    and g5782 ( n58 , n13572 , n12395 );
    or g5783 ( n8771 , n13531 , n8642 );
    or g5784 ( n4955 , n4065 , n8503 );
    or g5785 ( n3403 , n3777 , n7752 );
    and g5786 ( n9473 , n9238 , n7022 );
    or g5787 ( n2625 , n6263 , n12043 );
    and g5788 ( n2196 , n11816 , n11540 );
    or g5789 ( n12022 , n2181 , n9058 );
    not g5790 ( n2878 , n622 );
    or g5791 ( n4961 , n5266 , n4308 );
    or g5792 ( n323 , n3512 , n14479 );
    or g5793 ( n9761 , n12994 , n5439 );
    and g5794 ( n7958 , n2082 , n6160 );
    and g5795 ( n6713 , n13676 , n12399 );
    and g5796 ( n2198 , n333 , n12240 );
    or g5797 ( n13930 , n3914 , n8114 );
    and g5798 ( n4687 , n7041 , n5856 );
    and g5799 ( n13674 , n2445 , n9711 );
    not g5800 ( n5472 , n12394 );
    nor g5801 ( n10456 , n11580 , n9700 );
    and g5802 ( n6068 , n4722 , n4026 );
    not g5803 ( n1189 , n9580 );
    or g5804 ( n12597 , n9804 , n8875 );
    or g5805 ( n724 , n6085 , n12758 );
    not g5806 ( n8496 , n4105 );
    or g5807 ( n4431 , n12034 , n2941 );
    or g5808 ( n7731 , n11839 , n3864 );
    and g5809 ( n8097 , n9898 , n1536 );
    and g5810 ( n2351 , n14042 , n13058 );
    and g5811 ( n6591 , n6744 , n3115 );
    or g5812 ( n11526 , n5861 , n6082 );
    and g5813 ( n2941 , n3743 , n14355 );
    or g5814 ( n14220 , n4908 , n10792 );
    and g5815 ( n2524 , n4871 , n9587 );
    and g5816 ( n8520 , n646 , n9832 );
    and g5817 ( n880 , n7053 , n1475 );
    or g5818 ( n4036 , n4443 , n1347 );
    or g5819 ( n3363 , n10808 , n2270 );
    or g5820 ( n5372 , n2843 , n13303 );
    not g5821 ( n14320 , n7052 );
    nor g5822 ( n2030 , n10929 , n12964 );
    or g5823 ( n9428 , n9490 , n13514 );
    or g5824 ( n10076 , n5807 , n14078 );
    nor g5825 ( n5325 , n5897 , n4337 );
    not g5826 ( n501 , n5108 );
    or g5827 ( n11705 , n5861 , n10555 );
    and g5828 ( n12584 , n13147 , n9235 );
    or g5829 ( n4461 , n3815 , n13146 );
    and g5830 ( n13160 , n1266 , n13178 );
    or g5831 ( n12056 , n8980 , n1476 );
    and g5832 ( n1157 , n5092 , n1621 );
    not g5833 ( n9321 , n8798 );
    and g5834 ( n14253 , n9972 , n11997 );
    or g5835 ( n9382 , n1741 , n5290 );
    or g5836 ( n5955 , n14088 , n10210 );
    nor g5837 ( n13538 , n3602 , n11044 );
    not g5838 ( n1760 , n2040 );
    nor g5839 ( n1604 , n8701 , n9037 );
    and g5840 ( n13804 , n10367 , n14043 );
    or g5841 ( n13401 , n974 , n9219 );
    and g5842 ( n1980 , n7427 , n415 );
    or g5843 ( n12207 , n11171 , n12493 );
    and g5844 ( n9659 , n4692 , n9452 );
    not g5845 ( n9577 , n3345 );
    and g5846 ( n1069 , n8431 , n11873 );
    nor g5847 ( n4272 , n3768 , n10340 );
    and g5848 ( n12048 , n1117 , n8174 );
    or g5849 ( n26 , n2149 , n3303 );
    or g5850 ( n6078 , n11405 , n3605 );
    or g5851 ( n7690 , n5548 , n2007 );
    and g5852 ( n581 , n4525 , n181 );
    or g5853 ( n3634 , n8517 , n5003 );
    nor g5854 ( n3694 , n4313 , n10739 );
    and g5855 ( n290 , n2533 , n12529 );
    and g5856 ( n10392 , n9069 , n11271 );
    and g5857 ( n5778 , n8066 , n6886 );
    or g5858 ( n5752 , n7887 , n3677 );
    not g5859 ( n4162 , n6123 );
    or g5860 ( n14288 , n7888 , n12789 );
    or g5861 ( n7829 , n6867 , n7381 );
    and g5862 ( n8859 , n13379 , n7732 );
    and g5863 ( n3459 , n11028 , n7323 );
    nor g5864 ( n12670 , n1383 , n4375 );
    not g5865 ( n7618 , n702 );
    and g5866 ( n13872 , n9238 , n323 );
    not g5867 ( n11470 , n4296 );
    not g5868 ( n9494 , n674 );
    not g5869 ( n11704 , n8735 );
    or g5870 ( n4055 , n5861 , n9281 );
    or g5871 ( n3236 , n11542 , n4193 );
    and g5872 ( n14422 , n9188 , n4473 );
    not g5873 ( n4880 , n6990 );
    not g5874 ( n7900 , n9236 );
    and g5875 ( n13582 , n12542 , n8940 );
    nor g5876 ( n13947 , n13707 , n6813 );
    and g5877 ( n9470 , n2758 , n10982 );
    and g5878 ( n1743 , n10084 , n8278 );
    and g5879 ( n5355 , n10084 , n9861 );
    and g5880 ( n62 , n5348 , n8834 );
    and g5881 ( n13253 , n7443 , n12004 );
    and g5882 ( n11063 , n7443 , n1077 );
    or g5883 ( n2976 , n5139 , n1673 );
    and g5884 ( n4658 , n808 , n11061 );
    and g5885 ( n1794 , n10072 , n4431 );
    and g5886 ( n13302 , n4509 , n11705 );
    or g5887 ( n8608 , n782 , n325 );
    and g5888 ( n4604 , n8302 , n12440 );
    and g5889 ( n9023 , n8066 , n9670 );
    and g5890 ( n10692 , n7427 , n13680 );
    or g5891 ( n269 , n7249 , n10726 );
    not g5892 ( n10363 , n3742 );
    nor g5893 ( n10627 , n13675 , n7072 );
    or g5894 ( n10488 , n185 , n5503 );
    and g5895 ( n5187 , n5011 , n1386 );
    and g5896 ( n2298 , n4382 , n10830 );
    and g5897 ( n624 , n6343 , n10443 );
    or g5898 ( n9880 , n8210 , n1298 );
    and g5899 ( n1732 , n4614 , n2077 );
    or g5900 ( n11234 , n7912 , n12314 );
    or g5901 ( n2982 , n11909 , n9399 );
    and g5902 ( n8132 , n14351 , n10427 );
    nor g5903 ( n13661 , n5780 , n10106 );
    nor g5904 ( n6421 , n6428 , n7955 );
    or g5905 ( n1396 , n10024 , n11205 );
    not g5906 ( n11040 , n5195 );
    or g5907 ( n6074 , n8635 , n13814 );
    or g5908 ( n7017 , n6242 , n12649 );
    not g5909 ( n1881 , n6603 );
    nor g5910 ( n12165 , n2597 , n11915 );
    nor g5911 ( n11727 , n3287 , n3214 );
    not g5912 ( n9721 , n10400 );
    or g5913 ( n11448 , n6373 , n8546 );
    not g5914 ( n5695 , n10204 );
    and g5915 ( n8711 , n4546 , n14066 );
    or g5916 ( n6454 , n3134 , n13777 );
    or g5917 ( n3136 , n13130 , n14456 );
    or g5918 ( n9320 , n8304 , n4214 );
    and g5919 ( n13715 , n10247 , n13468 );
    or g5920 ( n1207 , n12821 , n11167 );
    or g5921 ( n9014 , n14337 , n12563 );
    or g5922 ( n4665 , n10383 , n14314 );
    nor g5923 ( n11023 , n12197 , n13474 );
    nor g5924 ( n12878 , n14166 , n2125 );
    or g5925 ( n13766 , n9111 , n1350 );
    not g5926 ( n8923 , n2432 );
    or g5927 ( n1510 , n12400 , n1969 );
    nor g5928 ( n186 , n4210 , n2695 );
    not g5929 ( n13641 , n5108 );
    or g5930 ( n4504 , n11285 , n6932 );
    and g5931 ( n10108 , n13230 , n398 );
    and g5932 ( n7786 , n12741 , n8226 );
    and g5933 ( n12408 , n965 , n6923 );
    nor g5934 ( n6833 , n4439 , n14333 );
    and g5935 ( n5149 , n14178 , n1850 );
    or g5936 ( n7189 , n3164 , n401 );
    or g5937 ( n9769 , n13420 , n10466 );
    not g5938 ( n9265 , n7621 );
    or g5939 ( n822 , n6730 , n2728 );
    and g5940 ( n6467 , n5062 , n1579 );
    nor g5941 ( n3859 , n13759 , n9615 );
    and g5942 ( n8587 , n1414 , n6494 );
    not g5943 ( n11435 , n12757 );
    nor g5944 ( n10014 , n9577 , n7437 );
    or g5945 ( n13762 , n3527 , n2143 );
    or g5946 ( n10993 , n4562 , n12293 );
    or g5947 ( n7402 , n6260 , n11930 );
    and g5948 ( n6332 , n6844 , n937 );
    and g5949 ( n14452 , n1520 , n1179 );
    or g5950 ( n5369 , n11739 , n2689 );
    and g5951 ( n7279 , n7419 , n5134 );
    nor g5952 ( n5720 , n13677 , n6760 );
    nor g5953 ( n8796 , n2057 , n12876 );
    and g5954 ( n10966 , n6507 , n2625 );
    nor g5955 ( n13352 , n7011 , n3719 );
    and g5956 ( n4538 , n222 , n6834 );
    or g5957 ( n3221 , n10245 , n10996 );
    not g5958 ( n4614 , n7808 );
    or g5959 ( n198 , n361 , n738 );
    and g5960 ( n12073 , n8768 , n3933 );
    not g5961 ( n9856 , n10985 );
    and g5962 ( n12719 , n4722 , n4667 );
    nor g5963 ( n7876 , n648 , n8603 );
    or g5964 ( n5523 , n12130 , n9223 );
    not g5965 ( n4851 , n14133 );
    not g5966 ( n12100 , n1966 );
    or g5967 ( n1933 , n4807 , n13241 );
    or g5968 ( n7562 , n7011 , n2121 );
    or g5969 ( n7559 , n11935 , n7777 );
    nor g5970 ( n4231 , n5569 , n9475 );
    or g5971 ( n1130 , n3273 , n455 );
    not g5972 ( n12248 , n7521 );
    and g5973 ( n11030 , n12425 , n6568 );
    or g5974 ( n4800 , n13854 , n25 );
    or g5975 ( n14315 , n9780 , n2568 );
    or g5976 ( n4062 , n4508 , n1316 );
    and g5977 ( n8759 , n6830 , n9988 );
    and g5978 ( n3155 , n2012 , n10079 );
    and g5979 ( n13480 , n8512 , n9068 );
    and g5980 ( n14307 , n6480 , n7631 );
    or g5981 ( n1819 , n8908 , n12715 );
    or g5982 ( n10764 , n7426 , n5262 );
    not g5983 ( n4289 , n2497 );
    and g5984 ( n10125 , n2983 , n7565 );
    or g5985 ( n14083 , n12622 , n14502 );
    or g5986 ( n3722 , n11542 , n7786 );
    and g5987 ( n7413 , n10302 , n10369 );
    and g5988 ( n14199 , n14327 , n9488 );
    nor g5989 ( n12330 , n11489 , n2623 );
    and g5990 ( n7071 , n14408 , n12708 );
    and g5991 ( n9609 , n4422 , n8437 );
    and g5992 ( n152 , n7079 , n1014 );
    and g5993 ( n6553 , n8432 , n4274 );
    and g5994 ( n8035 , n4692 , n6252 );
    or g5995 ( n13898 , n2645 , n3397 );
    or g5996 ( n8442 , n7697 , n6203 );
    and g5997 ( n4419 , n12037 , n5321 );
    or g5998 ( n3574 , n9269 , n9405 );
    or g5999 ( n979 , n4828 , n2935 );
    or g6000 ( n13757 , n9429 , n13138 );
    or g6001 ( n1816 , n523 , n11012 );
    nor g6002 ( n6246 , n1028 , n6488 );
    and g6003 ( n7770 , n12531 , n2546 );
    and g6004 ( n11514 , n11484 , n8270 );
    or g6005 ( n12050 , n4967 , n11215 );
    or g6006 ( n3562 , n12130 , n7540 );
    not g6007 ( n11935 , n11788 );
    or g6008 ( n7181 , n3512 , n2459 );
    or g6009 ( n13380 , n6288 , n9326 );
    or g6010 ( n883 , n10019 , n5109 );
    nor g6011 ( n14488 , n228 , n12891 );
    and g6012 ( n9796 , n10374 , n10757 );
    or g6013 ( n12302 , n5493 , n460 );
    not g6014 ( n1559 , n5467 );
    or g6015 ( n14470 , n6242 , n6823 );
    nor g6016 ( n1251 , n10973 , n10431 );
    or g6017 ( n8703 , n9211 , n3897 );
    and g6018 ( n4268 , n11313 , n1438 );
    and g6019 ( n1402 , n9724 , n8063 );
    and g6020 ( n4540 , n13359 , n3751 );
    and g6021 ( n5370 , n2904 , n10086 );
    or g6022 ( n1605 , n6711 , n4364 );
    or g6023 ( n6037 , n2897 , n4456 );
    or g6024 ( n9671 , n2562 , n1641 );
    and g6025 ( n10664 , n2064 , n4778 );
    and g6026 ( n13494 , n5471 , n7828 );
    nor g6027 ( n8090 , n8301 , n5599 );
    or g6028 ( n7048 , n6205 , n3306 );
    or g6029 ( n1815 , n13477 , n8953 );
    or g6030 ( n1936 , n1640 , n3972 );
    or g6031 ( n14274 , n8277 , n12520 );
    not g6032 ( n9111 , n2472 );
    or g6033 ( n3053 , n8825 , n3571 );
    nor g6034 ( n11745 , n9340 , n6087 );
    not g6035 ( n9724 , n3967 );
    nor g6036 ( n878 , n7756 , n3817 );
    and g6037 ( n1832 , n11636 , n3476 );
    and g6038 ( n13439 , n13520 , n2606 );
    nor g6039 ( n11543 , n4624 , n7372 );
    or g6040 ( n4557 , n4313 , n3632 );
    nor g6041 ( n489 , n7980 , n9059 );
    not g6042 ( n8197 , n7710 );
    not g6043 ( n10059 , n11605 );
    or g6044 ( n1983 , n13112 , n12309 );
    or g6045 ( n35 , n4407 , n6146 );
    or g6046 ( n4021 , n6607 , n3384 );
    or g6047 ( n11202 , n7736 , n13702 );
    or g6048 ( n1594 , n9151 , n1201 );
    and g6049 ( n10033 , n10930 , n5331 );
    not g6050 ( n3546 , n3046 );
    or g6051 ( n969 , n14188 , n13708 );
    and g6052 ( n13398 , n638 , n14317 );
    and g6053 ( n14440 , n10922 , n3554 );
    and g6054 ( n1148 , n10084 , n5424 );
    or g6055 ( n7376 , n2804 , n5009 );
    not g6056 ( n521 , n14011 );
    and g6057 ( n4541 , n5184 , n8051 );
    not g6058 ( n3876 , n10864 );
    and g6059 ( n10908 , n718 , n1207 );
    and g6060 ( n12140 , n11748 , n10040 );
    nor g6061 ( n13628 , n6000 , n3517 );
    and g6062 ( n2775 , n80 , n6272 );
    or g6063 ( n13830 , n12994 , n4457 );
    and g6064 ( n14207 , n8025 , n1661 );
    or g6065 ( n8203 , n9931 , n7279 );
    or g6066 ( n3662 , n1701 , n14050 );
    and g6067 ( n12769 , n5471 , n7342 );
    and g6068 ( n14085 , n12455 , n14266 );
    and g6069 ( n10925 , n1775 , n11632 );
    and g6070 ( n4891 , n5788 , n8682 );
    or g6071 ( n5200 , n4195 , n10570 );
    or g6072 ( n3051 , n769 , n12887 );
    or g6073 ( n6427 , n8897 , n11106 );
    nor g6074 ( n8861 , n14198 , n3848 );
    not g6075 ( n12636 , n13636 );
    or g6076 ( n5310 , n4684 , n5696 );
    not g6077 ( n9140 , n4203 );
    or g6078 ( n250 , n361 , n11124 );
    and g6079 ( n9056 , n231 , n11906 );
    not g6080 ( n8106 , n9924 );
    and g6081 ( n2632 , n8569 , n8316 );
    nor g6082 ( n9566 , n4771 , n11762 );
    and g6083 ( n2374 , n1924 , n10850 );
    not g6084 ( n11017 , n13206 );
    or g6085 ( n2072 , n4602 , n9947 );
    and g6086 ( n8839 , n13700 , n3109 );
    not g6087 ( n4347 , n6657 );
    and g6088 ( n13212 , n7391 , n2870 );
    and g6089 ( n653 , n3710 , n5910 );
    or g6090 ( n1885 , n11090 , n6301 );
    or g6091 ( n8031 , n573 , n3584 );
    or g6092 ( n8614 , n7812 , n7285 );
    not g6093 ( n1136 , n13295 );
    and g6094 ( n13126 , n9885 , n9278 );
    or g6095 ( n12458 , n12994 , n7939 );
    nor g6096 ( n3749 , n8877 , n1411 );
    or g6097 ( n7534 , n1582 , n5607 );
    or g6098 ( n3381 , n6428 , n516 );
    and g6099 ( n9510 , n11300 , n11288 );
    and g6100 ( n4034 , n7691 , n13051 );
    and g6101 ( n14181 , n14450 , n3996 );
    not g6102 ( n2738 , n7904 );
    or g6103 ( n402 , n8304 , n1779 );
    or g6104 ( n2968 , n13446 , n5685 );
    not g6105 ( n9941 , n12142 );
    and g6106 ( n7214 , n6744 , n13125 );
    or g6107 ( n10443 , n2562 , n1466 );
    nor g6108 ( n7207 , n1685 , n13300 );
    and g6109 ( n14505 , n11674 , n9055 );
    not g6110 ( n1911 , n10341 );
    and g6111 ( n7172 , n5475 , n7579 );
    not g6112 ( n13863 , n3313 );
    or g6113 ( n2264 , n2531 , n9104 );
    or g6114 ( n525 , n7914 , n3189 );
    nor g6115 ( n4368 , n10858 , n3996 );
    and g6116 ( n1665 , n7392 , n2356 );
    or g6117 ( n12402 , n6690 , n7951 );
    and g6118 ( n2215 , n3401 , n6740 );
    not g6119 ( n13154 , n2778 );
    not g6120 ( n7781 , n650 );
    or g6121 ( n2232 , n14472 , n9524 );
    or g6122 ( n10623 , n14107 , n3121 );
    and g6123 ( n1893 , n4358 , n3847 );
    and g6124 ( n10582 , n10815 , n7297 );
    or g6125 ( n13920 , n523 , n2084 );
    or g6126 ( n10772 , n1006 , n13851 );
    or g6127 ( n5854 , n329 , n10305 );
    and g6128 ( n13207 , n5591 , n8088 );
    and g6129 ( n9706 , n12475 , n7137 );
    or g6130 ( n5120 , n8748 , n10260 );
    or g6131 ( n8694 , n8490 , n2429 );
    or g6132 ( n9183 , n12549 , n7306 );
    and g6133 ( n7765 , n4354 , n13393 );
    and g6134 ( n5624 , n5092 , n4056 );
    and g6135 ( n7441 , n1076 , n1045 );
    and g6136 ( n13272 , n286 , n1746 );
    and g6137 ( n2717 , n8620 , n11473 );
    and g6138 ( n8836 , n14150 , n4560 );
    and g6139 ( n2464 , n986 , n969 );
    or g6140 ( n2921 , n10731 , n7400 );
    or g6141 ( n10442 , n12047 , n10085 );
    or g6142 ( n10298 , n7887 , n5584 );
    nor g6143 ( n1627 , n10368 , n4705 );
    not g6144 ( n10079 , n666 );
    or g6145 ( n13247 , n12494 , n10375 );
    or g6146 ( n8790 , n12625 , n3992 );
    not g6147 ( n3577 , n5631 );
    and g6148 ( n2391 , n11470 , n9120 );
    and g6149 ( n1214 , n7822 , n2609 );
    not g6150 ( n14260 , n7902 );
    nor g6151 ( n9690 , n355 , n3619 );
    and g6152 ( n13006 , n12721 , n11746 );
    and g6153 ( n7815 , n7419 , n9960 );
    not g6154 ( n14109 , n5268 );
    or g6155 ( n2208 , n2315 , n6845 );
    or g6156 ( n13277 , n9864 , n13703 );
    or g6157 ( n5302 , n5997 , n11912 );
    nor g6158 ( n8612 , n12069 , n8090 );
    or g6159 ( n3489 , n5695 , n6866 );
    and g6160 ( n12535 , n2201 , n12718 );
    or g6161 ( n11286 , n13432 , n505 );
    or g6162 ( n12663 , n555 , n5355 );
    or g6163 ( n12437 , n3193 , n3795 );
    or g6164 ( n12138 , n5266 , n4921 );
    or g6165 ( n14498 , n69 , n4642 );
    or g6166 ( n11921 , n12543 , n417 );
    or g6167 ( n1890 , n7697 , n5081 );
    and g6168 ( n9636 , n7443 , n14519 );
    or g6169 ( n13662 , n781 , n13763 );
    nor g6170 ( n13030 , n7886 , n5192 );
    not g6171 ( n8361 , n6714 );
    nor g6172 ( n11531 , n4988 , n1902 );
    and g6173 ( n210 , n11262 , n6087 );
    or g6174 ( n12263 , n9218 , n1848 );
    or g6175 ( n538 , n6629 , n3740 );
    not g6176 ( n6629 , n3284 );
    or g6177 ( n1755 , n9803 , n9830 );
    nor g6178 ( n4471 , n30 , n4704 );
    or g6179 ( n841 , n5007 , n10513 );
    or g6180 ( n7632 , n6695 , n4060 );
    or g6181 ( n7728 , n3877 , n4449 );
    or g6182 ( n3593 , n9035 , n11772 );
    or g6183 ( n3118 , n11090 , n13899 );
    or g6184 ( n12062 , n12139 , n10359 );
    and g6185 ( n5598 , n2058 , n7632 );
    or g6186 ( n6998 , n89 , n2359 );
    and g6187 ( n9872 , n5823 , n2499 );
    and g6188 ( n8236 , n406 , n13346 );
    and g6189 ( n6800 , n6343 , n11876 );
    and g6190 ( n3077 , n8047 , n5020 );
    and g6191 ( n6461 , n5053 , n367 );
    and g6192 ( n1408 , n7043 , n2765 );
    or g6193 ( n8981 , n14319 , n10057 );
    or g6194 ( n13654 , n11315 , n11976 );
    and g6195 ( n6942 , n10854 , n7671 );
    not g6196 ( n8021 , n11244 );
    nor g6197 ( n3730 , n4877 , n6712 );
    and g6198 ( n9431 , n3526 , n2896 );
    not g6199 ( n6471 , n4609 );
    not g6200 ( n13213 , n9987 );
    and g6201 ( n7730 , n9726 , n4942 );
    nor g6202 ( n9714 , n13087 , n10483 );
    and g6203 ( n4679 , n9297 , n3257 );
    and g6204 ( n4288 , n4844 , n11561 );
    and g6205 ( n6061 , n13252 , n5017 );
    nor g6206 ( n1822 , n1617 , n13810 );
    and g6207 ( n6308 , n6023 , n2475 );
    nor g6208 ( n7709 , n10036 , n1042 );
    or g6209 ( n13580 , n13501 , n10175 );
    nor g6210 ( n2813 , n827 , n6906 );
    and g6211 ( n4517 , n2583 , n3960 );
    or g6212 ( n441 , n7551 , n9566 );
    or g6213 ( n6982 , n12428 , n5241 );
    and g6214 ( n3643 , n8702 , n5097 );
    or g6215 ( n435 , n9111 , n4273 );
    and g6216 ( n6116 , n1136 , n2802 );
    or g6217 ( n14395 , n7438 , n9662 );
    or g6218 ( n8618 , n3047 , n13174 );
    or g6219 ( n5316 , n10626 , n12750 );
    and g6220 ( n7657 , n5434 , n12862 );
    or g6221 ( n2165 , n12091 , n13473 );
    and g6222 ( n6057 , n3952 , n9536 );
    not g6223 ( n7755 , n12658 );
    or g6224 ( n10261 , n6706 , n13907 );
    or g6225 ( n12244 , n11875 , n4117 );
    not g6226 ( n3926 , n11001 );
    and g6227 ( n860 , n428 , n13598 );
    or g6228 ( n384 , n12034 , n12731 );
    and g6229 ( n5696 , n14120 , n11450 );
    and g6230 ( n12874 , n1936 , n13270 );
    nor g6231 ( n2584 , n31 , n6502 );
    nor g6232 ( n10856 , n11558 , n1064 );
    or g6233 ( n14090 , n2318 , n5374 );
    nor g6234 ( n11766 , n14466 , n9295 );
    or g6235 ( n5781 , n7887 , n5593 );
    and g6236 ( n9357 , n12461 , n2032 );
    and g6237 ( n8508 , n3813 , n1647 );
    and g6238 ( n13729 , n2942 , n5390 );
    or g6239 ( n13216 , n12075 , n10906 );
    nor g6240 ( n7890 , n1458 , n6963 );
    not g6241 ( n3768 , n11308 );
    or g6242 ( n4864 , n8242 , n14343 );
    nor g6243 ( n11046 , n1628 , n9359 );
    nor g6244 ( n1472 , n8404 , n12021 );
    or g6245 ( n6587 , n7418 , n4283 );
    or g6246 ( n1916 , n12353 , n14391 );
    and g6247 ( n6939 , n3942 , n3469 );
    and g6248 ( n990 , n7970 , n4194 );
    and g6249 ( n12310 , n4502 , n9738 );
    not g6250 ( n7308 , n8397 );
    and g6251 ( n4351 , n4261 , n9293 );
    and g6252 ( n8371 , n6754 , n14211 );
    and g6253 ( n1110 , n5458 , n1654 );
    not g6254 ( n7345 , n11218 );
    nor g6255 ( n1017 , n3905 , n3321 );
    nor g6256 ( n6906 , n2790 , n12678 );
    not g6257 ( n957 , n6555 );
    or g6258 ( n6084 , n4045 , n720 );
    and g6259 ( n1619 , n3268 , n11877 );
    and g6260 ( n1529 , n13433 , n13052 );
    nor g6261 ( n13049 , n6041 , n14047 );
    and g6262 ( n3992 , n7327 , n790 );
    and g6263 ( n5773 , n12472 , n3288 );
    and g6264 ( n8579 , n13860 , n13973 );
    or g6265 ( n3337 , n12400 , n9073 );
    nor g6266 ( n4536 , n13707 , n9948 );
    or g6267 ( n5083 , n504 , n10242 );
    nor g6268 ( n9909 , n11980 , n10347 );
    and g6269 ( n12689 , n2998 , n4150 );
    not g6270 ( n12455 , n11870 );
    or g6271 ( n11473 , n5414 , n12270 );
    or g6272 ( n5865 , n9285 , n14346 );
    not g6273 ( n12087 , n10917 );
    and g6274 ( n7860 , n7370 , n3188 );
    or g6275 ( n14387 , n5647 , n735 );
    and g6276 ( n3818 , n1729 , n8549 );
    nor g6277 ( n11267 , n2017 , n6889 );
    or g6278 ( n3866 , n7076 , n8258 );
    or g6279 ( n3537 , n1602 , n12407 );
    and g6280 ( n5045 , n1074 , n13015 );
    or g6281 ( n7095 , n10394 , n13034 );
    and g6282 ( n8380 , n2281 , n3192 );
    nor g6283 ( n11791 , n12453 , n9239 );
    not g6284 ( n2281 , n2752 );
    and g6285 ( n11753 , n8358 , n3618 );
    nor g6286 ( n2396 , n1480 , n13519 );
    or g6287 ( n11519 , n7754 , n7889 );
    or g6288 ( n9851 , n4508 , n258 );
    or g6289 ( n3030 , n10396 , n3417 );
    and g6290 ( n6604 , n7063 , n3363 );
    and g6291 ( n12314 , n2064 , n7737 );
    or g6292 ( n6970 , n4239 , n3482 );
    and g6293 ( n2449 , n4880 , n9503 );
    not g6294 ( n13021 , n12345 );
    not g6295 ( n11033 , n9414 );
    or g6296 ( n8477 , n11176 , n13701 );
    and g6297 ( n4377 , n11748 , n2815 );
    and g6298 ( n1646 , n4546 , n8263 );
    and g6299 ( n9902 , n11316 , n9389 );
    and g6300 ( n5408 , n3635 , n9343 );
    and g6301 ( n9310 , n9853 , n423 );
    or g6302 ( n13100 , n3126 , n826 );
    or g6303 ( n12223 , n6271 , n8674 );
    and g6304 ( n13909 , n12250 , n1826 );
    and g6305 ( n8430 , n6724 , n12361 );
    not g6306 ( n7227 , n6264 );
    nor g6307 ( n2195 , n11481 , n1492 );
    and g6308 ( n12747 , n8923 , n5328 );
    and g6309 ( n9453 , n1421 , n298 );
    not g6310 ( n13978 , n3681 );
    or g6311 ( n12590 , n2149 , n11557 );
    and g6312 ( n2519 , n14313 , n6580 );
    and g6313 ( n12928 , n7026 , n11843 );
    or g6314 ( n2585 , n11090 , n8484 );
    and g6315 ( n5946 , n8147 , n13380 );
    and g6316 ( n10591 , n3910 , n1546 );
    nor g6317 ( n9787 , n8877 , n1859 );
    not g6318 ( n10647 , n1378 );
    and g6319 ( n5571 , n718 , n13027 );
    and g6320 ( n6069 , n5062 , n5099 );
    or g6321 ( n11598 , n5603 , n1948 );
    not g6322 ( n2924 , n5046 );
    or g6323 ( n10173 , n13547 , n607 );
    or g6324 ( n8233 , n9245 , n9110 );
    not g6325 ( n11614 , n6743 );
    or g6326 ( n133 , n4207 , n9135 );
    or g6327 ( n8987 , n2055 , n3103 );
    or g6328 ( n4945 , n9035 , n7393 );
    not g6329 ( n6753 , n7808 );
    and g6330 ( n1488 , n10855 , n3515 );
    and g6331 ( n12430 , n1011 , n4564 );
    not g6332 ( n7605 , n9677 );
    and g6333 ( n1515 , n103 , n12537 );
    not g6334 ( n2624 , n1908 );
    or g6335 ( n2203 , n4978 , n6151 );
    and g6336 ( n25 , n10566 , n11103 );
    not g6337 ( n1904 , n12697 );
    not g6338 ( n8183 , n8122 );
    and g6339 ( n12550 , n11411 , n1096 );
    and g6340 ( n14048 , n9345 , n12411 );
    or g6341 ( n12788 , n2694 , n10334 );
    and g6342 ( n12746 , n56 , n201 );
    not g6343 ( n11687 , n6114 );
    and g6344 ( n13057 , n6316 , n12495 );
    and g6345 ( n365 , n9745 , n50 );
    or g6346 ( n13985 , n11953 , n10119 );
    and g6347 ( n379 , n550 , n13539 );
    or g6348 ( n10674 , n11951 , n3919 );
    and g6349 ( n8308 , n6316 , n7848 );
    or g6350 ( n6812 , n850 , n10388 );
    and g6351 ( n7183 , n225 , n1692 );
    not g6352 ( n9913 , n5683 );
    and g6353 ( n4235 , n1193 , n6431 );
    not g6354 ( n2387 , n8272 );
    and g6355 ( n6863 , n11336 , n993 );
    and g6356 ( n12172 , n13823 , n10971 );
    and g6357 ( n3006 , n3743 , n4817 );
    and g6358 ( n4558 , n4788 , n14092 );
    or g6359 ( n8725 , n10083 , n12561 );
    and g6360 ( n6164 , n13780 , n1088 );
    or g6361 ( n5413 , n5480 , n3947 );
    or g6362 ( n10286 , n6690 , n13497 );
    and g6363 ( n5820 , n9275 , n13792 );
    not g6364 ( n9703 , n8672 );
    or g6365 ( n12950 , n3888 , n14353 );
    and g6366 ( n11330 , n7909 , n7858 );
    or g6367 ( n9200 , n1576 , n4731 );
    and g6368 ( n14206 , n9824 , n4717 );
    and g6369 ( n11172 , n4655 , n4140 );
    nor g6370 ( n12666 , n5118 , n1767 );
    or g6371 ( n2673 , n5936 , n2534 );
    and g6372 ( n2545 , n12397 , n6928 );
    nor g6373 ( n725 , n9806 , n14526 );
    or g6374 ( n14128 , n2057 , n9155 );
    and g6375 ( n2008 , n13641 , n6202 );
    and g6376 ( n14391 , n14327 , n9756 );
    not g6377 ( n1447 , n9921 );
    and g6378 ( n8195 , n8386 , n5909 );
    nor g6379 ( n8953 , n13394 , n3730 );
    nor g6380 ( n12447 , n4953 , n11068 );
    or g6381 ( n5426 , n4840 , n13065 );
    and g6382 ( n7470 , n8769 , n3098 );
    or g6383 ( n8362 , n8821 , n12123 );
    or g6384 ( n1490 , n11438 , n12834 );
    or g6385 ( n8718 , n1805 , n5592 );
    and g6386 ( n10270 , n11816 , n8038 );
    not g6387 ( n9541 , n4720 );
    and g6388 ( n8689 , n1354 , n745 );
    and g6389 ( n1007 , n7187 , n2481 );
    or g6390 ( n11037 , n10539 , n6470 );
    and g6391 ( n11156 , n6167 , n8951 );
    not g6392 ( n8213 , n10377 );
    or g6393 ( n11876 , n2562 , n6171 );
    or g6394 ( n13921 , n492 , n608 );
    or g6395 ( n12144 , n954 , n10708 );
    nor g6396 ( n9732 , n11628 , n6405 );
    not g6397 ( n8353 , n3572 );
    and g6398 ( n1868 , n6640 , n1203 );
    nor g6399 ( n9888 , n5977 , n3014 );
    not g6400 ( n4897 , n749 );
    or g6401 ( n13902 , n6867 , n3500 );
    nor g6402 ( n11977 , n3922 , n12116 );
    or g6403 ( n2013 , n11176 , n1150 );
    and g6404 ( n13200 , n1247 , n2441 );
    nor g6405 ( n789 , n906 , n8594 );
    and g6406 ( n1454 , n6013 , n5589 );
    or g6407 ( n1548 , n13882 , n6680 );
    nor g6408 ( n13530 , n2415 , n4438 );
    or g6409 ( n4253 , n3219 , n10631 );
    nor g6410 ( n9586 , n8580 , n11778 );
    and g6411 ( n11174 , n8786 , n1322 );
    nor g6412 ( n12099 , n10323 , n9612 );
    and g6413 ( n4237 , n9238 , n1034 );
    or g6414 ( n14217 , n4562 , n1723 );
    or g6415 ( n5984 , n5936 , n2295 );
    not g6416 ( n1613 , n4606 );
    nor g6417 ( n488 , n584 , n2999 );
    and g6418 ( n13427 , n2099 , n6458 );
    or g6419 ( n612 , n8620 , n2674 );
    or g6420 ( n2375 , n6046 , n11525 );
    or g6421 ( n998 , n8821 , n6612 );
    nor g6422 ( n8982 , n10254 , n3890 );
    or g6423 ( n12393 , n6596 , n2022 );
    or g6424 ( n10991 , n10245 , n10968 );
    or g6425 ( n9032 , n10857 , n13788 );
    and g6426 ( n1405 , n11213 , n13198 );
    or g6427 ( n925 , n12295 , n3746 );
    and g6428 ( n5311 , n13676 , n4950 );
    not g6429 ( n12779 , n10080 );
    and g6430 ( n4184 , n7852 , n1446 );
    nor g6431 ( n7913 , n7973 , n2303 );
    and g6432 ( n12373 , n13626 , n13578 );
    or g6433 ( n2050 , n14107 , n4081 );
    or g6434 ( n11098 , n1480 , n11069 );
    and g6435 ( n8366 , n5857 , n4814 );
    not g6436 ( n5936 , n3007 );
    and g6437 ( n13855 , n3952 , n6783 );
    or g6438 ( n7423 , n12820 , n13769 );
    or g6439 ( n2393 , n3826 , n8259 );
    and g6440 ( n756 , n14091 , n4883 );
    not g6441 ( n13968 , n13224 );
    and g6442 ( n8810 , n13745 , n6236 );
    and g6443 ( n6496 , n3277 , n452 );
    and g6444 ( n11477 , n2310 , n7341 );
    or g6445 ( n13861 , n3886 , n9651 );
    nor g6446 ( n8670 , n2969 , n9493 );
    and g6447 ( n14415 , n9726 , n10505 );
    or g6448 ( n10198 , n7171 , n5046 );
    not g6449 ( n1342 , n10603 );
    and g6450 ( n6095 , n12101 , n7984 );
    and g6451 ( n12003 , n2099 , n814 );
    nor g6452 ( n6221 , n6768 , n903 );
    and g6453 ( n10680 , n8432 , n13187 );
    not g6454 ( n10323 , n2320 );
    nor g6455 ( n5170 , n2781 , n9520 );
    not g6456 ( n7370 , n12872 );
    and g6457 ( n12577 , n12159 , n7082 );
    and g6458 ( n4553 , n3169 , n13724 );
    and g6459 ( n12610 , n687 , n3856 );
    or g6460 ( n4311 , n320 , n12927 );
    and g6461 ( n5422 , n1140 , n938 );
    or g6462 ( n4922 , n12019 , n10769 );
    and g6463 ( n14436 , n5582 , n13323 );
    not g6464 ( n3800 , n10069 );
    or g6465 ( n5596 , n13511 , n13364 );
    or g6466 ( n1243 , n10147 , n14464 );
    and g6467 ( n3812 , n12209 , n8134 );
    and g6468 ( n10780 , n13464 , n143 );
    or g6469 ( n3590 , n7438 , n7269 );
    and g6470 ( n12806 , n4803 , n2265 );
    nor g6471 ( n6449 , n7115 , n9031 );
    and g6472 ( n13750 , n12057 , n10195 );
    not g6473 ( n13190 , n739 );
    or g6474 ( n8016 , n9442 , n12434 );
    not g6475 ( n10622 , n10975 );
    and g6476 ( n10599 , n4098 , n2915 );
    and g6477 ( n5737 , n9811 , n1643 );
    or g6478 ( n11095 , n100 , n939 );
    or g6479 ( n9043 , n4602 , n2337 );
    nor g6480 ( n613 , n5468 , n12312 );
    not g6481 ( n5234 , n3455 );
    and g6482 ( n8079 , n7053 , n1992 );
    and g6483 ( n14247 , n10622 , n1581 );
    nor g6484 ( n11246 , n10837 , n6418 );
    or g6485 ( n9068 , n8726 , n5383 );
    and g6486 ( n13311 , n10084 , n1698 );
    or g6487 ( n9488 , n11360 , n5579 );
    or g6488 ( n4702 , n7888 , n14081 );
    and g6489 ( n9684 , n6531 , n8833 );
    and g6490 ( n8099 , n1100 , n10073 );
    or g6491 ( n4816 , n11438 , n10503 );
    or g6492 ( n40 , n12549 , n2622 );
    not g6493 ( n10179 , n7027 );
    or g6494 ( n8351 , n4162 , n5811 );
    not g6495 ( n14213 , n13219 );
    and g6496 ( n5269 , n3204 , n7728 );
    and g6497 ( n9987 , n12636 , n7811 );
    not g6498 ( n2218 , n9959 );
    not g6499 ( n6830 , n1771 );
    and g6500 ( n13459 , n10678 , n209 );
    and g6501 ( n10849 , n14038 , n6996 );
    nor g6502 ( n11910 , n5715 , n6667 );
    not g6503 ( n9956 , n10147 );
    or g6504 ( n12156 , n8527 , n12128 );
    nor g6505 ( n578 , n2766 , n3566 );
    and g6506 ( n13658 , n7282 , n1277 );
    and g6507 ( n7258 , n3628 , n8970 );
    nor g6508 ( n10390 , n7900 , n6279 );
    or g6509 ( n338 , n6695 , n4937 );
    or g6510 ( n5787 , n3512 , n3915 );
    or g6511 ( n1302 , n12622 , n4841 );
    and g6512 ( n8595 , n2772 , n1334 );
    and g6513 ( n2459 , n7026 , n5111 );
    not g6514 ( n12428 , n8148 );
    nor g6515 ( n7582 , n10402 , n3235 );
    and g6516 ( n9208 , n14227 , n507 );
    not g6517 ( n13722 , n4646 );
    and g6518 ( n4811 , n10516 , n4402 );
    or g6519 ( n9010 , n11576 , n12980 );
    and g6520 ( n909 , n11411 , n12555 );
    nor g6521 ( n4653 , n13675 , n12120 );
    and g6522 ( n7907 , n2177 , n5557 );
    nor g6523 ( n5006 , n9984 , n6124 );
    or g6524 ( n11119 , n13718 , n10578 );
    or g6525 ( n10971 , n8986 , n4758 );
    not g6526 ( n1312 , n11305 );
    or g6527 ( n11208 , n11036 , n182 );
    and g6528 ( n10724 , n129 , n7774 );
    not g6529 ( n3132 , n12776 );
    and g6530 ( n8848 , n7429 , n11785 );
    or g6531 ( n507 , n8748 , n9632 );
    and g6532 ( n11282 , n5489 , n9430 );
    and g6533 ( n7126 , n4806 , n13861 );
    and g6534 ( n7851 , n10457 , n12329 );
    and g6535 ( n4919 , n12475 , n3083 );
    nor g6536 ( n413 , n2417 , n10329 );
    and g6537 ( n5874 , n5458 , n12491 );
    not g6538 ( n8866 , n5077 );
    or g6539 ( n14121 , n1028 , n14172 );
    nor g6540 ( n7927 , n3354 , n13089 );
    nor g6541 ( n5469 , n1844 , n1527 );
    and g6542 ( n2589 , n4844 , n5025 );
    and g6543 ( n9246 , n12015 , n11734 );
    nor g6544 ( n8186 , n13081 , n13352 );
    nor g6545 ( n12155 , n7551 , n9630 );
    not g6546 ( n11647 , n2130 );
    or g6547 ( n3617 , n5234 , n14437 );
    and g6548 ( n3868 , n405 , n4992 );
    or g6549 ( n6293 , n12020 , n9661 );
    and g6550 ( n5580 , n1804 , n10741 );
    nor g6551 ( n3338 , n5118 , n878 );
    or g6552 ( n12908 , n2246 , n3945 );
    not g6553 ( n5997 , n751 );
    and g6554 ( n2372 , n1431 , n9000 );
    and g6555 ( n314 , n4546 , n9688 );
    or g6556 ( n11792 , n9119 , n2895 );
    or g6557 ( n1579 , n9780 , n11243 );
    nor g6558 ( n6444 , n4978 , n4760 );
    not g6559 ( n317 , n622 );
    not g6560 ( n14210 , n7941 );
    and g6561 ( n14003 , n5240 , n8050 );
    and g6562 ( n7016 , n5940 , n12319 );
    and g6563 ( n13301 , n12265 , n8175 );
    or g6564 ( n9670 , n4052 , n3180 );
    or g6565 ( n13982 , n1391 , n4332 );
    nor g6566 ( n10607 , n9984 , n9701 );
    and g6567 ( n13499 , n2224 , n2920 );
    nor g6568 ( n10492 , n3132 , n8473 );
    and g6569 ( n7509 , n2465 , n7901 );
    or g6570 ( n4179 , n1535 , n3000 );
    and g6571 ( n14026 , n11093 , n3221 );
    or g6572 ( n2079 , n9931 , n12859 );
    or g6573 ( n99 , n13509 , n2201 );
    nor g6574 ( n818 , n1693 , n2631 );
    and g6575 ( n11102 , n1427 , n9505 );
    or g6576 ( n4883 , n3273 , n6433 );
    and g6577 ( n4380 , n432 , n88 );
    and g6578 ( n8102 , n7053 , n1644 );
    nor g6579 ( n11410 , n4248 , n6268 );
    and g6580 ( n6394 , n13641 , n12793 );
    or g6581 ( n3301 , n387 , n2594 );
    or g6582 ( n4242 , n2181 , n9872 );
    or g6583 ( n3347 , n3134 , n12231 );
    not g6584 ( n10254 , n4966 );
    or g6585 ( n7741 , n8986 , n12684 );
    not g6586 ( n5977 , n382 );
    nor g6587 ( n12539 , n3873 , n705 );
    nor g6588 ( n4673 , n10593 , n7695 );
    and g6589 ( n9399 , n3607 , n1569 );
    and g6590 ( n9982 , n13107 , n3124 );
    and g6591 ( n9798 , n10969 , n7726 );
    or g6592 ( n4497 , n2412 , n9930 );
    or g6593 ( n2274 , n49 , n8275 );
    or g6594 ( n5097 , n49 , n2641 );
    or g6595 ( n3216 , n11047 , n6935 );
    or g6596 ( n187 , n7358 , n9648 );
    not g6597 ( n1804 , n10372 );
    or g6598 ( n13731 , n4602 , n7049 );
    not g6599 ( n1685 , n622 );
    or g6600 ( n1166 , n7684 , n2578 );
    or g6601 ( n3058 , n7359 , n14467 );
    or g6602 ( n832 , n1582 , n13564 );
    not g6603 ( n9226 , n5242 );
    not g6604 ( n7216 , n2454 );
    or g6605 ( n12722 , n6629 , n8414 );
    nor g6606 ( n2798 , n8825 , n1385 );
    or g6607 ( n9551 , n11171 , n4597 );
    nor g6608 ( n2036 , n14135 , n11757 );
    not g6609 ( n1520 , n10036 );
    or g6610 ( n12482 , n781 , n8430 );
    or g6611 ( n5903 , n3877 , n5244 );
    or g6612 ( n275 , n14430 , n10162 );
    or g6613 ( n5776 , n8828 , n9822 );
    nor g6614 ( n2390 , n7227 , n8199 );
    or g6615 ( n14305 , n3559 , n3872 );
    and g6616 ( n14467 , n10338 , n12214 );
    and g6617 ( n5374 , n6531 , n6896 );
    and g6618 ( n1228 , n11220 , n832 );
    or g6619 ( n13033 , n4502 , n2201 );
    nor g6620 ( n6630 , n4049 , n13183 );
    and g6621 ( n381 , n1225 , n11751 );
    or g6622 ( n11145 , n7527 , n11896 );
    and g6623 ( n1730 , n7677 , n7528 );
    or g6624 ( n8883 , n2510 , n10652 );
    not g6625 ( n11011 , n7404 );
    or g6626 ( n10500 , n1602 , n14034 );
    or g6627 ( n6004 , n1261 , n7994 );
    or g6628 ( n10018 , n568 , n2581 );
    or g6629 ( n3060 , n1494 , n2826 );
    or g6630 ( n9361 , n11459 , n5731 );
    and g6631 ( n7287 , n4289 , n3343 );
    not g6632 ( n9266 , n12506 );
    or g6633 ( n6241 , n11551 , n2119 );
    nor g6634 ( n4280 , n2098 , n6443 );
    not g6635 ( n6941 , n12322 );
    or g6636 ( n3985 , n4899 , n4249 );
    or g6637 ( n3687 , n11722 , n13144 );
    not g6638 ( n11440 , n12746 );
    not g6639 ( n14273 , n3893 );
    and g6640 ( n3744 , n12730 , n10764 );
    not g6641 ( n8232 , n8048 );
    or g6642 ( n4429 , n3193 , n3957 );
    or g6643 ( n4685 , n1137 , n5004 );
    and g6644 ( n13587 , n533 , n9095 );
    and g6645 ( n11043 , n12335 , n6587 );
    and g6646 ( n13075 , n1431 , n5079 );
    or g6647 ( n2765 , n49 , n11185 );
    and g6648 ( n8676 , n8111 , n704 );
    not g6649 ( n9450 , n6248 );
    and g6650 ( n3713 , n6724 , n3688 );
    or g6651 ( n7889 , n10765 , n4154 );
    and g6652 ( n6769 , n13489 , n4665 );
    or g6653 ( n14176 , n9747 , n13994 );
    or g6654 ( n12481 , n2897 , n2936 );
    or g6655 ( n2244 , n6891 , n3026 );
    not g6656 ( n1924 , n3344 );
    and g6657 ( n11962 , n8932 , n10916 );
    or g6658 ( n4717 , n13432 , n2939 );
    not g6659 ( n2017 , n13668 );
    and g6660 ( n6774 , n12475 , n6035 );
    or g6661 ( n6412 , n14029 , n6666 );
    and g6662 ( n6505 , n333 , n4006 );
    and g6663 ( n7246 , n13093 , n578 );
    nor g6664 ( n3177 , n2677 , n12667 );
    and g6665 ( n5529 , n12018 , n4823 );
    and g6666 ( n10932 , n12772 , n2043 );
    and g6667 ( n738 , n10589 , n6021 );
    and g6668 ( n11917 , n98 , n8325 );
    and g6669 ( n6784 , n8066 , n9791 );
    and g6670 ( n6339 , n4276 , n10884 );
    or g6671 ( n13483 , n5450 , n13170 );
    or g6672 ( n10538 , n11953 , n4127 );
    nor g6673 ( n6949 , n7739 , n8139 );
    and g6674 ( n213 , n4289 , n1800 );
    and g6675 ( n12961 , n10229 , n2263 );
    or g6676 ( n131 , n766 , n1543 );
    or g6677 ( n11320 , n12112 , n12327 );
    and g6678 ( n4937 , n13359 , n11263 );
    and g6679 ( n13243 , n12185 , n11133 );
    or g6680 ( n12344 , n7076 , n2721 );
    or g6681 ( n5114 , n4498 , n14129 );
    nor g6682 ( n1411 , n7660 , n6583 );
    or g6683 ( n14338 , n8575 , n4426 );
    not g6684 ( n6743 , n13725 );
    nor g6685 ( n12865 , n6953 , n10464 );
    and g6686 ( n1445 , n6135 , n2803 );
    nor g6687 ( n828 , n1820 , n3262 );
    or g6688 ( n5420 , n10913 , n570 );
    and g6689 ( n11958 , n4856 , n12662 );
    or g6690 ( n2131 , n7156 , n6708 );
    not g6691 ( n5144 , n426 );
    or g6692 ( n3892 , n1914 , n8137 );
    nor g6693 ( n13508 , n4233 , n13145 );
    and g6694 ( n12887 , n6354 , n569 );
    nor g6695 ( n13648 , n9818 , n13325 );
    nor g6696 ( n6476 , n14419 , n13538 );
    or g6697 ( n30 , n4659 , n12573 );
    or g6698 ( n9296 , n11121 , n8074 );
    and g6699 ( n14035 , n10678 , n4023 );
    and g6700 ( n10362 , n5764 , n5594 );
    not g6701 ( n12069 , n8927 );
    and g6702 ( n14122 , n1662 , n12307 );
    not g6703 ( n5855 , n13511 );
    and g6704 ( n11795 , n11336 , n633 );
    or g6705 ( n3684 , n361 , n4677 );
    and g6706 ( n3787 , n2367 , n6796 );
    and g6707 ( n9736 , n8213 , n1037 );
    and g6708 ( n10606 , n14109 , n6173 );
    not g6709 ( n1137 , n1041 );
    or g6710 ( n2237 , n13074 , n2616 );
    or g6711 ( n10543 , n6730 , n4139 );
    and g6712 ( n13423 , n5779 , n13797 );
    and g6713 ( n3142 , n5137 , n1005 );
    or g6714 ( n520 , n13220 , n8676 );
    and g6715 ( n3471 , n6838 , n12913 );
    nor g6716 ( n8547 , n2251 , n9376 );
    and g6717 ( n13701 , n9315 , n11049 );
    nor g6718 ( n13997 , n6797 , n7876 );
    and g6719 ( n10419 , n13700 , n10417 );
    and g6720 ( n9139 , n9824 , n6549 );
    and g6721 ( n13858 , n1278 , n1958 );
    and g6722 ( n6826 , n5038 , n13366 );
    and g6723 ( n10812 , n14327 , n5248 );
    not g6724 ( n4646 , n4135 );
    and g6725 ( n13395 , n11406 , n10614 );
    and g6726 ( n7553 , n14063 , n14438 );
    or g6727 ( n1903 , n5695 , n8556 );
    or g6728 ( n13955 , n8714 , n10685 );
    or g6729 ( n9676 , n172 , n7317 );
    and g6730 ( n9073 , n3565 , n7892 );
    and g6731 ( n12098 , n6016 , n5817 );
    not g6732 ( n8507 , n12885 );
    or g6733 ( n11378 , n10825 , n14422 );
    and g6734 ( n3584 , n3 , n980 );
    not g6735 ( n13081 , n12580 );
    not g6736 ( n6046 , n4149 );
    or g6737 ( n10976 , n12994 , n9409 );
    and g6738 ( n987 , n6023 , n1054 );
    or g6739 ( n6097 , n2784 , n8102 );
    or g6740 ( n1496 , n1189 , n5054 );
    or g6741 ( n10429 , n4840 , n6394 );
    not g6742 ( n11980 , n6978 );
    not g6743 ( n7250 , n3284 );
    and g6744 ( n13465 , n13246 , n7243 );
    and g6745 ( n6722 , n9232 , n1664 );
    and g6746 ( n4579 , n9052 , n641 );
    not g6747 ( n6052 , n6874 );
    and g6748 ( n11347 , n12391 , n6368 );
    or g6749 ( n13809 , n12211 , n4222 );
    not g6750 ( n1775 , n3402 );
    not g6751 ( n13226 , n1267 );
    or g6752 ( n6267 , n10024 , n397 );
    and g6753 ( n12033 , n2724 , n6503 );
    nor g6754 ( n9039 , n7887 , n13414 );
    not g6755 ( n4978 , n8695 );
    and g6756 ( n6960 , n12935 , n13191 );
    and g6757 ( n3613 , n11484 , n1599 );
    or g6758 ( n12729 , n10913 , n9949 );
    and g6759 ( n6759 , n11838 , n3842 );
    and g6760 ( n12509 , n11702 , n11897 );
    or g6761 ( n13888 , n2901 , n7235 );
    not g6762 ( n1086 , n4595 );
    and g6763 ( n2407 , n10147 , n4671 );
    not g6764 ( n12229 , n1843 );
    or g6765 ( n1562 , n2510 , n4029 );
    not g6766 ( n11180 , n8704 );
    or g6767 ( n12581 , n2946 , n5418 );
    not g6768 ( n7145 , n7291 );
    or g6769 ( n5863 , n6971 , n852 );
    or g6770 ( n8267 , n5144 , n8294 );
    or g6771 ( n6170 , n7116 , n13963 );
    or g6772 ( n8560 , n4435 , n5560 );
    or g6773 ( n13305 , n2518 , n13503 );
    or g6774 ( n3430 , n5732 , n6069 );
    and g6775 ( n736 , n13840 , n177 );
    not g6776 ( n3491 , n9818 );
    not g6777 ( n4713 , n2731 );
    and g6778 ( n10199 , n11838 , n2031 );
    or g6779 ( n10847 , n9230 , n4775 );
    or g6780 ( n12082 , n12543 , n6226 );
    and g6781 ( n7316 , n7081 , n2259 );
    or g6782 ( n11083 , n12844 , n12598 );
    or g6783 ( n10063 , n9375 , n14460 );
    and g6784 ( n12587 , n6899 , n689 );
    nor g6785 ( n3541 , n11111 , n165 );
    not g6786 ( n13413 , n9596 );
    and g6787 ( n9149 , n10247 , n14030 );
    not g6788 ( n2505 , n1763 );
    or g6789 ( n1328 , n7684 , n6995 );
    or g6790 ( n1692 , n8821 , n12277 );
    or g6791 ( n3550 , n4128 , n12735 );
    not g6792 ( n12193 , n10465 );
    nor g6793 ( n8590 , n7075 , n2844 );
    not g6794 ( n11576 , n1041 );
    or g6795 ( n1200 , n14058 , n6752 );
    not g6796 ( n49 , n9306 );
    nor g6797 ( n10287 , n10688 , n723 );
    not g6798 ( n7291 , n10803 );
    and g6799 ( n7925 , n6981 , n10672 );
    not g6800 ( n1417 , n3324 );
    and g6801 ( n10693 , n3424 , n14100 );
    not g6802 ( n6907 , n12580 );
    or g6803 ( n5858 , n7527 , n466 );
    and g6804 ( n10156 , n12038 , n4987 );
    or g6805 ( n5286 , n12295 , n7620 );
    and g6806 ( n5176 , n13069 , n13827 );
    and g6807 ( n7059 , n10763 , n1999 );
    or g6808 ( n4113 , n1112 , n7457 );
    nor g6809 ( n11987 , n14296 , n7791 );
    not g6810 ( n10834 , n751 );
    and g6811 ( n396 , n9705 , n7046 );
    and g6812 ( n936 , n222 , n9075 );
    or g6813 ( n3538 , n1202 , n1145 );
    and g6814 ( n11027 , n8401 , n3016 );
    not g6815 ( n7171 , n4039 );
    and g6816 ( n6105 , n13877 , n675 );
    not g6817 ( n11438 , n10346 );
    and g6818 ( n3950 , n12265 , n12049 );
    or g6819 ( n229 , n8304 , n9762 );
    or g6820 ( n10158 , n3120 , n3039 );
    not g6821 ( n3952 , n10828 );
    and g6822 ( n10874 , n13525 , n8541 );
    and g6823 ( n5054 , n1231 , n8367 );
    or g6824 ( n3929 , n14521 , n7832 );
    and g6825 ( n3821 , n14109 , n1921 );
    or g6826 ( n11511 , n7781 , n9252 );
    or g6827 ( n8667 , n2531 , n13066 );
    and g6828 ( n6940 , n11329 , n10671 );
    or g6829 ( n4814 , n283 , n4753 );
    and g6830 ( n10920 , n12461 , n4310 );
    and g6831 ( n4462 , n12101 , n5363 );
    or g6832 ( n7510 , n976 , n11201 );
    or g6833 ( n4533 , n14009 , n2048 );
    or g6834 ( n3150 , n7898 , n3111 );
    not g6835 ( n9046 , n2298 );
    and g6836 ( n12608 , n10032 , n291 );
    or g6837 ( n8814 , n9142 , n6460 );
    not g6838 ( n5647 , n4939 );
    not g6839 ( n4509 , n1178 );
    and g6840 ( n5102 , n11403 , n10853 );
    not g6841 ( n2973 , n9414 );
    or g6842 ( n5662 , n11704 , n120 );
    or g6843 ( n6725 , n6607 , n13812 );
    and g6844 ( n10547 , n12202 , n12413 );
    and g6845 ( n7645 , n1678 , n556 );
    and g6846 ( n7093 , n8855 , n10023 );
    not g6847 ( n9778 , n742 );
    or g6848 ( n9786 , n5454 , n8405 );
    or g6849 ( n12603 , n7736 , n8195 );
    or g6850 ( n8700 , n12047 , n6415 );
    or g6851 ( n2408 , n8821 , n7460 );
    and g6852 ( n3837 , n12953 , n7564 );
    or g6853 ( n7097 , n5493 , n12623 );
    not g6854 ( n12132 , n8302 );
    not g6855 ( n1610 , n2692 );
    or g6856 ( n1366 , n10154 , n831 );
    or g6857 ( n12559 , n13118 , n385 );
    and g6858 ( n3503 , n12105 , n5259 );
    or g6859 ( n2290 , n11360 , n4380 );
    or g6860 ( n13453 , n10781 , n14414 );
    or g6861 ( n7047 , n14198 , n9307 );
    or g6862 ( n855 , n12034 , n597 );
    and g6863 ( n5501 , n10209 , n8488 );
    and g6864 ( n13853 , n3367 , n2768 );
    or g6865 ( n4496 , n6428 , n2283 );
    and g6866 ( n12748 , n2547 , n4940 );
    and g6867 ( n10915 , n7667 , n12790 );
    or g6868 ( n7465 , n10871 , n1832 );
    nor g6869 ( n4654 , n6000 , n9552 );
    and g6870 ( n7821 , n11157 , n4480 );
    and g6871 ( n7328 , n9113 , n8610 );
    nor g6872 ( n13950 , n1944 , n9303 );
    nor g6873 ( n13124 , n12046 , n8312 );
    and g6874 ( n12624 , n12101 , n7151 );
    or g6875 ( n3251 , n14282 , n13744 );
    or g6876 ( n3646 , n10449 , n10490 );
    and g6877 ( n1583 , n8066 , n8477 );
    not g6878 ( n7043 , n10269 );
    and g6879 ( n13322 , n8702 , n1889 );
    not g6880 ( n4544 , n7875 );
    or g6881 ( n7373 , n69 , n1164 );
    or g6882 ( n961 , n5266 , n5061 );
    and g6883 ( n9179 , n11028 , n1845 );
    and g6884 ( n2700 , n1255 , n3183 );
    and g6885 ( n14190 , n3724 , n11690 );
    or g6886 ( n3699 , n4791 , n1583 );
    or g6887 ( n12839 , n3125 , n3513 );
    or g6888 ( n6032 , n13005 , n7698 );
    not g6889 ( n11315 , n7339 );
    or g6890 ( n556 , n7971 , n3576 );
    not g6891 ( n4092 , n565 );
    or g6892 ( n6376 , n1576 , n11398 );
    nor g6893 ( n5864 , n13394 , n8943 );
    and g6894 ( n5437 , n14388 , n3604 );
    and g6895 ( n2753 , n1678 , n12473 );
    or g6896 ( n1078 , n12077 , n6917 );
    not g6897 ( n748 , n2497 );
    and g6898 ( n11398 , n1100 , n9320 );
    and g6899 ( n1847 , n2378 , n12559 );
    not g6900 ( n10731 , n9846 );
    not g6901 ( n1140 , n11969 );
    and g6902 ( n6772 , n4486 , n7626 );
    or g6903 ( n2363 , n1821 , n5351 );
    or g6904 ( n3683 , n6730 , n13369 );
    and g6905 ( n4408 , n10909 , n1249 );
    or g6906 ( n13149 , n387 , n4001 );
    or g6907 ( n9964 , n7122 , n10174 );
    and g6908 ( n8823 , n13860 , n11720 );
    and g6909 ( n3849 , n5764 , n11658 );
    and g6910 ( n9513 , n12101 , n3811 );
    not g6911 ( n6829 , n4379 );
    or g6912 ( n6266 , n8552 , n9589 );
    and g6913 ( n2620 , n14446 , n13699 );
    and g6914 ( n5763 , n5348 , n4592 );
    not g6915 ( n5064 , n6978 );
    or g6916 ( n10881 , n817 , n6771 );
    or g6917 ( n8495 , n11379 , n6333 );
    and g6918 ( n3707 , n965 , n4204 );
    and g6919 ( n5027 , n3370 , n1562 );
    not g6920 ( n48 , n777 );
    and g6921 ( n8774 , n8358 , n9263 );
    or g6922 ( n11263 , n1198 , n3643 );
    or g6923 ( n2213 , n9151 , n8130 );
    and g6924 ( n10160 , n13555 , n3575 );
    and g6925 ( n2534 , n10822 , n13457 );
    nor g6926 ( n14047 , n1028 , n5712 );
    not g6927 ( n14525 , n11401 );
    and g6928 ( n4143 , n2564 , n3404 );
    and g6929 ( n9641 , n8401 , n5781 );
    or g6930 ( n433 , n1147 , n5743 );
    and g6931 ( n14232 , n15 , n10674 );
    and g6932 ( n9153 , n10399 , n5464 );
    or g6933 ( n1889 , n10396 , n3518 );
    and g6934 ( n1735 , n11313 , n4327 );
    or g6935 ( n1216 , n5641 , n2374 );
    and g6936 ( n8468 , n5317 , n9411 );
    or g6937 ( n11885 , n3449 , n650 );
    and g6938 ( n3841 , n6754 , n13277 );
    not g6939 ( n4602 , n7441 );
    or g6940 ( n10786 , n10461 , n3601 );
    and g6941 ( n5816 , n1610 , n5971 );
    and g6942 ( n9715 , n13338 , n11354 );
    and g6943 ( n10870 , n12449 , n4748 );
    and g6944 ( n1948 , n12389 , n5928 );
    nor g6945 ( n12170 , n11498 , n8551 );
    not g6946 ( n10828 , n210 );
    or g6947 ( n7442 , n5483 , n11030 );
    not g6948 ( n10231 , n13093 );
    or g6949 ( n1442 , n11572 , n3718 );
    or g6950 ( n6824 , n3809 , n1835 );
    and g6951 ( n13743 , n13484 , n9731 );
    or g6952 ( n927 , n3888 , n1326 );
    not g6953 ( n7011 , n7289 );
    or g6954 ( n6129 , n12764 , n1435 );
    and g6955 ( n11517 , n12620 , n11019 );
    or g6956 ( n11927 , n3271 , n74 );
    and g6957 ( n9467 , n3986 , n11598 );
    nor g6958 ( n1762 , n6052 , n602 );
    or g6959 ( n10435 , n4978 , n343 );
    and g6960 ( n9058 , n5823 , n4825 );
    and g6961 ( n6746 , n9885 , n2959 );
    and g6962 ( n2266 , n1876 , n5377 );
    or g6963 ( n1967 , n7803 , n7242 );
    or g6964 ( n1474 , n8480 , n7344 );
    or g6965 ( n10068 , n5625 , n8206 );
    and g6966 ( n6227 , n7943 , n7310 );
    not g6967 ( n6271 , n409 );
    nor g6968 ( n14508 , n8458 , n1344 );
    nor g6969 ( n3651 , n1929 , n6875 );
    and g6970 ( n8585 , n12105 , n1275 );
    or g6971 ( n4686 , n1711 , n2038 );
    and g6972 ( n4599 , n2322 , n8140 );
    or g6973 ( n11632 , n3871 , n11042 );
    and g6974 ( n1897 , n10330 , n14158 );
    and g6975 ( n8977 , n10166 , n1166 );
    not g6976 ( n350 , n8315 );
    and g6977 ( n4324 , n7934 , n1793 );
    or g6978 ( n6615 , n11704 , n4930 );
    nor g6979 ( n12966 , n8277 , n9606 );
    and g6980 ( n12958 , n3710 , n10412 );
    or g6981 ( n1357 , n10378 , n10080 );
    not g6982 ( n2949 , n5901 );
    nor g6983 ( n13266 , n5944 , n11862 );
    or g6984 ( n971 , n8332 , n7172 );
    nor g6985 ( n11069 , n11546 , n11812 );
    nor g6986 ( n4366 , n3394 , n4252 );
    and g6987 ( n3796 , n2006 , n3270 );
    or g6988 ( n3390 , n13413 , n6153 );
    or g6989 ( n12629 , n10624 , n12985 );
    not g6990 ( n4481 , n9846 );
    or g6991 ( n14147 , n13118 , n6250 );
    and g6992 ( n1169 , n12741 , n1020 );
    or g6993 ( n7398 , n390 , n11327 );
    and g6994 ( n6894 , n6486 , n12696 );
    not g6995 ( n9416 , n10115 );
    or g6996 ( n1139 , n6867 , n9659 );
    and g6997 ( n437 , n12475 , n6615 );
    and g6998 ( n6988 , n2904 , n4367 );
    and g6999 ( n14507 , n11153 , n1809 );
    and g7000 ( n8260 , n4581 , n10131 );
    or g7001 ( n10669 , n2149 , n4187 );
    not g7002 ( n12527 , n6254 );
    nor g7003 ( n2512 , n8656 , n9147 );
    and g7004 ( n6588 , n3586 , n11208 );
    or g7005 ( n5797 , n11360 , n11322 );
    and g7006 ( n4881 , n2998 , n9854 );
    and g7007 ( n1331 , n11737 , n10517 );
    and g7008 ( n7028 , n3204 , n1367 );
    or g7009 ( n13621 , n8304 , n4454 );
    not g7010 ( n10377 , n8003 );
    not g7011 ( n9388 , n2520 );
    not g7012 ( n11950 , n12503 );
    or g7013 ( n10903 , n4199 , n10602 );
    and g7014 ( n2482 , n3672 , n8032 );
    and g7015 ( n4465 , n11188 , n772 );
    and g7016 ( n2324 , n783 , n953 );
    not g7017 ( n11680 , n4786 );
    and g7018 ( n2782 , n15 , n12804 );
    and g7019 ( n1587 , n9745 , n5510 );
    or g7020 ( n11175 , n4967 , n11925 );
    not g7021 ( n7156 , n7339 );
    not g7022 ( n7327 , n12904 );
    not g7023 ( n12280 , n3587 );
    and g7024 ( n3478 , n2521 , n3843 );
    or g7025 ( n5699 , n11581 , n3209 );
    and g7026 ( n10448 , n8147 , n3073 );
    and g7027 ( n4783 , n783 , n3490 );
    and g7028 ( n1150 , n8183 , n9425 );
    not g7029 ( n10360 , n12782 );
    or g7030 ( n1683 , n2878 , n10691 );
    and g7031 ( n6255 , n9238 , n13563 );
    and g7032 ( n4539 , n13240 , n3979 );
    and g7033 ( n7054 , n6697 , n7034 );
    or g7034 ( n13716 , n6109 , n6359 );
    and g7035 ( n5151 , n6909 , n6185 );
    or g7036 ( n21 , n11839 , n9208 );
    and g7037 ( n11447 , n8213 , n503 );
    or g7038 ( n10221 , n13531 , n11893 );
    nor g7039 ( n11999 , n10289 , n1251 );
    not g7040 ( n5512 , n4659 );
    and g7041 ( n2794 , n5416 , n6705 );
    not g7042 ( n69 , n11055 );
    and g7043 ( n5862 , n428 , n4182 );
    not g7044 ( n6731 , n4708 );
    and g7045 ( n10525 , n8431 , n2216 );
    or g7046 ( n2839 , n13477 , n5034 );
    and g7047 ( n8011 , n7079 , n9758 );
    or g7048 ( n9777 , n13005 , n2806 );
    or g7049 ( n7984 , n5833 , n4903 );
    or g7050 ( n9894 , n10913 , n10695 );
    not g7051 ( n1401 , n10470 );
    not g7052 ( n3724 , n5618 );
    or g7053 ( n11769 , n14401 , n6759 );
    or g7054 ( n10000 , n14065 , n13944 );
    and g7055 ( n3502 , n1857 , n5749 );
    and g7056 ( n7733 , n14465 , n13524 );
    nor g7057 ( n558 , n7146 , n7281 );
    or g7058 ( n3083 , n1838 , n8070 );
    nor g7059 ( n9493 , n4195 , n5022 );
    not g7060 ( n6838 , n7902 );
    and g7061 ( n12863 , n3247 , n5369 );
    or g7062 ( n6688 , n5891 , n8836 );
    or g7063 ( n13900 , n7401 , n8873 );
    or g7064 ( n12709 , n3394 , n11432 );
    and g7065 ( n14414 , n10647 , n11448 );
    not g7066 ( n3922 , n2816 );
    nor g7067 ( n12912 , n3530 , n9707 );
    and g7068 ( n1449 , n5279 , n6581 );
    and g7069 ( n265 , n7673 , n6998 );
    and g7070 ( n5756 , n7612 , n14283 );
    or g7071 ( n189 , n5409 , n7214 );
    nor g7072 ( n10519 , n6088 , n10774 );
    or g7073 ( n14514 , n523 , n7680 );
    not g7074 ( n13784 , n14133 );
    not g7075 ( n1378 , n14071 );
    or g7076 ( n5615 , n8592 , n13462 );
    and g7077 ( n2864 , n12057 , n1922 );
    or g7078 ( n6983 , n511 , n7311 );
    not g7079 ( n2888 , n11331 );
    nor g7080 ( n1818 , n12999 , n11198 );
    or g7081 ( n14491 , n4357 , n502 );
    or g7082 ( n3763 , n2318 , n9381 );
    and g7083 ( n4448 , n5779 , n3699 );
    or g7084 ( n9599 , n1051 , n3064 );
    or g7085 ( n5331 , n5695 , n8426 );
    not g7086 ( n10399 , n5182 );
    or g7087 ( n14335 , n11909 , n7287 );
    or g7088 ( n1029 , n13531 , n10576 );
    or g7089 ( n6458 , n11722 , n7561 );
    not g7090 ( n10177 , n14071 );
    or g7091 ( n13783 , n12047 , n2365 );
    and g7092 ( n5687 , n4803 , n9020 );
    or g7093 ( n11941 , n13547 , n5933 );
    and g7094 ( n9942 , n14093 , n8284 );
    or g7095 ( n833 , n7426 , n11694 );
    and g7096 ( n13878 , n6243 , n12663 );
    or g7097 ( n1671 , n4092 , n1464 );
    or g7098 ( n7868 , n3062 , n6902 );
    or g7099 ( n4735 , n6629 , n10043 );
    nor g7100 ( n9439 , n11581 , n1463 );
    and g7101 ( n2705 , n533 , n13794 );
    or g7102 ( n6420 , n2694 , n11968 );
    and g7103 ( n8597 , n9890 , n10117 );
    or g7104 ( n3133 , n13707 , n9476 );
    not g7105 ( n3234 , n2788 );
    and g7106 ( n4227 , n5553 , n7446 );
    and g7107 ( n9469 , n1428 , n10957 );
    and g7108 ( n11808 , n12039 , n2399 );
    or g7109 ( n830 , n4807 , n10610 );
    or g7110 ( n14031 , n3608 , n12025 );
    nor g7111 ( n6887 , n2341 , n12099 );
    not g7112 ( n4018 , n2432 );
    or g7113 ( n3808 , n11171 , n3123 );
    nor g7114 ( n7661 , n5569 , n12666 );
    or g7115 ( n9876 , n12131 , n10101 );
    and g7116 ( n11817 , n3212 , n3304 );
    or g7117 ( n7749 , n6288 , n13025 );
    and g7118 ( n12551 , n4156 , n9781 );
    and g7119 ( n9889 , n6822 , n11380 );
    not g7120 ( n11412 , n13213 );
    and g7121 ( n1043 , n14042 , n13921 );
    or g7122 ( n3208 , n747 , n9023 );
    and g7123 ( n14191 , n1788 , n3023 );
    or g7124 ( n60 , n10224 , n3647 );
    or g7125 ( n1253 , n4162 , n13106 );
    and g7126 ( n4976 , n7961 , n9868 );
    nor g7127 ( n4664 , n9577 , n11796 );
    and g7128 ( n2865 , n7079 , n10218 );
    not g7129 ( n6990 , n4966 );
    or g7130 ( n7922 , n4822 , n7236 );
    not g7131 ( n3015 , n9810 );
    not g7132 ( n13476 , n3870 );
    not g7133 ( n11163 , n1955 );
    and g7134 ( n3455 , n6903 , n10751 );
    not g7135 ( n1339 , n9613 );
    and g7136 ( n10721 , n8630 , n6353 );
    or g7137 ( n13957 , n3320 , n11555 );
    and g7138 ( n14061 , n8300 , n7492 );
    not g7139 ( n5710 , n2794 );
    and g7140 ( n9883 , n2583 , n12803 );
    not g7141 ( n1414 , n6559 );
    and g7142 ( n1469 , n7963 , n11981 );
    or g7143 ( n8819 , n6428 , n5387 );
    and g7144 ( n4563 , n6649 , n10118 );
    or g7145 ( n9425 , n954 , n12145 );
    nor g7146 ( n12749 , n478 , n11747 );
    or g7147 ( n14148 , n7862 , n13054 );
    and g7148 ( n12924 , n1640 , n7590 );
    not g7149 ( n11852 , n3130 );
    or g7150 ( n8760 , n5362 , n13459 );
    and g7151 ( n12111 , n12852 , n9837 );
    not g7152 ( n11969 , n1079 );
    and g7153 ( n6295 , n14150 , n5804 );
    and g7154 ( n11499 , n9113 , n8266 );
    or g7155 ( n3067 , n820 , n9812 );
    nor g7156 ( n10475 , n3546 , n4782 );
    and g7157 ( n12258 , n432 , n1572 );
    and g7158 ( n4516 , n2445 , n3144 );
    not g7159 ( n8605 , n6829 );
    or g7160 ( n2546 , n2686 , n9348 );
    nor g7161 ( n7474 , n438 , n396 );
    nor g7162 ( n4848 , n1023 , n4090 );
    and g7163 ( n8978 , n7826 , n639 );
    and g7164 ( n1670 , n646 , n1971 );
    and g7165 ( n6185 , n9941 , n12126 );
    or g7166 ( n7412 , n11303 , n6836 );
    and g7167 ( n7163 , n6606 , n5689 );
    nor g7168 ( n13807 , n8816 , n13526 );
    and g7169 ( n8091 , n2099 , n13971 );
    or g7170 ( n1475 , n10713 , n2775 );
    and g7171 ( n5438 , n1278 , n14023 );
    nor g7172 ( n6513 , n11628 , n6300 );
    nor g7173 ( n312 , n1722 , n13993 );
    and g7174 ( n4298 , n8247 , n10995 );
    and g7175 ( n7032 , n3846 , n7805 );
    or g7176 ( n4748 , n7697 , n9383 );
    or g7177 ( n2217 , n3193 , n2364 );
    and g7178 ( n14041 , n533 , n14409 );
    and g7179 ( n5060 , n4806 , n5403 );
    not g7180 ( n3672 , n13383 );
    or g7181 ( n14291 , n9442 , n12660 );
    not g7182 ( n13072 , n12897 );
    or g7183 ( n3692 , n3134 , n9886 );
    and g7184 ( n7088 , n6957 , n12545 );
    or g7185 ( n9935 , n2510 , n10592 );
    and g7186 ( n1143 , n9275 , n9319 );
    and g7187 ( n892 , n8393 , n2507 );
    not g7188 ( n11259 , n6364 );
    nor g7189 ( n8334 , n9967 , n13842 );
    not g7190 ( n239 , n5306 );
    nor g7191 ( n10604 , n14466 , n8984 );
    or g7192 ( n652 , n12968 , n5126 );
    not g7193 ( n5278 , n7704 );
    and g7194 ( n543 , n5185 , n4035 );
    and g7195 ( n13554 , n4932 , n14008 );
    not g7196 ( n492 , n1010 );
    and g7197 ( n995 , n2006 , n10868 );
    and g7198 ( n3215 , n10820 , n11863 );
    and g7199 ( n6698 , n8183 , n12144 );
    nor g7200 ( n1553 , n2822 , n6456 );
    or g7201 ( n8461 , n12351 , n7251 );
    and g7202 ( n11684 , n4018 , n1229 );
    and g7203 ( n4214 , n6898 , n11692 );
    and g7204 ( n6314 , n6999 , n10290 );
    or g7205 ( n13449 , n4876 , n12110 );
    or g7206 ( n6523 , n10083 , n11740 );
    nor g7207 ( n5966 , n14466 , n3844 );
    nor g7208 ( n11165 , n9423 , n360 );
    and g7209 ( n3591 , n12611 , n13865 );
    nor g7210 ( n9631 , n8353 , n3510 );
    and g7211 ( n9773 , n9724 , n13431 );
    or g7212 ( n3096 , n11551 , n2385 );
    or g7213 ( n4623 , n3320 , n12465 );
    not g7214 ( n10099 , n14524 );
    nor g7215 ( n2543 , n4200 , n8671 );
    or g7216 ( n13643 , n14107 , n7547 );
    nor g7217 ( n2617 , n619 , n10481 );
    and g7218 ( n12422 , n8697 , n12732 );
    and g7219 ( n8483 , n10763 , n12429 );
    not g7220 ( n10760 , n10573 );
    not g7221 ( n11406 , n2497 );
    nor g7222 ( n8784 , n13435 , n1234 );
    nor g7223 ( n1004 , n1838 , n11280 );
    not g7224 ( n1539 , n1342 );
    or g7225 ( n13819 , n348 , n8439 );
    and g7226 ( n6150 , n12015 , n7019 );
    or g7227 ( n4246 , n317 , n365 );
    and g7228 ( n7857 , n11422 , n12518 );
    and g7229 ( n14402 , n1428 , n3430 );
    and g7230 ( n11537 , n9726 , n1605 );
    and g7231 ( n8120 , n1775 , n13288 );
    and g7232 ( n8523 , n646 , n9415 );
    or g7233 ( n3465 , n7609 , n4656 );
    or g7234 ( n6500 , n11123 , n4084 );
    and g7235 ( n1622 , n501 , n8478 );
    and g7236 ( n12011 , n10032 , n5254 );
    or g7237 ( n851 , n11510 , n13040 );
    or g7238 ( n11334 , n227 , n8972 );
    nor g7239 ( n1839 , n7809 , n7277 );
    and g7240 ( n8272 , n8822 , n5412 );
    and g7241 ( n1793 , n14521 , n659 );
    and g7242 ( n6825 , n9265 , n8416 );
    or g7243 ( n2613 , n11647 , n1799 );
    not g7244 ( n6909 , n3388 );
    or g7245 ( n12281 , n194 , n5565 );
    not g7246 ( n9972 , n10469 );
    not g7247 ( n9807 , n11813 );
    and g7248 ( n1406 , n3861 , n8170 );
    nor g7249 ( n2990 , n7662 , n7843 );
    nor g7250 ( n10542 , n12112 , n1798 );
    and g7251 ( n635 , n10854 , n9204 );
    and g7252 ( n4971 , n1222 , n2034 );
    or g7253 ( n1998 , n14366 , n9643 );
    and g7254 ( n5890 , n13404 , n1787 );
    not g7255 ( n5625 , n4550 );
    nor g7256 ( n2170 , n12651 , n2360 );
    or g7257 ( n11744 , n3164 , n14382 );
    or g7258 ( n1809 , n13991 , n926 );
    and g7259 ( n12843 , n8855 , n11334 );
    and g7260 ( n313 , n4806 , n4048 );
    not g7261 ( n13437 , n4535 );
    and g7262 ( n6455 , n11008 , n7121 );
    or g7263 ( n5390 , n9218 , n4315 );
    or g7264 ( n10266 , n1834 , n4224 );
    nor g7265 ( n2104 , n7365 , n8146 );
    or g7266 ( n13436 , n10394 , n9842 );
    or g7267 ( n13051 , n9289 , n3916 );
    not g7268 ( n12730 , n1813 );
    or g7269 ( n14223 , n2387 , n2273 );
    and g7270 ( n10388 , n10229 , n1864 );
    and g7271 ( n10783 , n9069 , n12618 );
    nor g7272 ( n11770 , n9124 , n3735 );
    or g7273 ( n11150 , n3025 , n12609 );
    or g7274 ( n7307 , n1741 , n4666 );
    not g7275 ( n1383 , n5242 );
    or g7276 ( n9298 , n7462 , n11781 );
    nor g7277 ( n2123 , n10977 , n11056 );
    or g7278 ( n5543 , n2111 , n7716 );
    not g7279 ( n11369 , n9971 );
    or g7280 ( n5789 , n2784 , n3767 );
    and g7281 ( n7599 , n4627 , n14138 );
    nor g7282 ( n12253 , n5024 , n5381 );
    or g7283 ( n3745 , n9211 , n9720 );
    and g7284 ( n7049 , n7081 , n6611 );
    not g7285 ( n12542 , n14501 );
    or g7286 ( n8103 , n12353 , n6281 );
    not g7287 ( n5525 , n1311 );
    and g7288 ( n2175 , n13890 , n9047 );
    not g7289 ( n1681 , n14512 );
    and g7290 ( n5819 , n9811 , n9164 );
    or g7291 ( n12552 , n4481 , n9666 );
    and g7292 ( n7368 , n8431 , n3678 );
    nor g7293 ( n7687 , n11713 , n9094 );
    nor g7294 ( n1283 , n11094 , n7962 );
    and g7295 ( n325 , n10302 , n5263 );
    or g7296 ( n856 , n4045 , n12153 );
    or g7297 ( n6872 , n5491 , n3151 );
    or g7298 ( n9926 , n9230 , n6895 );
    or g7299 ( n13833 , n251 , n213 );
    not g7300 ( n7708 , n6270 );
    or g7301 ( n2358 , n8517 , n2995 );
    or g7302 ( n5133 , n7436 , n3540 );
    or g7303 ( n7724 , n3126 , n7005 );
    or g7304 ( n3342 , n4684 , n9801 );
    not g7305 ( n9766 , n10050 );
    and g7306 ( n8894 , n1428 , n12631 );
    nor g7307 ( n13063 , n7660 , n5128 );
    or g7308 ( n13865 , n10808 , n8993 );
    nor g7309 ( n7601 , n12651 , n4212 );
    or g7310 ( n13808 , n6085 , n9179 );
    and g7311 ( n6408 , n8907 , n11660 );
    or g7312 ( n9389 , n3134 , n2145 );
    or g7313 ( n6734 , n13720 , n3673 );
    or g7314 ( n11561 , n13220 , n3141 );
    not g7315 ( n1784 , n12175 );
    or g7316 ( n3124 , n1838 , n285 );
    and g7317 ( n10473 , n4018 , n5661 );
    and g7318 ( n8642 , n11020 , n3650 );
    nor g7319 ( n3458 , n355 , n14476 );
    and g7320 ( n12810 , n2177 , n14322 );
    or g7321 ( n5160 , n14303 , n7667 );
    or g7322 ( n7849 , n7438 , n11289 );
    and g7323 ( n14111 , n2082 , n5067 );
    or g7324 ( n1048 , n10539 , n2516 );
    nor g7325 ( n2235 , n2790 , n3372 );
    and g7326 ( n1586 , n3672 , n8069 );
    and g7327 ( n6333 , n9972 , n208 );
    and g7328 ( n13490 , n1071 , n10976 );
    not g7329 ( n14238 , n4906 );
    or g7330 ( n10205 , n1051 , n7866 );
    and g7331 ( n11001 , n7798 , n12937 );
    and g7332 ( n9248 , n748 , n12534 );
    and g7333 ( n4139 , n13823 , n13424 );
    and g7334 ( n12195 , n10332 , n13599 );
    and g7335 ( n10210 , n1138 , n4386 );
    or g7336 ( n6108 , n7862 , n3637 );
    and g7337 ( n7379 , n9102 , n9775 );
    not g7338 ( n4821 , n11415 );
    or g7339 ( n2140 , n10234 , n8046 );
    and g7340 ( n4904 , n4844 , n921 );
    nor g7341 ( n12055 , n11713 , n13630 );
    nor g7342 ( n5669 , n742 , n8058 );
    and g7343 ( n10365 , n4261 , n5994 );
    not g7344 ( n12435 , n8799 );
    not g7345 ( n7971 , n2794 );
    and g7346 ( n9067 , n541 , n5415 );
    not g7347 ( n13359 , n13181 );
    and g7348 ( n294 , n8300 , n10393 );
    or g7349 ( n12307 , n9747 , n3116 );
    nor g7350 ( n809 , n8419 , n12785 );
    not g7351 ( n4359 , n4824 );
    or g7352 ( n4170 , n3011 , n8333 );
    or g7353 ( n1657 , n9423 , n10779 );
    and g7354 ( n12442 , n4525 , n13149 );
    and g7355 ( n8164 , n10969 , n8392 );
    and g7356 ( n9302 , n6822 , n463 );
    or g7357 ( n14453 , n2025 , n7461 );
    or g7358 ( n13215 , n11576 , n3052 );
    or g7359 ( n12345 , n12132 , n3166 );
    or g7360 ( n3330 , n13108 , n12065 );
    or g7361 ( n7148 , n7116 , n6317 );
    not g7362 ( n3273 , n12489 );
    or g7363 ( n1589 , n14400 , n13541 );
    or g7364 ( n13834 , n10136 , n3912 );
    not g7365 ( n12934 , n12588 );
    or g7366 ( n14495 , n3527 , n7516 );
    or g7367 ( n9125 , n12549 , n8775 );
    and g7368 ( n8271 , n9069 , n9539 );
    and g7369 ( n7503 , n5918 , n12239 );
    or g7370 ( n14242 , n8964 , n1032 );
    not g7371 ( n227 , n6274 );
    nor g7372 ( n12838 , n3443 , n5941 );
    and g7373 ( n8516 , n11674 , n5352 );
    nor g7374 ( n6677 , n10285 , n10641 );
    and g7375 ( n3806 , n7443 , n7526 );
    and g7376 ( n1364 , n13367 , n3254 );
    and g7377 ( n1518 , n10032 , n7976 );
    or g7378 ( n1217 , n9230 , n11940 );
    or g7379 ( n14202 , n8301 , n11696 );
    not g7380 ( n5268 , n11375 );
    not g7381 ( n13854 , n4891 );
    and g7382 ( n12493 , n5240 , n9926 );
    not g7383 ( n5951 , n2371 );
    or g7384 ( n8314 , n3099 , n3481 );
    and g7385 ( n14010 , n7693 , n13137 );
    not g7386 ( n11444 , n5217 );
    or g7387 ( n12464 , n2025 , n10899 );
    or g7388 ( n7300 , n48 , n9869 );
    or g7389 ( n13282 , n3800 , n13837 );
    or g7390 ( n4070 , n12295 , n8853 );
    or g7391 ( n6035 , n12149 , n7387 );
    and g7392 ( n12710 , n9198 , n4800 );
    and g7393 ( n13922 , n392 , n9212 );
    not g7394 ( n2857 , n10346 );
    and g7395 ( n14071 , n1011 , n9658 );
    or g7396 ( n6789 , n6111 , n5862 );
    and g7397 ( n126 , n4022 , n2664 );
    nor g7398 ( n1615 , n228 , n14228 );
    and g7399 ( n1154 , n392 , n216 );
    and g7400 ( n6235 , n5053 , n13088 );
    and g7401 ( n2806 , n11569 , n12839 );
    and g7402 ( n2796 , n4422 , n9331 );
    not g7403 ( n13877 , n7120 );
    and g7404 ( n10557 , n2961 , n12017 );
    or g7405 ( n11204 , n10857 , n8123 );
    nor g7406 ( n7783 , n5833 , n10001 );
    and g7407 ( n5030 , n9724 , n12337 );
    and g7408 ( n13696 , n9829 , n5148 );
    and g7409 ( n643 , n1193 , n13515 );
    not g7410 ( n12475 , n1571 );
    not g7411 ( n1920 , n9110 );
    or g7412 ( n13588 , n6695 , n13179 );
    or g7413 ( n3160 , n7462 , n290 );
    and g7414 ( n12438 , n12259 , n11807 );
    or g7415 ( n1593 , n13083 , n653 );
    and g7416 ( n1124 , n271 , n9765 );
    or g7417 ( n11831 , n387 , n11599 );
    or g7418 ( n7611 , n185 , n2324 );
    not g7419 ( n11636 , n13219 );
    and g7420 ( n27 , n12421 , n4770 );
    and g7421 ( n7674 , n1699 , n13032 );
    or g7422 ( n6208 , n1028 , n106 );
    or g7423 ( n8834 , n9864 , n5792 );
    or g7424 ( n13424 , n3168 , n9028 );
    and g7425 ( n12231 , n7057 , n14371 );
    or g7426 ( n6628 , n8581 , n5080 );
    and g7427 ( n2876 , n7779 , n7932 );
    or g7428 ( n12291 , n4684 , n14381 );
    or g7429 ( n13281 , n3120 , n12369 );
    or g7430 ( n11437 , n4739 , n4938 );
    not g7431 ( n7462 , n1060 );
    nor g7432 ( n9328 , n4741 , n1012 );
    nor g7433 ( n3920 , n10511 , n12283 );
    nor g7434 ( n4738 , n7223 , n3909 );
    and g7435 ( n10430 , n3715 , n8040 );
    or g7436 ( n3454 , n12139 , n3828 );
    and g7437 ( n539 , n7957 , n806 );
    or g7438 ( n8772 , n11710 , n9049 );
    or g7439 ( n1377 , n4320 , n11666 );
    nor g7440 ( n13070 , n1722 , n3639 );
    and g7441 ( n2261 , n4244 , n273 );
    and g7442 ( n9369 , n3861 , n1596 );
    or g7443 ( n862 , n4045 , n7451 );
    not g7444 ( n13489 , n4490 );
    or g7445 ( n13284 , n13142 , n11823 );
    and g7446 ( n12833 , n7267 , n13136 );
    or g7447 ( n2838 , n4255 , n9911 );
    not g7448 ( n4633 , n1544 );
    and g7449 ( n7349 , n8849 , n5514 );
    and g7450 ( n12834 , n2322 , n3071 );
    nor g7451 ( n9521 , n1769 , n86 );
    or g7452 ( n1645 , n13432 , n2659 );
    and g7453 ( n2361 , n3212 , n1817 );
    and g7454 ( n574 , n10399 , n4526 );
    nor g7455 ( n3816 , n11771 , n11275 );
    or g7456 ( n3316 , n7250 , n5737 );
    not g7457 ( n11674 , n6829 );
    or g7458 ( n11690 , n10713 , n1558 );
    or g7459 ( n5971 , n9780 , n2828 );
    and g7460 ( n2182 , n10855 , n4834 );
    and g7461 ( n7335 , n3405 , n3160 );
    not g7462 ( n6857 , n4720 );
    or g7463 ( n10439 , n11459 , n9510 );
    and g7464 ( n9662 , n10854 , n529 );
    and g7465 ( n835 , n9315 , n11806 );
    or g7466 ( n5220 , n1261 , n4567 );
    and g7467 ( n12787 , n12721 , n3827 );
    not g7468 ( n3457 , n7546 );
    or g7469 ( n10645 , n2181 , n13057 );
    not g7470 ( n1452 , n1843 );
    and g7471 ( n551 , n5240 , n5337 );
    and g7472 ( n6342 , n7911 , n9258 );
    or g7473 ( n5717 , n2057 , n13950 );
    not g7474 ( n12480 , n13364 );
    or g7475 ( n8783 , n1202 , n1736 );
    and g7476 ( n4721 , n1804 , n2980 );
    or g7477 ( n7665 , n695 , n1465 );
    and g7478 ( n2633 , n12935 , n1068 );
    and g7479 ( n8632 , n12592 , n5056 );
    and g7480 ( n232 , n5252 , n2430 );
    or g7481 ( n5305 , n7227 , n3999 );
    or g7482 ( n2867 , n6971 , n4470 );
    or g7483 ( n9782 , n11223 , n4952 );
    nor g7484 ( n6840 , n11580 , n7625 );
    or g7485 ( n10561 , n1258 , n2220 );
    and g7486 ( n3328 , n14388 , n2469 );
    and g7487 ( n10581 , n6316 , n3985 );
    and g7488 ( n3666 , n8020 , n5896 );
    or g7489 ( n13896 , n7430 , n7664 );
    not g7490 ( n919 , n8814 );
    and g7491 ( n2975 , n638 , n5699 );
    and g7492 ( n5388 , n13572 , n12996 );
    not g7493 ( n13361 , n7376 );
    and g7494 ( n13144 , n9113 , n12997 );
    not g7495 ( n5335 , n8963 );
    or g7496 ( n2450 , n2412 , n6733 );
    not g7497 ( n6311 , n5427 );
    and g7498 ( n5942 , n10678 , n11549 );
    nor g7499 ( n3148 , n10650 , n7567 );
    nor g7500 ( n1050 , n11259 , n4344 );
    nor g7501 ( n12433 , n4092 , n3971 );
    and g7502 ( n2722 , n10562 , n1645 );
    and g7503 ( n9527 , n5071 , n12849 );
    and g7504 ( n2701 , n12259 , n13410 );
    and g7505 ( n1543 , n986 , n12064 );
    not g7506 ( n3276 , n11668 );
    not g7507 ( n8821 , n622 );
    or g7508 ( n3701 , n9747 , n11736 );
    and g7509 ( n11382 , n1231 , n10009 );
    and g7510 ( n7311 , n8432 , n4241 );
    or g7511 ( n14127 , n5587 , n226 );
    and g7512 ( n14447 , n7529 , n13665 );
    or g7513 ( n1796 , n5997 , n13638 );
    or g7514 ( n370 , n4840 , n8371 );
    and g7515 ( n8246 , n904 , n6294 );
    or g7516 ( n8355 , n172 , n9902 );
    or g7517 ( n1248 , n1538 , n13289 );
    not g7518 ( n5317 , n7346 );
    not g7519 ( n2645 , n426 );
    and g7520 ( n1170 , n8147 , n9367 );
    not g7521 ( n13869 , n394 );
    and g7522 ( n8531 , n12592 , n2203 );
    and g7523 ( n1162 , n10209 , n7423 );
    or g7524 ( n13374 , n3025 , n11115 );
    and g7525 ( n13668 , n2967 , n12924 );
    nor g7526 ( n13596 , n9557 , n1953 );
    and g7527 ( n2028 , n6486 , n13801 );
    and g7528 ( n5983 , n4359 , n13451 );
    and g7529 ( n5224 , n5471 , n3330 );
    and g7530 ( n13241 , n8047 , n12653 );
    nor g7531 ( n7625 , n11988 , n4108 );
    or g7532 ( n6621 , n3219 , n10833 );
    and g7533 ( n6465 , n873 , n83 );
    and g7534 ( n8056 , n10763 , n284 );
    and g7535 ( n7640 , n103 , n11294 );
    or g7536 ( n7615 , n10534 , n2500 );
    and g7537 ( n6636 , n13863 , n7133 );
    not g7538 ( n12615 , n6193 );
    or g7539 ( n9756 , n10024 , n5578 );
    and g7540 ( n5169 , n11008 , n14090 );
    not g7541 ( n8250 , n230 );
    or g7542 ( n6811 , n14449 , n4948 );
    and g7543 ( n8754 , n6128 , n13482 );
    and g7544 ( n3374 , n1772 , n4106 );
    or g7545 ( n1156 , n6781 , n8823 );
    not g7546 ( n2432 , n10861 );
    nor g7547 ( n1274 , n4050 , n956 );
    or g7548 ( n614 , n11647 , n7411 );
    or g7549 ( n11601 , n10784 , n3289 );
    nor g7550 ( n5805 , n12075 , n2209 );
    and g7551 ( n686 , n12730 , n10551 );
    and g7552 ( n4271 , n3536 , n10139 );
    and g7553 ( n8519 , n7063 , n11346 );
    nor g7554 ( n10843 , n1860 , n7204 );
    or g7555 ( n14030 , n3527 , n1082 );
    and g7556 ( n1024 , n12421 , n10170 );
    and g7557 ( n2551 , n9315 , n11307 );
    not g7558 ( n6041 , n13779 );
    not g7559 ( n9232 , n10269 );
    and g7560 ( n1531 , n1610 , n14315 );
    or g7561 ( n12262 , n14435 , n4129 );
    or g7562 ( n4799 , n7527 , n4979 );
    or g7563 ( n6651 , n13847 , n14180 );
    and g7564 ( n8305 , n12250 , n5671 );
    and g7565 ( n13504 , n1125 , n1863 );
    nor g7566 ( n11538 , n5159 , n11657 );
    or g7567 ( n5327 , n11551 , n6592 );
    or g7568 ( n775 , n5507 , n10696 );
    and g7569 ( n12784 , n3813 , n190 );
    or g7570 ( n4992 , n3088 , n10337 );
    nor g7571 ( n6269 , n1681 , n6133 );
    not g7572 ( n13283 , n1073 );
    and g7573 ( n5440 , n12472 , n14053 );
    or g7574 ( n7656 , n5986 , n10306 );
    or g7575 ( n4605 , n7914 , n4736 );
    or g7576 ( n14298 , n12034 , n14010 );
    or g7577 ( n8658 , n8816 , n12313 );
    or g7578 ( n11633 , n13186 , n8439 );
    and g7579 ( n3468 , n10457 , n12085 );
    not g7580 ( n10342 , n2607 );
    and g7581 ( n774 , n11163 , n1470 );
    and g7582 ( n11255 , n3586 , n1330 );
    nor g7583 ( n2880 , n10289 , n6702 );
    or g7584 ( n7425 , n10913 , n551 );
    or g7585 ( n2731 , n3652 , n3799 );
    and g7586 ( n6737 , n12998 , n13344 );
    nor g7587 ( n11681 , n1685 , n10885 );
    and g7588 ( n7647 , n8147 , n12814 );
    and g7589 ( n3680 , n5948 , n8744 );
    or g7590 ( n12732 , n11647 , n5028 );
    or g7591 ( n7045 , n3062 , n64 );
    or g7592 ( n12496 , n9174 , n6367 );
    nor g7593 ( n5784 , n12191 , n4463 );
    or g7594 ( n9001 , n85 , n5820 );
    and g7595 ( n6895 , n9617 , n8760 );
    not g7596 ( n678 , n11969 );
    not g7597 ( n1458 , n14181 );
    or g7598 ( n6871 , n13941 , n3966 );
    or g7599 ( n8792 , n11472 , n3753 );
    or g7600 ( n11103 , n251 , n12843 );
    or g7601 ( n2817 , n11581 , n14117 );
    or g7602 ( n1957 , n6350 , n8205 );
    or g7603 ( n12136 , n4172 , n74 );
    and g7604 ( n11534 , n6436 , n8298 );
    and g7605 ( n8625 , n5948 , n5021 );
    nor g7606 ( n11772 , n13979 , n7207 );
    or g7607 ( n11638 , n4052 , n654 );
    or g7608 ( n13746 , n7358 , n4027 );
    and g7609 ( n10292 , n3286 , n1635 );
    or g7610 ( n5171 , n8450 , n10378 );
    or g7611 ( n307 , n4065 , n3732 );
    or g7612 ( n5157 , n7678 , n12405 );
    or g7613 ( n11692 , n4631 , n2586 );
    and g7614 ( n11513 , n1937 , n5770 );
    or g7615 ( n1477 , n4828 , n7986 );
    not g7616 ( n13981 , n4500 );
    and g7617 ( n4397 , n5071 , n3664 );
    not g7618 ( n3043 , n5023 );
    not g7619 ( n79 , n5795 );
    and g7620 ( n8092 , n10229 , n3761 );
    and g7621 ( n12646 , n2682 , n4097 );
    or g7622 ( n12538 , n12019 , n5165 );
    not g7623 ( n10864 , n2752 );
    and g7624 ( n10632 , n14042 , n113 );
    nor g7625 ( n708 , n7900 , n11267 );
    and g7626 ( n14412 , n2951 , n10403 );
    not g7627 ( n3424 , n6193 );
    not g7628 ( n3356 , n5761 );
    or g7629 ( n10411 , n9529 , n7100 );
    and g7630 ( n4548 , n7284 , n440 );
    or g7631 ( n11759 , n6654 , n4251 );
    or g7632 ( n10773 , n13698 , n13006 );
    or g7633 ( n4512 , n9507 , n5913 );
    and g7634 ( n10644 , n9890 , n12951 );
    and g7635 ( n7231 , n3986 , n4070 );
    and g7636 ( n12963 , n8250 , n175 );
    or g7637 ( n9350 , n7230 , n702 );
    and g7638 ( n157 , n6318 , n9491 );
    and g7639 ( n13073 , n3405 , n846 );
    and g7640 ( n1942 , n6343 , n9678 );
    or g7641 ( n5484 , n6848 , n12782 );
    and g7642 ( n3576 , n7203 , n13550 );
    and g7643 ( n9548 , n5317 , n2335 );
    nor g7644 ( n3475 , n1357 , n7184 );
    or g7645 ( n7574 , n8517 , n10581 );
    or g7646 ( n13429 , n3673 , n5023 );
    and g7647 ( n10403 , n10953 , n5226 );
    or g7648 ( n7215 , n8581 , n5814 );
    or g7649 ( n8830 , n974 , n1754 );
    and g7650 ( n8182 , n7187 , n11323 );
    and g7651 ( n1453 , n13626 , n13838 );
    nor g7652 ( n12979 , n3107 , n7234 );
    or g7653 ( n4680 , n6519 , n10665 );
    or g7654 ( n11326 , n11047 , n3004 );
    not g7655 ( n1480 , n5627 );
    not g7656 ( n2310 , n8008 );
    or g7657 ( n13699 , n5483 , n9064 );
    or g7658 ( n434 , n9490 , n9914 );
    not g7659 ( n6053 , n10254 );
    or g7660 ( n12696 , n8242 , n7288 );
    nor g7661 ( n10106 , n2236 , n13358 );
    not g7662 ( n4906 , n11628 );
    and g7663 ( n1142 , n13342 , n3998 );
    or g7664 ( n3656 , n14481 , n6505 );
    and g7665 ( n7326 , n4722 , n7688 );
    or g7666 ( n9602 , n12625 , n6735 );
    not g7667 ( n11581 , n11055 );
    and g7668 ( n4551 , n8569 , n3593 );
    or g7669 ( n4514 , n8748 , n3611 );
    not g7670 ( n2904 , n1495 );
    and g7671 ( n8307 , n11636 , n6190 );
    not g7672 ( n1225 , n10283 );
    or g7673 ( n8951 , n5362 , n2637 );
    nor g7674 ( n6324 , n6397 , n1519 );
    and g7675 ( n9526 , n11838 , n2114 );
    and g7676 ( n7288 , n11153 , n14443 );
    or g7677 ( n1863 , n11090 , n5534 );
    or g7678 ( n121 , n6519 , n880 );
    or g7679 ( n12228 , n10024 , n8098 );
    or g7680 ( n9738 , n2760 , n13509 );
    not g7681 ( n9803 , n7450 );
    and g7682 ( n11169 , n2058 , n625 );
    not g7683 ( n12226 , n6139 );
    not g7684 ( n12705 , n12691 );
    and g7685 ( n14125 , n3932 , n3241 );
    and g7686 ( n9443 , n5053 , n7646 );
    or g7687 ( n1569 , n1172 , n3567 );
    and g7688 ( n13911 , n8786 , n12954 );
    not g7689 ( n6013 , n9950 );
    or g7690 ( n11777 , n12400 , n4451 );
    and g7691 ( n3153 , n7284 , n4798 );
    or g7692 ( n13949 , n7803 , n14294 );
    nor g7693 ( n2899 , n13627 , n709 );
    or g7694 ( n3578 , n14282 , n7750 );
    not g7695 ( n9353 , n9169 );
    or g7696 ( n5087 , n3273 , n12787 );
    or g7697 ( n5063 , n8045 , n9548 );
    not g7698 ( n9113 , n5268 );
    and g7699 ( n4763 , n7708 , n1755 );
    nor g7700 ( n5069 , n5132 , n8101 );
    and g7701 ( n10498 , n706 , n10706 );
    not g7702 ( n9174 , n6332 );
    or g7703 ( n12322 , n10407 , n4659 );
    not g7704 ( n8386 , n9197 );
    or g7705 ( n7292 , n8581 , n3911 );
    not g7706 ( n14166 , n12687 );
    and g7707 ( n7302 , n706 , n10690 );
    nor g7708 ( n1390 , n12112 , n7985 );
    and g7709 ( n4939 , n9516 , n7336 );
    and g7710 ( n1773 , n4757 , n8095 );
    and g7711 ( n12563 , n6130 , n13100 );
    not g7712 ( n7219 , n6357 );
    or g7713 ( n1306 , n14419 , n12824 );
    or g7714 ( n6916 , n8332 , n105 );
    and g7715 ( n6225 , n7391 , n2708 );
    or g7716 ( n5238 , n11036 , n12003 );
    not g7717 ( n717 , n8291 );
    and g7718 ( n14267 , n5475 , n2773 );
    nor g7719 ( n5323 , n13072 , n9033 );
    not g7720 ( n200 , n8048 );
    and g7721 ( n10869 , n2521 , n6792 );
    and g7722 ( n14407 , n3028 , n6042 );
    or g7723 ( n5044 , n5800 , n13545 );
    and g7724 ( n13391 , n1962 , n10476 );
    and g7725 ( n1456 , n11803 , n12578 );
    and g7726 ( n2438 , n7529 , n8173 );
    or g7727 ( n8118 , n838 , n12921 );
    or g7728 ( n11218 , n11479 , n8463 );
    not g7729 ( n4417 , n93 );
    and g7730 ( n6482 , n7934 , n3929 );
    and g7731 ( n9251 , n646 , n5659 );
    or g7732 ( n11351 , n8821 , n12006 );
    not g7733 ( n6099 , n4656 );
    not g7734 ( n12994 , n1220 );
    nor g7735 ( n12758 , n10189 , n5299 );
    or g7736 ( n10155 , n11980 , n2574 );
    and g7737 ( n3731 , n6318 , n11955 );
    not g7738 ( n1278 , n4785 );
    and g7739 ( n7257 , n4722 , n2652 );
    and g7740 ( n9347 , n8111 , n8807 );
    nor g7741 ( n3235 , n1112 , n2579 );
    nor g7742 ( n12194 , n946 , n12940 );
    and g7743 ( n9842 , n3536 , n9935 );
    or g7744 ( n847 , n7481 , n2997 );
    or g7745 ( n12340 , n14107 , n5581 );
    or g7746 ( n9202 , n10523 , n1580 );
    not g7747 ( n1100 , n6326 );
    and g7748 ( n14441 , n638 , n10297 );
    and g7749 ( n11586 , n10622 , n6183 );
    nor g7750 ( n3997 , n7720 , n11353 );
    not g7751 ( n5675 , n13560 );
    and g7752 ( n11616 , n7015 , n11846 );
    or g7753 ( n5470 , n13547 , n6235 );
    nor g7754 ( n10200 , n13350 , n1472 );
    and g7755 ( n6336 , n8605 , n8560 );
    or g7756 ( n8040 , n7219 , n351 );
    or g7757 ( n14024 , n6989 , n30 );
    and g7758 ( n13164 , n1937 , n6576 );
    not g7759 ( n5459 , n10828 );
    nor g7760 ( n11418 , n8607 , n1056 );
    and g7761 ( n5115 , n10134 , n13217 );
    and g7762 ( n11136 , n13535 , n1973 );
    or g7763 ( n5103 , n6595 , n3796 );
    and g7764 ( n1437 , n7691 , n5487 );
    nor g7765 ( n6199 , n5480 , n2512 );
    and g7766 ( n4121 , n5779 , n1130 );
    nor g7767 ( n3735 , n48 , n11486 );
    and g7768 ( n6739 , n14063 , n14439 );
    and g7769 ( n12208 , n11093 , n5813 );
    and g7770 ( n680 , n3846 , n4863 );
    not g7771 ( n13038 , n6308 );
    and g7772 ( n1906 , n13252 , n8394 );
    and g7773 ( n9573 , n2527 , n14424 );
    not g7774 ( n2822 , n481 );
    not g7775 ( n12243 , n2009 );
    and g7776 ( n5736 , n9102 , n5039 );
    or g7777 ( n7820 , n85 , n12027 );
    and g7778 ( n13441 , n10815 , n8192 );
    and g7779 ( n5282 , n9890 , n2614 );
    or g7780 ( n891 , n13706 , n8109 );
    or g7781 ( n10575 , n3219 , n1454 );
    and g7782 ( n7964 , n7421 , n7356 );
    or g7783 ( n13095 , n769 , n4794 );
    and g7784 ( n7895 , n12445 , n10037 );
    and g7785 ( n2328 , n13240 , n12199 );
    and g7786 ( n9619 , n2367 , n1188 );
    or g7787 ( n9462 , n7249 , n3059 );
    not g7788 ( n7130 , n8446 );
    or g7789 ( n303 , n4365 , n7652 );
    nor g7790 ( n5849 , n9529 , n5741 );
    and g7791 ( n1129 , n12013 , n12419 );
    or g7792 ( n12861 , n2645 , n9534 );
    or g7793 ( n11026 , n11951 , n6366 );
    and g7794 ( n10818 , n13525 , n11075 );
    not g7795 ( n1391 , n9686 );
    and g7796 ( n14018 , n8247 , n11895 );
    not g7797 ( n700 , n201 );
    and g7798 ( n13702 , n8427 , n1276 );
    or g7799 ( n383 , n3826 , n7089 );
    or g7800 ( n6181 , n1061 , n5292 );
    or g7801 ( n6102 , n9211 , n3486 );
    and g7802 ( n4186 , n541 , n12246 );
    not g7803 ( n2781 , n6670 );
    or g7804 ( n12692 , n5569 , n11709 );
    and g7805 ( n4734 , n4289 , n6628 );
    and g7806 ( n11292 , n9052 , n332 );
    nor g7807 ( n12286 , n2017 , n237 );
    or g7808 ( n922 , n7700 , n12583 );
    nor g7809 ( n7894 , n4639 , n7355 );
    or g7810 ( n6021 , n7116 , n14432 );
    or g7811 ( n11773 , n10449 , n1016 );
    and g7812 ( n13914 , n4445 , n4068 );
    nor g7813 ( n3239 , n3255 , n7608 );
    or g7814 ( n12361 , n12695 , n11395 );
    or g7815 ( n11892 , n8332 , n8030 );
    not g7816 ( n7275 , n13765 );
    nor g7817 ( n11079 , n14058 , n322 );
    nor g7818 ( n1758 , n12334 , n9007 );
    not g7819 ( n12211 , n1220 );
    or g7820 ( n9533 , n11804 , n7025 );
    and g7821 ( n10088 , n5475 , n7307 );
    and g7822 ( n12959 , n12592 , n6530 );
    or g7823 ( n9160 , n6690 , n33 );
    nor g7824 ( n5748 , n9807 , n7136 );
    or g7825 ( n4293 , n7076 , n148 );
    or g7826 ( n8456 , n4822 , n8995 );
    or g7827 ( n10237 , n10089 , n11005 );
    and g7828 ( n2883 , n2521 , n11083 );
    not g7829 ( n10332 , n168 );
    not g7830 ( n13781 , n12970 );
    and g7831 ( n9946 , n1452 , n9363 );
    and g7832 ( n2004 , n12960 , n4378 );
    and g7833 ( n786 , n1937 , n649 );
    and g7834 ( n6470 , n7208 , n9797 );
    or g7835 ( n7966 , n3273 , n13122 );
    or g7836 ( n7193 , n6206 , n10206 );
    and g7837 ( n6201 , n12185 , n12458 );
    and g7838 ( n8070 , n2422 , n9518 );
    or g7839 ( n4716 , n6388 , n1568 );
    and g7840 ( n9447 , n12782 , n9276 );
    and g7841 ( n2308 , n9315 , n10716 );
    and g7842 ( n5130 , n9972 , n12464 );
    and g7843 ( n2060 , n4655 , n10533 );
    or g7844 ( n6580 , n11231 , n12877 );
    not g7845 ( n4791 , n12489 );
    and g7846 ( n9180 , n13421 , n4801 );
    or g7847 ( n345 , n13501 , n3020 );
    and g7848 ( n9642 , n3710 , n7033 );
    or g7849 ( n867 , n5144 , n3006 );
    or g7850 ( n13417 , n6672 , n7542 );
    and g7851 ( n7750 , n4422 , n1184 );
    and g7852 ( n8253 , n898 , n12783 );
    or g7853 ( n14056 , n172 , n3200 );
    and g7854 ( n2671 , n2021 , n14025 );
    and g7855 ( n11943 , n7909 , n10454 );
    nor g7856 ( n1694 , n5035 , n2028 );
    and g7857 ( n8937 , n1904 , n13341 );
    or g7858 ( n5838 , n12625 , n2458 );
    or g7859 ( n2226 , n3043 , n4225 );
    or g7860 ( n10998 , n1011 , n8800 );
    or g7861 ( n50 , n7219 , n10547 );
    and g7862 ( n12044 , n6606 , n29 );
    and g7863 ( n11364 , n5489 , n4119 );
    not g7864 ( n10245 , n3007 );
    or g7865 ( n139 , n6519 , n7738 );
    nor g7866 ( n6228 , n900 , n2314 );
    and g7867 ( n3199 , n8866 , n5576 );
    or g7868 ( n5304 , n5483 , n5161 );
    or g7869 ( n10770 , n11223 , n14234 );
    and g7870 ( n13570 , n7370 , n5309 );
    and g7871 ( n14299 , n6135 , n9162 );
    or g7872 ( n1367 , n838 , n2440 );
    not g7873 ( n8363 , n5690 );
    or g7874 ( n12889 , n13501 , n14272 );
    and g7875 ( n14275 , n5582 , n6154 );
    nor g7876 ( n11964 , n9078 , n12979 );
    not g7877 ( n2694 , n628 );
    not g7878 ( n8557 , n9214 );
    or g7879 ( n8196 , n8701 , n4959 );
    nor g7880 ( n13278 , n2575 , n1233 );
    not g7881 ( n4340 , n918 );
    or g7882 ( n5832 , n1278 , n730 );
    and g7883 ( n6929 , n4358 , n2821 );
    not g7884 ( n3967 , n5886 );
    not g7885 ( n10511 , n7291 );
    and g7886 ( n11865 , n6507 , n9964 );
    not g7887 ( n7779 , n2619 );
    or g7888 ( n9420 , n8592 , n11770 );
    not g7889 ( n5944 , n1979 );
    nor g7890 ( n8146 , n1623 , n1852 );
    and g7891 ( n4132 , n12185 , n4285 );
    or g7892 ( n7874 , n10154 , n12607 );
    or g7893 ( n76 , n4045 , n14021 );
    or g7894 ( n5928 , n8964 , n6095 );
    and g7895 ( n10483 , n7308 , n10518 );
    not g7896 ( n3196 , n4711 );
    or g7897 ( n2570 , n11620 , n3810 );
    not g7898 ( n11445 , n12189 );
    not g7899 ( n168 , n3331 );
    or g7900 ( n1290 , n5084 , n3580 );
    or g7901 ( n10017 , n3273 , n6180 );
    and g7902 ( n12507 , n7429 , n11372 );
    nor g7903 ( n3436 , n2086 , n302 );
    or g7904 ( n9594 , n3914 , n5657 );
    or g7905 ( n3902 , n8638 , n2650 );
    and g7906 ( n11925 , n5348 , n3187 );
    and g7907 ( n1146 , n2961 , n2702 );
    or g7908 ( n9540 , n8378 , n849 );
    or g7909 ( n11138 , n14481 , n1081 );
    or g7910 ( n2759 , n573 , n13448 );
    and g7911 ( n137 , n3724 , n8616 );
    or g7912 ( n12410 , n555 , n1148 );
    and g7913 ( n1476 , n8801 , n545 );
    nor g7914 ( n14341 , n5217 , n459 );
    and g7915 ( n2389 , n8769 , n470 );
    or g7916 ( n10307 , n1855 , n11404 );
    or g7917 ( n11878 , n3193 , n7789 );
    or g7918 ( n12491 , n7359 , n4376 );
    or g7919 ( n7194 , n5007 , n14146 );
    and g7920 ( n1224 , n3846 , n6143 );
    and g7921 ( n1235 , n8932 , n1281 );
    and g7922 ( n4223 , n4095 , n5868 );
    not g7923 ( n10637 , n10775 );
    or g7924 ( n2433 , n13226 , n4647 );
    and g7925 ( n2859 , n8412 , n9175 );
    and g7926 ( n1310 , n12531 , n13612 );
    or g7927 ( n2553 , n12401 , n6303 );
    or g7928 ( n3554 , n8210 , n6772 );
    nor g7929 ( n1344 , n2781 , n3924 );
    and g7930 ( n2853 , n5252 , n12290 );
    and g7931 ( n7248 , n12226 , n3337 );
    or g7932 ( n5189 , n4481 , n12806 );
    nor g7933 ( n10963 , n619 , n6419 );
    or g7934 ( n10844 , n14419 , n5821 );
    or g7935 ( n13787 , n2686 , n5000 );
    and g7936 ( n2504 , n10854 , n21 );
    and g7937 ( n10813 , n9811 , n5451 );
    or g7938 ( n6120 , n8034 , n14247 );
    or g7939 ( n7824 , n3168 , n5517 );
    and g7940 ( n1592 , n2709 , n4981 );
    nor g7941 ( n4671 , n10712 , n3231 );
    not g7942 ( n11123 , n7875 );
    or g7943 ( n14161 , n4840 , n3841 );
    nor g7944 ( n2317 , n3696 , n5645 );
    or g7945 ( n3484 , n3777 , n14179 );
    and g7946 ( n8137 , n4509 , n14398 );
    nor g7947 ( n10425 , n13276 , n1103 );
    and g7948 ( n12359 , n9890 , n2153 );
    or g7949 ( n14251 , n6090 , n8169 );
    or g7950 ( n1206 , n5997 , n2884 );
    or g7951 ( n594 , n13112 , n10279 );
    not g7952 ( n1423 , n12714 );
    or g7953 ( n3869 , n12169 , n3921 );
    and g7954 ( n10806 , n8932 , n3858 );
    or g7955 ( n4048 , n3886 , n2108 );
    and g7956 ( n7128 , n5137 , n9511 );
    or g7957 ( n11312 , n6629 , n10386 );
    and g7958 ( n10810 , n2330 , n13282 );
    and g7959 ( n11338 , n4289 , n2937 );
    not g7960 ( n4601 , n14408 );
    nor g7961 ( n9840 , n3845 , n8648 );
    or g7962 ( n3254 , n8378 , n4262 );
    or g7963 ( n14443 , n12695 , n2639 );
    or g7964 ( n12091 , n11519 , n10225 );
    and g7965 ( n11460 , n6527 , n1387 );
    or g7966 ( n4285 , n12211 , n9559 );
    not g7967 ( n10626 , n13234 );
    nor g7968 ( n14333 , n13477 , n5864 );
    and g7969 ( n12203 , n5999 , n5066 );
    and g7970 ( n3198 , n2846 , n308 );
    and g7971 ( n13456 , n3743 , n12873 );
    not g7972 ( n3126 , n4939 );
    nor g7973 ( n14228 , n4270 , n11727 );
    or g7974 ( n4946 , n7812 , n14378 );
    or g7975 ( n7138 , n930 , n9932 );
    or g7976 ( n2835 , n1006 , n7827 );
    or g7977 ( n12913 , n2761 , n3143 );
    nor g7978 ( n12513 , n8361 , n12005 );
    nor g7979 ( n9115 , n10936 , n8057 );
    nor g7980 ( n6572 , n6672 , n5243 );
    or g7981 ( n576 , n9442 , n1224 );
    and g7982 ( n14123 , n4690 , n8870 );
    or g7983 ( n2309 , n13754 , n2165 );
    not g7984 ( n8404 , n918 );
    and g7985 ( n11308 , n1932 , n5265 );
    not g7986 ( n11597 , n9465 );
    nor g7987 ( n5703 , n5977 , n2739 );
    or g7988 ( n10356 , n5807 , n9584 );
    and g7989 ( n5892 , n3861 , n800 );
    and g7990 ( n8176 , n6013 , n10992 );
    or g7991 ( n8053 , n5977 , n2764 );
    and g7992 ( n2825 , n9650 , n13747 );
    or g7993 ( n13521 , n6271 , n13242 );
    and g7994 ( n1398 , n10622 , n9660 );
    nor g7995 ( n3305 , n13557 , n10373 );
    or g7996 ( n7594 , n11724 , n4165 );
    not g7997 ( n8301 , n4939 );
    and g7998 ( n2333 , n14213 , n1542 );
    nor g7999 ( n10464 , n1820 , n10793 );
    and g8000 ( n2284 , n14358 , n7029 );
    or g8001 ( n5002 , n13518 , n10471 );
    not g8002 ( n13912 , n6517 );
    and g8003 ( n3601 , n2378 , n3067 );
    and g8004 ( n7361 , n3923 , n11866 );
    and g8005 ( n7769 , n10763 , n14127 );
    and g8006 ( n7165 , n11406 , n5096 );
    or g8007 ( n1849 , n5454 , n6066 );
    or g8008 ( n8744 , n5144 , n6207 );
    and g8009 ( n9812 , n9102 , n3508 );
    and g8010 ( n9407 , n286 , n12595 );
    not g8011 ( n930 , n3455 );
    and g8012 ( n3291 , n7779 , n13275 );
    or g8013 ( n13919 , n7430 , n719 );
    and g8014 ( n9790 , n1526 , n13094 );
    and g8015 ( n2778 , n8620 , n4975 );
    and g8016 ( n13775 , n3286 , n11769 );
    or g8017 ( n5415 , n1383 , n12901 );
    and g8018 ( n1918 , n12092 , n11077 );
    or g8019 ( n4373 , n9792 , n13992 );
    or g8020 ( n14046 , n3088 , n6826 );
    or g8021 ( n794 , n5570 , n2479 );
    and g8022 ( n8001 , n2643 , n1811 );
    or g8023 ( n7495 , n4791 , n11089 );
    and g8024 ( n10038 , n5088 , n9384 );
    or g8025 ( n1443 , n8908 , n114 );
    and g8026 ( n3406 , n11484 , n8718 );
    or g8027 ( n1484 , n10534 , n5973 );
    and g8028 ( n3082 , n13755 , n14152 );
    not g8029 ( n8581 , n6274 );
    and g8030 ( n6229 , n2564 , n3674 );
    and g8031 ( n9524 , n12472 , n7301 );
    not g8032 ( n10330 , n7802 );
    or g8033 ( n5993 , n8638 , n6346 );
    and g8034 ( n4700 , n6854 , n4100 );
    not g8035 ( n8332 , n4317 );
    or g8036 ( n660 , n2179 , n12287 );
    and g8037 ( n5546 , n5471 , n6017 );
    and g8038 ( n1220 , n10012 , n887 );
    and g8039 ( n784 , n2983 , n4946 );
    not g8040 ( n7767 , n7920 );
    or g8041 ( n9148 , n11405 , n4329 );
    or g8042 ( n3761 , n11105 , n274 );
    or g8043 ( n10716 , n11048 , n7847 );
    and g8044 ( n9326 , n12105 , n13374 );
    and g8045 ( n8328 , n5071 , n14192 );
    or g8046 ( n10339 , n476 , n13542 );
    not g8047 ( n10560 , n12588 );
    or g8048 ( n14014 , n5253 , n5501 );
    and g8049 ( n9138 , n4365 , n9270 );
    or g8050 ( n12372 , n13991 , n4989 );
    and g8051 ( n8566 , n13404 , n7226 );
    or g8052 ( n569 , n1044 , n6483 );
    or g8053 ( n7848 , n1576 , n5653 );
    nor g8054 ( n8352 , n14058 , n14434 );
    and g8055 ( n4442 , n8950 , n1512 );
    or g8056 ( n872 , n12500 , n6255 );
    or g8057 ( n1348 , n2201 , n6147 );
    or g8058 ( n616 , n4180 , n1688 );
    nor g8059 ( n2163 , n4771 , n9838 );
    and g8060 ( n14479 , n1414 , n7790 );
    and g8061 ( n6582 , n10399 , n5123 );
    or g8062 ( n9085 , n8458 , n2482 );
    not g8063 ( n974 , n6978 );
    nor g8064 ( n8459 , n7683 , n6195 );
    not g8065 ( n13867 , n11666 );
    and g8066 ( n11333 , n4289 , n4644 );
    nor g8067 ( n6667 , n4417 , n4185 );
    and g8068 ( n11243 , n14063 , n11850 );
    or g8069 ( n11265 , n3569 , n7473 );
    nor g8070 ( n13573 , n2684 , n9629 );
    nor g8071 ( n13595 , n7624 , n6840 );
    not g8072 ( n3062 , n4720 );
    and g8073 ( n8606 , n11422 , n11006 );
    or g8074 ( n1864 , n1494 , n5529 );
    or g8075 ( n12164 , n791 , n10095 );
    and g8076 ( n5517 , n7060 , n9825 );
    or g8077 ( n6977 , n2518 , n12701 );
    or g8078 ( n3842 , n14198 , n1413 );
    not g8079 ( n11688 , n11529 );
    not g8080 ( n9423 , n6274 );
    and g8081 ( n8935 , n12990 , n1029 );
    and g8082 ( n13261 , n1526 , n67 );
    or g8083 ( n13735 , n8638 , n13995 );
    and g8084 ( n1298 , n10302 , n1846 );
    or g8085 ( n7125 , n6111 , n603 );
    or g8086 ( n8194 , n2401 , n6868 );
    or g8087 ( n14177 , n7076 , n5927 );
    not g8088 ( n13885 , n12249 );
    or g8089 ( n13928 , n1875 , n1585 );
    and g8090 ( n9294 , n7693 , n12652 );
    or g8091 ( n8185 , n13978 , n11563 );
    or g8092 ( n13948 , n950 , n2662 );
    or g8093 ( n11035 , n13118 , n5490 );
    or g8094 ( n1355 , n10960 , n5882 );
    and g8095 ( n4030 , n10763 , n14231 );
    and g8096 ( n11665 , n7961 , n8351 );
    or g8097 ( n4190 , n8151 , n2267 );
    not g8098 ( n7756 , n8220 );
    and g8099 ( n10889 , n7871 , n3015 );
    not g8100 ( n3047 , n10108 );
    or g8101 ( n9341 , n48 , n7707 );
    or g8102 ( n7584 , n6517 , n6999 );
    or g8103 ( n10551 , n14188 , n13496 );
    and g8104 ( n2280 , n6167 , n870 );
    and g8105 ( n6995 , n8786 , n8713 );
    or g8106 ( n5559 , n12100 , n4384 );
    or g8107 ( n5866 , n1840 , n12646 );
    or g8108 ( n11881 , n7249 , n8188 );
    and g8109 ( n2033 , n8849 , n2254 );
    or g8110 ( n7139 , n6971 , n2120 );
    not g8111 ( n12034 , n426 );
    or g8112 ( n6691 , n6109 , n3334 );
    or g8113 ( n12257 , n820 , n5736 );
    or g8114 ( n14184 , n7227 , n3441 );
    nor g8115 ( n13632 , n6428 , n13844 );
    or g8116 ( n6549 , n4828 , n10849 );
    and g8117 ( n12036 , n8386 , n11729 );
    not g8118 ( n7920 , n5178 );
    not g8119 ( n1820 , n6804 );
    and g8120 ( n2225 , n3715 , n14316 );
    nor g8121 ( n9170 , n3546 , n9090 );
    and g8122 ( n13066 , n8250 , n1153 );
    and g8123 ( n2144 , n5312 , n4820 );
    or g8124 ( n8657 , n11117 , n3833 );
    and g8125 ( n3644 , n10922 , n13512 );
    and g8126 ( n10616 , n11329 , n10532 );
    and g8127 ( n4203 , n4744 , n8049 );
    or g8128 ( n13137 , n13501 , n7602 );
    and g8129 ( n13328 , n14063 , n11293 );
    and g8130 ( n4989 , n8427 , n7727 );
    or g8131 ( n7872 , n8513 , n12725 );
    and g8132 ( n6131 , n9102 , n2066 );
    not g8133 ( n1462 , n7533 );
    and g8134 ( n6351 , n9564 , n12496 );
    or g8135 ( n1831 , n1223 , n7674 );
    not g8136 ( n6527 , n11548 );
    and g8137 ( n6232 , n13555 , n4461 );
    and g8138 ( n4437 , n8044 , n11641 );
    and g8139 ( n4617 , n6838 , n2835 );
    or g8140 ( n13824 , n9620 , n5617 );
    not g8141 ( n5986 , n238 );
    not g8142 ( n5148 , n6266 );
    nor g8143 ( n1309 , n6313 , n10785 );
    nor g8144 ( n10641 , n5468 , n3928 );
    nor g8145 ( n1063 , n13061 , n115 );
    or g8146 ( n2696 , n2218 , n6227 );
    nor g8147 ( n12035 , n10179 , n13438 );
    not g8148 ( n2760 , n10426 );
    or g8149 ( n3759 , n9620 , n6980 );
    or g8150 ( n12473 , n6206 , n5760 );
    or g8151 ( n14420 , n4899 , n7107 );
    or g8152 ( n10821 , n5180 , n13319 );
    nor g8153 ( n3104 , n2624 , n8564 );
    and g8154 ( n12151 , n9052 , n5461 );
    not g8155 ( n6383 , n10407 );
    not g8156 ( n5414 , n5009 );
    and g8157 ( n9455 , n5948 , n14298 );
    nor g8158 ( n5022 , n2212 , n5735 );
    and g8159 ( n13099 , n12425 , n8584 );
    and g8160 ( n12859 , n3212 , n10063 );
    not g8161 ( n14029 , n565 );
    and g8162 ( n8074 , n4722 , n118 );
    not g8163 ( n848 , n1093 );
    nor g8164 ( n4696 , n2332 , n13371 );
    not g8165 ( n1722 , n11493 );
    or g8166 ( n7903 , n12353 , n2284 );
    or g8167 ( n1862 , n13806 , n7101 );
    not g8168 ( n12042 , n3309 );
    and g8169 ( n13320 , n5458 , n12379 );
    nor g8170 ( n4730 , n648 , n12315 );
    and g8171 ( n3244 , n5857 , n5754 );
    and g8172 ( n9273 , n11816 , n5666 );
    or g8173 ( n1503 , n8980 , n9451 );
    not g8174 ( n9218 , n4149 );
    and g8175 ( n2905 , n7961 , n8013 );
    or g8176 ( n1295 , n13446 , n13934 );
    or g8177 ( n6558 , n7436 , n9784 );
    or g8178 ( n819 , n12820 , n3573 );
    or g8179 ( n4192 , n12764 , n11602 );
    or g8180 ( n8584 , n390 , n10075 );
    and g8181 ( n958 , n3755 , n3885 );
    or g8182 ( n3756 , n2843 , n13562 );
    or g8183 ( n4583 , n3099 , n4434 );
    or g8184 ( n1995 , n1061 , n3503 );
    or g8185 ( n10226 , n5603 , n3731 );
    not g8186 ( n14472 , n1894 );
    not g8187 ( n7448 , n53 );
    and g8188 ( n9334 , n10197 , n6749 );
    or g8189 ( n9788 , n7229 , n8346 );
    or g8190 ( n7301 , n1258 , n180 );
    or g8191 ( n12690 , n317 , n7167 );
    or g8192 ( n4372 , n7914 , n9997 );
    and g8193 ( n5643 , n457 , n6508 );
    and g8194 ( n7716 , n10134 , n4113 );
    and g8195 ( n9817 , n7911 , n10840 );
    and g8196 ( n4621 , n9509 , n5103 );
    and g8197 ( n12523 , n9853 , n10415 );
    not g8198 ( n11967 , n2644 );
    nor g8199 ( n12143 , n8511 , n1307 );
    and g8200 ( n10165 , n1074 , n10838 );
    nor g8201 ( n6515 , n12280 , n6358 );
    and g8202 ( n5650 , n13520 , n1631 );
    or g8203 ( n7897 , n14107 , n178 );
    and g8204 ( n932 , n1699 , n11321 );
    and g8205 ( n9616 , n4573 , n5127 );
    not g8206 ( n5582 , n9046 );
    or g8207 ( n690 , n12712 , n13667 );
    or g8208 ( n8502 , n10936 , n1749 );
    or g8209 ( n3717 , n12100 , n12203 );
    and g8210 ( n4501 , n4359 , n12835 );
    and g8211 ( n1032 , n2180 , n10772 );
    and g8212 ( n6372 , n10458 , n10284 );
    or g8213 ( n14137 , n10191 , n2504 );
    or g8214 ( n11002 , n12353 , n8791 );
    and g8215 ( n6742 , n1447 , n14039 );
    and g8216 ( n95 , n11495 , n7098 );
    or g8217 ( n3322 , n11724 , n1349 );
    not g8218 ( n10428 , n12121 );
    or g8219 ( n696 , n10394 , n11451 );
    or g8220 ( n9588 , n8452 , n4206 );
    not g8221 ( n7802 , n6364 );
    and g8222 ( n11363 , n11411 , n9412 );
    and g8223 ( n6200 , n10166 , n4472 );
    not g8224 ( n13407 , n8555 );
    not g8225 ( n6657 , n5872 );
    or g8226 ( n8240 , n13706 , n14505 );
    and g8227 ( n211 , n6838 , n347 );
    and g8228 ( n2604 , n9953 , n2248 );
    or g8229 ( n9491 , n2086 , n10185 );
    and g8230 ( n12570 , n2709 , n9448 );
    or g8231 ( n3570 , n8172 , n14149 );
    and g8232 ( n9141 , n3169 , n5083 );
    or g8233 ( n5330 , n8452 , n188 );
    or g8234 ( n9048 , n3093 , n12762 );
    nor g8235 ( n2360 , n14133 , n4142 );
    not g8236 ( n8663 , n3587 );
    nor g8237 ( n13377 , n12483 , n13337 );
    or g8238 ( n5962 , n5986 , n6774 );
    or g8239 ( n12301 , n5815 , n6689 );
    or g8240 ( n10094 , n85 , n1143 );
    or g8241 ( n10187 , n10933 , n9579 );
    nor g8242 ( n795 , n5977 , n6887 );
    not g8243 ( n4788 , n10269 );
    not g8244 ( n7065 , n1357 );
    and g8245 ( n8166 , n11607 , n11887 );
    and g8246 ( n9584 , n3586 , n2787 );
    and g8247 ( n12856 , n10815 , n2340 );
    nor g8248 ( n7788 , n4046 , n3899 );
    or g8249 ( n1404 , n3093 , n254 );
    not g8250 ( n10091 , n8572 );
    and g8251 ( n5008 , n4095 , n7525 );
    or g8252 ( n3705 , n12494 , n3314 );
    or g8253 ( n12392 , n9285 , n4675 );
    and g8254 ( n3368 , n7429 , n10325 );
    or g8255 ( n12724 , n1840 , n8060 );
    and g8256 ( n1158 , n12018 , n2628 );
    and g8257 ( n10132 , n12918 , n12760 );
    or g8258 ( n5377 , n8575 , n4228 );
    and g8259 ( n10613 , n6128 , n1525 );
    not g8260 ( n450 , n14510 );
    or g8261 ( n13785 , n11953 , n557 );
    and g8262 ( n6915 , n12460 , n13655 );
    not g8263 ( n13840 , n5185 );
    not g8264 ( n1834 , n3070 );
    or g8265 ( n9156 , n3561 , n14163 );
    and g8266 ( n3140 , n8401 , n10298 );
    and g8267 ( n1959 , n348 , n4949 );
    and g8268 ( n1991 , n13535 , n4626 );
    or g8269 ( n11891 , n2016 , n7469 );
    and g8270 ( n3197 , n6822 , n12831 );
    or g8271 ( n11029 , n4128 , n6793 );
    and g8272 ( n7795 , n8111 , n1328 );
    and g8273 ( n8294 , n13433 , n13580 );
    and g8274 ( n13267 , n457 , n1097 );
    and g8275 ( n12145 , n7768 , n236 );
    or g8276 ( n12488 , n2272 , n10042 );
    or g8277 ( n9763 , n12870 , n3471 );
    or g8278 ( n13015 , n2750 , n1751 );
    and g8279 ( n8133 , n12389 , n11182 );
    and g8280 ( n1985 , n7230 , n7401 );
    or g8281 ( n2109 , n10713 , n7273 );
    and g8282 ( n4224 , n5926 , n6732 );
    not g8283 ( n12683 , n7575 );
    or g8284 ( n14054 , n9218 , n2033 );
    not g8285 ( n10913 , n2970 );
    and g8286 ( n11797 , n4276 , n11655 );
    and g8287 ( n9053 , n718 , n1882 );
    or g8288 ( n9011 , n839 , n2060 );
    and g8289 ( n6177 , n12449 , n4728 );
    and g8290 ( n5645 , n14357 , n5484 );
    nor g8291 ( n1534 , n4207 , n4652 );
    and g8292 ( n8343 , n5335 , n5835 );
    or g8293 ( n13403 , n11620 , n3509 );
    and g8294 ( n8311 , n2091 , n13990 );
    or g8295 ( n2704 , n553 , n10096 );
    nor g8296 ( n5914 , n6428 , n6622 );
    and g8297 ( n1905 , n1662 , n11193 );
    or g8298 ( n3770 , n10534 , n8228 );
    and g8299 ( n6439 , n7284 , n11892 );
    or g8300 ( n2265 , n14029 , n14048 );
    and g8301 ( n10927 , n776 , n10472 );
    and g8302 ( n1727 , n9188 , n3206 );
    and g8303 ( n6248 , n2091 , n11485 );
    or g8304 ( n12698 , n10781 , n13308 );
    or g8305 ( n780 , n4822 , n12974 );
    not g8306 ( n10556 , n9613 );
    or g8307 ( n9398 , n11036 , n13849 );
    and g8308 ( n10691 , n2820 , n2916 );
    nor g8309 ( n13993 , n478 , n1899 );
    not g8310 ( n9617 , n1436 );
    and g8311 ( n6361 , n2177 , n9243 );
    or g8312 ( n4710 , n7250 , n195 );
    nor g8313 ( n4582 , n8663 , n9847 );
    not g8314 ( n8942 , n1780 );
    or g8315 ( n6155 , n1494 , n10898 );
    or g8316 ( n6245 , n5454 , n4784 );
    not g8317 ( n14466 , n10204 );
    or g8318 ( n9655 , n4199 , n3266 );
    and g8319 ( n11252 , n536 , n6652 );
    not g8320 ( n8580 , n5549 );
    and g8321 ( n13600 , n8923 , n722 );
    not g8322 ( n14501 , n2257 );
    nor g8323 ( n13776 , n11445 , n14324 );
    not g8324 ( n474 , n5029 );
    or g8325 ( n9528 , n7481 , n11387 );
    or g8326 ( n2457 , n2694 , n14193 );
    not g8327 ( n6867 , n6978 );
    or g8328 ( n728 , n12295 , n1710 );
    or g8329 ( n1252 , n7249 , n10865 );
    nor g8330 ( n3351 , n2194 , n9888 );
    and g8331 ( n607 , n5053 , n8230 );
    and g8332 ( n455 , n12721 , n10249 );
    or g8333 ( n5949 , n13432 , n391 );
    nor g8334 ( n9629 , n1383 , n3621 );
    or g8335 ( n7447 , n2897 , n14372 );
    or g8336 ( n9358 , n9747 , n6624 );
    nor g8337 ( n8829 , n6011 , n6116 );
    and g8338 ( n5319 , n12018 , n9752 );
    and g8339 ( n6086 , n333 , n12942 );
    or g8340 ( n3690 , n11405 , n9728 );
    and g8341 ( n5568 , n6838 , n4043 );
    and g8342 ( n2444 , n2486 , n2673 );
    and g8343 ( n2647 , n12101 , n11571 );
    or g8344 ( n5363 , n2761 , n10265 );
    and g8345 ( n1514 , n12990 , n1156 );
    or g8346 ( n6495 , n2016 , n13595 );
    or g8347 ( n7343 , n6690 , n7293 );
    and g8348 ( n7080 , n4156 , n13211 );
    or g8349 ( n10040 , n13112 , n14454 );
    and g8350 ( n10236 , n1850 , n11852 );
    nor g8351 ( n5712 , n2000 , n9909 );
    nor g8352 ( n7371 , n9404 , n10811 );
    nor g8353 ( n8594 , n228 , n10391 );
    and g8354 ( n7457 , n2961 , n5156 );
    not g8355 ( n13650 , n14293 );
    nor g8356 ( n12060 , n4233 , n14080 );
    nor g8357 ( n2052 , n1838 , n12035 );
    nor g8358 ( n8645 , n11428 , n13986 );
    nor g8359 ( n10441 , n3959 , n8874 );
    or g8360 ( n9116 , n8301 , n378 );
    or g8361 ( n10919 , n6271 , n12001 );
    not g8362 ( n3107 , n1997 );
    or g8363 ( n14405 , n12576 , n7543 );
    and g8364 ( n7102 , n10556 , n2681 );
    nor g8365 ( n7281 , n5160 , n7811 );
    or g8366 ( n5812 , n2111 , n13500 );
    and g8367 ( n3520 , n11093 , n7593 );
    nor g8368 ( n6089 , n14198 , n1280 );
    and g8369 ( n7698 , n12404 , n8348 );
    and g8370 ( n13307 , n541 , n4556 );
    and g8371 ( n12661 , n8453 , n912 );
    or g8372 ( n1803 , n4195 , n10859 );
    and g8373 ( n3480 , n4880 , n1191 );
    nor g8374 ( n4651 , n6085 , n4944 );
    or g8375 ( n540 , n4468 , n1170 );
    and g8376 ( n3872 , n1876 , n8904 );
    and g8377 ( n6516 , n3419 , n11 );
    and g8378 ( n13024 , n3715 , n7435 );
    not g8379 ( n1769 , n10380 );
    or g8380 ( n13589 , n3826 , n13272 );
    not g8381 ( n5959 , n6387 );
    and g8382 ( n2159 , n10032 , n12325 );
    nor g8383 ( n5404 , n14106 , n14271 );
    and g8384 ( n10341 , n11362 , n1056 );
    nor g8385 ( n6529 , n9529 , n7701 );
    and g8386 ( n6655 , n10197 , n6843 );
    not g8387 ( n3813 , n1473 );
    not g8388 ( n10408 , n7275 );
    not g8389 ( n955 , n9272 );
    not g8390 ( n11329 , n13003 );
    and g8391 ( n14240 , n8213 , n4479 );
    and g8392 ( n6275 , n666 , n12627 );
    nor g8393 ( n12955 , n4313 , n14186 );
    not g8394 ( n6654 , n12588 );
    and g8395 ( n5034 , n13597 , n11175 );
    or g8396 ( n2898 , n5710 , n2827 );
    not g8397 ( n14521 , n11961 );
    or g8398 ( n10225 , n9107 , n2332 );
    and g8399 ( n2484 , n3623 , n235 );
    nor g8400 ( n6335 , n6030 , n7524 );
    or g8401 ( n1661 , n8490 , n6726 );
    or g8402 ( n804 , n4602 , n6479 );
    not g8403 ( n9188 , n6819 );
    or g8404 ( n2679 , n930 , n643 );
    and g8405 ( n12675 , n13507 , n4831 );
    or g8406 ( n6764 , n11472 , n574 );
    and g8407 ( n8634 , n7443 , n13955 );
    or g8408 ( n7996 , n1741 , n7968 );
    not g8409 ( n4824 , n241 );
    and g8410 ( n2059 , n11316 , n2288 );
    nor g8411 ( n7692 , n3577 , n12978 );
    not g8412 ( n9142 , n12025 );
    not g8413 ( n355 , n7915 );
    or g8414 ( n4241 , n10539 , n6850 );
    nor g8415 ( n3928 , n13255 , n4280 );
    or g8416 ( n2340 , n13978 , n12509 );
    and g8417 ( n12596 , n3485 , n5745 );
    and g8418 ( n6945 , n7961 , n7654 );
    nor g8419 ( n9277 , n1914 , n3823 );
    and g8420 ( n8599 , n5459 , n13643 );
    not g8421 ( n2461 , n9865 );
    and g8422 ( n136 , n8453 , n4750 );
    nor g8423 ( n1707 , n5018 , n11562 );
    and g8424 ( n2301 , n2643 , n73 );
    and g8425 ( n4456 , n12857 , n6930 );
    not g8426 ( n10191 , n628 );
    nor g8427 ( n10065 , n8424 , n14254 );
    nor g8428 ( n13244 , n5715 , n2245 );
    nor g8429 ( n9021 , n13429 , n8901 );
    not g8430 ( n10897 , n11325 );
    nor g8431 ( n14112 , n12244 , n10830 );
    and g8432 ( n12907 , n6531 , n1404 );
    or g8433 ( n7034 , n4899 , n7224 );
    or g8434 ( n4248 , n12927 , n10050 );
    and g8435 ( n517 , n4358 , n12114 );
    not g8436 ( n2910 , n7584 );
    or g8437 ( n8742 , n3709 , n1763 );
    not g8438 ( n1843 , n13425 );
    or g8439 ( n2680 , n930 , n10067 );
    or g8440 ( n9479 , n2901 , n13905 );
    not g8441 ( n12857 , n11771 );
    or g8442 ( n4820 , n11953 , n242 );
    nor g8443 ( n11125 , n234 , n3252 );
    not g8444 ( n6854 , n6807 );
    and g8445 ( n12327 , n12449 , n7225 );
    or g8446 ( n11179 , n11472 , n1437 );
    and g8447 ( n9158 , n1962 , n14274 );
    not g8448 ( n11697 , n1868 );
    not g8449 ( n10846 , n4225 );
    or g8450 ( n209 , n13978 , n2735 );
    or g8451 ( n3399 , n2111 , n272 );
    or g8452 ( n6402 , n11379 , n4425 );
    not g8453 ( n550 , n5502 );
    or g8454 ( n3627 , n12428 , n13866 );
    and g8455 ( n7831 , n3405 , n13974 );
    and g8456 ( n4838 , n11867 , n12628 );
    or g8457 ( n1275 , n5491 , n12769 );
    not g8458 ( n11336 , n2692 );
    and g8459 ( n6795 , n3169 , n1400 );
    and g8460 ( n13765 , n12528 , n1388 );
    and g8461 ( n13851 , n129 , n8593 );
    or g8462 ( n13599 , n2874 , n12217 );
    and g8463 ( n2636 , n2486 , n1457 );
    and g8464 ( n11283 , n3628 , n10307 );
    nor g8465 ( n12273 , n3394 , n8466 );
    or g8466 ( n545 , n11909 , n249 );
    or g8467 ( n10216 , n4899 , n3757 );
    or g8468 ( n4460 , n2531 , n14041 );
    or g8469 ( n1964 , n6288 , n8413 );
    not g8470 ( n1686 , n5195 );
    and g8471 ( n5387 , n1924 , n3236 );
    and g8472 ( n5685 , n4803 , n1671 );
    or g8473 ( n12682 , n12820 , n4161 );
    not g8474 ( n13394 , n10314 );
    and g8475 ( n2862 , n10408 , n3620 );
    or g8476 ( n12657 , n9742 , n13567 );
    or g8477 ( n13167 , n10523 , n11296 );
    not g8478 ( n582 , n4172 );
    nor g8479 ( n2515 , n11990 , n14101 );
    and g8480 ( n2572 , n3263 , n13334 );
    and g8481 ( n490 , n10615 , n10843 );
    and g8482 ( n12977 , n5582 , n1578 );
    nor g8483 ( n1513 , n6085 , n7024 );
    or g8484 ( n2271 , n5861 , n1318 );
    and g8485 ( n12755 , n9745 , n5133 );
    or g8486 ( n11521 , n11951 , n12733 );
    or g8487 ( n7570 , n13547 , n1735 );
    nor g8488 ( n9820 , n3395 , n11924 );
    or g8489 ( n9539 , n11542 , n14125 );
    or g8490 ( n9027 , n3161 , n7823 );
    and g8491 ( n11433 , n7691 , n8898 );
    and g8492 ( n8145 , n6243 , n3346 );
    not g8493 ( n10705 , n10400 );
    not g8494 ( n13118 , n13901 );
    and g8495 ( n7262 , n13520 , n11918 );
    not g8496 ( n11551 , n4847 );
    or g8497 ( n3801 , n619 , n9866 );
    and g8498 ( n4493 , n4932 , n9454 );
    not g8499 ( n9754 , n461 );
    not g8500 ( n12020 , n1010 );
    or g8501 ( n2655 , n4631 , n12716 );
    nor g8502 ( n12605 , n5278 , n5849 );
    or g8503 ( n13 , n2908 , n6329 );
    not g8504 ( n6525 , n1724 );
    and g8505 ( n7285 , n2820 , n1141 );
    or g8506 ( n4869 , n9111 , n1636 );
    or g8507 ( n1448 , n9403 , n8336 );
    and g8508 ( n1795 , n6531 , n4474 );
    or g8509 ( n13288 , n5570 , n11003 );
    nor g8510 ( n14130 , n11581 , n2543 );
    not g8511 ( n8569 , n9592 );
    and g8512 ( n14051 , n6157 , n11026 );
    nor g8513 ( n12274 , n2415 , n6572 );
    nor g8514 ( n454 , n3871 , n526 );
    or g8515 ( n7274 , n3877 , n6922 );
    or g8516 ( n59 , n8897 , n3754 );
    and g8517 ( n10424 , n12039 , n5637 );
    and g8518 ( n7540 , n13297 , n3495 );
    nor g8519 ( n989 , n8065 , n10425 );
    or g8520 ( n14302 , n12633 , n13622 );
    nor g8521 ( n8671 , n5715 , n5989 );
    not g8522 ( n11493 , n6326 );
    not g8523 ( n7970 , n7278 );
    and g8524 ( n5314 , n11313 , n9036 );
    and g8525 ( n13332 , n5471 , n895 );
    nor g8526 ( n6137 , n5435 , n6816 );
    not g8527 ( n4963 , n4953 );
    and g8528 ( n65 , n3485 , n5752 );
    and g8529 ( n11813 , n4786 , n4859 );
    not g8530 ( n438 , n12850 );
    or g8531 ( n8576 , n9977 , n13890 );
    or g8532 ( n12094 , n227 , n12863 );
    and g8533 ( n5332 , n6318 , n4416 );
    or g8534 ( n14237 , n9620 , n6280 );
    or g8535 ( n5273 , n13276 , n5227 );
    nor g8536 ( n4760 , n13722 , n2276 );
    or g8537 ( n14004 , n8881 , n7326 );
    and g8538 ( n2258 , n4525 , n11644 );
    and g8539 ( n12418 , n13103 , n1890 );
    or g8540 ( n8741 , n817 , n14085 );
    or g8541 ( n9758 , n9490 , n2004 );
    not g8542 ( n9747 , n81 );
    not g8543 ( n3277 , n11765 );
    and g8544 ( n1089 , n446 , n6663 );
    nor g8545 ( n11275 , n6544 , n5663 );
    and g8546 ( n401 , n9617 , n4746 );
    or g8547 ( n8946 , n14110 , n8516 );
    not g8548 ( n5026 , n11130 );
    or g8549 ( n11877 , n12139 , n7280 );
    nor g8550 ( n9239 , n1112 , n14390 );
    not g8551 ( n8528 , n2201 );
    or g8552 ( n423 , n9226 , n544 );
    or g8553 ( n4695 , n7359 , n7129 );
    or g8554 ( n14053 , n5732 , n11504 );
    and g8555 ( n6974 , n3 , n2858 );
    and g8556 ( n6287 , n13952 , n9368 );
    and g8557 ( n4500 , n3675 , n4763 );
    and g8558 ( n10576 , n11403 , n5316 );
    nor g8559 ( n3462 , n6422 , n7313 );
    or g8560 ( n12452 , n8747 , n11917 );
    or g8561 ( n7579 , n7426 , n107 );
    nor g8562 ( n11634 , n9388 , n1040 );
    or g8563 ( n10832 , n2246 , n9499 );
    or g8564 ( n11261 , n13991 , n6589 );
    not g8565 ( n12130 , n8272 );
    or g8566 ( n13134 , n8015 , n5440 );
    or g8567 ( n11396 , n14166 , n13018 );
    nor g8568 ( n11630 , n1112 , n7634 );
    not g8569 ( n5861 , n13165 );
    or g8570 ( n6947 , n11121 , n14073 );
    and g8571 ( n7511 , n3268 , n10658 );
    and g8572 ( n9869 , n13626 , n5838 );
    and g8573 ( n4873 , n5011 , n8639 );
    not g8574 ( n12483 , n746 );
    and g8575 ( n10013 , n8786 , n1057 );
    not g8576 ( n13350 , n11809 );
    or g8577 ( n12562 , n2874 , n2182 );
    nor g8578 ( n4889 , n7407 , n6327 );
    or g8579 ( n3606 , n781 , n11922 );
    and g8580 ( n10587 , n200 , n5420 );
    and g8581 ( n11942 , n11329 , n10990 );
    and g8582 ( n4221 , n80 , n6524 );
    and g8583 ( n3493 , n7308 , n14229 );
    and g8584 ( n2918 , n14118 , n736 );
    and g8585 ( n7908 , n7717 , n6412 );
    or g8586 ( n8142 , n7914 , n8761 );
    not g8587 ( n14446 , n10322 );
    or g8588 ( n4670 , n5569 , n5648 );
    and g8589 ( n6043 , n3370 , n6208 );
    or g8590 ( n4097 , n9285 , n7039 );
    and g8591 ( n5806 , n7652 , n11206 );
    and g8592 ( n6699 , n392 , n3701 );
    or g8593 ( n8278 , n9403 , n5174 );
    nor g8594 ( n8882 , n1152 , n1388 );
    and g8595 ( n9687 , n9724 , n12031 );
    not g8596 ( n11481 , n11967 );
    or g8597 ( n4530 , n8096 , n7541 );
    and g8598 ( n4996 , n6013 , n3420 );
    and g8599 ( n777 , n11743 , n6794 );
    and g8600 ( n2359 , n10072 , n2406 );
    and g8601 ( n8644 , n6724 , n8653 );
    and g8602 ( n1580 , n5012 , n12054 );
    not g8603 ( n6413 , n10403 );
    or g8604 ( n5694 , n7156 , n6719 );
    and g8605 ( n8052 , n5779 , n7966 );
    or g8606 ( n9364 , n77 , n7784 );
    or g8607 ( n7556 , n4162 , n4998 );
    and g8608 ( n11195 , n4365 , n6948 );
    not g8609 ( n10368 , n834 );
    and g8610 ( n902 , n3932 , n1484 );
    not g8611 ( n4525 , n304 );
    and g8612 ( n3092 , n7943 , n13453 );
    and g8613 ( n739 , n5574 , n3214 );
    and g8614 ( n4251 , n12039 , n7261 );
    or g8615 ( n5228 , n636 , n3506 );
    and g8616 ( n9801 , n14120 , n2131 );
    not g8617 ( n3332 , n5288 );
    nor g8618 ( n9066 , n7375 , n3170 );
    or g8619 ( n3839 , n12764 , n3078 );
    not g8620 ( n1875 , n630 );
    and g8621 ( n534 , n904 , n3371 );
    or g8622 ( n12786 , n4899 , n11058 );
    or g8623 ( n2638 , n10933 , n5619 );
    not g8624 ( n6899 , n2919 );
    or g8625 ( n4024 , n2949 , n4042 );
    not g8626 ( n1742 , n10115 );
    or g8627 ( n13831 , n2017 , n7028 );
    or g8628 ( n135 , n8045 , n10893 );
    and g8629 ( n7679 , n5252 , n7724 );
    or g8630 ( n6382 , n11739 , n13499 );
    nor g8631 ( n11096 , n7245 , n13498 );
    or g8632 ( n7833 , n4821 , n11388 );
    not g8633 ( n2409 , n2566 );
    or g8634 ( n4189 , n478 , n11695 );
    and g8635 ( n12232 , n13102 , n2690 );
    or g8636 ( n14398 , n9931 , n7815 );
    not g8637 ( n5848 , n11515 );
    and g8638 ( n1783 , n11153 , n9336 );
    or g8639 ( n3340 , n6824 , n3835 );
    or g8640 ( n499 , n3193 , n3792 );
    or g8641 ( n9713 , n13005 , n860 );
    or g8642 ( n7084 , n14370 , n11156 );
    not g8643 ( n5857 , n1724 );
    or g8644 ( n11522 , n13413 , n4186 );
    or g8645 ( n13886 , n2518 , n14393 );
    and g8646 ( n9737 , n13240 , n2565 );
    and g8647 ( n13189 , n4346 , n12585 );
    or g8648 ( n14189 , n69 , n6674 );
    or g8649 ( n5522 , n1805 , n3849 );
    and g8650 ( n11038 , n12986 , n7501 );
    nor g8651 ( n5518 , n6413 , n13989 );
    or g8652 ( n14059 , n11121 , n3806 );
    or g8653 ( n2842 , n5253 , n5701 );
    not g8654 ( n2405 , n5117 );
    and g8655 ( n191 , n4359 , n5742 );
    and g8656 ( n813 , n7284 , n2142 );
    not g8657 ( n1266 , n13139 );
    or g8658 ( n4107 , n10089 , n10635 );
    or g8659 ( n1972 , n13016 , n13409 );
    and g8660 ( n3740 , n12772 , n7465 );
    nor g8661 ( n12591 , n2644 , n9714 );
    not g8662 ( n11580 , n7339 );
    and g8663 ( n8282 , n12250 , n10343 );
    and g8664 ( n4641 , n13342 , n3202 );
    and g8665 ( n12851 , n3 , n7549 );
    and g8666 ( n9028 , n13626 , n11396 );
    not g8667 ( n5418 , n12279 );
    and g8668 ( n11764 , n12185 , n1888 );
    or g8669 ( n2068 , n2874 , n10904 );
    nor g8670 ( n12739 , n500 , n7725 );
    or g8671 ( n11413 , n1875 , n10444 );
    and g8672 ( n5401 , n8427 , n4423 );
    nor g8673 ( n9560 , n3870 , n4793 );
    not g8674 ( n9673 , n1702 );
    and g8675 ( n8369 , n1699 , n6799 );
    or g8676 ( n9797 , n13854 , n2275 );
    and g8677 ( n3725 , n13745 , n8243 );
    and g8678 ( n3017 , n12421 , n13521 );
    nor g8679 ( n1277 , n2571 , n7953 );
    and g8680 ( n1079 , n550 , n1307 );
    or g8681 ( n10999 , n10245 , n2620 );
    or g8682 ( n7142 , n11710 , n13460 );
    or g8683 ( n6504 , n6891 , n13771 );
    or g8684 ( n8665 , n2181 , n328 );
    and g8685 ( n281 , n7057 , n1796 );
    and g8686 ( n12498 , n6724 , n9725 );
    not g8687 ( n5628 , n5427 );
    nor g8688 ( n6816 , n13714 , n2524 );
    nor g8689 ( n3991 , n7352 , n488 );
    and g8690 ( n3700 , n11950 , n5691 );
    and g8691 ( n6509 , n2846 , n11214 );
    and g8692 ( n12917 , n13407 , n13834 );
    nor g8693 ( n6712 , n9703 , n8796 );
    and g8694 ( n11480 , n3607 , n11691 );
    or g8695 ( n13129 , n8476 , n445 );
    not g8696 ( n1857 , n8008 );
    or g8697 ( n9209 , n2387 , n7599 );
    not g8698 ( n6206 , n2794 );
    or g8699 ( n6398 , n9403 , n3880 );
    or g8700 ( n7597 , n5710 , n1905 );
    nor g8701 ( n1106 , n2969 , n13681 );
    not g8702 ( n8607 , n1334 );
    or g8703 ( n10552 , n3867 , n700 );
    and g8704 ( n6309 , n4445 , n5642 );
    not g8705 ( n8789 , n7808 );
    and g8706 ( n5061 , n2724 , n6779 );
    and g8707 ( n5630 , n3861 , n5049 );
    and g8708 ( n14212 , n12202 , n12818 );
    not g8709 ( n10855 , n11474 );
    nor g8710 ( n1546 , n162 , n7761 );
    and g8711 ( n12089 , n14373 , n2653 );
    or g8712 ( n7796 , n7527 , n1389 );
    and g8713 ( n1045 , n8812 , n2012 );
    and g8714 ( n5371 , n7745 , n7576 );
    and g8715 ( n2672 , n9977 , n3970 );
    or g8716 ( n14457 , n1147 , n11254 );
    and g8717 ( n14119 , n5317 , n366 );
    and g8718 ( n4962 , n4098 , n8820 );
    nor g8719 ( n9506 , n12107 , n11928 );
    and g8720 ( n14001 , n9080 , n1977 );
    or g8721 ( n12825 , n11011 , n7685 );
    and g8722 ( n11657 , n13860 , n4066 );
    or g8723 ( n13192 , n9285 , n13439 );
    and g8724 ( n4957 , n4346 , n5380 );
    and g8725 ( n4005 , n8372 , n7178 );
    or g8726 ( n4522 , n1223 , n12948 );
    and g8727 ( n13942 , n7677 , n10381 );
    and g8728 ( n1567 , n1414 , n5145 );
    or g8729 ( n6484 , n2874 , n7719 );
    and g8730 ( n2611 , n1059 , n8742 );
    or g8731 ( n4003 , n5833 , n8369 );
    and g8732 ( n2997 , n9920 , n240 );
    and g8733 ( n9903 , n9953 , n214 );
    not g8734 ( n10154 , n13901 );
    or g8735 ( n416 , n679 , n13109 );
    or g8736 ( n9854 , n7683 , n122 );
    and g8737 ( n2555 , n541 , n4260 );
    and g8738 ( n4446 , n5240 , n2 );
    nor g8739 ( n5722 , n9618 , n8578 );
    not g8740 ( n3247 , n12107 );
    or g8741 ( n9344 , n12712 , n8802 );
    and g8742 ( n5341 , n9232 , n4253 );
    and g8743 ( n12370 , n13103 , n8442 );
    nor g8744 ( n1064 , n1760 , n6997 );
    and g8745 ( n6735 , n7327 , n8992 );
    or g8746 ( n13450 , n1711 , n6839 );
    and g8747 ( n9100 , n4657 , n1250 );
    or g8748 ( n2966 , n8304 , n4405 );
    or g8749 ( n3843 , n2055 , n6785 );
    and g8750 ( n8060 , n2465 , n14386 );
    and g8751 ( n1928 , n1520 , n4648 );
    or g8752 ( n11801 , n6046 , n8848 );
    or g8753 ( n11944 , n568 , n9201 );
    and g8754 ( n7552 , n13433 , n2801 );
    and g8755 ( n3245 , n13379 , n2162 );
    nor g8756 ( n13306 , n4988 , n11634 );
    or g8757 ( n1163 , n8828 , n9105 );
    or g8758 ( n1561 , n7448 , n2923 );
    and g8759 ( n10656 , n7596 , n3782 );
    not g8760 ( n2098 , n12249 );
    not g8761 ( n6323 , n4465 );
    and g8762 ( n13534 , n14157 , n5698 );
    or g8763 ( n549 , n2874 , n3010 );
    or g8764 ( n12798 , n10857 , n2485 );
    and g8765 ( n1413 , n4757 , n2730 );
    and g8766 ( n13172 , n13863 , n13461 );
    and g8767 ( n2477 , n7427 , n368 );
    or g8768 ( n634 , n9716 , n2135 );
    and g8769 ( n8390 , n5458 , n3562 );
    and g8770 ( n4845 , n627 , n2685 );
    nor g8771 ( n8902 , n11040 , n2530 );
    and g8772 ( n14356 , n13096 , n311 );
    and g8773 ( n335 , n12412 , n5758 );
    and g8774 ( n13478 , n3710 , n12154 );
    or g8775 ( n8822 , n9766 , n4039 );
    and g8776 ( n7968 , n8769 , n10266 );
    nor g8777 ( n9177 , n7359 , n6072 );
    or g8778 ( n10098 , n12601 , n6417 );
    nor g8779 ( n9668 , n1820 , n3920 );
    nor g8780 ( n2726 , n8023 , n8360 );
    not g8781 ( n12202 , n14524 );
    not g8782 ( n13464 , n5795 );
    not g8783 ( n4828 , n8595 );
    and g8784 ( n13622 , n3424 , n11864 );
    or g8785 ( n113 , n9269 , n10540 );
    and g8786 ( n9306 , n12714 , n11444 );
    nor g8787 ( n2483 , n11285 , n9553 );
    not g8788 ( n4422 , n4618 );
    and g8789 ( n3417 , n12147 , n867 );
    and g8790 ( n5239 , n3635 , n3381 );
    not g8791 ( n4049 , n11016 );
    and g8792 ( n6948 , n6849 , n13857 );
    or g8793 ( n11567 , n5603 , n10681 );
    or g8794 ( n11177 , n12075 , n7548 );
    or g8795 ( n2453 , n3126 , n5251 );
    not g8796 ( n11498 , n12897 );
    not g8797 ( n5348 , n5108 );
    or g8798 ( n6202 , n7003 , n10692 );
    and g8799 ( n1919 , n5876 , n12944 );
    or g8800 ( n5637 , n3569 , n8619 );
    or g8801 ( n13634 , n11048 , n517 );
    or g8802 ( n9708 , n6695 , n6106 );
    or g8803 ( n9981 , n6242 , n4089 );
    and g8804 ( n4994 , n4803 , n6678 );
    or g8805 ( n7772 , n14401 , n9796 );
    or g8806 ( n801 , n5815 , n9290 );
    and g8807 ( n12877 , n10678 , n8299 );
    or g8808 ( n1249 , n2246 , n9889 );
    or g8809 ( n9075 , n9529 , n8696 );
    or g8810 ( n7830 , n2412 , n13502 );
    or g8811 ( n13917 , n6595 , n6687 );
    and g8812 ( n6777 , n7670 , n10277 );
    not g8813 ( n2401 , n12588 );
    and g8814 ( n5267 , n646 , n8502 );
    or g8815 ( n14295 , n4898 , n13385 );
    not g8816 ( n5131 , n5596 );
    or g8817 ( n2230 , n6857 , n2403 );
    and g8818 ( n9995 , n8358 , n6462 );
    or g8819 ( n2368 , n8575 , n11491 );
    not g8820 ( n7720 , n8672 );
    nor g8821 ( n13443 , n10289 , n8368 );
    or g8822 ( n7515 , n3088 , n10502 );
    nor g8823 ( n13916 , n2132 , n7837 );
    nor g8824 ( n12456 , n1820 , n5181 );
    nor g8825 ( n2623 , n12934 , n3380 );
    not g8826 ( n2154 , n2451 );
    or g8827 ( n7787 , n8582 , n3624 );
    and g8828 ( n9476 , n627 , n6181 );
    not g8829 ( n13365 , n12014 );
    and g8830 ( n13969 , n6838 , n6459 );
    or g8831 ( n3794 , n234 , n5778 );
    nor g8832 ( n12354 , n1423 , n5402 );
    or g8833 ( n12180 , n6111 , n9152 );
    and g8834 ( n8717 , n10622 , n1972 );
    or g8835 ( n2767 , n9931 , n12439 );
    or g8836 ( n2206 , n4498 , n5672 );
    and g8837 ( n12824 , n7391 , n5559 );
    or g8838 ( n6143 , n11739 , n12098 );
    nor g8839 ( n1026 , n8217 , n4231 );
    and g8840 ( n7006 , n12953 , n4429 );
    and g8841 ( n8283 , n1414 , n6842 );
    and g8842 ( n6592 , n1775 , n4596 );
    not g8843 ( n8304 , n3455 );
    and g8844 ( n3780 , n5940 , n1371 );
    or g8845 ( n2348 , n1261 , n7785 );
    or g8846 ( n11637 , n8034 , n1773 );
    and g8847 ( n13899 , n14388 , n6097 );
    or g8848 ( n4076 , n10062 , n9514 );
    or g8849 ( n13852 , n3320 , n14132 );
    or g8850 ( n10453 , n3011 , n8329 );
    or g8851 ( n4472 , n2531 , n3714 );
    or g8852 ( n2039 , n8404 , n6247 );
    and g8853 ( n11984 , n4851 , n10847 );
    or g8854 ( n2346 , n12695 , n8018 );
    not g8855 ( n4876 , n12776 );
    nor g8856 ( n3262 , n10511 , n7066 );
    not g8857 ( n12084 , n4830 );
    nor g8858 ( n4773 , n12483 , n9282 );
    nor g8859 ( n8135 , n8629 , n334 );
    and g8860 ( n13296 , n5092 , n2491 );
    or g8861 ( n7792 , n3886 , n10183 );
    nor g8862 ( n8324 , n239 , n12982 );
    and g8863 ( n3708 , n12611 , n9313 );
    or g8864 ( n1915 , n13226 , n12907 );
    or g8865 ( n2256 , n10523 , n13472 );
    or g8866 ( n944 , n6607 , n4215 );
    or g8867 ( n13845 , n5493 , n282 );
    nor g8868 ( n7702 , n6883 , n5827 );
    or g8869 ( n633 , n9780 , n5895 );
    or g8870 ( n3127 , n2747 , n9387 );
    and g8871 ( n2494 , n11422 , n8533 );
    and g8872 ( n7472 , n12404 , n10536 );
    not g8873 ( n13147 , n6787 );
    and g8874 ( n13790 , n783 , n13134 );
    and g8875 ( n9643 , n11313 , n4179 );
    not g8876 ( n7230 , n8439 );
    and g8877 ( n5110 , n9509 , n3529 );
    and g8878 ( n13880 , n3710 , n5106 );
    and g8879 ( n9354 , n3776 , n10276 );
    nor g8880 ( n9019 , n14466 , n3467 );
    nor g8881 ( n14384 , n9305 , n9634 );
    and g8882 ( n11859 , n11803 , n4120 );
    or g8883 ( n8589 , n2272 , n10105 );
    or g8884 ( n5334 , n329 , n4343 );
    or g8885 ( n12049 , n14430 , n1335 );
    nor g8886 ( n12021 , n10638 , n14517 );
    or g8887 ( n12469 , n6373 , n4538 );
    nor g8888 ( n7608 , n5833 , n12525 );
    and g8889 ( n6392 , n231 , n13110 );
    and g8890 ( n11490 , n7938 , n7838 );
    not g8891 ( n504 , n8595 );
    or g8892 ( n3917 , n7245 , n8867 );
    or g8893 ( n10489 , n9507 , n1606 );
    and g8894 ( n5743 , n3565 , n2740 );
    not g8895 ( n3667 , n5974 );
    and g8896 ( n9914 , n7063 , n6077 );
    or g8897 ( n4371 , n7551 , n6050 );
    nor g8898 ( n4808 , n9388 , n9685 );
    and g8899 ( n8678 , n12615 , n2560 );
    and g8900 ( n9256 , n6606 , n5122 );
    and g8901 ( n13385 , n13597 , n5684 );
    and g8902 ( n11949 , n12960 , n10295 );
    or g8903 ( n14383 , n2181 , n4900 );
    or g8904 ( n2601 , n8877 , n9672 );
    and g8905 ( n2479 , n2583 , n2982 );
    not g8906 ( n4631 , n3616 );
    or g8907 ( n8470 , n8210 , n4160 );
    and g8908 ( n12175 , n3366 , n2871 );
    or g8909 ( n7871 , n7484 , n6251 );
    not g8910 ( n1623 , n13696 );
    or g8911 ( n14256 , n492 , n7880 );
    and g8912 ( n8336 , n8789 , n8036 );
    or g8913 ( n4010 , n1701 , n4668 );
    or g8914 ( n2841 , n1031 , n3501 );
    and g8915 ( n8875 , n4163 , n9912 );
    or g8916 ( n5837 , n2111 , n11616 );
    and g8917 ( n6180 , n8066 , n3739 );
    and g8918 ( n7789 , n10595 , n8296 );
    and g8919 ( n14193 , n14042 , n583 );
    or g8920 ( n8833 , n4925 , n623 );
    and g8921 ( n10055 , n7938 , n1062 );
    and g8922 ( n802 , n14388 , n5260 );
    and g8923 ( n1384 , n8238 , n8985 );
    or g8924 ( n10530 , n8151 , n12053 );
    or g8925 ( n5389 , n116 , n3041 );
    and g8926 ( n9051 , n3097 , n8251 );
    nor g8927 ( n12525 , n3907 , n9969 );
    or g8928 ( n14062 , n11105 , n9006 );
    nor g8929 ( n1385 , n7575 , n9637 );
    or g8930 ( n13184 , n5472 , n6832 );
    and g8931 ( n9417 , n14446 , n819 );
    nor g8932 ( n6622 , n3344 , n5894 );
    nor g8933 ( n4344 , n7609 , n9373 );
    not g8934 ( n2315 , n2918 );
    not g8935 ( n4135 , n6534 );
    or g8936 ( n11615 , n10933 , n4957 );
    and g8937 ( n6082 , n536 , n1114 );
    and g8938 ( n8433 , n3586 , n10453 );
    nor g8939 ( n1196 , n2103 , n6439 );
    and g8940 ( n212 , n6157 , n1648 );
    or g8941 ( n4204 , n3815 , n4540 );
    or g8942 ( n6321 , n1805 , n2911 );
    or g8943 ( n5494 , n4508 , n6351 );
    nor g8944 ( n3771 , n12112 , n10122 );
    nor g8945 ( n8895 , n10309 , n13640 );
    and g8946 ( n3232 , n638 , n7856 );
    nor g8947 ( n4718 , n10363 , n10814 );
    and g8948 ( n10007 , n4788 , n12499 );
    or g8949 ( n11897 , n10626 , n10644 );
    or g8950 ( n659 , n4433 , n1222 );
    and g8951 ( n1825 , n5229 , n1479 );
    and g8952 ( n7978 , n11329 , n8912 );
    or g8953 ( n5492 , n8172 , n6653 );
    or g8954 ( n13857 , n8721 , n6680 );
    nor g8955 ( n13325 , n9806 , n2036 );
    or g8956 ( n5296 , n8096 , n2384 );
    or g8957 ( n1506 , n14273 , n8926 );
    or g8958 ( n5086 , n504 , n9891 );
    and g8959 ( n13381 , n9015 , n270 );
    not g8960 ( n10808 , n8148 );
    and g8961 ( n11589 , n11803 , n3935 );
    nor g8962 ( n5324 , n4741 , n1274 );
    not g8963 ( n5406 , n4609 );
    and g8964 ( n14389 , n9890 , n2205 );
    or g8965 ( n11228 , n14435 , n8321 );
    or g8966 ( n4047 , n14178 , n498 );
    and g8967 ( n4125 , n427 , n3104 );
    and g8968 ( n3592 , n1729 , n2211 );
    not g8969 ( n9275 , n5153 );
    or g8970 ( n13175 , n283 , n2671 );
    not g8971 ( n1409 , n5960 );
    or g8972 ( n63 , n5975 , n4022 );
    and g8973 ( n1949 , n7427 , n8690 );
    and g8974 ( n1931 , n7970 , n9633 );
    and g8975 ( n7009 , n748 , n7292 );
    and g8976 ( n14381 , n14120 , n12482 );
    or g8977 ( n4275 , n5575 , n12512 );
    and g8978 ( n8349 , n848 , n12992 );
    and g8979 ( n2520 , n3608 , n12932 );
    nor g8980 ( n10774 , n13276 , n9907 );
    and g8981 ( n6714 , n12357 , n4687 );
    not g8982 ( n446 , n6119 );
    not g8983 ( n6724 , n9994 );
    not g8984 ( n5153 , n8224 );
    or g8985 ( n257 , n14400 , n8164 );
    or g8986 ( n6852 , n10083 , n959 );
    not g8987 ( n10825 , n3284 );
    nor g8988 ( n2988 , n2919 , n537 );
    and g8989 ( n14474 , n4932 , n915 );
    and g8990 ( n11304 , n1074 , n11356 );
    nor g8991 ( n11233 , n10936 , n14250 );
    or g8992 ( n4393 , n12130 , n8978 );
    or g8993 ( n3783 , n12023 , n2336 );
    or g8994 ( n7933 , n3120 , n12619 );
    and g8995 ( n5934 , n7267 , n9487 );
    not g8996 ( n7518 , n6397 );
    and g8997 ( n13870 , n7972 , n8374 );
    or g8998 ( n12714 , n12435 , n411 );
    nor g8999 ( n2446 , n473 , n2186 );
    not g9000 ( n6254 , n11259 );
    or g9001 ( n4352 , n11379 , n8227 );
    and g9002 ( n3632 , n5104 , n9011 );
    nor g9003 ( n1375 , n1697 , n1652 );
    or g9004 ( n10004 , n8964 , n8198 );
    and g9005 ( n3760 , n11262 , n11885 );
    nor g9006 ( n11155 , n12084 , n10203 );
    nor g9007 ( n14104 , n8223 , n13584 );
    and g9008 ( n3496 , n4655 , n6992 );
    or g9009 ( n2847 , n10834 , n10102 );
    or g9010 ( n14185 , n6323 , n7853 );
    not g9011 ( n11667 , n3623 );
    or g9012 ( n12737 , n573 , n12879 );
    or g9013 ( n12377 , n1480 , n8084 );
    and g9014 ( n197 , n12425 , n12247 );
    not g9015 ( n8986 , n777 );
    and g9016 ( n8993 , n1788 , n1380 );
    and g9017 ( n12975 , n7041 , n10483 );
    and g9018 ( n12594 , n13484 , n661 );
    or g9019 ( n6142 , n11459 , n10272 );
    not g9020 ( n6660 , n7889 );
    not g9021 ( n8925 , n11232 );
    and g9022 ( n8318 , n7691 , n7651 );
    and g9023 ( n12589 , n4856 , n10984 );
    and g9024 ( n9108 , n9953 , n4832 );
    nor g9025 ( n7524 , n3445 , n13104 );
    or g9026 ( n684 , n4481 , n1240 );
    and g9027 ( n2809 , n6130 , n14202 );
    not g9028 ( n2057 , n9371 );
    or g9029 ( n10281 , n5625 , n12745 );
    or g9030 ( n12794 , n8210 , n1766 );
    not g9031 ( n14524 , n3331 );
    nor g9032 ( n526 , n3196 , n7663 );
    not g9033 ( n6159 , n6088 );
    or g9034 ( n14363 , n13516 , n3868 );
    and g9035 ( n249 , n3607 , n7215 );
    and g9036 ( n2756 , n7026 , n6809 );
    not g9037 ( n5840 , n10465 );
    nor g9038 ( n3156 , n10363 , n4693 );
    and g9039 ( n4042 , n6507 , n6276 );
    nor g9040 ( n8298 , n7605 , n11407 );
    and g9041 ( n6839 , n8250 , n4688 );
    or g9042 ( n2915 , n4898 , n5842 );
    not g9043 ( n13219 , n1984 );
    or g9044 ( n10662 , n8513 , n8979 );
    and g9045 ( n10541 , n13252 , n11301 );
    not g9046 ( n6498 , n8746 );
    or g9047 ( n5870 , n11438 , n10418 );
    or g9048 ( n6425 , n8476 , n1866 );
    or g9049 ( n6276 , n6263 , n10608 );
    or g9050 ( n1244 , n7003 , n6541 );
    or g9051 ( n2713 , n4828 , n7183 );
    and g9052 ( n4426 , n13078 , n12328 );
    and g9053 ( n8927 , n815 , n9022 );
    or g9054 ( n6259 , n3132 , n4927 );
    and g9055 ( n1173 , n9315 , n8736 );
    or g9056 ( n1446 , n5450 , n6105 );
    and g9057 ( n8010 , n8786 , n5465 );
    or g9058 ( n4688 , n13005 , n901 );
    or g9059 ( n913 , n9174 , n7860 );
    not g9060 ( n9375 , n4550 );
    and g9061 ( n9735 , n9811 , n7463 );
    nor g9062 ( n7746 , n12999 , n11678 );
    or g9063 ( n3840 , n11647 , n13405 );
    and g9064 ( n1487 , n406 , n11159 );
    not g9065 ( n8034 , n7322 );
    or g9066 ( n8724 , n13413 , n9108 );
    or g9067 ( n11717 , n10825 , n11768 );
    or g9068 ( n20 , n11739 , n260 );
    nor g9069 ( n5937 , n3907 , n2352 );
    not g9070 ( n6018 , n5001 );
    or g9071 ( n174 , n9529 , n2328 );
    and g9072 ( n391 , n2983 , n10320 );
    and g9073 ( n11781 , n2533 , n4980 );
    not g9074 ( n1639 , n10172 );
    not g9075 ( n14011 , n10485 );
    or g9076 ( n4208 , n6111 , n2152 );
    not g9077 ( n14063 , n2958 );
    and g9078 ( n13445 , n7852 , n8613 );
    and g9079 ( n12072 , n3565 , n11216 );
    and g9080 ( n2580 , n1452 , n1786 );
    or g9081 ( n3206 , n412 , n5105 );
    or g9082 ( n3618 , n13108 , n8499 );
    nor g9083 ( n2185 , n12075 , n12739 );
    or g9084 ( n5463 , n228 , n6164 );
    and g9085 ( n6305 , n10512 , n9611 );
    or g9086 ( n3298 , n9229 , n11684 );
    nor g9087 ( n3359 , n4913 , n4629 );
    and g9088 ( n14504 , n7961 , n10142 );
    not g9089 ( n13367 , n3361 );
    or g9090 ( n3243 , n3512 , n7770 );
    not g9091 ( n2367 , n10377 );
    or g9092 ( n2652 , n8714 , n10521 );
    and g9093 ( n5215 , n2533 , n12186 );
    or g9094 ( n12774 , n12295 , n8022 );
    and g9095 ( n8910 , n2177 , n1139 );
    nor g9096 ( n4330 , n11498 , n14485 );
    and g9097 ( n12041 , n14227 , n11429 );
    or g9098 ( n853 , n100 , n1333 );
    and g9099 ( n6926 , n10668 , n12182 );
    and g9100 ( n9933 , n3932 , n2072 );
    or g9101 ( n13230 , n10231 , n11902 );
    or g9102 ( n11714 , n5033 , n4172 );
    or g9103 ( n8506 , n820 , n10005 );
    or g9104 ( n13268 , n5977 , n8952 );
    nor g9105 ( n1121 , n13213 , n13097 );
    or g9106 ( n11850 , n7684 , n13911 );
    or g9107 ( n11830 , n12131 , n6187 );
    or g9108 ( n10729 , n12100 , n3829 );
    or g9109 ( n10275 , n10624 , n5939 );
    not g9110 ( n1812 , n6058 );
    nor g9111 ( n13104 , n4624 , n8352 );
    and g9112 ( n207 , n10134 , n6100 );
    or g9113 ( n1292 , n5570 , n9118 );
    not g9114 ( n3440 , n10380 );
    and g9115 ( n6836 , n333 , n8384 );
    and g9116 ( n1887 , n6649 , n3310 );
    or g9117 ( n13618 , n6857 , n8497 );
    and g9118 ( n6835 , n9015 , n8159 );
    or g9119 ( n8928 , n1356 , n9141 );
    and g9120 ( n2285 , n3932 , n4972 );
    or g9121 ( n9945 , n8582 , n7154 );
    and g9122 ( n6804 , n7929 , n11113 );
    and g9123 ( n13495 , n8789 , n4107 );
    and g9124 ( n8494 , n7677 , n11166 );
    or g9125 ( n7585 , n1741 , n11039 );
    nor g9126 ( n13358 , n3003 , n6404 );
    and g9127 ( n7942 , n5104 , n11249 );
    not g9128 ( n14227 , n11668 );
    and g9129 ( n8357 , n10310 , n6546 );
    or g9130 ( n7654 , n12543 , n1418 );
    nor g9131 ( n9700 , n4633 , n5748 );
    not g9132 ( n11097 , n13234 );
    or g9133 ( n5652 , n4340 , n5147 );
    or g9134 ( n10497 , n4267 , n10407 );
    nor g9135 ( n3321 , n13310 , n1552 );
    and g9136 ( n146 , n5899 , n5854 );
    nor g9137 ( n14290 , n6387 , n4831 );
    nor g9138 ( n6813 , n10400 , n11439 );
    or g9139 ( n13663 , n1669 , n5704 );
    and g9140 ( n14392 , n9726 , n10579 );
    and g9141 ( n5610 , n8427 , n4559 );
    not g9142 ( n4806 , n13447 );
    and g9143 ( n14444 , n1255 , n3729 );
    not g9144 ( n12086 , n4270 );
    or g9145 ( n8896 , n11231 , n5942 );
    or g9146 ( n3238 , n478 , n11848 );
    not g9147 ( n14091 , n1495 );
    nor g9148 ( n3719 , n3876 , n9365 );
    nor g9149 ( n3912 , n7739 , n10848 );
    or g9150 ( n11612 , n2949 , n12033 );
    and g9151 ( n3887 , n10330 , n530 );
    nor g9152 ( n13551 , n8701 , n8334 );
    and g9153 ( n1075 , n12990 , n1192 );
    not g9154 ( n10394 , n4465 );
    nor g9155 ( n4309 , n1686 , n8733 );
    and g9156 ( n6612 , n11220 , n3641 );
    or g9157 ( n3072 , n2877 , n12113 );
    or g9158 ( n311 , n10624 , n6920 );
    and g9159 ( n226 , n5252 , n8428 );
    or g9160 ( n7151 , n1223 , n2381 );
    and g9161 ( n5939 , n8697 , n3748 );
    not g9162 ( n1427 , n7346 );
    or g9163 ( n3884 , n9931 , n11817 );
    or g9164 ( n10232 , n8907 , n4895 );
    or g9165 ( n4416 , n2086 , n12612 );
    nor g9166 ( n1159 , n4924 , n8860 );
    or g9167 ( n10315 , n13130 , n9158 );
    not g9168 ( n4128 , n3046 );
    and g9169 ( n3059 , n13641 , n8871 );
    not g9170 ( n13078 , n13038 );
    and g9171 ( n6371 , n1427 , n7044 );
    or g9172 ( n6024 , n10808 , n9009 );
    or g9173 ( n9349 , n13016 , n5319 );
    nor g9174 ( n3734 , n6209 , n6755 );
    nor g9175 ( n10907 , n5977 , n3642 );
    or g9176 ( n9518 , n6046 , n10892 );
    not g9177 ( n163 , n12874 );
    not g9178 ( n13874 , n6903 );
    and g9179 ( n3453 , n12404 , n130 );
    and g9180 ( n14175 , n8043 , n10274 );
    nor g9181 ( n6583 , n3394 , n10597 );
    and g9182 ( n8930 , n12015 , n12266 );
    and g9183 ( n13545 , n12445 , n963 );
    or g9184 ( n9270 , n6849 , n3804 );
    not g9185 ( n13194 , n3367 );
    or g9186 ( n8616 , n10713 , n8719 );
    nor g9187 ( n7109 , n4313 , n6751 );
    nor g9188 ( n7606 , n4897 , n12955 );
    and g9189 ( n13105 , n1138 , n9669 );
    and g9190 ( n11266 , n11020 , n10026 );
    or g9191 ( n11827 , n9289 , n3131 );
    or g9192 ( n14262 , n390 , n9431 );
    and g9193 ( n13771 , n10556 , n4323 );
    not g9194 ( n6030 , n10406 );
    and g9195 ( n9576 , n2820 , n11203 );
    nor g9196 ( n1246 , n3333 , n10257 );
    or g9197 ( n5127 , n12357 , n666 );
    and g9198 ( n8317 , n5012 , n2015 );
    or g9199 ( n5496 , n10825 , n4297 );
    or g9200 ( n5788 , n7216 , n14293 );
    or g9201 ( n10536 , n7212 , n4157 );
    nor g9202 ( n5989 , n4417 , n2561 );
    and g9203 ( n3501 , n10330 , n9622 );
    not g9204 ( n100 , n9453 );
    nor g9205 ( n10776 , n12644 , n9963 );
    or g9206 ( n8274 , n11722 , n10212 );
    and g9207 ( n6418 , n8817 , n13862 );
    or g9208 ( n5017 , n13130 , n14098 );
    nor g9209 ( n1852 , n6731 , n3355 );
    or g9210 ( n9095 , n6111 , n767 );
    not g9211 ( n4484 , n760 );
    and g9212 ( n10513 , n12542 , n10221 );
    or g9213 ( n9752 , n12401 , n6942 );
    and g9214 ( n7738 , n7053 , n11567 );
    or g9215 ( n8316 , n13432 , n1069 );
    or g9216 ( n4531 , n14319 , n6496 );
    or g9217 ( n10009 , n11405 , n10901 );
    and g9218 ( n5616 , n2709 , n11868 );
    or g9219 ( n5809 , n5491 , n7917 );
    or g9220 ( n14403 , n2016 , n8732 );
    or g9221 ( n13887 , n7212 , n2536 );
    not g9222 ( n9119 , n5184 );
    not g9223 ( n3523 , n11227 );
    and g9224 ( n2156 , n2521 , n6257 );
    and g9225 ( n10888 , n9571 , n3756 );
    nor g9226 ( n12316 , n4549 , n11751 );
    or g9227 ( n13388 , n12353 , n2913 );
    or g9228 ( n13879 , n3025 , n3551 );
    or g9229 ( n7743 , n11105 , n6858 );
    or g9230 ( n4749 , n4988 , n8885 );
    or g9231 ( n9829 , n560 , n8486 );
    nor g9232 ( n5005 , n163 , n2446 );
    or g9233 ( n6773 , n1172 , n3830 );
    nor g9234 ( n9295 , n5990 , n14168 );
    and g9235 ( n5345 , n9191 , n7217 );
    nor g9236 ( n8178 , n5042 , n9639 );
    nor g9237 ( n13414 , n12522 , n2199 );
    nor g9238 ( n10114 , n13937 , n5810 );
    not g9239 ( n506 , n11412 );
    nor g9240 ( n7714 , n4342 , n987 );
    nor g9241 ( n4974 , n7362 , n2380 );
    or g9242 ( n6570 , n11576 , n10927 );
    or g9243 ( n3241 , n10534 , n3084 );
    and g9244 ( n12125 , n12730 , n13454 );
    and g9245 ( n3048 , n12039 , n8666 );
    and g9246 ( n8756 , n11163 , n12146 );
    and g9247 ( n10501 , n5053 , n9623 );
    not g9248 ( n11240 , n8424 );
    or g9249 ( n9121 , n4739 , n8009 );
    or g9250 ( n2042 , n8045 , n6371 );
    or g9251 ( n8862 , n5266 , n3256 );
    not g9252 ( n7717 , n1742 );
    and g9253 ( n6987 , n7429 , n2232 );
    nor g9254 ( n13569 , n1623 , n6841 );
    and g9255 ( n12656 , n4856 , n12645 );
    not g9256 ( n13041 , n7920 );
    nor g9257 ( n4610 , n12872 , n10495 );
    or g9258 ( n14144 , n3815 , n7168 );
    and g9259 ( n11200 , n6606 , n3119 );
    and g9260 ( n9402 , n10595 , n8403 );
    or g9261 ( n11100 , n14039 , n6791 );
    not g9262 ( n13155 , n6264 );
    nor g9263 ( n10401 , n1458 , n10746 );
    or g9264 ( n7878 , n6471 , n12457 );
    and g9265 ( n7870 , n678 , n14495 );
    or g9266 ( n8419 , n203 , n5184 );
    nor g9267 ( n9150 , n7418 , n9396 );
    and g9268 ( n12474 , n6531 , n559 );
    and g9269 ( n8258 , n1452 , n10666 );
    and g9270 ( n5261 , n6744 , n10438 );
    or g9271 ( n2511 , n1538 , n13444 );
    or g9272 ( n8962 , n1582 , n12195 );
    not g9273 ( n11809 , n4296 );
    not g9274 ( n11142 , n11861 );
    nor g9275 ( n933 , n8301 , n6515 );
    or g9276 ( n9832 , n6629 , n10419 );
    and g9277 ( n1871 , n10930 , n9992 );
    or g9278 ( n5774 , n4840 , n7598 );
    or g9279 ( n5322 , n14401 , n8508 );
    nor g9280 ( n4797 , n1685 , n13530 );
    and g9281 ( n6682 , n3506 , n1758 );
    or g9282 ( n13150 , n13854 , n9547 );
    or g9283 ( n12723 , n3062 , n5633 );
    not g9284 ( n4844 , n2692 );
    or g9285 ( n12306 , n4092 , n8872 );
    or g9286 ( n1181 , n13130 , n5688 );
    and g9287 ( n6624 , n10458 , n4130 );
    and g9288 ( n10137 , n13359 , n246 );
    and g9289 ( n723 , n6909 , n7816 );
    and g9290 ( n13331 , n4722 , n2049 );
    or g9291 ( n9729 , n974 , n11883 );
    and g9292 ( n4391 , n1414 , n11904 );
    or g9293 ( n13077 , n6596 , n13554 );
    and g9294 ( n908 , n8789 , n13372 );
    or g9295 ( n6390 , n8581 , n9989 );
    or g9296 ( n4339 , n11459 , n8083 );
    not g9297 ( n4098 , n304 );
    and g9298 ( n4029 , n11950 , n13818 );
    not g9299 ( n523 , n12776 );
    or g9300 ( n3080 , n3164 , n10835 );
    not g9301 ( n129 , n742 );
    or g9302 ( n9896 , n7527 , n13906 );
    or g9303 ( n10788 , n12712 , n431 );
    or g9304 ( n10994 , n5226 , n13625 );
    nor g9305 ( n4547 , n1623 , n10133 );
    or g9306 ( n9036 , n1535 , n8434 );
    and g9307 ( n12952 , n3785 , n305 );
    not g9308 ( n8816 , n7600 );
    and g9309 ( n1060 , n4341 , n6319 );
    and g9310 ( n4900 , n6316 , n3049 );
    and g9311 ( n9805 , n6527 , n7479 );
    or g9312 ( n12519 , n6706 , n631 );
    and g9313 ( n4903 , n129 , n9815 );
    or g9314 ( n10120 , n4199 , n336 );
    or g9315 ( n1965 , n1840 , n4958 );
    or g9316 ( n9585 , n9078 , n9727 );
    not g9317 ( n7691 , n5182 );
    and g9318 ( n3163 , n10457 , n8225 );
    not g9319 ( n7940 , n11401 );
    and g9320 ( n1533 , n3097 , n2629 );
    or g9321 ( n7537 , n647 , n3244 );
    or g9322 ( n14016 , n2012 , n6810 );
    and g9323 ( n2383 , n4373 , n6941 );
    and g9324 ( n13007 , n14109 , n13919 );
    or g9325 ( n12529 , n954 , n11141 );
    not g9326 ( n8650 , n5257 );
    or g9327 ( n8069 , n12351 , n4699 );
    or g9328 ( n144 , n6350 , n8519 );
    and g9329 ( n14180 , n9069 , n2992 );
    and g9330 ( n292 , n3672 , n12163 );
    nor g9331 ( n8180 , n9423 , n2726 );
    and g9332 ( n138 , n10457 , n3902 );
    not g9333 ( n3248 , n6806 );
    not g9334 ( n3394 , n13234 );
    or g9335 ( n3375 , n14472 , n8155 );
    not g9336 ( n14239 , n14510 );
    not g9337 ( n12593 , n9550 );
    and g9338 ( n13540 , n11495 , n13976 );
    or g9339 ( n13903 , n11438 , n6370 );
    or g9340 ( n13864 , n14110 , n1300 );
    and g9341 ( n13708 , n5628 , n9884 );
    nor g9342 ( n13260 , n12934 , n681 );
    not g9343 ( n5306 , n14367 );
    and g9344 ( n10985 , n1908 , n8750 );
    or g9345 ( n1296 , n2318 , n12474 );
    and g9346 ( n13031 , n10015 , n9349 );
    not g9347 ( n194 , n3357 );
    not g9348 ( n6486 , n1120 );
    or g9349 ( n8804 , n7364 , n4781 );
    not g9350 ( n2925 , n13944 );
    or g9351 ( n10805 , n7003 , n10613 );
    or g9352 ( n7298 , n2055 , n9443 );
    or g9353 ( n6603 , n11776 , n6873 );
    and g9354 ( n13444 , n7060 , n13864 );
    nor g9355 ( n5041 , n163 , n1126 );
    not g9356 ( n2188 , n9186 );
    and g9357 ( n13345 , n10595 , n11830 );
    or g9358 ( n5664 , n13035 , n9186 );
    nor g9359 ( n13844 , n6434 , n5400 );
    not g9360 ( n13700 , n6819 );
    and g9361 ( n10087 , n5475 , n12811 );
    and g9362 ( n3353 , n13147 , n5002 );
    and g9363 ( n5499 , n2486 , n8071 );
    and g9364 ( n10652 , n2564 , n1761 );
    nor g9365 ( n3325 , n1686 , n3658 );
    or g9366 ( n5089 , n10808 , n2636 );
    or g9367 ( n5846 , n12633 , n10693 );
    or g9368 ( n13004 , n13537 , n5730 );
    not g9369 ( n3742 , n12522 );
    and g9370 ( n288 , n501 , n14128 );
    or g9371 ( n11516 , n10035 , n4911 );
    or g9372 ( n14209 , n6654 , n5191 );
    and g9373 ( n426 , n5668 , n7546 );
    not g9374 ( n12101 , n7902 );
    and g9375 ( n5222 , n2758 , n13247 );
    or g9376 ( n252 , n9429 , n5744 );
    nor g9377 ( n5075 , n1028 , n1553 );
    or g9378 ( n7867 , n5007 , n5803 );
    or g9379 ( n13185 , n10300 , n14225 );
    or g9380 ( n845 , n12414 , n9939 );
    and g9381 ( n10183 , n327 , n14458 );
    or g9382 ( n1 , n2843 , n12864 );
    and g9383 ( n8845 , n5062 , n262 );
    and g9384 ( n10361 , n6130 , n9121 );
    and g9385 ( n4401 , n1247 , n11339 );
    or g9386 ( n7135 , n13547 , n6461 );
    not g9387 ( n5613 , n7258 );
    nor g9388 ( n8441 , n2919 , n10782 );
    not g9389 ( n4050 , n7931 );
    nor g9390 ( n10811 , n7551 , n1338 );
    nor g9391 ( n66 , n8887 , n9317 );
    and g9392 ( n10182 , n5940 , n5774 );
    and g9393 ( n11855 , n8213 , n7639 );
    and g9394 ( n676 , n9275 , n9575 );
    or g9395 ( n1419 , n1628 , n8099 );
    and g9396 ( n2026 , n5876 , n13113 );
    and g9397 ( n2027 , n4615 , n13980 );
    and g9398 ( n3969 , n13240 , n5721 );
    or g9399 ( n10409 , n5084 , n6014 );
    or g9400 ( n13825 , n387 , n8409 );
    or g9401 ( n7351 , n523 , n7747 );
    and g9402 ( n9772 , n2998 , n10301 );
    not g9403 ( n6135 , n7621 );
    or g9404 ( n6249 , n5891 , n9741 );
    and g9405 ( n2311 , n3804 , n7757 );
    and g9406 ( n6577 , n5348 , n8364 );
    not g9407 ( n13734 , n11347 );
    not g9408 ( n9078 , n4149 );
    or g9409 ( n6387 , n3833 , n6436 );
    or g9410 ( n2605 , n5144 , n12007 );
    not g9411 ( n11300 , n12697 );
    and g9412 ( n8739 , n7717 , n7665 );
    or g9413 ( n2882 , n10035 , n7480 );
    and g9414 ( n12217 , n10855 , n10348 );
    not g9415 ( n1178 , n11324 );
    or g9416 ( n4017 , n4562 , n2319 );
    or g9417 ( n5094 , n820 , n7379 );
    or g9418 ( n2249 , n11223 , n3712 );
    or g9419 ( n8911 , n14337 , n6805 );
    and g9420 ( n7531 , n4844 , n10978 );
    or g9421 ( n13039 , n12844 , n10501 );
    or g9422 ( n3228 , n930 , n13914 );
    not g9423 ( n9269 , n1010 );
    or g9424 ( n11104 , n7156 , n2071 );
    not g9425 ( n3569 , n8272 );
    or g9426 ( n10249 , n8096 , n1381 );
    or g9427 ( n4754 , n5641 , n8554 );
    or g9428 ( n6136 , n3667 , n1753 );
    not g9429 ( n6388 , n8635 );
    and g9430 ( n7747 , n6830 , n408 );
    or g9431 ( n8914 , n13516 , n5511 );
    nor g9432 ( n9065 , n9871 , n13566 );
    or g9433 ( n7635 , n4908 , n3548 );
    nor g9434 ( n9653 , n3905 , n1733 );
    not g9435 ( n6316 , n3926 );
    not g9436 ( n11213 , n6426 );
    not g9437 ( n12772 , n5944 );
    and g9438 ( n5231 , n12615 , n6178 );
    or g9439 ( n12095 , n648 , n6401 );
    or g9440 ( n12117 , n7282 , n13944 );
    or g9441 ( n938 , n9230 , n10150 );
    and g9442 ( n11089 , n12721 , n6140 );
    and g9443 ( n9963 , n13236 , n11573 );
    or g9444 ( n461 , n1203 , n10426 );
    not g9445 ( n2521 , n6193 );
    and g9446 ( n9980 , n678 , n13285 );
    and g9447 ( n12973 , n12449 , n8031 );
    or g9448 ( n11429 , n647 , n8683 );
    and g9449 ( n9292 , n13362 , n12540 );
    not g9450 ( n2727 , n9041 );
    and g9451 ( n195 , n9188 , n7304 );
    or g9452 ( n4023 , n7700 , n8136 );
    not g9453 ( n6556 , n9555 );
    and g9454 ( n13286 , n8431 , n12148 );
    or g9455 ( n6466 , n13364 , n2061 );
    and g9456 ( n2305 , n3276 , n1901 );
    or g9457 ( n13285 , n9111 , n13678 );
    or g9458 ( n173 , n5861 , n4709 );
    and g9459 ( n3913 , n10678 , n14329 );
    or g9460 ( n2592 , n3193 , n9500 );
    not g9461 ( n12866 , n8822 );
    and g9462 ( n2160 , n3672 , n6669 );
    not g9463 ( n2790 , n14354 );
    or g9464 ( n11244 , n13194 , n9543 );
    nor g9465 ( n5058 , n11285 , n1403 );
    and g9466 ( n5519 , n12105 , n10981 );
    or g9467 ( n13475 , n5266 , n3691 );
    or g9468 ( n10533 , n6730 , n9627 );
    and g9469 ( n3084 , n7081 , n1891 );
    or g9470 ( n6156 , n185 , n4783 );
    and g9471 ( n10636 , n14351 , n9057 );
    and g9472 ( n12234 , n11737 , n12984 );
    or g9473 ( n13686 , n387 , n7587 );
    or g9474 ( n12811 , n7426 , n12752 );
    not g9475 ( n13270 , n4561 );
    and g9476 ( n8989 , n8386 , n3791 );
    and g9477 ( n7259 , n11020 , n9974 );
    nor g9478 ( n8126 , n12765 , n12388 );
    and g9479 ( n7424 , n2310 , n11358 );
    or g9480 ( n3623 , n13132 , n5960 );
    or g9481 ( n5211 , n4828 , n4779 );
    and g9482 ( n64 , n1678 , n12971 );
    or g9483 ( n10389 , n49 , n8176 );
    or g9484 ( n4827 , n8897 , n14191 );
    and g9485 ( n570 , n10247 , n3080 );
    and g9486 ( n3349 , n13362 , n9327 );
    or g9487 ( n6514 , n11440 , n6910 );
    or g9488 ( n11091 , n4407 , n5261 );
    or g9489 ( n9626 , n839 , n10947 );
    and g9490 ( n9016 , n2021 , n10493 );
    nor g9491 ( n1293 , n13154 , n3716 );
    and g9492 ( n9900 , n12404 , n1483 );
    and g9493 ( n13040 , n225 , n2599 );
    or g9494 ( n13713 , n8575 , n10468 );
    and g9495 ( n1324 , n9323 , n10161 );
    and g9496 ( n8611 , n8950 , n1285 );
    and g9497 ( n42 , n3268 , n1873 );
    or g9498 ( n5808 , n3871 , n6782 );
    and g9499 ( n6806 , n11824 , n1447 );
    and g9500 ( n10129 , n6606 , n6648 );
    not g9501 ( n2099 , n8008 );
    and g9502 ( n11618 , n12475 , n9802 );
    and g9503 ( n13987 , n9726 , n8542 );
    not g9504 ( n13557 , n670 );
    or g9505 ( n8202 , n2877 , n13212 );
    and g9506 ( n10902 , n14109 , n2945 );
    or g9507 ( n4726 , n1711 , n2382 );
    or g9508 ( n11700 , n14400 , n14261 );
    not g9509 ( n14075 , n4324 );
    and g9510 ( n8447 , n200 , n5775 );
    or g9511 ( n11188 , n3364 , n6007 );
    not g9512 ( n1223 , n1676 );
    not g9513 ( n4207 , n2130 );
    not g9514 ( n4210 , n8809 );
    or g9515 ( n5096 , n9442 , n5765 );
    or g9516 ( n11845 , n3320 , n13529 );
    not g9517 ( n12576 , n11415 );
    and g9518 ( n472 , n13379 , n7240 );
    and g9519 ( n9661 , n3276 , n8623 );
    not g9520 ( n8277 , n14412 );
    or g9521 ( n13974 , n7462 , n914 );
    and g9522 ( n8755 , n12185 , n7591 );
    not g9523 ( n3019 , n6196 );
    or g9524 ( n2259 , n1147 , n10557 );
    nor g9525 ( n360 , n12107 , n11745 );
    not g9526 ( n2766 , n5668 );
    and g9527 ( n11377 , n9890 , n14056 );
    and g9528 ( n11556 , n8692 , n11629 );
    or g9529 ( n14013 , n14088 , n9241 );
    or g9530 ( n8722 , n13485 , n5598 );
    and g9531 ( n1585 , n11950 , n9449 );
    nor g9532 ( n12220 , n14106 , n11050 );
    and g9533 ( n9809 , n9705 , n1448 );
    or g9534 ( n1080 , n6690 , n5538 );
    or g9535 ( n6173 , n7888 , n5423 );
    or g9536 ( n73 , n1697 , n5371 );
    or g9537 ( n5158 , n4162 , n9254 );
    and g9538 ( n9385 , n10566 , n11880 );
    not g9539 ( n7392 , n300 );
    or g9540 ( n23 , n3826 , n10851 );
    and g9541 ( n2135 , n432 , n4020 );
    and g9542 ( n1736 , n2281 , n10786 );
    and g9543 ( n10028 , n7691 , n5996 );
    nor g9544 ( n374 , n7229 , n9380 );
    not g9545 ( n12823 , n736 );
    not g9546 ( n10715 , n13779 );
    or g9547 ( n9597 , n10731 , n11943 );
    and g9548 ( n5308 , n1662 , n14176 );
    or g9549 ( n2960 , n4255 , n11099 );
    or g9550 ( n1317 , n10534 , n662 );
    or g9551 ( n6112 , n2761 , n12938 );
    not g9552 ( n3871 , n4891 );
    or g9553 ( n13617 , n2645 , n7147 );
    or g9554 ( n10384 , n1920 , n7104 );
    and g9555 ( n11888 , n3097 , n3318 );
    or g9556 ( n11787 , n13130 , n253 );
    and g9557 ( n1049 , n13338 , n6328 );
    nor g9558 ( n11662 , n8404 , n75 );
    and g9559 ( n3324 , n11688 , n6268 );
    and g9560 ( n24 , n9705 , n1442 );
    or g9561 ( n895 , n7227 , n12605 );
    and g9562 ( n2569 , n1428 , n12981 );
    or g9563 ( n369 , n2179 , n2725 );
    not g9564 ( n7961 , n7808 );
    or g9565 ( n840 , n10461 , n6310 );
    or g9566 ( n657 , n1820 , n10020 );
    or g9567 ( n3625 , n9541 , n90 );
    and g9568 ( n8279 , n1266 , n7118 );
    and g9569 ( n14141 , n8386 , n11478 );
    and g9570 ( n11270 , n8232 , n6681 );
    or g9571 ( n10246 , n11223 , n14356 );
    or g9572 ( n11989 , n11303 , n13749 );
    nor g9573 ( n4259 , n12568 , n1524 );
    and g9574 ( n11599 , n6192 , n12050 );
    or g9575 ( n8226 , n12414 , n319 );
    and g9576 ( n10515 , n4154 , n1180 );
    or g9577 ( n6620 , n7358 , n1018 );
    nor g9578 ( n4035 , n11761 , n1297 );
    and g9579 ( n10436 , n4347 , n12671 );
    or g9580 ( n12419 , n12428 , n5356 );
    not g9581 ( n3914 , n1214 );
    not g9582 ( n2473 , n10803 );
    or g9583 ( n910 , n1875 , n11092 );
    nor g9584 ( n14285 , n13350 , n8729 );
    or g9585 ( n7178 , n8458 , n7233 );
    not g9586 ( n6957 , n6139 );
    and g9587 ( n10078 , n5628 , n8831 );
    or g9588 ( n12997 , n2888 , n2855 );
    nor g9589 ( n9400 , n8277 , n5396 );
    and g9590 ( n4040 , n8238 , n2290 );
    and g9591 ( n1272 , n13781 , n7447 );
    or g9592 ( n11373 , n13108 , n2859 );
    or g9593 ( n6886 , n11176 , n6698 );
    or g9594 ( n13123 , n9429 , n539 );
    and g9595 ( n3703 , n10399 , n4370 );
    or g9596 ( n9610 , n1914 , n2950 );
    and g9597 ( n10635 , n14145 , n5258 );
    and g9598 ( n14055 , n14446 , n12777 );
    or g9599 ( n1940 , n11576 , n6445 );
    or g9600 ( n5498 , n6039 , n3733 );
    and g9601 ( n3331 , n10619 , n4419 );
    nor g9602 ( n14136 , n5418 , n6643 );
    or g9603 ( n12078 , n6323 , n10397 );
    and g9604 ( n5196 , n13867 , n4515 );
    and g9605 ( n13556 , n6525 , n716 );
    or g9606 ( n175 , n9507 , n11931 );
    nor g9607 ( n13964 , n1838 , n4363 );
    or g9608 ( n8525 , n4481 , n3980 );
    or g9609 ( n13156 , n8881 , n13253 );
    or g9610 ( n12567 , n11105 , n2243 );
    and g9611 ( n10894 , n873 , n10561 );
    not g9612 ( n6883 , n3094 );
    or g9613 ( n6581 , n14466 , n13221 );
    nor g9614 ( n3414 , n7551 , n299 );
    not g9615 ( n10457 , n7802 );
    nor g9616 ( n5057 , n882 , n12198 );
    and g9617 ( n12514 , n7673 , n10798 );
    or g9618 ( n6635 , n361 , n289 );
    nor g9619 ( n9683 , n10121 , n12755 );
    not g9620 ( n8855 , n13190 );
    and g9621 ( n10743 , n9275 , n12068 );
    not g9622 ( n5591 , n10278 );
    or g9623 ( n10827 , n9507 , n2100 );
    or g9624 ( n3396 , n1198 , n2190 );
    and g9625 ( n6993 , n13338 , n9054 );
    and g9626 ( n12867 , n3405 , n4530 );
    or g9627 ( n2894 , n89 , n5162 );
    and g9628 ( n5326 , n10705 , n3138 );
    or g9629 ( n8245 , n9078 , n12507 );
    nor g9630 ( n3863 , n12568 , n3779 );
    and g9631 ( n9045 , n7911 , n3096 );
    or g9632 ( n10282 , n7502 , n6758 );
    and g9633 ( n14330 , n5725 , n2856 );
    and g9634 ( n2134 , n7691 , n13517 );
    or g9635 ( n11118 , n1044 , n604 );
    not g9636 ( n6243 , n2566 );
    nor g9637 ( n7210 , n11633 , n13207 );
    or g9638 ( n5397 , n9218 , n7134 );
    nor g9639 ( n685 , n8959 , n7865 );
    and g9640 ( n3535 , n9745 , n5072 );
    and g9641 ( n10752 , n10710 , n10886 );
    not g9642 ( n6807 , n11441 );
    nor g9643 ( n14236 , n5569 , n3338 );
    or g9644 ( n9574 , n12994 , n2831 );
    and g9645 ( n11235 , n3565 , n1279 );
    nor g9646 ( n3308 , n1023 , n13471 );
    not g9647 ( n9052 , n1086 );
    nor g9648 ( n13816 , n8458 , n5170 );
    or g9649 ( n3891 , n5180 , n8402 );
    not g9650 ( n13991 , n11813 );
    or g9651 ( n10640 , n1613 , n714 );
    and g9652 ( n4060 , n13850 , n12156 );
    or g9653 ( n3112 , n1112 , n7928 );
    and g9654 ( n13001 , n11142 , n11717 );
    or g9655 ( n11458 , n11315 , n14507 );
    or g9656 ( n7350 , n3888 , n6511 );
    and g9657 ( n13546 , n11403 , n2630 );
    and g9658 ( n9410 , n7826 , n13746 );
    and g9659 ( n2751 , n4422 , n6291 );
    not g9660 ( n1061 , n9959 );
    nor g9661 ( n1530 , n8209 , n9631 );
    or g9662 ( n6792 , n12844 , n3862 );
    or g9663 ( n9114 , n8404 , n3502 );
    not g9664 ( n839 , n2794 );
    nor g9665 ( n13528 , n7227 , n4636 );
    nor g9666 ( n9147 , n1548 , n2193 );
    and g9667 ( n10901 , n200 , n4360 );
    or g9668 ( n12793 , n12764 , n14306 );
    nor g9669 ( n7252 , n3418 , n3033 );
    and g9670 ( n11441 , n9245 , n356 );
    and g9671 ( n1082 , n2330 , n724 );
    and g9672 ( n12564 , n2587 , n10639 );
    nor g9673 ( n1859 , n12193 , n4366 );
    or g9674 ( n1416 , n4207 , n1309 );
    and g9675 ( n5600 , n8769 , n12478 );
    not g9676 ( n185 , n4149 );
    or g9677 ( n14049 , n7862 , n4400 );
    or g9678 ( n2989 , n5641 , n5280 );
    and g9679 ( n485 , n14446 , n6692 );
    or g9680 ( n7528 , n14472 , n3362 );
    not g9681 ( n6953 , n1312 );
    or g9682 ( n4564 , n13650 , n8044 );
    nor g9683 ( n6964 , n14166 , n6221 );
    or g9684 ( n12595 , n12549 , n7896 );
    or g9685 ( n1421 , n3820 , n674 );
    and g9686 ( n3834 , n9650 , n13430 );
    and g9687 ( n3063 , n11093 , n1537 );
    and g9688 ( n10861 , n2760 , n2717 );
    or g9689 ( n3230 , n6680 , n3804 );
    nor g9690 ( n11898 , n5468 , n3774 );
    or g9691 ( n14519 , n850 , n8092 );
    and g9692 ( n13876 , n8183 , n12950 );
    and g9693 ( n9625 , n13555 , n13229 );
    not g9694 ( n10302 , n1120 );
    or g9695 ( n2168 , n14319 , n8770 );
    not g9696 ( n5391 , n2369 );
    nor g9697 ( n13603 , n10620 , n8443 );
    nor g9698 ( n1524 , n13072 , n12433 );
    not g9699 ( n4104 , n6397 );
    or g9700 ( n1097 , n492 , n6955 );
    and g9701 ( n4240 , n904 , n8819 );
    and g9702 ( n3266 , n55 , n1555 );
    or g9703 ( n4150 , n10300 , n1601 );
    and g9704 ( n8853 , n12389 , n10004 );
    and g9705 ( n3294 , n9265 , n6299 );
    and g9706 ( n13176 , n3923 , n4319 );
    or g9707 ( n4338 , n3768 , n1897 );
    or g9708 ( n1068 , n7364 , n4611 );
    and g9709 ( n7042 , n2820 , n10500 );
    and g9710 ( n3391 , n1857 , n2621 );
    and g9711 ( n6370 , n2322 , n3825 );
    and g9712 ( n13141 , n4147 , n14096 );
    nor g9713 ( n8876 , n393 , n10880 );
    or g9714 ( n13747 , n3025 , n5101 );
    or g9715 ( n372 , n13446 , n8708 );
    or g9716 ( n7676 , n8655 , n11143 );
    or g9717 ( n7367 , n13885 , n786 );
    or g9718 ( n4526 , n1061 , n2907 );
    nor g9719 ( n11767 , n5172 , n6290 );
    not g9720 ( n3449 , n11902 );
    or g9721 ( n3748 , n8828 , n7394 );
    or g9722 ( n6767 , n11176 , n10193 );
    and g9723 ( n11602 , n7427 , n12798 );
    or g9724 ( n3128 , n8242 , n6762 );
    and g9725 ( n1688 , n9824 , n1477 );
    and g9726 ( n12617 , n1140 , n435 );
    nor g9727 ( n7775 , n2171 , n2396 );
    and g9728 ( n5581 , n11607 , n218 );
    or g9729 ( n301 , n480 , n7906 );
    or g9730 ( n9274 , n550 , n9544 );
    or g9731 ( n5745 , n3877 , n1009 );
    and g9732 ( n13101 , n11153 , n5935 );
    and g9733 ( n4122 , n7284 , n12227 );
    and g9734 ( n2715 , n11816 , n2933 );
    or g9735 ( n3739 , n8096 , n2184 );
    not g9736 ( n12580 , n5990 );
    not g9737 ( n3820 , n3910 );
    and g9738 ( n5490 , n6527 , n2079 );
    or g9739 ( n4770 , n6271 , n17 );
    and g9740 ( n10792 , n6753 , n13491 );
    or g9741 ( n6908 , n568 , n11991 );
    not g9742 ( n2103 , n7929 );
    and g9743 ( n10157 , n5574 , n5228 );
    and g9744 ( n6602 , n3743 , n7097 );
    and g9745 ( n11289 , n10854 , n8990 );
    nor g9746 ( n3639 , n478 , n2707 );
    nor g9747 ( n5015 , n14332 , n13826 );
    or g9748 ( n2293 , n13413 , n12282 );
    not g9749 ( n9967 , n11264 );
    and g9750 ( n6578 , n13780 , n13982 );
    or g9751 ( n10586 , n8983 , n5750 );
    nor g9752 ( n7742 , n2875 , n3226 );
    not g9753 ( n7660 , n4991 );
    not g9754 ( n7364 , n7086 );
    or g9755 ( n4100 , n10808 , n2444 );
    nor g9756 ( n4142 , n14370 , n13945 );
    or g9757 ( n6992 , n11459 , n9495 );
    not g9758 ( n13432 , n8595 );
    and g9759 ( n9985 , n2760 , n612 );
    or g9760 ( n1988 , n10637 , n8218 );
    and g9761 ( n1467 , n718 , n14397 );
    and g9762 ( n2070 , n8232 , n4202 );
    and g9763 ( n12598 , n2461 , n3805 );
    nor g9764 ( n7422 , n7023 , n1004 );
    or g9765 ( n11821 , n5253 , n10484 );
    and g9766 ( n6882 , n11313 , n8456 );
    and g9767 ( n918 , n9677 , n2269 );
    or g9768 ( n3253 , n2562 , n1726 );
    or g9769 ( n3172 , n2857 , n11501 );
    nor g9770 ( n5289 , n12872 , n10263 );
    not g9771 ( n7407 , n14461 );
    nor g9772 ( n13389 , n2799 , n12431 );
    and g9773 ( n2277 , n11316 , n8536 );
    not g9774 ( n13518 , n10775 );
    nor g9775 ( n4523 , n2236 , n7580 );
    or g9776 ( n6022 , n10310 , n2061 );
    or g9777 ( n3671 , n14319 , n4312 );
    or g9778 ( n6093 , n14400 , n11536 );
    and g9779 ( n864 , n13107 , n11238 );
    and g9780 ( n4279 , n10736 , n10921 );
    nor g9781 ( n12275 , n1342 , n858 );
    or g9782 ( n4258 , n2925 , n7941 );
    and g9783 ( n11296 , n5012 , n4787 );
    not g9784 ( n2251 , n9829 );
    or g9785 ( n13454 , n1741 , n6851 );
    and g9786 ( n13956 , n11422 , n8460 );
    or g9787 ( n12146 , n2747 , n6658 );
    not g9788 ( n2451 , n7223 );
    and g9789 ( n7106 , n12721 , n11638 );
    not g9790 ( n6424 , n11654 );
    or g9791 ( n11640 , n13991 , n6492 );
    nor g9792 ( n10653 , n4195 , n3676 );
    not g9793 ( n7943 , n4589 );
    nor g9794 ( n7105 , n2405 , n9779 );
    not g9795 ( n1575 , n5690 );
    or g9796 ( n10510 , n14110 , n155 );
    and g9797 ( n2582 , n14260 , n8234 );
    and g9798 ( n2971 , n4856 , n134 );
    not g9799 ( n10269 , n10219 );
    nor g9800 ( n6349 , n7809 , n10353 );
    or g9801 ( n7948 , n2747 , n7993 );
    or g9802 ( n29 , n8404 , n10097 );
    or g9803 ( n3661 , n12023 , n11144 );
    or g9804 ( n4780 , n227 , n14447 );
    nor g9805 ( n8257 , n1480 , n8249 );
    and g9806 ( n11721 , n12421 , n561 );
    and g9807 ( n2596 , n4261 , n711 );
    nor g9808 ( n2707 , n3521 , n6374 );
    and g9809 ( n2365 , n1266 , n6961 );
    or g9810 ( n9247 , n5144 , n3896 );
    nor g9811 ( n13688 , n8353 , n6584 );
    and g9812 ( n5457 , n4276 , n8506 );
    or g9813 ( n10 , n9423 , n7263 );
    and g9814 ( n8952 , n13952 , n12505 );
    and g9815 ( n12299 , n6243 , n4600 );
    or g9816 ( n13336 , n3076 , n10937 );
    and g9817 ( n10371 , n12018 , n5836 );
    not g9818 ( n9228 , n8552 );
    and g9819 ( n11055 , n5683 , n1985 );
    and g9820 ( n6174 , n1193 , n540 );
    and g9821 ( n6472 , n1193 , n11179 );
    or g9822 ( n14421 , n10191 , n8303 );
    or g9823 ( n10995 , n2057 , n2598 );
    or g9824 ( n1420 , n11647 , n5623 );
    and g9825 ( n8493 , n2021 , n9821 );
    or g9826 ( n10016 , n12324 , n4603 );
    and g9827 ( n9989 , n11411 , n8957 );
    and g9828 ( n3117 , n1074 , n14182 );
    not g9829 ( n11422 , n13360 );
    or g9830 ( n8889 , n4340 , n8444 );
    and g9831 ( n5439 , n7745 , n11057 );
    nor g9832 ( n8231 , n2946 , n11485 );
    and g9833 ( n10279 , n1452 , n14498 );
    not g9834 ( n13276 , n1966 );
    or g9835 ( n3791 , n12934 , n1235 );
    and g9836 ( n9648 , n11748 , n1609 );
    and g9837 ( n4550 , n12102 , n12533 );
    or g9838 ( n13366 , n1701 , n9418 );
    nor g9839 ( n8633 , n8015 , n13387 );
    or g9840 ( n7330 , n1669 , n5485 );
    or g9841 ( n2423 , n9807 , n9834 );
    or g9842 ( n3057 , n3815 , n2912 );
    and g9843 ( n9279 , n12250 , n3722 );
    and g9844 ( n11132 , n79 , n6504 );
    and g9845 ( n3039 , n11336 , n12632 );
    not g9846 ( n4346 , n13908 );
    not g9847 ( n2064 , n261 );
    or g9848 ( n9366 , n1582 , n9332 );
    nor g9849 ( n8153 , n4207 , n5343 );
    nor g9850 ( n10006 , n2057 , n344 );
    nor g9851 ( n6345 , n1623 , n2733 );
    and g9852 ( n6853 , n11345 , n4580 );
    and g9853 ( n1374 , n3743 , n779 );
    or g9854 ( n248 , n2878 , n9739 );
    or g9855 ( n3469 , n4967 , n2008 );
    not g9856 ( n2158 , n1911 );
    not g9857 ( n8908 , n2970 );
    or g9858 ( n10583 , n3914 , n11712 );
    not g9859 ( n4313 , n4720 );
    or g9860 ( n10472 , n5409 , n4681 );
    and g9861 ( n7092 , n5999 , n12066 );
    and g9862 ( n4831 , n11117 , n13390 );
    not g9863 ( n8828 , n2130 );
    not g9864 ( n12391 , n5430 );
    and g9865 ( n4812 , n11838 , n6120 );
    and g9866 ( n378 , n2643 , n13830 );
    not g9867 ( n286 , n82 );
    and g9868 ( n2071 , n6724 , n2346 );
    and g9869 ( n4858 , n3652 , n9683 );
    and g9870 ( n6087 , n3449 , n6162 );
    and g9871 ( n4612 , n986 , n6605 );
    and g9872 ( n8903 , n1059 , n1765 );
    or g9873 ( n13187 , n10331 , n1619 );
    not g9874 ( n10318 , n3442 );
    or g9875 ( n12880 , n4821 , n10124 );
    or g9876 ( n3087 , n14435 , n12174 );
    or g9877 ( n10393 , n8172 , n10642 );
    and g9878 ( n10152 , n13342 , n11189 );
    and g9879 ( n11201 , n3365 , n4497 );
    or g9880 ( n11454 , n11011 , n2227 );
    and g9881 ( n11387 , n12229 , n2217 );
    or g9882 ( n5554 , n11621 , n6118 );
    or g9883 ( n12536 , n8821 , n13024 );
    nor g9884 ( n10859 , n11508 , n4607 );
    and g9885 ( n6597 , n446 , n2293 );
    and g9886 ( n810 , n11008 , n4171 );
    and g9887 ( n33 , n2985 , n3484 );
    or g9888 ( n11970 , n2412 , n10268 );
    not g9889 ( n9136 , n8049 );
    and g9890 ( n6858 , n10506 , n11402 );
    and g9891 ( n12583 , n11020 , n13210 );
    nor g9892 ( n8368 , n10730 , n374 );
    or g9893 ( n625 , n6695 , n9474 );
    or g9894 ( n8864 , n12601 , n4321 );
    and g9895 ( n12348 , n11737 , n8347 );
    not g9896 ( n7502 , n4147 );
    or g9897 ( n3727 , n6205 , n14389 );
    and g9898 ( n5544 , n2461 , n8255 );
    or g9899 ( n12753 , n13155 , n5394 );
    not g9900 ( n3003 , n11582 );
    and g9901 ( n6639 , n11803 , n11373 );
    or g9902 ( n11229 , n11935 , n146 );
    or g9903 ( n1912 , n14370 , n8135 );
    and g9904 ( n2418 , n8232 , n9746 );
    or g9905 ( n1105 , n8575 , n12809 );
    not g9906 ( n5182 , n12925 );
    or g9907 ( n8558 , n11420 , n710 );
    or g9908 ( n5444 , n12100 , n10008 );
    or g9909 ( n9367 , n3161 , n11507 );
    not g9910 ( n4276 , n13360 );
    nor g9911 ( n2488 , n11832 , n9100 );
    or g9912 ( n6219 , n361 , n3274 );
    and g9913 ( n5399 , n2527 , n133 );
    or g9914 ( n11107 , n1576 , n8515 );
    and g9915 ( n6771 , n5088 , n8526 );
    and g9916 ( n9559 , n7745 , n14187 );
    or g9917 ( n10139 , n1875 , n9242 );
    nor g9918 ( n11903 , n5986 , n1101 );
    nor g9919 ( n6386 , n1577 , n10627 );
    and g9920 ( n9534 , n12986 , n13742 );
    and g9921 ( n1145 , n2281 , n7113 );
    or g9922 ( n4220 , n3011 , n4811 );
    or g9923 ( n3636 , n2025 , n10311 );
    or g9924 ( n1921 , n2888 , n11992 );
    or g9925 ( n8610 , n7888 , n12973 );
    nor g9926 ( n4252 , n7919 , n3158 );
    and g9927 ( n8235 , n3755 , n3759 );
    not g9928 ( n2000 , n481 );
    not g9929 ( n5918 , n2405 );
    nor g9930 ( n6072 , n14239 , n13807 );
    not g9931 ( n8849 , n8168 );
    nor g9932 ( n3964 , n6018 , n8880 );
    or g9933 ( n7549 , n8980 , n5203 );
    or g9934 ( n8254 , n14319 , n13203 );
    or g9935 ( n5929 , n1669 , n8052 );
    not g9936 ( n5509 , n1780 );
    or g9937 ( n10747 , n10245 , n5934 );
    nor g9938 ( n1611 , n1112 , n5057 );
    or g9939 ( n6406 , n116 , n10199 );
    or g9940 ( n4061 , n817 , n8067 );
    and g9941 ( n5981 , n5137 , n1080 );
    not g9942 ( n5104 , n1812 );
    or g9943 ( n7492 , n695 , n8322 );
    and g9944 ( n11230 , n8923 , n917 );
    and g9945 ( n1269 , n14091 , n10017 );
    and g9946 ( n8188 , n8247 , n2063 );
    and g9947 ( n1563 , n1427 , n13156 );
    or g9948 ( n13666 , n4199 , n326 );
    or g9949 ( n463 , n11935 , n8097 );
    or g9950 ( n7416 , n1576 , n12847 );
    and g9951 ( n9723 , n7211 , n2508 );
    and g9952 ( n868 , n13359 , n13312 );
    and g9953 ( n2911 , n4525 , n712 );
    and g9954 ( n11080 , n986 , n7996 );
    and g9955 ( n9372 , n9494 , n2357 );
    or g9956 ( n11985 , n4435 , n6926 );
    or g9957 ( n9633 , n4602 , n9355 );
    or g9958 ( n4211 , n7912 , n6038 );
    not g9959 ( n10917 , n10036 );
    not g9960 ( n9931 , n13165 );
    and g9961 ( n13866 , n1788 , n7434 );
    or g9962 ( n8985 , n10024 , n4277 );
    and g9963 ( n7454 , n6354 , n8891 );
    or g9964 ( n5668 , n400 , n8073 );
    or g9965 ( n12518 , n820 , n7090 );
    not g9966 ( n12311 , n11515 );
    or g9967 ( n2066 , n5861 , n6380 );
    and g9968 ( n642 , n2998 , n11045 );
    nor g9969 ( n3285 , n7418 , n3816 );
    and g9970 ( n5193 , n783 , n3213 );
    not g9971 ( n34 , n7466 );
    not g9972 ( n4624 , n8291 );
    and g9973 ( n14399 , n10765 , n13916 );
    and g9974 ( n1779 , n4973 , n11134 );
    not g9975 ( n1059 , n12009 );
    and g9976 ( n13730 , n11674 , n7935 );
    and g9977 ( n12932 , n14074 , n11726 );
    or g9978 ( n5487 , n9289 , n5947 );
    and g9979 ( n6002 , n13575 , n5093 );
    and g9980 ( n8776 , n5038 , n13129 );
    or g9981 ( n9485 , n12625 , n1461 );
    nor g9982 ( n2395 , n14419 , n10459 );
    or g9983 ( n7169 , n4923 , n7983 );
    nor g9984 ( n11088 , n10318 , n13075 );
    and g9985 ( n1018 , n11748 , n1983 );
    not g9986 ( n9315 , n8122 );
    and g9987 ( n4591 , n2310 , n7491 );
    or g9988 ( n9503 , n228 , n47 );
    nor g9989 ( n6047 , n7023 , n12447 );
    and g9990 ( n591 , n8630 , n2408 );
    and g9991 ( n7086 , n9182 , n14060 );
    nor g9992 ( n9307 , n4299 , n7475 );
    nor g9993 ( n1101 , n6052 , n5361 );
    and g9994 ( n7819 , n1053 , n13298 );
    or g9995 ( n5036 , n3888 , n3173 );
    and g9996 ( n10416 , n1138 , n7522 );
    and g9997 ( n3334 , n3028 , n9894 );
    nor g9998 ( n5142 , n2194 , n795 );
    or g9999 ( n8050 , n9230 , n1215 );
    or g10000 ( n6391 , n5986 , n4080 );
    not g10001 ( n3193 , n11055 );
    and g10002 ( n10905 , n13147 , n14077 );
    not g10003 ( n4195 , n7064 );
    not g10004 ( n10458 , n12697 );
    or g10005 ( n14509 , n8908 , n5277 );
    not g10006 ( n3364 , n271 );
    or g10007 ( n4274 , n10539 , n6234 );
    nor g10008 ( n11277 , n228 , n5536 );
    or g10009 ( n3460 , n511 , n6025 );
    or g10010 ( n14187 , n1628 , n5375 );
    or g10011 ( n8338 , n4313 , n8611 );
    or g10012 ( n1578 , n10834 , n1797 );
    or g10013 ( n7535 , n9403 , n6945 );
    and g10014 ( n5116 , n13700 , n10974 );
    not g10015 ( n7255 , n7354 );
    not g10016 ( n13362 , n7802 );
    and g10017 ( n4379 , n4447 , n8901 );
    and g10018 ( n10679 , n2985 , n8651 );
    not g10019 ( n7484 , n14072 );
    not g10020 ( n5504 , n210 );
    nor g10021 ( n3446 , n9567 , n12396 );
    and g10022 ( n9316 , n10562 , n1359 );
    and g10023 ( n11311 , n6507 , n10253 );
    or g10024 ( n7304 , n412 , n12836 );
    or g10025 ( n8071 , n568 , n9417 );
    and g10026 ( n4376 , n7826 , n8998 );
    not g10027 ( n2942 , n13447 );
    or g10028 ( n14155 , n11472 , n11433 );
    and g10029 ( n7879 , n815 , n1013 );
    nor g10030 ( n3171 , n7359 , n7946 );
    or g10031 ( n13022 , n8881 , n7967 );
    and g10032 ( n7293 , n2985 , n5888 );
    not g10033 ( n3846 , n4266 );
    nor g10034 ( n13945 , n14011 , n8882 );
    and g10035 ( n3447 , n13379 , n7337 );
    and g10036 ( n9451 , n8801 , n1768 );
    or g10037 ( n12205 , n11739 , n4737 );
    not g10038 ( n13005 , n2320 );
    or g10039 ( n1104 , n9174 , n7464 );
    or g10040 ( n3300 , n7438 , n4751 );
    not g10041 ( n7053 , n5618 );
    not g10042 ( n9924 , n6516 );
    nor g10043 ( n6302 , n8920 , n14508 );
    not g10044 ( n1962 , n7346 );
    and g10045 ( n1960 , n13421 , n13023 );
    and g10046 ( n4325 , n14164 , n8540 );
    or g10047 ( n6352 , n2017 , n4795 );
    or g10048 ( n8408 , n2218 , n11018 );
    and g10049 ( n8901 , n13720 , n14031 );
    or g10050 ( n13761 , n5562 , n1168 );
    or g10051 ( n3149 , n6242 , n4599 );
    and g10052 ( n2100 , n11569 , n12471 );
    or g10053 ( n8479 , n9151 , n1445 );
    or g10054 ( n13254 , n976 , n4874 );
    nor g10055 ( n6457 , n3457 , n14204 );
    not g10056 ( n12986 , n11425 );
    or g10057 ( n12290 , n4739 , n3237 );
    and g10058 ( n5303 , n2724 , n5716 );
    and g10059 ( n5726 , n1854 , n4529 );
    and g10060 ( n10817 , n748 , n1657 );
    not g10061 ( n6695 , n5901 );
    nor g10062 ( n14284 , n1638 , n2917 );
    and g10063 ( n14325 , n10032 , n1128 );
    and g10064 ( n2706 , n638 , n12241 );
    or g10065 ( n14124 , n13108 , n10165 );
    and g10066 ( n0 , n8605 , n11884 );
    or g10067 ( n12397 , n4404 , n10112 );
    or g10068 ( n5055 , n13531 , n5143 );
    or g10069 ( n2289 , n13978 , n12176 );
    or g10070 ( n8116 , n5007 , n5622 );
    and g10071 ( n5109 , n12998 , n11320 );
    and g10072 ( n8838 , n6854 , n11914 );
    or g10073 ( n12081 , n172 , n11707 );
    and g10074 ( n4775 , n9617 , n2093 );
    or g10075 ( n5666 , n6323 , n13846 );
    and g10076 ( n12868 , n1708 , n12889 );
    and g10077 ( n2496 , n678 , n6750 );
    not g10078 ( n8476 , n10775 );
    or g10079 ( n12742 , n8527 , n8324 );
    not g10080 ( n3428 , n13544 );
    or g10081 ( n13690 , n12844 , n12903 );
    nor g10082 ( n1899 , n2468 , n13947 );
    not g10083 ( n5048 , n6088 );
    or g10084 ( n9212 , n8592 , n2618 );
    or g10085 ( n11655 , n13118 , n13126 );
    and g10086 ( n7777 , n5899 , n10852 );
    nor g10087 ( n5098 , n234 , n4818 );
    nor g10088 ( n11971 , n4633 , n159 );
    or g10089 ( n11644 , n9856 , n13591 );
    or g10090 ( n12582 , n4967 , n9070 );
    or g10091 ( n1913 , n5569 , n11076 );
    nor g10092 ( n1065 , n7345 , n1167 );
    or g10093 ( n83 , n5732 , n2589 );
    and g10094 ( n12964 , n14065 , n6134 );
    nor g10095 ( n3676 , n11508 , n12681 );
    and g10096 ( n13796 , n8786 , n14079 );
    and g10097 ( n7347 , n2158 , n4670 );
    not g10098 ( n8398 , n10688 );
    or g10099 ( n771 , n10191 , n4078 );
    not g10100 ( n5118 , n2250 );
    or g10101 ( n12760 , n2315 , n9273 );
    not g10102 ( n6697 , n7091 );
    nor g10103 ( n4580 , n5026 , n10088 );
    and g10104 ( n5485 , n5779 , n1909 );
    and g10105 ( n8033 , n12802 , n9300 );
    and g10106 ( n5759 , n2669 , n5270 );
    and g10107 ( n3911 , n7529 , n20 );
    not g10108 ( n13656 , n13139 );
    nor g10109 ( n8286 , n13941 , n9352 );
    not g10110 ( n11008 , n6829 );
    nor g10111 ( n2631 , n11581 , n8330 );
    not g10112 ( n8555 , n2298 );
    and g10113 ( n720 , n748 , n5655 );
    or g10114 ( n6272 , n12019 , n13800 );
    and g10115 ( n14073 , n4722 , n13059 );
    and g10116 ( n3224 , n286 , n10584 );
    nor g10117 ( n7500 , n12322 , n12937 );
    and g10118 ( n1989 , n1610 , n12566 );
    not g10119 ( n14430 , n12588 );
    or g10120 ( n7892 , n13413 , n14162 );
    not g10121 ( n12957 , n14433 );
    and g10122 ( n1115 , n7911 , n3348 );
    and g10123 ( n5462 , n1699 , n6495 );
    or g10124 ( n4479 , n4925 , n1898 );
    or g10125 ( n7241 , n6981 , n427 );
    nor g10126 ( n8312 , n9984 , n6 );
    or g10127 ( n2800 , n5472 , n7018 );
    or g10128 ( n8014 , n13016 , n7959 );
    not g10129 ( n10300 , n9878 );
    or g10130 ( n347 , n10035 , n191 );
    not g10131 ( n9124 , n5921 );
    and g10132 ( n13131 , n10969 , n2173 );
    and g10133 ( n11627 , n9186 , n12423 );
    not g10134 ( n13354 , n203 );
    and g10135 ( n13988 , n1489 , n5523 );
    and g10136 ( n9332 , n1125 , n3118 );
    or g10137 ( n5719 , n8964 , n4617 );
    or g10138 ( n9356 , n7812 , n7721 );
    not g10139 ( n7223 , n10055 );
    not g10140 ( n13522 , n13784 );
    and g10141 ( n6014 , n13489 , n4676 );
    and g10142 ( n10987 , n4973 , n6870 );
    or g10143 ( n7935 , n10351 , n5222 );
    and g10144 ( n1900 , n730 , n9444 );
    and g10145 ( n5353 , n13850 , n10873 );
    and g10146 ( n9846 , n513 , n34 );
    or g10147 ( n3835 , n611 , n2309 );
    or g10148 ( n9362 , n11804 , n9051 );
    nor g10149 ( n12030 , n8825 , n6335 );
    and g10150 ( n11257 , n7693 , n9976 );
    and g10151 ( n2957 , n5312 , n10544 );
    and g10152 ( n11003 , n2583 , n13833 );
    nor g10153 ( n13274 , n6672 , n9653 );
    and g10154 ( n8787 , n6016 , n13177 );
    or g10155 ( n11779 , n11420 , n8680 );
    and g10156 ( n564 , n7673 , n3176 );
    or g10157 ( n6042 , n11171 , n12919 );
    not g10158 ( n7596 , n11628 );
    or g10159 ( n13665 , n3047 , n8377 );
    and g10160 ( n3470 , n225 , n998 );
    nor g10161 ( n386 , n10637 , n14174 );
    or g10162 ( n4335 , n3126 , n8382 );
    or g10163 ( n12206 , n5815 , n8493 );
    or g10164 ( n7626 , n11315 , n5709 );
    not g10165 ( n9172 , n2417 );
    and g10166 ( n296 , n7529 , n8574 );
    or g10167 ( n6930 , n3134 , n13615 );
    and g10168 ( n3280 , n11117 , n12298 );
    not g10169 ( n8453 , n13219 );
    and g10170 ( n14160 , n13520 , n10586 );
    and g10171 ( n1176 , n4347 , n13604 );
    or g10172 ( n13951 , n13706 , n6455 );
    or g10173 ( n11880 , n11909 , n7009 );
    and g10174 ( n13182 , n10506 , n5107 );
    nor g10175 ( n14170 , n13153 , n3990 );
    and g10176 ( n8922 , n11157 , n13716 );
    or g10177 ( n14100 , n12844 , n11310 );
    or g10178 ( n12674 , n11183 , n11292 );
    nor g10179 ( n8727 , n12127 , n11283 );
    nor g10180 ( n8158 , n4572 , n6278 );
    or g10181 ( n3925 , n2874 , n1025 );
    or g10182 ( n1837 , n1535 , n10600 );
    and g10183 ( n7220 , n4244 , n3347 );
    and g10184 ( n337 , n1140 , n1360 );
    and g10185 ( n179 , n7963 , n5654 );
    not g10186 ( n14106 , n9863 );
    or g10187 ( n12085 , n9804 , n581 );
    not g10188 ( n7027 , n8361 );
    or g10189 ( n5686 , n3546 , n1563 );
    not g10190 ( n4527 , n10630 );
    nor g10191 ( n10317 , n8767 , n5214 );
    and g10192 ( n6845 , n11816 , n7817 );
    or g10193 ( n1330 , n11036 , n7424 );
    and g10194 ( n9667 , n2158 , n9480 );
    or g10195 ( n11608 , n3815 , n6578 );
    not g10196 ( n6531 , n10377 );
    and g10197 ( n2634 , n7267 , n13330 );
    or g10198 ( n3589 , n4631 , n9153 );
    nor g10199 ( n9862 , n6933 , n7459 );
    not g10200 ( n3011 , n918 );
    nor g10201 ( n11353 , n2057 , n3446 );
    or g10202 ( n14244 , n1701 , n2442 );
    or g10203 ( n2801 , n1356 , n9917 );
    and g10204 ( n7613 , n13464 , n2244 );
    not g10205 ( n10035 , n1676 );
    or g10206 ( n8350 , n13991 , n8989 );
    or g10207 ( n12342 , n8490 , n14474 );
    nor g10208 ( n14250 , n5944 , n10355 );
    and g10209 ( n11210 , n7267 , n6179 );
    or g10210 ( n11629 , n8210 , n1689 );
    and g10211 ( n9860 , n12250 , n6566 );
    or g10212 ( n13299 , n11090 , n10382 );
    and g10213 ( n4794 , n6354 , n4571 );
    not g10214 ( n788 , n2226 );
    and g10215 ( n5163 , n10330 , n9210 );
    or g10216 ( n10720 , n4357 , n970 );
    and g10217 ( n7157 , n11153 , n2423 );
    nor g10218 ( n13062 , n14198 , n11512 );
    not g10219 ( n5092 , n5606 );
    and g10220 ( n7254 , n10566 , n7149 );
    and g10221 ( n5731 , n13823 , n1430 );
    or g10222 ( n1700 , n11011 , n2782 );
    or g10223 ( n9561 , n13885 , n1397 );
    or g10224 ( n8063 , n619 , n1368 );
    not g10225 ( n9620 , n9596 );
    or g10226 ( n12804 , n2877 , n2676 );
    or g10227 ( n4254 , n12292 , n14452 );
    nor g10228 ( n2834 , n2098 , n6315 );
    and g10229 ( n11635 , n2564 , n11527 );
    nor g10230 ( n2739 , n2651 , n11535 );
    and g10231 ( n13166 , n12039 , n4776 );
    and g10232 ( n3426 , n8147 , n1964 );
    or g10233 ( n7056 , n6147 , n11842 );
    not g10234 ( n1231 , n5197 );
    and g10235 ( n5360 , n1857 , n7351 );
    and g10236 ( n12985 , n14321 , n5567 );
    or g10237 ( n2657 , n2229 , n10164 );
    not g10238 ( n1741 , n7404 );
    and g10239 ( n1270 , n6128 , n7945 );
    and g10240 ( n4921 , n6507 , n7405 );
    not g10241 ( n3565 , n1462 );
    or g10242 ( n14477 , n954 , n2861 );
    and g10243 ( n8457 , n13597 , n1252 );
    or g10244 ( n10451 , n13432 , n10721 );
    or g10245 ( n1229 , n9140 , n14309 );
    or g10246 ( n513 , n582 , n4774 );
    or g10247 ( n11593 , n13005 , n3453 );
    or g10248 ( n1680 , n6323 , n4764 );
    nor g10249 ( n1652 , n7091 , n11469 );
    not g10250 ( n8020 , n7223 );
    not g10251 ( n5139 , n9580 );
    and g10252 ( n1240 , n4803 , n7578 );
    or g10253 ( n2937 , n1172 , n909 );
    nor g10254 ( n6798 , n7364 , n14385 );
    and g10255 ( n54 , n11814 , n9184 );
    and g10256 ( n5287 , n12461 , n6304 );
    not g10257 ( n7438 , n628 );
    or g10258 ( n4936 , n10234 , n6728 );
    or g10259 ( n10537 , n317 , n11524 );
    or g10260 ( n9384 , n1840 , n7509 );
    not g10261 ( n13682 , n10061 );
    or g10262 ( n11355 , n974 , n4725 );
    or g10263 ( n11894 , n3559 , n12977 );
    and g10264 ( n901 , n98 , n4275 );
    and g10265 ( n13769 , n1937 , n7398 );
    or g10266 ( n11965 , n11620 , n4004 );
    and g10267 ( n10941 , n2758 , n2338 );
    and g10268 ( n6920 , n14321 , n10611 );
    and g10269 ( n6010 , n3743 , n11509 );
    not g10270 ( n2006 , n10177 );
    nor g10271 ( n9475 , n5365 , n2185 );
    and g10272 ( n3278 , n12226 , n10288 );
    nor g10273 ( n11446 , n8527 , n6386 );
    and g10274 ( n11851 , n9853 , n11735 );
    not g10275 ( n8047 , n920 );
    not g10276 ( n4741 , n7819 );
    and g10277 ( n12355 , n14464 , n12766 );
    or g10278 ( n6162 , n1361 , n13093 );
    or g10279 ( n14484 , n5575 , n10675 );
    or g10280 ( n924 , n10461 , n3326 );
    and g10281 ( n4998 , n14145 , n484 );
    and g10282 ( n6411 , n2527 , n614 );
    not g10283 ( n3675 , n3166 );
    or g10284 ( n3549 , n14210 , n8649 );
    and g10285 ( n4089 , n2322 , n992 );
    and g10286 ( n6658 , n7026 , n2088 );
    not g10287 ( n4435 , n1267 );
    and g10288 ( n4842 , n13252 , n8421 );
    or g10289 ( n14350 , n2531 , n2557 );
    or g10290 ( n8659 , n492 , n10636 );
    not g10291 ( n12294 , n3704 );
    and g10292 ( n4427 , n7957 , n12178 );
    or g10293 ( n12212 , n7436 , n9224 );
    and g10294 ( n13744 , n4354 , n3086 );
    and g10295 ( n5081 , n9198 , n2051 );
    and g10296 ( n816 , n1074 , n223 );
    or g10297 ( n12840 , n553 , n3738 );
    and g10298 ( n1041 , n7814 , n8398 );
    and g10299 ( n9091 , n13850 , n10220 );
    or g10300 ( n2508 , n9140 , n9093 );
    not g10301 ( n4929 , n13981 );
    not g10302 ( n7443 , n8451 );
    and g10303 ( n5633 , n5104 , n1415 );
    and g10304 ( n9013 , n12412 , n10747 );
    or g10305 ( n13482 , n14088 , n10522 );
    or g10306 ( n6968 , n1820 , n7409 );
    nor g10307 ( n9875 , n1612 , n11051 );
    and g10308 ( n12987 , n783 , n9117 );
    or g10309 ( n10550 , n5997 , n497 );
    or g10310 ( n1088 , n6263 , n13821 );
    or g10311 ( n6215 , n8096 , n835 );
    not g10312 ( n12139 , n4891 );
    and g10313 ( n13203 , n14091 , n9459 );
    or g10314 ( n10798 , n10396 , n10742 );
    and g10315 ( n10602 , n13096 , n7123 );
    or g10316 ( n4120 , n13155 , n4868 );
    not g10317 ( n11771 , n3280 );
    or g10318 ( n3622 , n4199 , n10905 );
    not g10319 ( n14465 , n8963 );
    nor g10320 ( n1714 , n9754 , n2233 );
    and g10321 ( n3174 , n5048 , n1986 );
    not g10322 ( n2058 , n10254 );
    not g10323 ( n14296 , n9182 );
    or g10324 ( n6802 , n1728 , n3022 );
    not g10325 ( n10646 , n10378 );
    and g10326 ( n6348 , n2583 , n11065 );
    and g10327 ( n3962 , n11157 , n2779 );
    and g10328 ( n6001 , n13641 , n149 );
    or g10329 ( n10890 , n6595 , n6865 );
    or g10330 ( n12854 , n1189 , n7863 );
    or g10331 ( n1109 , n5873 , n10255 );
    or g10332 ( n11874 , n3667 , n10577 );
    and g10333 ( n8808 , n3904 , n2237 );
    and g10334 ( n12604 , n10815 , n8185 );
    not g10335 ( n3191 , n12403 );
    and g10336 ( n12735 , n3286 , n7772 );
    not g10337 ( n5159 , n1365 );
    and g10338 ( n1895 , n10197 , n3728 );
    nor g10339 ( n516 , n6434 , n10963 );
    and g10340 ( n3879 , n1409 , n2316 );
    and g10341 ( n10375 , n2473 , n8743 );
    or g10342 ( n12478 , n1834 , n3174 );
    and g10343 ( n8954 , n9944 , n14428 );
    or g10344 ( n2558 , n1494 , n10718 );
    and g10345 ( n12219 , n14358 , n12228 );
    not g10346 ( n12765 , n10047 );
    or g10347 ( n12942 , n3134 , n5753 );
    or g10348 ( n13721 , n14366 , n5314 );
    or g10349 ( n586 , n1391 , n9308 );
    nor g10350 ( n4185 , n5986 , n12508 );
    and g10351 ( n5214 , n3861 , n4318 );
    nor g10352 ( n4747 , n3768 , n9395 );
    and g10353 ( n1715 , n11163 , n5925 );
    or g10354 ( n7521 , n888 , n12829 );
    not g10355 ( n12630 , n7846 );
    nor g10356 ( n2881 , n7584 , n609 );
    or g10357 ( n11966 , n13354 , n737 );
    and g10358 ( n4715 , n13017 , n3817 );
    or g10359 ( n5478 , n553 , n2460 );
    or g10360 ( n6925 , n4313 , n13628 );
    and g10361 ( n11034 , n5335 , n7420 );
    and g10362 ( n10970 , n4347 , n9876 );
    or g10363 ( n6809 , n2686 , n6659 );
    and g10364 ( n14429 , n1254 , n13836 );
    not g10365 ( n14358 , n7507 );
    not g10366 ( n9190 , n1417 );
    and g10367 ( n637 , n5414 , n310 );
    and g10368 ( n10717 , n12159 , n2249 );
    not g10369 ( n12450 , n10055 );
    or g10370 ( n11663 , n3886 , n13942 );
    nor g10371 ( n5385 , n12548 , n13672 );
    or g10372 ( n9427 , n5480 , n11023 );
    or g10373 ( n4226 , n791 , n9961 );
    and g10374 ( n8809 , n10059 , n13259 );
    not g10375 ( n5011 , n168 );
    and g10376 ( n1759 , n4276 , n6108 );
    and g10377 ( n9222 , n6609 , n9433 );
    not g10378 ( n6559 , n11264 );
    or g10379 ( n1971 , n7250 , n5819 );
    not g10380 ( n10294 , n426 );
    and g10381 ( n8094 , n9952 , n8327 );
    or g10382 ( n7226 , n7481 , n13171 );
    or g10383 ( n5219 , n3025 , n5546 );
    and g10384 ( n10174 , n7043 , n4855 );
    or g10385 ( n10455 , n5084 , n8765 );
    or g10386 ( n2746 , n2784 , n137 );
    not g10387 ( n5795 , n6534 );
    not g10388 ( n898 , n442 );
    and g10389 ( n11018 , n12105 , n5809 );
    and g10390 ( n9464 , n12472 , n9301 );
    and g10391 ( n10685 , n10015 , n4578 );
    or g10392 ( n7883 , n3914 , n2266 );
    and g10393 ( n13793 , n7421 , n2287 );
    nor g10394 ( n3040 , n5288 , n1534 );
    or g10395 ( n12261 , n10913 , n9149 );
    and g10396 ( n14287 , n9297 , n7731 );
    nor g10397 ( n7234 , n8015 , n4110 );
    not g10398 ( n1854 , n304 );
    or g10399 ( n4487 , n10871 , n8307 );
    and g10400 ( n9022 , n12528 , n1557 );
    and g10401 ( n11368 , n5335 , n6635 );
    or g10402 ( n3249 , n782 , n9873 );
    and g10403 ( n1353 , n6016 , n5697 );
    and g10404 ( n9281 , n8372 , n13832 );
    not g10405 ( n2877 , n3070 );
    not g10406 ( n3025 , n5627 );
    or g10407 ( n9857 , n3800 , n13441 );
    or g10408 ( n10335 , n2597 , n3063 );
    or g10409 ( n9681 , n11183 , n854 );
    or g10410 ( n5988 , n12169 , n6381 );
    or g10411 ( n4683 , n9229 , n9723 );
    nor g10412 ( n9768 , n1769 , n10349 );
    and g10413 ( n6329 , n8965 , n1493 );
    or g10414 ( n12996 , n8242 , n14489 );
    not g10415 ( n4320 , n4117 );
    and g10416 ( n13269 , n10710 , n10702 );
    and g10417 ( n2831 , n7068 , n1313 );
    and g10418 ( n5853 , n13781 , n9970 );
    and g10419 ( n10657 , n3401 , n9435 );
    and g10420 ( n13067 , n14373 , n6967 );
    not g10421 ( n10121 , n7979 );
    and g10422 ( n11120 , n8507 , n5196 );
    not g10423 ( n8189 , n496 );
    or g10424 ( n12463 , n11572 , n14032 );
    and g10425 ( n8281 , n11748 , n3207 );
    nor g10426 ( n14246 , n1623 , n14384 );
    not g10427 ( n10036 , n1938 );
    and g10428 ( n2656 , n9853 , n9533 );
    or g10429 ( n9800 , n361 , n3814 );
    or g10430 ( n4529 , n13477 , n3954 );
    and g10431 ( n13064 , n13246 , n3298 );
    and g10432 ( n6385 , n7421 , n8479 );
    and g10433 ( n7020 , n873 , n11173 );
    not g10434 ( n11515 , n300 );
    and g10435 ( n4051 , n13404 , n14177 );
    or g10436 ( n11585 , n4065 , n8235 );
    and g10437 ( n11324 , n4698 , n1395 );
    and g10438 ( n2721 , n1452 , n5494 );
    or g10439 ( n10725 , n5064 , n4374 );
    or g10440 ( n3192 , n10461 , n2494 );
    or g10441 ( n12154 , n3099 , n1308 );
    and g10442 ( n7369 , n12101 , n1831 );
    or g10443 ( n14413 , n12543 , n7800 );
    not g10444 ( n12568 , n9846 );
    not g10445 ( n782 , n12746 );
    or g10446 ( n11087 , n12139 , n7877 );
    not g10447 ( n6787 , n885 );
    and g10448 ( n829 , n4525 , n9168 );
    or g10449 ( n415 , n14337 , n2435 );
    or g10450 ( n5758 , n568 , n11210 );
    nor g10451 ( n12002 , n5569 , n1851 );
    and g10452 ( n5003 , n7068 , n1419 );
    and g10453 ( n3111 , n55 , n5526 );
    and g10454 ( n4084 , n3861 , n3411 );
    not g10455 ( n3434 , n2029 );
    or g10456 ( n11402 , n7438 , n5091 );
    not g10457 ( n2082 , n7681 );
    or g10458 ( n1648 , n11951 , n9324 );
    nor g10459 ( n858 , n11047 , n3645 );
    not g10460 ( n7693 , n11425 );
    and g10461 ( n3175 , n6753 , n1187 );
    not g10462 ( n12922 , n7077 );
    and g10463 ( n7315 , n3485 , n11840 );
    nor g10464 ( n10814 , n12968 , n10200 );
    or g10465 ( n154 , n4435 , n2710 );
    or g10466 ( n2142 , n11953 , n3744 );
    nor g10467 ( n10793 , n7145 , n8818 );
    and g10468 ( n120 , n4806 , n7611 );
    not g10469 ( n8726 , n2545 );
    or g10470 ( n10427 , n12023 , n8177 );
    nor g10471 ( n12024 , n8363 , n6477 );
    and g10472 ( n8136 , n11020 , n13758 );
    or g10473 ( n10852 , n6350 , n907 );
    not g10474 ( n8288 , n1086 );
    or g10475 ( n12837 , n8825 , n5141 );
    or g10476 ( n280 , n10784 , n13913 );
    or g10477 ( n5713 , n8209 , n13470 );
    and g10478 ( n9547 , n8801 , n2687 );
    or g10479 ( n3594 , n12034 , n9250 );
    nor g10480 ( n8101 , n1813 , n12316 );
    and g10481 ( n914 , n2533 , n5417 );
    or g10482 ( n11189 , n10083 , n10336 );
    and g10483 ( n4846 , n7211 , n14442 );
    not g10484 ( n6318 , n13723 );
    and g10485 ( n2639 , n8427 , n11759 );
    and g10486 ( n8220 , n2529 , n13840 );
    not g10487 ( n7007 , n4210 );
    nor g10488 ( n2879 , n4544 , n10980 );
    or g10489 ( n6903 , n13682 , n12885 );
    nor g10490 ( n9990 , n717 , n4201 );
    and g10491 ( n5398 , n1225 , n11062 );
    or g10492 ( n890 , n5762 , n5441 );
    and g10493 ( n14482 , n11803 , n14124 );
    or g10494 ( n6134 , n8866 , n7282 );
    not g10495 ( n3419 , n2573 );
    and g10496 ( n12938 , n1699 , n3249 );
    and g10497 ( n1770 , n12986 , n7353 );
    and g10498 ( n13440 , n10015 , n12567 );
    or g10499 ( n3343 , n1172 , n7032 );
    or g10500 ( n181 , n387 , n380 );
    or g10501 ( n14499 , n3099 , n8838 );
    nor g10502 ( n7658 , n8544 , n2666 );
    and g10503 ( n12660 , n3247 , n8685 );
    not g10504 ( n13755 , n11369 );
    or g10505 ( n12413 , n2874 , n2327 );
    and g10506 ( n182 , n2099 , n5528 );
    nor g10507 ( n7372 , n14058 , n5902 );
    and g10508 ( n7388 , n98 , n449 );
    or g10509 ( n2456 , n2747 , n4167 );
    and g10510 ( n3147 , n904 , n2989 );
    and g10511 ( n3090 , n650 , n14222 );
    nor g10512 ( n322 , n5509 , n2170 );
    not g10513 ( n2474 , n5014 );
    or g10514 ( n11394 , n3512 , n11701 );
    and g10515 ( n3691 , n6507 , n3002 );
    and g10516 ( n3918 , n6848 , n9031 );
    or g10517 ( n6562 , n2908 , n3533 );
    or g10518 ( n11983 , n5997 , n4257 );
    or g10519 ( n11126 , n12034 , n6010 );
    or g10520 ( n10683 , n412 , n13795 );
    not g10521 ( n12209 , n7104 );
    and g10522 ( n7451 , n3607 , n14425 );
    or g10523 ( n1781 , n11440 , n5388 );
    or g10524 ( n10614 , n227 , n7813 );
    and g10525 ( n12106 , n5734 , n13002 );
    not g10526 ( n3461 , n9563 );
    and g10527 ( n13798 , n5899 , n6115 );
    and g10528 ( n2239 , n14157 , n7653 );
    not g10529 ( n11988 , n10358 );
    and g10530 ( n11122 , n8649 , n7124 );
    not g10531 ( n7973 , n7177 );
    and g10532 ( n12338 , n8697 , n10768 );
    not g10533 ( n8450 , n6758 );
    or g10534 ( n7309 , n13728 , n13102 );
    or g10535 ( n950 , n3287 , n8419 );
    and g10536 ( n8381 , n12531 , n9083 );
    not g10537 ( n3219 , n9306 );
    or g10538 ( n11256 , n10624 , n1716 );
    or g10539 ( n9516 , n1401 , n6693 );
    nor g10540 ( n7806 , n4299 , n12672 );
    or g10541 ( n3106 , n8404 , n7894 );
    and g10542 ( n2490 , n6744 , n9427 );
    not g10543 ( n12548 , n11435 );
    or g10544 ( n7082 , n7898 , n7324 );
    or g10545 ( n12537 , n14188 , n10078 );
    or g10546 ( n3329 , n11647 , n5679 );
    and g10547 ( n6106 , n6507 , n111 );
    and g10548 ( n5402 , n6013 , n7595 );
    not g10549 ( n3402 , n14365 );
    and g10550 ( n589 , n3952 , n2050 );
    and g10551 ( n13162 , n2820 , n3537 );
    not g10552 ( n8212 , n7007 );
    or g10553 ( n13368 , n12576 , n2449 );
    and g10554 ( n6066 , n13379 , n3350 );
    not g10555 ( n3395 , n9740 );
    or g10556 ( n6286 , n3527 , n5535 );
    or g10557 ( n493 , n10136 , n12773 );
    and g10558 ( n5607 , n889 , n10940 );
    not g10559 ( n14319 , n12394 );
    or g10560 ( n8681 , n12169 , n7881 );
    or g10561 ( n4727 , n647 , n7659 );
    and g10562 ( n1641 , n4289 , n6803 );
    or g10563 ( n13457 , n12820 , n11513 );
    or g10564 ( n2043 , n7527 , n5545 );
    or g10565 ( n10748 , n10323 , n7472 );
    and g10566 ( n622 , n7979 , n4713 );
    and g10567 ( n8375 , n428 , n11550 );
    and g10568 ( n10359 , n9944 , n856 );
    not g10569 ( n12870 , n12444 );
    and g10570 ( n13651 , n55 , n7111 );
    and g10571 ( n8832 , n5275 , n11197 );
    or g10572 ( n4068 , n13707 , n7687 );
    and g10573 ( n3279 , n2587 , n3801 );
    or g10574 ( n12756 , n10035 , n4099 );
    nor g10575 ( n4693 , n12968 , n6551 );
    or g10576 ( n13655 , n7527 , n3614 );
    and g10577 ( n12176 , n11702 , n6356 );
    and g10578 ( n6415 , n7284 , n10538 );
    not g10579 ( n8023 , n5738 );
    and g10580 ( n9242 , n2564 , n414 );
    not g10581 ( n12601 , n13165 );
    or g10582 ( n6599 , n11231 , n1075 );
    and g10583 ( n9233 , n405 , n10829 );
    and g10584 ( n10043 , n13700 , n3711 );
    or g10585 ( n2480 , n1031 , n3349 );
    and g10586 ( n7467 , n13147 , n7384 );
    not g10587 ( n10516 , n8008 );
    and g10588 ( n9103 , n7429 , n362 );
    not g10589 ( n10062 , n13668 );
    not g10590 ( n2137 , n12136 );
    not g10591 ( n98 , n11547 );
    and g10592 ( n7464 , n14093 , n896 );
    or g10593 ( n2065 , n8425 , n6938 );
    or g10594 ( n5658 , n1031 , n668 );
    and g10595 ( n7547 , n11607 , n5496 );
    or g10596 ( n1412 , n10713 , n157 );
    or g10597 ( n7513 , n10024 , n7734 );
    or g10598 ( n9622 , n9804 , n11290 );
    and g10599 ( n8440 , n3846 , n2268 );
    and g10600 ( n10116 , n3942 , n14161 );
    nor g10601 ( n5941 , n7466 , n7397 );
    not g10602 ( n4988 , n9354 );
    or g10603 ( n10142 , n10089 , n13712 );
    not g10604 ( n12807 , n9769 );
    or g10605 ( n12187 , n8480 , n13828 );
    or g10606 ( n8036 , n11047 , n5425 );
    and g10607 ( n6182 , n1804 , n3172 );
    or g10608 ( n6965 , n9562 , n6586 );
    or g10609 ( n9511 , n5715 , n10192 );
    or g10610 ( n61 , n5603 , n6377 );
    or g10611 ( n8248 , n647 , n7329 );
    and g10612 ( n2204 , n2583 , n3398 );
    and g10613 ( n13815 , n3485 , n2393 );
    and g10614 ( n9308 , n9232 , n295 );
    nor g10615 ( n6217 , n11980 , n430 );
    and g10616 ( n5082 , n7717 , n9882 );
    and g10617 ( n477 , n898 , n3403 );
    or g10618 ( n2035 , n3164 , n10810 );
    or g10619 ( n5138 , n2218 , n11245 );
    or g10620 ( n2994 , n9716 , n65 );
    and g10621 ( n3994 , n3904 , n2563 );
    or g10622 ( n3786 , n1535 , n3220 );
    and g10623 ( n8434 , n14465 , n6078 );
    or g10624 ( n10111 , n10351 , n5347 );
    and g10625 ( n2257 , n6556 , n10880 );
    and g10626 ( n10699 , n10820 , n173 );
    and g10627 ( n12684 , n13489 , n3341 );
    not g10628 ( n7334 , n3191 );
    or g10629 ( n1359 , n13432 , n7368 );
    or g10630 ( n2514 , n4923 , n2864 );
    and g10631 ( n5090 , n7596 , n7325 );
    and g10632 ( n13304 , n4300 , n5357 );
    or g10633 ( n9272 , n13869 , n8892 );
    or g10634 ( n797 , n523 , n13799 );
    and g10635 ( n2594 , n6192 , n12582 );
    not g10636 ( n14196 , n752 );
    and g10637 ( n6447 , n8372 , n6161 );
    and g10638 ( n662 , n7015 , n6685 );
    not g10639 ( n5921 , n4928 );
    or g10640 ( n6669 , n7683 , n9446 );
    and g10641 ( n4343 , n7063 , n6024 );
    and g10642 ( n8061 , n5876 , n7142 );
    or g10643 ( n3885 , n9620 , n11851 );
    nor g10644 ( n13892 , n8816 , n12238 );
    and g10645 ( n2525 , n1775 , n794 );
    or g10646 ( n5113 , n9856 , n7016 );
    or g10647 ( n7176 , n5236 , n4729 );
    or g10648 ( n11919 , n2179 , n11618 );
    and g10649 ( n4181 , n7810 , n6341 );
    or g10650 ( n3903 , n6046 , n7131 );
    nor g10651 ( n11911 , n6989 , n12298 );
    and g10652 ( n2442 , n14321 , n14302 );
    or g10653 ( n12534 , n9442 , n296 );
    or g10654 ( n12814 , n3161 , n4015 );
    not g10655 ( n13055 , n937 );
    or g10656 ( n5154 , n2149 , n10167 );
    or g10657 ( n10218 , n9490 , n1129 );
    and g10658 ( n9850 , n4574 , n256 );
    nor g10659 ( n8138 , n1706 , n14057 );
    or g10660 ( n2691 , n2218 , n7775 );
    and g10661 ( n5383 , n1588 , n11312 );
    or g10662 ( n5684 , n6706 , n10259 );
    or g10663 ( n13323 , n8575 , n10797 );
    not g10664 ( n10678 , n14501 );
    and g10665 ( n5657 , n7057 , n9554 );
    not g10666 ( n13153 , n4007 );
    and g10667 ( n6726 , n4932 , n9163 );
    not g10668 ( n6649 , n7621 );
    not g10669 ( n8721 , n5943 );
    or g10670 ( n12545 , n1147 , n1089 );
    and g10671 ( n11457 , n9745 , n5875 );
    and g10672 ( n13165 , n11052 , n9751 );
    and g10673 ( n6793 , n3286 , n9194 );
    not g10674 ( n12047 , n6804 );
    and g10675 ( n4854 , n8007 , n12122 );
    nor g10676 ( n956 , n9035 , n2302 );
    and g10677 ( n10965 , n3709 , n8794 );
    not g10678 ( n172 , n11456 );
    nor g10679 ( n3517 , n7971 , n8643 );
    not g10680 ( n4973 , n13003 );
    not g10681 ( n13531 , n3681 );
    or g10682 ( n8364 , n7003 , n2477 );
    and g10683 ( n4114 , n10822 , n5304 );
    or g10684 ( n3376 , n2877 , n10888 );
    not g10685 ( n2224 , n4618 );
    or g10686 ( n6605 , n7426 , n12711 );
    not g10687 ( n11574 , n4050 );
    or g10688 ( n11358 , n4876 , n9918 );
    or g10689 ( n38 , n10960 , n8937 );
    not g10690 ( n7523 , n13102 );
    not g10691 ( n8817 , n737 );
    or g10692 ( n12121 , n13912 , n12218 );
    and g10693 ( n9286 , n6525 , n12301 );
    or g10694 ( n4264 , n12549 , n4590 );
    or g10695 ( n11182 , n12870 , n9798 );
    or g10696 ( n7710 , n2188 , n6114 );
    nor g10697 ( n10655 , n7359 , n4455 );
    not g10698 ( n8372 , n1478 );
    and g10699 ( n9099 , n14388 , n5789 );
    not g10700 ( n7003 , n9371 );
    not g10701 ( n6819 , n1979 );
    and g10702 ( n4985 , n7081 , n14457 );
    or g10703 ( n2563 , n13074 , n12952 );
    not g10704 ( n13248 , n9231 );
    nor g10705 ( n8991 , n13874 , n12224 );
    and g10706 ( n409 , n12850 , n13257 );
    or g10707 ( n10740 , n511 , n1115 );
    not g10708 ( n10803 , n3544 );
    and g10709 ( n10943 , n3435 , n14292 );
    and g10710 ( n6885 , n7043 , n3030 );
    and g10711 ( n6837 , n7208 , n12056 );
    and g10712 ( n13470 , n2224 , n2127 );
    or g10713 ( n9260 , n5625 , n4881 );
    and g10714 ( n10071 , n13069 , n6947 );
    not g10715 ( n6139 , n3493 );
    and g10716 ( n124 , n10589 , n6170 );
    and g10717 ( n13492 , n10506 , n9734 );
    nor g10718 ( n3272 , n10091 , n9400 );
    or g10719 ( n3031 , n2229 , n6564 );
    or g10720 ( n8992 , n10351 , n3539 );
    or g10721 ( n9868 , n12543 , n13382 );
    and g10722 ( n3941 , n1354 , n5885 );
    nor g10723 ( n8518 , n3211 , n13121 );
    and g10724 ( n4668 , n10197 , n6720 );
    nor g10725 ( n1219 , n2171 , n14116 );
    and g10726 ( n7191 , n8111 , n8667 );
    not g10727 ( n1258 , n9354 );
    or g10728 ( n7636 , n5132 , n5313 );
    and g10729 ( n8465 , n5434 , n1212 );
    nor g10730 ( n2467 , n11017 , n1432 );
    and g10731 ( n11525 , n7429 , n508 );
    or g10732 ( n11658 , n387 , n6939 );
    or g10733 ( n6814 , n555 , n10440 );
    and g10734 ( n5378 , n2985 , n6391 );
    and g10735 ( n1625 , n5899 , n5334 );
    or g10736 ( n7929 , n9228 , n1637 );
    and g10737 ( n5291 , n10930 , n13805 );
    not g10738 ( n12691 , n1812 );
    or g10739 ( n11972 , n7426 , n212 );
    not g10740 ( n7621 , n637 );
    not g10741 ( n1713 , n8899 );
    and g10742 ( n398 , n7781 , n12435 );
    or g10743 ( n3100 , n2315 , n1517 );
    and g10744 ( n4112 , n12615 , n1939 );
    and g10745 ( n8206 , n9080 , n4178 );
    nor g10746 ( n14168 , n99 , n9985 );
    or g10747 ( n6801 , n6596 , n13064 );
    and g10748 ( n7602 , n9015 , n11642 );
    or g10749 ( n4245 , n12400 , n12905 );
    or g10750 ( n7213 , n12034 , n13456 );
    nor g10751 ( n13826 , n13055 , n12272 );
    and g10752 ( n5705 , n3491 , n1500 );
    or g10753 ( n2197 , n85 , n7321 );
    and g10754 ( n11196 , n1699 , n10258 );
    not g10755 ( n5480 , n2545 );
    or g10756 ( n9130 , n13718 , n552 );
    and g10757 ( n10779 , n1729 , n8618 );
    and g10758 ( n12812 , n12147 , n610 );
    and g10759 ( n10386 , n13700 , n12281 );
    nor g10760 ( n9092 , n4535 , n3285 );
    and g10761 ( n4389 , n405 , n14046 );
    not g10762 ( n13181 , n12409 );
    or g10763 ( n5456 , n12568 , n6197 );
    and g10764 ( n2143 , n14313 , n8896 );
    not g10765 ( n283 , n8695 );
    or g10766 ( n3144 , n14435 , n1440 );
    not g10767 ( n7365 , n12096 );
    or g10768 ( n4956 , n1356 , n14206 );
    and g10769 ( n3915 , n4901 , n13738 );
    and g10770 ( n11536 , n10969 , n2882 );
    or g10771 ( n13196 , n329 , n3807 );
    or g10772 ( n3998 , n12351 , n7499 );
    or g10773 ( n5691 , n4205 , n2876 );
    nor g10774 ( n5177 , n11597 , n12103 );
    and g10775 ( n14087 , n4276 , n10842 );
    nor g10776 ( n11730 , n3400 , n7209 );
    nor g10777 ( n1552 , n2005 , n6798 );
    or g10778 ( n13523 , n28 , n6560 );
    nor g10779 ( n8080 , n12527 , n13279 );
    and g10780 ( n11215 , n5348 , n12204 );
    not g10781 ( n2067 , n6693 );
    nor g10782 ( n6760 , n9806 , n1226 );
    or g10783 ( n10493 , n13080 , n3706 );
    nor g10784 ( n5366 , n14239 , n13892 );
    not g10785 ( n13555 , n6990 );
    not g10786 ( n2341 , n13041 );
    and g10787 ( n7411 , n7221 , n7298 );
    and g10788 ( n12150 , n3904 , n1680 );
    or g10789 ( n150 , n89 , n6579 );
    and g10790 ( n8400 , n1074 , n6570 );
    and g10791 ( n603 , n6899 , n2480 );
    not g10792 ( n2415 , n14461 );
    and g10793 ( n13837 , n10678 , n1651 );
    and g10794 ( n11290 , n4163 , n4013 );
    and g10795 ( n11205 , n10408 , n23 );
    nor g10796 ( n11114 , n7624 , n9519 );
    or g10797 ( n14156 , n11572 , n3175 );
    nor g10798 ( n12390 , n14419 , n7965 );
    not g10799 ( n2587 , n3967 );
    or g10800 ( n371 , n5548 , n8310 );
    not g10801 ( n3572 , n8798 );
    or g10802 ( n13512 , n11440 , n196 );
    and g10803 ( n9224 , n889 , n8391 );
    or g10804 ( n2020 , n5807 , n7163 );
    or g10805 ( n7525 , n11094 , n13881 );
    nor g10806 ( n13442 , n1812 , n7834 );
    not g10807 ( n2932 , n5438 );
    nor g10808 ( n11578 , n4333 , n12060 );
    or g10809 ( n5564 , n1660 , n982 );
    not g10810 ( n11223 , n13696 );
    and g10811 ( n8538 , n3028 , n11719 );
    or g10812 ( n5122 , n3011 , n5785 );
    nor g10813 ( n1426 , n7146 , n11630 );
    not g10814 ( n817 , n6264 );
    and g10815 ( n11623 , n4346 , n9626 );
    or g10816 ( n10316 , n11704 , n14374 );
    not g10817 ( n1805 , n8813 );
    and g10818 ( n4362 , n4788 , n3516 );
    not g10819 ( n13360 , n4830 );
    or g10820 ( n8736 , n12075 , n13455 );
    or g10821 ( n985 , n13220 , n3386 );
    and g10822 ( n10775 , n11100 , n12593 );
    and g10823 ( n7721 , n11220 , n6558 );
    and g10824 ( n12141 , n3586 , n5238 );
    or g10825 ( n5917 , n10784 , n6127 );
    or g10826 ( n3207 , n13112 , n4565 );
    and g10827 ( n8765 , n7060 , n10031 );
    or g10828 ( n3858 , n12130 , n6921 );
    nor g10829 ( n1327 , n7589 , n9848 );
    or g10830 ( n1828 , n11558 , n14410 );
    or g10831 ( n7560 , n1685 , n12274 );
    nor g10832 ( n86 , n4877 , n554 );
    or g10833 ( n6718 , n10394 , n9123 );
    nor g10834 ( n1460 , n11148 , n2851 );
    or g10835 ( n4054 , n12494 , n13160 );
    or g10836 ( n585 , n4615 , n730 );
    and g10837 ( n3162 , n14157 , n10140 );
    not g10838 ( n10372 , n13047 );
    not g10839 ( n11628 , n6212 );
    and g10840 ( n4015 , n9650 , n3317 );
    nor g10841 ( n2688 , n234 , n1026 );
    or g10842 ( n3393 , n12019 , n3473 );
    and g10843 ( n11922 , n2547 , n7586 );
    nor g10844 ( n6644 , n8942 , n5626 );
    not g10845 ( n8959 , n5218 );
    not g10846 ( n7529 , n4266 );
    and g10847 ( n3303 , n9811 , n11072 );
    and g10848 ( n3151 , n5471 , n13962 );
    and g10849 ( n2675 , n11422 , n9582 );
    not g10850 ( n13908 , n6058 );
    and g10851 ( n5814 , n7529 , n3578 );
    and g10852 ( n6008 , n9509 , n10890 );
    and g10853 ( n6034 , n12250 , n10509 );
    not g10854 ( n13507 , n2699 );
    or g10855 ( n8004 , n8897 , n8851 );
    or g10856 ( n3045 , n7530 , n6103 );
    or g10857 ( n6938 , n9134 , n2041 );
    and g10858 ( n13034 , n9191 , n7690 );
    or g10859 ( n8624 , n11472 , n9081 );
    or g10860 ( n12526 , n4631 , n11221 );
    and g10861 ( n8474 , n783 , n13318 );
    and g10862 ( n11291 , n4447 , n6734 );
    or g10863 ( n11981 , n9673 , n14072 );
    or g10864 ( n7814 , n9280 , n3388 );
    and g10865 ( n2381 , n1699 , n8608 );
    and g10866 ( n1046 , n7267 , n71 );
    and g10867 ( n6683 , n11220 , n6463 );
    or g10868 ( n5068 , n13142 , n8583 );
    and g10869 ( n2626 , n8605 , n4849 );
    nor g10870 ( n5250 , n4233 , n13049 );
    or g10871 ( n2032 , n10523 , n14173 );
    nor g10872 ( n75 , n4639 , n10492 );
    or g10873 ( n8973 , n9780 , n4188 );
    or g10874 ( n13180 , n8458 , n13924 );
    and g10875 ( n10206 , n11495 , n10034 );
    or g10876 ( n5682 , n5548 , n10944 );
    or g10877 ( n1668 , n14430 , n11808 );
    and g10878 ( n7880 , n3276 , n10010 );
    and g10879 ( n12989 , n3893 , n12253 );
    and g10880 ( n988 , n748 , n11319 );
    or g10881 ( n11530 , n11551 , n12710 );
    and g10882 ( n3432 , n10854 , n13197 );
    nor g10883 ( n6893 , n9807 , n1293 );
    and g10884 ( n9508 , n13535 , n13579 );
    not g10885 ( n12953 , n1843 );
    or g10886 ( n530 , n1805 , n10362 );
    or g10887 ( n10732 , n10834 , n8810 );
    and g10888 ( n6298 , n4527 , n12738 );
    and g10889 ( n943 , n10357 , n9143 );
    and g10890 ( n8110 , n8569 , n5949 );
    not g10891 ( n13952 , n230 );
    and g10892 ( n7380 , n6854 , n4623 );
    and g10893 ( n1256 , n8020 , n8415 );
    nor g10894 ( n8729 , n8404 , n10480 );
    and g10895 ( n3939 , n8697 , n2613 );
    or g10896 ( n7078 , n7426 , n1674 );
    not g10897 ( n9654 , n8044 );
    and g10898 ( n3397 , n3743 , n12668 );
    and g10899 ( n6733 , n4690 , n11801 );
    not g10900 ( n6607 , n9846 );
    and g10901 ( n13369 , n10458 , n1290 );
    or g10902 ( n11728 , n7418 , n2198 );
    and g10903 ( n12969 , n14351 , n4727 );
    and g10904 ( n4729 , n79 , n11067 );
    nor g10905 ( n9639 , n14419 , n989 );
    and g10906 ( n10095 , n6625 , n370 );
    or g10907 ( n12077 , n11086 , n10552 );
    or g10908 ( n2697 , n9269 , n2305 );
    not g10909 ( n9231 , n5944 );
    and g10910 ( n11939 , n2942 , n1990 );
    and g10911 ( n14002 , n3277 , n6149 );
    and g10912 ( n11790 , n776 , n11588 );
    and g10913 ( n6274 , n3989 , n6660 );
    or g10914 ( n11540 , n11620 , n981 );
    and g10915 ( n8879 , n12531 , n5453 );
    and g10916 ( n3603 , n3130 , n6081 );
    or g10917 ( n10509 , n5406 , n4850 );
    nor g10918 ( n14116 , n1480 , n3685 );
    and g10919 ( n2485 , n2445 , n2805 );
    and g10920 ( n3494 , n7211 , n840 );
    or g10921 ( n12222 , n4876 , n3821 );
    nor g10922 ( n3302 , n11581 , n7702 );
    nor g10923 ( n2928 , n3546 , n5247 );
    nor g10924 ( n1468 , n4897 , n3694 );
    or g10925 ( n8773 , n5891 , n4520 );
    and g10926 ( n8918 , n8250 , n4208 );
    not g10927 ( n8825 , n4777 );
    and g10928 ( n4677 , n200 , n1819 );
    nor g10929 ( n9205 , n6971 , n10588 );
    and g10930 ( n3580 , n7060 , n12416 );
    not g10931 ( n2370 , n5504 );
    or g10932 ( n1901 , n647 , n8465 );
    or g10933 ( n7266 , n14286 , n3893 );
    nor g10934 ( n554 , n11975 , n12143 );
    or g10935 ( n2819 , n11183 , n10643 );
    or g10936 ( n5689 , n4340 , n4591 );
    and g10937 ( n12427 , n13359 , n4432 );
    and g10938 ( n12267 , n9890 , n12767 );
    and g10939 ( n13089 , n5279 , n4176 );
    or g10940 ( n12163 , n12759 , n13931 );
    or g10941 ( n10181 , n4631 , n1259 );
    or g10942 ( n5980 , n13466 , n1702 );
    or g10943 ( n4701 , n3088 , n10874 );
    and g10944 ( n4958 , n2682 , n12688 );
    and g10945 ( n5105 , n12918 , n4934 );
    or g10946 ( n408 , n511 , n1987 );
    and g10947 ( n8778 , n3672 , n11170 );
    nor g10948 ( n6613 , n7120 , n4348 );
    not g10949 ( n8458 , n4550 );
    or g10950 ( n4031 , n14166 , n11533 );
    or g10951 ( n6026 , n3088 , n11872 );
    or g10952 ( n2933 , n6323 , n11187 );
    or g10953 ( n10997 , n8964 , n13131 );
    and g10954 ( n10553 , n4261 , n10550 );
    or g10955 ( n11287 , n12401 , n13267 );
    or g10956 ( n11197 , n9403 , n13841 );
    or g10957 ( n5382 , n10224 , n10273 );
    and g10958 ( n2814 , n2445 , n10385 );
    not g10959 ( n8007 , n11428 );
    and g10960 ( n3757 , n5229 , n2679 );
    and g10961 ( n1830 , n13240 , n2595 );
    and g10962 ( n1717 , n11213 , n14257 );
    or g10963 ( n14008 , n9229 , n10473 );
    not g10964 ( n9564 , n6657 );
    and g10965 ( n5798 , n13407 , n2745 );
    or g10966 ( n12182 , n4925 , n9916 );
    and g10967 ( n4777 , n12658 , n482 );
    not g10968 ( n231 , n5871 );
    or g10969 ( n10858 , n7667 , n10147 );
    and g10970 ( n14379 , n14373 , n7574 );
    and g10971 ( n3451 , n8453 , n7787 );
    not g10972 ( n4765 , n8487 );
    not g10973 ( n2820 , n3356 );
    not g10974 ( n4486 , n1120 );
    or g10975 ( n14079 , n13005 , n9900 );
    not g10976 ( n10648 , n1109 );
    or g10977 ( n583 , n12020 , n403 );
    and g10978 ( n5674 , n3332 , n12300 );
    or g10979 ( n10476 , n14401 , n9722 );
    or g10980 ( n7858 , n8172 , n5843 );
    or g10981 ( n11007 , n2181 , n10800 );
    not g10982 ( n10331 , n4847 );
    not g10983 ( n481 , n7120 );
    and g10984 ( n10162 , n718 , n11265 );
    and g10985 ( n11856 , n9069 , n1058 );
    nor g10986 ( n4152 , n1348 , n12310 );
    or g10987 ( n3187 , n9864 , n10749 );
    not g10988 ( n9507 , n2320 );
    and g10989 ( n765 , n7768 , n9593 );
    not g10990 ( n12039 , n5525 );
    not g10991 ( n8431 , n13734 );
    or g10992 ( n7333 , n12494 , n3723 );
    not g10993 ( n13220 , n7875 );
    not g10994 ( n1332 , n6703 );
    and g10995 ( n6820 , n1772 , n1589 );
    or g10996 ( n3113 , n5634 , n8552 );
    and g10997 ( n7603 , n7961 , n11672 );
    and g10998 ( n1511 , n8412 , n5866 );
    and g10999 ( n11226 , n3635 , n4496 );
    or g11000 ( n9986 , n13080 , n4838 );
    or g11001 ( n978 , n10294 , n14279 );
    or g11002 ( n7182 , n10300 , n1108 );
    nor g11003 ( n11802 , n7418 , n13661 );
    nor g11004 ( n2352 , n2016 , n11114 );
    or g11005 ( n5556 , n7697 , n11689 );
    and g11006 ( n5300 , n4433 , n7313 );
    and g11007 ( n13620 , n9650 , n12698 );
    nor g11008 ( n4133 , n7362 , n7197 );
    and g11009 ( n14294 , n1047 , n6363 );
    and g11010 ( n2648 , n5948 , n4886 );
    not g11011 ( n11832 , n12949 );
    nor g11012 ( n9207 , n12757 , n8138 );
    or g11013 ( n7629 , n850 , n6450 );
    and g11014 ( n5590 , n2224 , n5929 );
    or g11015 ( n9855 , n8897 , n9578 );
    or g11016 ( n8843 , n2272 , n3162 );
    or g11017 ( n12346 , n7697 , n6598 );
    or g11018 ( n1659 , n4357 , n11721 );
    or g11019 ( n1508 , n10619 , n11776 );
    or g11020 ( n1664 , n89 , n339 );
    nor g11021 ( n8900 , n7145 , n352 );
    or g11022 ( n11793 , n12900 , n2164 );
    nor g11023 ( n9922 , n4608 , n11446 );
    and g11024 ( n4392 , n4932 , n13167 );
    or g11025 ( n3809 , n7744 , n2065 );
    or g11026 ( n8095 , n1494 , n13182 );
    not g11027 ( n11153 , n9994 );
    and g11028 ( n8239 , n5312 , n9844 );
    and g11029 ( n11501 , n3635 , n11834 );
    or g11030 ( n10584 , n12549 , n13592 );
    and g11031 ( n8851 , n1788 , n9227 );
    and g11032 ( n10569 , n10330 , n12235 );
    and g11033 ( n3706 , n10357 , n7045 );
    nor g11034 ( n5128 , n2808 , n6673 );
    not g11035 ( n1047 , n11474 );
    nor g11036 ( n14297 , n4829 , n2660 );
    and g11037 ( n1740 , n718 , n1970 );
    or g11038 ( n1160 , n8452 , n11622 );
    not g11039 ( n1660 , n4325 );
    or g11040 ( n8609 , n1261 , n10028 );
    or g11041 ( n12726 , n6111 , n8375 );
    or g11042 ( n12555 , n1821 , n6927 );
    or g11043 ( n4444 , n6519 , n6489 );
    not g11044 ( n3875 , n5160 );
    and g11045 ( n13566 , n1802 , n5171 );
    not g11046 ( n14135 , n13560 );
    not g11047 ( n7267 , n10322 );
    or g11048 ( n306 , n5587 , n2809 );
    or g11049 ( n13679 , n839 , n13540 );
    nor g11050 ( n7577 , n5509 , n10244 );
    nor g11051 ( n6721 , n7696 , n1719 );
    and g11052 ( n2559 , n7832 , n1694 );
    or g11053 ( n8292 , n11551 , n12851 );
    or g11054 ( n8385 , n1576 , n9079 );
    not g11055 ( n3870 , n9608 );
    and g11056 ( n5183 , n350 , n12308 );
    and g11057 ( n4892 , n12935 , n2746 );
    and g11058 ( n2528 , n7079 , n2711 );
    or g11059 ( n3317 , n6595 , n6639 );
    or g11060 ( n11214 , n7684 , n11174 );
    and g11061 ( n2689 , n6016 , n13965 );
    or g11062 ( n5655 , n9423 , n5037 );
    not g11063 ( n12037 , n6007 );
    and g11064 ( n14411 , n11163 , n11760 );
    nor g11065 ( n12965 , n11492 , n6189 );
    not g11066 ( n13420 , n6680 );
    or g11067 ( n12171 , n6909 , n4154 );
    not g11068 ( n1127 , n5294 );
    nor g11069 ( n3889 , n6030 , n13060 );
    or g11070 ( n9536 , n8726 , n5267 );
    not g11071 ( n8980 , n4891 );
    not g11072 ( n12259 , n4210 );
    nor g11073 ( n6443 , n14075 , n11766 );
    and g11074 ( n12341 , n9853 , n4441 );
    or g11075 ( n6896 , n3093 , n11799 );
    or g11076 ( n1052 , n1202 , n3494 );
    or g11077 ( n5040 , n7219 , n4369 );
    or g11078 ( n4006 , n3559 , n14275 );
    or g11079 ( n13726 , n13108 , n4281 );
    not g11080 ( n9206 , n13814 );
    and g11081 ( n3482 , n11336 , n5660 );
    nor g11082 ( n3798 , n6700 , n8390 );
    nor g11083 ( n13168 , n13875 , n11977 );
    and g11084 ( n11491 , n13078 , n12557 );
    and g11085 ( n12236 , n11867 , n4557 );
    and g11086 ( n8356 , n3526 , n7650 );
    nor g11087 ( n7843 , n7683 , n8857 );
    nor g11088 ( n7475 , n10289 , n7094 );
    nor g11089 ( n11566 , n12323 , n4419 );
    or g11090 ( n7225 , n7697 , n6837 );
    not g11091 ( n7684 , n382 );
    and g11092 ( n11475 , n7057 , n493 );
    or g11093 ( n1656 , n11262 , n8799 );
    and g11094 ( n3200 , n11316 , n11773 );
    or g11095 ( n9368 , n10323 , n4002 );
    nor g11096 ( n14271 , n9423 , n9694 );
    or g11097 ( n5473 , n10245 , n9710 );
    and g11098 ( n12571 , n8453 , n10328 );
    and g11099 ( n8601 , n12460 , n9896 );
    not g11100 ( n8767 , n3765 );
    or g11101 ( n5446 , n3164 , n3437 );
    not g11102 ( n6507 , n13181 );
    and g11103 ( n7273 , n1772 , n6175 );
    or g11104 ( n639 , n5891 , n2981 );
    or g11105 ( n8421 , n2025 , n5176 );
    nor g11106 ( n1945 , n4424 , n13013 );
    or g11107 ( n3805 , n3445 , n9990 );
    or g11108 ( n11085 , n6891 , n9322 );
    or g11109 ( n3595 , n12019 , n4462 );
    and g11110 ( n4611 , n3766 , n4745 );
    and g11111 ( n5394 , n8412 , n13111 );
    nor g11112 ( n13505 , n1628 , n312 );
    or g11113 ( n3265 , n8332 , n6244 );
    and g11114 ( n13772 , n10556 , n968 );
    or g11115 ( n2297 , n12139 , n363 );
    and g11116 ( n11707 , n4244 , n8878 );
    not g11117 ( n2996 , n14135 );
    or g11118 ( n4588 , n9353 , n4326 );
    and g11119 ( n9558 , n7419 , n9260 );
    or g11120 ( n11895 , n2057 , n4030 );
    or g11121 ( n1691 , n7430 , n12370 );
    and g11122 ( n13646 , n1431 , n11424 );
    and g11123 ( n4350 , n9885 , n8567 );
    or g11124 ( n1483 , n7212 , n10569 );
    nor g11125 ( n8860 , n4741 , n7512 );
    not g11126 ( n8856 , n10617 );
    and g11127 ( n3250 , n3526 , n5078 );
    nor g11128 ( n6634 , n9529 , n9185 );
    or g11129 ( n5998 , n4925 , n8279 );
    nor g11130 ( n7965 , n6088 , n10554 );
    not g11131 ( n3766 , n5618 );
    and g11132 ( n10910 , n13240 , n11119 );
    and g11133 ( n1363 , n11008 , n2433 );
    and g11134 ( n7409 , n7284 , n13985 );
    and g11135 ( n3180 , n309 , n8686 );
    or g11136 ( n13341 , n1538 , n14347 );
    or g11137 ( n698 , n4898 , n14230 );
    and g11138 ( n6092 , n14465 , n198 );
    or g11139 ( n6183 , n11105 , n7158 );
    not g11140 ( n5807 , n2383 );
    and g11141 ( n13848 , n11020 , n8193 );
    or g11142 ( n2439 , n12549 , n10048 );
    nor g11143 ( n4629 , n12765 , n6828 );
    or g11144 ( n436 , n12020 , n10433 );
    nor g11145 ( n7437 , n1480 , n11427 );
    and g11146 ( n12881 , n1428 , n11786 );
    not g11147 ( n1044 , n409 );
    or g11148 ( n12251 , n13806 , n14190 );
    and g11149 ( n8426 , n3526 , n11279 );
    and g11150 ( n14103 , n4574 , n3838 );
    nor g11151 ( n13334 , n13376 , n11209 );
    and g11152 ( n7987 , n4300 , n7017 );
    not g11153 ( n11117 , n11933 );
    nor g11154 ( n13422 , n8825 , n424 );
    or g11155 ( n12495 , n4899 , n1825 );
    and g11156 ( n12805 , n6135 , n771 );
    and g11157 ( n2943 , n13367 , n3745 );
    and g11158 ( n10265 , n129 , n5232 );
    and g11159 ( n380 , n6192 , n11004 );
    or g11160 ( n2153 , n11303 , n2277 );
    and g11161 ( n8734 , n5275 , n2404 );
    and g11162 ( n11820 , n13850 , n13883 );
    and g11163 ( n7394 , n12521 , n10168 );
    nor g11164 ( n6075 , n4174 , n3528 );
    and g11165 ( n831 , n10820 , n3884 );
    and g11166 ( n127 , n2064 , n11794 );
    and g11167 ( n12381 , n13525 , n12629 );
    or g11168 ( n1800 , n227 , n3818 );
    nor g11169 ( n266 , n2086 , n3239 );
    nor g11170 ( n13630 , n2218 , n10014 );
    and g11171 ( n1081 , n2082 , n13927 );
    or g11172 ( n11564 , n6271 , n3898 );
    or g11173 ( n5465 , n10323 , n9908 );
    not g11174 ( n14373 , n11715 );
    and g11175 ( n3260 , n10025 , n456 );
    and g11176 ( n9484 , n7370 , n369 );
    or g11177 ( n10722 , n12211 , n7320 );
    or g11178 ( n8478 , n7003 , n94 );
    nor g11179 ( n1092 , n8656 , n11233 );
    not g11180 ( n12827 , n5980 );
    or g11181 ( n4398 , n3886 , n1603 );
    and g11182 ( n5262 , n8769 , n1789 );
    or g11183 ( n13579 , n5483 , n3069 );
    or g11184 ( n5020 , n10394 , n5345 );
    or g11185 ( n2745 , n2518 , n54 );
    and g11186 ( n9958 , n10338 , n1021 );
    and g11187 ( n9006 , n9265 , n14395 );
    and g11188 ( n7546 , n10231 , n7781 );
    not g11189 ( n11990 , n5354 );
    and g11190 ( n1316 , n13421 , n10911 );
    nor g11191 ( n7799 , n12800 , n9097 );
    and g11192 ( n8563 , n7211 , n11643 );
    nor g11193 ( n7557 , n4439 , n8127 );
    not g11194 ( n14357 , n7272 );
    and g11195 ( n10422 , n6167 , n8827 );
    not g11196 ( n8210 , n12746 );
    and g11197 ( n5194 , n3247 , n542 );
    and g11198 ( n7947 , n5071 , n1734 );
    or g11199 ( n13023 , n12131 , n9942 );
    or g11200 ( n2339 , n10351 , n8268 );
    and g11201 ( n9542 , n12960 , n9261 );
    or g11202 ( n4980 , n12500 , n1893 );
    or g11203 ( n14334 , n8828 , n5119 );
    or g11204 ( n8211 , n8277 , n4740 );
    and g11205 ( n6118 , n4018 , n1560 );
    and g11206 ( n7445 , n2006 , n9794 );
    or g11207 ( n12278 , n5225 , n9977 );
    and g11208 ( n10598 , n6531 , n8700 );
    not g11209 ( n2091 , n11143 );
    not g11210 ( n533 , n230 );
    or g11211 ( n562 , n12100 , n8145 );
    nor g11212 ( n1323 , n48 , n13009 );
    or g11213 ( n4176 , n390 , n4867 );
    nor g11214 ( n9395 , n6788 , n13669 );
    and g11215 ( n9337 , n12986 , n12115 );
    or g11216 ( n2621 , n3132 , n13673 );
    nor g11217 ( n9253 , n8592 , n3524 );
    or g11218 ( n12541 , n5833 , n12853 );
    and g11219 ( n595 , n11142 , n5154 );
    nor g11220 ( n3844 , n5990 , n11299 );
    and g11221 ( n5351 , n2224 , n13184 );
    or g11222 ( n4146 , n10079 , n11756 );
    or g11223 ( n2951 , n13037 , n1027 );
    or g11224 ( n2481 , n6629 , n5010 );
    and g11225 ( n8454 , n11614 , n13617 );
    and g11226 ( n1676 , n13426 , n9793 );
    or g11227 ( n8347 , n2908 , n12044 );
    or g11228 ( n519 , n6090 , n8165 );
    nor g11229 ( n467 , n7004 , n8841 );
    and g11230 ( n14022 , n13367 , n1351 );
    and g11231 ( n7550 , n2473 , n3265 );
    or g11232 ( n11380 , n584 , n2865 );
    nor g11233 ( n9440 , n12084 , n9277 );
    or g11234 ( n3261 , n2510 , n4143 );
    or g11235 ( n6285 , n3126 , n6684 );
    or g11236 ( n13411 , n1538 , n12135 );
    not g11237 ( n5333 , n12084 );
    and g11238 ( n3441 , n12455 , n1940 );
    or g11239 ( n9679 , n2002 , n11933 );
    or g11240 ( n5867 , n10560 , n1824 );
    nor g11241 ( n13300 , n7407 , n13274 );
    and g11242 ( n78 , n13700 , n12972 );
    or g11243 ( n2887 , n13706 , n1363 );
    and g11244 ( n7713 , n8427 , n1668 );
    or g11245 ( n13818 , n4205 , n7622 );
    and g11246 ( n389 , n2061 , n7913 );
    and g11247 ( n4736 , n8043 , n7169 );
    not g11248 ( n316 , n6426 );
    and g11249 ( n11751 , n6537 , n5832 );
    and g11250 ( n9003 , n13700 , n12364 );
    or g11251 ( n9505 , n8277 , n3857 );
    nor g11252 ( n11994 , n2752 , n10700 );
    or g11253 ( n14007 , n504 , n7440 );
    and g11254 ( n770 , n8213 , n44 );
    or g11255 ( n8472 , n6937 , n10470 );
    not g11256 ( n10624 , n10775 );
    and g11257 ( n13703 , n4929 , n14013 );
    and g11258 ( n5906 , n13342 , n8461 );
    and g11259 ( n8966 , n4788 , n13998 );
    or g11260 ( n12557 , n12576 , n1238 );
    and g11261 ( n254 , n13656 , n131 );
    and g11262 ( n4772 , n1125 , n13299 );
    or g11263 ( n7141 , n11676 , n8780 );
    nor g11264 ( n5368 , n11325 , n9318 );
    or g11265 ( n5888 , n3777 , n315 );
    not g11266 ( n5634 , n8486 );
    or g11267 ( n9607 , n6730 , n9040 );
    and g11268 ( n6687 , n2006 , n6710 );
    and g11269 ( n13704 , n10374 , n11637 );
    or g11270 ( n14280 , n3164 , n10422 );
    or g11271 ( n5260 , n2784 , n8947 );
    not g11272 ( n5265 , n585 );
    not g11273 ( n13324 , n5333 );
    and g11274 ( n746 , n1802 , n7184 );
    and g11275 ( n2797 , n11503 , n6107 );
    nor g11276 ( n6158 , n2218 , n1219 );
    and g11277 ( n7265 , n1776 , n7927 );
    and g11278 ( n12256 , n11028 , n3422 );
    and g11279 ( n5802 , n11336 , n10052 );
    nor g11280 ( n13893 , n14058 , n5513 );
    not g11281 ( n458 , n4373 );
    nor g11282 ( n1865 , n4284 , n4272 );
    or g11283 ( n7493 , n9353 , n1487 );
    and g11284 ( n4077 , n11008 , n1752 );
    and g11285 ( n6127 , n9571 , n3051 );
    and g11286 ( n3214 , n636 , n12171 );
    nor g11287 ( n10876 , n10637 , n1945 );
    and g11288 ( n7960 , n5475 , n12825 );
    and g11289 ( n3010 , n1047 , n2893 );
    nor g11290 ( n6914 , n48 , n1121 );
    not g11291 ( n2531 , n382 );
    nor g11292 ( n709 , n8592 , n1707 );
    or g11293 ( n13211 , n839 , n11172 );
    and g11294 ( n6123 , n12909 , n12358 );
    not g11295 ( n5562 , n7600 );
    nor g11296 ( n4247 , n10648 , n6582 );
    not g11297 ( n10593 , n2370 );
    or g11298 ( n6176 , n5562 , n7471 );
    not g11299 ( n3710 , n871 );
    not g11300 ( n3561 , n8550 );
    or g11301 ( n515 , n8828 , n2883 );
    and g11302 ( n14353 , n4358 , n1808 );
    or g11303 ( n8429 , n2901 , n6761 );
    and g11304 ( n13846 , n3370 , n910 );
    or g11305 ( n13027 , n7359 , n5366 );
    not g11306 ( n8544 , n4216 );
    not g11307 ( n7842 , n8576 );
    or g11308 ( n1748 , n11837 , n2454 );
    and g11309 ( n1907 , n12421 , n12410 );
    not g11310 ( n11839 , n1010 );
    and g11311 ( n4890 , n4422 , n5230 );
    or g11312 ( n12585 , n480 , n10819 );
    or g11313 ( n7956 , n492 , n8132 );
    and g11314 ( n10577 , n12013 , n11703 );
    or g11315 ( n3575 , n228 , n5353 );
    or g11316 ( n9393 , n6857 , n12606 );
    nor g11317 ( n14126 , n8217 , n7661 );
    or g11318 ( n11651 , n10309 , n2603 );
    and g11319 ( n2081 , n4359 , n6514 );
    and g11320 ( n2108 , n8849 , n9925 );
    not g11321 ( n1473 , n5300 );
    and g11322 ( n14131 , n1857 , n1816 );
    or g11323 ( n7793 , n28 , n6339 );
    or g11324 ( n13642 , n7430 , n7180 );
    and g11325 ( n10444 , n687 , n13401 );
    or g11326 ( n3659 , n3088 , n13651 );
    and g11327 ( n7794 , n12461 , n13079 );
    and g11328 ( n3293 , n6838 , n13581 );
    not g11329 ( n7912 , n9371 );
    nor g11330 ( n2733 , n6731 , n4059 );
    and g11331 ( n9405 , n14227 , n8248 );
    not g11332 ( n1495 , n407 );
    not g11333 ( n13069 , n13458 );
    and g11334 ( n5947 , n9650 , n5219 );
    not g11335 ( n976 , n238 );
    or g11336 ( n5417 , n12500 , n1715 );
    and g11337 ( n5933 , n2461 , n10563 );
    or g11338 ( n10304 , n1875 , n3700 );
    or g11339 ( n9859 , n10871 , n6847 );
    and g11340 ( n14448 , n687 , n10155 );
    and g11341 ( n5516 , n5011 , n11409 );
    and g11342 ( n2435 , n5092 , n3087 );
    nor g11343 ( n9841 , n1473 , n4152 );
    and g11344 ( n5844 , n8965 , n8012 );
    and g11345 ( n5431 , n8238 , n7513 );
    and g11346 ( n1315 , n12449 , n5556 );
    or g11347 ( n11397 , n10234 , n9347 );
    or g11348 ( n4656 , n6480 , n3263 );
    and g11349 ( n7734 , n432 , n4588 );
    and g11350 ( n5907 , n6697 , n14083 );
    and g11351 ( n9911 , n7053 , n12967 );
    and g11352 ( n13347 , n14109 , n7637 );
    and g11353 ( n11031 , n8768 , n10202 );
    nor g11354 ( n6210 , n2866 , n12736 );
    not g11355 ( n13297 , n6113 );
    and g11356 ( n4281 , n222 , n3282 );
    or g11357 ( n2076 , n8151 , n1221 );
    or g11358 ( n2993 , n11647 , n14089 );
    or g11359 ( n13664 , n10449 , n4506 );
    and g11360 ( n609 , n7997 , n7241 );
    nor g11361 ( n1372 , n151 , n2688 );
    and g11362 ( n14417 , n9297 , n436 );
    not g11363 ( n1494 , n14154 );
    and g11364 ( n1171 , n80 , n257 );
    nor g11365 ( n9969 , n2016 , n7030 );
    nor g11366 ( n2540 , n3445 , n9213 );
    nor g11367 ( n12920 , n11489 , n13260 );
    nor g11368 ( n7921 , n3882 , n13508 );
    nor g11369 ( n11671 , n7245 , n8645 );
    and g11370 ( n10141 , n4358 , n2456 );
    nor g11371 ( n7153 , n13399 , n13644 );
    or g11372 ( n13157 , n3125 , n12490 );
    and g11373 ( n14346 , n13520 , n9588 );
    or g11374 ( n6369 , n10309 , n14284 );
    not g11375 ( n3354 , n10994 );
    and g11376 ( n13629 , n5458 , n13653 );
    and g11377 ( n1696 , n14351 , n12544 );
    and g11378 ( n2101 , n12802 , n1317 );
    nor g11379 ( n13400 , n11094 , n789 );
    and g11380 ( n12118 , n1354 , n14486 );
    or g11381 ( n284 , n163 , n707 );
    or g11382 ( n8160 , n12543 , n5431 );
    or g11383 ( n11203 , n7436 , n7764 );
    or g11384 ( n10558 , n11303 , n12685 );
    or g11385 ( n10690 , n2017 , n11027 );
    and g11386 ( n3311 , n14373 , n2900 );
    or g11387 ( n6663 , n9620 , n13307 );
    or g11388 ( n610 , n10294 , n6602 );
    and g11389 ( n1190 , n7187 , n3316 );
    or g11390 ( n1346 , n28 , n5457 );
    and g11391 ( n5974 , n8163 , n10801 );
    and g11392 ( n6538 , n3169 , n14007 );
    and g11393 ( n11274 , n12455 , n4685 );
    or g11394 ( n2288 , n3559 , n5798 );
    or g11395 ( n10417 , n412 , n6931 );
    and g11396 ( n6357 , n11244 , n1881 );
    or g11397 ( n14418 , n3888 , n774 );
    and g11398 ( n12515 , n12449 , n6241 );
    and g11399 ( n12931 , n8923 , n377 );
    and g11400 ( n14264 , n1854 , n2837 );
    not g11401 ( n10609 , n2967 );
    not g11402 ( n4534 , n4646 );
    or g11403 ( n12204 , n7912 , n10664 );
    and g11404 ( n13042 , n8569 , n2713 );
    or g11405 ( n11603 , n9620 , n14270 );
    or g11406 ( n8487 , n8746 , n8550 );
    nor g11407 ( n9927 , n12968 , n1460 );
    nor g11408 ( n5902 , n8942 , n8121 );
    not g11409 ( n1669 , n12394 );
    or g11410 ( n1555 , n1701 , n6655 );
    or g11411 ( n9161 , n10857 , n2814 );
    and g11412 ( n7132 , n11590 , n6430 );
    not g11413 ( n10224 , n8735 );
    not g11414 ( n13977 , n2973 );
    not g11415 ( n3527 , n2472 );
    and g11416 ( n11673 , n3942 , n11881 );
    and g11417 ( n805 , n3846 , n6382 );
    not g11418 ( n2747 , n2484 );
    and g11419 ( n7232 , n12018 , n4941 );
    not g11420 ( n1254 , n2906 );
    nor g11421 ( n10733 , n3394 , n2123 );
    or g11422 ( n13026 , n791 , n9996 );
    nor g11423 ( n3857 , n4637 , n13062 );
    and g11424 ( n10370 , n2082 , n2683 );
    or g11425 ( n5636 , n10089 , n2219 );
    and g11426 ( n3883 , n4346 , n13679 );
    or g11427 ( n11006 , n10154 , n10699 );
    and g11428 ( n10689 , n9745 , n13417 );
    nor g11429 ( n4836 , n239 , n10387 );
    and g11430 ( n8423 , n5489 , n11035 );
    nor g11431 ( n3581 , n12568 , n12010 );
    and g11432 ( n1168 , n14150 , n572 );
    not g11433 ( n12528 , n10945 );
    or g11434 ( n13344 , n7888 , n1665 );
    nor g11435 ( n3560 , n12957 , n13657 );
    or g11436 ( n12566 , n10234 , n13328 );
    or g11437 ( n2047 , n7212 , n3887 );
    nor g11438 ( n3450 , n8021 , n8679 );
    not g11439 ( n7060 , n4490 );
    or g11440 ( n1554 , n9804 , n1720 );
    or g11441 ( n10274 , n4033 , n2656 );
    not g11442 ( n1138 , n12069 );
    nor g11443 ( n5970 , n2000 , n2541 );
    and g11444 ( n10074 , n2961 , n11295 );
    and g11445 ( n2429 , n12461 , n3689 );
    or g11446 ( n11579 , n2518 , n9569 );
    and g11447 ( n12264 , n5317 , n14004 );
    or g11448 ( n1909 , n3273 , n524 );
    not g11449 ( n6326 , n6248 );
    and g11450 ( n9118 , n8801 , n2698 );
    and g11451 ( n4938 , n2643 , n5898 );
    or g11452 ( n11659 , n4822 , n8029 );
    or g11453 ( n1761 , n6867 , n3498 );
    and g11454 ( n7641 , n2983 , n6878 );
    nor g11455 ( n7377 , n8798 , n13340 );
    or g11456 ( n5963 , n9747 , n11031 );
    or g11457 ( n4056 , n5647 , n13343 );
    or g11458 ( n1845 , n7700 , n7259 );
    not g11459 ( n850 , n7322 );
    not g11460 ( n3445 , n9580 );
    and g11461 ( n12006 , n11240 , n4008 );
    and g11462 ( n10346 , n12506 , n5221 );
    or g11463 ( n1099 , n1198 , n12946 );
    and g11464 ( n6534 , n13209 , n10697 );
    or g11465 ( n11957 , n13537 , n8133 );
    and g11466 ( n11670 , n10922 , n1781 );
    or g11467 ( n8141 , n5625 , n10738 );
    nor g11468 ( n7160 , n8798 , n6121 );
    and g11469 ( n13777 , n7057 , n7545 );
    or g11470 ( n6996 , n317 , n10689 );
    and g11471 ( n5050 , n3923 , n6402 );
    or g11472 ( n13652 , n5762 , n4011 );
    nor g11473 ( n10305 , n11040 , n12165 );
    not g11474 ( n1011 , n8204 );
    or g11475 ( n11062 , n6537 , n9921 );
    nor g11476 ( n537 , n585 , n14023 );
    or g11477 ( n12300 , n8828 , n13205 );
    nor g11478 ( n10257 , n6971 , n5573 );
    nor g11479 ( n5208 , n8216 , n7925 );
    or g11480 ( n2714 , n839 , n8208 );
    or g11481 ( n2037 , n5641 , n1402 );
    or g11482 ( n11708 , n12211 , n3336 );
    and g11483 ( n2397 , n12620 , n13896 );
    and g11484 ( n3864 , n14351 , n9681 );
    or g11485 ( n3472 , n4821 , n3772 );
    nor g11486 ( n2189 , n4135 , n7210 );
    not g11487 ( n13083 , n11788 );
    not g11488 ( n6205 , n13234 );
    not g11489 ( n8975 , n10736 );
    and g11490 ( n10395 , n4601 , n14249 );
    or g11491 ( n5134 , n12324 , n4475 );
    and g11492 ( n13343 , n12185 , n11819 );
    and g11493 ( n4137 , n6311 , n11601 );
    and g11494 ( n7664 , n13103 , n11037 );
    and g11495 ( n11115 , n10647 , n7718 );
    not g11496 ( n13310 , n10629 );
    and g11497 ( n8169 , n7670 , n7495 );
    or g11498 ( n1808 , n2747 , n8879 );
    or g11499 ( n5274 , n781 , n726 );
    or g11500 ( n140 , n8821 , n13895 );
    and g11501 ( n12906 , n8183 , n7350 );
    and g11502 ( n6573 , n3861 , n13803 );
    and g11503 ( n11343 , n3449 , n14204 );
    not g11504 ( n4299 , n10897 );
    or g11505 ( n7726 , n1223 , n2081 );
    or g11506 ( n6356 , n3076 , n5282 );
    and g11507 ( n11451 , n9191 , n8883 );
    not g11508 ( n6937 , n12829 );
    and g11509 ( n7847 , n9238 , n6936 );
    and g11510 ( n12517 , n7673 , n11952 );
    and g11511 ( n1381 , n13236 , n927 );
    not g11512 ( n1946 , n8649 );
    or g11513 ( n8869 , n3011 , n9881 );
    or g11514 ( n8647 , n5046 , n394 );
    or g11515 ( n4745 , n13537 , n11032 );
    and g11516 ( n12076 , n405 , n7490 );
    and g11517 ( n8208 , n11495 , n5963 );
    nor g11518 ( n9968 , n12403 , n199 );
    or g11519 ( n8207 , n4876 , n7328 );
    not g11520 ( n3418 , n8521 );
    or g11521 ( n1536 , n6350 , n3591 );
    not g11522 ( n8672 , n11975 );
    and g11523 ( n4584 , n898 , n8331 );
    and g11524 ( n4511 , n13555 , n11923 );
    or g11525 ( n2491 , n14435 , n13490 );
    nor g11526 ( n9185 , n6905 , n3414 );
    not g11527 ( n442 , n3918 );
    and g11528 ( n514 , n4018 , n10877 );
    and g11529 ( n9437 , n12614 , n12354 );
    and g11530 ( n13678 , n2330 , n4009 );
    or g11531 ( n11294 , n11011 , n2389 );
    and g11532 ( n10540 , n14227 , n4390 );
    or g11533 ( n3073 , n3161 , n2824 );
    and g11534 ( n7101 , n3724 , n14496 );
    or g11535 ( n10951 , n2645 , n1770 );
    and g11536 ( n9109 , n11503 , n2208 );
    not g11537 ( n5641 , n3021 );
    not g11538 ( n31 , n14134 );
    and g11539 ( n7785 , n8147 , n3865 );
    nor g11540 ( n8057 , n13248 , n1257 );
    not g11541 ( n4549 , n6742 );
    and g11542 ( n11331 , n12168 , n12192 );
    nor g11543 ( n10480 , n10638 , n592 );
    or g11544 ( n6842 , n2686 , n8011 );
    or g11545 ( n10277 , n13698 , n10758 );
    nor g11546 ( n7954 , n4682 , n8311 );
    or g11547 ( n8062 , n10825 , n1727 );
    not g11548 ( n6596 , n10204 );
    and g11549 ( n10069 , n6067 , n4769 );
    and g11550 ( n2136 , n3846 , n1792 );
    and g11551 ( n13583 , n4445 , n12526 );
    and g11552 ( n43 , n13338 , n119 );
    or g11553 ( n6973 , n12351 , n9086 );
    or g11554 ( n2421 , n817 , n936 );
    and g11555 ( n9241 , n6130 , n4058 );
    and g11556 ( n4719 , n8047 , n4158 );
    and g11557 ( n331 , n13755 , n9978 );
    or g11558 ( n1658 , n12149 , n166 );
    nor g11559 ( n5164 , n2932 , n9408 );
    not g11560 ( n9289 , n9959 );
    or g11561 ( n10842 , n13118 , n881 );
    not g11562 ( n3607 , n2497 );
    or g11563 ( n7479 , n9931 , n2922 );
    and g11564 ( n5953 , n10134 , n3553 );
    and g11565 ( n12374 , n9190 , n2649 );
    or g11566 ( n14219 , n3895 , n760 );
    or g11567 ( n6161 , n77 , n2160 );
    not g11568 ( n2468 , n11120 );
    or g11569 ( n8749 , n8714 , n14480 );
    or g11570 ( n11653 , n11360 , n8745 );
    or g11571 ( n6569 , n7618 , n844 );
    and g11572 ( n1350 , n6167 , n3229 );
    and g11573 ( n1070 , n8768 , n7741 );
    or g11574 ( n9598 , n10394 , n8936 );
    or g11575 ( n5407 , n14435 , n13067 );
    or g11576 ( n4981 , n11704 , n12477 );
    or g11577 ( n12054 , n10461 , n11282 );
    and g11578 ( n3061 , n889 , n3925 );
    not g11579 ( n8480 , n11415 );
    nor g11580 ( n12356 , n11445 , n5978 );
    or g11581 ( n677 , n12149 , n3186 );
    nor g11582 ( n12643 , n5505 , n5824 );
    and g11583 ( n6818 , n231 , n8738 );
    or g11584 ( n377 , n28 , n11797 );
    and g11585 ( n12929 , n9650 , n10923 );
    nor g11586 ( n4458 , n4978 , n13140 );
    and g11587 ( n11524 , n9745 , n1810 );
    or g11588 ( n11019 , n2888 , n1315 );
    or g11589 ( n3310 , n12401 , n14487 );
    not g11590 ( n2412 , n8735 );
    nor g11591 ( n13616 , n5977 , n10029 );
    and g11592 ( n12919 , n10247 , n2035 );
    and g11593 ( n1704 , n11316 , n14305 );
    not g11594 ( n5507 , n382 );
    and g11595 ( n12640 , n2486 , n8411 );
    not g11596 ( n8513 , n4317 );
    not g11597 ( n4508 , n11055 );
    and g11598 ( n5614 , n3365 , n12090 );
    or g11599 ( n7150 , n1701 , n184 );
    and g11600 ( n8805 , n4690 , n4398 );
    and g11601 ( n1564 , n2158 , n13767 );
    and g11602 ( n5277 , n5240 , n5446 );
    not g11603 ( n11547 , n381 );
    or g11604 ( n9753 , n4739 , n8001 );
    or g11605 ( n984 , n10224 , n4209 );
    and g11606 ( n9923 , n4394 , n147 );
    or g11607 ( n4810 , n5710 , n6478 );
    not g11608 ( n7284 , n13139 );
    and g11609 ( n11699 , n8431 , n4246 );
    not g11610 ( n4213 , n8572 );
    or g11611 ( n10916 , n12130 , n2930 );
    nor g11612 ( n13986 , n1383 , n7981 );
    or g11613 ( n14076 , n14074 , n3130 );
    and g11614 ( n2509 , n8855 , n2110 );
    and g11615 ( n7655 , n13882 , n8214 );
    and g11616 ( n10507 , n7852 , n14121 );
    and g11617 ( n2749 , n12425 , n1903 );
    and g11618 ( n10796 , n12772 , n10790 );
    or g11619 ( n273 , n3914 , n8865 );
    not g11620 ( n7812 , n622 );
    and g11621 ( n141 , n8043 , n6766 );
    or g11622 ( n8827 , n11231 , n9106 );
    and g11623 ( n1340 , n309 , n14477 );
    or g11624 ( n2019 , n2908 , n6222 );
    or g11625 ( n13056 , n8881 , n9181 );
    and g11626 ( n6511 , n4358 , n7948 );
    or g11627 ( n3205 , n7812 , n1228 );
    and g11628 ( n12754 , n12039 , n13553 );
    and g11629 ( n5771 , n446 , n3917 );
    or g11630 ( n414 , n6867 , n9852 );
    not g11631 ( n1855 , n10750 );
    nor g11632 ( n10700 , n10309 , n11155 );
    or g11633 ( n4825 , n12622 , n2642 );
    and g11634 ( n12502 , n11316 , n6331 );
    or g11635 ( n4882 , n12295 , n4221 );
    not g11636 ( n6625 , n3440 );
    or g11637 ( n9002 , n4357 , n3663 );
    and g11638 ( n952 , n10209 , n5155 );
    and g11639 ( n1334 , n3561 , n12900 );
    or g11640 ( n12949 , n4887 , n6054 );
    or g11641 ( n1485 , n9229 , n13294 );
    or g11642 ( n8448 , n1051 , n8626 );
    and g11643 ( n2437 , n6898 , n6764 );
    or g11644 ( n7286 , n6867 , n2718 );
    or g11645 ( n2436 , n3125 , n7851 );
    or g11646 ( n7396 , n5861 , n7010 );
    not g11647 ( n11508 , n11453 );
    and g11648 ( n2084 , n9113 , n1343 );
    nor g11649 ( n7100 , n4174 , n12155 );
    and g11650 ( n4543 , n12741 , n845 );
    nor g11651 ( n6475 , n2236 , n3963 );
    and g11652 ( n2227 , n6157 , n13602 );
    and g11653 ( n907 , n12611 , n4910 );
    or g11654 ( n11959 , n13446 , n294 );
    and g11655 ( n7397 , n3271 , n2262 );
    and g11656 ( n10336 , n4300 , n5870 );
    or g11657 ( n7453 , n13016 , n12188 );
    not g11658 ( n6373 , n6264 );
    or g11659 ( n4360 , n10913 , n13028 );
    and g11660 ( n7541 , n13236 , n9730 );
    nor g11661 ( n7355 , n3132 , n12965 );
    or g11662 ( n6641 , n5986 , n13751 );
    and g11663 ( n8852 , n13421 , n10574 );
    nor g11664 ( n3619 , n11227 , n10157 );
    or g11665 ( n14497 , n10857 , n11219 );
    nor g11666 ( n9436 , n9967 , n13249 );
    and g11667 ( n3385 , n80 , n10149 );
    not g11668 ( n1772 , n13723 );
    not g11669 ( n510 , n11714 );
    and g11670 ( n2278 , n4690 , n9954 );
    or g11671 ( n10491 , n9490 , n3708 );
    nor g11672 ( n6189 , n12112 , n12626 );
    or g11673 ( n8858 , n769 , n1024 );
    and g11674 ( n14084 , n12038 , n11841 );
    and g11675 ( n8972 , n1729 , n2938 );
    not g11676 ( n1860 , n1936 );
    not g11677 ( n13096 , n6787 );
    and g11678 ( n2243 , n6135 , n1358 );
    and g11679 ( n9312 , n12592 , n13175 );
    not g11680 ( n2445 , n5606 );
    and g11681 ( n14114 , n11607 , n11774 );
    nor g11682 ( n13214 , n4928 , n6914 );
    and g11683 ( n1984 , n4484 , n6116 );
    and g11684 ( n13684 , n103 , n11454 );
    or g11685 ( n11424 , n11183 , n5186 );
    not g11686 ( n11231 , n10069 );
    and g11687 ( n3947 , n7187 , n12590 );
    not g11688 ( n7530 , n2130 );
    and g11689 ( n9959 , n11792 , n8115 );
    not g11690 ( n8631 , n5435 );
    nor g11691 ( n13657 , n900 , n1818 );
    nor g11692 ( n5181 , n10803 , n5069 );
    or g11693 ( n9325 , n976 , n11390 );
    not g11694 ( n1602 , n6357 );
    not g11695 ( n12888 , n4715 );
    nor g11696 ( n6448 , n3182 , n5293 );
    nor g11697 ( n6124 , n3290 , n828 );
    or g11698 ( n12284 , n6706 , n3737 );
    and g11699 ( n5126 , n8965 , n10205 );
    or g11700 ( n12849 , n13118 , n11194 );
    or g11701 ( n9962 , n1834 , n13820 );
    and g11702 ( n6073 , n1481 , n14241 );
    or g11703 ( n11075 , n10624 , n3939 );
    not g11704 ( n13080 , n4325 );
    nor g11705 ( n5299 , n8877 , n6501 );
    or g11706 ( n3119 , n3011 , n7686 );
    nor g11707 ( n13644 , n8378 , n803 );
    or g11708 ( n3259 , n9490 , n12296 );
    or g11709 ( n6524 , n12870 , n9157 );
    or g11710 ( n2869 , n10936 , n10932 );
    or g11711 ( n4990 , n12324 , n8917 );
    and g11712 ( n565 , n12949 , n10239 );
    or g11713 ( n7310 , n6595 , n12650 );
    or g11714 ( n3938 , n8825 , n3889 );
    or g11715 ( n11238 , n1838 , n14000 );
    or g11716 ( n12862 , n5236 , n472 );
    or g11717 ( n12850 , n10646 , n4282 );
    and g11718 ( n2854 , n5634 , n13791 );
    and g11719 ( n5004 , n13240 , n4371 );
    and g11720 ( n14489 , n13484 , n11936 );
    not g11721 ( n7041 , n12012 );
    not g11722 ( n9490 , n5974 );
    or g11723 ( n10126 , n1582 , n13946 );
    or g11724 ( n147 , n11405 , n8447 );
    not g11725 ( n4255 , n7086 );
    or g11726 ( n8335 , n4162 , n7302 );
    or g11727 ( n12831 , n11935 , n1405 );
    and g11728 ( n10097 , n10516 , n11462 );
    or g11729 ( n12618 , n2229 , n8640 );
    and g11730 ( n6541 , n6128 , n4819 );
    not g11731 ( n13626 , n4490 );
    nor g11732 ( n343 , n13722 , n2610 );
    or g11733 ( n11004 , n4967 , n8290 );
    or g11734 ( n3287 , n3506 , n6703 );
    and g11735 ( n7989 , n5335 , n1200 );
    and g11736 ( n13151 , n2064 , n9497 );
    or g11737 ( n1177 , n77 , n14001 );
    or g11738 ( n2478 , n930 , n2437 );
    or g11739 ( n8687 , n4468 , n5946 );
    and g11740 ( n3916 , n9509 , n8571 );
    or g11741 ( n1313 , n12622 , n6063 );
    not g11742 ( n9994 , n1544 );
    not g11743 ( n6263 , n9686 );
    or g11744 ( n3604 , n2784 , n6320 );
    nor g11745 ( n4438 , n6672 , n12643 );
    and g11746 ( n12687 , n6965 , n359 );
    and g11747 ( n9079 , n5229 , n9287 );
    or g11748 ( n1598 , n11580 , n13373 );
    or g11749 ( n11611 , n1362 , n13793 );
    and g11750 ( n10695 , n10247 , n7084 );
    and g11751 ( n9223 , n13297 , n6249 );
    nor g11752 ( n1616 , n12866 , n842 );
    or g11753 ( n1153 , n13005 , n6763 );
    and g11754 ( n6539 , n6744 , n1926 );
    and g11755 ( n11221 , n10399 , n11718 );
    or g11756 ( n9734 , n10191 , n14417 );
    or g11757 ( n9187 , n11722 , n13601 );
    or g11758 ( n176 , n5491 , n5224 );
    or g11759 ( n3371 , n5315 , n894 );
    and g11760 ( n10005 , n10820 , n11780 );
    and g11761 ( n10478 , n10166 , n4686 );
    or g11762 ( n14266 , n2750 , n3969 );
    and g11763 ( n5842 , n5940 , n6904 );
    or g11764 ( n745 , n3777 , n4197 );
    or g11765 ( n1870 , n11036 , n3075 );
    and g11766 ( n106 , n687 , n11355 );
    and g11767 ( n3996 , n12636 , n5059 );
    and g11768 ( n6027 , n9190 , n8323 );
    and g11769 ( n4699 , n9726 , n11731 );
    and g11770 ( n2873 , n12202 , n8558 );
    and g11771 ( n3957 , n13421 , n7343 );
    and g11772 ( n5534 , n1047 , n8793 );
    or g11773 ( n12744 , n8714 , n1407 );
    and g11774 ( n3052 , n2682 , n10789 );
    not g11775 ( n4102 , n9388 );
    or g11776 ( n9831 , n2181 , n6545 );
    not g11777 ( n1801 , n11776 );
    or g11778 ( n5528 , n523 , n13347 );
    nor g11779 ( n14500 , n14367 , n14341 );
    or g11780 ( n8904 , n10834 , n7675 );
    and g11781 ( n12349 , n8630 , n10537 );
    and g11782 ( n5257 , n13720 , n13999 );
    not g11783 ( n7436 , n6357 );
    and g11784 ( n7881 , n9564 , n12402 );
    and g11785 ( n351 , n10332 , n160 );
    nor g11786 ( n10481 , n2644 , n9390 );
    and g11787 ( n10259 , n8247 , n3995 );
    not g11788 ( n3944 , n6874 );
    not g11789 ( n6891 , n4325 );
    or g11790 ( n7022 , n8701 , n9302 );
    and g11791 ( n4852 , n7745 , n1302 );
    and g11792 ( n713 , n4300 , n9981 );
    and g11793 ( n2907 , n12105 , n12462 );
    nor g11794 ( n8818 , n5132 , n6944 );
    not g11795 ( n82 , n6055 );
    and g11796 ( n13500 , n12226 , n4245 );
    and g11797 ( n5964 , n6354 , n11828 );
    or g11798 ( n12339 , n4205 , n4353 );
    or g11799 ( n11301 , n4128 , n8468 );
    not g11800 ( n14286 , n11269 );
    or g11801 ( n12468 , n6857 , n7942 );
    not g11802 ( n12403 , n2011 );
    and g11803 ( n3795 , n4347 , n1441 );
    or g11804 ( n10090 , n11804 , n12076 );
    or g11805 ( n12158 , n1172 , n2136 );
    and g11806 ( n1721 , n13240 , n11810 );
    or g11807 ( n7572 , n14188 , n12801 );
    not g11808 ( n9238 , n1955 );
    and g11809 ( n10754 , n12990 , n2289 );
    and g11810 ( n8085 , n8800 , n57 );
    not g11811 ( n799 , n7871 );
    not g11812 ( n13132 , n2334 );
    or g11813 ( n5976 , n6690 , n8689 );
    and g11814 ( n12648 , n3932 , n3770 );
    or g11815 ( n6497 , n11551 , n13527 );
    and g11816 ( n1238 , n4880 , n975 );
    or g11817 ( n8815 , n1202 , n514 );
    nor g11818 ( n10122 , n300 , n6277 );
    not g11819 ( n10883 , n4744 );
    or g11820 ( n3751 , n1391 , n5341 );
    nor g11821 ( n14044 , n8856 , n32 );
    or g11822 ( n9892 , n769 , n5964 );
    nor g11823 ( n7209 , n10936 , n13266 );
    nor g11824 ( n12956 , n7971 , n1382 );
    and g11825 ( n5210 , n12935 , n2838 );
    not g11826 ( n4739 , n4939 );
    nor g11827 ( n1703 , n11017 , n10934 );
    or g11828 ( n8806 , n10294 , n1374 );
    and g11829 ( n9376 , n13147 , n9674 );
    or g11830 ( n9483 , n4092 , n1434 );
    or g11831 ( n620 , n4340 , n11258 );
    nor g11832 ( n699 , n13811 , n2928 );
    and g11833 ( n7855 , n11163 , n8196 );
    nor g11834 ( n11482 , n2566 , n6070 );
    or g11835 ( n2787 , n11036 , n8091 );
    or g11836 ( n5557 , n974 , n321 );
    or g11837 ( n14224 , n5641 , n12564 );
    not g11838 ( n11975 , n179 );
    not g11839 ( n5236 , n8695 );
    or g11840 ( n6341 , n10731 , n7908 );
    and g11841 ( n13339 , n8047 , n104 );
    or g11842 ( n13645 , n8476 , n4678 );
    not g11843 ( n14367 , n10219 );
    and g11844 ( n5301 , n501 , n13258 );
    nor g11845 ( n3789 , n8378 , n8670 );
    not g11846 ( n8025 , n9456 );
    and g11847 ( n9666 , n3923 , n8495 );
    and g11848 ( n10397 , n9191 , n14364 );
    or g11849 ( n362 , n8015 , n483 );
    or g11850 ( n7218 , n14029 , n12641 );
    and g11851 ( n11485 , n13507 , n8657 );
    and g11852 ( n7186 , n7970 , n13954 );
    not g11853 ( n5434 , n1724 );
    nor g11854 ( n9779 , n1697 , n1111 );
    and g11855 ( n431 , n13227 , n9217 );
    and g11856 ( n10239 , n2505 , n14252 );
    or g11857 ( n3825 , n13847 , n8271 );
    or g11858 ( n5931 , n13537 , n3374 );
    or g11859 ( n67 , n14110 , n8161 );
    or g11860 ( n4823 , n2694 , n7539 );
    and g11861 ( n13086 , n5434 , n1849 );
    or g11862 ( n7099 , n1189 , n3267 );
    and g11863 ( n4451 , n446 , n9339 );
    or g11864 ( n7778 , n317 , n3535 );
    and g11865 ( n5441 , n7015 , n763 );
    and g11866 ( n11847 , n203 , n1065 );
    and g11867 ( n9288 , n10562 , n645 );
    or g11868 ( n5868 , n13485 , n6232 );
    or g11869 ( n1599 , n5180 , n11212 );
    or g11870 ( n13111 , n1137 , n4951 );
    not g11871 ( n1780 , n13365 );
    or g11872 ( n4635 , n2179 , n6499 );
    and g11873 ( n773 , n9953 , n4290 );
    or g11874 ( n9235 , n13518 , n3931 );
    and g11875 ( n9699 , n2904 , n3794 );
    or g11876 ( n5072 , n7219 , n5561 );
    and g11877 ( n12817 , n6625 , n12284 );
    and g11878 ( n2275 , n9944 , n2331 );
    and g11879 ( n11167 , n4627 , n4217 );
    or g11880 ( n8175 , n6654 , n6601 );
    nor g11881 ( n12010 , n1742 , n2420 );
    and g11882 ( n12776 , n1377 , n9406 );
    and g11883 ( n10948 , n9015 , n5086 );
    not g11884 ( n4095 , n13038 );
    or g11885 ( n10940 , n11420 , n4970 );
    and g11886 ( n10904 , n10855 , n4444 );
    and g11887 ( n2830 , n14091 , n3208 );
    or g11888 ( n8878 , n3914 , n2129 );
    or g11889 ( n11955 , n14400 , n2523 );
    nor g11890 ( n6966 , n8015 , n8784 );
    nor g11891 ( n8885 , n12569 , n9378 );
    not g11892 ( n7352 , n5354 );
    not g11893 ( n946 , n1506 );
    and g11894 ( n710 , n7596 , n6994 );
    and g11895 ( n14522 , n3861 , n10420 );
    not g11896 ( n14327 , n7507 );
    or g11897 ( n6218 , n10534 , n4985 );
    and g11898 ( n4188 , n2846 , n3382 );
    and g11899 ( n12864 , n5999 , n8475 );
    or g11900 ( n10220 , n7122 , n84 );
    and g11901 ( n12905 , n2961 , n14221 );
    and g11902 ( n9951 , n6167 , n3269 );
    or g11903 ( n2599 , n1685 , n4809 );
    and g11904 ( n13183 , n446 , n11656 );
    or g11905 ( n4969 , n747 , n3190 );
    and g11906 ( n5474 , n13404 , n1853 );
    or g11907 ( n1891 , n4065 , n13559 );
    not g11908 ( n2318 , n1267 );
    not g11909 ( n8462 , n11188 );
    or g11910 ( n11573 , n11048 , n14411 );
    not g11911 ( n7358 , n7600 );
    not g11912 ( n304 , n2040 );
    and g11913 ( n962 , n3766 , n12647 );
    and g11914 ( n5646 , n6343 , n9671 );
    and g11915 ( n5811 , n14327 , n12436 );
    and g11916 ( n1036 , n13342 , n6852 );
    and g11917 ( n11577 , n7063 , n7859 );
    or g11918 ( n171 , n11572 , n486 );
    and g11919 ( n2603 , n5489 , n7874 );
    and g11920 ( n8156 , n3766 , n61 );
    not g11921 ( n11765 , n407 );
    and g11922 ( n11092 , n687 , n12339 );
    and g11923 ( n4761 , n13362 , n1554 );
    not g11924 ( n8907 , n1265 );
    not g11925 ( n11455 , n11743 );
    or g11926 ( n8354 , n1821 , n4890 );
    not g11927 ( n10247 , n11969 );
    or g11928 ( n5156 , n13413 , n2604 );
    and g11929 ( n2776 , n5137 , n12051 );
    and g11930 ( n4567 , n10705 , n9983 );
    not g11931 ( n3094 , n14332 );
    not g11932 ( n11816 , n920 );
    and g11933 ( n12574 , n4614 , n11002 );
    not g11934 ( n11542 , n4609 );
    nor g11935 ( n424 , n12191 , n2540 );
    nor g11936 ( n5573 , n12888 , n8751 );
    and g11937 ( n14149 , n13252 , n2678 );
    and g11938 ( n2388 , n13147 , n4010 );
    or g11939 ( n905 , n3527 , n9024 );
    or g11940 ( n10688 , n4154 , n3506 );
    or g11941 ( n13461 , n6205 , n11377 );
    and g11942 ( n12871 , n10072 , n855 );
    and g11943 ( n3336 , n7068 , n11107 );
    and g11944 ( n6103 , n12521 , n7570 );
    or g11945 ( n1786 , n4508 , n2291 );
    and g11946 ( n2167 , n7810 , n8712 );
    and g11947 ( n524 , n8066 , n12692 );
    and g11948 ( n1894 , n2226 , n10395 );
    or g11949 ( n722 , n14449 , n9527 );
    and g11950 ( n2463 , n11484 , n4356 );
    or g11951 ( n10003 , n9541 , n4442 );
    and g11952 ( n7705 , n428 , n13737 );
    or g11953 ( n11151 , n4895 , n8780 );
    nor g11954 ( n2434 , n5468 , n4133 );
    or g11955 ( n893 , n7912 , n8754 );
    not g11956 ( n11148 , n11809 );
    not g11957 ( n11870 , n10172 );
    not g11958 ( n8983 , n2545 );
    and g11959 ( n3141 , n10166 , n14350 );
    nor g11960 ( n13097 , n6044 , n11291 );
    not g11961 ( n4205 , n6978 );
    or g11962 ( n7240 , n1660 , n12236 );
    nor g11963 ( n1767 , n12075 , n14310 );
    or g11964 ( n10381 , n85 , n429 );
    nor g11965 ( n11041 , n7223 , n8286 );
    or g11966 ( n9336 , n7736 , n12036 );
    not g11967 ( n12185 , n11715 );
    or g11968 ( n778 , n13310 , n11500 );
    or g11969 ( n9821 , n13875 , n11109 );
    and g11970 ( n6148 , n10822 , n7367 );
    and g11971 ( n11947 , n7187 , n11359 );
    nor g11972 ( n7432 , n7011 , n11000 );
    or g11973 ( n13623 , n4821 , n12408 );
    or g11974 ( n7325 , n4255 , n12438 );
    or g11975 ( n1883 , n14188 , n5338 );
    or g11976 ( n6463 , n7219 , n2873 );
    not g11977 ( n4657 , n10469 );
    not g11978 ( n8704 , n9546 );
    and g11979 ( n7917 , n11803 , n1422 );
    not g11980 ( n3204 , n5429 );
    not g11981 ( n12425 , n9456 );
    or g11982 ( n6710 , n817 , n5045 );
    or g11983 ( n1188 , n3093 , n3433 );
    or g11984 ( n6616 , n8726 , n10633 );
    and g11985 ( n10749 , n2064 , n14492 );
    and g11986 ( n1867 , n11814 , n13368 );
    and g11987 ( n12282 , n541 , n2161 );
    or g11988 ( n9940 , n7551 , n10682 );
    and g11989 ( n1094 , n6555 , n3296 );
    not g11990 ( n13252 , n10469 );
    and g11991 ( n460 , n8569 , n10590 );
    not g11992 ( n4365 , n10112 );
    or g11993 ( n9538 , n8816 , n6295 );
    and g11994 ( n11015 , n6318 , n3595 );
    or g11995 ( n6675 , n4908 , n4976 );
    or g11996 ( n4648 , n12019 , n224 );
    or g11997 ( n8712 , n12568 , n5687 );
    and g11998 ( n11648 , n10302 , n11104 );
    not g11999 ( n5852 , n11441 );
    and g12000 ( n12943 , n8025 , n3657 );
    or g12001 ( n10240 , n5548 , n8910 );
    or g12002 ( n10579 , n6711 , n8660 );
    nor g12003 ( n12283 , n5132 , n1703 );
    nor g12004 ( n13313 , n6971 , n8154 );
    and g12005 ( n4315 , n8849 , n8149 );
    or g12006 ( n233 , n1685 , n1587 );
    not g12007 ( n10396 , n9306 );
    or g12008 ( n9825 , n14166 , n5799 );
    and g12009 ( n7598 , n501 , n7845 );
    and g12010 ( n10020 , n2473 , n10662 );
    or g12011 ( n13970 , n4484 , n8746 );
    and g12012 ( n4193 , n3932 , n7406 );
    not g12013 ( n9618 , n14433 );
    or g12014 ( n806 , n478 , n8668 );
    and g12015 ( n12946 , n8702 , n1205 );
    not g12016 ( n10539 , n4847 );
    or g12017 ( n11683 , n1613 , n6741 );
    or g12018 ( n11478 , n14430 , n1740 );
    and g12019 ( n5746 , n6128 , n358 );
    or g12020 ( n208 , n2025 , n6083 );
    or g12021 ( n7885 , n14110 , n10243 );
    not g12022 ( n10357 , n9613 );
    not g12023 ( n827 , n4711 );
    or g12024 ( n7247 , n9742 , n6186 );
    or g12025 ( n14158 , n1805 , n5608 );
    not g12026 ( n2908 , n2383 );
    and g12027 ( n5593 , n11737 , n4264 );
    not g12028 ( n13201 , n11606 );
    not g12029 ( n5024 , n13012 );
    nor g12030 ( n7804 , n3873 , n3789 );
    or g12031 ( n1635 , n14401 , n7295 );
    not g12032 ( n9291 , n749 );
    or g12033 ( n5079 , n12023 , n14036 );
    and g12034 ( n12446 , n4929 , n5955 );
    and g12035 ( n854 , n5857 , n37 );
    and g12036 ( n13953 , n11158 , n3177 );
    or g12037 ( n8571 , n5491 , n11859 );
    not g12038 ( n10229 , n10975 );
    or g12039 ( n7366 , n4739 , n12089 );
    and g12040 ( n10819 , n1662 , n9361 );
    or g12041 ( n9234 , n10449 , n2596 );
    and g12042 ( n6763 , n98 , n11483 );
    or g12043 ( n8996 , n5472 , n9076 );
    or g12044 ( n456 , n1059 , n5033 );
    not g12045 ( n14139 , n9516 );
    and g12046 ( n7456 , n12015 , n3965 );
    or g12047 ( n13202 , n4199 , n9063 );
    and g12048 ( n13615 , n5582 , n6977 );
    or g12049 ( n6473 , n1805 , n6661 );
    or g12050 ( n3674 , n5064 , n12161 );
    nor g12051 ( n13148 , n13941 , n13997 );
    not g12052 ( n12935 , n11474 );
    or g12053 ( n2567 , n5807 , n5844 );
    and g12054 ( n11978 , n9564 , n5976 );
    or g12055 ( n2306 , n6695 , n868 );
    not g12056 ( n14282 , n10108 );
    or g12057 ( n6803 , n8581 , n11363 );
    not g12058 ( n13501 , n7819 );
    nor g12059 ( n6277 , n573 , n3951 );
    and g12060 ( n4528 , n7745 , n13370 );
    or g12061 ( n14492 , n5587 , n13105 );
    or g12062 ( n6716 , n9490 , n9542 );
    not g12063 ( n4535 , n10423 );
    or g12064 ( n4494 , n4468 , n9504 );
    or g12065 ( n8653 , n2272 , n9955 );
    and g12066 ( n3792 , n4347 , n14205 );
    or g12067 ( n9430 , n7862 , n6532 );
    not g12068 ( n10953 , n1222 );
    not g12069 ( n12644 , n4341 );
    and g12070 ( n5550 , n5046 , n1616 );
    not g12071 ( n8151 , n2383 );
    or g12072 ( n11672 , n10089 , n11367 );
    or g12073 ( n2552 , n974 , n2413 );
    or g12074 ( n12235 , n5180 , n2258 );
    not g12075 ( n10322 , n6516 );
    and g12076 ( n4847 , n11966 , n5839 );
    or g12077 ( n14277 , n5315 , n3373 );
    and g12078 ( n11436 , n12615 , n5470 );
    or g12079 ( n5233 , n2747 , n8108 );
    and g12080 ( n11264 , n1409 , n12103 );
    not g12081 ( n8697 , n9583 );
    and g12082 ( n11788 , n2029 , n7842 );
    or g12083 ( n10296 , n5936 , n14055 );
    not g12084 ( n6085 , n10069 );
    and g12085 ( n13174 , n4354 , n1379 );
    and g12086 ( n12333 , n6744 , n6442 );
    and g12087 ( n3181 , n3526 , n9556 );
    and g12088 ( n205 , n10556 , n2638 );
    not g12089 ( n12768 , n656 );
    nor g12090 ( n11073 , n5762 , n330 );
    or g12091 ( n7270 , n14401 , n7257 );
    not g12092 ( n14200 , n2061 );
    or g12093 ( n13873 , n5732 , n6467 );
    not g12094 ( n4266 , n11426 );
    or g12095 ( n3778 , n13518 , n10153 );
    not g12096 ( n13107 , n1571 );
    or g12097 ( n11086 , n13356 , n8647 );
    and g12098 ( n1221 , n2783 , n7558 );
    nor g12099 ( n4524 , n6971 , n7921 );
    and g12100 ( n9783 , n12265 , n6438 );
    or g12101 ( n694 , n1875 , n7907 );
    nor g12102 ( n1304 , n10730 , n13910 );
    and g12103 ( n5125 , n13407 , n2847 );
    and g12104 ( n6585 , n13338 , n7497 );
    or g12105 ( n2737 , n9229 , n9502 );
    not g12106 ( n10309 , n4203 );
    not g12107 ( n1937 , n9456 );
    nor g12108 ( n2398 , n7905 , n5703 );
    and g12109 ( n14279 , n13433 , n6490 );
    nor g12110 ( n101 , n10571 , n9513 );
    and g12111 ( n14374 , n2422 , n9585 );
    and g12112 ( n2296 , n3952 , n9268 );
    or g12113 ( n13349 , n1362 , n11886 );
    or g12114 ( n7198 , n5362 , n1514 );
    and g12115 ( n7850 , n7957 , n13621 );
    and g12116 ( n8890 , n3485 , n14068 );
    and g12117 ( n11190 , n11362 , n4894 );
    or g12118 ( n5887 , n4195 , n908 );
    or g12119 ( n295 , n13675 , n1655 );
    or g12120 ( n4342 , n13814 , n4022 );
    or g12121 ( n2187 , n7584 , n3248 );
    and g12122 ( n10744 , n11679 , n14220 );
    or g12123 ( n8032 , n12351 , n13304 );
    not g12124 ( n4163 , n1760 );
    and g12125 ( n3386 , n10166 , n13450 );
    or g12126 ( n4644 , n1172 , n8440 );
    nor g12127 ( n5810 , n9035 , n3139 );
    not g12128 ( n406 , n82 );
    and g12129 ( n10564 , n4156 , n6827 );
    or g12130 ( n4314 , n6471 , n7117 );
    nor g12131 ( n10353 , n194 , n14362 );
    or g12132 ( n5777 , n7888 , n11342 );
    not g12133 ( n5899 , n871 );
    or g12134 ( n10320 , n2878 , n395 );
    or g12135 ( n3114 , n13885 , n7762 );
    or g12136 ( n8295 , n2510 , n7992 );
    nor g12137 ( n11112 , n7905 , n10907 );
    and g12138 ( n1886 , n1904 , n5482 );
    not g12139 ( n4925 , n6804 );
    or g12140 ( n13932 , n976 , n9982 );
    and g12141 ( n3732 , n3755 , n2514 );
    and g12142 ( n6969 , n8512 , n6616 );
    and g12143 ( n9696 , n2367 , n7333 );
    not g12144 ( n8963 , n1861 );
    not g12145 ( n7476 , n13882 );
    not g12146 ( n5782 , n8419 );
    or g12147 ( n14095 , n12500 , n7159 );
    or g12148 ( n5751 , n8581 , n2438 );
    not g12149 ( n3427 , n9640 );
    or g12150 ( n9677 , n12167 , n2699 );
    or g12151 ( n2902 , n7011 , n5447 );
    and g12152 ( n10628 , n4581 , n11272 );
    not g12153 ( n2848 , n6422 );
    nor g12154 ( n2183 , n3234 , n5755 );
    nor g12155 ( n5912 , n1178 , n3359 );
    or g12156 ( n10092 , n4877 , n12177 );
    nor g12157 ( n3685 , n6020 , n13528 );
    or g12158 ( n11807 , n10713 , n4136 );
    not g12159 ( n3762 , n2895 );
    or g12160 ( n7485 , n6090 , n1269 );
    or g12161 ( n2965 , n6471 , n990 );
    and g12162 ( n4758 , n13489 , n8710 );
    and g12163 ( n5411 , n6724 , n8843 );
    or g12164 ( n13197 , n9269 , n12041 );
    not g12165 ( n2985 , n442 );
    and g12166 ( n9070 , n5348 , n487 );
    not g12167 ( n10351 , n1267 );
    nor g12168 ( n6132 , n5480 , n8628 );
    or g12169 ( n6766 , n4923 , n5276 );
    nor g12170 ( n5957 , n3290 , n9668 );
    not g12171 ( n89 , n9306 );
    or g12172 ( n7264 , n7116 , n3203 );
    or g12173 ( n3653 , n2229 , n2550 );
    or g12174 ( n6821 , n4562 , n1002 );
    not g12175 ( n9865 , n8565 );
    or g12176 ( n8140 , n5315 , n10392 );
    not g12177 ( n4354 , n4618 );
    or g12178 ( n7108 , n8748 , n7729 );
    or g12179 ( n4689 , n2111 , n7088 );
    or g12180 ( n1073 , n14006 , n4785 );
    and g12181 ( n14410 , n4163 , n5113 );
    and g12182 ( n1370 , n4244 , n7883 );
    and g12183 ( n2267 , n2783 , n6694 );
    and g12184 ( n3908 , n7596 , n12251 );
    and g12185 ( n9904 , n12038 , n4485 );
    or g12186 ( n8636 , n13310 , n10528 );
    and g12187 ( n2303 , n13107 , n12470 );
    and g12188 ( n2670 , n11033 , n5296 );
    not g12189 ( n333 , n7681 );
    or g12190 ( n134 , n5409 , n9760 );
    nor g12191 ( n7512 , n13937 , n14028 );
    or g12192 ( n11248 , n1602 , n9749 );
    or g12193 ( n1884 , n1258 , n11795 );
    and g12194 ( n3598 , n5489 , n9610 );
    and g12195 ( n682 , n5033 , n101 );
    and g12196 ( n4361 , n14063 , n13268 );
    and g12197 ( n13624 , n2322 , n6756 );
    and g12198 ( n8028 , n4757 , n7453 );
    and g12199 ( n4660 , n9102 , n7247 );
    and g12200 ( n5136 , n13755 , n5444 );
    or g12201 ( n863 , n12130 , n9410 );
    not g12202 ( n6313 , n496 );
    not g12203 ( n7700 , n3681 );
    and g12204 ( n12224 , n4973 , n2655 );
    nor g12205 ( n14310 , n7200 , n4759 );
    or g12206 ( n2614 , n172 , n2261 );
    not g12207 ( n10871 , n3357 );
    and g12208 ( n14339 , n6649 , n6253 );
    and g12209 ( n1987 , n12449 , n10659 );
    not g12210 ( n7426 , n7404 );
    and g12211 ( n6231 , n13575 , n10499 );
    and g12212 ( n2321 , n8025 , n9082 );
    not g12213 ( n5065 , n9863 );
    not g12214 ( n7997 , n9893 );
    or g12215 ( n5285 , n3512 , n7175 );
    and g12216 ( n2222 , n7419 , n8141 );
    or g12217 ( n12873 , n13501 , n4553 );
    or g12218 ( n6360 , n7249 , n7383 );
    or g12219 ( n368 , n14337 , n2668 );
    and g12220 ( n8078 , n3276 , n3661 );
    and g12221 ( n7506 , n4289 , n9025 );
    and g12222 ( n14343 , n11153 , n8600 );
    nor g12223 ( n6551 , n4296 , n6365 );
    or g12224 ( n7564 , n11581 , n2776 );
    nor g12225 ( n8104 , n11151 , n6408 );
    and g12226 ( n3737 , n501 , n6561 );
    and g12227 ( n13529 , n2486 , n11944 );
    or g12228 ( n10837 , n5184 , n8635 );
    not g12229 ( n12802 , n7278 );
    or g12230 ( n5070 , n5562 , n8566 );
    not g12231 ( n10668 , n11305 );
    or g12232 ( n12884 , n89 , n13333 );
    not g12233 ( n7200 , n6305 );
    not g12234 ( n11453 , n1342 );
    or g12235 ( n14317 , n12169 , n13345 );
    not g12236 ( n555 , n409 );
    not g12237 ( n6606 , n10303 );
    or g12238 ( n10735 , n480 , n1872 );
    and g12239 ( n11798 , n1610 , n13321 );
    not g12240 ( n9601 , n11574 );
    not g12241 ( n11093 , n6975 );
    and g12242 ( n11723 , n11816 , n11965 );
    and g12243 ( n8602 , n7421 , n1594 );
    and g12244 ( n6153 , n9953 , n5044 );
    or g12245 ( n2114 , n8714 , n1398 );
    or g12246 ( n10580 , n1728 , n4391 );
    not g12247 ( n10660 , n14483 );
    and g12248 ( n14359 , n4790 , n2680 );
    and g12249 ( n495 , n8358 , n4061 );
    or g12250 ( n13965 , n6039 , n4121 );
    nor g12251 ( n10565 , n2355 , n13116 );
    or g12252 ( n7477 , n7250 , n5140 );
    or g12253 ( n2967 , n8975 , n10945 );
    not g12254 ( n7091 , n11001 );
    or g12255 ( n9304 , n10019 , n10606 );
    not g12256 ( n2804 , n8780 );
    nor g12257 ( n8443 , n12292 , n11078 );
    not g12258 ( n6426 , n9757 );
    and g12259 ( n2935 , n2983 , n7778 );
    or g12260 ( n7121 , n13226 , n3787 );
    not g12261 ( n1522 , n4415 );
    not g12262 ( n11362 , n14163 );
    nor g12263 ( n10082 , n8543 , n2431 );
    nor g12264 ( n9637 , n3445 , n10447 );
    or g12265 ( n3018 , n3161 , n5110 );
    and g12266 ( n4127 , n8393 , n8921 );
    nor g12267 ( n7066 , n5132 , n247 );
    and g12268 ( n7561 , n12620 , n3460 );
    not g12269 ( n14449 , n4203 );
    and g12270 ( n1434 , n12832 , n10634 );
    and g12271 ( n6240 , n8569 , n979 );
    not g12272 ( n11420 , n10629 );
    and g12273 ( n13712 , n706 , n13831 );
    and g12274 ( n1502 , n8950 , n9937 );
    and g12275 ( n2500 , n7015 , n433 );
    nor g12276 ( n8857 , n9818 , n2317 );
    not g12277 ( n12472 , n8223 );
    and g12278 ( n9531 , n8950 , n3038 );
    or g12279 ( n12173 , n11804 , n5428 );
    and g12280 ( n2121 , n2281 , n1346 );
    or g12281 ( n968 , n6857 , n12551 );
    and g12282 ( n12007 , n12986 , n3781 );
    not g12283 ( n5053 , n9865 );
    and g12284 ( n5822 , n2180 , n11516 );
    not g12285 ( n8512 , n5504 );
    or g12286 ( n4855 , n10396 , n935 );
    and g12287 ( n12901 , n3097 , n10903 );
    or g12288 ( n5878 , n10300 , n5705 );
    not g12289 ( n13718 , n1833 );
    or g12290 ( n4395 , n4631 , n5739 );
    nor g12291 ( n5192 , n329 , n4309 );
    and g12292 ( n2116 , n10457 , n3463 );
    nor g12293 ( n1393 , n5621 , n11681 );
    not g12294 ( n1678 , n13908 );
    and g12295 ( n4470 , n3904 , n7095 );
    and g12296 ( n13502 , n4690 , n10816 );
    not g12297 ( n11706 , n9406 );
    and g12298 ( n14480 , n7421 , n2558 );
    or g12299 ( n217 , n317 , n6683 );
    or g12300 ( n8740 , n12994 , n7002 );
    or g12301 ( n9522 , n7245 , n4243 );
    not g12302 ( n13627 , n14134 );
    not g12303 ( n9650 , n2906 );
    or g12304 ( n675 , n974 , n836 );
    or g12305 ( n5329 , n10062 , n12258 );
    or g12306 ( n5979 , n12576 , n11169 );
    or g12307 ( n3495 , n8816 , n9572 );
    not g12308 ( n12543 , n6123 );
    not g12309 ( n7527 , n3357 );
    not g12310 ( n4433 , n1027 );
    or g12311 ( n13071 , n4481 , n5050 );
    or g12312 ( n12560 , n4435 , n10967 );
    not g12313 ( n2729 , n12168 );
    and g12314 ( n626 , n6531 , n3389 );
    and g12315 ( n9445 , n3435 , n13588 );
    and g12316 ( n5609 , n1254 , n11150 );
    and g12317 ( n1877 , n9323 , n6312 );
    and g12318 ( n4837 , n1339 , n12468 );
    and g12319 ( n13548 , n406 , n6623 );
    and g12320 ( n14369 , n5628 , n3056 );
    not g12321 ( n4573 , n11756 );
    and g12322 ( n13098 , n13850 , n1099 );
    and g12323 ( n9693 , n2445 , n11437 );
    not g12324 ( n4046 , n10917 );
    nor g12325 ( n13060 , n3445 , n11543 );
    and g12326 ( n11212 , n4098 , n11835 );
    and g12327 ( n1259 , n10399 , n9027 );
    or g12328 ( n4723 , n2949 , n13613 );
    or g12329 ( n3229 , n6085 , n10949 );
    not g12330 ( n14107 , n2545 );
    or g12331 ( n4744 , n14360 , n8598 );
    or g12332 ( n10831 , n10626 , n3159 );
    or g12333 ( n9711 , n5647 , n8755 );
    not g12334 ( n6256 , n7282 );
    or g12335 ( n6844 , n14245 , n4292 );
    and g12336 ( n10570 , n1539 , n14413 );
    or g12337 ( n5900 , n1582 , n4772 );
    not g12338 ( n8877 , n3681 );
    and g12339 ( n2586 , n10399 , n5138 );
    nor g12340 ( n6315 , n14075 , n3462 );
    or g12341 ( n5671 , n11542 , n9933 );
    not g12342 ( n2212 , n11453 );
    and g12343 ( n1807 , n9188 , n5858 );
    and g12344 ( n6346 , n1854 , n2532 );
    or g12345 ( n10706 , n11360 , n8890 );
    and g12346 ( n7073 , n5023 , n6210 );
    or g12347 ( n4926 , n10560 , n5571 );
    or g12348 ( n2678 , n3546 , n287 );
    or g12349 ( n13355 , n2897 , n1370 );
    not g12350 ( n11715 , n5117 );
    and g12351 ( n7314 , n7079 , n144 );
    not g12352 ( n13467 , n3976 );
    and g12353 ( n5761 , n4527 , n13434 );
    and g12354 ( n13717 , n12858 , n12063 );
    or g12355 ( n6328 , n5139 , n12828 );
    nor g12356 ( n665 , n2462 , n8868 );
    nor g12357 ( n6918 , n14011 , n7069 );
    or g12358 ( n7353 , n4741 , n11844 );
    and g12359 ( n7331 , n7211 , n11651 );
    and g12360 ( n14099 , n4525 , n11831 );
    or g12361 ( n3620 , n3877 , n1331 );
    not g12362 ( n13158 , n10973 );
    or g12363 ( n9928 , n1031 , n12026 );
    and g12364 ( n11686 , n9898 , n4583 );
    or g12365 ( n13631 , n4876 , n10902 );
    not g12366 ( n348 , n11854 );
    and g12367 ( n10256 , n10399 , n2696 );
    or g12368 ( n470 , n14419 , n5612 );
    not g12369 ( n8045 , n3046 );
    not g12370 ( n7208 , n3402 );
    or g12371 ( n518 , n11047 , n14199 );
    and g12372 ( n579 , n1255 , n11570 );
    and g12373 ( n2373 , n9323 , n13202 );
    or g12374 ( n11642 , n504 , n12245 );
    nor g12375 ( n4287 , n1771 , n1390 );
    nor g12376 ( n1806 , n4313 , n4654 );
    and g12377 ( n2349 , n3365 , n469 );
    nor g12378 ( n10952 , n1697 , n8730 );
    not g12379 ( n3715 , n3356 );
    and g12380 ( n4597 , n1140 , n11744 );
    or g12381 ( n11298 , n8908 , n12617 );
    or g12382 ( n10618 , n1697 , n7054 );
    or g12383 ( n4559 , n14430 , n10908 );
    and g12384 ( n7566 , n12802 , n890 );
    or g12385 ( n4767 , n9807 , n13481 );
    or g12386 ( n11045 , n10300 , n13987 );
    or g12387 ( n716 , n5815 , n9581 );
    and g12388 ( n5162 , n5948 , n8806 );
    and g12389 ( n14153 , n406 , n10327 );
    and g12390 ( n1764 , n2461 , n12210 );
    and g12391 ( n10119 , n103 , n12962 );
    or g12392 ( n10590 , n504 , n7641 );
    or g12393 ( n1768 , n4045 , n14086 );
    or g12394 ( n6510 , n5180 , n14099 );
    and g12395 ( n2040 , n9819 , n10900 );
    or g12396 ( n5106 , n3099 , n3752 );
    and g12397 ( n13018 , n2669 , n154 );
    and g12398 ( n13121 , n3526 , n8287 );
    and g12399 ( n11443 , n7693 , n6676 );
    and g12400 ( n2299 , n10357 , n8913 );
    not g12401 ( n2750 , n1041 );
    or g12402 ( n9268 , n5480 , n13697 );
    or g12403 ( n5698 , n2401 , n9053 );
    or g12404 ( n13357 , n2562 , n7165 );
    nor g12405 ( n9553 , n1693 , n14130 );
    not g12406 ( n8801 , n12930 );
    not g12407 ( n8393 , n5951 );
    and g12408 ( n13552 , n4486 , n663 );
    nor g12409 ( n5956 , n2727 , n1046 );
    not g12410 ( n13477 , n10985 );
    and g12411 ( n1982 , n2099 , n13920 );
    not g12412 ( n887 , n30 );
    and g12413 ( n2774 , n3370 , n10962 );
    not g12414 ( n5275 , n10376 );
    and g12415 ( n4454 , n4445 , n3133 );
    or g12416 ( n8192 , n13531 , n5455 );
    and g12417 ( n630 , n4036 , n5549 );
    nor g12418 ( n12133 , n4656 , n5398 );
    or g12419 ( n11956 , n782 , n10958 );
    and g12420 ( n1195 , n3365 , n13786 );
    not g12421 ( n2354 , n11765 );
    not g12422 ( n11837 , n8926 );
    nor g12423 ( n10306 , n3944 , n13964 );
    nor g12424 ( n4759 , n11901 , n3879 );
    or g12425 ( n983 , n11090 , n3851 );
    and g12426 ( n6708 , n3401 , n219 );
    and g12427 ( n5765 , n7529 , n10058 );
    and g12428 ( n272 , n12226 , n3112 );
    and g12429 ( n12797 , n4574 , n13436 );
    and g12430 ( n688 , n12990 , n2601 );
    not g12431 ( n4546 , n8048 );
    or g12432 ( n4950 , n5936 , n1879 );
    or g12433 ( n3002 , n6263 , n1941 );
    not g12434 ( n2269 , n2946 );
    not g12435 ( n13016 , n14154 );
    or g12436 ( n8219 , n2089 , n7936 );
    or g12437 ( n13827 , n116 , n7563 );
    or g12438 ( n12984 , n12968 , n8777 );
    or g12439 ( n547 , n6781 , n1482 );
    or g12440 ( n12471 , n3125 , n2463 );
    and g12441 ( n12701 , n11814 , n14263 );
    or g12442 ( n1614 , n6466 , n11633 );
    not g12443 ( n13485 , n11415 );
    nor g12444 ( n14248 , n11232 , n4984 );
    nor g12445 ( n7452 , n3640 , n2150 );
    and g12446 ( n7583 , n7677 , n3375 );
    and g12447 ( n407 , n6849 , n5166 );
    and g12448 ( n10102 , n13745 , n4151 );
    and g12449 ( n13173 , n10710 , n2037 );
    and g12450 ( n8785 , n1481 , n6860 );
    nor g12451 ( n10340 , n12527 , n12700 );
    not g12452 ( n6705 , n6466 );
    and g12453 ( n2295 , n10822 , n7442 );
    not g12454 ( n261 , n4500 );
    or g12455 ( n4071 , n5710 , n8326 );
    and g12456 ( n3362 , n12038 , n4302 );
    not g12457 ( n2330 , n1436 );
    and g12458 ( n4032 , n6753 , n1253 );
    and g12459 ( n11487 , n7060 , n2292 );
    or g12460 ( n218 , n10825 , n1807 );
    and g12461 ( n9463 , n9113 , n4168 );
    and g12462 ( n13487 , n2058 , n11070 );
    and g12463 ( n6264 , n13012 , n8345 );
    or g12464 ( n3085 , n4180 , n6671 );
    or g12465 ( n1379 , n1669 , n4448 );
    and g12466 ( n941 , n4095 , n11430 );
    or g12467 ( n8533 , n1914 , n12052 );
    or g12468 ( n1179 , n12870 , n13969 );
    or g12469 ( n5424 , n4908 , n9257 );
    nor g12470 ( n2663 , n500 , n8573 );
    not g12471 ( n10209 , n9924 );
    or g12472 ( n1470 , n2246 , n2756 );
    or g12473 ( n945 , n8983 , n12899 );
    nor g12474 ( n142 , n9136 , n310 );
    or g12475 ( n9397 , n2387 , n13717 );
    or g12476 ( n11726 , n3628 , n4175 );
    and g12477 ( n1969 , n3755 , n12896 );
    and g12478 ( n843 , n8300 , n7882 );
    not g12479 ( n7421 , n10975 );
    or g12480 ( n5059 , n10660 , n14303 );
    and g12481 ( n8405 , n79 , n8693 );
    not g12482 ( n473 , n13408 );
    and g12483 ( n12059 , n309 , n7619 );
    and g12484 ( n2720 , n8043 , n8724 );
    not g12485 ( n9885 , n11548 );
    or g12486 ( n13068 , n8513 , n1515 );
    and g12487 ( n12937 , n4267 , n8498 );
    not g12488 ( n9340 , n398 );
    and g12489 ( n6900 , n4844 , n985 );
    and g12490 ( n7573 , n12092 , n9271 );
    or g12491 ( n4632 , n6711 , n8061 );
    nor g12492 ( n7538 , n12254 , n3610 );
    and g12493 ( n2828 , n10166 , n14471 );
    and g12494 ( n5688 , n5317 , n14067 );
    and g12495 ( n4569 , n10822 , n3114 );
    not g12496 ( n1361 , n8073 );
    or g12497 ( n8600 , n2272 , n9783 );
    or g12498 ( n3781 , n4741 , n12230 );
    and g12499 ( n1297 , n11816 , n10066 );
    or g12500 ( n934 , n3132 , n8759 );
    or g12501 ( n5754 , n5815 , n13694 );
    or g12502 ( n12126 , n5640 , n12614 );
    and g12503 ( n2550 , n12802 , n13652 );
    and g12504 ( n1273 , n13489 , n9485 );
    or g12505 ( n14268 , n5562 , n4377 );
    or g12506 ( n4914 , n14449 , n318 );
    and g12507 ( n6244 , n5475 , n8399 );
    and g12508 ( n4206 , n11607 , n3525 );
    or g12509 ( n12894 , n100 , n3837 );
    nor g12510 ( n6944 , n911 , n5469 );
    or g12511 ( n6520 , n1776 , n13102 );
    or g12512 ( n1634 , n6205 , n12267 );
    nor g12513 ( n8591 , n10715 , n651 );
    nor g12514 ( n6423 , n14198 , n5368 );
    and g12515 ( n3814 , n10589 , n7264 );
    and g12516 ( n5702 , n1946 , n1705 );
    or g12517 ( n11272 , n10383 , n3988 );
    or g12518 ( n2469 , n13806 , n9467 );
    or g12519 ( n12362 , n2877 , n14331 );
    nor g12520 ( n3823 , n1178 , n11410 );
    and g12521 ( n11520 , n5279 , n3489 );
    and g12522 ( n10193 , n13236 , n14418 );
    and g12523 ( n8346 , n457 , n7956 );
    and g12524 ( n3564 , n1610 , n11164 );
    not g12525 ( n9583 , n13593 );
    or g12526 ( n2870 , n12100 , n7092 );
    or g12527 ( n1192 , n7700 , n6636 );
    not g12528 ( n5007 , n10069 );
    and g12529 ( n9858 , n2820 , n9366 );
    or g12530 ( n546 , n10351 , n9736 );
    and g12531 ( n1376 , n12611 , n8004 );
    and g12532 ( n8144 , n8780 , n6897 );
    or g12533 ( n10877 , n10309 , n1847 );
    or g12534 ( n10957 , n1258 , n1531 );
    nor g12535 ( n4663 , n6426 , n6567 );
    and g12536 ( n10567 , n10015 , n11591 );
    or g12537 ( n5259 , n6595 , n11589 );
    or g12538 ( n1737 , n10936 , n78 );
    or g12539 ( n11997 , n13130 , n9131 );
    and g12540 ( n8640 , n7970 , n7615 );
    not g12541 ( n14404 , n2918 );
    nor g12542 ( n803 , n6018 , n10653 );
    and g12543 ( n10867 , n8066 , n4630 );
    and g12544 ( n6009 , n10302 , n3128 );
    and g12545 ( n1956 , n5011 , n51 );
    or g12546 ( n2779 , n14058 , n14426 );
    and g12547 ( n4935 , n6527 , n8203 );
    not g12548 ( n13847 , n3021 );
    not g12549 ( n13084 , n8656 );
    and g12550 ( n8515 , n4790 , n4189 );
    and g12551 ( n2734 , n6703 , n11805 );
    or g12552 ( n13553 , n3569 , n12915 );
    and g12553 ( n8320 , n8300 , n9483 );
    and g12554 ( n2371 , n494 , n12111 );
    or g12555 ( n8107 , n12695 , n14141 );
    nor g12556 ( n522 , n7011 , n11994 );
    or g12557 ( n3965 , n2857 , n5239 );
    or g12558 ( n2748 , n7156 , n12498 );
    and g12559 ( n14265 , n10302 , n12343 );
    and g12560 ( n1814 , n3204 , n2755 );
    and g12561 ( n7204 , n6130 , n4532 );
    and g12562 ( n13821 , n4788 , n2789 );
    and g12563 ( n3600 , n718 , n14233 );
    or g12564 ( n6554 , n12933 , n5502 );
    or g12565 ( n13370 , n1628 , n8464 );
    not g12566 ( n13676 , n6975 );
    and g12567 ( n6881 , n14321 , n13926 );
    not g12568 ( n5197 , n1861 );
    not g12569 ( n14058 , n4606 );
    nor g12570 ( n3439 , n7940 , n1501 );
    or g12571 ( n12063 , n5562 , n4051 );
    not g12572 ( n13139 , n3544 );
    and g12573 ( n5681 , n5012 , n7793 );
    or g12574 ( n11016 , n4601 , n14483 );
    or g12575 ( n7930 , n6288 , n14429 );
    not g12576 ( n10568 , n10239 );
    not g12577 ( n3586 , n10303 );
    and g12578 ( n4069 , n2709 , n2450 );
    nor g12579 ( n2024 , n8629 , n1513 );
    and g12580 ( n734 , n7211 , n12420 );
    or g12581 ( n9587 , n494 , n11345 );
    and g12582 ( n1591 , n1266 , n5466 );
    and g12583 ( n10801 , n1920 , n13968 );
    not g12584 ( n6747 , n13230 );
    nor g12585 ( n3410 , n13021 , n8483 );
    or g12586 ( n5482 , n1538 , n3803 );
    and g12587 ( n4986 , n8453 , n9005 );
    or g12588 ( n1970 , n12130 , n11646 );
    nor g12589 ( n3970 , n3434 , n7314 );
    not g12590 ( n4144 , n11412 );
    and g12591 ( n5704 , n7670 , n5769 );
    and g12592 ( n11931 , n11569 , n658 );
    and g12593 ( n11696 , n5918 , n9831 );
    not g12594 ( n12764 , n9371 );
    and g12595 ( n4230 , n6192 , n10151 );
    not g12596 ( n10710 , n5675 );
    and g12597 ( n2926 , n13252 , n5686 );
    or g12598 ( n7979 , n13840 , n10630 );
    or g12599 ( n10745 , n11580 , n13101 );
    nor g12600 ( n12718 , n1677 , n10567 );
    and g12601 ( n6065 , n536 , n9364 );
    or g12602 ( n1621 , n3126 , n667 );
    nor g12603 ( n13910 , n7229 , n1712 );
    and g12604 ( n11954 , n79 , n5478 );
    and g12605 ( n242 , n8393 , n8835 );
    nor g12606 ( n6565 , n8592 , n1392 );
    and g12607 ( n6499 , n2709 , n5831 );
    or g12608 ( n5925 , n2246 , n3197 );
    and g12609 ( n7305 , n8250 , n10827 );
    or g12610 ( n7722 , n7678 , n9600 );
    and g12611 ( n12448 , n748 , n5751 );
    nor g12612 ( n12120 , n6743 , n6457 );
    not g12613 ( n4357 , n1966 );
    nor g12614 ( n3252 , n9414 , n8829 );
    nor g12615 ( n7386 , n5833 , n5937 );
    not g12616 ( n9890 , n12970 );
    or g12617 ( n10201 , n1548 , n2009 );
    and g12618 ( n417 , n14358 , n4724 );
    or g12619 ( n11162 , n8747 , n7705 );
    or g12620 ( n6870 , n13707 , n5326 );
    or g12621 ( n7807 , n954 , n765 );
    and g12622 ( n6079 , n6957 , n4605 );
    not g12623 ( n11403 , n7660 );
    and g12624 ( n6489 , n7053 , n4882 );
    or g12625 ( n11164 , n10234 , n3504 );
    not g12626 ( n5940 , n3440 );
    and g12627 ( n6805 , n5252 , n4335 );
    not g12628 ( n646 , n11861 );
    and g12629 ( n12650 , n2006 , n8654 );
    not g12630 ( n7192 , n1421 );
    and g12631 ( n6110 , n5940 , n6360 );
    and g12632 ( n14372 , n12857 , n9594 );
    and g12633 ( n13472 , n5012 , n6869 );
    and g12634 ( n9097 , n10247 , n4869 );
    or g12635 ( n6869 , n9140 , n2956 );
    or g12636 ( n9976 , n4180 , n13381 );
    or g12637 ( n8539 , n1820 , n1591 );
    and g12638 ( n7813 , n1729 , n2363 );
    and g12639 ( n13462 , n11300 , n3474 );
    nor g12640 ( n3774 , n9924 , n4064 );
    nor g12641 ( n6456 , n11980 , n3145 );
    and g12642 ( n8955 , n309 , n12124 );
    nor g12643 ( n9799 , n1628 , n7742 );
    and g12644 ( n11317 , n6389 , n7 );
    or g12645 ( n8435 , n7736 , n13727 );
    and g12646 ( n8775 , n3586 , n13856 );
    nor g12647 ( n4375 , n448 , n14246 );
    or g12648 ( n10482 , n1623 , n6125 );
    nor g12649 ( n6400 , n14166 , n1791 );
    not g12650 ( n12820 , n12249 );
    nor g12651 ( n12238 , n14455 , n10344 );
    or g12652 ( n11550 , n3125 , n6073 );
    or g12653 ( n5056 , n4978 , n7206 );
    or g12654 ( n10860 , n14466 , n3181 );
    not g12655 ( n8702 , n14367 );
    and g12656 ( n8241 , n10166 , n4726 );
    and g12657 ( n8022 , n80 , n11700 );
    not g12658 ( n12930 , n7915 );
    and g12659 ( n9517 , n6625 , n109 );
    or g12660 ( n11066 , n7818 , n5014 );
    nor g12661 ( n8621 , n12311 , n10180 );
    nor g12662 ( n11116 , n6397 , n13193 );
    not g12663 ( n4216 , n11428 );
    or g12664 ( n1325 , n2908 , n1841 );
    or g12665 ( n7633 , n6595 , n995 );
    or g12666 ( n5594 , n9856 , n4230 );
    or g12667 ( n2287 , n9151 , n12805 );
    not g12668 ( n7810 , n2619 );
    and g12669 ( n8709 , n3276 , n6506 );
    or g12670 ( n7838 , n4698 , n394 );
    and g12671 ( n5085 , n3755 , n9929 );
    and g12672 ( n6776 , n6525 , n7176 );
    and g12673 ( n13232 , n3923 , n8105 );
    not g12674 ( n5471 , n10177 );
    or g12675 ( n4406 , n14029 , n4842 );
    and g12676 ( n3897 , n11679 , n1684 );
    not g12677 ( n5491 , n5627 );
    or g12678 ( n4402 , n4876 , n13007 );
    or g12679 ( n11906 , n11285 , n6296 );
    or g12680 ( n6704 , n10289 , n4563 );
    and g12681 ( n7983 , n12057 , n9362 );
    or g12682 ( n9794 , n13155 , n11304 );
    not g12683 ( n10822 , n10322 );
    and g12684 ( n10759 , n2942 , n9413 );
    and g12685 ( n359 , n3043 , n4601 );
    and g12686 ( n8244 , n898 , n9325 );
    or g12687 ( n13549 , n13531 , n13172 );
    or g12688 ( n2238 , n10933 , n11623 );
    and g12689 ( n10762 , n5252 , n14387 );
    or g12690 ( n2410 , n9174 , n8253 );
    or g12691 ( n8263 , n7116 , n4446 );
    or g12692 ( n7098 , n10960 , n11559 );
    or g12693 ( n4420 , n7462 , n12906 );
    and g12694 ( n13560 , n14357 , n12272 );
    nor g12695 ( n2191 , n7364 , n186 );
    nor g12696 ( n6828 , n12117 , n3199 );
    or g12697 ( n3976 , n1801 , n10912 );
    or g12698 ( n3420 , n12034 , n11257 );
    and g12699 ( n11191 , n8372 , n13392 );
    not g12700 ( n12759 , n9878 );
    not g12701 ( n687 , n12503 );
    not g12702 ( n4840 , n10889 );
    nor g12703 ( n10934 , n1844 , n4503 );
    or g12704 ( n2903 , n13854 , n6348 );
    not g12705 ( n2087 , n8288 );
    and g12706 ( n12161 , n5553 , n684 );
    or g12707 ( n12926 , n5432 , n10858 );
    or g12708 ( n267 , n5695 , n13465 );
    not g12709 ( n9818 , n13047 );
    or g12710 ( n8673 , n12169 , n1960 );
    or g12711 ( n9132 , n2857 , n4240 );
    or g12712 ( n13290 , n1602 , n14269 );
    and g12713 ( n156 , n2058 , n5481 );
    or g12714 ( n10291 , n11315 , n13743 );
    or g12715 ( n1566 , n766 , n14394 );
    and g12716 ( n1927 , n8737 , n7252 );
    or g12717 ( n11571 , n2761 , n4501 );
    not g12718 ( n12695 , n11813 );
    and g12719 ( n4418 , n13572 , n13654 );
    nor g12720 ( n5392 , n4978 , n740 );
    nor g12721 ( n10109 , n2889 , n7536 );
    or g12722 ( n13739 , n4828 , n13286 );
    not g12723 ( n8066 , n1911 );
    and g12724 ( n8333 , n2099 , n797 );
    and g12725 ( n10382 , n14388 , n5052 );
    or g12726 ( n11022 , n8969 , n10694 );
    or g12727 ( n14043 , n8151 , n9523 );
    and g12728 ( n3637 , n10820 , n4519 );
    or g12729 ( n13832 , n9375 , n1586 );
    or g12730 ( n12497 , n5562 , n9056 );
    and g12731 ( n13592 , n8965 , n2039 );
    not g12732 ( n11459 , n81 );
    or g12733 ( n4560 , n7076 , n3232 );
    and g12734 ( n10215 , n13407 , n11579 );
    and g12735 ( n7875 , n3765 , n5149 );
    or g12736 ( n11281 , n3546 , n13076 );
    and g12737 ( n14204 , n1361 , n303 );
    or g12738 ( n440 , n5132 , n14267 );
    not g12739 ( n5042 , n3461 );
    not g12740 ( n7362 , n8106 );
    not g12741 ( n5458 , n5525 );
    and g12742 ( n9178 , n3785 , n8295 );
    or g12743 ( n6652 , n12324 , n10152 );
    not g12744 ( n2684 , n4216 );
    or g12745 ( n1175 , n12622 , n1030 );
    nor g12746 ( n4792 , n648 , n1672 );
    and g12747 ( n2327 , n12935 , n121 );
    not g12748 ( n6343 , n12930 );
    not g12749 ( n8920 , n4007 );
    and g12750 ( n9645 , n1904 , n2511 );
    or g12751 ( n13971 , n11722 , n9463 );
    and g12752 ( n3012 , n14321 , n2096 );
    nor g12753 ( n2950 , n9657 , n3670 );
    or g12754 ( n2300 , n6046 , n13802 );
    not g12755 ( n3802 , n9350 );
    and g12756 ( n3966 , n9190 , n7537 );
    or g12757 ( n9287 , n8304 , n11335 );
    nor g12758 ( n9359 , n6326 , n12749 );
    not g12759 ( n2090 , n74 );
    nor g12760 ( n4793 , n7056 , n2871 );
    or g12761 ( n10845 , n7229 , n10632 );
    and g12762 ( n9338 , n1193 , n11948 );
    not g12763 ( n12453 , n12088 );
    and g12764 ( n3862 , n13338 , n11383 );
    and g12765 ( n2097 , n11674 , n1915 );
    not g12766 ( n787 , n3506 );
    nor g12767 ( n11924 , n648 , n1509 );
    and g12768 ( n10185 , n14260 , n9012 );
    or g12769 ( n4260 , n9226 , n655 );
    or g12770 ( n8193 , n10626 , n1629 );
    and g12771 ( n8568 , n2709 , n9899 );
    and g12772 ( n4674 , n4614 , n5198 );
    or g12773 ( n8256 , n2098 , n1871 );
    and g12774 ( n8130 , n9265 , n7849 );
    not g12775 ( n7507 , n13544 );
    and g12776 ( n1091 , n11636 , n1725 );
    nor g12777 ( n4818 , n13977 , n9087 );
    or g12778 ( n3188 , n976 , n7070 );
    or g12779 ( n3505 , n11510 , n823 );
    and g12780 ( n628 , n9272 , n12694 );
    nor g12781 ( n2344 , n3959 , n10456 );
    nor g12782 ( n302 , n9546 , n13996 );
    not g12783 ( n1198 , n9686 );
    or g12784 ( n12890 , n4481 , n6076 );
    or g12785 ( n8844 , n1198 , n12517 );
    or g12786 ( n4041 , n13080 , n11853 );
    nor g12787 ( n9685 , n5904 , n8970 );
    not g12788 ( n12533 , n12117 );
    not g12789 ( n619 , n4609 );
    or g12790 ( n9960 , n77 , n3387 );
    not g12791 ( n12292 , n12106 );
    nor g12792 ( n10848 , n11094 , n9458 );
    and g12793 ( n6036 , n8007 , n11698 );
    or g12794 ( n5352 , n9984 , n14240 );
    nor g12795 ( n247 , n1813 , n10321 );
    or g12796 ( n12352 , n6706 , n1622 );
    and g12797 ( n7025 , n3097 , n10482 );
    not g12798 ( n9567 , n11302 );
    not g12799 ( n12494 , n6804 );
    and g12800 ( n2517 , n3424 , n5632 );
    or g12801 ( n10946 , n9541 , n108 );
    or g12802 ( n11864 , n12844 , n5168 );
    not g12803 ( n14510 , n3577 );
    and g12804 ( n7520 , n6354 , n2535 );
    not g12805 ( n9751 , n4248 );
    or g12806 ( n2702 , n4923 , n9903 );
    or g12807 ( n4620 , n4561 , n9810 );
    and g12808 ( n9076 , n7670 , n12317 );
    and g12809 ( n9290 , n13464 , n1424 );
    or g12810 ( n5995 , n3126 , n3597 );
    and g12811 ( n4666 , n6311 , n10844 );
    not g12812 ( n10589 , n8048 );
    or g12813 ( n3194 , n7436 , n8641 );
    or g12814 ( n1144 , n8575 , n3725 );
    and g12815 ( n3954 , n6625 , n5223 );
    nor g12816 ( n10737 , n573 , n8006 );
    not g12817 ( n1203 , n2674 );
    and g12818 ( n2394 , n14260 , n12541 );
    or g12819 ( n2304 , n9742 , n1133 );
    and g12820 ( n13237 , n3607 , n10 );
    nor g12821 ( n2929 , n9557 , n9215 );
    not g12822 ( n2843 , n1966 );
    or g12823 ( n12914 , n4898 , n11673 );
    or g12824 ( n7463 , n10871 , n11314 );
    nor g12825 ( n9087 , n5569 , n3305 );
    and g12826 ( n8114 , n13407 , n5547 );
    not g12827 ( n2470 , n1473 );
    or g12828 ( n2542 , n8480 , n10943 );
    and g12829 ( n10687 , n8183 , n10064 );
    not g12830 ( n177 , n3652 );
    not g12831 ( n9920 , n2889 );
    or g12832 ( n6178 , n14366 , n2214 );
    nor g12833 ( n852 , n3882 , n5250 );
    or g12834 ( n2254 , n9422 , n14084 );
    or g12835 ( n5749 , n523 , n7884 );
    and g12836 ( n2270 , n1788 , n10296 );
    and g12837 ( n5344 , n965 , n768 );
    not g12838 ( n10933 , n4720 );
    nor g12839 ( n1733 , n13310 , n11024 );
    or g12840 ( n353 , n12576 , n6487 );
    or g12841 ( n9391 , n12494 , n2957 );
    or g12842 ( n11430 , n13485 , n9445 );
    and g12843 ( n7236 , n14465 , n2466 );
    and g12844 ( n4927 , n14109 , n4669 );
    and g12845 ( n3614 , n12918 , n2046 );
    and g12846 ( n8152 , n8250 , n10489 );
    or g12847 ( n12308 , n10059 , n5225 );
    and g12848 ( n926 , n1255 , n6233 );
    or g12849 ( n193 , n3193 , n10436 );
    nor g12850 ( n11051 , n6039 , n1185 );
    nor g12851 ( n3488 , n9618 , n5577 );
    or g12852 ( n11385 , n6023 , n13814 );
    not g12853 ( n3886 , n4149 );
    or g12854 ( n7718 , n6373 , n11274 );
    or g12855 ( n7648 , n12759 , n9966 );
    not g12856 ( n10977 , n13437 );
    nor g12857 ( n1107 , n10479 , n14026 );
    not g12858 ( n5240 , n11969 );
    or g12859 ( n13680 , n14337 , n10345 );
    or g12860 ( n2377 , n13083 , n3629 );
    or g12861 ( n975 , n6695 , n13098 );
    or g12862 ( n11973 , n6263 , n4362 );
    not g12863 ( n11328 , n11345 );
    not g12864 ( n2969 , n5001 );
    or g12865 ( n4905 , n3877 , n13548 );
    and g12866 ( n7482 , n11674 , n10612 );
    or g12867 ( n9974 , n10626 , n6618 );
    and g12868 ( n14347 , n4581 , n13951 );
    and g12869 ( n13609 , n5764 , n6168 );
    or g12870 ( n12443 , n9716 , n2862 );
    not g12871 ( n14145 , n3428 );
    not g12872 ( n6192 , n3440 );
    or g12873 ( n8913 , n9541 , n741 );
    or g12874 ( n13938 , n11379 , n4839 );
    nor g12875 ( n2664 , n2729 , n12515 );
    not g12876 ( n12694 , n12097 );
    or g12877 ( n12104 , n2877 , n6225 );
    not g12878 ( n6706 , n10889 );
    or g12879 ( n8399 , n1844 , n10676 );
    or g12880 ( n4556 , n1383 , n2104 );
    and g12881 ( n4598 , n5471 , n5305 );
    not g12882 ( n6113 , n5631 );
    not g12883 ( n8111 , n2958 );
    and g12884 ( n13333 , n10072 , n9050 );
    not g12885 ( n3888 , n11152 );
    or g12886 ( n8179 , n8812 , n12012 );
    or g12887 ( n7 , n9229 , n8380 );
    or g12888 ( n11923 , n3815 , n11211 );
    or g12889 ( n1400 , n11510 , n11699 );
    or g12890 ( n2173 , n1223 , n7581 );
    and g12891 ( n7195 , n10668 , n2362 );
    and g12892 ( n4301 , n1854 , n7776 );
    and g12893 ( n9999 , n10589 , n10841 );
    or g12894 ( n2833 , n1044 , n2221 );
    or g12895 ( n11216 , n4033 , n6036 );
    nor g12896 ( n13980 , n11251 , n9292 );
    or g12897 ( n13539 , n3675 , n12321 );
    or g12898 ( n11052 , n1946 , n5950 );
    not g12899 ( n11503 , n6765 );
    and g12900 ( n6955 , n3276 , n12095 );
    and g12901 ( n10527 , n5764 , n3301 );
    and g12902 ( n12103 , n5188 , n22 );
    and g12903 ( n4263 , n12229 , n2592 );
    not g12904 ( n263 , n4154 );
    and g12905 ( n1016 , n4261 , n6414 );
    nor g12906 ( n9215 , n14370 , n13894 );
    and g12907 ( n6910 , n6486 , n4638 );
    nor g12908 ( n5364 , n9984 , n12865 );
    not g12909 ( n5312 , n13139 );
    and g12910 ( n12635 , n6957 , n7861 );
    or g12911 ( n9227 , n5468 , n4974 );
    nor g12912 ( n13672 , n3546 , n3272 );
    or g12913 ( n3585 , n2510 , n3195 );
    or g12914 ( n10031 , n10383 , n4077 );
    not g12915 ( n2901 , n11788 );
    or g12916 ( n2499 , n4899 , n12048 );
    or g12917 ( n4013 , n791 , n13008 );
    and g12918 ( n3131 , n9509 , n10703 );
    or g12919 ( n6149 , n747 , n2670 );
    or g12920 ( n2818 , n2089 , n1878 );
    and g12921 ( n6540 , n1140 , n8976 );
    or g12922 ( n2392 , n2857 , n1919 );
    and g12923 ( n3817 , n10512 , n1508 );
    and g12924 ( n1633 , n9198 , n7505 );
    not g12925 ( n4650 , n13561 );
    or g12926 ( n11340 , n13310 , n4892 );
    and g12927 ( n5653 , n5229 , n6330 );
    and g12928 ( n2978 , n1962 , n13056 );
    or g12929 ( n5049 , n1711 , n6287 );
    or g12930 ( n4269 , n11621 , n8707 );
    or g12931 ( n9549 , n8983 , n8157 );
    or g12932 ( n5813 , n5468 , n9351 );
    not g12933 ( n5948 , n9950 );
    or g12934 ( n14192 , n13118 , n11460 );
    and g12935 ( n2291 , n9564 , n13685 );
    and g12936 ( n5753 , n7057 , n11983 );
    not g12937 ( n10136 , n751 );
    or g12938 ( n9000 , n8748 , n13556 );
    and g12939 ( n6560 , n4276 , n259 );
    or g12940 ( n8163 , n8112 , n13231 );
    or g12941 ( n5067 , n3914 , n10215 );
    or g12942 ( n9244 , n7803 , n10656 );
    and g12943 ( n10423 , n2474 , n8311 );
    and g12944 ( n9502 , n4018 , n3352 );
    not g12945 ( n1261 , n3616 );
    and g12946 ( n1874 , n13362 , n5522 );
    and g12947 ( n321 , n7810 , n3836 );
    or g12948 ( n7395 , n12209 , n13224 );
    and g12949 ( n3733 , n3277 , n9998 );
    or g12950 ( n10853 , n3076 , n10169 );
    or g12951 ( n10873 , n1198 , n4558 );
    or g12952 ( n357 , n13547 , n13169 );
    or g12953 ( n6561 , n12764 , n13151 );
    and g12954 ( n1963 , n2669 , n12781 );
    nor g12955 ( n12988 , n14524 , n5177 );
    and g12956 ( n14050 , n8697 , n3840 );
    not g12957 ( n8252 , n8463 );
    and g12958 ( n13289 , n1526 , n7885 );
    and g12959 ( n10380 , n6981 , n13566 );
    and g12960 ( n4111 , n14042 , n5073 );
    and g12961 ( n6250 , n9885 , n10756 );
    nor g12962 ( n11512 , n6062 , n13443 );
    or g12963 ( n645 , n11510 , n10264 );
    nor g12964 ( n287 , n10091 , n12119 );
    or g12965 ( n10195 , n13516 , n2347 );
    or g12966 ( n14329 , n7700 , n2665 );
    nor g12967 ( n4110 , n1522 , n13306 );
    not g12968 ( n747 , n12489 );
    and g12969 ( n70 , n5823 , n11889 );
    nor g12970 ( n8249 , n1378 , n3148 );
    and g12971 ( n9084 , n4932 , n8815 );
    and g12972 ( n7458 , n1254 , n10056 );
    and g12973 ( n6689 , n13464 , n11502 );
    nor g12974 ( n8006 , n1575 , n3089 );
    and g12975 ( n793 , n3923 , n3327 );
    not g12976 ( n11285 , n9453 );
    or g12977 ( n419 , n7684 , n6645 );
    and g12978 ( n13409 , n12018 , n14137 );
    or g12979 ( n364 , n1137 , n1551 );
    nor g12980 ( n3158 , n7418 , n297 );
    nor g12981 ( n2010 , n10280 , n1530 );
    or g12982 ( n12068 , n3120 , n7623 );
    not g12983 ( n8015 , n1894 );
    not g12984 ( n6690 , n6332 );
    or g12985 ( n11735 , n1383 , n10717 );
    not g12986 ( n12549 , n2383 );
    not g12987 ( n2923 , n10801 );
    nor g12988 ( n14243 , n2236 , n1595 );
    or g12989 ( n8392 , n10035 , n4294 );
    and g12990 ( n5584 , n10767 , n10530 );
    and g12991 ( n439 , n10357 , n3693 );
    and g12992 ( n9823 , n4346 , n2886 );
    nor g12993 ( n7631 , n12200 , n1756 );
    or g12994 ( n13473 , n11818 , n1561 );
    nor g12995 ( n8201 , n7364 , n8691 );
    or g12996 ( n13738 , n2686 , n1717 );
    and g12997 ( n105 , n12730 , n11139 );
    and g12998 ( n7763 , n13147 , n1000 );
    and g12999 ( n2934 , n11016 , n3875 );
    and g13000 ( n12184 , n12404 , n4338 );
    and g13001 ( n5179 , n7026 , n8429 );
    nor g13002 ( n11560 , n13627 , n6565 );
    or g13003 ( n5107 , n12401 , n8485 );
    and g13004 ( n9570 , n4172 , n1107 );
    or g13005 ( n5039 , n12601 , n10524 );
    or g13006 ( n11819 , n8517 , n4528 );
    or g13007 ( n1209 , n4631 , n2134 );
    nor g13008 ( n3797 , n3019 , n10542 );
    and g13009 ( n11886 , n10622 , n6289 );
    and g13010 ( n8679 , n10332 , n192 );
    and g13011 ( n5565 , n11636 , n9702 );
    not g13012 ( n3313 , n4991 );
    and g13013 ( n1349 , n12918 , n4826 );
    or g13014 ( n663 , n11315 , n12594 );
    or g13015 ( n2260 , n7418 , n11442 );
    nor g13016 ( n5932 , n2731 , n6298 );
    not g13017 ( n12832 , n12757 );
    nor g13018 ( n4108 , n9807 , n12936 );
    and g13019 ( n9267 , n8393 , n833 );
    or g13020 ( n14516 , n14029 , n4467 );
    or g13021 ( n9159 , n8096 , n1173 );
    and g13022 ( n13448 , n9198 , n10961 );
    or g13023 ( n1747 , n10083 , n4721 );
    nor g13024 ( n2646 , n7887 , n3156 );
    or g13025 ( n11857 , n7430 , n10680 );
    nor g13026 ( n14174 , n4424 , n8153 );
    or g13027 ( n5768 , n9804 , n1227 );
    and g13028 ( n5913 , n11569 , n14484 );
    and g13029 ( n4126 , n2006 , n2421 );
    and g13030 ( n14331 , n5926 , n3319 );
    or g13031 ( n1829 , n5144 , n4804 );
    or g13032 ( n8313 , n6085 , n2107 );
    or g13033 ( n6213 , n2412 , n8805 );
    not g13034 ( n7346 , n14406 );
    and g13035 ( n11825 , n1431 , n2819 );
    not g13036 ( n9198 , n3402 );
    not g13037 ( n11379 , n565 );
    or g13038 ( n11077 , n10083 , n5580 );
    nor g13039 ( n4984 , n8557 , n5756 );
    and g13040 ( n12655 , n9275 , n2593 );
    and g13041 ( n13749 , n4244 , n7672 );
    and g13042 ( n10103 , n8111 , n775 );
    nor g13043 ( n3658 , n2597 , n6677 );
    nor g13044 ( n2245 , n1262 , n2947 );
    or g13045 ( n4638 , n11580 , n12748 );
    or g13046 ( n6190 , n14404 , n9850 );
    or g13047 ( n1285 , n5710 , n7995 );
    or g13048 ( n10217 , n12759 , n3154 );
    and g13049 ( n7542 , n10332 , n2112 );
    and g13050 ( n1880 , n5088 , n13711 );
    and g13051 ( n8409 , n3942 , n9462 );
    and g13052 ( n12052 , n9102 , n12657 );
    or g13053 ( n8958 , n6205 , n3855 );
    and g13054 ( n8229 , n8213 , n8539 );
    nor g13055 ( n18 , n13707 , n580 );
    not g13056 ( n4684 , n12746 );
    or g13057 ( n9781 , n5710 , n95 );
    and g13058 ( n2413 , n7810 , n12890 );
    or g13059 ( n1532 , n9269 , n8078 );
    or g13060 ( n1003 , n10512 , n6873 );
    or g13061 ( n1647 , n8714 , n2210 );
    nor g13062 ( n10597 , n4535 , n14290 );
    or g13063 ( n3050 , n1613 , n11270 );
    and g13064 ( n12600 , n13096 , n3662 );
    and g13065 ( n13133 , n5312 , n13785 );
    and g13066 ( n12045 , n9724 , n3031 );
    and g13067 ( n278 , n12025 , n123 );
    or g13068 ( n4067 , n8817 , n5184 );
    or g13069 ( n7666 , n13112 , n12367 );
    nor g13070 ( n2209 , n6122 , n4093 );
    and g13071 ( n9611 , n10619 , n2001 );
    or g13072 ( n2803 , n2694 , n3432 );
    and g13073 ( n8341 , n7818 , n9792 );
    or g13074 ( n1021 , n7358 , n5890 );
    and g13075 ( n13904 , n10332 , n9244 );
    not g13076 ( n3755 , n6119 );
    and g13077 ( n732 , n1231 , n6691 );
    or g13078 ( n14486 , n2179 , n8960 );
    and g13079 ( n796 , n12335 , n12360 );
    or g13080 ( n754 , n13806 , n5358 );
    and g13081 ( n8695 , n13900 , n931 );
    not g13082 ( n11309 , n14219 );
    and g13083 ( n5656 , n12229 , n8673 );
    and g13084 ( n128 , n13103 , n11530 );
    or g13085 ( n8884 , n9008 , n8002 );
    and g13086 ( n1311 , n8907 , n11490 );
    nor g13087 ( n7277 , n194 , n1246 );
    or g13088 ( n14025 , n13875 , n1468 );
    nor g13089 ( n1790 , n8527 , n14500 );
    or g13090 ( n2356 , n10331 , n8120 );
    or g13091 ( n5693 , n8881 , n3588 );
    and g13092 ( n11352 , n7026 , n2023 );
    or g13093 ( n10923 , n3025 , n7445 );
    and g13094 ( n4681 , n5459 , n3974 );
    and g13095 ( n11419 , n12615 , n7706 );
    and g13096 ( n997 , n3485 , n8652 );
    and g13097 ( n8664 , n2082 , n11894 );
    and g13098 ( n13607 , n1775 , n2903 );
    or g13099 ( n4020 , n9353 , n13804 );
    not g13100 ( n3958 , n1268 );
    nor g13101 ( n14311 , n8816 , n3557 );
    not g13102 ( n3497 , n7676 );
    or g13103 ( n7123 , n10624 , n12338 );
    and g13104 ( n10851 , n10367 , n10356 );
    and g13105 ( n9219 , n7810 , n1471 );
    and g13106 ( n2812 , n200 , n10494 );
    and g13107 ( n4249 , n1117 , n4044 );
    nor g13108 ( n13279 , n11558 , n6833 );
    and g13109 ( n1333 , n9920 , n12437 );
    and g13110 ( n3764 , n13096 , n14244 );
    or g13111 ( n443 , n6654 , n2538 );
    and g13112 ( n4457 , n5823 , n10216 );
    or g13113 ( n8994 , n1006 , n349 );
    not g13114 ( n4052 , n1060 );
    or g13115 ( n3327 , n11379 , n6224 );
    or g13116 ( n14201 , n2318 , n11365 );
    or g13117 ( n1873 , n12139 , n6410 );
    not g13118 ( n5587 , n12874 );
    or g13119 ( n8536 , n3559 , n11475 );
    or g13120 ( n4594 , n5807 , n6588 );
    or g13121 ( n2681 , n3062 , n12504 );
    not g13122 ( n10402 , n12088 );
    nor g13123 ( n8407 , n1299 , n379 );
    or g13124 ( n11652 , n13847 , n10783 );
    and g13125 ( n10642 , n12832 , n10956 );
    and g13126 ( n4294 , n4359 , n5310 );
    or g13127 ( n6422 , n11842 , n1222 );
    or g13128 ( n12653 , n6323 , n14165 );
    nor g13129 ( n13438 , n9078 , n10401 );
    and g13130 ( n11327 , n13246 , n8783 );
    not g13131 ( n703 , n6844 );
    or g13132 ( n10045 , n11231 , n14035 );
    and g13133 ( n1797 , n11814 , n12187 );
    and g13134 ( n2202 , n4502 , n9985 );
    or g13135 ( n1541 , n8172 , n5869 );
    or g13136 ( n704 , n5507 , n5644 );
    nor g13137 ( n8330 , n14332 , n3146 );
    nor g13138 ( n6897 , n10883 , n7857 );
    or g13139 ( n1014 , n3667 , n8824 );
    nor g13140 ( n6646 , n11546 , n12008 );
    not g13141 ( n5209 , n9236 );
    not g13142 ( n2780 , n10864 );
    and g13143 ( n3157 , n3212 , n10016 );
    and g13144 ( n5283 , n4788 , n10575 );
    not g13145 ( n7736 , n11813 );
    and g13146 ( n12586 , n5489 , n5094 );
    not g13147 ( n14401 , n14412 );
    or g13148 ( n13318 , n14472 , n158 );
    and g13149 ( n3943 , n5312 , n11181 );
    or g13150 ( n7688 , n8034 , n6396 );
    not g13151 ( n7179 , n2951 );
    nor g13152 ( n10431 , n12097 , n11490 );
    or g13153 ( n192 , n11420 , n11682 );
    and g13154 ( n8758 , n7670 , n4999 );
    or g13155 ( n7944 , n12633 , n4112 );
    or g13156 ( n4390 , n647 , n8366 );
    and g13157 ( n7827 , n10922 , n12794 );
    not g13158 ( n4899 , n11541 );
    and g13159 ( n8148 , n2791 , n2137 );
    nor g13160 ( n4278 , n2016 , n9560 );
    and g13161 ( n601 , n333 , n13664 );
    and g13162 ( n3663 , n6354 , n2833 );
    not g13163 ( n5762 , n7441 );
    and g13164 ( n1326 , n11163 , n5393 );
    or g13165 ( n12546 , n4791 , n7335 );
    nor g13166 ( n4096 , n9078 , n8359 );
    and g13167 ( n7387 , n2942 , n12263 );
    and g13168 ( n10608 , n4788 , n7174 );
    or g13169 ( n240 , n69 , n10970 );
    nor g13170 ( n4409 , n7887 , n9614 );
    and g13171 ( n12679 , n5088 , n3281 );
    nor g13172 ( n3296 , n14139 , n4132 );
    and g13173 ( n11058 , n5229 , n8661 );
    not g13174 ( n9305 , n885 );
    and g13175 ( n10057 , n5779 , n866 );
    and g13176 ( n11504 , n5062 , n3682 );
    and g13177 ( n5190 , n3942 , n10092 );
    nor g13178 ( n9498 , n2868 , n14488 );
    or g13179 ( n9512 , n9984 , n5957 );
    not g13180 ( n3904 , n12888 );
    and g13181 ( n8522 , n7068 , n8782 );
    and g13182 ( n9722 , n10374 , n7047 );
    not g13183 ( n4608 , n12086 );
    or g13184 ( n14257 , n6350 , n5 );
    and g13185 ( n12439 , n7419 , n12616 );
    or g13186 ( n4202 , n12651 , n13715 );
    not g13187 ( n9102 , n11548 );
    and g13188 ( n10594 , n2682 , n9130 );
    not g13189 ( n14461 , n8424 );
    or g13190 ( n8076 , n11011 , n4295 );
    and g13191 ( n2119 , n9198 , n761 );
    and g13192 ( n6643 , n6937 , n5256 );
    nor g13193 ( n9037 , n11990 , n14520 );
    nor g13194 ( n10290 , n10428 , n2943 );
    not g13195 ( n9323 , n5613 );
    and g13196 ( n2242 , n10854 , n1199 );
    not g13197 ( n5489 , n13360 );
    or g13198 ( n2549 , n4791 , n6784 );
    nor g13199 ( n11916 , n3768 , n11371 );
    or g13200 ( n5775 , n8908 , n2240 );
    nor g13201 ( n5585 , n2236 , n8158 );
    and g13202 ( n11466 , n13641 , n6129 );
    or g13203 ( n12102 , n1559 , n5077 );
    or g13204 ( n4964 , n9864 , n2169 );
    nor g13205 ( n7580 , n4572 , n928 );
    and g13206 ( n4466 , n4346 , n7766 );
    not g13207 ( n5847 , n11966 );
    and g13208 ( n751 , n4716 , n11938 );
    nor g13209 ( n3464 , n2241 , n5076 );
    or g13210 ( n1037 , n12494 , n9038 );
    nor g13211 ( n3610 , n13477 , n3466 );
    not g13212 ( n10406 , n7575 );
    not g13213 ( n11028 , n11232 );
    or g13214 ( n14425 , n227 , n13090 );
    and g13215 ( n10631 , n11614 , n384 );
    nor g13216 ( n12678 , n5065 , n12637 );
    and g13217 ( n9500 , n5137 , n913 );
    not g13218 ( n387 , n10985 );
    and g13219 ( n10524 , n536 , n11084 );
    and g13220 ( n4405 , n1193 , n10181 );
    or g13221 ( n2338 , n4925 , n10673 );
    not g13222 ( n2322 , n5675 );
    not g13223 ( n2272 , n11813 );
    and g13224 ( n12575 , n11867 , n3679 );
    and g13225 ( n7532 , n10815 , n5055 );
    or g13226 ( n8284 , n7678 , n8568 );
    and g13227 ( n4862 , n9315 , n13634 );
    and g13228 ( n6197 , n8300 , n9492 );
    and g13229 ( n11273 , n2310 , n9187 );
    or g13230 ( n5204 , n1728 , n13695 );
    and g13231 ( n12941 , n11316 , n3692 );
    or g13232 ( n12271 , n12712 , n6563 );
    and g13233 ( n13639 , n12927 , n1744 );
    and g13234 ( n1084 , n13404 , n12894 );
    or g13235 ( n2112 , n7803 , n10804 );
    or g13236 ( n110 , n3132 , n3797 );
    and g13237 ( n4997 , n11157 , n7773 );
    nor g13238 ( n2952 , n2154 , n11946 );
    or g13239 ( n8990 , n11839 , n9867 );
    nor g13240 ( n453 , n6933 , n4536 );
    or g13241 ( n5856 , n7308 , n14464 );
    and g13242 ( n14162 , n9853 , n632 );
    or g13243 ( n13773 , n11804 , n6322 );
    or g13244 ( n6717 , n8517 , n5907 );
    or g13245 ( n529 , n11839 , n12969 );
    not g13246 ( n13379 , n5795 );
    not g13247 ( n6350 , n5974 );
    and g13248 ( n9709 , n6609 , n4399 );
    and g13249 ( n13994 , n11300 , n11554 );
    and g13250 ( n4322 , n1489 , n12680 );
    or g13251 ( n6799 , n8210 , n7413 );
    and g13252 ( n12110 , n12998 , n10809 );
    and g13253 ( n6618 , n12335 , n6037 );
    or g13254 ( n12225 , n9353 , n3224 );
    and g13255 ( n10694 , n12038 , n92 );
    and g13256 ( n7222 , n1117 , n13884 );
    or g13257 ( n6154 , n2518 , n1294 );
    not g13258 ( n80 , n13723 );
    and g13259 ( n13460 , n9724 , n3747 );
    and g13260 ( n3046 , n3542 , n2850 );
    nor g13261 ( n13681 , n4195 , n6141 );
    and g13262 ( n4129 , n14373 , n3741 );
    and g13263 ( n8068 , n13363 , n5956 );
    not g13264 ( n8065 , n6159 );
    or g13265 ( n12319 , n7249 , n5301 );
    or g13266 ( n11841 , n4239 , n11476 );
    and g13267 ( n5147 , n4104 , n883 );
    or g13268 ( n566 , n14481 , n7220 );
    and g13269 ( n12773 , n12042 , n12880 );
    and g13270 ( n9651 , n7677 , n13943 );
    or g13271 ( n5859 , n11724 , n3850 );
    nor g13272 ( n11496 , n12112 , n8504 );
    and g13273 ( n4273 , n6167 , n6223 );
    not g13274 ( n5362 , n10069 );
    nor g13275 ( n10133 , n10649 , n10876 );
    nor g13276 ( n6590 , n2742 , n9652 );
    and g13277 ( n6608 , n13781 , n6727 );
    and g13278 ( n6598 , n3268 , n5121 );
    and g13279 ( n1547 , n12615 , n599 );
    or g13280 ( n11389 , n4033 , n7486 );
    and g13281 ( n8329 , n2310 , n8274 );
    and g13282 ( n13741 , n4276 , n12257 );
    and g13283 ( n821 , n8247 , n893 );
    or g13284 ( n8019 , n5253 , n1991 );
    or g13285 ( n2791 , n14252 , n4755 );
    and g13286 ( n8290 , n5348 , n2712 );
    or g13287 ( n1738 , n4340 , n13048 );
    and g13288 ( n6780 , n7427 , n12233 );
    nor g13289 ( n8628 , n12197 , n9115 );
    or g13290 ( n11049 , n954 , n10141 );
    nor g13291 ( n11131 , n3922 , n6449 );
    or g13292 ( n5495 , n504 , n591 );
    and g13293 ( n13425 , n9494 , n13116 );
    and g13294 ( n258 , n13421 , n8219 );
    not g13295 ( n13227 , n5871 );
    or g13296 ( n9998 , n13698 , n9379 );
    and g13297 ( n7393 , n225 , n12536 );
    nor g13298 ( n13740 , n7589 , n5098 );
    or g13299 ( n1184 , n6090 , n8758 );
    not g13300 ( n5294 , n9818 );
    and g13301 ( n13778 , n4692 , n2964 );
    or g13302 ( n14194 , n116 , n9060 );
    nor g13303 ( n4959 , n7352 , n6817 );
    or g13304 ( n13486 , n10062 , n14033 );
    or g13305 ( n9988 , n7430 , n128 );
    and g13306 ( n10214 , n14227 , n7780 );
    not g13307 ( n6193 , n5438 );
    nor g13308 ( n4645 , n12075 , n2663 );
    nor g13309 ( n3466 , n3210 , n3421 );
    or g13310 ( n1523 , n8969 , n8894 );
    and g13311 ( n8436 , n6157 , n5917 );
    and g13312 ( n6943 , n7943 , n7604 );
    nor g13313 ( n12431 , n7887 , n1033 );
    not g13314 ( n1006 , n1676 );
    or g13315 ( n4762 , n13446 , n3055 );
    and g13316 ( n3448 , n10705 , n7749 );
    and g13317 ( n7675 , n13745 , n3472 );
    and g13318 ( n112 , n11157 , n12792 );
    not g13319 ( n12886 , n7115 );
    and g13320 ( n13225 , n13464 , n11085 );
    not g13321 ( n12461 , n1784 );
    nor g13322 ( n5718 , n11305 , n8999 );
    and g13323 ( n13326 , n14465 , n9148 );
    not g13324 ( n8517 , n1220 );
    and g13325 ( n13568 , n7043 , n8669 );
    not g13326 ( n7375 , n11967 );
    and g13327 ( n502 , n12421 , n8797 );
    and g13328 ( n2107 , n12990 , n13396 );
    not g13329 ( n3877 , n9169 );
    and g13330 ( n12606 , n8950 , n301 );
    and g13331 ( n3339 , n2583 , n6610 );
    not g13332 ( n4742 , n10529 );
    not g13333 ( n7681 , n3280 );
    and g13334 ( n11417 , n12683 , n1837 );
    not g13335 ( n7957 , n9450 );
    or g13336 ( n2073 , n13659 , n12926 );
    nor g13337 ( n12423 , n474 , n12045 );
    or g13338 ( n8871 , n9864 , n7769 );
    or g13339 ( n5201 , n390 , n3773 );
    and g13340 ( n11883 , n5825 , n944 );
    or g13341 ( n11810 , n7551 , n2176 );
    and g13342 ( n1335 , n1489 , n14223 );
    or g13343 ( n755 , n12625 , n5169 );
    and g13344 ( n8198 , n14260 , n598 );
    not g13345 ( n4445 , n13003 );
    or g13346 ( n3776 , n11852 , n13000 );
    or g13347 ( n8537 , n11738 , n2615 );
    or g13348 ( n11483 , n5575 , n6745 );
    or g13349 ( n12835 , n782 , n6894 );
    and g13350 ( n3901 , n12573 , n11538 );
    or g13351 ( n7166 , n2318 , n11447 );
    or g13352 ( n4386 , n5647 , n13243 );
    or g13353 ( n6059 , n2055 , n5544 );
    not g13354 ( n7909 , n9416 );
    nor g13355 ( n10723 , n5209 , n12286 );
    or g13356 ( n4105 , n2061 , n9186 );
    or g13357 ( n598 , n1006 , n11670 );
    or g13358 ( n5318 , n2236 , n6474 );
    or g13359 ( n2886 , n6206 , n3179 );
    not g13360 ( n2758 , n10377 );
    and g13361 ( n11799 , n5312 , n10211 );
    or g13362 ( n3865 , n9289 , n14518 );
    nor g13363 ( n13085 , n717 , n11079 );
    nor g13364 ( n11535 , n10323 , n2115 );
    nor g13365 ( n8984 , n6907 , n522 );
    and g13366 ( n4414 , n11163 , n5787 );
    or g13367 ( n9750 , n13537 , n1171 );
    or g13368 ( n824 , n5253 , n5384 );
    or g13369 ( n1118 , n3099 , n6642 );
    or g13370 ( n14342 , n10560 , n12939 );
    and g13371 ( n2523 , n14260 , n12756 );
    or g13372 ( n2041 , n4953 , n13055 );
    or g13373 ( n2719 , n6607 , n11330 );
    nor g13374 ( n3874 , n8301 , n3937 );
    and g13375 ( n10326 , n9803 , n13091 );
    nor g13376 ( n341 , n12904 , n11624 );
    or g13377 ( n9319 , n4988 , n5816 );
    and g13378 ( n9038 , n2473 , n6916 );
    or g13379 ( n3389 , n4925 , n11381 );
    or g13380 ( n4250 , n1660 , n4453 );
    nor g13381 ( n2579 , n1462 , n11096 );
    and g13382 ( n7175 , n12531 , n13888 );
    and g13383 ( n4839 , n9345 , n6770 );
    or g13384 ( n9050 , n10294 , n1529 );
    and g13385 ( n310 , n11676 , n10232 );
    or g13386 ( n762 , n9226 , n5992 );
    or g13387 ( n3352 , n9140 , n3598 );
    and g13388 ( n224 , n2180 , n3790 );
    or g13389 ( n1015 , n4239 , n12895 );
    or g13390 ( n5258 , n10062 , n5269 );
    and g13391 ( n6399 , n2224 , n9689 );
    not g13392 ( n8162 , n13154 );
    not g13393 ( n13780 , n4270 );
    or g13394 ( n8666 , n12821 , n999 );
    and g13395 ( n8680 , n12935 , n1608 );
    and g13396 ( n1233 , n6167 , n1925 );
    and g13397 ( n2981 , n231 , n4504 );
    and g13398 ( n3629 , n5899 , n3852 );
    and g13399 ( n12174 , n14373 , n11284 );
    not g13400 ( n6794 , n10858 );
    not g13401 ( n1628 , n11541 );
    or g13402 ( n12297 , n3088 , n7467 );
    or g13403 ( n12399 , n10245 , n11136 );
    and g13404 ( n8824 , n7063 , n4074 );
    or g13405 ( n5742 , n11440 , n3948 );
    or g13406 ( n10170 , n555 , n9167 );
    or g13407 ( n12669 , n12414 , n207 );
    or g13408 ( n9098 , n5891 , n874 );
    nor g13409 ( n3510 , n6039 , n1327 );
    not g13410 ( n478 , n3455 );
    or g13411 ( n1165 , n11687 , n12336 );
    and g13412 ( n10228 , n327 , n7067 );
    nor g13413 ( n1595 , n9046 , n10548 );
    or g13414 ( n4878 , n14435 , n14379 );
    nor g13415 ( n4218 , n2098 , n5597 );
    and g13416 ( n3753 , n627 , n1995 );
    or g13417 ( n9660 , n10289 , n1158 );
    and g13418 ( n9169 , n7521 , n12279 );
    not g13419 ( n4404 , n3804 );
    not g13420 ( n11489 , n8162 );
    nor g13421 ( n14101 , n584 , n5540 );
    or g13422 ( n8387 , n11909 , n11333 );
    or g13423 ( n10514 , n6039 , n5370 );
    or g13424 ( n6936 , n3512 , n13966 );
    and g13425 ( n14235 , n1193 , n346 );
    or g13426 ( n5909 , n12934 , n2640 );
    and g13427 ( n6410 , n6343 , n14335 );
    not g13428 ( n911 , n13206 );
    not g13429 ( n1262 , n93 );
    and g13430 ( n14423 , n392 , n3630 );
    and g13431 ( n1723 , n1539 , n8335 );
    not g13432 ( n12569 , n264 );
    or g13433 ( n11889 , n12622 , n7222 );
    and g13434 ( n8181 , n3536 , n10250 );
    or g13435 ( n8976 , n14370 , n8117 );
    and g13436 ( n13768 , n11814 , n14405 );
    and g13437 ( n2129 , n4261 , n1206 );
    or g13438 ( n8743 , n766 , n10087 );
    or g13439 ( n2127 , n5472 , n2743 );
    or g13440 ( n8545 , n4357 , n7969 );
    and g13441 ( n6823 , n10710 , n3167 );
    or g13442 ( n9263 , n817 , n7616 );
    and g13443 ( n9167 , n11679 , n2849 );
    or g13444 ( n8159 , n13432 , n10125 );
    or g13445 ( n8793 , n6519 , n7231 );
    nor g13446 ( n11024 , n2005 , n2191 );
    and g13447 ( n4099 , n8692 , n11186 );
    nor g13448 ( n2044 , n2684 , n12670 );
    nor g13449 ( n10192 , n1262 , n11903 );
    and g13450 ( n6952 , n13109 , n12761 );
    and g13451 ( n12736 , n2669 , n7628 );
    and g13452 ( n5245 , n5459 , n12109 );
    not g13453 ( n7914 , n2934 );
    nor g13454 ( n792 , n14198 , n7806 );
    and g13455 ( n5783 , n333 , n10583 );
    and g13456 ( n13416 , n1962 , n5389 );
    or g13457 ( n7196 , n7076 , n5419 );
    or g13458 ( n5379 , n14435 , n3311 );
    or g13459 ( n5898 , n12211 , n2792 );
    and g13460 ( n2735 , n13863 , n87 );
    or g13461 ( n2216 , n7812 , n13162 );
    and g13462 ( n14432 , n678 , n1217 );
    or g13463 ( n5567 , n7530 , n12699 );
    or g13464 ( n2200 , n3168 , n1453 );
    and g13465 ( n9581 , n79 , n1119 );
    or g13466 ( n7790 , n584 , n527 );
    and g13467 ( n12135 , n1526 , n1556 );
    not g13468 ( n14400 , n12444 );
    or g13469 ( n13925 , n10062 , n13815 );
    and g13470 ( n14142 , n2486 , n10333 );
    or g13471 ( n9764 , n648 , n4579 );
    or g13472 ( n8339 , n7250 , n9735 );
    and g13473 ( n3292 , n12683 , n1496 );
    and g13474 ( n2891 , n12147 , n11341 );
    and g13475 ( n8646 , n1428 , n7933 );
    nor g13476 ( n705 , n8378 , n4773 );
    and g13477 ( n8707 , n8923 , n13523 );
    or g13478 ( n10866 , n13531 , n13848 );
    or g13479 ( n5135 , n14400 , n12624 );
    or g13480 ( n779 , n13501 , n6835 );
    or g13481 ( n7774 , n782 , n4418 );
    or g13482 ( n5506 , n747 , n1564 );
    and g13483 ( n14272 , n3169 , n7949 );
    not g13484 ( n8451 , n5300 );
    and g13485 ( n4606 , n10282 , n7065 );
    nor g13486 ( n10663 , n11998 , n8548 );
    and g13487 ( n6728 , n8111 , n2264 );
    and g13488 ( n7514 , n457 , n6293 );
    and g13489 ( n5037 , n3247 , n9877 );
    or g13490 ( n2900 , n12211 , n2741 );
    or g13491 ( n10123 , n4544 , n5892 );
    and g13492 ( n12813 , n13520 , n5330 );
    nor g13493 ( n6875 , n7683 , n5720 );
    or g13494 ( n13426 , n7523 , n10573 );
    and g13495 ( n10212 , n9113 , n5777 );
    and g13496 ( n8583 , n4445 , n1209 );
    and g13497 ( n2130 , n1073 , n6806 );
    not g13498 ( n1693 , n2577 );
    or g13499 ( n6958 , n4877 , n9192 );
    not g13500 ( n432 , n7275 );
    not g13501 ( n13246 , n1784 );
    nor g13502 ( n9284 , n10323 , n8441 );
    and g13503 ( n11160 , n8358 , n6637 );
    not g13504 ( n4443 , n9977 );
    and g13505 ( n4159 , n4856 , n441 );
    and g13506 ( n8414 , n12460 , n9859 );
    or g13507 ( n921 , n10234 , n13574 );
    or g13508 ( n14283 , n7798 , n4659 );
    or g13509 ( n6912 , n10309 , n13956 );
    not g13510 ( n2486 , n6975 );
    or g13511 ( n6662 , n5491 , n4126 );
    and g13512 ( n9580 , n6096 , n2910 );
    and g13513 ( n9255 , n8147 , n3018 );
    and g13514 ( n14098 , n1962 , n9360 );
    or g13515 ( n10836 , n8980 , n2204 );
    and g13516 ( n4436 , n12159 , n3622 );
    and g13517 ( n3896 , n7693 , n733 );
    not g13518 ( n5493 , n7819 );
    and g13519 ( n14023 , n4650 , n1260 );
    nor g13520 ( n14434 , n13365 , n7601 );
    or g13521 ( n6292 , n4255 , n8079 );
    and g13522 ( n9128 , n1254 , n6872 );
    or g13523 ( n13217 , n1147 , n14175 );
    or g13524 ( n366 , n11121 , n12719 );
    not g13525 ( n12389 , n13723 );
    or g13526 ( n7975 , n4065 , n2720 );
    not g13527 ( n3602 , n6159 );
    and g13528 ( n8484 , n1047 , n754 );
    and g13529 ( n7825 , n11404 , n10317 );
    and g13530 ( n1345 , n7909 , n6632 );
    or g13531 ( n2653 , n12211 , n4815 );
    or g13532 ( n1134 , n5234 , n9171 );
    and g13533 ( n4412 , n7911 , n2759 );
    or g13534 ( n7357 , n6350 , n1376 );
    and g13535 ( n11012 , n14109 , n2513 );
    or g13536 ( n8437 , n5472 , n6777 );
    or g13537 ( n13032 , n8210 , n9835 );
    nor g13538 ( n6997 , n13477 , n9768 );
    or g13539 ( n11528 , n6109 , n1620 );
    not g13540 ( n5001 , n12483 );
    and g13541 ( n11858 , n4627 , n12029 );
    and g13542 ( n12216 , n4486 , n10745 );
    and g13543 ( n8402 , n4098 , n698 );
    or g13544 ( n4306 , n8582 , n45 );
    not g13545 ( n4296 , n9537 );
    nor g13546 ( n8603 , n2087 , n8586 );
    and g13547 ( n5545 , n12918 , n3100 );
    not g13548 ( n480 , n2794 );
    or g13549 ( n13386 , n4162 , n11207 );
    and g13550 ( n9460 , n8047 , n12078 );
    or g13551 ( n11554 , n8986 , n13683 );
    or g13552 ( n3319 , n13276 , n12318 );
    and g13553 ( n9181 , n10374 , n8749 );
    not g13554 ( n12633 , n2130 );
    not g13555 ( n8238 , n7507 );
    and g13556 ( n7969 , n5999 , n11564 );
    not g13557 ( n8575 , n751 );
    or g13558 ( n10044 , n12625 , n13730 );
    or g13559 ( n8757 , n4205 , n3201 );
    or g13560 ( n12947 , n3366 , n11842 );
    nor g13561 ( n6702 , n10973 , n11449 );
    and g13562 ( n5000 , n5899 , n6716 );
    or g13563 ( n10887 , n3800 , n7532 );
    or g13564 ( n8266 , n7888 , n4037 );
    and g13565 ( n10661 , n12404 , n9928 );
    nor g13566 ( n2062 , n10285 , n13273 );
    or g13567 ( n1734 , n10154 , n6746 );
    not g13568 ( n9864 , n9371 );
    and g13569 ( n12641 , n4657 , n11281 );
    not g13570 ( n6260 , n7667 );
    and g13571 ( n7782 , n2942 , n8699 );
    or g13572 ( n6442 , n8726 , n11947 );
    or g13573 ( n6017 , n6373 , n5047 );
    not g13574 ( n2518 , n751 );
    or g13575 ( n9134 , n5904 , n9461 );
    or g13576 ( n14451 , n13080 , n11400 );
    and g13577 ( n9096 , n6680 , n3541 );
    nor g13578 ( n14028 , n9035 , n1393 );
    and g13579 ( n2693 , n6243 , n6102 );
    and g13580 ( n3540 , n889 , n778 );
    or g13581 ( n11014 , n8034 , n6060 );
    or g13582 ( n3847 , n1728 , n11352 );
    and g13583 ( n3431 , n10330 , n13428 );
    and g13584 ( n3588 , n10374 , n593 );
    not g13585 ( n10024 , n13668 );
    or g13586 ( n13348 , n4739 , n2940 );
    or g13587 ( n6493 , n3826 , n11421 );
    or g13588 ( n12717 , n13885 , n13164 );
    or g13589 ( n7651 , n9289 , n4691 );
    nor g13590 ( n8578 , n900 , n13163 );
    and g13591 ( n9145 , n5475 , n807 );
    nor g13592 ( n9694 , n10280 , n5945 );
    or g13593 ( n2411 , n3062 , n9531 );
    and g13594 ( n6671 , n8569 , n9471 );
    and g13595 ( n11314 , n14213 , n12991 );
    not g13596 ( n6051 , n2644 );
    not g13597 ( n9230 , n2472 );
    or g13598 ( n9692 , n6111 , n1540 );
    or g13599 ( n2207 , n4255 , n10728 );
    and g13600 ( n2763 , n7677 , n2197 );
    and g13601 ( n11646 , n4627 , n5070 );
    and g13602 ( n6664 , n2547 , n12603 );
    not g13603 ( n6167 , n1436 );
    and g13604 ( n12511 , n8697 , n14334 );
    and g13605 ( n12609 , n10647 , n13726 );
    not g13606 ( n12625 , n12687 );
    not g13607 ( n3401 , n9994 );
    nor g13608 ( n2764 , n2651 , n12860 );
    not g13609 ( n8881 , n14412 );
    or g13610 ( n12061 , n13108 , n12679 );
    and g13611 ( n10164 , n12741 , n5812 );
    or g13612 ( n2789 , n49 , n3680 );
    and g13613 ( n1993 , n9509 , n13239 );
    or g13614 ( n691 , n10396 , n2891 );
    nor g13615 ( n11695 , n3521 , n18 );
    not g13616 ( n5271 , n3583 );
    and g13617 ( n6378 , n3435 , n11612 );
    or g13618 ( n8373 , n283 , n10413 );
    not g13619 ( n7551 , n1833 );
    not g13620 ( n10083 , n9878 );
    not g13621 ( n10712 , n7402 );
    nor g13622 ( n13669 , n11558 , n8417 );
    and g13623 ( n11575 , n11008 , n13036 );
    not g13624 ( n3435 , n6990 );
    and g13625 ( n6038 , n10763 , n5298 );
    and g13626 ( n10967 , n2758 , n657 );
    and g13627 ( n12504 , n1678 , n669 );
    and g13628 ( n7152 , n9830 , n13278 );
    or g13629 ( n8184 , n930 , n10987 );
    or g13630 ( n3474 , n5084 , n12255 );
    nor g13631 ( n13235 , n7238 , n2544 );
    or g13632 ( n13770 , n9507 , n11357 );
    and g13633 ( n11826 , n286 , n4388 );
    and g13634 ( n7990 , n2422 , n7792 );
    and g13635 ( n8945 , n8569 , n3505 );
    or g13636 ( n3008 , n7041 , n12976 );
    and g13637 ( n5729 , n7779 , n9144 );
    and g13638 ( n7233 , n9080 , n1747 );
    not g13639 ( n10025 , n4755 );
    or g13640 ( n9899 , n10224 , n7126 );
    and g13641 ( n644 , n4354 , n14251 );
    not g13642 ( n12741 , n7278 );
    not g13643 ( n2378 , n12084 );
    and g13644 ( n1827 , n394 , n6184 );
    and g13645 ( n5241 , n11093 , n8019 );
    and g13646 ( n753 , n986 , n13418 );
    and g13647 ( n10085 , n1266 , n7636 );
    or g13648 ( n2708 , n12100 , n12299 );
    not g13649 ( n2002 , n9154 );
    or g13650 ( n4073 , n11123 , n7795 );
    and g13651 ( n12487 , n2082 , n12659 );
    or g13652 ( n4861 , n4602 , n6631 );
    and g13653 ( n4977 , n13297 , n3668 );
    nor g13654 ( n7801 , n4742 , n2617 );
    not g13655 ( n12040 , n9156 );
    or g13656 ( n2049 , n8034 , n4918 );
    or g13657 ( n9669 , n5647 , n7503 );
    not g13658 ( n2577 , n2889 );
    not g13659 ( n3882 , n9604 );
    and g13660 ( n8485 , n457 , n12703 );
    nor g13661 ( n13958 , n13276 , n11482 );
    not g13662 ( n7076 , n9453 );
    and g13663 ( n397 , n432 , n12225 );
    and g13664 ( n10260 , n5857 , n12305 );
    and g13665 ( n13488 , n1876 , n10732 );
    and g13666 ( n8345 , n14273 , n7216 );
    or g13667 ( n9702 , n4807 , n9709 );
    or g13668 ( n8105 , n695 , n5130 );
    and g13669 ( n6366 , n9571 , n1659 );
    not g13670 ( n648 , n12331 );
    or g13671 ( n4630 , n7462 , n10687 );
    nor g13672 ( n2424 , n2057 , n5883 );
    not g13673 ( n12460 , n6819 );
    nor g13674 ( n1672 , n1086 , n5958 );
    nor g13675 ( n8190 , n11580 , n11971 );
    nor g13676 ( n6488 , n7120 , n7161 );
    and g13677 ( n13571 , n13096 , n13645 );
    not g13678 ( n10960 , n81 );
    not g13679 ( n3512 , n2484 );
    and g13680 ( n9466 , n13096 , n6778 );
    and g13681 ( n6855 , n3762 , n6418 );
    and g13682 ( n8082 , n9953 , n9 );
    and g13683 ( n13614 , n11470 , n8869 );
    and g13684 ( n2247 , n8358 , n12061 );
    or g13685 ( n3553 , n1112 , n3308 );
    not g13686 ( n3088 , n13696 );
    and g13687 ( n238 , n7177 , n8496 );
    or g13688 ( n3257 , n12020 , n4896 );
    and g13689 ( n13562 , n13367 , n11118 );
    nor g13690 ( n13474 , n10936 , n9675 );
    nor g13691 ( n5741 , n9404 , n8840 );
    and g13692 ( n13375 , n9898 , n13733 );
    and g13693 ( n9387 , n7026 , n13412 );
    and g13694 ( n3712 , n13525 , n5207 );
    or g13695 ( n9593 , n2747 , n8381 );
    and g13696 ( n3878 , n11950 , n1632 );
    or g13697 ( n4987 , n1258 , n3564 );
    or g13698 ( n12842 , n11097 , n13200 );
    or g13699 ( n4009 , n5362 , n12256 );
    not g13700 ( n13404 , n5871 );
    and g13701 ( n4355 , n10330 , n4219 );
    and g13702 ( n2912 , n2724 , n10432 );
    and g13703 ( n2376 , n5434 , n2829 );
    and g13704 ( n5785 , n2310 , n6593 );
    not g13705 ( n2132 , n3989 );
    nor g13706 ( n297 , n11771 , n6475 );
    and g13707 ( n9478 , n10330 , n13735 );
    not g13708 ( n1705 , n12927 );
    not g13709 ( n8358 , n10177 );
    and g13710 ( n12287 , n3365 , n984 );
    or g13711 ( n4378 , n10808 , n6265 );
    and g13712 ( n13223 , n7211 , n6369 );
    or g13713 ( n6732 , n13276 , n7153 );
    or g13714 ( n4473 , n10871 , n12571 );
    not g13715 ( n871 , n9757 );
    nor g13716 ( n12162 , n2752 , n142 );
    or g13717 ( n9225 , n9285 , n5650 );
    and g13718 ( n13959 , n2334 , n8577 );
    or g13719 ( n11067 , n553 , n13772 );
    not g13720 ( n14332 , n5872 );
    and g13721 ( n13127 , n11748 , n3079 );
    or g13722 ( n11656 , n4033 , n9067 );
    and g13723 ( n879 , n7745 , n10350 );
    not g13724 ( n14313 , n1436 );
    nor g13725 ( n1033 , n12288 , n9927 );
    and g13726 ( n4149 , n7402 , n5129 );
    nor g13727 ( n9838 , n5480 , n11730 );
    not g13728 ( n8209 , n10108 );
    not g13729 ( n10189 , n8925 );
    and g13730 ( n7190 , n4554 , n4103 );
    or g13731 ( n7491 , n10019 , n11544 );
    and g13732 ( n9472 , n11213 , n5700 );
    not g13733 ( n3743 , n11425 );
    or g13734 ( n2419 , n5603 , n10299 );
    and g13735 ( n5503 , n327 , n10094 );
    or g13736 ( n4153 , n13226 , n11583 );
    and g13737 ( n1966 , n12121 , n11606 );
    or g13738 ( n10324 , n2949 , n1451 );
    and g13739 ( n4835 , n8866 , n9372 );
    nor g13740 ( n10878 , n7229 , n11041 );
    and g13741 ( n7299 , n1071 , n13764 );
    and g13742 ( n11995 , n11495 , n13915 );
    nor g13743 ( n7136 , n13154 , n8104 );
    and g13744 ( n2927 , n11316 , n375 );
    and g13745 ( n7363 , n10820 , n2984 );
    or g13746 ( n11936 , n12695 , n5401 );
    or g13747 ( n2262 , n10025 , n4172 );
    nor g13748 ( n3467 , n6907 , n7432 );
    and g13749 ( n8382 , n2643 , n4242 );
    and g13750 ( n9499 , n4901 , n4714 );
    and g13751 ( n6564 , n7970 , n4421 );
    and g13752 ( n4321 , n536 , n8766 );
    or g13753 ( n12647 , n12292 , n6650 );
    or g13754 ( n11168 , n10784 , n9018 );
    or g13755 ( n11698 , n13516 , n9233 );
    or g13756 ( n9034 , n2949 , n215 );
    or g13757 ( n2105 , n6695 , n11820 );
    not g13758 ( n588 , n10384 );
    or g13759 ( n9815 , n4684 , n7569 );
    not g13760 ( n8540 , n11633 );
    and g13761 ( n1606 , n98 , n11661 );
    and g13762 ( n11161 , n13433 , n345 );
    and g13763 ( n7918 , n2758 , n3705 );
    not g13764 ( n1771 , n11375 );
    and g13765 ( n3209 , n4347 , n1836 );
    and g13766 ( n11025 , n9323 , n10770 );
    nor g13767 ( n1341 , n1844 , n13011 );
    and g13768 ( n8503 , n8043 , n4499 );
    not g13769 ( n8147 , n5182 );
    nor g13770 ( n10980 , n5435 , n13616 );
    and g13771 ( n5579 , n432 , n8118 );
    nor g13772 ( n3721 , n2154 , n1858 );
    nor g13773 ( n8688 , n8363 , n13975 );
    or g13774 ( n1371 , n4967 , n5763 );
    or g13775 ( n3065 , n4898 , n2018 );
    and g13776 ( n3738 , n10556 , n9220 );
    not g13777 ( n5891 , n7600 );
    or g13778 ( n11276 , n10560 , n4322 );
    and g13779 ( n1731 , n10562 , n1433 );
    not g13780 ( n2343 , n12244 );
    and g13781 ( n552 , n5459 , n12340 );
    and g13782 ( n8321 , n1071 , n12022 );
    nor g13783 ( n13013 , n4207 , n5164 );
    or g13784 ( n12242 , n12139 , n5646 );
    nor g13785 ( n2345 , n13458 , n5518 );
    and g13786 ( n5221 , n2080 , n11392 );
    not g13787 ( n3286 , n7346 );
    not g13788 ( n6354 , n3361 );
    or g13789 ( n3109 , n412 , n6668 );
    or g13790 ( n1977 , n12759 , n4177 );
    and g13791 ( n3988 , n8605 , n4019 );
    or g13792 ( n10634 , n4128 , n7112 );
    or g13793 ( n14292 , n5266 , n8854 );
    and g13794 ( n11596 , n7670 , n12546 );
    and g13795 ( n9465 , n13132 , n3364 );
    nor g13796 ( n14222 , n6747 , n8787 );
    not g13797 ( n1711 , n382 );
    and g13798 ( n9579 , n4346 , n7193 );
    and g13799 ( n2871 , n11384 , n13033 );
    nor g13800 ( n6932 , n1218 , n9439 );
    or g13801 ( n10504 , n838 , n1132 );
    and g13802 ( n11408 , n2643 , n2358 );
    or g13803 ( n10415 , n1383 , n6709 );
    or g13804 ( n12686 , n5253 , n7937 );
    or g13805 ( n10034 , n9747 , n1070 );
    not g13806 ( n6888 , n2607 );
    and g13807 ( n916 , n865 , n6821 );
    nor g13808 ( n2302 , n5665 , n5932 );
    and g13809 ( n3070 , n8521 , n3977 );
    not g13810 ( n13745 , n13038 );
    or g13811 ( n6610 , n2562 , n11338 );
    and g13812 ( n13800 , n12101 , n5969 );
    not g13813 ( n749 , n3922 );
    and g13814 ( n11800 , n10367 , n3552 );
    not g13815 ( n4581 , n4490 );
    and g13816 ( n12065 , n5088 , n12816 );
    or g13817 ( n6233 , n2401 , n11962 );
    or g13818 ( n10666 , n4508 , n9719 );
    and g13819 ( n12775 , n13952 , n590 );
    and g13820 ( n6650 , n1772 , n5719 );
    not g13821 ( n13537 , n12106 );
    or g13822 ( n8669 , n10396 , n13748 );
    not g13823 ( n9863 , n13190 );
    and g13824 ( n8715 , n11607 , n7477 );
    and g13825 ( n12815 , n2533 , n9335 );
    or g13826 ( n452 , n4791 , n10190 );
    or g13827 ( n2840 , n2645 , n9337 );
    and g13828 ( n4853 , n2021 , n169 );
    not g13829 ( n10763 , n261 );
    not g13830 ( n2607 , n3443 );
    not g13831 ( n12088 , n7146 );
    and g13832 ( n9030 , n6318 , n6093 );
    not g13833 ( n6428 , n3021 );
    or g13834 ( n12893 , n480 , n6699 );
    nor g13835 ( n12923 , n9563 , n4101 );
    not g13836 ( n5132 , n4317 );
    and g13837 ( n7251 , n1804 , n9132 );
    not g13838 ( n12250 , n3967 );
    or g13839 ( n4182 , n3768 , n4761 );
    and g13840 ( n4568 , n1854 , n13825 );
    not g13841 ( n5833 , n1676 );
    and g13842 ( n13419 , n11737 , n9183 );
    nor g13843 ( n13984 , n12757 , n13159 );
    and g13844 ( n7000 , n2533 , n3507 );
    not g13845 ( n12521 , n6193 );
    nor g13846 ( n13378 , n6788 , n10856 );
    or g13847 ( n12763 , n13516 , n11888 );
    and g13848 ( n13405 , n2521 , n12837 );
    nor g13849 ( n1392 , n5018 , n3568 );
    and g13850 ( n8677 , n2158 , n9159 );
    or g13851 ( n9249 , n4822 , n9042 );
    and g13852 ( n7953 , n2998 , n6340 );
    nor g13853 ( n10959 , n7229 , n2952 );
    or g13854 ( n10026 , n3076 , n2159 );
    or g13855 ( n11137 , n2387 , n12183 );
    nor g13856 ( n11434 , n1522 , n11531 );
    and g13857 ( n8205 , n7063 , n9855 );
    nor g13858 ( n1103 , n13399 , n164 );
    or g13859 ( n973 , n8747 , n13660 );
    nor g13860 ( n3951 , n14216 , n5112 );
    or g13861 ( n5359 , n1152 , n1299 );
    or g13862 ( n729 , n9931 , n2222 );
    or g13863 ( n10863 , n7219 , n7162 );
    and g13864 ( n4317 , n11130 , n2548 );
    and g13865 ( n6985 , n7909 , n4406 );
    and g13866 ( n253 , n1962 , n13022 );
    and g13867 ( n6864 , n1678 , n10735 );
    not g13868 ( n4807 , n2918 );
    or g13869 ( n7644 , n5574 , n6703 );
    or g13870 ( n2535 , n555 , n4545 );
    or g13871 ( n12971 , n6206 , n8041 );
    not g13872 ( n8748 , n12331 );
    nor g13873 ( n4455 , n450 , n14311 );
    and g13874 ( n3633 , n8965 , n620 );
    not g13875 ( n8217 , n2973 );
    not g13876 ( n4490 , n9987 );
    not g13877 ( n1844 , n7404 );
    or g13878 ( n9210 , n11558 , n10527 );
    and g13879 ( n4731 , n1100 , n13284 );
    and g13880 ( n1550 , n5275 , n171 );
    nor g13881 ( n159 , n3867 , n2717 );
    and g13882 ( n14081 , n7911 , n12737 );
    and g13883 ( n2425 , n8849 , n7820 );
    nor g13884 ( n4636 , n11870 , n6529 );
    nor g13885 ( n10391 , n6211 , n117 );
    not g13886 ( n14133 , n1079 );
    or g13887 ( n4733 , n8480 , n9680 );
    or g13888 ( n2178 , n11223 , n10818 );
    and g13889 ( n268 , n12147 , n8267 );
    and g13890 ( n14057 , n13728 , n929 );
    and g13891 ( n5143 , n11702 , n12709 );
    and g13892 ( n10872 , n1788 , n10999 );
    or g13893 ( n12364 , n11724 , n4986 );
    or g13894 ( n4008 , n7436 , n14212 );
    or g13895 ( n10659 , n10331 , n1633 );
    not g13896 ( n10367 , n82 );
    and g13897 ( n4643 , n2985 , n6641 );
    or g13898 ( n8270 , n5180 , n5173 );
    or g13899 ( n13329 , n6781 , n12993 );
    and g13900 ( n2936 , n333 , n5318 );
    not g13901 ( n7278 , n2723 );
    nor g13902 ( n11862 , n194 , n10271 );
    and g13903 ( n11335 , n4973 , n8792 );
    or g13904 ( n2630 , n10626 , n5853 );
    or g13905 ( n13293 , n6596 , n354 );
    and g13906 ( n13048 , n1857 , n13631 );
    and g13907 ( n4138 , n7767 , n7125 );
    and g13908 ( n13271 , n392 , n10439 );
    and g13909 ( n5095 , n12092 , n13185 );
    and g13910 ( n9515 , n4358 , n1934 );
    and g13911 ( n8215 , n10407 , n10128 );
    not g13912 ( n13342 , n13383 );
    and g13913 ( n11401 , n14376 , n9616 );
    or g13914 ( n12368 , n8513 , n13684 );
    and g13915 ( n8627 , n12858 , n1892 );
    or g13916 ( n764 , n4128 , n12264 );
    and g13917 ( n6146 , n3952 , n5413 );
    or g13918 ( n9759 , n3161 , n3092 );
    or g13919 ( n6163 , n6266 , n13429 );
    or g13920 ( n1695 , n85 , n6859 );
    and g13921 ( n12320 , n8453 , n7139 );
    and g13922 ( n90 , n1678 , n4482 );
    and g13923 ( n14426 , n4546 , n12207 );
    and g13924 ( n5654 , n9673 , n9274 );
    nor g13925 ( n12978 , n8816 , n413 );
    not g13926 ( n13128 , n421 );
    not g13927 ( n8412 , n1639 );
    or g13928 ( n10208 , n1602 , n12252 );
    or g13929 ( n10348 , n4255 , n5206 );
    or g13930 ( n4234 , n10933 , n5563 );
    nor g13931 ( n8733 , n2597 , n7841 );
    and g13932 ( n6696 , n6517 , n2054 );
    nor g13933 ( n2234 , n4928 , n4368 );
    nor g13934 ( n3686 , n14367 , n4653 );
    or g13935 ( n7410 , n185 , n5193 );
    and g13936 ( n6381 , n5137 , n9160 );
    and g13937 ( n13029 , n13297 , n14268 );
    or g13938 ( n11568 , n12870 , n14215 );
    and g13939 ( n11619 , n1699 , n11518 );
    and g13940 ( n5623 , n3424 , n10173 );
    and g13941 ( n8395 , n5038 , n10275 );
    or g13942 ( n4304 , n11980 , n2979 );
    nor g13943 ( n10548 , n10136 , n9126 );
    and g13944 ( n14354 , n13633 , n3523 );
    and g13945 ( n4027 , n231 , n7196 );
    nor g13946 ( n3014 , n2341 , n9284 );
    or g13947 ( n5576 , n9494 , n5467 );
    or g13948 ( n14040 , n5587 , n10416 );
    not g13949 ( n6898 , n2468 );
    not g13950 ( n1577 , n5306 );
    not g13951 ( n9529 , n1041 );
    and g13952 ( n4037 , n8432 , n5175 );
    and g13953 ( n2823 , n10367 , n2076 );
    and g13954 ( n8228 , n6957 , n13469 );
    and g13955 ( n5080 , n3846 , n10585 );
    or g13956 ( n12436 , n9716 , n1814 );
    not g13957 ( n815 , n3972 );
    and g13958 ( n1649 , n4354 , n2168 );
    or g13959 ( n2406 , n10294 , n7552 );
    or g13960 ( n1925 , n3800 , n9905 );
    not g13961 ( n8122 , n2250 );
    not g13962 ( n7068 , n3926 );
    and g13963 ( n96 , n6830 , n12910 );
    not g13964 ( n11425 , n13135 );
    and g13965 ( n6083 , n1427 , n6406 );
    and g13966 ( n13544 , n7708 , n10326 );
    not g13967 ( n560 , n5786 );
    or g13968 ( n3056 , n11951 , n6019 );
    and g13969 ( n4236 , n10710 , n13218 );
    and g13970 ( n1133 , n3212 , n13536 );
    not g13971 ( n10186 , n3461 );
    not g13972 ( n8965 , n10303 );
    not g13973 ( n10534 , n7441 );
    and g13974 ( n3479 , n638 , n5349 );
    and g13975 ( n3306 , n13781 , n7412 );
    and g13976 ( n7600 , n4258 , n5702 );
    or g13977 ( n1322 , n10323 , n4521 );
    and g13978 ( n1650 , n3424 , n10054 );
    or g13979 ( n6984 , n3492 , n13882 );
    or g13980 ( n13923 , n5406 , n8033 );
    and g13981 ( n3987 , n4851 , n12869 );
    or g13982 ( n4349 , n6519 , n5801 );
    or g13983 ( n7998 , n5891 , n6392 );
    and g13984 ( n11471 , n898 , n1778 );
    and g13985 ( n4918 , n10622 , n6155 );
    or g13986 ( n9480 , n4052 , n7000 );
    or g13987 ( n12819 , n5908 , n14024 );
    and g13988 ( n3831 , n3370 , n10304 );
    nor g13989 ( n7161 , n11980 , n12838 );
    or g13990 ( n13998 , n10396 , n268 );
    not g13991 ( n7673 , n10269 );
    or g13992 ( n3129 , n4908 , n11665 );
    not g13993 ( n11305 , n8003 );
    not g13994 ( n13728 , n14475 );
    and g13995 ( n10223 , n5459 , n3264 );
    and g13996 ( n5206 , n3986 , n2109 );
    and g13997 ( n1305 , n11300 , n5757 );
    nor g13998 ( n4059 , n10637 , n3040 );
    nor g13999 ( n4063 , n13255 , n4218 );
    not g14000 ( n1120 , n9608 );
    or g14001 ( n3824 , n13698 , n6557 );
    or g14002 ( n5207 , n8476 , n10144 );
    or g14003 ( n8912 , n4631 , n5520 );
    or g14004 ( n4863 , n3047 , n14276 );
    nor g14005 ( n6405 , n7364 , n532 );
    or g14006 ( n5217 , n12614 , n10765 );
    not g14007 ( n5640 , n411 );
    and g14008 ( n6627 , n3755 , n10178 );
    or g14009 ( n13088 , n5139 , n10766 );
    not g14010 ( n5108 , n179 );
    not g14011 ( n10303 , n9537 );
    and g14012 ( n7508 , n873 , n1035 );
    or g14013 ( n8593 , n782 , n4585 );
    not g14014 ( n5315 , n3021 );
    nor g14015 ( n9672 , n12193 , n12273 );
    or g14016 ( n5697 , n14319 , n4954 );
    and g14017 ( n4833 , n3724 , n9750 );
    and g14018 ( n6846 , n5434 , n14005 );
    nor g14019 ( n1226 , n14135 , n5914 );
    not g14020 ( n7911 , n8524 );
    and g14021 ( n3437 , n14313 , n8438 );
    or g14022 ( n12995 , n12852 , n3263 );
    or g14023 ( n2526 , n1535 , n13326 );
    and g14024 ( n6674 , n5137 , n11784 );
    and g14025 ( n3123 , n5240 , n1444 );
    or g14026 ( n4993 , n5454 , n2658 );
    nor g14027 ( n9704 , n13276 , n7804 );
    not g14028 ( n9806 , n10346 );
    nor g14029 ( n10235 , n7971 , n2899 );
    and g14030 ( n4305 , n2454 , n12194 );
    and g14031 ( n11494 , n9265 , n3590 );
    not g14032 ( n8932 , n2241 );
    not g14033 ( n10535 , n6096 );
    or g14034 ( n10021 , n13446 , n3483 );
    and g14035 ( n14032 , n8789 , n5158 );
    and g14036 ( n13841 , n1539 , n7556 );
    or g14037 ( n7646 , n1535 , n8922 );
    or g14038 ( n837 , n2315 , n10270 );
    not g14039 ( n14419 , n3070 );
    or g14040 ( n7668 , n4684 , n7415 );
    not g14041 ( n5012 , n2432 );
    or g14042 ( n5911 , n1223 , n932 );
    and g14043 ( n14456 , n13069 , n14194 );
    and g14044 ( n10176 , n8453 , n837 );
    not g14045 ( n12105 , n2906 );
    or g14046 ( n6462 , n6373 , n1880 );
    or g14047 ( n1757 , n1840 , n12589 );
    and g14048 ( n4400 , n4509 , n12728 );
    and g14049 ( n8123 , n2445 , n2890 );
    and g14050 ( n6203 , n7208 , n3454 );
    not g14051 ( n7401 , n844 );
    or g14052 ( n14068 , n9353 , n14153 );
    nor g14053 ( n9496 , n6679 , n7444 );
    not g14054 ( n14088 , n12874 );
    and g14055 ( n12921 , n286 , n9125 );
    or g14056 ( n13330 , n13885 , n10033 );
    and g14057 ( n2152 , n428 , n8938 );
    nor g14058 ( n5945 , n8209 , n7377 );
    not g14059 ( n4757 , n11325 );
    not g14060 ( n12013 , n6807 );
    nor g14061 ( n11486 , n4144 , n10625 );
    or g14062 ( n2001 , n12037 , n3367 );
    not g14063 ( n6600 , n1776 );
    or g14064 ( n10545 , n8480 , n6647 );
    or g14065 ( n4085 , n2401 , n11306 );
    not g14066 ( n9442 , n6274 );
    or g14067 ( n13889 , n5548 , n13222 );
    or g14068 ( n9623 , n3445 , n11382 );
    or g14069 ( n6160 , n3559 , n12917 );
    not g14070 ( n2547 , n4633 );
    nor g14071 ( n117 , n8527 , n3686 );
    or g14072 ( n2268 , n14282 , n1649 );
    or g14073 ( n3429 , n9747 , n13314 );
    or g14074 ( n13188 , n11724 , n1197 );
    or g14075 ( n4886 , n900 , n11443 );
    nor g14076 ( n8691 , n8212 , n3032 );
    and g14077 ( n2792 , n7068 , n9200 );
    and g14078 ( n14314 , n11008 , n14201 );
    or g14079 ( n6144 , n10760 , n7354 );
    and g14080 ( n1113 , n3401 , n12486 );
    not g14081 ( n13675 , n9306 );
    and g14082 ( n8619 , n4627 , n9344 );
    and g14083 ( n9173 , n12531 , n13787 );
    or g14084 ( n899 , n695 , n1906 );
    not g14085 ( n1436 , n10485 );
    not g14086 ( n965 , n6990 );
    or g14087 ( n11372 , n9422 , n12881 );
    nor g14088 ( n4118 , n11148 , n11662 );
    or g14089 ( n4302 , n5732 , n14151 );
    nor g14090 ( n4348 , n10651 , n13259 );
    or g14091 ( n14113 , n4205 , n7012 );
    nor g14092 ( n14183 , n14166 , n341 );
    or g14093 ( n8530 , n5569 , n1340 );
    or g14094 ( n9874 , n4877 , n821 );
    or g14095 ( n1975 , n9429 , n11523 );
    or g14096 ( n2292 , n14110 , n11575 );
    and g14097 ( n9749 , n5011 , n11932 );
    and g14098 ( n10681 , n6318 , n11568 );
    nor g14099 ( n13053 , n10637 , n12743 );
    or g14100 ( n8396 , n13948 , n5583 );
    and g14101 ( n4868 , n8412 , n1757 );
    or g14102 ( n9992 , n8490 , n10410 );
    not g14103 ( n5690 , n14216 );
    or g14104 ( n3615 , n4508 , n11833 );
    nor g14105 ( n3973 , n2017 , n13389 );
    and g14106 ( n2658 , n13379 , n4250 );
    and g14107 ( n1182 , n14313 , n841 );
    not g14108 ( n1997 , n1458 );
    and g14109 ( n8117 , n2330 , n10045 );
    or g14110 ( n12186 , n11048 , n4414 );
    not g14111 ( n1617 , n264 );
    or g14112 ( n14442 , n10461 , n4397 );
    or g14113 ( n6067 , n957 , n9555 );
    nor g14114 ( n1126 , n12069 , n8876 );
    or g14115 ( n1725 , n2315 , n4586 );
    and g14116 ( n4369 , n889 , n10077 );
    and g14117 ( n9324 , n13755 , n9122 );
    and g14118 ( n6364 , n4650 , n4385 );
    and g14119 ( n4165 , n11636 , n5013 );
    or g14120 ( n6815 , n13226 , n9684 );
    and g14121 ( n13242 , n11679 , n6675 );
    or g14122 ( n125 , n2401 , n13629 );
    and g14123 ( n13694 , n2021 , n5564 );
    and g14124 ( n823 , n14038 , n13590 );
    nor g14125 ( n8121 , n12651 , n1174 );
    nor g14126 ( n10447 , n5197 , n3475 );
    not g14127 ( n9726 , n10372 );
    and g14128 ( n7751 , n10922 , n14403 );
    not g14129 ( n9811 , n6819 );
    or g14130 ( n1119 , n13080 , n14478 );
    or g14131 ( n4173 , n7678 , n13868 );
    and g14132 ( n3921 , n9564 , n8422 );
    or g14133 ( n1343 , n7430 , n1083 );
    not g14134 ( n11350 , n5665 );
    or g14135 ( n7297 , n8877 , n5102 );
    or g14136 ( n2661 , n4822 , n4334 );
    not g14137 ( n7590 , n10615 );
    and g14138 ( n9640 , n7401 , n3820 );
    or g14139 ( n1679 , n5575 , n2116 );
    or g14140 ( n3415 , n12821 , n2095 );
    not g14141 ( n4394 , n8963 );
    or g14142 ( n2849 , n11572 , n3377 );
    or g14143 ( n11133 , n1697 , n12751 );
    and g14144 ( n13906 , n12918 , n1933 );
    or g14145 ( n10741 , n2857 , n13269 );
    or g14146 ( n7737 , n163 , n11945 );
    and g14147 ( n14306 , n7427 , n9032 );
    not g14148 ( n13112 , n9453 );
    and g14149 ( n13849 , n2099 , n9304 );
    and g14150 ( n245 , n2310 , n9836 );
    and g14151 ( n3547 , n4880 , n11608 );
    and g14152 ( n12298 , n8507 , n8847 );
    not g14153 ( n10857 , n12874 );
    and g14154 ( n459 , n5640 , n1656 );
    or g14155 ( n6757 , n8726 , n1190 );
    or g14156 ( n1034 , n2246 , n1505 );
    nor g14157 ( n9137 , n10233 , n6634 );
    and g14158 ( n6542 , n12615 , n13721 );
    nor g14159 ( n8051 , n5847 , n5791 );
    and g14160 ( n2022 , n3526 , n7562 );
    or g14161 ( n5373 , n1669 , n13608 );
    not g14162 ( n1788 , n6975 );
    or g14163 ( n1990 , n6046 , n7349 );
    and g14164 ( n1108 , n3491 , n4632 );
    not g14165 ( n3255 , n8704 );
    not g14166 ( n11111 , n1053 );
    or g14167 ( n12214 , n12712 , n7256 );
    and g14168 ( n14261 , n10969 , n2944 );
    or g14169 ( n3283 , n976 , n4919 );
    nor g14170 ( n6282 , n8544 , n1090 );
    and g14171 ( n14478 , n11867 , n2230 );
    not g14172 ( n13706 , n12687 );
    nor g14173 ( n5894 , n5596 , n9616 );
    or g14174 ( n8693 , n553 , n5524 );
    and g14175 ( n81 , n8179 , n3155 );
    or g14176 ( n12628 , n4313 , n2753 );
    or g14177 ( n1054 , n3762 , n8635 );
    and g14178 ( n5651 , n4790 , n229 );
    and g14179 ( n9342 , n8439 , n4164 );
    or g14180 ( n2591 , n7481 , n2706 );
    and g14181 ( n664 , n6013 , n3594 );
    and g14182 ( n14034 , n1125 , n549 );
    and g14183 ( n857 , n10310 , n4072 );
    and g14184 ( n4187 , n9188 , n11145 );
    or g14185 ( n3529 , n5491 , n10486 );
    and g14186 ( n2148 , n748 , n576 );
    or g14187 ( n9691 , n8045 , n14119 );
    and g14188 ( n9697 , n7693 , n7649 );
    not g14189 ( n5605 , n13633 );
    and g14190 ( n3509 , n3785 , n11979 );
    or g14191 ( n11140 , n3800 , n12604 );
    nor g14192 ( n8449 , n648 , n5216 );
    nor g14193 ( n2811 , n1612 , n1486 );
    or g14194 ( n11774 , n10825 , n4028 );
    nor g14195 ( n3940 , n506 , n6964 );
    and g14196 ( n9259 , n2422 , n8245 );
    or g14197 ( n9300 , n12414 , n5115 );
    and g14198 ( n8683 , n5857 , n6245 );
    not g14199 ( n7427 , n261 );
    or g14200 ( n10352 , n4052 , n2308 );
    and g14201 ( n2233 , n4018 , n10159 );
    or g14202 ( n11591 , n1494 , n10896 );
    and g14203 ( n4732 , n13489 , n10044 );
    and g14204 ( n2151 , n4973 , n6004 );
    and g14205 ( n5016 , n8183 , n4875 );
    and g14206 ( n167 , n4619 , n3625 );
    and g14207 ( n5648 , n13236 , n8916 );
    or g14208 ( n11339 , n11303 , n14111 );
    and g14209 ( n3773 , n3526 , n3538 );
    or g14210 ( n10496 , n13142 , n14235 );
    or g14211 ( n4488 , n9804 , n4885 );
    and g14212 ( n11896 , n14213 , n10698 );
    or g14213 ( n14097 , n13485 , n10160 );
    or g14214 ( n3425 , n6263 , n8966 );
    and g14215 ( n1056 , n12391 , n13970 );
    not g14216 ( n12445 , n5613 );
    nor g14217 ( n14052 , n8212 , n11101 );
    or g14218 ( n1542 , n8582 , n7711 );
    and g14219 ( n9870 , n6625 , n5426 );
    not g14220 ( n4967 , n10889 );
    or g14221 ( n3269 , n11231 , n10754 );
    not g14222 ( n12651 , n2970 );
    or g14223 ( n9682 , n9289 , n12929 );
    not g14224 ( n4574 , n920 );
    not g14225 ( n3867 , n4859 );
    and g14226 ( n12638 , n13078 , n4995 );
    and g14227 ( n12845 , n11737 , n2020 );
    and g14228 ( n1098 , n11569 , n2841 );
    and g14229 ( n10022 , n3635 , n615 );
    and g14230 ( n750 , n7391 , n8545 );
    not g14231 ( n808 , n8361 );
    or g14232 ( n6261 , n4988 , n4328 );
    or g14233 ( n12323 , n3367 , n11776 );
    or g14234 ( n14515 , n8151 , n12196 );
    nor g14235 ( n4002 , n11488 , n4747 );
    and g14236 ( n10958 , n4486 , n3606 );
    and g14237 ( n8089 , n13246 , n4269 );
    or g14238 ( n3049 , n1576 , n5651 );
    or g14239 ( n658 , n3125 , n9478 );
    and g14240 ( n1718 , n11674 , n9512 );
    and g14241 ( n5566 , n12038 , n9477 );
    and g14242 ( n12394 , n9769 , n4134 );
    or g14243 ( n13758 , n11097 , n373 );
    or g14244 ( n5923 , n11090 , n9099 );
    and g14245 ( n10243 , n7327 , n2339 );
    or g14246 ( n7703 , n69 , n11900 );
    or g14247 ( n1271 , n2318 , n1795 );
    and g14248 ( n4595 , n14065 , n3199 );
    or g14249 ( n9435 , n7736 , n8893 );
    nor g14250 ( n13975 , n3871 , n3458 );
    nor g14251 ( n9834 , n512 , n2757 );
    or g14252 ( n1076 , n9956 , n8397 );
    or g14253 ( n5670 , n11011 , n14369 );
    and g14254 ( n13316 , n5467 , n886 );
    or g14255 ( n12241 , n11581 , n3312 );
    and g14256 ( n940 , n10229 , n3110 );
    and g14257 ( n5850 , n3846 , n1284 );
    or g14258 ( n6435 , n7736 , n1745 );
    nor g14259 ( n10180 , n573 , n12024 );
    or g14260 ( n1882 , n2387 , n7715 );
    not g14261 ( n6319 , n6011 );
    and g14262 ( n1710 , n12389 , n13291 );
    and g14263 ( n12255 , n4581 , n5954 );
    or g14264 ( n2063 , n7912 , n951 );
    or g14265 ( n1429 , n5507 , n7305 );
    and g14266 ( n14036 , n6525 , n3982 );
    nor g14267 ( n9365 , n10309 , n9440 );
    not g14268 ( n536 , n1478 );
    or g14269 ( n5757 , n3168 , n4057 );
    and g14270 ( n3438 , n12057 , n10090 );
endmodule
