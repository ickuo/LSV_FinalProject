module top( n36 , n147 , n697 , n800 , n830 , n835 , n848 , n1178 , n1217 , 
n1275 , n1336 , n1715 , n1836 , n1842 , n1858 , n1950 , n2001 , n2104 , n2172 , 
n2366 , n2479 , n2764 , n3205 , n3222 , n3694 , n3741 , n3946 , n4288 , n4461 , 
n4519 , n4758 , n4772 , n4788 , n4878 , n4885 , n4960 , n4962 , n5067 , n5287 , 
n5335 , n5738 , n6226 , n6542 , n6875 , n7153 , n7540 , n7647 , n7759 , n7910 , 
n8431 , n8432 , n8594 , n9194 , n9291 , n9495 , n9568 , n9658 , n9789 , n9793 , 
n10297 , n10298 , n10682 , n10768 , n10852 , n10894 , n11046 , n11190 , n11218 , n11243 , 
n11455 , n11833 , n11961 , n12062 , n12183 , n12264 , n13159 , n13179 , n13217 , n13413 , 
n13455 , n13553 , n13967 , n14261 , n14263 , n14488 , n15095 , n15097 , n15131 , n15299 , 
n15357 , n15403 , n15464 , n15497 , n15570 , n15886 , n16135 , n16524 , n16620 , n16700 , 
n16817 , n16895 , n16899 , n16912 , n16922 , n16961 , n17485 , n17568 , n17702 , n17751 , 
n17829 , n17871 , n17982 , n18379 , n18477 , n18841 , n18912 , n18986 , n19084 , n19182 , 
n19418 , n19421 , n19454 , n19458 , n19484 , n19551 , n19984 , n20010 , n20210 , n20318 , 
n20358 , n20432 , n20466 , n20812 , n20979 , n21027 , n21281 , n21364 , n21426 , n21644 , 
n21673 , n21737 , n21996 , n22291 , n22322 , n22781 , n22980 , n23011 , n23222 , n23320 , 
n23426 , n23604 , n23953 , n24047 , n24259 , n24332 , n24356 , n24371 , n24434 , n25036 , 
n25174 , n25255 , n25355 , n25447 , n25602 , n25631 , n25694 , n25767 , n25831 , n26329 , 
n26336 , n26659 , n26695 , n26801 , n26984 , n27009 , n27226 , n27291 , n27447 , n27467 , 
n27489 , n27501 , n27627 , n27641 , n28093 , n28563 , n28667 , n28946 , n28958 , n28969 , 
n29037 , n29261 , n29649 , n29713 , n29731 , n29744 , n29788 , n29839 , n29884 , n30009 , 
n30016 , n30141 , n30181 , n30204 , n30292 , n30306 , n30507 , n30553 , n30578 , n30625 , 
n30646 , n30742 , n30986 , n31054 , n31056 , n31215 , n31272 , n31289 , n31419 , n31559 , 
n31606 , n31799 , n31803 , n32095 , n32205 , n32329 , n32584 , n32665 , n32675 , n32697 , 
n32715 , n32857 , n33004 , n33041 , n33116 , n33248 , n33524 , n33588 , n33650 , n33890 , 
n34201 , n34245 , n34269 , n34484 , n34571 , n34677 , n34820 , n34903 , n34923 , n35029 , 
n35111 , n35372 , n35479 , n35618 , n35924 , n35927 , n35950 );
    input n147 , n830 , n835 , n1178 , n1217 , n1836 , n1842 , n1950 , n2172 , 
n2764 , n3205 , n3222 , n3741 , n3946 , n4288 , n4461 , n4519 , n4758 , n4878 , 
n4960 , n4962 , n5067 , n5287 , n5335 , n5738 , n6226 , n7540 , n7759 , n8431 , 
n8432 , n9291 , n9568 , n9658 , n9789 , n9793 , n10298 , n10768 , n10852 , n10894 , 
n11046 , n11190 , n11455 , n12062 , n12264 , n13159 , n13179 , n13413 , n13553 , n15095 , 
n15097 , n15299 , n15403 , n15464 , n15886 , n16135 , n16620 , n16922 , n17485 , n17568 , 
n17702 , n17751 , n17982 , n18379 , n18912 , n19182 , n19418 , n19458 , n19551 , n19984 , 
n21281 , n21737 , n22291 , n22980 , n23604 , n23953 , n24332 , n24371 , n24434 , n25174 , 
n25602 , n25767 , n26695 , n26801 , n27009 , n27226 , n27291 , n27489 , n27627 , n28563 , 
n28958 , n29037 , n29649 , n29713 , n29731 , n29839 , n29884 , n30009 , n30016 , n30141 , 
n30181 , n30306 , n30553 , n30578 , n30742 , n31054 , n31056 , n31215 , n31272 , n31289 , 
n31419 , n31559 , n31799 , n32095 , n32584 , n32675 , n32715 , n32857 , n33041 , n33524 , 
n33588 , n33650 , n33890 , n34269 , n34677 , n35372 , n35479 , n35927 , n35950 ;
    output n36 , n697 , n800 , n848 , n1275 , n1336 , n1715 , n1858 , n2001 , 
n2104 , n2366 , n2479 , n3694 , n4772 , n4788 , n4885 , n6542 , n6875 , n7153 , 
n7647 , n7910 , n8594 , n9194 , n9495 , n10297 , n10682 , n11218 , n11243 , n11833 , 
n11961 , n12183 , n13217 , n13455 , n13967 , n14261 , n14263 , n14488 , n15131 , n15357 , 
n15497 , n15570 , n16524 , n16700 , n16817 , n16895 , n16899 , n16912 , n16961 , n17829 , 
n17871 , n18477 , n18841 , n18986 , n19084 , n19421 , n19454 , n19484 , n20010 , n20210 , 
n20318 , n20358 , n20432 , n20466 , n20812 , n20979 , n21027 , n21364 , n21426 , n21644 , 
n21673 , n21996 , n22322 , n22781 , n23011 , n23222 , n23320 , n23426 , n24047 , n24259 , 
n24356 , n25036 , n25255 , n25355 , n25447 , n25631 , n25694 , n25831 , n26329 , n26336 , 
n26659 , n26984 , n27447 , n27467 , n27501 , n27641 , n28093 , n28667 , n28946 , n28969 , 
n29261 , n29744 , n29788 , n30204 , n30292 , n30507 , n30625 , n30646 , n30986 , n31606 , 
n31803 , n32205 , n32329 , n32665 , n32697 , n33004 , n33116 , n33248 , n34201 , n34245 , 
n34484 , n34571 , n34820 , n34903 , n34923 , n35029 , n35111 , n35618 , n35924 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , 
n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , 
n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , 
n29 , n30 , n31 , n32 , n33 , n34 , n35 , n37 , n38 , n39 , 
n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
n140 , n141 , n142 , n143 , n144 , n145 , n146 , n148 , n149 , n150 , 
n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , 
n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , 
n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , 
n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , 
n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , 
n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , 
n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , 
n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , 
n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , 
n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , 
n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , 
n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , 
n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , 
n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , 
n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , 
n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , 
n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , 
n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , 
n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , 
n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , 
n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , 
n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , 
n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , 
n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , 
n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , 
n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , 
n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , 
n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , 
n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , 
n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , 
n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , 
n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , 
n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , 
n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , 
n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , 
n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , 
n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , 
n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , 
n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , 
n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , 
n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , 
n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , 
n691 , n692 , n693 , n694 , n695 , n696 , n698 , n699 , n700 , n701 , 
n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , 
n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , 
n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , 
n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , 
n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , 
n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , 
n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , 
n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , 
n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , 
n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n801 , n802 , 
n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , 
n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , 
n823 , n824 , n825 , n826 , n827 , n828 , n829 , n831 , n832 , n833 , 
n834 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , 
n845 , n846 , n847 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , 
n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , 
n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , 
n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , 
n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , 
n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , 
n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , 
n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , 
n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , 
n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , 
n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , 
n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , 
n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , 
n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , 
n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , 
n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , 
n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , 
n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , 
n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , 
n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , 
n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , 
n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , 
n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , 
n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , 
n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , 
n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , 
n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , 
n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , 
n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , 
n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , 
n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , 
n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , 
n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , 
n1176 , n1177 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , 
n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , 
n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , 
n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , 
n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , 
n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , 
n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , 
n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , 
n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , 
n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1276 , n1277 , n1278 , 
n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , 
n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , 
n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , 
n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , 
n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , 
n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1337 , n1338 , n1339 , 
n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
n1710 , n1711 , n1712 , n1713 , n1714 , n1716 , n1717 , n1718 , n1719 , n1720 , 
n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , 
n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , 
n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , 
n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , 
n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , 
n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , 
n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , 
n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , 
n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , 
n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , 
n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , 
n1831 , n1832 , n1833 , n1834 , n1835 , n1837 , n1838 , n1839 , n1840 , n1841 , 
n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , 
n1853 , n1854 , n1855 , n1856 , n1857 , n1859 , n1860 , n1861 , n1862 , n1863 , 
n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , 
n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , 
n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , 
n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , 
n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , 
n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , 
n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , 
n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , 
n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1951 , n1952 , n1953 , n1954 , 
n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , 
n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , 
n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , 
n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , 
n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2002 , n2003 , n2004 , n2005 , 
n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , 
n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , 
n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , 
n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , 
n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , 
n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , 
n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , 
n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , 
n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , 
n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2105 , n2106 , 
n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , 
n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , 
n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , 
n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , 
n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , 
n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , 
n2167 , n2168 , n2169 , n2170 , n2171 , n2173 , n2174 , n2175 , n2176 , n2177 , 
n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , 
n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , 
n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , 
n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , 
n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , 
n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , 
n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , 
n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , 
n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , 
n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , 
n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , 
n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , 
n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , 
n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , 
n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , 
n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , 
n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , 
n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , 
n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2367 , n2368 , 
n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , 
n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , 
n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , 
n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , 
n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , 
n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , 
n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , 
n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , 
n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , 
n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , 
n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , 
n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
n2760 , n2761 , n2762 , n2763 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , 
n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , 
n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , 
n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , 
n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , 
n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , 
n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , 
n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , 
n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , 
n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , 
n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , 
n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , 
n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , 
n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , 
n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , 
n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , 
n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , 
n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , 
n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , 
n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , 
n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , 
n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , 
n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , 
n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , 
n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , 
n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , 
n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , 
n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , 
n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , 
n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , 
n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , 
n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , 
n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , 
n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , 
n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , 
n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , 
n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , 
n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , 
n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , 
n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , 
n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , 
n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , 
n3201 , n3202 , n3203 , n3204 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , 
n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , 
n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , 
n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , 
n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , 
n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , 
n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , 
n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , 
n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , 
n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , 
n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , 
n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , 
n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , 
n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , 
n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , 
n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , 
n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , 
n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , 
n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , 
n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , 
n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , 
n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , 
n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , 
n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , 
n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , 
n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , 
n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , 
n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , 
n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , 
n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , 
n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , 
n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , 
n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , 
n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , 
n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , 
n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , 
n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , 
n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , 
n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , 
n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , 
n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , 
n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , 
n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , 
n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , 
n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , 
n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , 
n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , 
n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , 
n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , 
n3693 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , 
n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , 
n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , 
n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , 
n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3742 , n3743 , n3744 , 
n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , 
n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , 
n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , 
n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , 
n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , 
n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , 
n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , 
n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , 
n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , 
n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , 
n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , 
n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , 
n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , 
n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , 
n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , 
n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , 
n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , 
n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , 
n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , 
n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , 
n3945 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , 
n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , 
n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , 
n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , 
n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , 
n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , 
n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , 
n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , 
n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , 
n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , 
n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , 
n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , 
n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , 
n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , 
n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , 
n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , 
n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , 
n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , 
n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , 
n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , 
n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , 
n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , 
n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , 
n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , 
n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , 
n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , 
n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , 
n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , 
n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , 
n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , 
n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , 
n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , 
n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , 
n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , 
n4286 , n4287 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , 
n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , 
n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , 
n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , 
n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , 
n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , 
n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , 
n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , 
n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , 
n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , 
n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , 
n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , 
n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , 
n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , 
n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , 
n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , 
n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , 
n4457 , n4458 , n4459 , n4460 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , 
n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , 
n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , 
n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , 
n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , 
n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , 
n4518 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , 
n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , 
n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , 
n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , 
n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , 
n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , 
n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , 
n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , 
n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , 
n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , 
n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , 
n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , 
n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , 
n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , 
n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , 
n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , 
n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , 
n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , 
n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , 
n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , 
n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , 
n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , 
n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , 
n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4759 , 
n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , 
n4770 , n4771 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4789 , n4790 , n4791 , 
n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , 
n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , 
n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , 
n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , 
n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , 
n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , 
n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , 
n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , 
n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4879 , n4880 , n4881 , n4882 , 
n4883 , n4884 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , 
n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , 
n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , 
n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , 
n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , 
n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , 
n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , 
n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4961 , n4963 , n4964 , n4965 , 
n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , 
n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , 
n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , 
n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , 
n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , 
n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , 
n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , 
n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , 
n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , 
n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , 
n5066 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , 
n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , 
n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , 
n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , 
n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , 
n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , 
n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , 
n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , 
n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , 
n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , 
n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , 
n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , 
n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , 
n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , 
n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , 
n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , 
n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , 
n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , 
n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , 
n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , 
n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , 
n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , 
n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , 
n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , 
n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , 
n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , 
n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5336 , n5337 , n5338 , 
n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , 
n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , 
n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , 
n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , 
n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , 
n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , 
n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , 
n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , 
n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , 
n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , 
n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , 
n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , 
n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , 
n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , 
n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , 
n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , 
n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , 
n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , 
n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , 
n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , 
n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , 
n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , 
n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , 
n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , 
n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , 
n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , 
n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , 
n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , 
n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , 
n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , 
n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , 
n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , 
n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , 
n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , 
n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , 
n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , 
n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , 
n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , 
n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , 
n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5739 , 
n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , 
n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , 
n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , 
n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , 
n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , 
n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , 
n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , 
n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , 
n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , 
n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , 
n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , 
n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , 
n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , 
n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , 
n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , 
n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , 
n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , 
n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , 
n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , 
n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , 
n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , 
n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , 
n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , 
n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , 
n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , 
n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , 
n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , 
n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , 
n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , 
n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , 
n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , 
n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , 
n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , 
n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , 
n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , 
n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , 
n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , 
n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , 
n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , 
n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , 
n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , 
n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , 
n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , 
n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , 
n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , 
n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , 
n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , 
n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , 
n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6227 , n6228 , n6229 , n6230 , 
n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , 
n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , 
n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , 
n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , 
n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , 
n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , 
n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , 
n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , 
n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , 
n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , 
n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , 
n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , 
n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , 
n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , 
n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , 
n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , 
n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , 
n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , 
n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , 
n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , 
n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , 
n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , 
n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , 
n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , 
n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , 
n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , 
n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , 
n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , 
n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , 
n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , 
n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , 
n6541 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , 
n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , 
n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , 
n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , 
n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , 
n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , 
n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , 
n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , 
n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , 
n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , 
n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , 
n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , 
n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , 
n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , 
n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , 
n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , 
n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , 
n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , 
n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , 
n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , 
n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , 
n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , 
n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , 
n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , 
n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , 
n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , 
n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , 
n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , 
n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , 
n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , 
n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , 
n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , 
n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , 
n6872 , n6873 , n6874 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , 
n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , 
n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , 
n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , 
n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , 
n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , 
n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , 
n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , 
n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , 
n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , 
n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , 
n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , 
n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , 
n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , 
n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , 
n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , 
n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , 
n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , 
n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , 
n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , 
n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , 
n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , 
n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , 
n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , 
n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , 
n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , 
n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , 
n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , 
n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , 
n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , 
n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , 
n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , 
n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , 
n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , 
n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , 
n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , 
n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , 
n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , 
n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , 
n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , 
n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , 
n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , 
n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , 
n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , 
n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , 
n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , 
n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , 
n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , 
n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , 
n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , 
n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , 
n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , 
n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , 
n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , 
n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , 
n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , 
n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , 
n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , 
n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , 
n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , 
n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , 
n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , 
n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , 
n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , 
n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , 
n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , 
n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7541 , n7542 , n7543 , n7544 , 
n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , 
n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , 
n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , 
n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , 
n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , 
n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , 
n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , 
n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , 
n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , 
n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , 
n7645 , n7646 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , 
n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , 
n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , 
n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , 
n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , 
n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , 
n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , 
n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , 
n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , 
n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , 
n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , 
n7756 , n7757 , n7758 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , 
n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , 
n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , 
n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , 
n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , 
n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , 
n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , 
n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , 
n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , 
n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , 
n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , 
n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , 
n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , 
n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , 
n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , 
n7907 , n7908 , n7909 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , 
n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , 
n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , 
n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , 
n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , 
n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , 
n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , 
n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , 
n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , 
n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , 
n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , 
n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , 
n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , 
n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , 
n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , 
n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , 
n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , 
n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , 
n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , 
n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , 
n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , 
n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , 
n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , 
n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , 
n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , 
n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , 
n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , 
n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , 
n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , 
n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , 
n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , 
n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , 
n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , 
n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , 
n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , 
n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , 
n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , 
n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , 
n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , 
n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , 
n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , 
n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , 
n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , 
n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , 
n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , 
n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , 
n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , 
n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , 
n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , 
n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , 
n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , 
n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , 
n8428 , n8429 , n8430 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , 
n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , 
n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , 
n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , 
n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , 
n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , 
n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , 
n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , 
n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , 
n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , 
n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , 
n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , 
n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , 
n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , 
n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , 
n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , 
n8590 , n8591 , n8592 , n8593 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , 
n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , 
n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , 
n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , 
n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , 
n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , 
n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , 
n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , 
n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , 
n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , 
n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , 
n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , 
n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , 
n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , 
n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , 
n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , 
n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , 
n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , 
n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , 
n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , 
n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , 
n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , 
n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , 
n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , 
n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , 
n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , 
n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , 
n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , 
n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , 
n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , 
n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , 
n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , 
n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , 
n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , 
n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , 
n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , 
n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , 
n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , 
n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , 
n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , 
n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , 
n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , 
n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , 
n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , 
n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , 
n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , 
n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , 
n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , 
n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , 
n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , 
n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , 
n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , 
n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , 
n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , 
n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , 
n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , 
n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , 
n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , 
n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , 
n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , 
n9191 , n9192 , n9193 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , 
n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , 
n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , 
n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , 
n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , 
n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , 
n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , 
n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , 
n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , 
n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9292 , 
n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , 
n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , 
n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , 
n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , 
n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , 
n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , 
n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , 
n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , 
n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , 
n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , 
n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , 
n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , 
n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , 
n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , 
n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , 
n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , 
n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , 
n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , 
n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , 
n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , 
n9493 , n9494 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , 
n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , 
n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , 
n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , 
n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , 
n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , 
n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , 
n9564 , n9565 , n9566 , n9567 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , 
n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , 
n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , 
n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , 
n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , 
n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , 
n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , 
n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , 
n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , 
n9655 , n9656 , n9657 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , 
n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , 
n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , 
n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , 
n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , 
n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , 
n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , 
n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , 
n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , 
n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , 
n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , 
n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , 
n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , 
n9786 , n9787 , n9788 , n9790 , n9791 , n9792 , n9794 , n9795 , n9796 , n9797 , 
n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , 
n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , 
n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , 
n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , 
n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , 
n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , 
n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , 
n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , 
n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , 
n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , 
n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , 
n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , 
n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , 
n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , 
n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , 
n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , 
n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , 
n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , 
n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , 
n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , 
n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , 
n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , 
n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , 
n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , 
n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , 
n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , 
n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , 
n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , 
n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , 
n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , 
n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , 
n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , 
n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , 
n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , 
n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , 
n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , 
n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , 
n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , 
n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , 
n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , 
n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , 
n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , 
n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , 
n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , 
n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , 
n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , 
n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , 
n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , 
n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , 
n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10299 , 
n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , 
n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , 
n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , 
n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , 
n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , 
n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , 
n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , 
n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , 
n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , 
n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , 
n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , 
n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , 
n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , 
n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , 
n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , 
n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , 
n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , 
n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , 
n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , 
n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , 
n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , 
n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , 
n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , 
n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , 
n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , 
n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , 
n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , 
n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , 
n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , 
n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , 
n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , 
n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , 
n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , 
n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , 
n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , 
n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , 
n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , 
n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , 
n10680 , n10681 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , 
n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , 
n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , 
n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , 
n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , 
n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , 
n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , 
n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , 
n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10769 , n10770 , n10771 , 
n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , 
n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , 
n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , 
n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , 
n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , 
n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , 
n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , 
n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , 
n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , 
n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , 
n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , 
n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , 
n10893 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , 
n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , 
n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , 
n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , 
n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , 
n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , 
n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , 
n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , 
n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , 
n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , 
n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , 
n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , 
n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , 
n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , 
n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , 
n11044 , n11045 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , 
n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , 
n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , 
n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , 
n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , 
n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , 
n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , 
n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , 
n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , 
n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , 
n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , 
n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , 
n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , 
n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , 
n11185 , n11186 , n11187 , n11188 , n11189 , n11191 , n11192 , n11193 , n11194 , n11195 , 
n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , 
n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , 
n11216 , n11217 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , 
n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , 
n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11244 , n11245 , n11246 , n11247 , 
n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , 
n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , 
n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , 
n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , 
n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , 
n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , 
n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , 
n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , 
n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , 
n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , 
n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , 
n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , 
n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , 
n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , 
n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , 
n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , 
n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , 
n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , 
n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , 
n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , 
n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11456 , n11457 , n11458 , 
n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , 
n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , 
n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , 
n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , 
n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , 
n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , 
n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , 
n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , 
n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , 
n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , 
n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , 
n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , 
n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , 
n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , 
n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , 
n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , 
n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , 
n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , 
n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , 
n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , 
n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , 
n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , 
n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , 
n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , 
n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , 
n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , 
n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , 
n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , 
n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , 
n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , 
n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , 
n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , 
n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , 
n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , 
n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , 
n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , 
n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , 
n11829 , n11830 , n11831 , n11832 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , 
n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , 
n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , 
n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , 
n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , 
n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , 
n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , 
n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , 
n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , 
n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , 
n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , 
n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , 
n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , 
n11960 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , 
n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , 
n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , 
n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , 
n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , 
n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , 
n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , 
n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , 
n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , 
n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , 
n12061 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , 
n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , 
n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , 
n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , 
n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , 
n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , 
n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , 
n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , 
n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , 
n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , 
n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , 
n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , 
n12182 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , 
n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , 
n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , 
n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , 
n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , 
n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , 
n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , 
n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , 
n12263 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , 
n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , 
n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , 
n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , 
n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , 
n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , 
n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , 
n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , 
n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , 
n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , 
n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , 
n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , 
n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , 
n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , 
n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , 
n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , 
n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , 
n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , 
n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , 
n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , 
n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , 
n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , 
n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , 
n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , 
n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , 
n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , 
n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , 
n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , 
n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , 
n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , 
n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , 
n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , 
n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , 
n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , 
n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , 
n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , 
n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , 
n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , 
n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , 
n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , 
n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , 
n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , 
n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , 
n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , 
n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , 
n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , 
n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , 
n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , 
n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , 
n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , 
n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , 
n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , 
n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , 
n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , 
n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , 
n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , 
n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , 
n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , 
n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , 
n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , 
n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , 
n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , 
n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , 
n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , 
n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , 
n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , 
n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , 
n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , 
n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , 
n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , 
n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , 
n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , 
n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , 
n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , 
n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , 
n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , 
n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , 
n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , 
n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , 
n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , 
n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , 
n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , 
n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , 
n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , 
n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , 
n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , 
n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , 
n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , 
n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , 
n13154 , n13155 , n13156 , n13157 , n13158 , n13160 , n13161 , n13162 , n13163 , n13164 , 
n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , 
n13175 , n13176 , n13177 , n13178 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , 
n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , 
n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , 
n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , 
n13216 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , 
n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , 
n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , 
n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , 
n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , 
n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , 
n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , 
n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , 
n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , 
n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , 
n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , 
n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , 
n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , 
n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , 
n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , 
n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , 
n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , 
n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , 
n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , 
n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13414 , n13415 , n13416 , n13417 , 
n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , 
n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , 
n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , 
n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13456 , n13457 , n13458 , 
n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , 
n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , 
n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , 
n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , 
n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , 
n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , 
n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , 
n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , 
n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , 
n13549 , n13550 , n13551 , n13552 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , 
n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , 
n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , 
n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , 
n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , 
n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , 
n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , 
n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , 
n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , 
n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , 
n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , 
n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , 
n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , 
n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , 
n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , 
n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , 
n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , 
n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , 
n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , 
n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , 
n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , 
n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , 
n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , 
n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , 
n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , 
n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , 
n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , 
n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , 
n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , 
n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , 
n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , 
n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , 
n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , 
n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , 
n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , 
n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , 
n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , 
n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , 
n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , 
n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , 
n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , 
n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13968 , n13969 , n13970 , 
n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , 
n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , 
n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , 
n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , 
n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , 
n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , 
n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , 
n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , 
n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , 
n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , 
n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , 
n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , 
n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , 
n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , 
n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , 
n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , 
n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , 
n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , 
n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , 
n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , 
n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , 
n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , 
n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , 
n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , 
n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , 
n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , 
n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , 
n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , 
n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , 
n14262 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , 
n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , 
n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , 
n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , 
n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , 
n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , 
n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , 
n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , 
n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , 
n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , 
n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , 
n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , 
n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , 
n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , 
n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , 
n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , 
n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , 
n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , 
n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , 
n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , 
n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , 
n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , 
n14483 , n14484 , n14485 , n14486 , n14487 , n14489 , n14490 , n14491 , n14492 , n14493 , 
n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , 
n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , 
n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , 
n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , 
n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , 
n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , 
n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , 
n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , 
n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , 
n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , 
n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , 
n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , 
n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , 
n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , 
n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , 
n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , 
n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , 
n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , 
n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , 
n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , 
n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , 
n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , 
n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , 
n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , 
n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , 
n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , 
n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , 
n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , 
n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , 
n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , 
n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , 
n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , 
n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , 
n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , 
n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , 
n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , 
n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , 
n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , 
n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , 
n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , 
n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , 
n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , 
n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , 
n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , 
n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , 
n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , 
n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , 
n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , 
n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , 
n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , 
n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , 
n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , 
n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , 
n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , 
n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , 
n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , 
n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , 
n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , 
n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , 
n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , 
n15094 , n15096 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , 
n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , 
n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , 
n15126 , n15127 , n15128 , n15129 , n15130 , n15132 , n15133 , n15134 , n15135 , n15136 , 
n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , 
n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , 
n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , 
n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , 
n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , 
n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , 
n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , 
n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , 
n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , 
n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , 
n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , 
n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , 
n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , 
n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , 
n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , 
n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , 
n15297 , n15298 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , 
n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , 
n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , 
n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , 
n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , 
n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15358 , 
n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , 
n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , 
n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , 
n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , 
n15399 , n15400 , n15401 , n15402 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , 
n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , 
n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , 
n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , 
n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , 
n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , 
n15460 , n15461 , n15462 , n15463 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , 
n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , 
n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , 
n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15498 , n15499 , n15500 , n15501 , 
n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , 
n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , 
n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , 
n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , 
n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , 
n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , 
n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15571 , n15572 , 
n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , 
n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , 
n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , 
n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , 
n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , 
n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , 
n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , 
n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , 
n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , 
n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , 
n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , 
n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , 
n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , 
n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , 
n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , 
n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , 
n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , 
n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , 
n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , 
n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , 
n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , 
n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , 
n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , 
n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , 
n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , 
n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , 
n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , 
n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , 
n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , 
n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , 
n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , 
n15883 , n15884 , n15885 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , 
n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , 
n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , 
n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , 
n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , 
n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , 
n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , 
n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , 
n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , 
n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , 
n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , 
n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , 
n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , 
n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , 
n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , 
n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , 
n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , 
n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , 
n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , 
n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , 
n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , 
n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , 
n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , 
n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , 
n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , 
n16134 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , 
n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , 
n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , 
n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , 
n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , 
n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , 
n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , 
n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , 
n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , 
n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , 
n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , 
n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , 
n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , 
n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , 
n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , 
n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , 
n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , 
n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , 
n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , 
n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , 
n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , 
n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , 
n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , 
n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , 
n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , 
n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , 
n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , 
n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , 
n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , 
n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , 
n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , 
n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , 
n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , 
n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , 
n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , 
n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , 
n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , 
n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , 
n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16525 , 
n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , 
n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , 
n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , 
n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , 
n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , 
n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , 
n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , 
n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , 
n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , 
n16616 , n16617 , n16618 , n16619 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , 
n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , 
n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , 
n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , 
n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , 
n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , 
n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , 
n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , 
n16697 , n16698 , n16699 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , 
n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , 
n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , 
n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , 
n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , 
n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , 
n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , 
n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , 
n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , 
n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , 
n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , 
n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16818 , 
n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , 
n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , 
n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , 
n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , 
n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , 
n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , 
n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , 
n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16896 , n16897 , n16898 , n16900 , 
n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , 
n16911 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , 
n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , 
n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , 
n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , 
n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16962 , n16963 , 
n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , 
n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , 
n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , 
n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , 
n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , 
n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , 
n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , 
n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , 
n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , 
n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , 
n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , 
n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , 
n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , 
n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , 
n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , 
n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , 
n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , 
n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , 
n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , 
n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , 
n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , 
n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , 
n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , 
n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , 
n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , 
n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , 
n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , 
n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , 
n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , 
n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , 
n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , 
n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , 
n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , 
n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , 
n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , 
n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , 
n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , 
n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , 
n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , 
n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , 
n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , 
n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , 
n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , 
n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , 
n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , 
n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , 
n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , 
n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , 
n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , 
n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , 
n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , 
n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , 
n17484 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , 
n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , 
n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , 
n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , 
n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , 
n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , 
n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , 
n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , 
n17565 , n17566 , n17567 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , 
n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , 
n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , 
n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , 
n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , 
n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , 
n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , 
n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , 
n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , 
n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , 
n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , 
n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , 
n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , 
n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17703 , n17704 , n17705 , n17706 , 
n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , 
n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , 
n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , 
n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , 
n17747 , n17748 , n17749 , n17750 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , 
n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , 
n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , 
n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , 
n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , 
n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , 
n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , 
n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , 
n17828 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , 
n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , 
n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , 
n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , 
n17869 , n17870 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , 
n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , 
n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , 
n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , 
n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , 
n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , 
n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , 
n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , 
n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , 
n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , 
n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , 
n17980 , n17981 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , 
n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , 
n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , 
n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , 
n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , 
n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , 
n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , 
n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , 
n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , 
n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , 
n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , 
n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , 
n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , 
n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , 
n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , 
n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , 
n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , 
n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , 
n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , 
n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , 
n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , 
n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , 
n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , 
n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , 
n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , 
n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , 
n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , 
n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , 
n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , 
n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , 
n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , 
n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , 
n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , 
n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , 
n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , 
n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , 
n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , 
n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , 
n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , 
n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18380 , n18381 , 
n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , 
n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , 
n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , 
n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , 
n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , 
n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , 
n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , 
n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , 
n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , 
n18472 , n18473 , n18474 , n18475 , n18476 , n18478 , n18479 , n18480 , n18481 , n18482 , 
n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , 
n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , 
n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , 
n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , 
n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , 
n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , 
n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , 
n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , 
n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , 
n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , 
n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , 
n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , 
n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , 
n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , 
n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , 
n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , 
n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , 
n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , 
n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , 
n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , 
n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , 
n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , 
n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , 
n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , 
n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , 
n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , 
n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , 
n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , 
n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , 
n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , 
n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , 
n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , 
n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , 
n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , 
n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , 
n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18842 , n18843 , 
n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , 
n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , 
n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , 
n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , 
n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , 
n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , 
n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18913 , n18914 , 
n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , 
n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , 
n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , 
n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , 
n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , 
n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , 
n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , 
n18985 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , 
n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , 
n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , 
n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , 
n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , 
n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , 
n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , 
n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , 
n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , 
n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19085 , n19086 , 
n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , 
n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , 
n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , 
n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , 
n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , 
n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , 
n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , 
n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , 
n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , 
n19177 , n19178 , n19179 , n19180 , n19181 , n19183 , n19184 , n19185 , n19186 , n19187 , 
n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , 
n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , 
n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , 
n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , 
n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , 
n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , 
n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , 
n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , 
n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , 
n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , 
n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , 
n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , 
n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , 
n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , 
n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , 
n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , 
n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , 
n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , 
n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , 
n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , 
n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , 
n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , 
n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , 
n19419 , n19420 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , 
n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , 
n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , 
n19450 , n19451 , n19452 , n19453 , n19455 , n19456 , n19457 , n19459 , n19460 , n19461 , 
n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , 
n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , 
n19482 , n19483 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , 
n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , 
n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , 
n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , 
n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , 
n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , 
n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19552 , n19553 , 
n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , 
n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , 
n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , 
n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , 
n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , 
n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , 
n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , 
n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , 
n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , 
n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , 
n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , 
n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , 
n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , 
n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , 
n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , 
n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , 
n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , 
n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , 
n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , 
n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , 
n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , 
n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , 
n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , 
n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , 
n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , 
n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , 
n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , 
n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , 
n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , 
n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , 
n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , 
n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , 
n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , 
n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , 
n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , 
n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , 
n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , 
n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , 
n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , 
n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , 
n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , 
n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , 
n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , 
n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , 
n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , 
n20005 , n20006 , n20007 , n20008 , n20009 , n20011 , n20012 , n20013 , n20014 , n20015 , 
n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , 
n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , 
n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , 
n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , 
n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , 
n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , 
n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , 
n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , 
n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , 
n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , 
n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , 
n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , 
n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , 
n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , 
n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , 
n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , 
n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , 
n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , 
n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , 
n20206 , n20207 , n20208 , n20209 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , 
n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , 
n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , 
n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , 
n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , 
n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , 
n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , 
n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , 
n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , 
n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , 
n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , 
n20317 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , 
n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , 
n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , 
n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , 
n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , 
n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , 
n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , 
n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , 
n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , 
n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , 
n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , 
n20429 , n20430 , n20431 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , 
n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , 
n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , 
n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20467 , n20468 , n20469 , n20470 , 
n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , 
n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , 
n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , 
n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , 
n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , 
n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , 
n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , 
n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , 
n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , 
n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , 
n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , 
n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , 
n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , 
n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , 
n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , 
n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , 
n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , 
n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , 
n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , 
n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , 
n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , 
n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , 
n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , 
n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , 
n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , 
n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , 
n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , 
n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , 
n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , 
n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , 
n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , 
n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , 
n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , 
n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , 
n20811 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , 
n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , 
n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , 
n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , 
n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , 
n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , 
n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , 
n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , 
n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , 
n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , 
n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , 
n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , 
n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , 
n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , 
n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , 
n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , 
n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20980 , n20981 , n20982 , 
n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , 
n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , 
n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , 
n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , 
n21023 , n21024 , n21025 , n21026 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , 
n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , 
n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , 
n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , 
n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , 
n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , 
n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , 
n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , 
n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , 
n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , 
n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , 
n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , 
n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , 
n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , 
n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , 
n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , 
n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , 
n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , 
n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , 
n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , 
n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , 
n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , 
n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , 
n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , 
n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , 
n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21282 , n21283 , n21284 , 
n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , 
n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , 
n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , 
n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , 
n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , 
n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , 
n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , 
n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21365 , 
n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , 
n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , 
n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , 
n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , 
n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , 
n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , 
n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , 
n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , 
n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , 
n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , 
n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , 
n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , 
n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , 
n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , 
n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , 
n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , 
n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , 
n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , 
n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , 
n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , 
n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , 
n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , 
n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , 
n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , 
n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , 
n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , 
n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , 
n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21645 , n21646 , n21647 , 
n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , 
n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , 
n21668 , n21669 , n21670 , n21671 , n21672 , n21674 , n21675 , n21676 , n21677 , n21678 , 
n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , 
n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , 
n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , 
n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , 
n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , 
n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21738 , n21739 , 
n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , 
n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , 
n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , 
n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , 
n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , 
n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , 
n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , 
n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , 
n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , 
n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , 
n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , 
n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , 
n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , 
n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , 
n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , 
n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , 
n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , 
n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , 
n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , 
n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , 
n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , 
n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , 
n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , 
n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , 
n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , 
n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21997 , n21998 , n21999 , n22000 , 
n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , 
n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , 
n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , 
n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , 
n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , 
n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , 
n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , 
n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , 
n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , 
n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , 
n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , 
n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , 
n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , 
n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , 
n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , 
n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , 
n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , 
n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , 
n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , 
n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , 
n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , 
n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , 
n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , 
n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , 
n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , 
n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , 
n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , 
n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , 
n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , 
n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , 
n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , 
n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , 
n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , 
n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , 
n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , 
n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , 
n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , 
n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , 
n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , 
n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , 
n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , 
n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , 
n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , 
n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , 
n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , 
n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , 
n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , 
n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , 
n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , 
n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , 
n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , 
n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , 
n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , 
n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , 
n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , 
n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , 
n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , 
n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , 
n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , 
n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , 
n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , 
n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , 
n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , 
n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , 
n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , 
n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , 
n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , 
n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , 
n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , 
n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , 
n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , 
n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , 
n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , 
n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , 
n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , 
n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , 
n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , 
n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22782 , n22783 , 
n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , 
n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , 
n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , 
n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , 
n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , 
n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , 
n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , 
n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , 
n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , 
n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , 
n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , 
n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , 
n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , 
n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , 
n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , 
n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , 
n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , 
n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , 
n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , 
n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22981 , n22982 , n22983 , n22984 , 
n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , 
n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , 
n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23012 , n23013 , n23014 , n23015 , 
n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , 
n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , 
n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , 
n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , 
n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , 
n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , 
n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , 
n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , 
n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , 
n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , 
n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , 
n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , 
n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , 
n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , 
n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , 
n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , 
n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , 
n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , 
n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , 
n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , 
n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23223 , n23224 , n23225 , n23226 , 
n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , 
n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , 
n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , 
n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , 
n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , 
n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , 
n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , 
n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , 
n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , 
n23317 , n23318 , n23319 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , 
n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , 
n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , 
n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , 
n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , 
n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , 
n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , 
n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , 
n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , 
n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , 
n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23427 , n23428 , 
n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , 
n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , 
n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , 
n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , 
n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , 
n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , 
n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , 
n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , 
n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , 
n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , 
n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , 
n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , 
n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , 
n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , 
n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , 
n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , 
n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , 
n23599 , n23600 , n23601 , n23602 , n23603 , n23605 , n23606 , n23607 , n23608 , n23609 , 
n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , 
n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , 
n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , 
n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , 
n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , 
n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , 
n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , 
n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , 
n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , 
n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , 
n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , 
n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , 
n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , 
n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , 
n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , 
n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , 
n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , 
n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , 
n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , 
n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , 
n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , 
n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , 
n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , 
n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , 
n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , 
n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , 
n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , 
n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , 
n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , 
n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , 
n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , 
n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , 
n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , 
n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , 
n23950 , n23951 , n23952 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , 
n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , 
n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , 
n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , 
n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , 
n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , 
n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , 
n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , 
n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , 
n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24048 , n24049 , n24050 , n24051 , 
n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , 
n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , 
n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , 
n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , 
n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , 
n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , 
n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , 
n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , 
n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , 
n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , 
n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , 
n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , 
n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , 
n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , 
n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , 
n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , 
n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , 
n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , 
n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , 
n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , 
n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24260 , n24261 , n24262 , 
n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , 
n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , 
n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , 
n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , 
n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , 
n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , 
n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24333 , 
n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , 
n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , 
n24354 , n24355 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , 
n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24372 , n24373 , n24374 , n24375 , 
n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , 
n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , 
n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , 
n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , 
n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , 
n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24435 , n24436 , 
n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , 
n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , 
n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , 
n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , 
n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , 
n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , 
n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , 
n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , 
n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , 
n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , 
n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , 
n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , 
n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , 
n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , 
n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , 
n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , 
n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , 
n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , 
n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , 
n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , 
n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , 
n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , 
n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , 
n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , 
n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , 
n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , 
n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , 
n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , 
n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , 
n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , 
n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , 
n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , 
n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , 
n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , 
n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , 
n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , 
n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , 
n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , 
n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , 
n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , 
n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , 
n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , 
n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , 
n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , 
n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , 
n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , 
n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , 
n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , 
n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , 
n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , 
n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , 
n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , 
n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , 
n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , 
n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , 
n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , 
n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , 
n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , 
n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , 
n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25037 , 
n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , 
n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , 
n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , 
n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , 
n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , 
n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , 
n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , 
n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , 
n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , 
n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , 
n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , 
n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , 
n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , 
n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25175 , n25176 , n25177 , n25178 , 
n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , 
n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , 
n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , 
n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , 
n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , 
n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , 
n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , 
n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25256 , n25257 , n25258 , n25259 , 
n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , 
n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , 
n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , 
n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , 
n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , 
n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , 
n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , 
n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , 
n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , 
n25350 , n25351 , n25352 , n25353 , n25354 , n25356 , n25357 , n25358 , n25359 , n25360 , 
n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , 
n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , 
n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , 
n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , 
n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , 
n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , 
n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , 
n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , 
n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25448 , n25449 , n25450 , n25451 , 
n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , 
n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , 
n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , 
n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , 
n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , 
n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , 
n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , 
n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , 
n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , 
n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , 
n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , 
n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , 
n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , 
n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , 
n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , 
n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , 
n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , 
n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25632 , n25633 , 
n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , 
n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , 
n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , 
n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , 
n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , 
n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , 
n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , 
n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , 
n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , 
n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , 
n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , 
n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , 
n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , 
n25765 , n25766 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , 
n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , 
n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , 
n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , 
n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , 
n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , 
n25826 , n25827 , n25828 , n25829 , n25830 , n25832 , n25833 , n25834 , n25835 , n25836 , 
n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , 
n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , 
n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , 
n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , 
n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , 
n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , 
n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , 
n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , 
n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , 
n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , 
n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , 
n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , 
n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , 
n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , 
n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , 
n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , 
n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , 
n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , 
n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , 
n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , 
n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , 
n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , 
n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , 
n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , 
n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , 
n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , 
n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , 
n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , 
n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , 
n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , 
n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , 
n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , 
n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , 
n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , 
n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , 
n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , 
n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , 
n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , 
n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , 
n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , 
n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , 
n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , 
n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , 
n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , 
n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , 
n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , 
n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , 
n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , 
n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , 
n26327 , n26328 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26337 , n26338 , 
n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , 
n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , 
n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , 
n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , 
n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , 
n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , 
n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , 
n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , 
n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , 
n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , 
n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , 
n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , 
n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , 
n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , 
n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , 
n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , 
n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , 
n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , 
n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , 
n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , 
n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , 
n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , 
n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , 
n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , 
n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , 
n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , 
n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , 
n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , 
n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , 
n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , 
n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , 
n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , 
n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , 
n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , 
n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , 
n26690 , n26691 , n26692 , n26693 , n26694 , n26696 , n26697 , n26698 , n26699 , n26700 , 
n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , 
n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , 
n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , 
n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , 
n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , 
n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , 
n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , 
n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , 
n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , 
n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , 
n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , 
n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , 
n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , 
n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , 
n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , 
n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , 
n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , 
n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , 
n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , 
n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , 
n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , 
n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , 
n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , 
n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , 
n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , 
n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , 
n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , 
n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , 
n26982 , n26983 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , 
n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , 
n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27010 , n27011 , n27012 , n27013 , 
n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , 
n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , 
n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , 
n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , 
n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , 
n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , 
n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , 
n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , 
n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , 
n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , 
n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , 
n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , 
n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , 
n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , 
n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , 
n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , 
n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , 
n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , 
n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , 
n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , 
n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , 
n27224 , n27225 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , 
n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , 
n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , 
n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , 
n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , 
n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , 
n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27292 , n27293 , n27294 , n27295 , 
n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , 
n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , 
n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , 
n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , 
n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , 
n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , 
n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , 
n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , 
n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , 
n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , 
n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , 
n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , 
n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , 
n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , 
n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , 
n27446 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , 
n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , 
n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , 
n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , 
n27488 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , 
n27499 , n27500 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , 
n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , 
n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , 
n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , 
n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , 
n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , 
n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , 
n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , 
n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , 
n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , 
n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , 
n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , 
n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27628 , n27629 , n27630 , 
n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , 
n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , 
n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , 
n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , 
n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , 
n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , 
n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , 
n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , 
n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , 
n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , 
n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , 
n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , 
n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , 
n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , 
n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , 
n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , 
n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , 
n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , 
n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , 
n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , 
n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , 
n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , 
n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , 
n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , 
n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , 
n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , 
n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , 
n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , 
n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , 
n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , 
n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , 
n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , 
n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , 
n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , 
n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , 
n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , 
n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , 
n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , 
n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , 
n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , 
n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , 
n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , 
n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , 
n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , 
n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , 
n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , 
n28092 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , 
n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , 
n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , 
n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , 
n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , 
n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , 
n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , 
n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , 
n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , 
n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , 
n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , 
n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , 
n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , 
n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , 
n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , 
n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , 
n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , 
n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , 
n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , 
n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , 
n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , 
n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , 
n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , 
n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , 
n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , 
n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , 
n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , 
n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , 
n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , 
n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , 
n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , 
n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , 
n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , 
n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , 
n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , 
n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , 
n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , 
n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , 
n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , 
n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , 
n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , 
n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , 
n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , 
n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , 
n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , 
n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , 
n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , 
n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , 
n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , 
n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , 
n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , 
n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , 
n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , 
n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , 
n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , 
n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , 
n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , 
n28664 , n28665 , n28666 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , 
n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , 
n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , 
n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , 
n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , 
n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , 
n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , 
n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , 
n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , 
n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , 
n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , 
n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , 
n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , 
n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , 
n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , 
n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , 
n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , 
n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , 
n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , 
n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , 
n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , 
n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , 
n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , 
n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , 
n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , 
n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , 
n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , 
n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , 
n28945 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , 
n28956 , n28957 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , 
n28967 , n28968 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , 
n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , 
n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , 
n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , 
n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , 
n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , 
n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29038 , 
n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , 
n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , 
n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , 
n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , 
n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , 
n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , 
n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , 
n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , 
n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , 
n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , 
n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , 
n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , 
n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , 
n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , 
n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , 
n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , 
n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , 
n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , 
n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , 
n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , 
n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , 
n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , 
n29259 , n29260 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , 
n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , 
n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , 
n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , 
n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , 
n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , 
n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , 
n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , 
n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , 
n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , 
n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , 
n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , 
n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , 
n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , 
n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , 
n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , 
n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , 
n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , 
n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , 
n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , 
n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , 
n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , 
n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , 
n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , 
n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , 
n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , 
n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , 
n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , 
n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , 
n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , 
n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , 
n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , 
n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , 
n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , 
n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , 
n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , 
n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , 
n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , 
n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29650 , 
n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , 
n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , 
n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , 
n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , 
n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , 
n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , 
n29711 , n29712 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , 
n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29732 , 
n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , 
n29743 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , 
n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , 
n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , 
n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , 
n29784 , n29785 , n29786 , n29787 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , 
n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , 
n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , 
n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , 
n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , 
n29835 , n29836 , n29837 , n29838 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , 
n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , 
n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , 
n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , 
n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29885 , n29886 , 
n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , 
n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , 
n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , 
n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , 
n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , 
n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , 
n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , 
n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , 
n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , 
n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , 
n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , 
n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , 
n30007 , n30008 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30017 , n30018 , 
n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , 
n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , 
n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , 
n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , 
n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , 
n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , 
n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , 
n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , 
n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , 
n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , 
n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , 
n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , 
n30139 , n30140 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , 
n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , 
n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , 
n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , 
n30180 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , 
n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , 
n30201 , n30202 , n30203 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , 
n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , 
n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , 
n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , 
n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , 
n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , 
n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , 
n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , 
n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , 
n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , 
n30303 , n30304 , n30305 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , 
n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , 
n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , 
n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , 
n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , 
n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , 
n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , 
n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , 
n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , 
n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , 
n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , 
n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , 
n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , 
n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , 
n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , 
n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , 
n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , 
n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , 
n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , 
n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , 
n30504 , n30505 , n30506 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , 
n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , 
n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , 
n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , 
n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30554 , n30555 , 
n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , 
n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , 
n30576 , n30577 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , 
n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , 
n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , 
n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , 
n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30626 , n30627 , 
n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , 
n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30647 , n30648 , 
n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , 
n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , 
n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , 
n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , 
n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , 
n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , 
n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , 
n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , 
n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , 
n30739 , n30740 , n30741 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , 
n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , 
n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , 
n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , 
n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , 
n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , 
n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , 
n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , 
n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , 
n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , 
n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , 
n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , 
n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , 
n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , 
n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , 
n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , 
n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , 
n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , 
n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , 
n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , 
n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , 
n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , 
n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , 
n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , 
n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30987 , n30988 , n30989 , n30990 , 
n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , 
n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , 
n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , 
n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , 
n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , 
n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , 
n31051 , n31052 , n31053 , n31055 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , 
n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , 
n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , 
n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , 
n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , 
n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , 
n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , 
n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , 
n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , 
n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , 
n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , 
n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , 
n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , 
n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , 
n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , 
n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , 
n31213 , n31214 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , 
n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , 
n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , 
n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , 
n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , 
n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31273 , n31274 , 
n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , 
n31285 , n31286 , n31287 , n31288 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , 
n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , 
n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , 
n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , 
n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , 
n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , 
n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , 
n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , 
n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , 
n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , 
n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , 
n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , 
n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , 
n31416 , n31417 , n31418 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , 
n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , 
n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , 
n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , 
n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , 
n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , 
n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , 
n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , 
n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , 
n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , 
n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , 
n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , 
n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , 
n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , 
n31557 , n31558 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , 
n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , 
n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , 
n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , 
n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31607 , n31608 , 
n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , 
n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , 
n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , 
n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , 
n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , 
n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , 
n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , 
n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , 
n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , 
n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , 
n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , 
n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , 
n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , 
n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , 
n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , 
n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , 
n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , 
n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , 
n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , 
n31800 , n31801 , n31802 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , 
n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , 
n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , 
n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , 
n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , 
n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , 
n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , 
n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , 
n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , 
n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , 
n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , 
n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , 
n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , 
n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , 
n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , 
n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , 
n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , 
n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , 
n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , 
n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , 
n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , 
n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , 
n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , 
n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , 
n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , 
n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , 
n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , 
n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , 
n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , 
n32091 , n32092 , n32093 , n32094 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , 
n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , 
n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , 
n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , 
n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , 
n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , 
n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , 
n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , 
n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , 
n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , 
n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , 
n32202 , n32203 , n32204 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , 
n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , 
n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , 
n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , 
n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , 
n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , 
n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , 
n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , 
n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , 
n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , 
n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , 
n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , 
n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32330 , n32331 , n32332 , n32333 , 
n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , 
n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , 
n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , 
n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , 
n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , 
n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , 
n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , 
n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , 
n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , 
n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , 
n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , 
n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , 
n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , 
n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , 
n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , 
n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , 
n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , 
n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , 
n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , 
n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , 
n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , 
n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , 
n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , 
n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , 
n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , 
n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , 
n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , 
n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , 
n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , 
n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , 
n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , 
n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , 
n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , 
n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32676 , 
n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , 
n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , 
n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , 
n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32716 , n32717 , n32718 , 
n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , 
n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , 
n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , 
n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , 
n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , 
n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , 
n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , 
n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , 
n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , 
n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , 
n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , 
n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , 
n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , 
n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32858 , n32859 , 
n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , 
n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , 
n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , 
n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , 
n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , 
n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , 
n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , 
n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , 
n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , 
n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , 
n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , 
n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , 
n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , 
n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , 
n33000 , n33001 , n33002 , n33003 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , 
n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , 
n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , 
n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , 
n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , 
n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , 
n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , 
n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , 
n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , 
n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , 
n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , 
n33112 , n33113 , n33114 , n33115 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , 
n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , 
n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , 
n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , 
n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , 
n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , 
n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , 
n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , 
n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , 
n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , 
n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , 
n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , 
n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , 
n33243 , n33244 , n33245 , n33246 , n33247 , n33249 , n33250 , n33251 , n33252 , n33253 , 
n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , 
n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , 
n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , 
n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , 
n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , 
n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , 
n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , 
n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , 
n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , 
n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , 
n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , 
n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , 
n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , 
n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , 
n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , 
n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , 
n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , 
n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , 
n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , 
n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , 
n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , 
n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , 
n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , 
n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , 
n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , 
n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , 
n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , 
n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , 
n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , 
n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , 
n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , 
n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , 
n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , 
n33585 , n33586 , n33587 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , 
n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , 
n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , 
n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , 
n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , 
n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , 
n33646 , n33647 , n33648 , n33649 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , 
n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , 
n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , 
n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , 
n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , 
n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , 
n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , 
n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , 
n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , 
n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , 
n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , 
n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , 
n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , 
n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , 
n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , 
n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , 
n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , 
n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , 
n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , 
n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , 
n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , 
n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , 
n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , 
n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , 
n33887 , n33888 , n33889 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , 
n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , 
n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , 
n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , 
n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , 
n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , 
n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , 
n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , 
n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , 
n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , 
n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , 
n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , 
n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , 
n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , 
n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , 
n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , 
n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , 
n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , 
n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , 
n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , 
n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , 
n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , 
n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , 
n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , 
n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , 
n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , 
n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , 
n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , 
n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , 
n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , 
n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , 
n34198 , n34199 , n34200 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , 
n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , 
n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , 
n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , 
n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34246 , n34247 , n34248 , n34249 , 
n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , 
n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34270 , 
n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , 
n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , 
n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , 
n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , 
n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , 
n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , 
n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , 
n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , 
n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , 
n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , 
n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , 
n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , 
n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , 
n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , 
n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , 
n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , 
n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , 
n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , 
n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , 
n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , 
n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , 
n34481 , n34482 , n34483 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , 
n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , 
n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , 
n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , 
n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , 
n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , 
n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , 
n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , 
n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34572 , 
n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , 
n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , 
n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , 
n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , 
n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , 
n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , 
n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , 
n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , 
n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , 
n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , 
n34673 , n34674 , n34675 , n34676 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , 
n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , 
n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , 
n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , 
n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , 
n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , 
n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , 
n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , 
n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , 
n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , 
n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , 
n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , 
n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , 
n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , 
n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34821 , n34822 , n34823 , n34824 , 
n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , 
n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , 
n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , 
n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , 
n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , 
n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , 
n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , 
n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34904 , n34905 , 
n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , 
n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34924 , n34925 , n34926 , 
n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , 
n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , 
n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , 
n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , 
n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , 
n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , 
n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , 
n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , 
n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , 
n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , 
n35027 , n35028 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , 
n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , 
n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , 
n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , 
n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , 
n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , 
n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , 
n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , 
n35108 , n35109 , n35110 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , 
n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , 
n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , 
n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , 
n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , 
n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , 
n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , 
n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , 
n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , 
n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , 
n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , 
n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , 
n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , 
n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , 
n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , 
n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , 
n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , 
n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , 
n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , 
n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , 
n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , 
n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , 
n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , 
n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , 
n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , 
n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , 
n35369 , n35370 , n35371 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , 
n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , 
n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , 
n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , 
n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , 
n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , 
n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , 
n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , 
n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , 
n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , 
n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35480 , 
n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , 
n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , 
n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , 
n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , 
n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , 
n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , 
n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , 
n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , 
n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , 
n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , 
n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , 
n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , 
n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , 
n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35619 , n35620 , n35621 , 
n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , 
n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , 
n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , 
n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , 
n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , 
n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , 
n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , 
n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , 
n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , 
n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , 
n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , 
n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , 
n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , 
n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , 
n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , 
n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , 
n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , 
n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , 
n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , 
n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , 
n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , 
n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , 
n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , 
n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , 
n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , 
n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , 
n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , 
n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , 
n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , 
n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , 
n35922 , n35923 , n35925 , n35926 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , 
n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , 
n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35951 , n35952 , n35953 , n35954 , 
n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , 
n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , 
n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , 
n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , 
n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , 
n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , 
n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , 
n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , 
n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , 
n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , 
n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , 
n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , 
n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , 
n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 ;
    and g0 ( n34347 , n19596 , n12943 );
    or g1 ( n34076 , n25436 , n6705 );
    or g2 ( n23999 , n17918 , n27643 );
    or g3 ( n12475 , n30742 , n22313 );
    and g4 ( n28859 , n31904 , n14576 );
    or g5 ( n32279 , n29713 , n32989 );
    or g6 ( n31197 , n19272 , n25355 );
    and g7 ( n14617 , n11030 , n1292 );
    or g8 ( n34732 , n24627 , n4132 );
    xnor g9 ( n17219 , n2795 , n34801 );
    and g10 ( n18158 , n23141 , n7886 );
    nor g11 ( n13788 , n33717 , n13267 );
    nor g12 ( n14345 , n25602 , n5172 );
    buf g13 ( n34537 , n30877 );
    or g14 ( n14433 , n3946 , n15305 );
    or g15 ( n32599 , n6038 , n16919 );
    xnor g16 ( n15 , n35459 , n16747 );
    or g17 ( n21254 , n31215 , n3498 );
    or g18 ( n27047 , n13794 , n26089 );
    or g19 ( n29325 , n20244 , n18255 );
    xnor g20 ( n17637 , n1033 , n11772 );
    and g21 ( n19559 , n5786 , n912 );
    and g22 ( n23046 , n13756 , n30143 );
    or g23 ( n12325 , n3202 , n32135 );
    xnor g24 ( n14081 , n684 , n9658 );
    and g25 ( n481 , n13054 , n19408 );
    and g26 ( n16600 , n15423 , n1770 );
    and g27 ( n24468 , n18690 , n34893 );
    not g28 ( n34852 , n25392 );
    or g29 ( n16340 , n16065 , n25567 );
    or g30 ( n26923 , n24647 , n4996 );
    not g31 ( n9352 , n22980 );
    and g32 ( n6624 , n5325 , n24983 );
    and g33 ( n18353 , n4306 , n9662 );
    and g34 ( n8080 , n104 , n13530 );
    or g35 ( n8361 , n21648 , n27580 );
    and g36 ( n713 , n16828 , n7935 );
    not g37 ( n36048 , n9725 );
    xnor g38 ( n32705 , n4536 , n961 );
    or g39 ( n28537 , n3205 , n28397 );
    xnor g40 ( n9892 , n72 , n35468 );
    or g41 ( n32048 , n13858 , n3964 );
    or g42 ( n8458 , n34195 , n3634 );
    or g43 ( n30810 , n25668 , n3581 );
    or g44 ( n32977 , n13002 , n30555 );
    or g45 ( n22671 , n5945 , n30826 );
    or g46 ( n17289 , n24371 , n29163 );
    xnor g47 ( n24376 , n11656 , n891 );
    or g48 ( n28391 , n19476 , n16817 );
    nor g49 ( n15940 , n11166 , n20797 );
    or g50 ( n28409 , n29108 , n28574 );
    or g51 ( n25669 , n13194 , n17190 );
    and g52 ( n2037 , n33266 , n13968 );
    or g53 ( n14408 , n4962 , n33902 );
    and g54 ( n7472 , n30272 , n10406 );
    or g55 ( n21793 , n21247 , n19732 );
    or g56 ( n12265 , n12013 , n2769 );
    and g57 ( n32717 , n10578 , n33072 );
    and g58 ( n3240 , n28149 , n13297 );
    or g59 ( n26656 , n3529 , n34189 );
    or g60 ( n28936 , n4585 , n373 );
    xnor g61 ( n32544 , n22115 , n15782 );
    or g62 ( n23705 , n15657 , n28240 );
    nor g63 ( n34905 , n9658 , n19499 );
    or g64 ( n22562 , n23652 , n28160 );
    and g65 ( n32739 , n1838 , n28626 );
    xnor g66 ( n23807 , n163 , n35211 );
    not g67 ( n33379 , n29999 );
    or g68 ( n13921 , n761 , n6553 );
    and g69 ( n8043 , n25038 , n11777 );
    nor g70 ( n8559 , n4960 , n18871 );
    or g71 ( n22307 , n35012 , n16456 );
    or g72 ( n21191 , n33927 , n26365 );
    or g73 ( n11367 , n32106 , n7315 );
    xnor g74 ( n9191 , n16489 , n13451 );
    or g75 ( n21632 , n17568 , n28070 );
    and g76 ( n30334 , n11884 , n12978 );
    xnor g77 ( n18339 , n21022 , n18233 );
    not g78 ( n24647 , n31551 );
    and g79 ( n13610 , n24696 , n24383 );
    xnor g80 ( n20587 , n10951 , n24150 );
    nor g81 ( n17611 , n33541 , n12852 );
    xnor g82 ( n12028 , n35436 , n27152 );
    nor g83 ( n15288 , n16922 , n24422 );
    xnor g84 ( n19274 , n24121 , n17568 );
    xnor g85 ( n29891 , n2907 , n22834 );
    not g86 ( n27057 , n29659 );
    or g87 ( n29711 , n32139 , n2044 );
    or g88 ( n17993 , n19551 , n27158 );
    or g89 ( n12882 , n6762 , n1856 );
    and g90 ( n12612 , n31457 , n26740 );
    or g91 ( n28946 , n12324 , n23763 );
    and g92 ( n34874 , n7678 , n4061 );
    and g93 ( n5103 , n30690 , n17209 );
    or g94 ( n13352 , n10063 , n35840 );
    and g95 ( n4334 , n26993 , n29013 );
    or g96 ( n31654 , n34223 , n25366 );
    or g97 ( n17148 , n1330 , n14554 );
    not g98 ( n29460 , n21894 );
    or g99 ( n17036 , n4957 , n22316 );
    xnor g100 ( n25025 , n19186 , n10847 );
    xnor g101 ( n364 , n12237 , n15107 );
    xor g102 ( n21280 , n17891 , n14693 );
    and g103 ( n32866 , n5646 , n12182 );
    and g104 ( n12581 , n23523 , n3085 );
    and g105 ( n31239 , n10518 , n5649 );
    or g106 ( n20560 , n10429 , n4081 );
    and g107 ( n7921 , n8565 , n3460 );
    or g108 ( n30845 , n16922 , n5396 );
    xnor g109 ( n4380 , n10966 , n13797 );
    xnor g110 ( n27297 , n13349 , n1458 );
    or g111 ( n18987 , n20683 , n33155 );
    nor g112 ( n4327 , n147 , n17297 );
    or g113 ( n21628 , n25008 , n31786 );
    or g114 ( n2681 , n17378 , n20576 );
    or g115 ( n11352 , n24272 , n2251 );
    and g116 ( n10847 , n12865 , n2759 );
    buf g117 ( n13305 , n4354 );
    xnor g118 ( n1944 , n10761 , n7540 );
    or g119 ( n11299 , n32940 , n7861 );
    or g120 ( n272 , n7397 , n21494 );
    not g121 ( n5081 , n29801 );
    or g122 ( n7145 , n6898 , n585 );
    xnor g123 ( n10939 , n4346 , n32632 );
    and g124 ( n11927 , n23479 , n20657 );
    xnor g125 ( n30380 , n22153 , n16620 );
    and g126 ( n29529 , n5514 , n33318 );
    or g127 ( n32251 , n32095 , n1295 );
    or g128 ( n13652 , n29839 , n35169 );
    xnor g129 ( n17624 , n16467 , n16736 );
    not g130 ( n5560 , n30934 );
    or g131 ( n8744 , n9850 , n25392 );
    xnor g132 ( n25696 , n14977 , n14911 );
    not g133 ( n21786 , n15464 );
    or g134 ( n565 , n30180 , n29214 );
    or g135 ( n6476 , n421 , n32697 );
    and g136 ( n8970 , n14432 , n16968 );
    or g137 ( n10987 , n7408 , n35457 );
    not g138 ( n14745 , n20840 );
    or g139 ( n9610 , n16848 , n21210 );
    or g140 ( n12005 , n13345 , n24381 );
    and g141 ( n30357 , n31901 , n3105 );
    xnor g142 ( n20881 , n24539 , n4878 );
    xnor g143 ( n35059 , n16737 , n2531 );
    or g144 ( n26496 , n26315 , n27085 );
    and g145 ( n35282 , n34871 , n10274 );
    and g146 ( n19216 , n8331 , n17989 );
    and g147 ( n24919 , n13876 , n33775 );
    or g148 ( n13219 , n14883 , n2384 );
    xnor g149 ( n18341 , n13681 , n35927 );
    or g150 ( n33159 , n4599 , n5618 );
    and g151 ( n17487 , n27306 , n11327 );
    or g152 ( n22107 , n23762 , n4994 );
    or g153 ( n24516 , n17972 , n28291 );
    or g154 ( n31118 , n32857 , n2646 );
    and g155 ( n2010 , n20287 , n30503 );
    and g156 ( n23098 , n7904 , n1258 );
    and g157 ( n13747 , n16029 , n14638 );
    not g158 ( n21305 , n3205 );
    and g159 ( n16177 , n6671 , n19431 );
    xnor g160 ( n11378 , n2232 , n19551 );
    and g161 ( n31957 , n10126 , n22674 );
    nor g162 ( n21176 , n13031 , n35643 );
    and g163 ( n34591 , n28344 , n1991 );
    xnor g164 ( n1161 , n12191 , n34922 );
    and g165 ( n9141 , n15862 , n32870 );
    or g166 ( n22473 , n24371 , n4707 );
    xnor g167 ( n21538 , n27978 , n8432 );
    and g168 ( n32989 , n13946 , n3777 );
    xnor g169 ( n7565 , n12318 , n16620 );
    and g170 ( n31984 , n6522 , n18401 );
    xnor g171 ( n11551 , n10112 , n29839 );
    xnor g172 ( n31330 , n29361 , n573 );
    or g173 ( n14686 , n26821 , n2168 );
    and g174 ( n26287 , n34818 , n33903 );
    or g175 ( n133 , n31289 , n25139 );
    nor g176 ( n35297 , n2826 , n6151 );
    or g177 ( n29171 , n26001 , n21956 );
    xnor g178 ( n9426 , n863 , n15403 );
    or g179 ( n30625 , n19523 , n32309 );
    or g180 ( n33709 , n20017 , n3188 );
    xnor g181 ( n16664 , n15813 , n3222 );
    xnor g182 ( n20065 , n22621 , n4962 );
    xnor g183 ( n6541 , n25118 , n16073 );
    and g184 ( n9580 , n19508 , n25118 );
    or g185 ( n33514 , n10265 , n26411 );
    or g186 ( n17943 , n21533 , n1511 );
    or g187 ( n11847 , n2176 , n24710 );
    and g188 ( n34614 , n22683 , n6944 );
    or g189 ( n17452 , n10325 , n1763 );
    or g190 ( n13080 , n13298 , n14841 );
    and g191 ( n13056 , n25187 , n31561 );
    and g192 ( n900 , n29749 , n28673 );
    and g193 ( n28981 , n27173 , n14302 );
    and g194 ( n3778 , n7013 , n33667 );
    or g195 ( n27347 , n9793 , n13364 );
    or g196 ( n17833 , n31336 , n12950 );
    xnor g197 ( n25862 , n33138 , n3222 );
    and g198 ( n25350 , n15023 , n28204 );
    or g199 ( n11160 , n5096 , n16659 );
    and g200 ( n17288 , n29286 , n4502 );
    or g201 ( n18004 , n24371 , n16644 );
    or g202 ( n10193 , n15213 , n23209 );
    not g203 ( n3552 , n26604 );
    or g204 ( n29944 , n14270 , n10960 );
    xnor g205 ( n29029 , n34208 , n31832 );
    nor g206 ( n34110 , n27513 , n2132 );
    or g207 ( n1006 , n10894 , n28308 );
    or g208 ( n15907 , n6384 , n3437 );
    or g209 ( n12390 , n15454 , n28438 );
    xnor g210 ( n18162 , n35880 , n8210 );
    and g211 ( n2118 , n13534 , n9018 );
    and g212 ( n3964 , n34065 , n3684 );
    and g213 ( n26049 , n35367 , n2094 );
    xnor g214 ( n34037 , n19925 , n15515 );
    xnor g215 ( n6773 , n34246 , n8273 );
    xnor g216 ( n35773 , n21147 , n17568 );
    or g217 ( n8508 , n32095 , n30132 );
    not g218 ( n27514 , n10802 );
    not g219 ( n7081 , n15886 );
    and g220 ( n4929 , n8120 , n30055 );
    nor g221 ( n18656 , n29167 , n34117 );
    not g222 ( n22445 , n3805 );
    or g223 ( n29618 , n5335 , n26046 );
    and g224 ( n26580 , n2835 , n3452 );
    or g225 ( n35295 , n7056 , n11364 );
    or g226 ( n16299 , n23429 , n32777 );
    or g227 ( n30730 , n5287 , n34398 );
    xnor g228 ( n8243 , n18778 , n32289 );
    and g229 ( n26514 , n32582 , n9653 );
    xnor g230 ( n675 , n11296 , n26705 );
    or g231 ( n3200 , n13963 , n18373 );
    or g232 ( n16700 , n2218 , n30222 );
    or g233 ( n28025 , n17568 , n24953 );
    nor g234 ( n10979 , n35927 , n2684 );
    or g235 ( n4721 , n16620 , n32611 );
    not g236 ( n27667 , n18296 );
    xnor g237 ( n14482 , n28717 , n13262 );
    or g238 ( n25670 , n20794 , n8674 );
    xnor g239 ( n15956 , n24880 , n32199 );
    not g240 ( n1624 , n6653 );
    or g241 ( n1445 , n4072 , n29393 );
    and g242 ( n9553 , n6248 , n845 );
    and g243 ( n31182 , n31635 , n1872 );
    nor g244 ( n27143 , n25416 , n3501 );
    or g245 ( n12170 , n32857 , n21124 );
    or g246 ( n22762 , n25098 , n19939 );
    or g247 ( n5453 , n20169 , n920 );
    or g248 ( n28749 , n19915 , n25392 );
    or g249 ( n12471 , n16168 , n9832 );
    and g250 ( n21638 , n32706 , n8569 );
    or g251 ( n18789 , n13799 , n25744 );
    and g252 ( n25673 , n2594 , n5903 );
    xnor g253 ( n31169 , n1355 , n29848 );
    nor g254 ( n11392 , n29839 , n2733 );
    not g255 ( n446 , n7540 );
    nor g256 ( n10928 , n5736 , n19834 );
    and g257 ( n2769 , n16325 , n19670 );
    or g258 ( n4121 , n24248 , n2798 );
    and g259 ( n4196 , n12283 , n2891 );
    and g260 ( n13407 , n15622 , n16218 );
    nor g261 ( n29143 , n24286 , n29366 );
    or g262 ( n25791 , n18061 , n34971 );
    not g263 ( n29771 , n31559 );
    and g264 ( n6128 , n19482 , n12696 );
    xnor g265 ( n24322 , n3294 , n24213 );
    or g266 ( n11358 , n17568 , n21040 );
    and g267 ( n23722 , n7362 , n23995 );
    and g268 ( n10660 , n3606 , n18865 );
    or g269 ( n8880 , n34317 , n21691 );
    xnor g270 ( n15257 , n12848 , n21935 );
    xnor g271 ( n25757 , n25215 , n16620 );
    or g272 ( n892 , n5908 , n31333 );
    or g273 ( n13721 , n2879 , n15344 );
    or g274 ( n6536 , n11760 , n24000 );
    nor g275 ( n19305 , n9833 , n7448 );
    nor g276 ( n7337 , n7928 , n17177 );
    xnor g277 ( n15626 , n24623 , n2513 );
    or g278 ( n13388 , n12844 , n34537 );
    and g279 ( n34670 , n25497 , n19406 );
    and g280 ( n35465 , n4877 , n19847 );
    and g281 ( n1591 , n6284 , n12037 );
    and g282 ( n26926 , n20483 , n390 );
    or g283 ( n22670 , n6941 , n28225 );
    or g284 ( n25362 , n15403 , n21990 );
    nor g285 ( n14820 , n29011 , n13045 );
    and g286 ( n35841 , n2747 , n12310 );
    or g287 ( n8759 , n20273 , n17125 );
    and g288 ( n18208 , n15232 , n6346 );
    nor g289 ( n12638 , n25602 , n9820 );
    and g290 ( n19515 , n10904 , n16779 );
    or g291 ( n17989 , n3005 , n27447 );
    or g292 ( n21033 , n15150 , n27625 );
    nor g293 ( n6670 , n31559 , n33878 );
    xnor g294 ( n11910 , n12185 , n23211 );
    and g295 ( n28719 , n8061 , n22053 );
    nor g296 ( n31838 , n7631 , n15645 );
    or g297 ( n21948 , n11046 , n17415 );
    not g298 ( n35050 , n17885 );
    or g299 ( n2043 , n25801 , n23790 );
    or g300 ( n10505 , n14078 , n11601 );
    and g301 ( n580 , n14804 , n3079 );
    or g302 ( n10347 , n1950 , n25282 );
    and g303 ( n26851 , n6654 , n1382 );
    and g304 ( n31437 , n15355 , n21763 );
    and g305 ( n16169 , n19527 , n31259 );
    and g306 ( n7355 , n22436 , n13819 );
    xnor g307 ( n1694 , n12838 , n35324 );
    nor g308 ( n1806 , n32857 , n2167 );
    or g309 ( n24207 , n18310 , n23798 );
    not g310 ( n33279 , n22980 );
    xnor g311 ( n25978 , n6606 , n31799 );
    xnor g312 ( n3783 , n32536 , n22258 );
    and g313 ( n12039 , n9336 , n2172 );
    or g314 ( n8839 , n14456 , n12879 );
    or g315 ( n21257 , n28922 , n25397 );
    xor g316 ( n26763 , n24694 , n17967 );
    xnor g317 ( n19715 , n13148 , n32095 );
    buf g318 ( n1856 , n3805 );
    or g319 ( n17275 , n18564 , n32634 );
    xnor g320 ( n20995 , n10158 , n4960 );
    xnor g321 ( n34176 , n5908 , n31333 );
    xnor g322 ( n26704 , n35980 , n31175 );
    xnor g323 ( n10547 , n27995 , n34011 );
    or g324 ( n32333 , n3587 , n13307 );
    not g325 ( n11837 , n12096 );
    xnor g326 ( n20017 , n23432 , n20854 );
    xnor g327 ( n4391 , n21562 , n5287 );
    and g328 ( n29687 , n9581 , n15231 );
    or g329 ( n19381 , n19099 , n33435 );
    or g330 ( n15217 , n1288 , n11749 );
    or g331 ( n26170 , n7521 , n14854 );
    or g332 ( n12878 , n32095 , n35197 );
    not g333 ( n24555 , n2433 );
    or g334 ( n32783 , n1304 , n508 );
    or g335 ( n17048 , n21227 , n25447 );
    or g336 ( n23488 , n9720 , n17111 );
    or g337 ( n3062 , n16619 , n24696 );
    and g338 ( n20948 , n5603 , n13730 );
    xnor g339 ( n12414 , n29964 , n4495 );
    and g340 ( n22399 , n20005 , n16613 );
    or g341 ( n16942 , n31634 , n11295 );
    or g342 ( n15357 , n21567 , n36024 );
    and g343 ( n26621 , n8086 , n24787 );
    and g344 ( n11600 , n33599 , n4985 );
    and g345 ( n28329 , n17236 , n20128 );
    or g346 ( n9356 , n2325 , n22501 );
    not g347 ( n18798 , n22980 );
    xnor g348 ( n26493 , n27777 , n12069 );
    and g349 ( n30902 , n5847 , n7037 );
    and g350 ( n1643 , n23615 , n30653 );
    xnor g351 ( n14957 , n13803 , n23228 );
    or g352 ( n34308 , n5067 , n3649 );
    or g353 ( n22592 , n9757 , n24262 );
    nor g354 ( n11017 , n9793 , n31336 );
    or g355 ( n35263 , n11046 , n9961 );
    or g356 ( n12157 , n35614 , n28357 );
    or g357 ( n2153 , n32095 , n6790 );
    or g358 ( n34495 , n32036 , n24115 );
    xnor g359 ( n20334 , n19255 , n32584 );
    nor g360 ( n17058 , n30742 , n34883 );
    or g361 ( n654 , n31799 , n27195 );
    and g362 ( n15621 , n5969 , n33583 );
    not g363 ( n14097 , n22980 );
    xnor g364 ( n20972 , n19482 , n5287 );
    xnor g365 ( n832 , n15231 , n9581 );
    and g366 ( n35782 , n28481 , n9644 );
    not g367 ( n252 , n1154 );
    or g368 ( n9851 , n34986 , n19245 );
    or g369 ( n21617 , n22025 , n5752 );
    or g370 ( n9973 , n31087 , n20797 );
    and g371 ( n31781 , n14235 , n21505 );
    nor g372 ( n12130 , n31799 , n20090 );
    xnor g373 ( n4582 , n34052 , n21386 );
    and g374 ( n29639 , n9000 , n5055 );
    and g375 ( n7312 , n29530 , n23202 );
    and g376 ( n814 , n6587 , n1526 );
    or g377 ( n19913 , n26540 , n1474 );
    or g378 ( n15147 , n22399 , n24710 );
    not g379 ( n4348 , n30333 );
    or g380 ( n25614 , n29164 , n32959 );
    or g381 ( n10332 , n25097 , n3593 );
    and g382 ( n8074 , n19703 , n33336 );
    and g383 ( n28601 , n12985 , n9606 );
    xnor g384 ( n30199 , n5351 , n25602 );
    xnor g385 ( n1302 , n8716 , n31799 );
    or g386 ( n21542 , n8432 , n1421 );
    or g387 ( n12718 , n27773 , n21644 );
    not g388 ( n6366 , n16594 );
    nor g389 ( n14001 , n3222 , n5770 );
    not g390 ( n8084 , n31419 );
    and g391 ( n15066 , n1445 , n15879 );
    or g392 ( n9669 , n35777 , n17068 );
    and g393 ( n19440 , n23881 , n13977 );
    and g394 ( n14363 , n31716 , n9304 );
    or g395 ( n21274 , n13277 , n25061 );
    nor g396 ( n10825 , n11046 , n9612 );
    or g397 ( n26420 , n3174 , n11712 );
    and g398 ( n25795 , n16130 , n12264 );
    and g399 ( n34585 , n25704 , n34453 );
    and g400 ( n11338 , n35835 , n28235 );
    or g401 ( n15591 , n22013 , n16961 );
    xnor g402 ( n28340 , n10647 , n25602 );
    and g403 ( n32160 , n11302 , n29281 );
    or g404 ( n29970 , n32726 , n6802 );
    or g405 ( n35368 , n25198 , n11177 );
    or g406 ( n19482 , n7882 , n21887 );
    and g407 ( n6233 , n14925 , n22976 );
    or g408 ( n11799 , n24324 , n19105 );
    not g409 ( n20379 , n2029 );
    xnor g410 ( n32656 , n35282 , n3481 );
    and g411 ( n29231 , n186 , n32213 );
    xnor g412 ( n24600 , n12355 , n33683 );
    and g413 ( n11808 , n34489 , n12983 );
    or g414 ( n16614 , n21261 , n4439 );
    xnor g415 ( n15858 , n12685 , n15942 );
    xnor g416 ( n33268 , n18334 , n32095 );
    and g417 ( n24112 , n33202 , n28140 );
    xnor g418 ( n19360 , n12253 , n28580 );
    or g419 ( n903 , n27291 , n169 );
    and g420 ( n6215 , n3558 , n5448 );
    xnor g421 ( n3930 , n12286 , n3222 );
    not g422 ( n3593 , n8746 );
    and g423 ( n13965 , n28316 , n35341 );
    or g424 ( n31144 , n35347 , n25594 );
    or g425 ( n28437 , n10951 , n24150 );
    or g426 ( n2910 , n17344 , n21315 );
    nor g427 ( n17191 , n8343 , n2458 );
    or g428 ( n32430 , n11455 , n20492 );
    and g429 ( n17152 , n22727 , n16753 );
    and g430 ( n16915 , n21768 , n27842 );
    xnor g431 ( n12695 , n33268 , n2778 );
    xnor g432 ( n36069 , n17950 , n2323 );
    or g433 ( n22436 , n30943 , n35046 );
    xnor g434 ( n16517 , n15832 , n35265 );
    and g435 ( n23852 , n21383 , n16588 );
    and g436 ( n16930 , n30388 , n19759 );
    xnor g437 ( n10071 , n27992 , n8071 );
    and g438 ( n21732 , n26496 , n23664 );
    or g439 ( n6687 , n21114 , n21616 );
    or g440 ( n15694 , n1749 , n32570 );
    or g441 ( n22806 , n11636 , n13341 );
    or g442 ( n36031 , n1175 , n6649 );
    or g443 ( n2142 , n8088 , n20797 );
    and g444 ( n15151 , n16535 , n27471 );
    and g445 ( n22177 , n24705 , n34998 );
    not g446 ( n12098 , n30865 );
    and g447 ( n214 , n21033 , n26494 );
    and g448 ( n4072 , n1008 , n28821 );
    and g449 ( n32443 , n16764 , n19873 );
    or g450 ( n22595 , n29037 , n28123 );
    or g451 ( n9537 , n7972 , n24479 );
    xnor g452 ( n23114 , n23612 , n4998 );
    buf g453 ( n8637 , n4526 );
    xnor g454 ( n4396 , n35732 , n4960 );
    or g455 ( n15348 , n29884 , n19145 );
    or g456 ( n12737 , n34159 , n4912 );
    nor g457 ( n12520 , n14106 , n6548 );
    xnor g458 ( n698 , n28560 , n30451 );
    not g459 ( n9257 , n32803 );
    or g460 ( n13150 , n18558 , n5868 );
    and g461 ( n25422 , n33378 , n7833 );
    and g462 ( n21687 , n8867 , n6367 );
    or g463 ( n17239 , n4869 , n31354 );
    xnor g464 ( n19777 , n7063 , n830 );
    or g465 ( n32956 , n7049 , n21042 );
    or g466 ( n2951 , n17180 , n6374 );
    or g467 ( n25709 , n3618 , n6950 );
    and g468 ( n8062 , n7044 , n20361 );
    xnor g469 ( n8409 , n14541 , n18588 );
    and g470 ( n29823 , n17147 , n23732 );
    or g471 ( n19075 , n26206 , n24672 );
    xnor g472 ( n4504 , n34383 , n32968 );
    and g473 ( n31572 , n17154 , n8414 );
    or g474 ( n10551 , n18336 , n14072 );
    xnor g475 ( n3186 , n35257 , n25837 );
    or g476 ( n5311 , n31686 , n23046 );
    and g477 ( n30983 , n24175 , n22981 );
    not g478 ( n29850 , n22980 );
    and g479 ( n4712 , n4203 , n25260 );
    or g480 ( n22098 , n94 , n3634 );
    or g481 ( n20989 , n25602 , n14291 );
    not g482 ( n18475 , n27291 );
    nor g483 ( n30302 , n30742 , n29009 );
    or g484 ( n12620 , n15464 , n103 );
    or g485 ( n5511 , n28125 , n35043 );
    and g486 ( n28315 , n7099 , n25290 );
    xnor g487 ( n11944 , n18377 , n32897 );
    and g488 ( n3338 , n11748 , n2033 );
    and g489 ( n8965 , n11219 , n16590 );
    and g490 ( n29987 , n12198 , n19959 );
    xnor g491 ( n28033 , n42 , n21256 );
    or g492 ( n28754 , n15578 , n7375 );
    nor g493 ( n34170 , n11190 , n1656 );
    and g494 ( n35979 , n3474 , n28979 );
    not g495 ( n844 , n17952 );
    and g496 ( n26306 , n27700 , n12988 );
    or g497 ( n33247 , n27473 , n27053 );
    xnor g498 ( n21003 , n8712 , n21486 );
    xnor g499 ( n17875 , n33753 , n35927 );
    xnor g500 ( n672 , n19302 , n5516 );
    or g501 ( n26791 , n17479 , n854 );
    or g502 ( n23680 , n28443 , n27728 );
    xnor g503 ( n35167 , n26448 , n29607 );
    or g504 ( n25325 , n29839 , n11569 );
    and g505 ( n15675 , n3022 , n20123 );
    not g506 ( n6831 , n13568 );
    or g507 ( n11097 , n13925 , n10264 );
    xnor g508 ( n33432 , n14765 , n7122 );
    or g509 ( n25959 , n18156 , n27743 );
    or g510 ( n15337 , n26136 , n23521 );
    and g511 ( n19867 , n7770 , n34828 );
    not g512 ( n1454 , n30732 );
    xnor g513 ( n26410 , n26550 , n30456 );
    or g514 ( n9422 , n12080 , n11921 );
    or g515 ( n13532 , n32715 , n23013 );
    not g516 ( n11755 , n26112 );
    or g517 ( n21663 , n35787 , n23829 );
    and g518 ( n12055 , n2424 , n32990 );
    or g519 ( n10652 , n4980 , n1796 );
    and g520 ( n18231 , n19780 , n2526 );
    or g521 ( n1432 , n21148 , n578 );
    or g522 ( n26123 , n2451 , n13015 );
    or g523 ( n1036 , n8085 , n21042 );
    nor g524 ( n13635 , n381 , n24213 );
    not g525 ( n34181 , n3281 );
    and g526 ( n448 , n26490 , n33922 );
    or g527 ( n10980 , n11685 , n16326 );
    or g528 ( n567 , n13336 , n29913 );
    xnor g529 ( n23262 , n21721 , n34154 );
    or g530 ( n24966 , n25376 , n581 );
    or g531 ( n27134 , n4962 , n10596 );
    xnor g532 ( n23314 , n4840 , n31559 );
    and g533 ( n24801 , n8166 , n35488 );
    or g534 ( n2553 , n3696 , n22946 );
    xnor g535 ( n14078 , n18906 , n26290 );
    or g536 ( n9425 , n17885 , n24489 );
    and g537 ( n30107 , n35011 , n27935 );
    nor g538 ( n32503 , n1234 , n28669 );
    or g539 ( n35781 , n24598 , n26002 );
    and g540 ( n18265 , n2279 , n27522 );
    buf g541 ( n30519 , n24307 );
    xnor g542 ( n9001 , n16857 , n15064 );
    and g543 ( n21237 , n31545 , n4721 );
    and g544 ( n409 , n30782 , n32652 );
    or g545 ( n15221 , n11323 , n18111 );
    or g546 ( n8799 , n17737 , n19258 );
    or g547 ( n34282 , n15277 , n4914 );
    xnor g548 ( n24276 , n89 , n26979 );
    and g549 ( n18395 , n23016 , n28150 );
    or g550 ( n23289 , n28011 , n25036 );
    and g551 ( n11478 , n6253 , n9638 );
    xnor g552 ( n30710 , n35717 , n15464 );
    and g553 ( n4827 , n22642 , n3189 );
    and g554 ( n35097 , n8894 , n6697 );
    xnor g555 ( n35163 , n27211 , n31289 );
    xnor g556 ( n15320 , n34475 , n29461 );
    xnor g557 ( n10333 , n23322 , n4288 );
    or g558 ( n9300 , n22137 , n139 );
    or g559 ( n23584 , n28139 , n20308 );
    and g560 ( n28835 , n23686 , n26088 );
    and g561 ( n32843 , n33095 , n23303 );
    or g562 ( n16134 , n16922 , n20516 );
    xnor g563 ( n13583 , n23309 , n17438 );
    nor g564 ( n31250 , n17659 , n18169 );
    or g565 ( n35133 , n2921 , n30095 );
    xnor g566 ( n3943 , n18094 , n17167 );
    or g567 ( n5672 , n14101 , n31554 );
    or g568 ( n14091 , n15559 , n25831 );
    xnor g569 ( n28220 , n29807 , n19391 );
    xnor g570 ( n19894 , n11172 , n30917 );
    and g571 ( n7282 , n8856 , n12706 );
    or g572 ( n8014 , n20237 , n31627 );
    xnor g573 ( n17571 , n19948 , n12775 );
    nor g574 ( n24652 , n7540 , n4109 );
    nor g575 ( n24162 , n24371 , n21142 );
    xnor g576 ( n31298 , n31040 , n34902 );
    and g577 ( n25717 , n24976 , n7358 );
    and g578 ( n16528 , n35035 , n7790 );
    or g579 ( n20471 , n18043 , n30204 );
    or g580 ( n9845 , n6361 , n557 );
    not g581 ( n18839 , n27277 );
    buf g582 ( n14554 , n5724 );
    xor g583 ( n30214 , n5377 , n33702 );
    xnor g584 ( n15282 , n9564 , n23707 );
    and g585 ( n11684 , n31871 , n5494 );
    or g586 ( n5305 , n12127 , n128 );
    or g587 ( n26837 , n15197 , n26336 );
    and g588 ( n27476 , n28897 , n10613 );
    or g589 ( n35563 , n31799 , n24810 );
    and g590 ( n7907 , n21053 , n31367 );
    xnor g591 ( n17343 , n13438 , n27420 );
    or g592 ( n15741 , n13437 , n21868 );
    or g593 ( n24238 , n22866 , n31321 );
    or g594 ( n12255 , n14966 , n5926 );
    xnor g595 ( n24875 , n29202 , n753 );
    and g596 ( n25569 , n4481 , n20397 );
    or g597 ( n31828 , n17031 , n2131 );
    xnor g598 ( n3256 , n25852 , n18993 );
    or g599 ( n15434 , n17899 , n33435 );
    nor g600 ( n5617 , n32715 , n10688 );
    or g601 ( n24975 , n32214 , n19490 );
    or g602 ( n4139 , n16620 , n652 );
    or g603 ( n3418 , n4288 , n18610 );
    and g604 ( n17223 , n15384 , n5035 );
    or g605 ( n16251 , n32095 , n456 );
    or g606 ( n13571 , n7002 , n2457 );
    or g607 ( n13356 , n18231 , n3437 );
    or g608 ( n7561 , n25024 , n14746 );
    or g609 ( n16393 , n27226 , n25836 );
    nor g610 ( n21155 , n31641 , n17753 );
    or g611 ( n17454 , n30578 , n21224 );
    xnor g612 ( n2752 , n33245 , n7712 );
    and g613 ( n3502 , n8281 , n4466 );
    or g614 ( n10865 , n5915 , n20911 );
    or g615 ( n15152 , n21639 , n26480 );
    xnor g616 ( n23581 , n18270 , n533 );
    buf g617 ( n29366 , n6548 );
    and g618 ( n14336 , n15640 , n22630 );
    or g619 ( n5047 , n9417 , n13210 );
    xnor g620 ( n572 , n1848 , n12391 );
    or g621 ( n15071 , n863 , n27053 );
    and g622 ( n31392 , n23635 , n13190 );
    nor g623 ( n16068 , n830 , n29059 );
    xnor g624 ( n19545 , n26729 , n16922 );
    or g625 ( n16511 , n17568 , n30761 );
    or g626 ( n16902 , n6584 , n18972 );
    and g627 ( n15333 , n17199 , n9857 );
    not g628 ( n16302 , n27337 );
    xnor g629 ( n11730 , n29103 , n10894 );
    xnor g630 ( n19424 , n15590 , n8781 );
    or g631 ( n29916 , n4940 , n28257 );
    or g632 ( n21571 , n9640 , n28248 );
    and g633 ( n25018 , n28620 , n12371 );
    or g634 ( n17841 , n10894 , n28720 );
    and g635 ( n20931 , n23463 , n5796 );
    xnor g636 ( n18897 , n3365 , n14049 );
    and g637 ( n16461 , n19111 , n25949 );
    xnor g638 ( n17749 , n9919 , n31740 );
    buf g639 ( n1763 , n21579 );
    and g640 ( n22334 , n5004 , n28244 );
    or g641 ( n26507 , n17682 , n3437 );
    or g642 ( n24726 , n10210 , n26728 );
    nor g643 ( n31319 , n2781 , n28283 );
    not g644 ( n17396 , n10191 );
    or g645 ( n2948 , n29309 , n15536 );
    xnor g646 ( n26548 , n25561 , n26393 );
    not g647 ( n21553 , n3205 );
    nor g648 ( n7460 , n16620 , n27571 );
    or g649 ( n15441 , n28901 , n19464 );
    not g650 ( n5694 , n27263 );
    and g651 ( n21774 , n28424 , n5175 );
    or g652 ( n3083 , n35088 , n27225 );
    xnor g653 ( n14965 , n6755 , n16773 );
    xnor g654 ( n32486 , n679 , n14297 );
    nor g655 ( n32984 , n22162 , n24027 );
    or g656 ( n24029 , n11143 , n4081 );
    and g657 ( n12829 , n34222 , n26383 );
    and g658 ( n17554 , n30213 , n3060 );
    xnor g659 ( n2226 , n21464 , n16135 );
    xnor g660 ( n32844 , n1093 , n4878 );
    nor g661 ( n6617 , n35321 , n36057 );
    and g662 ( n12693 , n28522 , n26702 );
    or g663 ( n22938 , n15886 , n31069 );
    nor g664 ( n13419 , n16135 , n11892 );
    or g665 ( n25739 , n24654 , n2823 );
    and g666 ( n14281 , n25132 , n586 );
    or g667 ( n29773 , n21214 , n17598 );
    or g668 ( n22744 , n23807 , n31549 );
    or g669 ( n27569 , n30277 , n28985 );
    nor g670 ( n12022 , n17485 , n34991 );
    buf g671 ( n30287 , n32837 );
    xnor g672 ( n28415 , n19715 , n3961 );
    xnor g673 ( n30907 , n29859 , n6537 );
    or g674 ( n6149 , n9790 , n9675 );
    or g675 ( n16520 , n7605 , n28680 );
    or g676 ( n16151 , n5287 , n17984 );
    and g677 ( n29686 , n9569 , n24369 );
    nor g678 ( n18349 , n9980 , n13352 );
    or g679 ( n7492 , n18257 , n35757 );
    or g680 ( n2087 , n18132 , n35660 );
    or g681 ( n30909 , n11455 , n6976 );
    nor g682 ( n15216 , n27870 , n1176 );
    or g683 ( n13741 , n3624 , n13850 );
    nor g684 ( n2877 , n22376 , n15835 );
    and g685 ( n24545 , n14913 , n15664 );
    or g686 ( n7099 , n34710 , n31067 );
    and g687 ( n30865 , n28274 , n3304 );
    xnor g688 ( n34637 , n34770 , n1910 );
    and g689 ( n10008 , n12232 , n24845 );
    or g690 ( n23673 , n31745 , n14754 );
    and g691 ( n4482 , n20777 , n27244 );
    or g692 ( n7414 , n4387 , n31514 );
    or g693 ( n23866 , n24231 , n21210 );
    xnor g694 ( n2399 , n26978 , n33261 );
    or g695 ( n11256 , n15804 , n11833 );
    xnor g696 ( n14561 , n5888 , n14192 );
    or g697 ( n22781 , n14193 , n25915 );
    or g698 ( n4806 , n17166 , n27420 );
    not g699 ( n31604 , n9568 );
    or g700 ( n8055 , n28735 , n5094 );
    nor g701 ( n32657 , n2878 , n33157 );
    or g702 ( n20969 , n12491 , n27860 );
    or g703 ( n2163 , n18303 , n11532 );
    or g704 ( n24578 , n19790 , n11593 );
    nor g705 ( n18051 , n3946 , n24968 );
    or g706 ( n18295 , n32098 , n30732 );
    or g707 ( n7641 , n2370 , n25466 );
    xnor g708 ( n30473 , n13010 , n31799 );
    or g709 ( n2866 , n22909 , n24905 );
    or g710 ( n6030 , n29298 , n17125 );
    and g711 ( n23369 , n21848 , n19046 );
    or g712 ( n18996 , n9226 , n20228 );
    or g713 ( n2071 , n22291 , n18196 );
    and g714 ( n10688 , n25784 , n31196 );
    nor g715 ( n27956 , n15704 , n9439 );
    xnor g716 ( n7599 , n32368 , n715 );
    not g717 ( n9910 , n12507 );
    xnor g718 ( n6960 , n10604 , n29754 );
    or g719 ( n20650 , n18083 , n25421 );
    or g720 ( n618 , n31413 , n10412 );
    xnor g721 ( n27161 , n17031 , n2131 );
    or g722 ( n18122 , n17811 , n14684 );
    or g723 ( n32891 , n20072 , n2814 );
    not g724 ( n29407 , n19633 );
    or g725 ( n29961 , n7774 , n18075 );
    and g726 ( n22115 , n15322 , n5143 );
    or g727 ( n25011 , n17499 , n33034 );
    or g728 ( n27809 , n9312 , n29049 );
    xnor g729 ( n23155 , n10981 , n31964 );
    or g730 ( n7216 , n26539 , n908 );
    xnor g731 ( n26712 , n26519 , n15714 );
    and g732 ( n16463 , n11541 , n28674 );
    xnor g733 ( n12289 , n9576 , n35927 );
    xnor g734 ( n18823 , n8068 , n24955 );
    and g735 ( n21058 , n17242 , n11190 );
    xnor g736 ( n8715 , n10601 , n8376 );
    and g737 ( n7828 , n5858 , n6313 );
    and g738 ( n19874 , n11137 , n13614 );
    buf g739 ( n32697 , n18088 );
    or g740 ( n20757 , n21275 , n19113 );
    and g741 ( n25080 , n31918 , n26625 );
    or g742 ( n22468 , n8875 , n21579 );
    xnor g743 ( n20461 , n18867 , n6341 );
    xnor g744 ( n35669 , n24312 , n11046 );
    not g745 ( n7357 , n33272 );
    or g746 ( n6356 , n16972 , n14903 );
    and g747 ( n2714 , n34122 , n21035 );
    or g748 ( n19209 , n25964 , n7582 );
    or g749 ( n21493 , n14258 , n35941 );
    or g750 ( n16436 , n31245 , n20291 );
    or g751 ( n18444 , n7540 , n21758 );
    nor g752 ( n20680 , n22291 , n32170 );
    or g753 ( n2249 , n16889 , n33742 );
    or g754 ( n31252 , n9306 , n5590 );
    not g755 ( n9924 , n10678 );
    and g756 ( n13955 , n10113 , n18759 );
    or g757 ( n5133 , n19029 , n6075 );
    xnor g758 ( n18677 , n6272 , n29839 );
    or g759 ( n21895 , n24685 , n34087 );
    or g760 ( n921 , n31685 , n13320 );
    or g761 ( n6562 , n23047 , n7673 );
    xnor g762 ( n16780 , n23171 , n7303 );
    xnor g763 ( n6396 , n14299 , n7672 );
    xnor g764 ( n12459 , n13875 , n9214 );
    xnor g765 ( n5194 , n28996 , n19551 );
    and g766 ( n4557 , n32839 , n30103 );
    or g767 ( n19372 , n32715 , n13036 );
    xnor g768 ( n13913 , n11426 , n32857 );
    not g769 ( n2333 , n30688 );
    xnor g770 ( n2434 , n27049 , n16311 );
    nor g771 ( n2760 , n35927 , n10339 );
    not g772 ( n9135 , n4878 );
    or g773 ( n13226 , n20039 , n16898 );
    nor g774 ( n7237 , n20997 , n10267 );
    nor g775 ( n9312 , n4960 , n25558 );
    not g776 ( n2366 , n9361 );
    or g777 ( n19782 , n830 , n1403 );
    and g778 ( n21562 , n8427 , n3996 );
    and g779 ( n1650 , n18484 , n15464 );
    or g780 ( n31576 , n10194 , n3634 );
    xnor g781 ( n7939 , n7828 , n29839 );
    and g782 ( n27125 , n31963 , n34825 );
    nor g783 ( n16521 , n17751 , n29408 );
    nor g784 ( n31025 , n7741 , n18115 );
    xnor g785 ( n19908 , n21916 , n19551 );
    or g786 ( n23957 , n27472 , n27903 );
    and g787 ( n24517 , n5933 , n28880 );
    or g788 ( n22615 , n4778 , n22783 );
    not g789 ( n27878 , n17568 );
    and g790 ( n35693 , n34854 , n12248 );
    or g791 ( n31833 , n22197 , n13426 );
    or g792 ( n2362 , n22282 , n3438 );
    or g793 ( n16320 , n35030 , n15663 );
    xnor g794 ( n19112 , n13717 , n9793 );
    and g795 ( n2254 , n24723 , n22980 );
    and g796 ( n8469 , n22953 , n12696 );
    or g797 ( n6688 , n7540 , n29311 );
    or g798 ( n12900 , n3069 , n17204 );
    nor g799 ( n9275 , n34391 , n20579 );
    nor g800 ( n15028 , n8992 , n4508 );
    not g801 ( n9929 , n9489 );
    and g802 ( n21771 , n17472 , n34579 );
    or g803 ( n1263 , n32715 , n17622 );
    xnor g804 ( n33772 , n33681 , n7177 );
    or g805 ( n28657 , n4596 , n4829 );
    or g806 ( n29190 , n3222 , n35507 );
    or g807 ( n21065 , n26693 , n34923 );
    and g808 ( n14319 , n21697 , n30909 );
    or g809 ( n8645 , n34205 , n9930 );
    and g810 ( n13033 , n32771 , n4843 );
    buf g811 ( n25306 , n9297 );
    or g812 ( n11899 , n4841 , n19173 );
    not g813 ( n14070 , n27148 );
    nor g814 ( n10444 , n9789 , n11728 );
    and g815 ( n9053 , n666 , n14206 );
    and g816 ( n22824 , n2383 , n35601 );
    or g817 ( n5563 , n15795 , n16577 );
    and g818 ( n3296 , n19486 , n26363 );
    and g819 ( n2352 , n9742 , n19744 );
    or g820 ( n26422 , n13776 , n10140 );
    nor g821 ( n24198 , n25602 , n18946 );
    or g822 ( n25259 , n15464 , n12393 );
    xnor g823 ( n11814 , n7774 , n18075 );
    xnor g824 ( n28986 , n28335 , n8872 );
    and g825 ( n7901 , n32971 , n8135 );
    nor g826 ( n28739 , n30709 , n4661 );
    or g827 ( n24498 , n13114 , n19678 );
    or g828 ( n7241 , n692 , n22322 );
    and g829 ( n25588 , n1483 , n21737 );
    not g830 ( n415 , n7588 );
    xnor g831 ( n8374 , n14696 , n19551 );
    nor g832 ( n17922 , n4566 , n32730 );
    not g833 ( n23613 , n9032 );
    and g834 ( n5598 , n9521 , n17476 );
    nor g835 ( n16927 , n33457 , n30858 );
    and g836 ( n15796 , n26685 , n22290 );
    or g837 ( n25571 , n664 , n20576 );
    buf g838 ( n16594 , n14112 );
    or g839 ( n17377 , n25602 , n152 );
    or g840 ( n13404 , n18225 , n36000 );
    xnor g841 ( n17094 , n29767 , n21097 );
    or g842 ( n4812 , n33286 , n28248 );
    and g843 ( n7029 , n24638 , n16792 );
    or g844 ( n27958 , n10716 , n11805 );
    not g845 ( n27583 , n6288 );
    and g846 ( n16324 , n27256 , n31866 );
    and g847 ( n22823 , n32977 , n13536 );
    and g848 ( n19469 , n3131 , n939 );
    xnor g849 ( n18846 , n26364 , n28953 );
    xnor g850 ( n23940 , n1845 , n3946 );
    and g851 ( n1050 , n13827 , n24693 );
    or g852 ( n389 , n20587 , n5208 );
    and g853 ( n23213 , n7723 , n23998 );
    or g854 ( n17969 , n11329 , n8472 );
    and g855 ( n11690 , n34712 , n10666 );
    or g856 ( n16695 , n4389 , n5996 );
    xnor g857 ( n33708 , n11904 , n35848 );
    xnor g858 ( n7419 , n34205 , n4962 );
    or g859 ( n18860 , n2811 , n31927 );
    buf g860 ( n16223 , n27816 );
    nor g861 ( n3752 , n12413 , n31411 );
    xnor g862 ( n27025 , n25463 , n7540 );
    or g863 ( n27848 , n18569 , n28574 );
    xnor g864 ( n29675 , n25015 , n28236 );
    or g865 ( n20549 , n30328 , n4595 );
    and g866 ( n9920 , n2867 , n12040 );
    buf g867 ( n30708 , n24719 );
    or g868 ( n19096 , n33357 , n2712 );
    or g869 ( n11399 , n25068 , n27625 );
    not g870 ( n5818 , n29452 );
    nor g871 ( n28332 , n8129 , n35290 );
    or g872 ( n33078 , n34162 , n25447 );
    or g873 ( n19310 , n6844 , n11484 );
    not g874 ( n24382 , n32095 );
    and g875 ( n20838 , n6048 , n6942 );
    and g876 ( n29015 , n34020 , n29386 );
    or g877 ( n9170 , n25721 , n32959 );
    and g878 ( n17345 , n24335 , n27847 );
    or g879 ( n18543 , n1625 , n26931 );
    or g880 ( n11932 , n26194 , n33444 );
    or g881 ( n32817 , n13048 , n35822 );
    or g882 ( n5448 , n7326 , n25648 );
    or g883 ( n33002 , n1848 , n12391 );
    and g884 ( n16264 , n9464 , n10899 );
    or g885 ( n28499 , n12921 , n27728 );
    or g886 ( n15775 , n10869 , n6374 );
    or g887 ( n5731 , n20372 , n25019 );
    or g888 ( n2662 , n5033 , n8203 );
    not g889 ( n35625 , n30764 );
    or g890 ( n34157 , n29713 , n10087 );
    xnor g891 ( n5062 , n34805 , n24585 );
    xnor g892 ( n21520 , n14840 , n9658 );
    or g893 ( n13761 , n16353 , n8153 );
    or g894 ( n33846 , n22089 , n27625 );
    nor g895 ( n3369 , n2380 , n29373 );
    nor g896 ( n11933 , n18379 , n7365 );
    or g897 ( n17644 , n25602 , n26356 );
    xnor g898 ( n25383 , n17027 , n3222 );
    and g899 ( n31484 , n3935 , n9264 );
    xnor g900 ( n1813 , n4947 , n4206 );
    and g901 ( n32935 , n8896 , n35095 );
    or g902 ( n5659 , n27226 , n17422 );
    nor g903 ( n14335 , n24371 , n34132 );
    nor g904 ( n29698 , n8432 , n9446 );
    or g905 ( n35775 , n5754 , n26239 );
    and g906 ( n22791 , n24577 , n25881 );
    or g907 ( n9907 , n34965 , n21002 );
    and g908 ( n18163 , n26527 , n28923 );
    or g909 ( n470 , n23983 , n4081 );
    nor g910 ( n16987 , n32857 , n28011 );
    or g911 ( n2896 , n24371 , n33976 );
    or g912 ( n11226 , n9559 , n17604 );
    xnor g913 ( n10326 , n11373 , n35157 );
    or g914 ( n15309 , n7950 , n27747 );
    xnor g915 ( n23670 , n19139 , n5711 );
    xnor g916 ( n12075 , n16857 , n21869 );
    xnor g917 ( n25195 , n3258 , n33020 );
    xnor g918 ( n29428 , n17958 , n5477 );
    and g919 ( n14662 , n13443 , n1189 );
    or g920 ( n312 , n14327 , n4595 );
    and g921 ( n22429 , n35114 , n28741 );
    nor g922 ( n19167 , n22677 , n16348 );
    xnor g923 ( n25934 , n5044 , n22291 );
    and g924 ( n18366 , n20108 , n26045 );
    nor g925 ( n9503 , n16620 , n17091 );
    xnor g926 ( n34827 , n14200 , n10139 );
    or g927 ( n6048 , n23045 , n2384 );
    xnor g928 ( n14085 , n25821 , n4621 );
    or g929 ( n33627 , n29839 , n14885 );
    or g930 ( n24641 , n3222 , n23276 );
    and g931 ( n31702 , n14635 , n30273 );
    xnor g932 ( n11422 , n7028 , n23254 );
    xnor g933 ( n35955 , n32838 , n8432 );
    or g934 ( n9336 , n25370 , n11643 );
    nor g935 ( n14966 , n4962 , n12968 );
    xnor g936 ( n1790 , n3877 , n19733 );
    not g937 ( n22246 , n32795 );
    nor g938 ( n18458 , n16922 , n23864 );
    or g939 ( n11759 , n16922 , n3942 );
    and g940 ( n6802 , n22295 , n29396 );
    or g941 ( n14321 , n4758 , n9838 );
    xnor g942 ( n17663 , n13355 , n17294 );
    xnor g943 ( n30888 , n9183 , n4288 );
    or g944 ( n14456 , n3741 , n29850 );
    not g945 ( n2247 , n1996 );
    or g946 ( n5109 , n21707 , n11833 );
    and g947 ( n21332 , n19053 , n12224 );
    or g948 ( n4070 , n20419 , n32878 );
    or g949 ( n19842 , n27669 , n216 );
    and g950 ( n33197 , n9182 , n30291 );
    and g951 ( n32673 , n34696 , n13553 );
    or g952 ( n19637 , n12227 , n23471 );
    and g953 ( n21679 , n14091 , n27247 );
    xnor g954 ( n21688 , n19873 , n16764 );
    or g955 ( n10354 , n27748 , n33778 );
    xnor g956 ( n23963 , n8771 , n15464 );
    or g957 ( n710 , n16620 , n25375 );
    or g958 ( n19503 , n7111 , n16919 );
    and g959 ( n1215 , n8354 , n35062 );
    or g960 ( n1095 , n2483 , n20021 );
    or g961 ( n35106 , n18437 , n9731 );
    and g962 ( n3512 , n25724 , n22239 );
    and g963 ( n18927 , n15748 , n2280 );
    xnor g964 ( n13987 , n26348 , n26852 );
    xnor g965 ( n24127 , n26101 , n7858 );
    nor g966 ( n16663 , n23604 , n7265 );
    and g967 ( n12824 , n27481 , n14159 );
    or g968 ( n7782 , n3522 , n35164 );
    or g969 ( n17287 , n15289 , n27728 );
    or g970 ( n14948 , n26989 , n12254 );
    or g971 ( n3772 , n7684 , n12465 );
    and g972 ( n12464 , n22845 , n33836 );
    nor g973 ( n21000 , n15464 , n25987 );
    and g974 ( n28355 , n14453 , n21966 );
    and g975 ( n31381 , n18550 , n23831 );
    or g976 ( n20052 , n16387 , n12996 );
    xnor g977 ( n28520 , n3887 , n10709 );
    or g978 ( n2788 , n7540 , n28242 );
    and g979 ( n13672 , n23584 , n31166 );
    and g980 ( n6980 , n20456 , n25693 );
    or g981 ( n34683 , n35392 , n9930 );
    or g982 ( n30307 , n11455 , n28927 );
    or g983 ( n20212 , n35460 , n7354 );
    or g984 ( n3726 , n4962 , n14837 );
    or g985 ( n34459 , n6527 , n1715 );
    xnor g986 ( n28781 , n13878 , n32857 );
    xnor g987 ( n7416 , n2230 , n17568 );
    or g988 ( n11634 , n22262 , n33505 );
    or g989 ( n7810 , n11244 , n9081 );
    and g990 ( n11929 , n23905 , n4031 );
    or g991 ( n14261 , n24855 , n16459 );
    or g992 ( n18184 , n26386 , n5868 );
    xnor g993 ( n34596 , n1487 , n10381 );
    or g994 ( n18166 , n9658 , n8498 );
    nor g995 ( n22555 , n31559 , n24698 );
    xnor g996 ( n11049 , n10878 , n5335 );
    or g997 ( n4040 , n6431 , n11750 );
    xnor g998 ( n2899 , n18196 , n22291 );
    and g999 ( n6012 , n2968 , n32421 );
    and g1000 ( n5648 , n16136 , n22956 );
    or g1001 ( n9468 , n31056 , n28962 );
    and g1002 ( n25536 , n33846 , n15815 );
    xnor g1003 ( n16575 , n30233 , n6383 );
    or g1004 ( n25785 , n33295 , n22079 );
    or g1005 ( n1136 , n31072 , n33416 );
    xnor g1006 ( n23189 , n7027 , n18985 );
    and g1007 ( n28857 , n5492 , n24020 );
    not g1008 ( n18873 , n4878 );
    or g1009 ( n22825 , n19551 , n29942 );
    and g1010 ( n19115 , n27241 , n17867 );
    xnor g1011 ( n25192 , n24520 , n12705 );
    or g1012 ( n15685 , n14762 , n316 );
    not g1013 ( n12659 , n23887 );
    or g1014 ( n17994 , n33176 , n8203 );
    and g1015 ( n1734 , n6669 , n19488 );
    or g1016 ( n4256 , n12488 , n7553 );
    not g1017 ( n30555 , n16299 );
    or g1018 ( n27752 , n4878 , n14883 );
    or g1019 ( n1058 , n27309 , n25255 );
    xnor g1020 ( n3975 , n28550 , n11190 );
    and g1021 ( n498 , n5656 , n15058 );
    xnor g1022 ( n34415 , n18594 , n2549 );
    or g1023 ( n5843 , n15292 , n34600 );
    xnor g1024 ( n922 , n247 , n32095 );
    or g1025 ( n31313 , n17114 , n22589 );
    nor g1026 ( n27040 , n18513 , n813 );
    not g1027 ( n270 , n27226 );
    or g1028 ( n9381 , n358 , n18811 );
    buf g1029 ( n8924 , n21691 );
    nor g1030 ( n35123 , n32857 , n26609 );
    and g1031 ( n8187 , n29180 , n2850 );
    xnor g1032 ( n33188 , n33183 , n34621 );
    or g1033 ( n1398 , n5287 , n21884 );
    and g1034 ( n20032 , n1136 , n11793 );
    xnor g1035 ( n18549 , n25731 , n24716 );
    or g1036 ( n27797 , n16176 , n151 );
    or g1037 ( n3079 , n20869 , n9601 );
    and g1038 ( n10339 , n3150 , n1116 );
    and g1039 ( n14840 , n17036 , n22900 );
    and g1040 ( n32170 , n17833 , n22288 );
    or g1041 ( n21053 , n22649 , n25392 );
    or g1042 ( n29506 , n15692 , n28248 );
    or g1043 ( n2925 , n24332 , n14489 );
    and g1044 ( n19430 , n23159 , n29067 );
    or g1045 ( n33855 , n30638 , n2119 );
    xnor g1046 ( n21068 , n26643 , n32095 );
    and g1047 ( n25878 , n35636 , n2498 );
    or g1048 ( n17019 , n30967 , n7647 );
    nor g1049 ( n5685 , n16620 , n14537 );
    or g1050 ( n30011 , n2521 , n12996 );
    or g1051 ( n33566 , n16620 , n14211 );
    or g1052 ( n8520 , n29090 , n35944 );
    or g1053 ( n21818 , n16709 , n19748 );
    xnor g1054 ( n15617 , n1244 , n32095 );
    not g1055 ( n22449 , n29469 );
    xnor g1056 ( n29202 , n22236 , n4878 );
    and g1057 ( n12057 , n18740 , n25726 );
    xnor g1058 ( n17193 , n4841 , n1700 );
    not g1059 ( n115 , n22471 );
    and g1060 ( n17498 , n33356 , n33055 );
    or g1061 ( n15092 , n7895 , n16919 );
    or g1062 ( n31085 , n31747 , n34660 );
    and g1063 ( n15641 , n22235 , n27772 );
    or g1064 ( n30196 , n4904 , n20143 );
    or g1065 ( n3330 , n32095 , n27472 );
    or g1066 ( n19713 , n24682 , n17861 );
    xnor g1067 ( n28534 , n29433 , n30048 );
    or g1068 ( n3474 , n33591 , n35986 );
    or g1069 ( n21515 , n10306 , n2712 );
    or g1070 ( n3894 , n23604 , n29225 );
    or g1071 ( n28024 , n11926 , n15138 );
    or g1072 ( n31849 , n25613 , n36000 );
    and g1073 ( n11254 , n2041 , n11902 );
    nor g1074 ( n16689 , n6763 , n21955 );
    or g1075 ( n25818 , n19723 , n3842 );
    xnor g1076 ( n22373 , n25612 , n4758 );
    not g1077 ( n34094 , n13374 );
    or g1078 ( n6444 , n851 , n29953 );
    or g1079 ( n2067 , n7079 , n3235 );
    or g1080 ( n22844 , n23795 , n12034 );
    or g1081 ( n14731 , n19378 , n8203 );
    or g1082 ( n26322 , n7875 , n1763 );
    not g1083 ( n7803 , n12235 );
    or g1084 ( n4544 , n7538 , n4823 );
    or g1085 ( n25925 , n830 , n33529 );
    xnor g1086 ( n16832 , n24731 , n23554 );
    xnor g1087 ( n25244 , n23946 , n6498 );
    buf g1088 ( n17829 , n29592 );
    or g1089 ( n27281 , n594 , n34560 );
    and g1090 ( n32198 , n19862 , n34354 );
    or g1091 ( n25827 , n23604 , n22774 );
    not g1092 ( n18708 , n15403 );
    or g1093 ( n2716 , n20157 , n7897 );
    not g1094 ( n5991 , n30858 );
    xnor g1095 ( n26028 , n16143 , n32510 );
    and g1096 ( n26398 , n15315 , n10501 );
    and g1097 ( n33261 , n22820 , n32347 );
    or g1098 ( n17842 , n6845 , n22998 );
    or g1099 ( n34731 , n25945 , n30514 );
    and g1100 ( n29241 , n34750 , n20088 );
    and g1101 ( n30028 , n18188 , n20658 );
    and g1102 ( n3219 , n26873 , n5939 );
    xnor g1103 ( n18202 , n26321 , n24371 );
    and g1104 ( n14856 , n4083 , n20129 );
    xnor g1105 ( n9117 , n17188 , n24586 );
    xnor g1106 ( n17427 , n1578 , n5067 );
    nor g1107 ( n25075 , n10221 , n27954 );
    and g1108 ( n1252 , n20254 , n26986 );
    xnor g1109 ( n13893 , n10843 , n22144 );
    and g1110 ( n4905 , n9156 , n7526 );
    or g1111 ( n5046 , n17568 , n28594 );
    nor g1112 ( n16005 , n4225 , n17135 );
    xnor g1113 ( n35247 , n28982 , n6086 );
    and g1114 ( n27624 , n30021 , n7257 );
    or g1115 ( n5180 , n7407 , n15030 );
    or g1116 ( n34380 , n7585 , n22062 );
    and g1117 ( n10072 , n12362 , n22980 );
    nor g1118 ( n29135 , n19551 , n14533 );
    xnor g1119 ( n20574 , n14802 , n30769 );
    xnor g1120 ( n230 , n2035 , n16097 );
    or g1121 ( n13214 , n14229 , n27203 );
    or g1122 ( n32380 , n7074 , n2955 );
    or g1123 ( n20933 , n5034 , n25295 );
    xnor g1124 ( n34983 , n31133 , n17568 );
    xnor g1125 ( n15863 , n23723 , n14778 );
    and g1126 ( n759 , n22662 , n12982 );
    xnor g1127 ( n21285 , n996 , n24371 );
    or g1128 ( n26650 , n9952 , n19464 );
    xnor g1129 ( n22425 , n35596 , n9877 );
    nor g1130 ( n23192 , n8007 , n7042 );
    nor g1131 ( n19863 , n33144 , n12569 );
    xnor g1132 ( n1422 , n4073 , n3502 );
    or g1133 ( n18990 , n33268 , n2778 );
    not g1134 ( n32928 , n6613 );
    xnor g1135 ( n31357 , n22594 , n2438 );
    or g1136 ( n13697 , n5585 , n27704 );
    and g1137 ( n6937 , n21265 , n14020 );
    xnor g1138 ( n8147 , n5299 , n22291 );
    or g1139 ( n3434 , n14428 , n10622 );
    xnor g1140 ( n14630 , n18410 , n29207 );
    xnor g1141 ( n23688 , n124 , n12958 );
    or g1142 ( n7389 , n23262 , n10762 );
    not g1143 ( n17376 , n4960 );
    or g1144 ( n4099 , n32770 , n22194 );
    or g1145 ( n22116 , n5539 , n22951 );
    xnor g1146 ( n14761 , n2815 , n6447 );
    and g1147 ( n31762 , n3826 , n16826 );
    xnor g1148 ( n10349 , n6605 , n34970 );
    or g1149 ( n27526 , n25271 , n4478 );
    or g1150 ( n25071 , n31211 , n5709 );
    and g1151 ( n21028 , n29365 , n21336 );
    and g1152 ( n16462 , n16301 , n34613 );
    nor g1153 ( n8233 , n20949 , n7877 );
    nor g1154 ( n30521 , n19984 , n21907 );
    or g1155 ( n325 , n11046 , n6807 );
    xnor g1156 ( n13820 , n4273 , n23604 );
    or g1157 ( n18830 , n12029 , n28410 );
    nor g1158 ( n30348 , n8582 , n18151 );
    nor g1159 ( n23976 , n22512 , n23921 );
    or g1160 ( n19562 , n11714 , n29872 );
    xnor g1161 ( n23540 , n12455 , n34235 );
    and g1162 ( n4421 , n4575 , n25853 );
    and g1163 ( n15695 , n35571 , n28313 );
    or g1164 ( n26617 , n15356 , n16345 );
    or g1165 ( n11766 , n19551 , n14882 );
    and g1166 ( n21077 , n20233 , n13481 );
    xnor g1167 ( n4325 , n29027 , n14483 );
    and g1168 ( n9692 , n3336 , n28164 );
    xnor g1169 ( n8577 , n20709 , n18556 );
    or g1170 ( n35611 , n24608 , n20762 );
    or g1171 ( n5104 , n8780 , n27728 );
    or g1172 ( n14922 , n29713 , n27370 );
    buf g1173 ( n19241 , n25761 );
    nor g1174 ( n6693 , n24332 , n28871 );
    or g1175 ( n3275 , n17715 , n22868 );
    or g1176 ( n35160 , n34286 , n29349 );
    or g1177 ( n20393 , n5087 , n15144 );
    xnor g1178 ( n13271 , n19635 , n31173 );
    not g1179 ( n33494 , n1950 );
    or g1180 ( n14525 , n29713 , n24458 );
    not g1181 ( n15011 , n29574 );
    or g1182 ( n238 , n15372 , n20930 );
    or g1183 ( n1182 , n35052 , n14286 );
    xnor g1184 ( n10434 , n212 , n4288 );
    or g1185 ( n26780 , n11215 , n10289 );
    or g1186 ( n35140 , n21054 , n10057 );
    and g1187 ( n29783 , n29257 , n15408 );
    or g1188 ( n33445 , n11882 , n5972 );
    not g1189 ( n7167 , n30204 );
    not g1190 ( n5171 , n22291 );
    or g1191 ( n8006 , n22972 , n763 );
    or g1192 ( n16221 , n7612 , n25658 );
    xnor g1193 ( n25813 , n21680 , n4288 );
    xnor g1194 ( n22285 , n3443 , n24332 );
    or g1195 ( n10511 , n27807 , n28438 );
    nor g1196 ( n4607 , n20790 , n4514 );
    nor g1197 ( n31997 , n32857 , n14458 );
    or g1198 ( n22388 , n8299 , n8950 );
    not g1199 ( n11718 , n14289 );
    or g1200 ( n4594 , n35676 , n24357 );
    or g1201 ( n21833 , n27763 , n15256 );
    xnor g1202 ( n4991 , n3776 , n17751 );
    xnor g1203 ( n28529 , n17643 , n12781 );
    and g1204 ( n397 , n35117 , n2806 );
    or g1205 ( n27390 , n18535 , n23490 );
    or g1206 ( n32004 , n28070 , n13480 );
    and g1207 ( n503 , n6292 , n13622 );
    xnor g1208 ( n12102 , n34676 , n24332 );
    nor g1209 ( n7056 , n31215 , n25026 );
    or g1210 ( n10113 , n35280 , n7844 );
    xnor g1211 ( n22979 , n1581 , n9592 );
    nor g1212 ( n32516 , n10568 , n10065 );
    xnor g1213 ( n32975 , n9150 , n16216 );
    or g1214 ( n28274 , n23522 , n20427 );
    xnor g1215 ( n28001 , n8325 , n2860 );
    or g1216 ( n15810 , n17063 , n22780 );
    nor g1217 ( n6069 , n14749 , n35699 );
    and g1218 ( n11241 , n670 , n26565 );
    or g1219 ( n30596 , n28882 , n2712 );
    not g1220 ( n8866 , n25602 );
    xnor g1221 ( n11574 , n30777 , n79 );
    nor g1222 ( n24775 , n16620 , n33325 );
    nor g1223 ( n17837 , n6120 , n28739 );
    nor g1224 ( n9825 , n31804 , n34869 );
    and g1225 ( n27631 , n21346 , n6407 );
    and g1226 ( n8585 , n8765 , n3123 );
    or g1227 ( n27087 , n25923 , n25219 );
    or g1228 ( n33187 , n21867 , n23323 );
    or g1229 ( n30245 , n30246 , n3239 );
    nor g1230 ( n22550 , n9014 , n6017 );
    or g1231 ( n31092 , n10783 , n34723 );
    not g1232 ( n21508 , n16620 );
    and g1233 ( n11846 , n35251 , n28977 );
    and g1234 ( n18388 , n23962 , n35137 );
    xnor g1235 ( n28692 , n29038 , n3205 );
    or g1236 ( n24540 , n35927 , n9816 );
    or g1237 ( n4319 , n32404 , n20074 );
    xnor g1238 ( n30768 , n18137 , n25757 );
    or g1239 ( n7837 , n30748 , n7381 );
    xnor g1240 ( n23756 , n29696 , n7964 );
    or g1241 ( n17679 , n10433 , n27447 );
    xnor g1242 ( n29329 , n2455 , n721 );
    and g1243 ( n20285 , n32121 , n18070 );
    or g1244 ( n5858 , n30658 , n33416 );
    or g1245 ( n31527 , n31289 , n20626 );
    and g1246 ( n17016 , n23251 , n28386 );
    and g1247 ( n12221 , n8003 , n33576 );
    or g1248 ( n27535 , n4288 , n28770 );
    or g1249 ( n1531 , n13027 , n26365 );
    or g1250 ( n30889 , n21499 , n28438 );
    and g1251 ( n11855 , n1473 , n35733 );
    xnor g1252 ( n5683 , n28822 , n10894 );
    or g1253 ( n32613 , n30742 , n9418 );
    and g1254 ( n23450 , n4535 , n15712 );
    xnor g1255 ( n34830 , n31220 , n27291 );
    or g1256 ( n19684 , n16253 , n7703 );
    and g1257 ( n32190 , n1023 , n25365 );
    or g1258 ( n4466 , n4878 , n16666 );
    or g1259 ( n5622 , n14811 , n26002 );
    or g1260 ( n24739 , n30505 , n3374 );
    xnor g1261 ( n1918 , n11808 , n4878 );
    or g1262 ( n14460 , n22701 , n20797 );
    or g1263 ( n34872 , n22313 , n13900 );
    or g1264 ( n21719 , n33529 , n22206 );
    nor g1265 ( n36020 , n10894 , n2721 );
    and g1266 ( n34096 , n14795 , n16947 );
    or g1267 ( n19250 , n30786 , n34862 );
    and g1268 ( n23924 , n4731 , n23200 );
    or g1269 ( n6390 , n33162 , n6998 );
    not g1270 ( n12371 , n31289 );
    not g1271 ( n17793 , n28404 );
    and g1272 ( n26356 , n5511 , n11278 );
    or g1273 ( n14878 , n7496 , n7118 );
    xnor g1274 ( n8188 , n9913 , n22161 );
    xnor g1275 ( n7286 , n34640 , n35532 );
    and g1276 ( n13857 , n22521 , n27938 );
    or g1277 ( n26906 , n24511 , n5968 );
    not g1278 ( n3430 , n4275 );
    not g1279 ( n4928 , n8432 );
    or g1280 ( n18454 , n33311 , n22946 );
    or g1281 ( n5387 , n34013 , n10960 );
    xnor g1282 ( n14831 , n28096 , n28398 );
    or g1283 ( n17439 , n1660 , n26737 );
    or g1284 ( n27845 , n2232 , n908 );
    or g1285 ( n28871 , n27196 , n34559 );
    xnor g1286 ( n28394 , n25873 , n20852 );
    and g1287 ( n33042 , n6467 , n20047 );
    and g1288 ( n27743 , n24500 , n6598 );
    or g1289 ( n646 , n9261 , n19091 );
    or g1290 ( n25689 , n5257 , n10762 );
    xnor g1291 ( n26083 , n22570 , n4878 );
    or g1292 ( n15840 , n9658 , n35328 );
    and g1293 ( n7065 , n31441 , n9189 );
    not g1294 ( n26286 , n25909 );
    and g1295 ( n19678 , n387 , n29637 );
    and g1296 ( n28211 , n5373 , n26554 );
    not g1297 ( n18808 , n30711 );
    and g1298 ( n27201 , n12327 , n22625 );
    or g1299 ( n16362 , n12423 , n20817 );
    or g1300 ( n9337 , n27027 , n3461 );
    xnor g1301 ( n33702 , n6591 , n4962 );
    and g1302 ( n24920 , n5589 , n18147 );
    or g1303 ( n14359 , n18181 , n26112 );
    and g1304 ( n28246 , n2244 , n16429 );
    xnor g1305 ( n2357 , n34664 , n11046 );
    xnor g1306 ( n24689 , n10454 , n27870 );
    and g1307 ( n13685 , n11127 , n15735 );
    nor g1308 ( n10723 , n9789 , n12984 );
    and g1309 ( n30504 , n16645 , n4586 );
    or g1310 ( n21023 , n29829 , n5252 );
    xnor g1311 ( n24902 , n12594 , n21787 );
    xnor g1312 ( n25074 , n5376 , n32715 );
    xnor g1313 ( n9116 , n1082 , n13117 );
    or g1314 ( n24178 , n27261 , n13117 );
    xnor g1315 ( n338 , n35579 , n31289 );
    and g1316 ( n35506 , n5050 , n21194 );
    or g1317 ( n33860 , n3937 , n5619 );
    or g1318 ( n15189 , n11935 , n9555 );
    and g1319 ( n20584 , n20800 , n7012 );
    or g1320 ( n13318 , n6085 , n24701 );
    xnor g1321 ( n32573 , n17890 , n11089 );
    or g1322 ( n7131 , n15886 , n35212 );
    or g1323 ( n17704 , n16200 , n28248 );
    and g1324 ( n26374 , n26065 , n29297 );
    nor g1325 ( n13322 , n3946 , n27397 );
    not g1326 ( n13878 , n10504 );
    or g1327 ( n19699 , n413 , n5457 );
    xnor g1328 ( n15343 , n35684 , n5232 );
    not g1329 ( n11785 , n21971 );
    or g1330 ( n13725 , n16023 , n3805 );
    nor g1331 ( n12451 , n9658 , n23427 );
    xnor g1332 ( n31533 , n31538 , n32095 );
    xnor g1333 ( n19309 , n32705 , n35221 );
    or g1334 ( n28588 , n35381 , n11258 );
    and g1335 ( n12165 , n28079 , n28708 );
    not g1336 ( n28788 , n3239 );
    nor g1337 ( n2821 , n15166 , n11029 );
    or g1338 ( n5492 , n26563 , n18423 );
    and g1339 ( n22604 , n17630 , n23295 );
    xnor g1340 ( n26362 , n12447 , n27226 );
    xnor g1341 ( n11911 , n29390 , n3205 );
    and g1342 ( n22945 , n7031 , n18444 );
    or g1343 ( n29564 , n17619 , n14746 );
    and g1344 ( n13936 , n13519 , n4115 );
    or g1345 ( n1521 , n19948 , n16533 );
    nor g1346 ( n9726 , n31289 , n11391 );
    xnor g1347 ( n12815 , n22822 , n21701 );
    or g1348 ( n25765 , n4097 , n18275 );
    or g1349 ( n16899 , n17814 , n30318 );
    or g1350 ( n5051 , n20841 , n17429 );
    or g1351 ( n30984 , n24457 , n10634 );
    and g1352 ( n16875 , n10250 , n12765 );
    and g1353 ( n14770 , n7231 , n29618 );
    xor g1354 ( n30416 , n32619 , n12167 );
    nor g1355 ( n20161 , n30742 , n27773 );
    or g1356 ( n25130 , n7759 , n18655 );
    and g1357 ( n2876 , n20769 , n17266 );
    and g1358 ( n13062 , n8626 , n18511 );
    nor g1359 ( n33899 , n15464 , n24707 );
    nor g1360 ( n5697 , n25174 , n20517 );
    buf g1361 ( n25592 , n34395 );
    nor g1362 ( n11598 , n28938 , n19137 );
    xnor g1363 ( n29161 , n27822 , n830 );
    nor g1364 ( n9546 , n13527 , n11077 );
    or g1365 ( n35759 , n33487 , n3968 );
    and g1366 ( n27010 , n33722 , n3244 );
    xnor g1367 ( n33666 , n33280 , n16876 );
    xnor g1368 ( n28862 , n9556 , n31289 );
    not g1369 ( n25197 , n22471 );
    and g1370 ( n21798 , n14430 , n3764 );
    or g1371 ( n15177 , n28494 , n26429 );
    or g1372 ( n3025 , n9849 , n3378 );
    not g1373 ( n34440 , n17568 );
    nor g1374 ( n14784 , n25677 , n19834 );
    or g1375 ( n9330 , n11625 , n10081 );
    or g1376 ( n27072 , n8737 , n25683 );
    or g1377 ( n11835 , n14986 , n31034 );
    xnor g1378 ( n24210 , n13332 , n3222 );
    and g1379 ( n18402 , n30837 , n12422 );
    or g1380 ( n13180 , n21038 , n15439 );
    and g1381 ( n34829 , n8916 , n5254 );
    or g1382 ( n26122 , n17791 , n7726 );
    or g1383 ( n17229 , n13940 , n27262 );
    xnor g1384 ( n10098 , n24617 , n436 );
    not g1385 ( n31227 , n3222 );
    xnor g1386 ( n925 , n17886 , n9550 );
    or g1387 ( n21292 , n838 , n21956 );
    xor g1388 ( n31788 , n22186 , n4700 );
    or g1389 ( n16406 , n29467 , n35961 );
    and g1390 ( n26849 , n4202 , n33308 );
    and g1391 ( n2416 , n23692 , n24116 );
    and g1392 ( n20626 , n5125 , n7911 );
    or g1393 ( n34124 , n28254 , n2168 );
    or g1394 ( n33377 , n34586 , n8910 );
    and g1395 ( n11447 , n15685 , n10916 );
    or g1396 ( n26987 , n33929 , n14506 );
    xnor g1397 ( n23743 , n28708 , n28079 );
    xnor g1398 ( n7393 , n29082 , n16041 );
    buf g1399 ( n14699 , n9006 );
    xnor g1400 ( n1533 , n30042 , n20605 );
    not g1401 ( n31477 , n10894 );
    or g1402 ( n24036 , n33520 , n35043 );
    nor g1403 ( n28894 , n21545 , n27363 );
    and g1404 ( n5615 , n6836 , n19961 );
    and g1405 ( n10765 , n22515 , n2763 );
    and g1406 ( n1155 , n17112 , n1385 );
    and g1407 ( n1172 , n16782 , n15392 );
    or g1408 ( n28233 , n7112 , n10400 );
    not g1409 ( n31429 , n29713 );
    or g1410 ( n30420 , n689 , n19490 );
    or g1411 ( n27369 , n24132 , n20797 );
    not g1412 ( n9358 , n11440 );
    and g1413 ( n35587 , n15681 , n16306 );
    xnor g1414 ( n18365 , n28534 , n30196 );
    xnor g1415 ( n28556 , n17532 , n7540 );
    or g1416 ( n22998 , n22440 , n17401 );
    and g1417 ( n6956 , n14205 , n32824 );
    xnor g1418 ( n35811 , n28470 , n32123 );
    or g1419 ( n21831 , n22113 , n19983 );
    xnor g1420 ( n26375 , n6973 , n16110 );
    or g1421 ( n30837 , n10157 , n30732 );
    and g1422 ( n29629 , n28722 , n27524 );
    nor g1423 ( n23559 , n25351 , n17825 );
    and g1424 ( n29225 , n5454 , n3868 );
    and g1425 ( n36035 , n33855 , n24632 );
    xor g1426 ( n17398 , n22369 , n32340 );
    and g1427 ( n10345 , n34572 , n19436 );
    or g1428 ( n16052 , n13553 , n3251 );
    and g1429 ( n9499 , n728 , n25579 );
    xnor g1430 ( n20685 , n33947 , n32095 );
    and g1431 ( n10656 , n28570 , n4620 );
    xnor g1432 ( n30785 , n24847 , n2315 );
    not g1433 ( n13905 , n34923 );
    or g1434 ( n28874 , n22237 , n4363 );
    or g1435 ( n19416 , n12872 , n12511 );
    not g1436 ( n2533 , n22850 );
    and g1437 ( n20808 , n15309 , n22465 );
    or g1438 ( n1984 , n32584 , n1801 );
    xnor g1439 ( n29469 , n10389 , n11190 );
    xnor g1440 ( n17295 , n15056 , n1950 );
    and g1441 ( n21802 , n5347 , n10047 );
    or g1442 ( n8120 , n33804 , n11982 );
    xnor g1443 ( n23796 , n13326 , n15886 );
    nor g1444 ( n35181 , n11924 , n19619 );
    or g1445 ( n13506 , n23722 , n30204 );
    or g1446 ( n5444 , n27084 , n20690 );
    or g1447 ( n29689 , n12459 , n5752 );
    or g1448 ( n30176 , n7540 , n24626 );
    nor g1449 ( n3466 , n33977 , n14375 );
    xnor g1450 ( n18797 , n19011 , n26419 );
    xnor g1451 ( n23255 , n32719 , n4962 );
    xnor g1452 ( n15330 , n15105 , n27116 );
    and g1453 ( n16622 , n11779 , n3037 );
    or g1454 ( n11804 , n5 , n14361 );
    nor g1455 ( n17773 , n7024 , n25197 );
    xnor g1456 ( n23817 , n24959 , n21735 );
    and g1457 ( n10410 , n17943 , n28432 );
    xnor g1458 ( n5179 , n21615 , n7221 );
    and g1459 ( n34029 , n21403 , n19250 );
    or g1460 ( n14576 , n830 , n18958 );
    or g1461 ( n23600 , n17564 , n23410 );
    and g1462 ( n5696 , n9177 , n16712 );
    xnor g1463 ( n4370 , n20713 , n30151 );
    or g1464 ( n35382 , n14789 , n24431 );
    or g1465 ( n5951 , n17415 , n13217 );
    xnor g1466 ( n35365 , n7428 , n29098 );
    xnor g1467 ( n34802 , n13020 , n4719 );
    or g1468 ( n18241 , n16180 , n2524 );
    nor g1469 ( n12174 , n14540 , n12926 );
    xnor g1470 ( n9068 , n91 , n9789 );
    or g1471 ( n24572 , n26922 , n12622 );
    and g1472 ( n9429 , n34026 , n778 );
    xnor g1473 ( n28419 , n22259 , n30024 );
    xnor g1474 ( n2439 , n33186 , n9236 );
    or g1475 ( n22187 , n25174 , n32493 );
    or g1476 ( n6201 , n20240 , n14723 );
    nor g1477 ( n3693 , n20067 , n27501 );
    or g1478 ( n11945 , n31215 , n22544 );
    and g1479 ( n20681 , n27641 , n20370 );
    nor g1480 ( n14118 , n10894 , n5111 );
    xnor g1481 ( n30231 , n16244 , n17140 );
    and g1482 ( n3923 , n28670 , n33242 );
    xnor g1483 ( n12312 , n12590 , n32649 );
    and g1484 ( n15611 , n27248 , n28687 );
    xnor g1485 ( n33195 , n31601 , n4962 );
    or g1486 ( n7134 , n18260 , n7647 );
    not g1487 ( n26282 , n18296 );
    or g1488 ( n30644 , n29884 , n27465 );
    or g1489 ( n32306 , n5937 , n27053 );
    and g1490 ( n20310 , n23357 , n21290 );
    xnor g1491 ( n22022 , n17912 , n32435 );
    or g1492 ( n16370 , n34311 , n18230 );
    nor g1493 ( n31982 , n26028 , n19834 );
    and g1494 ( n23854 , n30329 , n34032 );
    and g1495 ( n19263 , n35129 , n1128 );
    or g1496 ( n1773 , n9885 , n564 );
    and g1497 ( n27310 , n24481 , n9199 );
    or g1498 ( n21872 , n9460 , n15416 );
    xnor g1499 ( n34242 , n21354 , n22291 );
    or g1500 ( n30447 , n19192 , n1520 );
    xnor g1501 ( n9246 , n8643 , n27440 );
    or g1502 ( n28885 , n23628 , n16570 );
    buf g1503 ( n11601 , n2609 );
    xnor g1504 ( n15173 , n13135 , n8539 );
    xor g1505 ( n23589 , n15769 , n25079 );
    or g1506 ( n9324 , n28220 , n7726 );
    buf g1507 ( n33956 , n29203 );
    xnor g1508 ( n14730 , n7797 , n16264 );
    or g1509 ( n18425 , n34013 , n8025 );
    xnor g1510 ( n17175 , n20887 , n27226 );
    xnor g1511 ( n8829 , n1801 , n32584 );
    or g1512 ( n630 , n28831 , n23921 );
    not g1513 ( n22467 , n28756 );
    or g1514 ( n10520 , n7756 , n1245 );
    or g1515 ( n9869 , n2710 , n8090 );
    or g1516 ( n9691 , n33040 , n5290 );
    and g1517 ( n11355 , n18987 , n32786 );
    and g1518 ( n2191 , n33081 , n24748 );
    and g1519 ( n27947 , n22516 , n17770 );
    or g1520 ( n23472 , n1191 , n12703 );
    xnor g1521 ( n32519 , n6309 , n30742 );
    not g1522 ( n9723 , n4487 );
    xnor g1523 ( n8170 , n35154 , n7664 );
    not g1524 ( n35627 , n28865 );
    and g1525 ( n9796 , n35755 , n25257 );
    or g1526 ( n34508 , n28414 , n13307 );
    and g1527 ( n27343 , n32606 , n19511 );
    xnor g1528 ( n15007 , n17016 , n33629 );
    and g1529 ( n16423 , n32161 , n18342 );
    or g1530 ( n13655 , n831 , n4172 );
    not g1531 ( n18893 , n4250 );
    and g1532 ( n24853 , n29697 , n30411 );
    and g1533 ( n4981 , n9084 , n20309 );
    nor g1534 ( n13384 , n9837 , n25508 );
    or g1535 ( n19492 , n4598 , n28969 );
    nor g1536 ( n26891 , n17484 , n12001 );
    and g1537 ( n10995 , n20728 , n31102 );
    and g1538 ( n8845 , n12722 , n13434 );
    not g1539 ( n12234 , n31647 );
    nor g1540 ( n25421 , n15380 , n13643 );
    not g1541 ( n22001 , n6927 );
    or g1542 ( n20658 , n10894 , n9413 );
    xnor g1543 ( n15397 , n15048 , n27405 );
    and g1544 ( n28021 , n9272 , n6841 );
    or g1545 ( n22878 , n28163 , n16543 );
    or g1546 ( n2465 , n25174 , n17869 );
    and g1547 ( n35717 , n60 , n15118 );
    and g1548 ( n5080 , n32159 , n27510 );
    not g1549 ( n13649 , n11810 );
    and g1550 ( n19087 , n10658 , n27357 );
    xnor g1551 ( n11339 , n11377 , n29571 );
    or g1552 ( n21900 , n29094 , n2798 );
    xnor g1553 ( n30746 , n17806 , n30742 );
    and g1554 ( n33167 , n4145 , n24883 );
    xnor g1555 ( n24476 , n1888 , n28804 );
    or g1556 ( n19138 , n21629 , n11601 );
    xnor g1557 ( n24439 , n21544 , n17413 );
    or g1558 ( n17205 , n19554 , n21569 );
    or g1559 ( n36011 , n24371 , n26283 );
    or g1560 ( n1532 , n29782 , n22858 );
    nor g1561 ( n20199 , n3222 , n15813 );
    or g1562 ( n30291 , n2152 , n9951 );
    nor g1563 ( n29167 , n22153 , n7153 );
    and g1564 ( n4522 , n4093 , n15421 );
    buf g1565 ( n19125 , n26388 );
    xnor g1566 ( n26582 , n19841 , n19061 );
    and g1567 ( n10288 , n21789 , n19803 );
    xnor g1568 ( n16202 , n6884 , n30851 );
    xnor g1569 ( n2564 , n35325 , n11060 );
    and g1570 ( n32679 , n31515 , n3305 );
    or g1571 ( n14305 , n22383 , n8090 );
    or g1572 ( n19753 , n13122 , n26077 );
    and g1573 ( n17438 , n32320 , n9788 );
    and g1574 ( n16944 , n18666 , n32301 );
    or g1575 ( n26435 , n10168 , n9731 );
    or g1576 ( n35896 , n19015 , n16762 );
    and g1577 ( n17101 , n34562 , n17801 );
    nor g1578 ( n30237 , n15886 , n7618 );
    xnor g1579 ( n3654 , n23030 , n19551 );
    not g1580 ( n22850 , n11714 );
    not g1581 ( n28384 , n22119 );
    nor g1582 ( n24274 , n11392 , n2581 );
    xnor g1583 ( n35673 , n26678 , n18253 );
    and g1584 ( n3093 , n15039 , n23941 );
    or g1585 ( n21911 , n19139 , n5711 );
    and g1586 ( n32176 , n14152 , n10638 );
    not g1587 ( n10159 , n22980 );
    and g1588 ( n26179 , n24384 , n1493 );
    and g1589 ( n4609 , n15970 , n25358 );
    and g1590 ( n28700 , n7631 , n3125 );
    and g1591 ( n27176 , n18386 , n18619 );
    buf g1592 ( n32507 , n30047 );
    and g1593 ( n13910 , n7201 , n4614 );
    xnor g1594 ( n11162 , n7560 , n28533 );
    and g1595 ( n852 , n26945 , n9666 );
    and g1596 ( n26686 , n24378 , n29673 );
    and g1597 ( n5917 , n13403 , n17502 );
    xnor g1598 ( n4310 , n9161 , n31799 );
    or g1599 ( n17489 , n25602 , n9349 );
    and g1600 ( n4955 , n30966 , n19749 );
    not g1601 ( n21531 , n7540 );
    or g1602 ( n30910 , n26966 , n22206 );
    not g1603 ( n6819 , n18333 );
    and g1604 ( n19875 , n23223 , n11217 );
    xnor g1605 ( n5236 , n15168 , n16922 );
    or g1606 ( n21973 , n4288 , n10445 );
    or g1607 ( n24503 , n25602 , n27505 );
    and g1608 ( n4467 , n16677 , n9221 );
    or g1609 ( n6955 , n20137 , n25560 );
    or g1610 ( n30458 , n25250 , n32843 );
    not g1611 ( n29011 , n31056 );
    xnor g1612 ( n13005 , n29389 , n23757 );
    or g1613 ( n27156 , n22291 , n1797 );
    or g1614 ( n2204 , n17393 , n740 );
    or g1615 ( n14020 , n28419 , n28248 );
    and g1616 ( n17356 , n34033 , n15069 );
    or g1617 ( n26378 , n27994 , n22206 );
    or g1618 ( n26663 , n4962 , n19106 );
    xnor g1619 ( n18578 , n30626 , n34185 );
    or g1620 ( n9532 , n4004 , n23627 );
    or g1621 ( n27117 , n30742 , n6309 );
    or g1622 ( n8297 , n913 , n27625 );
    or g1623 ( n14454 , n18559 , n34862 );
    or g1624 ( n7120 , n29967 , n20762 );
    nor g1625 ( n10561 , n25602 , n24873 );
    xnor g1626 ( n32472 , n3859 , n19896 );
    not g1627 ( n8302 , n25245 );
    or g1628 ( n26216 , n6352 , n27580 );
    or g1629 ( n17464 , n24537 , n11712 );
    and g1630 ( n20053 , n8256 , n29 );
    or g1631 ( n24052 , n3548 , n12996 );
    or g1632 ( n24848 , n6369 , n40 );
    or g1633 ( n29344 , n26320 , n35422 );
    and g1634 ( n3356 , n32869 , n20524 );
    and g1635 ( n7720 , n21262 , n24994 );
    and g1636 ( n21532 , n2761 , n8794 );
    or g1637 ( n20649 , n15886 , n8748 );
    nor g1638 ( n24855 , n11672 , n18115 );
    or g1639 ( n3286 , n32584 , n24552 );
    and g1640 ( n32295 , n16765 , n17927 );
    or g1641 ( n25919 , n5127 , n2712 );
    xnor g1642 ( n21440 , n32040 , n28189 );
    or g1643 ( n17397 , n10894 , n10965 );
    xnor g1644 ( n33424 , n11838 , n27213 );
    and g1645 ( n6812 , n8812 , n25738 );
    not g1646 ( n17768 , n33810 );
    not g1647 ( n25183 , n36066 );
    not g1648 ( n17056 , n29409 );
    not g1649 ( n30898 , n20933 );
    or g1650 ( n4062 , n16394 , n21042 );
    xnor g1651 ( n15734 , n34132 , n3481 );
    xnor g1652 ( n14971 , n11693 , n14197 );
    not g1653 ( n26214 , n23093 );
    or g1654 ( n16963 , n13036 , n9930 );
    xnor g1655 ( n7300 , n8186 , n830 );
    nor g1656 ( n20085 , n18578 , n24505 );
    and g1657 ( n18610 , n14131 , n29523 );
    xnor g1658 ( n25320 , n13979 , n24497 );
    or g1659 ( n14413 , n30511 , n20300 );
    or g1660 ( n28427 , n6392 , n1557 );
    xnor g1661 ( n20904 , n11048 , n35927 );
    xnor g1662 ( n25239 , n21822 , n31289 );
    or g1663 ( n6471 , n28 , n20812 );
    buf g1664 ( n20762 , n35237 );
    or g1665 ( n9 , n16469 , n32572 );
    or g1666 ( n33873 , n9269 , n15805 );
    or g1667 ( n27835 , n9658 , n33993 );
    nor g1668 ( n8058 , n11046 , n21890 );
    xnor g1669 ( n19051 , n23919 , n3205 );
    or g1670 ( n11563 , n16240 , n32697 );
    xnor g1671 ( n35793 , n25329 , n20194 );
    and g1672 ( n12086 , n29107 , n22702 );
    xnor g1673 ( n6053 , n27431 , n10314 );
    or g1674 ( n16859 , n10615 , n20784 );
    and g1675 ( n28633 , n16142 , n8458 );
    or g1676 ( n7695 , n22063 , n17068 );
    and g1677 ( n20733 , n1013 , n33985 );
    and g1678 ( n21405 , n31940 , n29825 );
    xnor g1679 ( n31679 , n34041 , n3946 );
    nor g1680 ( n19642 , n33535 , n19834 );
    or g1681 ( n17142 , n7142 , n33557 );
    not g1682 ( n22992 , n5335 );
    xnor g1683 ( n11208 , n9525 , n10440 );
    or g1684 ( n650 , n35830 , n26503 );
    nor g1685 ( n17531 , n8094 , n27096 );
    or g1686 ( n9686 , n18924 , n26442 );
    not g1687 ( n7214 , n11712 );
    or g1688 ( n701 , n32857 , n28181 );
    not g1689 ( n29672 , n35289 );
    not g1690 ( n34563 , n10897 );
    and g1691 ( n22916 , n23472 , n20702 );
    nor g1692 ( n23518 , n9793 , n32255 );
    or g1693 ( n1188 , n19038 , n11833 );
    or g1694 ( n19484 , n26134 , n10094 );
    and g1695 ( n32255 , n14935 , n35207 );
    nor g1696 ( n4904 , n3205 , n32911 );
    and g1697 ( n35589 , n21333 , n10056 );
    xnor g1698 ( n358 , n17479 , n854 );
    and g1699 ( n9328 , n4272 , n6751 );
    or g1700 ( n18450 , n27937 , n20817 );
    or g1701 ( n6507 , n17425 , n21207 );
    or g1702 ( n20884 , n11555 , n4081 );
    and g1703 ( n25322 , n1309 , n19108 );
    xnor g1704 ( n12712 , n21029 , n34909 );
    and g1705 ( n25610 , n14186 , n22187 );
    or g1706 ( n30606 , n30742 , n17081 );
    xnor g1707 ( n4869 , n6504 , n29839 );
    xnor g1708 ( n28772 , n29133 , n9617 );
    and g1709 ( n25744 , n24426 , n14036 );
    or g1710 ( n18909 , n3946 , n8890 );
    or g1711 ( n17924 , n30742 , n30515 );
    or g1712 ( n19347 , n27905 , n63 );
    xor g1713 ( n6423 , n22176 , n1918 );
    not g1714 ( n895 , n17751 );
    and g1715 ( n4464 , n12625 , n2322 );
    or g1716 ( n15773 , n5067 , n30807 );
    or g1717 ( n33651 , n5335 , n30054 );
    or g1718 ( n30464 , n13748 , n22577 );
    or g1719 ( n11410 , n35927 , n23173 );
    not g1720 ( n33464 , n11833 );
    or g1721 ( n17029 , n19245 , n1731 );
    nor g1722 ( n7714 , n20047 , n21757 );
    or g1723 ( n11803 , n4960 , n20838 );
    or g1724 ( n24340 , n32826 , n28191 );
    not g1725 ( n28655 , n20558 );
    and g1726 ( n20517 , n32195 , n8141 );
    buf g1727 ( n13967 , n22876 );
    or g1728 ( n30079 , n23934 , n1306 );
    or g1729 ( n135 , n25602 , n34192 );
    and g1730 ( n24758 , n19016 , n35578 );
    or g1731 ( n10110 , n29885 , n2488 );
    xnor g1732 ( n23886 , n21169 , n22357 );
    or g1733 ( n14814 , n22944 , n13015 );
    xnor g1734 ( n2560 , n31156 , n17093 );
    or g1735 ( n8605 , n31215 , n34002 );
    not g1736 ( n12731 , n13016 );
    or g1737 ( n13819 , n20159 , n12332 );
    and g1738 ( n9265 , n22133 , n28378 );
    nor g1739 ( n19634 , n12779 , n34084 );
    or g1740 ( n31410 , n21798 , n128 );
    xnor g1741 ( n31630 , n35704 , n19169 );
    buf g1742 ( n3188 , n905 );
    not g1743 ( n2827 , n12747 );
    or g1744 ( n28508 , n4288 , n17075 );
    or g1745 ( n16214 , n8938 , n4523 );
    nor g1746 ( n24889 , n11046 , n14239 );
    or g1747 ( n12642 , n3440 , n33543 );
    xnor g1748 ( n26716 , n29902 , n24332 );
    nor g1749 ( n29090 , n29713 , n27995 );
    xnor g1750 ( n3976 , n9222 , n20780 );
    nor g1751 ( n1175 , n22291 , n34334 );
    or g1752 ( n2011 , n2726 , n4912 );
    nor g1753 ( n11005 , n2457 , n1402 );
    xor g1754 ( n14993 , n3380 , n26212 );
    xnor g1755 ( n21451 , n12768 , n8636 );
    or g1756 ( n4927 , n17568 , n31582 );
    or g1757 ( n24712 , n8156 , n20595 );
    or g1758 ( n27904 , n31875 , n21490 );
    and g1759 ( n27707 , n1318 , n1702 );
    or g1760 ( n12755 , n1195 , n18542 );
    and g1761 ( n25526 , n8730 , n30184 );
    or g1762 ( n2923 , n3623 , n6958 );
    or g1763 ( n26546 , n31272 , n14039 );
    or g1764 ( n7821 , n35434 , n34727 );
    or g1765 ( n11072 , n8604 , n12791 );
    xnor g1766 ( n31426 , n17718 , n10089 );
    xnor g1767 ( n11806 , n18861 , n19631 );
    or g1768 ( n20195 , n12894 , n3736 );
    and g1769 ( n30023 , n4403 , n34914 );
    xnor g1770 ( n20627 , n13046 , n29977 );
    buf g1771 ( n6075 , n16910 );
    or g1772 ( n13105 , n4762 , n12206 );
    or g1773 ( n17797 , n23996 , n16464 );
    or g1774 ( n754 , n29886 , n16768 );
    and g1775 ( n12753 , n36018 , n32372 );
    or g1776 ( n33026 , n9775 , n21691 );
    and g1777 ( n34272 , n1949 , n29920 );
    and g1778 ( n30149 , n16334 , n16713 );
    or g1779 ( n12948 , n18379 , n32491 );
    nor g1780 ( n2832 , n29141 , n7943 );
    or g1781 ( n22785 , n7599 , n25067 );
    xnor g1782 ( n2493 , n19249 , n15548 );
    nor g1783 ( n14144 , n32715 , n21372 );
    and g1784 ( n19328 , n5834 , n26202 );
    xnor g1785 ( n17660 , n14846 , n35490 );
    or g1786 ( n17251 , n21906 , n35977 );
    or g1787 ( n25630 , n32019 , n25075 );
    or g1788 ( n15712 , n22291 , n13745 );
    not g1789 ( n28130 , n4758 );
    and g1790 ( n11193 , n22905 , n7059 );
    and g1791 ( n10873 , n28129 , n9250 );
    or g1792 ( n25782 , n16061 , n21343 );
    or g1793 ( n4618 , n5664 , n21964 );
    and g1794 ( n23786 , n7602 , n28012 );
    xnor g1795 ( n26436 , n29802 , n29839 );
    or g1796 ( n17528 , n9413 , n19421 );
    or g1797 ( n35560 , n22275 , n3188 );
    and g1798 ( n24704 , n10580 , n28319 );
    nor g1799 ( n31138 , n830 , n20368 );
    or g1800 ( n30534 , n25174 , n20870 );
    or g1801 ( n12893 , n11246 , n11218 );
    xnor g1802 ( n31851 , n8920 , n18379 );
    xnor g1803 ( n26596 , n14619 , n1592 );
    or g1804 ( n31639 , n16261 , n18542 );
    xnor g1805 ( n411 , n10173 , n9602 );
    or g1806 ( n16029 , n18920 , n26225 );
    xnor g1807 ( n3475 , n3803 , n96 );
    xnor g1808 ( n20894 , n7997 , n29050 );
    xnor g1809 ( n8994 , n18087 , n4960 );
    xnor g1810 ( n28325 , n26571 , n3110 );
    or g1811 ( n31856 , n32735 , n25786 );
    xnor g1812 ( n28658 , n1428 , n5335 );
    or g1813 ( n4153 , n14786 , n13900 );
    or g1814 ( n21733 , n35330 , n23205 );
    not g1815 ( n24043 , n29243 );
    nor g1816 ( n22492 , n32584 , n29949 );
    or g1817 ( n25869 , n21538 , n33964 );
    not g1818 ( n961 , n31559 );
    and g1819 ( n19930 , n19130 , n28413 );
    and g1820 ( n27735 , n33340 , n2709 );
    xnor g1821 ( n29908 , n5391 , n18998 );
    nor g1822 ( n10974 , n17568 , n9800 );
    and g1823 ( n12830 , n31873 , n8791 );
    or g1824 ( n16449 , n203 , n24529 );
    nor g1825 ( n20711 , n24583 , n32130 );
    and g1826 ( n18850 , n26288 , n35428 );
    xnor g1827 ( n34587 , n33929 , n14506 );
    xnor g1828 ( n31423 , n10544 , n25602 );
    or g1829 ( n9319 , n11569 , n4318 );
    or g1830 ( n16443 , n7896 , n2168 );
    xnor g1831 ( n34524 , n16584 , n23236 );
    or g1832 ( n29233 , n10731 , n19939 );
    xnor g1833 ( n23482 , n35778 , n25663 );
    not g1834 ( n27177 , n4878 );
    and g1835 ( n31740 , n1324 , n31870 );
    xnor g1836 ( n16205 , n785 , n36049 );
    and g1837 ( n24082 , n7490 , n8664 );
    or g1838 ( n2888 , n19675 , n9817 );
    or g1839 ( n24493 , n5021 , n25592 );
    or g1840 ( n18967 , n1885 , n1796 );
    and g1841 ( n25990 , n3318 , n16853 );
    not g1842 ( n25369 , n3858 );
    and g1843 ( n34555 , n27170 , n31452 );
    or g1844 ( n5781 , n24406 , n11548 );
    or g1845 ( n14385 , n29715 , n27437 );
    not g1846 ( n22061 , n28273 );
    xnor g1847 ( n14557 , n15601 , n13106 );
    buf g1848 ( n32808 , n15344 );
    or g1849 ( n14443 , n11096 , n139 );
    and g1850 ( n19267 , n2550 , n25800 );
    and g1851 ( n4948 , n15866 , n33594 );
    or g1852 ( n10741 , n26214 , n26082 );
    or g1853 ( n35581 , n14266 , n544 );
    xnor g1854 ( n25227 , n34143 , n12607 );
    xnor g1855 ( n33858 , n30701 , n9658 );
    or g1856 ( n8973 , n11190 , n22882 );
    or g1857 ( n20224 , n20804 , n10960 );
    not g1858 ( n11013 , n16620 );
    nor g1859 ( n23763 , n29187 , n28230 );
    not g1860 ( n22189 , n27489 );
    and g1861 ( n12487 , n28999 , n15467 );
    or g1862 ( n11221 , n11331 , n2005 );
    or g1863 ( n25718 , n33533 , n5868 );
    xnor g1864 ( n35940 , n5422 , n13230 );
    and g1865 ( n15677 , n9129 , n17103 );
    or g1866 ( n2741 , n22115 , n15144 );
    or g1867 ( n34592 , n15308 , n17962 );
    xnor g1868 ( n33186 , n34761 , n14278 );
    or g1869 ( n16861 , n675 , n12791 );
    or g1870 ( n2873 , n11747 , n13900 );
    or g1871 ( n5649 , n32390 , n29953 );
    xnor g1872 ( n1331 , n34813 , n787 );
    xnor g1873 ( n14797 , n18260 , n31215 );
    xnor g1874 ( n21716 , n4287 , n17775 );
    and g1875 ( n30096 , n17936 , n26694 );
    or g1876 ( n24256 , n4707 , n1557 );
    xnor g1877 ( n3785 , n33369 , n4249 );
    and g1878 ( n26055 , n25283 , n19651 );
    or g1879 ( n25210 , n2803 , n9809 );
    xnor g1880 ( n29150 , n34159 , n4962 );
    xnor g1881 ( n5959 , n12372 , n19799 );
    or g1882 ( n7440 , n21153 , n30519 );
    buf g1883 ( n33034 , n14611 );
    or g1884 ( n4579 , n15240 , n18477 );
    and g1885 ( n28305 , n30631 , n29906 );
    or g1886 ( n11865 , n13578 , n13900 );
    nor g1887 ( n9082 , n32008 , n7720 );
    or g1888 ( n16687 , n23907 , n22961 );
    or g1889 ( n22452 , n31624 , n20812 );
    or g1890 ( n29708 , n24371 , n24419 );
    or g1891 ( n22221 , n22948 , n16456 );
    or g1892 ( n3630 , n12535 , n33429 );
    xnor g1893 ( n2544 , n19820 , n11455 );
    xnor g1894 ( n23464 , n14344 , n26308 );
    or g1895 ( n11219 , n14680 , n15256 );
    or g1896 ( n697 , n32312 , n11676 );
    or g1897 ( n11793 , n25938 , n25940 );
    and g1898 ( n11812 , n950 , n11192 );
    or g1899 ( n33323 , n30944 , n8392 );
    or g1900 ( n29879 , n371 , n16328 );
    xnor g1901 ( n3220 , n369 , n21909 );
    or g1902 ( n12323 , n8429 , n3892 );
    or g1903 ( n13304 , n11056 , n12808 );
    or g1904 ( n28298 , n30742 , n31302 );
    xnor g1905 ( n5581 , n20488 , n15403 );
    buf g1906 ( n26002 , n20840 );
    not g1907 ( n17767 , n22980 );
    not g1908 ( n15250 , n16326 );
    or g1909 ( n27799 , n2320 , n26023 );
    or g1910 ( n29021 , n13566 , n25887 );
    and g1911 ( n21965 , n30584 , n17347 );
    nor g1912 ( n34284 , n4950 , n23037 );
    or g1913 ( n6534 , n21179 , n33871 );
    nor g1914 ( n12503 , n1178 , n1247 );
    or g1915 ( n15708 , n4842 , n26346 );
    or g1916 ( n2088 , n9501 , n24489 );
    nor g1917 ( n25420 , n16620 , n24353 );
    xnor g1918 ( n9884 , n25809 , n33869 );
    and g1919 ( n3058 , n883 , n919 );
    xnor g1920 ( n14168 , n925 , n7740 );
    or g1921 ( n32741 , n25336 , n17612 );
    xnor g1922 ( n22362 , n4678 , n22291 );
    or g1923 ( n32759 , n24332 , n4369 );
    or g1924 ( n4237 , n8611 , n9928 );
    nor g1925 ( n32495 , n33601 , n26022 );
    or g1926 ( n756 , n16620 , n33811 );
    or g1927 ( n3015 , n26745 , n34280 );
    xnor g1928 ( n29878 , n27710 , n11046 );
    not g1929 ( n12658 , n21622 );
    xnor g1930 ( n26194 , n17984 , n5287 );
    or g1931 ( n9807 , n483 , n10889 );
    and g1932 ( n34664 , n31308 , n5443 );
    or g1933 ( n22636 , n7043 , n25762 );
    nor g1934 ( n25678 , n26600 , n13963 );
    or g1935 ( n34944 , n13046 , n15497 );
    or g1936 ( n218 , n32857 , n22686 );
    or g1937 ( n8134 , n16819 , n21977 );
    and g1938 ( n8657 , n16783 , n27052 );
    xnor g1939 ( n1003 , n113 , n10894 );
    or g1940 ( n18889 , n22127 , n32697 );
    and g1941 ( n31927 , n8863 , n30529 );
    or g1942 ( n5652 , n8142 , n17446 );
    nor g1943 ( n35460 , n14829 , n33956 );
    xnor g1944 ( n5503 , n12093 , n9658 );
    and g1945 ( n3671 , n35966 , n32343 );
    or g1946 ( n33030 , n4962 , n5530 );
    not g1947 ( n6665 , n11046 );
    or g1948 ( n28277 , n20793 , n6748 );
    or g1949 ( n26279 , n21452 , n4490 );
    xnor g1950 ( n34879 , n11468 , n32095 );
    or g1951 ( n26552 , n17568 , n21147 );
    or g1952 ( n12971 , n15951 , n9117 );
    not g1953 ( n31822 , n24880 );
    and g1954 ( n29163 , n18081 , n14169 );
    not g1955 ( n1479 , n4960 );
    xnor g1956 ( n30407 , n19948 , n8486 );
    xnor g1957 ( n13389 , n8337 , n25602 );
    or g1958 ( n2101 , n17076 , n33098 );
    and g1959 ( n17173 , n29230 , n15703 );
    nor g1960 ( n24002 , n33811 , n25831 );
    or g1961 ( n11582 , n29935 , n28837 );
    or g1962 ( n12469 , n4098 , n16039 );
    and g1963 ( n33821 , n2116 , n76 );
    and g1964 ( n2646 , n6170 , n33779 );
    or g1965 ( n4159 , n29059 , n19058 );
    and g1966 ( n4090 , n6638 , n23817 );
    or g1967 ( n10004 , n13234 , n15144 );
    and g1968 ( n21935 , n14714 , n7816 );
    and g1969 ( n6743 , n24753 , n23804 );
    xnor g1970 ( n26830 , n15277 , n4914 );
    or g1971 ( n25572 , n30766 , n30611 );
    and g1972 ( n14949 , n12395 , n7391 );
    xnor g1973 ( n35881 , n7900 , n12209 );
    xnor g1974 ( n25873 , n23986 , n3222 );
    xnor g1975 ( n12632 , n18027 , n8866 );
    and g1976 ( n25695 , n6171 , n10680 );
    and g1977 ( n1524 , n6882 , n4456 );
    or g1978 ( n30618 , n4960 , n10433 );
    or g1979 ( n31933 , n9658 , n29829 );
    xnor g1980 ( n1330 , n11329 , n8472 );
    or g1981 ( n7401 , n4976 , n9930 );
    not g1982 ( n11587 , n30742 );
    or g1983 ( n14469 , n4314 , n17829 );
    or g1984 ( n30782 , n5743 , n35043 );
    and g1985 ( n23257 , n17035 , n26345 );
    or g1986 ( n14933 , n17417 , n22776 );
    and g1987 ( n14387 , n1417 , n2497 );
    and g1988 ( n14239 , n12361 , n18450 );
    nor g1989 ( n12491 , n31799 , n9926 );
    and g1990 ( n32718 , n36070 , n9824 );
    xnor g1991 ( n18658 , n5761 , n11781 );
    nor g1992 ( n32312 , n1564 , n18115 );
    or g1993 ( n1791 , n17568 , n28014 );
    xnor g1994 ( n31741 , n21030 , n22079 );
    xnor g1995 ( n3569 , n24985 , n26577 );
    or g1996 ( n35343 , n9658 , n7762 );
    xnor g1997 ( n20787 , n4113 , n31799 );
    xnor g1998 ( n22110 , n7779 , n4878 );
    not g1999 ( n24741 , n4962 );
    xnor g2000 ( n34296 , n7956 , n25611 );
    or g2001 ( n7352 , n5348 , n34225 );
    or g2002 ( n1927 , n26632 , n12996 );
    or g2003 ( n15355 , n12485 , n4952 );
    not g2004 ( n32842 , n10266 );
    and g2005 ( n2323 , n28209 , n30668 );
    xnor g2006 ( n7542 , n5095 , n27760 );
    and g2007 ( n14059 , n3801 , n9727 );
    nor g2008 ( n442 , n30525 , n4722 );
    not g2009 ( n15790 , n8432 );
    nor g2010 ( n29272 , n29693 , n6548 );
    or g2011 ( n33805 , n1683 , n21126 );
    and g2012 ( n16304 , n10507 , n35517 );
    nor g2013 ( n40 , n16946 , n6800 );
    or g2014 ( n22016 , n24414 , n19890 );
    xnor g2015 ( n11111 , n17771 , n19551 );
    or g2016 ( n3515 , n8338 , n35205 );
    or g2017 ( n13408 , n3347 , n21977 );
    or g2018 ( n25646 , n24552 , n6459 );
    xnor g2019 ( n26033 , n31625 , n12826 );
    or g2020 ( n16291 , n23992 , n32197 );
    xnor g2021 ( n20752 , n33999 , n33685 );
    and g2022 ( n34530 , n6811 , n34617 );
    nor g2023 ( n11171 , n25602 , n31906 );
    and g2024 ( n28927 , n34594 , n5682 );
    and g2025 ( n31677 , n13003 , n17485 );
    nor g2026 ( n23870 , n9929 , n13426 );
    or g2027 ( n31515 , n26876 , n6091 );
    nor g2028 ( n15785 , n4878 , n22399 );
    not g2029 ( n16863 , n1942 );
    or g2030 ( n8034 , n35390 , n18510 );
    xnor g2031 ( n7623 , n35933 , n3205 );
    xnor g2032 ( n33518 , n26461 , n11497 );
    and g2033 ( n19997 , n35889 , n28068 );
    and g2034 ( n21045 , n19832 , n9134 );
    xnor g2035 ( n1698 , n9734 , n5287 );
    xnor g2036 ( n29709 , n1349 , n10550 );
    or g2037 ( n9221 , n19984 , n12351 );
    or g2038 ( n24223 , n30975 , n1942 );
    xnor g2039 ( n20880 , n32217 , n3946 );
    or g2040 ( n3709 , n30098 , n11646 );
    nor g2041 ( n25302 , n24228 , n7453 );
    or g2042 ( n17198 , n2224 , n10915 );
    and g2043 ( n34610 , n13442 , n26227 );
    or g2044 ( n34601 , n31289 , n17812 );
    or g2045 ( n34729 , n9901 , n30127 );
    or g2046 ( n9402 , n26792 , n33764 );
    not g2047 ( n28213 , n2010 );
    and g2048 ( n30780 , n34227 , n34126 );
    xnor g2049 ( n10728 , n6199 , n32563 );
    or g2050 ( n7317 , n35927 , n3362 );
    and g2051 ( n28385 , n4034 , n16978 );
    nor g2052 ( n12103 , n1396 , n22628 );
    and g2053 ( n2825 , n7970 , n22478 );
    or g2054 ( n29555 , n26119 , n27907 );
    xnor g2055 ( n24413 , n17435 , n17568 );
    xnor g2056 ( n14449 , n1691 , n19187 );
    or g2057 ( n15866 , n8719 , n11312 );
    and g2058 ( n18558 , n31160 , n16551 );
    not g2059 ( n35358 , n19746 );
    xnor g2060 ( n23070 , n28941 , n10894 );
    or g2061 ( n8284 , n23754 , n31255 );
    nor g2062 ( n28334 , n3990 , n318 );
    or g2063 ( n29168 , n717 , n28751 );
    and g2064 ( n18962 , n20623 , n9271 );
    not g2065 ( n9479 , n31924 );
    and g2066 ( n7140 , n3965 , n35470 );
    xnor g2067 ( n3397 , n20460 , n9658 );
    nor g2068 ( n35214 , n31799 , n16249 );
    xnor g2069 ( n26754 , n32023 , n27381 );
    xnor g2070 ( n29822 , n12084 , n34625 );
    xnor g2071 ( n180 , n10288 , n32857 );
    xnor g2072 ( n33096 , n15509 , n35927 );
    or g2073 ( n2068 , n21411 , n28455 );
    and g2074 ( n21220 , n3678 , n21222 );
    or g2075 ( n25202 , n8544 , n4739 );
    and g2076 ( n27113 , n20892 , n11410 );
    and g2077 ( n9698 , n11753 , n541 );
    and g2078 ( n4841 , n13640 , n25114 );
    nor g2079 ( n7425 , n19551 , n27696 );
    buf g2080 ( n3979 , n5952 );
    or g2081 ( n23239 , n9658 , n20518 );
    or g2082 ( n19375 , n9385 , n5222 );
    nor g2083 ( n34718 , n3946 , n12775 );
    or g2084 ( n16067 , n25432 , n19435 );
    or g2085 ( n26602 , n453 , n25404 );
    or g2086 ( n33071 , n19557 , n5900 );
    or g2087 ( n33282 , n33886 , n1414 );
    xnor g2088 ( n31844 , n28133 , n11741 );
    xnor g2089 ( n18096 , n25379 , n24392 );
    and g2090 ( n3596 , n35711 , n14046 );
    or g2091 ( n8536 , n16620 , n17892 );
    not g2092 ( n26275 , n23918 );
    and g2093 ( n28995 , n459 , n398 );
    xnor g2094 ( n26519 , n9647 , n10894 );
    or g2095 ( n271 , n7265 , n3352 );
    and g2096 ( n10914 , n25186 , n8557 );
    and g2097 ( n18083 , n805 , n16656 );
    and g2098 ( n6538 , n4933 , n9515 );
    or g2099 ( n28577 , n5173 , n26023 );
    nor g2100 ( n2680 , n34118 , n3537 );
    or g2101 ( n10936 , n31089 , n5197 );
    xnor g2102 ( n32017 , n5106 , n32075 );
    or g2103 ( n31244 , n35404 , n25392 );
    and g2104 ( n4399 , n2668 , n16205 );
    not g2105 ( n2487 , n35770 );
    nor g2106 ( n16042 , n32973 , n282 );
    xnor g2107 ( n32234 , n28361 , n4962 );
    or g2108 ( n15588 , n4878 , n10076 );
    xnor g2109 ( n32629 , n25474 , n23399 );
    xnor g2110 ( n4638 , n19772 , n25174 );
    or g2111 ( n26400 , n4962 , n32719 );
    or g2112 ( n15571 , n6040 , n32572 );
    xnor g2113 ( n4151 , n17482 , n188 );
    xnor g2114 ( n32727 , n13333 , n14805 );
    or g2115 ( n15076 , n9658 , n26423 );
    not g2116 ( n3757 , n147 );
    or g2117 ( n17547 , n3205 , n32227 );
    or g2118 ( n19961 , n32095 , n247 );
    or g2119 ( n18199 , n4288 , n29661 );
    or g2120 ( n27610 , n9814 , n25350 );
    or g2121 ( n25540 , n21132 , n859 );
    and g2122 ( n7978 , n31607 , n5063 );
    and g2123 ( n3707 , n26107 , n22927 );
    and g2124 ( n15463 , n24913 , n23367 );
    xnor g2125 ( n24298 , n448 , n9789 );
    xnor g2126 ( n20746 , n20126 , n24371 );
    or g2127 ( n2476 , n31505 , n22682 );
    xnor g2128 ( n20404 , n3416 , n4878 );
    or g2129 ( n7412 , n6043 , n15164 );
    or g2130 ( n6187 , n22189 , n5164 );
    and g2131 ( n34174 , n9708 , n18708 );
    xnor g2132 ( n24311 , n4223 , n20909 );
    and g2133 ( n23819 , n34158 , n26118 );
    and g2134 ( n17302 , n25252 , n8464 );
    and g2135 ( n4507 , n3993 , n25787 );
    buf g2136 ( n19084 , n5784 );
    xnor g2137 ( n30943 , n25222 , n22172 );
    xnor g2138 ( n9949 , n21311 , n29839 );
    and g2139 ( n5949 , n19623 , n30315 );
    or g2140 ( n14049 , n28615 , n15796 );
    or g2141 ( n3074 , n34827 , n27704 );
    and g2142 ( n26267 , n18673 , n22904 );
    xnor g2143 ( n18738 , n14999 , n19721 );
    xnor g2144 ( n9388 , n27362 , n9658 );
    and g2145 ( n9427 , n19159 , n28730 );
    and g2146 ( n13792 , n8631 , n9519 );
    xnor g2147 ( n23888 , n19026 , n8549 );
    not g2148 ( n4919 , n22291 );
    or g2149 ( n33164 , n24579 , n27600 );
    not g2150 ( n18059 , n35244 );
    and g2151 ( n5794 , n10323 , n34215 );
    or g2152 ( n19022 , n4878 , n30233 );
    and g2153 ( n23489 , n10831 , n21442 );
    and g2154 ( n15987 , n14198 , n22476 );
    or g2155 ( n24692 , n19821 , n29626 );
    nor g2156 ( n3303 , n4878 , n13162 );
    xnor g2157 ( n28462 , n16775 , n30553 );
    nor g2158 ( n34427 , n1996 , n28574 );
    and g2159 ( n7964 , n8010 , n32047 );
    or g2160 ( n15203 , n19551 , n6512 );
    xnor g2161 ( n9279 , n19894 , n35412 );
    not g2162 ( n10542 , n10876 );
    nor g2163 ( n21173 , n21281 , n858 );
    nor g2164 ( n30791 , n29713 , n11245 );
    or g2165 ( n25676 , n26044 , n26468 );
    or g2166 ( n35932 , n13263 , n29267 );
    and g2167 ( n9819 , n29416 , n16746 );
    xnor g2168 ( n10533 , n16951 , n16620 );
    nor g2169 ( n10535 , n13973 , n10872 );
    and g2170 ( n4047 , n3098 , n8117 );
    xnor g2171 ( n22864 , n19693 , n2720 );
    or g2172 ( n11255 , n24044 , n33551 );
    or g2173 ( n10863 , n10737 , n13015 );
    xnor g2174 ( n25379 , n8026 , n8092 );
    nor g2175 ( n23484 , n35878 , n7019 );
    and g2176 ( n29499 , n28083 , n9029 );
    and g2177 ( n30689 , n1074 , n23473 );
    or g2178 ( n30412 , n17910 , n4478 );
    and g2179 ( n35977 , n33246 , n7148 );
    or g2180 ( n34993 , n8656 , n16919 );
    not g2181 ( n18013 , n35372 );
    not g2182 ( n35009 , n27297 );
    or g2183 ( n13483 , n19551 , n21193 );
    or g2184 ( n31270 , n15567 , n4478 );
    or g2185 ( n34936 , n17338 , n21870 );
    xnor g2186 ( n4597 , n3937 , n5619 );
    and g2187 ( n6735 , n28499 , n10223 );
    and g2188 ( n7342 , n25950 , n10938 );
    or g2189 ( n19903 , n866 , n1411 );
    not g2190 ( n3834 , n32526 );
    or g2191 ( n30439 , n29839 , n20344 );
    xnor g2192 ( n21795 , n34238 , n2977 );
    or g2193 ( n7264 , n4884 , n25953 );
    xnor g2194 ( n13497 , n7670 , n24371 );
    and g2195 ( n16288 , n26948 , n17130 );
    or g2196 ( n21763 , n9517 , n23187 );
    nor g2197 ( n2126 , n23514 , n16357 );
    nor g2198 ( n24465 , n26800 , n12143 );
    nor g2199 ( n25983 , n3254 , n17196 );
    or g2200 ( n8809 , n30008 , n3756 );
    and g2201 ( n3278 , n12994 , n15461 );
    xnor g2202 ( n16200 , n19012 , n9619 );
    not g2203 ( n12364 , n28733 );
    or g2204 ( n35857 , n15505 , n12464 );
    xnor g2205 ( n21590 , n24820 , n4288 );
    and g2206 ( n8623 , n19375 , n10196 );
    and g2207 ( n31125 , n34243 , n34728 );
    and g2208 ( n13732 , n22609 , n2158 );
    and g2209 ( n26342 , n27838 , n15405 );
    or g2210 ( n1456 , n346 , n25332 );
    or g2211 ( n26668 , n5036 , n4172 );
    and g2212 ( n19728 , n297 , n11043 );
    or g2213 ( n6871 , n6704 , n14554 );
    and g2214 ( n12053 , n2566 , n6536 );
    and g2215 ( n9792 , n16515 , n24062 );
    or g2216 ( n16010 , n9576 , n26659 );
    xnor g2217 ( n24477 , n13472 , n3273 );
    or g2218 ( n4343 , n6746 , n10762 );
    xnor g2219 ( n23703 , n10269 , n4962 );
    or g2220 ( n24642 , n23646 , n22783 );
    or g2221 ( n21768 , n31377 , n28438 );
    or g2222 ( n8248 , n4636 , n725 );
    or g2223 ( n6522 , n30932 , n5820 );
    nor g2224 ( n26380 , n32675 , n33031 );
    nor g2225 ( n15798 , n2583 , n1859 );
    not g2226 ( n15707 , n32095 );
    or g2227 ( n24217 , n24151 , n10872 );
    nor g2228 ( n7878 , n22291 , n24361 );
    or g2229 ( n34559 , n8209 , n21417 );
    and g2230 ( n22637 , n15026 , n2937 );
    or g2231 ( n9666 , n22697 , n3188 );
    xnor g2232 ( n33932 , n13862 , n15403 );
    or g2233 ( n29028 , n30806 , n544 );
    not g2234 ( n14383 , n25992 );
    or g2235 ( n12807 , n23929 , n12252 );
    and g2236 ( n16562 , n19753 , n32627 );
    xnor g2237 ( n7064 , n107 , n23726 );
    not g2238 ( n26174 , n17568 );
    xnor g2239 ( n29732 , n21677 , n17682 );
    and g2240 ( n24537 , n10148 , n28460 );
    and g2241 ( n550 , n6708 , n8667 );
    not g2242 ( n26032 , n10689 );
    and g2243 ( n26308 , n20007 , n20988 );
    nor g2244 ( n5671 , n13620 , n17711 );
    nor g2245 ( n3954 , n33199 , n1366 );
    nor g2246 ( n16111 , n32095 , n7572 );
    xnor g2247 ( n32890 , n26833 , n35927 );
    or g2248 ( n27510 , n17751 , n25414 );
    and g2249 ( n16874 , n19208 , n25409 );
    or g2250 ( n10413 , n35652 , n22961 );
    and g2251 ( n12453 , n6460 , n7850 );
    not g2252 ( n29920 , n34503 );
    xnor g2253 ( n2027 , n12545 , n8432 );
    xnor g2254 ( n30938 , n6384 , n19551 );
    or g2255 ( n3760 , n5335 , n30368 );
    or g2256 ( n777 , n3511 , n15344 );
    and g2257 ( n3701 , n35953 , n8047 );
    or g2258 ( n11984 , n34694 , n995 );
    or g2259 ( n25206 , n23872 , n29872 );
    or g2260 ( n15901 , n17292 , n29643 );
    or g2261 ( n9542 , n5335 , n22261 );
    or g2262 ( n17212 , n21410 , n7293 );
    nor g2263 ( n27284 , n15294 , n17450 );
    or g2264 ( n460 , n29939 , n19756 );
    and g2265 ( n33411 , n20063 , n15447 );
    and g2266 ( n28475 , n2486 , n24802 );
    and g2267 ( n19668 , n31689 , n20182 );
    or g2268 ( n11129 , n9793 , n26074 );
    or g2269 ( n1945 , n22672 , n10336 );
    xnor g2270 ( n968 , n30976 , n16566 );
    or g2271 ( n32325 , n4378 , n10986 );
    not g2272 ( n8582 , n23604 );
    or g2273 ( n10750 , n25616 , n31464 );
    or g2274 ( n23952 , n16922 , n33853 );
    or g2275 ( n3133 , n11533 , n26927 );
    and g2276 ( n2230 , n10467 , n13684 );
    xnor g2277 ( n23550 , n20678 , n3946 );
    or g2278 ( n4295 , n26928 , n15086 );
    or g2279 ( n30450 , n13271 , n5779 );
    xnor g2280 ( n5899 , n31194 , n35927 );
    or g2281 ( n9084 , n36046 , n11712 );
    not g2282 ( n1151 , n19551 );
    or g2283 ( n20737 , n12263 , n2042 );
    and g2284 ( n35657 , n21131 , n20020 );
    or g2285 ( n35391 , n19551 , n32370 );
    nor g2286 ( n28646 , n24128 , n9921 );
    or g2287 ( n3820 , n7540 , n575 );
    and g2288 ( n10860 , n9704 , n2316 );
    xnor g2289 ( n22100 , n9094 , n29988 );
    nor g2290 ( n15689 , n33470 , n4844 );
    or g2291 ( n24070 , n18216 , n16456 );
    or g2292 ( n2616 , n32095 , n5773 );
    or g2293 ( n19804 , n23888 , n5208 );
    nor g2294 ( n14110 , n26695 , n35545 );
    or g2295 ( n12472 , n830 , n2118 );
    or g2296 ( n11451 , n23270 , n30708 );
    or g2297 ( n25497 , n15050 , n32288 );
    and g2298 ( n1117 , n15647 , n23048 );
    nor g2299 ( n35535 , n33743 , n621 );
    or g2300 ( n15932 , n31043 , n11361 );
    and g2301 ( n18623 , n23656 , n6593 );
    or g2302 ( n21368 , n15464 , n12947 );
    xnor g2303 ( n18326 , n10425 , n32857 );
    xnor g2304 ( n22529 , n27550 , n19353 );
    and g2305 ( n1933 , n14360 , n13256 );
    or g2306 ( n2772 , n35085 , n33157 );
    xnor g2307 ( n14710 , n9725 , n31593 );
    or g2308 ( n28018 , n16990 , n23090 );
    and g2309 ( n31696 , n10156 , n10972 );
    and g2310 ( n7583 , n33589 , n20134 );
    nor g2311 ( n11711 , n15966 , n10490 );
    or g2312 ( n15205 , n10866 , n32932 );
    not g2313 ( n9554 , n30317 );
    or g2314 ( n26746 , n17518 , n21439 );
    and g2315 ( n3028 , n5819 , n2159 );
    and g2316 ( n21799 , n3524 , n10846 );
    or g2317 ( n9704 , n34913 , n21691 );
    xnor g2318 ( n6184 , n30337 , n3928 );
    not g2319 ( n6028 , n4878 );
    nor g2320 ( n28521 , n4288 , n1639 );
    and g2321 ( n26125 , n13892 , n10188 );
    or g2322 ( n2759 , n31289 , n9690 );
    xnor g2323 ( n12914 , n18527 , n31289 );
    and g2324 ( n677 , n24110 , n2796 );
    or g2325 ( n9914 , n31799 , n28457 );
    nor g2326 ( n2694 , n22844 , n18115 );
    xnor g2327 ( n14165 , n4673 , n23604 );
    or g2328 ( n22060 , n17522 , n24479 );
    or g2329 ( n221 , n9657 , n24025 );
    and g2330 ( n27783 , n8342 , n29351 );
    xor g2331 ( n9441 , n6505 , n8265 );
    or g2332 ( n4199 , n33658 , n591 );
    or g2333 ( n31835 , n22299 , n20748 );
    or g2334 ( n2151 , n17672 , n21162 );
    or g2335 ( n23806 , n31724 , n13493 );
    nor g2336 ( n18275 , n321 , n19387 );
    xnor g2337 ( n27215 , n6468 , n4878 );
    and g2338 ( n25858 , n27846 , n35735 );
    nor g2339 ( n16470 , n10074 , n17684 );
    or g2340 ( n31644 , n35128 , n15497 );
    xnor g2341 ( n8265 , n20815 , n16620 );
    or g2342 ( n20305 , n10063 , n2849 );
    or g2343 ( n29905 , n9761 , n13058 );
    or g2344 ( n26171 , n7739 , n28716 );
    or g2345 ( n24138 , n16922 , n31205 );
    and g2346 ( n28808 , n22603 , n35149 );
    or g2347 ( n27207 , n23059 , n35141 );
    and g2348 ( n10644 , n13569 , n33414 );
    or g2349 ( n5432 , n22888 , n9030 );
    and g2350 ( n23643 , n14334 , n5710 );
    or g2351 ( n33050 , n28485 , n29643 );
    nor g2352 ( n27719 , n15886 , n31275 );
    or g2353 ( n10938 , n1106 , n6374 );
    or g2354 ( n34625 , n34210 , n27174 );
    or g2355 ( n6896 , n3222 , n7200 );
    and g2356 ( n28356 , n15219 , n26133 );
    or g2357 ( n16235 , n10858 , n18395 );
    or g2358 ( n20781 , n13050 , n24479 );
    and g2359 ( n32772 , n27957 , n34569 );
    or g2360 ( n35872 , n14953 , n21659 );
    and g2361 ( n29006 , n20561 , n9353 );
    or g2362 ( n22018 , n4157 , n15144 );
    nor g2363 ( n11477 , n5071 , n11471 );
    and g2364 ( n16937 , n1636 , n4752 );
    xnor g2365 ( n15997 , n33411 , n11954 );
    and g2366 ( n22226 , n32583 , n19898 );
    xnor g2367 ( n8516 , n34983 , n30384 );
    or g2368 ( n20706 , n4288 , n15230 );
    xnor g2369 ( n3885 , n16671 , n19708 );
    not g2370 ( n4708 , n1079 );
    xnor g2371 ( n7223 , n28356 , n32095 );
    or g2372 ( n18068 , n5287 , n21562 );
    or g2373 ( n23982 , n26823 , n20797 );
    xnor g2374 ( n30637 , n8698 , n31252 );
    or g2375 ( n8773 , n11046 , n17756 );
    and g2376 ( n6509 , n22933 , n26484 );
    or g2377 ( n21166 , n11975 , n16608 );
    not g2378 ( n5912 , n2965 );
    and g2379 ( n10001 , n34658 , n4121 );
    or g2380 ( n8764 , n19984 , n21965 );
    and g2381 ( n196 , n29239 , n28689 );
    and g2382 ( n30034 , n23206 , n5722 );
    or g2383 ( n20254 , n29665 , n11878 );
    xnor g2384 ( n13446 , n5678 , n16152 );
    xnor g2385 ( n23577 , n4045 , n19551 );
    or g2386 ( n18460 , n8625 , n7883 );
    or g2387 ( n14884 , n13176 , n10862 );
    not g2388 ( n11078 , n35100 );
    nor g2389 ( n33474 , n24703 , n7784 );
    and g2390 ( n4065 , n20940 , n14722 );
    or g2391 ( n30847 , n34848 , n25594 );
    or g2392 ( n8199 , n13276 , n34852 );
    or g2393 ( n35065 , n31289 , n23177 );
    nor g2394 ( n25555 , n16620 , n22340 );
    not g2395 ( n6181 , n9975 );
    xnor g2396 ( n24665 , n25518 , n9053 );
    or g2397 ( n9302 , n2654 , n32507 );
    or g2398 ( n9805 , n5566 , n25831 );
    and g2399 ( n5580 , n14355 , n32901 );
    or g2400 ( n4894 , n9599 , n27724 );
    and g2401 ( n29058 , n15575 , n10055 );
    and g2402 ( n34607 , n3538 , n34078 );
    and g2403 ( n10341 , n24484 , n10105 );
    xnor g2404 ( n15619 , n26515 , n32095 );
    xnor g2405 ( n27530 , n33858 , n17434 );
    or g2406 ( n24466 , n19531 , n33443 );
    xnor g2407 ( n25455 , n12023 , n5663 );
    or g2408 ( n26657 , n5101 , n26002 );
    xnor g2409 ( n35419 , n31438 , n14077 );
    xnor g2410 ( n6143 , n11280 , n25405 );
    and g2411 ( n7831 , n29388 , n35120 );
    and g2412 ( n9809 , n11610 , n34823 );
    or g2413 ( n16122 , n4962 , n23052 );
    or g2414 ( n17414 , n28052 , n31184 );
    or g2415 ( n11400 , n28021 , n13215 );
    or g2416 ( n17137 , n28397 , n25255 );
    and g2417 ( n454 , n18725 , n24990 );
    not g2418 ( n13758 , n24240 );
    or g2419 ( n15224 , n18018 , n22858 );
    xnor g2420 ( n16936 , n32437 , n5287 );
    or g2421 ( n2200 , n33070 , n11640 );
    not g2422 ( n1485 , n3563 );
    xnor g2423 ( n13473 , n34608 , n36002 );
    and g2424 ( n32350 , n9805 , n21584 );
    or g2425 ( n8887 , n24371 , n1833 );
    or g2426 ( n35798 , n28628 , n18269 );
    xnor g2427 ( n30976 , n6348 , n24371 );
    xnor g2428 ( n21696 , n23878 , n18168 );
    or g2429 ( n1714 , n3046 , n24274 );
    and g2430 ( n32680 , n22698 , n24113 );
    not g2431 ( n29577 , n16083 );
    xnor g2432 ( n19064 , n24302 , n4878 );
    not g2433 ( n21921 , n5729 );
    xnor g2434 ( n34329 , n20818 , n20547 );
    and g2435 ( n8988 , n27323 , n9230 );
    or g2436 ( n5425 , n5206 , n17203 );
    or g2437 ( n14635 , n2252 , n17068 );
    xnor g2438 ( n7895 , n12712 , n6723 );
    xnor g2439 ( n6535 , n28208 , n31544 );
    or g2440 ( n3692 , n28123 , n2194 );
    not g2441 ( n29120 , n21405 );
    nor g2442 ( n6981 , n6759 , n6456 );
    xnor g2443 ( n3444 , n25637 , n3923 );
    not g2444 ( n7447 , n8668 );
    or g2445 ( n12918 , n23710 , n11996 );
    or g2446 ( n22478 , n17751 , n14943 );
    or g2447 ( n21623 , n27291 , n31038 );
    or g2448 ( n22830 , n30141 , n12413 );
    or g2449 ( n16730 , n16922 , n8191 );
    xnor g2450 ( n27292 , n1204 , n32857 );
    and g2451 ( n32735 , n9522 , n20056 );
    and g2452 ( n18949 , n24965 , n4547 );
    or g2453 ( n31873 , n25236 , n25447 );
    and g2454 ( n2451 , n13017 , n8518 );
    or g2455 ( n14153 , n32834 , n9915 );
    or g2456 ( n22696 , n32095 , n31538 );
    or g2457 ( n1309 , n28863 , n19267 );
    or g2458 ( n19316 , n6127 , n8392 );
    nor g2459 ( n23260 , n22818 , n24389 );
    or g2460 ( n28729 , n18870 , n19441 );
    or g2461 ( n20502 , n20125 , n20346 );
    and g2462 ( n7582 , n24238 , n27153 );
    or g2463 ( n5404 , n14290 , n34644 );
    xnor g2464 ( n8505 , n13796 , n3946 );
    and g2465 ( n18127 , n15560 , n28753 );
    nor g2466 ( n11197 , n27238 , n33796 );
    or g2467 ( n34077 , n4758 , n20506 );
    not g2468 ( n34260 , n20760 );
    and g2469 ( n23191 , n2353 , n1151 );
    and g2470 ( n26183 , n9887 , n29564 );
    and g2471 ( n30150 , n25509 , n16472 );
    or g2472 ( n21314 , n23531 , n29872 );
    nor g2473 ( n261 , n5635 , n4595 );
    nor g2474 ( n15021 , n27009 , n25347 );
    and g2475 ( n30608 , n30797 , n15758 );
    and g2476 ( n21627 , n33894 , n11139 );
    and g2477 ( n19394 , n15643 , n33375 );
    xnor g2478 ( n35242 , n14047 , n2223 );
    or g2479 ( n9616 , n16685 , n5779 );
    nor g2480 ( n31864 , n1751 , n27801 );
    nor g2481 ( n19219 , n19050 , n31411 );
    xnor g2482 ( n4080 , n18958 , n830 );
    not g2483 ( n13165 , n8326 );
    and g2484 ( n2132 , n33512 , n32334 );
    not g2485 ( n9511 , n30016 );
    xnor g2486 ( n3160 , n22952 , n12389 );
    xnor g2487 ( n14220 , n18102 , n32857 );
    nor g2488 ( n10364 , n35927 , n15209 );
    xnor g2489 ( n30308 , n7820 , n19705 );
    or g2490 ( n2677 , n9583 , n24643 );
    or g2491 ( n32920 , n13818 , n30287 );
    xnor g2492 ( n10268 , n12351 , n19984 );
    not g2493 ( n5990 , n1334 );
    not g2494 ( n11307 , n27561 );
    xor g2495 ( n28048 , n4192 , n33613 );
    or g2496 ( n34267 , n23176 , n26220 );
    and g2497 ( n6194 , n27324 , n34953 );
    and g2498 ( n22202 , n32035 , n32013 );
    or g2499 ( n906 , n4670 , n19336 );
    not g2500 ( n29752 , n9020 );
    xnor g2501 ( n35467 , n9247 , n22312 );
    or g2502 ( n21185 , n17756 , n12950 );
    or g2503 ( n33137 , n25978 , n11801 );
    xnor g2504 ( n30152 , n3229 , n30216 );
    not g2505 ( n17184 , n1528 );
    or g2506 ( n6599 , n3387 , n25036 );
    nor g2507 ( n30885 , n7540 , n20869 );
    and g2508 ( n3514 , n21253 , n15076 );
    and g2509 ( n34219 , n29042 , n15016 );
    or g2510 ( n11328 , n4900 , n1583 );
    xnor g2511 ( n15953 , n14593 , n9793 );
    or g2512 ( n18628 , n6832 , n2119 );
    nor g2513 ( n31735 , n420 , n8950 );
    or g2514 ( n31987 , n2431 , n16145 );
    xnor g2515 ( n7111 , n14769 , n18176 );
    and g2516 ( n21420 , n27862 , n26444 );
    or g2517 ( n29076 , n15403 , n33515 );
    and g2518 ( n35404 , n18497 , n23641 );
    xnor g2519 ( n26755 , n4335 , n11046 );
    and g2520 ( n16995 , n18368 , n17010 );
    xnor g2521 ( n30398 , n22030 , n30432 );
    or g2522 ( n29332 , n27291 , n12749 );
    or g2523 ( n206 , n4365 , n22823 );
    and g2524 ( n28396 , n20491 , n32131 );
    not g2525 ( n29098 , n15886 );
    nor g2526 ( n31797 , n35927 , n22274 );
    buf g2527 ( n9731 , n11240 );
    or g2528 ( n35285 , n14387 , n27501 );
    or g2529 ( n28301 , n19429 , n8098 );
    and g2530 ( n29048 , n23557 , n20614 );
    not g2531 ( n16611 , n34060 );
    nor g2532 ( n20326 , n8432 , n10418 );
    and g2533 ( n4785 , n506 , n27529 );
    or g2534 ( n22622 , n19471 , n28759 );
    and g2535 ( n31481 , n5686 , n5238 );
    and g2536 ( n20255 , n33747 , n3358 );
    not g2537 ( n28230 , n22200 );
    and g2538 ( n19099 , n16542 , n5340 );
    or g2539 ( n17847 , n29713 , n35555 );
    or g2540 ( n34736 , n24727 , n27813 );
    or g2541 ( n25237 , n29593 , n8924 );
    or g2542 ( n11086 , n15876 , n27973 );
    and g2543 ( n30423 , n12215 , n24387 );
    or g2544 ( n6195 , n21881 , n34811 );
    xnor g2545 ( n6100 , n20872 , n17568 );
    and g2546 ( n30109 , n16270 , n19411 );
    or g2547 ( n167 , n18847 , n9037 );
    and g2548 ( n16365 , n31842 , n3740 );
    nor g2549 ( n5061 , n2676 , n9071 );
    and g2550 ( n19866 , n567 , n35617 );
    or g2551 ( n15651 , n16258 , n30028 );
    or g2552 ( n22039 , n12487 , n34971 );
    or g2553 ( n7852 , n32285 , n19490 );
    or g2554 ( n8529 , n29884 , n12907 );
    and g2555 ( n6786 , n8363 , n8790 );
    or g2556 ( n1818 , n17431 , n16345 );
    or g2557 ( n27017 , n3205 , n27868 );
    and g2558 ( n18263 , n22203 , n28611 );
    or g2559 ( n522 , n22247 , n139 );
    or g2560 ( n2792 , n5224 , n17298 );
    or g2561 ( n26260 , n6939 , n3420 );
    xnor g2562 ( n1477 , n19038 , n17568 );
    or g2563 ( n10631 , n11919 , n29102 );
    and g2564 ( n27803 , n34416 , n1110 );
    and g2565 ( n3389 , n36062 , n23742 );
    or g2566 ( n12919 , n19551 , n35741 );
    or g2567 ( n30593 , n4268 , n3006 );
    nor g2568 ( n36024 , n16015 , n7648 );
    or g2569 ( n18069 , n22547 , n29953 );
    xnor g2570 ( n19936 , n10132 , n23546 );
    or g2571 ( n18288 , n29222 , n24115 );
    and g2572 ( n14129 , n14133 , n26073 );
    or g2573 ( n12308 , n4878 , n9379 );
    or g2574 ( n1685 , n9890 , n17612 );
    not g2575 ( n18679 , n5978 );
    or g2576 ( n33208 , n17568 , n13638 );
    and g2577 ( n28108 , n30984 , n26384 );
    and g2578 ( n4342 , n19109 , n17512 );
    xnor g2579 ( n11830 , n4449 , n6383 );
    and g2580 ( n2432 , n15390 , n213 );
    xnor g2581 ( n29904 , n22829 , n30767 );
    or g2582 ( n4092 , n6172 , n30646 );
    or g2583 ( n8115 , n12815 , n4203 );
    and g2584 ( n4889 , n29109 , n25427 );
    xnor g2585 ( n34113 , n29655 , n2392 );
    and g2586 ( n5160 , n34343 , n11658 );
    or g2587 ( n15322 , n21696 , n15496 );
    or g2588 ( n7471 , n3043 , n25423 );
    or g2589 ( n35134 , n23171 , n7303 );
    nor g2590 ( n7548 , n33856 , n982 );
    or g2591 ( n35723 , n10073 , n31887 );
    xnor g2592 ( n3332 , n424 , n29839 );
    or g2593 ( n711 , n26389 , n30091 );
    or g2594 ( n13146 , n9793 , n14990 );
    and g2595 ( n2148 , n5575 , n19987 );
    or g2596 ( n22716 , n8045 , n17974 );
    or g2597 ( n19370 , n27984 , n4478 );
    or g2598 ( n18056 , n28596 , n3184 );
    and g2599 ( n25201 , n25211 , n15524 );
    not g2600 ( n24034 , n4758 );
    and g2601 ( n27199 , n9224 , n31660 );
    and g2602 ( n27652 , n3207 , n34385 );
    or g2603 ( n2897 , n24985 , n15497 );
    and g2604 ( n12481 , n27610 , n30644 );
    or g2605 ( n21761 , n18664 , n5779 );
    xnor g2606 ( n16776 , n11572 , n20743 );
    xnor g2607 ( n5932 , n10454 , n17141 );
    xnor g2608 ( n2554 , n12743 , n8677 );
    xnor g2609 ( n24682 , n6122 , n34270 );
    xnor g2610 ( n31177 , n32546 , n6909 );
    or g2611 ( n1720 , n25792 , n16339 );
    and g2612 ( n22138 , n4831 , n840 );
    xnor g2613 ( n13153 , n18470 , n26457 );
    and g2614 ( n7204 , n23804 , n10454 );
    and g2615 ( n17153 , n27136 , n4168 );
    or g2616 ( n3293 , n4962 , n27250 );
    and g2617 ( n19734 , n1588 , n23114 );
    or g2618 ( n19737 , n21830 , n27887 );
    and g2619 ( n28065 , n19508 , n31562 );
    or g2620 ( n24075 , n27959 , n8153 );
    nor g2621 ( n32171 , n32095 , n17525 );
    or g2622 ( n12038 , n1950 , n14789 );
    or g2623 ( n6526 , n5503 , n11067 );
    or g2624 ( n23948 , n1466 , n10292 );
    and g2625 ( n17815 , n29228 , n9465 );
    or g2626 ( n11819 , n9793 , n20061 );
    and g2627 ( n33396 , n21110 , n15587 );
    or g2628 ( n5320 , n11390 , n21239 );
    or g2629 ( n3872 , n14619 , n25392 );
    xnor g2630 ( n24460 , n16750 , n31272 );
    and g2631 ( n20987 , n31959 , n4027 );
    or g2632 ( n35496 , n27123 , n3979 );
    and g2633 ( n22499 , n18435 , n12110 );
    or g2634 ( n6045 , n31272 , n18348 );
    xnor g2635 ( n6539 , n1340 , n1950 );
    or g2636 ( n35073 , n30742 , n28981 );
    xnor g2637 ( n8037 , n35967 , n22291 );
    or g2638 ( n5199 , n1221 , n12128 );
    or g2639 ( n9903 , n9986 , n26143 );
    or g2640 ( n18966 , n3739 , n2386 );
    or g2641 ( n35320 , n2128 , n15497 );
    or g2642 ( n26721 , n23640 , n5457 );
    xnor g2643 ( n33995 , n8234 , n13492 );
    not g2644 ( n4874 , n4526 );
    or g2645 ( n6876 , n10564 , n26220 );
    and g2646 ( n6286 , n5576 , n2266 );
    or g2647 ( n34180 , n35927 , n11091 );
    xnor g2648 ( n34612 , n849 , n27291 );
    buf g2649 ( n26659 , n28539 );
    nor g2650 ( n4552 , n10894 , n16671 );
    xnor g2651 ( n5259 , n32469 , n10894 );
    or g2652 ( n11591 , n13791 , n22946 );
    and g2653 ( n10620 , n16241 , n4451 );
    and g2654 ( n22879 , n22019 , n16352 );
    or g2655 ( n23882 , n3222 , n13678 );
    xnor g2656 ( n21337 , n16186 , n23456 );
    or g2657 ( n455 , n20450 , n6712 );
    and g2658 ( n17711 , n35275 , n16599 );
    xnor g2659 ( n22275 , n17542 , n33448 );
    nor g2660 ( n29283 , n32857 , n33245 );
    or g2661 ( n28944 , n28188 , n14841 );
    and g2662 ( n1403 , n32151 , n7356 );
    and g2663 ( n174 , n20412 , n13310 );
    xnor g2664 ( n13138 , n29994 , n3222 );
    xnor g2665 ( n28637 , n35553 , n1950 );
    or g2666 ( n24722 , n24940 , n8366 );
    xnor g2667 ( n20215 , n29586 , n9551 );
    or g2668 ( n25859 , n12794 , n13541 );
    or g2669 ( n25967 , n22533 , n31549 );
    or g2670 ( n16551 , n5412 , n17337 );
    or g2671 ( n7077 , n19551 , n27804 );
    not g2672 ( n19036 , n4350 );
    or g2673 ( n19238 , n9184 , n16399 );
    and g2674 ( n20044 , n10169 , n17290 );
    nor g2675 ( n24720 , n16922 , n27601 );
    or g2676 ( n11200 , n29135 , n9162 );
    xnor g2677 ( n972 , n13409 , n15894 );
    and g2678 ( n28023 , n21577 , n14213 );
    and g2679 ( n19281 , n20523 , n18331 );
    or g2680 ( n6669 , n22434 , n33125 );
    not g2681 ( n35281 , n8230 );
    and g2682 ( n5627 , n29996 , n9374 );
    and g2683 ( n21169 , n16260 , n12335 );
    or g2684 ( n14111 , n21950 , n18749 );
    not g2685 ( n30767 , n24371 );
    and g2686 ( n30804 , n18608 , n16977 );
    or g2687 ( n23416 , n12018 , n1060 );
    nor g2688 ( n18680 , n4878 , n27746 );
    and g2689 ( n6685 , n27661 , n20860 );
    or g2690 ( n31493 , n7245 , n15757 );
    or g2691 ( n3970 , n12282 , n17964 );
    and g2692 ( n14485 , n25237 , n13589 );
    not g2693 ( n3090 , n10840 );
    and g2694 ( n11802 , n8837 , n17309 );
    xnor g2695 ( n35972 , n2443 , n13563 );
    or g2696 ( n3283 , n25139 , n33416 );
    and g2697 ( n6721 , n19356 , n8622 );
    not g2698 ( n34013 , n31472 );
    nor g2699 ( n13991 , n21706 , n26590 );
    nor g2700 ( n18214 , n35817 , n32562 );
    or g2701 ( n8894 , n35267 , n1856 );
    xnor g2702 ( n18500 , n25994 , n5431 );
    xnor g2703 ( n4004 , n21502 , n8432 );
    xnor g2704 ( n32326 , n11014 , n3627 );
    xnor g2705 ( n36034 , n25918 , n17568 );
    not g2706 ( n9146 , n29839 );
    and g2707 ( n16752 , n32800 , n9419 );
    xnor g2708 ( n35267 , n31551 , n5147 );
    xnor g2709 ( n9296 , n10514 , n17384 );
    nor g2710 ( n23282 , n10581 , n21240 );
    or g2711 ( n34033 , n4154 , n16919 );
    or g2712 ( n22015 , n8340 , n19732 );
    xnor g2713 ( n28776 , n21861 , n26718 );
    nor g2714 ( n3399 , n22291 , n2217 );
    and g2715 ( n29800 , n18997 , n27945 );
    or g2716 ( n17530 , n21209 , n6075 );
    xnor g2717 ( n22149 , n13624 , n12987 );
    xnor g2718 ( n357 , n29637 , n387 );
    or g2719 ( n26810 , n12234 , n20866 );
    nor g2720 ( n10856 , n15886 , n14299 );
    or g2721 ( n35461 , n2619 , n20797 );
    or g2722 ( n17523 , n5283 , n12596 );
    xnor g2723 ( n21069 , n29631 , n30742 );
    or g2724 ( n15652 , n15044 , n26815 );
    or g2725 ( n6246 , n15359 , n23921 );
    nor g2726 ( n26642 , n21523 , n25695 );
    xnor g2727 ( n19712 , n33604 , n4288 );
    and g2728 ( n30520 , n27702 , n1303 );
    not g2729 ( n2496 , n16568 );
    xnor g2730 ( n31141 , n5190 , n19984 );
    and g2731 ( n4681 , n17774 , n4960 );
    or g2732 ( n20382 , n1485 , n30604 );
    or g2733 ( n22796 , n9793 , n14099 );
    or g2734 ( n29781 , n18784 , n24479 );
    or g2735 ( n30122 , n1992 , n7448 );
    or g2736 ( n26142 , n31867 , n7344 );
    xnor g2737 ( n8407 , n3171 , n26972 );
    xor g2738 ( n17119 , n8454 , n4359 );
    xor g2739 ( n6990 , n1455 , n7528 );
    or g2740 ( n31030 , n31799 , n11488 );
    or g2741 ( n12945 , n35681 , n13161 );
    and g2742 ( n319 , n28458 , n11903 );
    not g2743 ( n14112 , n8869 );
    or g2744 ( n12343 , n16973 , n12428 );
    and g2745 ( n29589 , n30014 , n12356 );
    or g2746 ( n10187 , n33803 , n27625 );
    or g2747 ( n1887 , n16922 , n24759 );
    and g2748 ( n10709 , n31201 , n15407 );
    or g2749 ( n32035 , n25448 , n15290 );
    or g2750 ( n11082 , n29713 , n30107 );
    and g2751 ( n28208 , n35655 , n7633 );
    nor g2752 ( n19197 , n28266 , n33956 );
    and g2753 ( n32260 , n35577 , n10993 );
    or g2754 ( n20401 , n11266 , n21723 );
    and g2755 ( n1063 , n21163 , n22554 );
    and g2756 ( n12259 , n25886 , n15554 );
    and g2757 ( n24552 , n22587 , n2993 );
    or g2758 ( n7116 , n15178 , n8360 );
    xor g2759 ( n13679 , n19515 , n34786 );
    or g2760 ( n23371 , n4960 , n35732 );
    or g2761 ( n31171 , n26291 , n27704 );
    xnor g2762 ( n32639 , n19858 , n4774 );
    xnor g2763 ( n24430 , n22400 , n8405 );
    and g2764 ( n4749 , n19055 , n20826 );
    nor g2765 ( n11364 , n35753 , n35696 );
    xnor g2766 ( n18572 , n18937 , n10235 );
    not g2767 ( n11607 , n24996 );
    and g2768 ( n18377 , n33549 , n33861 );
    or g2769 ( n32987 , n30878 , n2613 );
    or g2770 ( n11875 , n3222 , n29994 );
    or g2771 ( n22140 , n3222 , n26622 );
    or g2772 ( n19111 , n22540 , n11499 );
    and g2773 ( n12288 , n11549 , n10095 );
    or g2774 ( n20275 , n24934 , n13480 );
    nor g2775 ( n4303 , n31126 , n20467 );
    or g2776 ( n9577 , n28086 , n31946 );
    or g2777 ( n6313 , n3750 , n17046 );
    and g2778 ( n18219 , n20080 , n31468 );
    and g2779 ( n15266 , n27331 , n15059 );
    not g2780 ( n34699 , n14727 );
    and g2781 ( n25499 , n29312 , n10226 );
    and g2782 ( n1810 , n26233 , n13539 );
    nor g2783 ( n6804 , n20093 , n29203 );
    xnor g2784 ( n27865 , n14117 , n12321 );
    and g2785 ( n421 , n1361 , n25333 );
    and g2786 ( n20484 , n31092 , n34198 );
    and g2787 ( n25812 , n24009 , n3222 );
    xnor g2788 ( n4276 , n348 , n35927 );
    xnor g2789 ( n13690 , n8528 , n489 );
    and g2790 ( n3679 , n8596 , n7737 );
    xnor g2791 ( n4709 , n31276 , n6397 );
    or g2792 ( n5946 , n17052 , n13967 );
    not g2793 ( n13084 , n34476 );
    and g2794 ( n27231 , n27338 , n30086 );
    or g2795 ( n7067 , n21598 , n34537 );
    and g2796 ( n7115 , n31427 , n13471 );
    nor g2797 ( n9998 , n3687 , n19432 );
    or g2798 ( n13032 , n4797 , n19732 );
    nor g2799 ( n9772 , n9318 , n23149 );
    xnor g2800 ( n19205 , n31433 , n22291 );
    xnor g2801 ( n7217 , n25584 , n11074 );
    and g2802 ( n31083 , n6794 , n7984 );
    or g2803 ( n18071 , n33129 , n34727 );
    and g2804 ( n21313 , n12596 , n10147 );
    xnor g2805 ( n9735 , n15818 , n33196 );
    or g2806 ( n33994 , n9658 , n13177 );
    or g2807 ( n28237 , n22598 , n14356 );
    or g2808 ( n7143 , n22291 , n31109 );
    or g2809 ( n6426 , n12007 , n4478 );
    xnor g2810 ( n2305 , n6500 , n31006 );
    xnor g2811 ( n13020 , n3596 , n31215 );
    xnor g2812 ( n22567 , n18815 , n7469 );
    or g2813 ( n16883 , n9789 , n15658 );
    or g2814 ( n33576 , n24371 , n30944 );
    xnor g2815 ( n29145 , n17288 , n12357 );
    xnor g2816 ( n34813 , n16093 , n3725 );
    nor g2817 ( n12399 , n1305 , n33416 );
    or g2818 ( n10198 , n8432 , n16048 );
    and g2819 ( n17346 , n27013 , n4118 );
    not g2820 ( n15743 , n9361 );
    xnor g2821 ( n1974 , n16654 , n9520 );
    and g2822 ( n19687 , n25036 , n108 );
    xnor g2823 ( n35573 , n35034 , n22315 );
    and g2824 ( n15962 , n28115 , n7266 );
    or g2825 ( n12777 , n18757 , n27801 );
    and g2826 ( n33864 , n2428 , n6949 );
    or g2827 ( n400 , n15498 , n17905 );
    or g2828 ( n9098 , n3946 , n28917 );
    or g2829 ( n16682 , n12345 , n12128 );
    and g2830 ( n35374 , n27314 , n27762 );
    xnor g2831 ( n27379 , n8804 , n17568 );
    xnor g2832 ( n10843 , n31302 , n30742 );
    not g2833 ( n6323 , n35848 );
    or g2834 ( n27677 , n5287 , n13565 );
    not g2835 ( n15623 , n30742 );
    xnor g2836 ( n20539 , n5631 , n7571 );
    or g2837 ( n11972 , n12424 , n30287 );
    or g2838 ( n12395 , n13624 , n12987 );
    xnor g2839 ( n2674 , n21392 , n11455 );
    nor g2840 ( n21583 , n4878 , n23133 );
    not g2841 ( n2549 , n16620 );
    not g2842 ( n419 , n456 );
    or g2843 ( n17728 , n24326 , n23939 );
    or g2844 ( n13456 , n1750 , n8185 );
    xnor g2845 ( n32463 , n14275 , n31559 );
    or g2846 ( n22239 , n31799 , n12653 );
    xnor g2847 ( n19850 , n900 , n32715 );
    and g2848 ( n2717 , n32956 , n16720 );
    or g2849 ( n18302 , n17786 , n2621 );
    and g2850 ( n21354 , n29450 , n5750 );
    or g2851 ( n25321 , n34762 , n1942 );
    or g2852 ( n8073 , n34793 , n32259 );
    xnor g2853 ( n3994 , n11015 , n9025 );
    or g2854 ( n3684 , n31272 , n365 );
    and g2855 ( n7679 , n35798 , n28535 );
    or g2856 ( n25462 , n30232 , n26220 );
    or g2857 ( n30552 , n32857 , n296 );
    xnor g2858 ( n5091 , n5739 , n10901 );
    xnor g2859 ( n12019 , n32911 , n1430 );
    xnor g2860 ( n21425 , n28393 , n27402 );
    nor g2861 ( n22298 , n25602 , n1891 );
    or g2862 ( n820 , n11455 , n32580 );
    or g2863 ( n30044 , n8926 , n34373 );
    not g2864 ( n27989 , n32637 );
    xnor g2865 ( n1313 , n34535 , n31251 );
    xnor g2866 ( n203 , n29614 , n9793 );
    or g2867 ( n20943 , n35323 , n7673 );
    xor g2868 ( n35739 , n32620 , n28794 );
    not g2869 ( n12666 , n26263 );
    or g2870 ( n25246 , n14915 , n25099 );
    or g2871 ( n5583 , n15170 , n28675 );
    not g2872 ( n25404 , n25392 );
    or g2873 ( n18368 , n16265 , n15172 );
    or g2874 ( n11624 , n5287 , n32437 );
    xnor g2875 ( n7239 , n3924 , n10373 );
    xnor g2876 ( n4969 , n25113 , n16321 );
    and g2877 ( n9482 , n1542 , n4992 );
    or g2878 ( n32353 , n29862 , n18371 );
    not g2879 ( n9860 , n4288 );
    xnor g2880 ( n29888 , n31415 , n18930 );
    or g2881 ( n17149 , n10894 , n5855 );
    xnor g2882 ( n14520 , n28809 , n35374 );
    or g2883 ( n4397 , n2277 , n24292 );
    and g2884 ( n3099 , n27023 , n6641 );
    xnor g2885 ( n19201 , n28561 , n22517 );
    not g2886 ( n2472 , n17568 );
    not g2887 ( n20239 , n12053 );
    or g2888 ( n26000 , n14267 , n15439 );
    xnor g2889 ( n14084 , n1155 , n33863 );
    not g2890 ( n29052 , n9361 );
    or g2891 ( n12085 , n32916 , n28404 );
    xnor g2892 ( n28833 , n11378 , n27635 );
    or g2893 ( n3952 , n20872 , n8392 );
    or g2894 ( n33502 , n33669 , n19861 );
    or g2895 ( n18980 , n15886 , n33357 );
    xnor g2896 ( n8711 , n2208 , n24498 );
    or g2897 ( n30465 , n32857 , n35494 );
    or g2898 ( n9466 , n2072 , n29033 );
    and g2899 ( n16285 , n14060 , n33230 );
    xnor g2900 ( n6970 , n22330 , n31960 );
    xnor g2901 ( n26624 , n35854 , n30742 );
    not g2902 ( n5701 , n16620 );
    or g2903 ( n7690 , n2259 , n18794 );
    or g2904 ( n27374 , n9309 , n13217 );
    xnor g2905 ( n12247 , n25317 , n4962 );
    or g2906 ( n35407 , n22664 , n33781 );
    nor g2907 ( n30383 , n11997 , n4076 );
    or g2908 ( n27132 , n19059 , n27590 );
    and g2909 ( n23701 , n9746 , n27478 );
    xnor g2910 ( n28913 , n25312 , n31370 );
    and g2911 ( n10839 , n31876 , n22179 );
    and g2912 ( n9020 , n35908 , n27222 );
    or g2913 ( n14772 , n35927 , n1312 );
    or g2914 ( n32971 , n27505 , n5868 );
    xnor g2915 ( n12014 , n34424 , n13062 );
    and g2916 ( n15272 , n21667 , n8235 );
    or g2917 ( n15970 , n17300 , n27501 );
    and g2918 ( n28219 , n28612 , n13700 );
    and g2919 ( n28636 , n12992 , n32523 );
    xnor g2920 ( n19897 , n23063 , n13786 );
    or g2921 ( n207 , n32858 , n11224 );
    xnor g2922 ( n12748 , n18099 , n29713 );
    not g2923 ( n13088 , n16980 );
    or g2924 ( n71 , n26915 , n26931 );
    or g2925 ( n23749 , n606 , n25262 );
    xnor g2926 ( n19459 , n21590 , n12499 );
    not g2927 ( n5475 , n28603 );
    nor g2928 ( n14360 , n29468 , n16642 );
    or g2929 ( n15504 , n21063 , n26002 );
    or g2930 ( n13184 , n12684 , n32441 );
    and g2931 ( n6439 , n32236 , n12484 );
    or g2932 ( n14248 , n7104 , n26365 );
    xor g2933 ( n31189 , n35710 , n14217 );
    or g2934 ( n28140 , n9793 , n555 );
    or g2935 ( n1401 , n35870 , n32038 );
    or g2936 ( n18854 , n26115 , n20300 );
    xnor g2937 ( n13577 , n13790 , n28246 );
    not g2938 ( n35339 , n16594 );
    xnor g2939 ( n30664 , n18558 , n22291 );
    and g2940 ( n8472 , n34200 , n35391 );
    xnor g2941 ( n21986 , n15005 , n17568 );
    xnor g2942 ( n25109 , n22844 , n15676 );
    xnor g2943 ( n4427 , n23212 , n29713 );
    and g2944 ( n22679 , n21007 , n15650 );
    nor g2945 ( n9966 , n6665 , n7198 );
    nor g2946 ( n4066 , n3810 , n29062 );
    xnor g2947 ( n15183 , n28066 , n7540 );
    not g2948 ( n13643 , n31712 );
    or g2949 ( n27131 , n7932 , n29411 );
    not g2950 ( n19601 , n29370 );
    or g2951 ( n19321 , n16339 , n8839 );
    and g2952 ( n27592 , n33696 , n6239 );
    and g2953 ( n10125 , n34211 , n35138 );
    or g2954 ( n6642 , n14438 , n21691 );
    nor g2955 ( n32053 , n11046 , n17565 );
    xnor g2956 ( n34568 , n1619 , n3205 );
    nor g2957 ( n22067 , n31996 , n29203 );
    xnor g2958 ( n10044 , n34762 , n4878 );
    xnor g2959 ( n298 , n6051 , n830 );
    xnor g2960 ( n8258 , n30186 , n2491 );
    and g2961 ( n7347 , n7426 , n27480 );
    nor g2962 ( n17721 , n7540 , n19476 );
    and g2963 ( n22997 , n24726 , n2368 );
    xnor g2964 ( n22418 , n20043 , n1165 );
    or g2965 ( n23180 , n21820 , n17314 );
    xnor g2966 ( n15996 , n31393 , n3434 );
    or g2967 ( n21187 , n11683 , n25786 );
    or g2968 ( n33710 , n35741 , n8392 );
    not g2969 ( n31744 , n4962 );
    nor g2970 ( n13785 , n13419 , n31514 );
    or g2971 ( n29724 , n819 , n6374 );
    or g2972 ( n20187 , n35299 , n35217 );
    and g2973 ( n11354 , n2249 , n1062 );
    buf g2974 ( n23187 , n4772 );
    nor g2975 ( n10253 , n21922 , n17968 );
    not g2976 ( n35631 , n5335 );
    not g2977 ( n13455 , n11996 );
    xnor g2978 ( n7985 , n683 , n822 );
    and g2979 ( n8197 , n9322 , n4408 );
    or g2980 ( n8449 , n7540 , n3876 );
    and g2981 ( n26856 , n35087 , n33431 );
    or g2982 ( n2623 , n6115 , n17162 );
    xnor g2983 ( n10012 , n13701 , n19866 );
    and g2984 ( n27232 , n25010 , n279 );
    and g2985 ( n27658 , n3982 , n18825 );
    or g2986 ( n34748 , n17568 , n23334 );
    or g2987 ( n16276 , n15846 , n1715 );
    nor g2988 ( n34602 , n12916 , n18115 );
    not g2989 ( n29854 , n3805 );
    xnor g2990 ( n34004 , n17571 , n18882 );
    not g2991 ( n12794 , n29353 );
    xnor g2992 ( n3636 , n14211 , n16620 );
    and g2993 ( n23278 , n6633 , n21921 );
    xnor g2994 ( n28188 , n33704 , n25789 );
    or g2995 ( n33165 , n27226 , n17682 );
    or g2996 ( n7862 , n25159 , n18488 );
    xnor g2997 ( n19973 , n31874 , n3640 );
    and g2998 ( n17701 , n12071 , n22411 );
    xnor g2999 ( n9655 , n22821 , n28511 );
    and g3000 ( n6995 , n4591 , n1335 );
    or g3001 ( n2703 , n31884 , n2057 );
    and g3002 ( n16536 , n2286 , n4166 );
    xnor g3003 ( n10097 , n34053 , n19451 );
    not g3004 ( n22417 , n22369 );
    not g3005 ( n31707 , n33611 );
    not g3006 ( n26388 , n21624 );
    and g3007 ( n14655 , n10342 , n1886 );
    and g3008 ( n27470 , n20599 , n26470 );
    or g3009 ( n10156 , n8534 , n31550 );
    xnor g3010 ( n9652 , n34606 , n24673 );
    or g3011 ( n931 , n10894 , n18801 );
    or g3012 ( n31343 , n16725 , n26124 );
    or g3013 ( n7855 , n4960 , n14788 );
    not g3014 ( n2826 , n27039 );
    nor g3015 ( n28285 , n25311 , n22293 );
    and g3016 ( n30025 , n21646 , n27368 );
    or g3017 ( n17949 , n19879 , n27973 );
    and g3018 ( n18192 , n2779 , n6899 );
    or g3019 ( n20777 , n11015 , n9025 );
    and g3020 ( n14184 , n11556 , n32462 );
    and g3021 ( n29453 , n12304 , n21769 );
    or g3022 ( n12350 , n25602 , n22180 );
    or g3023 ( n23523 , n367 , n9194 );
    or g3024 ( n34122 , n25208 , n12791 );
    nor g3025 ( n23663 , n11618 , n3106 );
    buf g3026 ( n16345 , n3243 );
    xnor g3027 ( n35491 , n22255 , n24371 );
    xnor g3028 ( n35019 , n31460 , n22522 );
    or g3029 ( n12291 , n10620 , n3738 );
    or g3030 ( n27714 , n21440 , n3805 );
    or g3031 ( n28371 , n19551 , n21213 );
    or g3032 ( n18243 , n28608 , n4254 );
    xnor g3033 ( n5739 , n14437 , n15403 );
    xnor g3034 ( n19148 , n8311 , n4288 );
    and g3035 ( n28135 , n32646 , n27951 );
    and g3036 ( n32259 , n9968 , n30301 );
    or g3037 ( n17001 , n5366 , n35402 );
    and g3038 ( n25272 , n23806 , n21897 );
    xnor g3039 ( n13280 , n23040 , n17751 );
    and g3040 ( n12797 , n21743 , n6602 );
    or g3041 ( n7686 , n13961 , n3307 );
    or g3042 ( n26434 , n32452 , n25355 );
    not g3043 ( n22071 , n591 );
    or g3044 ( n8811 , n14999 , n19721 );
    xnor g3045 ( n23035 , n24537 , n23604 );
    xnor g3046 ( n9599 , n27309 , n32857 );
    or g3047 ( n26392 , n20687 , n19084 );
    xnor g3048 ( n22822 , n1505 , n17568 );
    or g3049 ( n19193 , n786 , n11601 );
    or g3050 ( n33664 , n12517 , n3239 );
    or g3051 ( n32456 , n32095 , n9373 );
    or g3052 ( n6964 , n3536 , n30200 );
    or g3053 ( n22196 , n26126 , n28866 );
    or g3054 ( n5792 , n4962 , n1352 );
    xnor g3055 ( n6481 , n7229 , n31559 );
    not g3056 ( n25713 , n29713 );
    or g3057 ( n26977 , n31559 , n25174 );
    nor g3058 ( n26488 , n35927 , n19628 );
    or g3059 ( n7486 , n14481 , n23626 );
    or g3060 ( n30300 , n5955 , n3842 );
    and g3061 ( n10878 , n21670 , n3074 );
    and g3062 ( n16744 , n11486 , n7450 );
    xnor g3063 ( n13592 , n32133 , n22291 );
    xnor g3064 ( n19269 , n9333 , n7567 );
    xnor g3065 ( n20610 , n27332 , n17865 );
    and g3066 ( n22217 , n7042 , n8007 );
    xnor g3067 ( n17492 , n12406 , n13906 );
    xnor g3068 ( n27549 , n10450 , n12705 );
    and g3069 ( n8766 , n8046 , n15236 );
    not g3070 ( n30870 , n34865 );
    or g3071 ( n22148 , n688 , n908 );
    and g3072 ( n3751 , n10343 , n5860 );
    or g3073 ( n10327 , n33417 , n4033 );
    or g3074 ( n24661 , n19249 , n26659 );
    nor g3075 ( n22543 , n7482 , n30159 );
    and g3076 ( n12702 , n5288 , n26820 );
    or g3077 ( n14806 , n10894 , n15982 );
    and g3078 ( n301 , n11707 , n21855 );
    xnor g3079 ( n28568 , n11672 , n7540 );
    and g3080 ( n4561 , n6771 , n8828 );
    xnor g3081 ( n35397 , n21774 , n32095 );
    and g3082 ( n29317 , n31754 , n11183 );
    or g3083 ( n5185 , n33990 , n62 );
    xnor g3084 ( n18118 , n8654 , n13132 );
    or g3085 ( n7358 , n27954 , n18712 );
    xnor g3086 ( n35104 , n15298 , n25602 );
    or g3087 ( n10708 , n16851 , n6075 );
    and g3088 ( n34018 , n28251 , n32813 );
    and g3089 ( n27679 , n15993 , n15960 );
    xnor g3090 ( n34238 , n8980 , n5287 );
    or g3091 ( n34880 , n17169 , n1942 );
    or g3092 ( n18802 , n26960 , n21379 );
    and g3093 ( n8950 , n19417 , n24440 );
    nor g3094 ( n14633 , n11264 , n9921 );
    not g3095 ( n7700 , n31411 );
    xnor g3096 ( n19813 , n1939 , n4871 );
    xnor g3097 ( n24136 , n21404 , n25602 );
    or g3098 ( n20634 , n24332 , n5565 );
    and g3099 ( n33642 , n31328 , n31154 );
    nor g3100 ( n17940 , n30742 , n31793 );
    or g3101 ( n22046 , n21613 , n34727 );
    and g3102 ( n511 , n31600 , n25046 );
    or g3103 ( n8067 , n173 , n30419 );
    and g3104 ( n16113 , n31103 , n9904 );
    or g3105 ( n23974 , n32976 , n16797 );
    or g3106 ( n13552 , n24991 , n4175 );
    and g3107 ( n28656 , n5778 , n26574 );
    xnor g3108 ( n3360 , n9065 , n21754 );
    or g3109 ( n23168 , n19551 , n34482 );
    and g3110 ( n8642 , n9603 , n30788 );
    xnor g3111 ( n20955 , n25234 , n9789 );
    or g3112 ( n17108 , n28521 , n35119 );
    xnor g3113 ( n24684 , n32559 , n31289 );
    and g3114 ( n34999 , n28801 , n27229 );
    xnor g3115 ( n24544 , n6615 , n30223 );
    and g3116 ( n15375 , n33727 , n2107 );
    or g3117 ( n29522 , n6782 , n12837 );
    or g3118 ( n31166 , n15141 , n31514 );
    xnor g3119 ( n22045 , n29955 , n9450 );
    and g3120 ( n33976 , n356 , n618 );
    or g3121 ( n21461 , n35337 , n13305 );
    or g3122 ( n6801 , n18123 , n35402 );
    xnor g3123 ( n17299 , n22127 , n15886 );
    or g3124 ( n5589 , n29891 , n13307 );
    or g3125 ( n11430 , n4951 , n31815 );
    not g3126 ( n17235 , n4448 );
    and g3127 ( n8956 , n31565 , n35362 );
    xnor g3128 ( n12802 , n27263 , n4455 );
    and g3129 ( n7955 , n17799 , n27227 );
    or g3130 ( n33552 , n24157 , n16762 );
    xnor g3131 ( n27227 , n22668 , n32046 );
    and g3132 ( n22348 , n509 , n27841 );
    xnor g3133 ( n11506 , n20685 , n30089 );
    xnor g3134 ( n35767 , n1652 , n24371 );
    xnor g3135 ( n391 , n27239 , n7992 );
    or g3136 ( n2150 , n21353 , n16263 );
    or g3137 ( n34087 , n31355 , n27973 );
    and g3138 ( n14192 , n24877 , n7489 );
    nor g3139 ( n34210 , n31215 , n26879 );
    and g3140 ( n21787 , n18746 , n22644 );
    xnor g3141 ( n25766 , n2221 , n22831 );
    or g3142 ( n28691 , n24510 , n15109 );
    or g3143 ( n7941 , n1337 , n24636 );
    and g3144 ( n32782 , n1917 , n26869 );
    nor g3145 ( n18197 , n4288 , n1174 );
    xnor g3146 ( n21702 , n10461 , n35633 );
    or g3147 ( n10925 , n21840 , n17111 );
    and g3148 ( n5284 , n494 , n21281 );
    or g3149 ( n16360 , n9124 , n27728 );
    or g3150 ( n13124 , n25377 , n11996 );
    or g3151 ( n25704 , n14958 , n22322 );
    and g3152 ( n16331 , n13750 , n33686 );
    and g3153 ( n31749 , n20710 , n18167 );
    nor g3154 ( n30633 , n10834 , n29203 );
    and g3155 ( n568 , n17264 , n31320 );
    xnor g3156 ( n9226 , n17746 , n4960 );
    and g3157 ( n2690 , n16529 , n9368 );
    or g3158 ( n18322 , n30149 , n20797 );
    xnor g3159 ( n5522 , n1785 , n29884 );
    xnor g3160 ( n6372 , n7488 , n9793 );
    or g3161 ( n2290 , n3218 , n24025 );
    xnor g3162 ( n23049 , n15208 , n32310 );
    or g3163 ( n10395 , n31588 , n28668 );
    or g3164 ( n15600 , n31289 , n1256 );
    xnor g3165 ( n35875 , n27841 , n509 );
    or g3166 ( n11554 , n28243 , n12428 );
    not g3167 ( n14265 , n5335 );
    xnor g3168 ( n8148 , n21981 , n9793 );
    not g3169 ( n5120 , n31924 );
    or g3170 ( n56 , n22208 , n18264 );
    or g3171 ( n32941 , n18067 , n24672 );
    or g3172 ( n8518 , n31395 , n8233 );
    and g3173 ( n1103 , n21818 , n35842 );
    xnor g3174 ( n21857 , n22336 , n3222 );
    or g3175 ( n2371 , n4390 , n1414 );
    and g3176 ( n18838 , n10511 , n17348 );
    and g3177 ( n14837 , n20060 , n944 );
    or g3178 ( n25776 , n15020 , n2771 );
    or g3179 ( n16076 , n9793 , n13717 );
    and g3180 ( n30481 , n14642 , n11978 );
    and g3181 ( n6992 , n145 , n1776 );
    xnor g3182 ( n25165 , n30529 , n8863 );
    not g3183 ( n22376 , n32667 );
    and g3184 ( n21457 , n26434 , n33187 );
    or g3185 ( n18560 , n16922 , n20604 );
    not g3186 ( n27261 , n1082 );
    or g3187 ( n7034 , n23483 , n4912 );
    or g3188 ( n26560 , n18234 , n3556 );
    not g3189 ( n30048 , n25602 );
    buf g3190 ( n33157 , n29203 );
    or g3191 ( n6668 , n34328 , n18474 );
    or g3192 ( n1711 , n14371 , n25345 );
    and g3193 ( n3279 , n6201 , n16906 );
    or g3194 ( n32835 , n11467 , n17068 );
    nor g3195 ( n26294 , n15886 , n17345 );
    or g3196 ( n4025 , n18659 , n23323 );
    or g3197 ( n3213 , n24630 , n12566 );
    and g3198 ( n5780 , n6419 , n35670 );
    or g3199 ( n30914 , n16922 , n9357 );
    or g3200 ( n20998 , n28479 , n17974 );
    xnor g3201 ( n18581 , n10777 , n1950 );
    xnor g3202 ( n18050 , n11508 , n6035 );
    and g3203 ( n19933 , n4064 , n33970 );
    not g3204 ( n3856 , n1491 );
    nor g3205 ( n22218 , n31559 , n6586 );
    xnor g3206 ( n6674 , n2700 , n22291 );
    and g3207 ( n406 , n22839 , n17289 );
    nor g3208 ( n3323 , n13679 , n13222 );
    xor g3209 ( n10310 , n33088 , n24276 );
    not g3210 ( n20238 , n15941 );
    or g3211 ( n23174 , n16991 , n10770 );
    or g3212 ( n21017 , n10819 , n22419 );
    and g3213 ( n14962 , n17317 , n6241 );
    and g3214 ( n16133 , n22724 , n9093 );
    and g3215 ( n8891 , n10089 , n17718 );
    not g3216 ( n29676 , n35422 );
    not g3217 ( n28477 , n32095 );
    xnor g3218 ( n31556 , n10410 , n3205 );
    or g3219 ( n35026 , n25857 , n30896 );
    or g3220 ( n13174 , n27291 , n4026 );
    xnor g3221 ( n16342 , n918 , n29884 );
    or g3222 ( n21933 , n34061 , n20812 );
    xnor g3223 ( n18906 , n27722 , n9658 );
    and g3224 ( n4045 , n27463 , n11132 );
    xnor g3225 ( n34143 , n12205 , n28236 );
    and g3226 ( n30483 , n13855 , n4504 );
    xnor g3227 ( n3429 , n5460 , n8432 );
    and g3228 ( n704 , n32562 , n23697 );
    xnor g3229 ( n22178 , n15821 , n24282 );
    or g3230 ( n27499 , n24346 , n6683 );
    and g3231 ( n32266 , n29221 , n1871 );
    or g3232 ( n20075 , n24885 , n29953 );
    and g3233 ( n21372 , n18942 , n11011 );
    and g3234 ( n10942 , n11045 , n10805 );
    and g3235 ( n1122 , n8308 , n21683 );
    not g3236 ( n18536 , n33815 );
    or g3237 ( n14147 , n5287 , n22035 );
    and g3238 ( n32804 , n8839 , n24770 );
    or g3239 ( n32812 , n34531 , n30327 );
    or g3240 ( n13100 , n13681 , n12950 );
    or g3241 ( n5319 , n16684 , n3842 );
    xnor g3242 ( n21267 , n24590 , n22142 );
    or g3243 ( n35037 , n1273 , n13952 );
    and g3244 ( n13615 , n2058 , n13727 );
    xnor g3245 ( n32560 , n23722 , n25713 );
    xnor g3246 ( n19404 , n30634 , n23139 );
    or g3247 ( n5314 , n5593 , n4912 );
    or g3248 ( n29775 , n1830 , n7151 );
    or g3249 ( n24524 , n27226 , n3191 );
    nor g3250 ( n12790 , n35927 , n14855 );
    or g3251 ( n24233 , n9205 , n908 );
    or g3252 ( n35620 , n365 , n2299 );
    not g3253 ( n33840 , n32715 );
    not g3254 ( n34814 , n915 );
    or g3255 ( n6129 , n26926 , n128 );
    xnor g3256 ( n7159 , n11802 , n32857 );
    and g3257 ( n29118 , n17462 , n23345 );
    and g3258 ( n3565 , n197 , n389 );
    xnor g3259 ( n19554 , n4186 , n25174 );
    nor g3260 ( n13904 , n1962 , n17067 );
    or g3261 ( n32882 , n5335 , n32020 );
    or g3262 ( n11655 , n14211 , n8392 );
    or g3263 ( n6065 , n18906 , n26290 );
    not g3264 ( n13113 , n31289 );
    not g3265 ( n14278 , n4878 );
    or g3266 ( n16386 , n19950 , n3805 );
    or g3267 ( n17959 , n32095 , n1739 );
    and g3268 ( n30134 , n3434 , n31393 );
    and g3269 ( n28103 , n30869 , n10810 );
    nor g3270 ( n25604 , n3205 , n7112 );
    or g3271 ( n25370 , n1236 , n25659 );
    or g3272 ( n9753 , n3379 , n9731 );
    nor g3273 ( n24368 , n4962 , n29767 );
    or g3274 ( n7494 , n1334 , n32505 );
    or g3275 ( n24369 , n19984 , n30006 );
    or g3276 ( n16985 , n9726 , n3824 );
    xnor g3277 ( n13501 , n10125 , n4962 );
    or g3278 ( n15943 , n4878 , n26242 );
    xnor g3279 ( n32940 , n7363 , n4962 );
    or g3280 ( n21685 , n23138 , n17191 );
    not g3281 ( n34521 , n1529 );
    or g3282 ( n18480 , n25651 , n26480 );
    or g3283 ( n31217 , n18458 , n745 );
    or g3284 ( n6337 , n29158 , n17872 );
    and g3285 ( n11613 , n33612 , n13200 );
    and g3286 ( n11878 , n29193 , n23506 );
    xnor g3287 ( n9048 , n32227 , n3205 );
    nor g3288 ( n16021 , n25829 , n26054 );
    or g3289 ( n11480 , n28798 , n14918 );
    or g3290 ( n48 , n13714 , n24333 );
    and g3291 ( n13397 , n25965 , n6396 );
    or g3292 ( n18392 , n9045 , n16345 );
    and g3293 ( n21822 , n24650 , n14149 );
    or g3294 ( n25089 , n3384 , n23921 );
    or g3295 ( n9099 , n10072 , n16797 );
    and g3296 ( n28610 , n11754 , n35597 );
    xnor g3297 ( n8951 , n33669 , n19861 );
    xnor g3298 ( n7016 , n31177 , n27069 );
    xnor g3299 ( n15722 , n21528 , n26805 );
    or g3300 ( n7791 , n11401 , n8412 );
    xnor g3301 ( n10157 , n4216 , n36039 );
    nor g3302 ( n25070 , n5067 , n8002 );
    xnor g3303 ( n32492 , n12907 , n29884 );
    and g3304 ( n31006 , n18056 , n8995 );
    and g3305 ( n32133 , n26857 , n35781 );
    and g3306 ( n8632 , n6433 , n22011 );
    xnor g3307 ( n17218 , n2061 , n30742 );
    xnor g3308 ( n31377 , n14793 , n25394 );
    or g3309 ( n27460 , n29942 , n20812 );
    xnor g3310 ( n21717 , n19471 , n28759 );
    xnor g3311 ( n3064 , n16061 , n21343 );
    or g3312 ( n3934 , n5335 , n21297 );
    or g3313 ( n3163 , n32565 , n22467 );
    or g3314 ( n23291 , n23846 , n19058 );
    or g3315 ( n19826 , n18037 , n3352 );
    or g3316 ( n16121 , n5658 , n27172 );
    or g3317 ( n27220 , n9380 , n32425 );
    not g3318 ( n24946 , n27632 );
    or g3319 ( n21620 , n2225 , n16594 );
    not g3320 ( n35877 , n29921 );
    or g3321 ( n26463 , n4032 , n10415 );
    or g3322 ( n34958 , n17127 , n14699 );
    or g3323 ( n19212 , n13563 , n29393 );
    or g3324 ( n1490 , n23116 , n15439 );
    and g3325 ( n30763 , n16866 , n18911 );
    or g3326 ( n27063 , n14464 , n15290 );
    or g3327 ( n11169 , n22943 , n29604 );
    or g3328 ( n26471 , n24783 , n28668 );
    and g3329 ( n12801 , n14012 , n5808 );
    xnor g3330 ( n33183 , n19019 , n15403 );
    not g3331 ( n17709 , n4455 );
    xnor g3332 ( n33920 , n28808 , n4288 );
    or g3333 ( n10877 , n5335 , n10878 );
    and g3334 ( n12837 , n724 , n35939 );
    xnor g3335 ( n1140 , n29159 , n32715 );
    or g3336 ( n7174 , n8205 , n33098 );
    or g3337 ( n16453 , n17466 , n36000 );
    or g3338 ( n8968 , n13303 , n21652 );
    or g3339 ( n13410 , n1790 , n6374 );
    nor g3340 ( n5513 , n1488 , n22061 );
    and g3341 ( n7961 , n9889 , n19177 );
    buf g3342 ( n20601 , n18088 );
    or g3343 ( n25620 , n32857 , n22947 );
    or g3344 ( n22349 , n20219 , n23090 );
    xnor g3345 ( n28587 , n34704 , n35852 );
    not g3346 ( n5213 , n31085 );
    or g3347 ( n34952 , n7295 , n26662 );
    or g3348 ( n17867 , n32584 , n2489 );
    xnor g3349 ( n19528 , n30833 , n6435 );
    or g3350 ( n23700 , n1505 , n26659 );
    or g3351 ( n21835 , n1950 , n16858 );
    or g3352 ( n15995 , n18106 , n23187 );
    xnor g3353 ( n23310 , n31091 , n25281 );
    not g3354 ( n26336 , n22245 );
    or g3355 ( n12583 , n1413 , n4254 );
    xnor g3356 ( n17416 , n12699 , n6668 );
    xnor g3357 ( n25257 , n16937 , n32851 );
    or g3358 ( n3516 , n25510 , n25812 );
    xnor g3359 ( n28794 , n5533 , n4878 );
    and g3360 ( n20273 , n17464 , n27054 );
    not g3361 ( n26890 , n12811 );
    or g3362 ( n22587 , n30241 , n2119 );
    xnor g3363 ( n1811 , n29529 , n35927 );
    or g3364 ( n26118 , n31559 , n33146 );
    or g3365 ( n29239 , n1723 , n27437 );
    or g3366 ( n19239 , n26751 , n9317 );
    or g3367 ( n29685 , n17897 , n24672 );
    and g3368 ( n12553 , n17216 , n15938 );
    not g3369 ( n14611 , n19952 );
    or g3370 ( n19233 , n26667 , n978 );
    or g3371 ( n29966 , n830 , n10411 );
    xnor g3372 ( n20289 , n1795 , n31272 );
    xnor g3373 ( n19461 , n9607 , n20337 );
    xnor g3374 ( n29396 , n5877 , n28711 );
    nor g3375 ( n21484 , n1950 , n34383 );
    not g3376 ( n9210 , n341 );
    not g3377 ( n33936 , n16620 );
    and g3378 ( n18970 , n34736 , n1875 );
    or g3379 ( n27593 , n11489 , n14652 );
    not g3380 ( n6785 , n11046 );
    or g3381 ( n19870 , n33918 , n12996 );
    or g3382 ( n15354 , n7540 , n23245 );
    or g3383 ( n12027 , n31238 , n12128 );
    and g3384 ( n30097 , n7445 , n26835 );
    xnor g3385 ( n16956 , n15081 , n27251 );
    not g3386 ( n31287 , n22291 );
    xnor g3387 ( n1872 , n8614 , n4687 );
    or g3388 ( n4411 , n23670 , n19939 );
    or g3389 ( n34520 , n10894 , n23118 );
    nor g3390 ( n29096 , n29824 , n22279 );
    xnor g3391 ( n24906 , n1525 , n2326 );
    xnor g3392 ( n33259 , n9703 , n721 );
    not g3393 ( n9195 , n4962 );
    or g3394 ( n31286 , n337 , n23032 );
    or g3395 ( n32607 , n7393 , n28324 );
    xnor g3396 ( n29030 , n15740 , n14264 );
    nor g3397 ( n702 , n28563 , n32528 );
    and g3398 ( n4702 , n14247 , n23649 );
    or g3399 ( n16589 , n7591 , n10725 );
    and g3400 ( n14132 , n8690 , n11303 );
    nor g3401 ( n18409 , n4498 , n20621 );
    xnor g3402 ( n25774 , n23864 , n26779 );
    or g3403 ( n3896 , n11534 , n7755 );
    xnor g3404 ( n20363 , n27066 , n1950 );
    or g3405 ( n19520 , n4878 , n22873 );
    not g3406 ( n11826 , n9828 );
    or g3407 ( n10536 , n34463 , n25831 );
    and g3408 ( n15875 , n588 , n6700 );
    and g3409 ( n5465 , n9714 , n11803 );
    or g3410 ( n9746 , n11001 , n27501 );
    xnor g3411 ( n6514 , n31659 , n13777 );
    not g3412 ( n7055 , n10894 );
    xnor g3413 ( n23029 , n2167 , n14931 );
    or g3414 ( n27106 , n11455 , n12135 );
    or g3415 ( n35879 , n28170 , n7123 );
    or g3416 ( n35373 , n15975 , n18686 );
    or g3417 ( n2332 , n25912 , n10432 );
    xnor g3418 ( n8467 , n22166 , n35866 );
    not g3419 ( n4230 , n23614 );
    xnor g3420 ( n24623 , n10783 , n31215 );
    xnor g3421 ( n31703 , n19736 , n15299 );
    or g3422 ( n27486 , n34334 , n22322 );
    and g3423 ( n16311 , n24838 , n12041 );
    and g3424 ( n31736 , n17917 , n13006 );
    or g3425 ( n12828 , n3227 , n8707 );
    xnor g3426 ( n25204 , n15483 , n34392 );
    or g3427 ( n18856 , n29161 , n21164 );
    or g3428 ( n32238 , n15999 , n17612 );
    xnor g3429 ( n14864 , n6182 , n34997 );
    xnor g3430 ( n26210 , n11485 , n18964 );
    xnor g3431 ( n24211 , n8434 , n31799 );
    or g3432 ( n2756 , n5179 , n8312 );
    or g3433 ( n5219 , n30838 , n7417 );
    or g3434 ( n31021 , n16981 , n35402 );
    and g3435 ( n29397 , n34486 , n2306 );
    and g3436 ( n4835 , n6103 , n22387 );
    or g3437 ( n22677 , n22379 , n17888 );
    or g3438 ( n31721 , n34836 , n1583 );
    or g3439 ( n35860 , n19984 , n970 );
    xnor g3440 ( n33422 , n1173 , n35920 );
    or g3441 ( n3326 , n10669 , n23085 );
    or g3442 ( n34502 , n20842 , n35559 );
    xnor g3443 ( n34059 , n34455 , n30421 );
    not g3444 ( n13262 , n31799 );
    and g3445 ( n2791 , n27497 , n29577 );
    or g3446 ( n28626 , n26706 , n2117 );
    not g3447 ( n5742 , n26003 );
    and g3448 ( n27016 , n16150 , n30439 );
    xnor g3449 ( n31306 , n26472 , n7540 );
    and g3450 ( n30297 , n11482 , n2599 );
    xnor g3451 ( n25057 , n29856 , n27199 );
    or g3452 ( n31241 , n31559 , n7229 );
    or g3453 ( n34919 , n4352 , n22138 );
    nor g3454 ( n24285 , n18652 , n33956 );
    or g3455 ( n31790 , n19216 , n34923 );
    or g3456 ( n35632 , n14405 , n7417 );
    and g3457 ( n10623 , n31877 , n12670 );
    or g3458 ( n5767 , n35717 , n26365 );
    and g3459 ( n1204 , n13581 , n35452 );
    or g3460 ( n23366 , n28902 , n29322 );
    and g3461 ( n25465 , n31340 , n29591 );
    or g3462 ( n35850 , n31289 , n120 );
    or g3463 ( n27403 , n27226 , n12554 );
    or g3464 ( n10376 , n7777 , n29048 );
    or g3465 ( n27982 , n26812 , n24696 );
    and g3466 ( n26703 , n23969 , n35320 );
    or g3467 ( n16282 , n29884 , n19368 );
    or g3468 ( n4658 , n4105 , n15439 );
    or g3469 ( n36050 , n10460 , n29953 );
    nor g3470 ( n25560 , n16731 , n3129 );
    xnor g3471 ( n23822 , n24930 , n11587 );
    nor g3472 ( n10893 , n35927 , n26126 );
    nor g3473 ( n24686 , n31799 , n35584 );
    xnor g3474 ( n20823 , n20059 , n32715 );
    and g3475 ( n30883 , n7694 , n22832 );
    or g3476 ( n3823 , n11970 , n3805 );
    or g3477 ( n5787 , n767 , n27053 );
    or g3478 ( n17264 , n13418 , n4095 );
    xnor g3479 ( n17830 , n3995 , n14931 );
    xnor g3480 ( n32232 , n1195 , n19984 );
    xnor g3481 ( n17566 , n25816 , n15612 );
    or g3482 ( n31352 , n1950 , n10563 );
    xnor g3483 ( n3865 , n19605 , n2523 );
    nor g3484 ( n20069 , n16620 , n35995 );
    or g3485 ( n13680 , n20214 , n7726 );
    xnor g3486 ( n15105 , n23185 , n31799 );
    or g3487 ( n18048 , n22777 , n8392 );
    xnor g3488 ( n6393 , n16944 , n18379 );
    or g3489 ( n26913 , n35419 , n3979 );
    or g3490 ( n17653 , n18824 , n17357 );
    or g3491 ( n5666 , n6525 , n26480 );
    xnor g3492 ( n11862 , n28163 , n9793 );
    or g3493 ( n17055 , n6386 , n19732 );
    xnor g3494 ( n21454 , n9862 , n7540 );
    nor g3495 ( n4967 , n16996 , n15689 );
    or g3496 ( n20061 , n14633 , n2460 );
    or g3497 ( n5198 , n34471 , n5338 );
    and g3498 ( n3832 , n31555 , n22459 );
    or g3499 ( n34131 , n8008 , n763 );
    xnor g3500 ( n30554 , n29470 , n6283 );
    nor g3501 ( n2536 , n5081 , n31945 );
    or g3502 ( n28801 , n11490 , n27728 );
    xnor g3503 ( n26909 , n4480 , n36085 );
    or g3504 ( n1861 , n13716 , n15393 );
    or g3505 ( n16640 , n34776 , n1063 );
    or g3506 ( n32550 , n26013 , n10694 );
    and g3507 ( n9647 , n14478 , n7180 );
    or g3508 ( n2466 , n29989 , n28837 );
    or g3509 ( n28474 , n9793 , n29462 );
    xnor g3510 ( n16860 , n26257 , n29879 );
    or g3511 ( n19080 , n4962 , n19951 );
    or g3512 ( n13147 , n34121 , n24518 );
    or g3513 ( n32420 , n9789 , n5127 );
    or g3514 ( n29005 , n5335 , n15874 );
    xnor g3515 ( n30112 , n11248 , n32095 );
    or g3516 ( n30906 , n23342 , n5881 );
    xnor g3517 ( n28067 , n10948 , n30179 );
    not g3518 ( n822 , n17568 );
    and g3519 ( n29796 , n30671 , n31226 );
    not g3520 ( n11407 , n18876 );
    or g3521 ( n22023 , n27226 , n19413 );
    xnor g3522 ( n3394 , n5026 , n28846 );
    and g3523 ( n34250 , n32223 , n249 );
    and g3524 ( n6021 , n25410 , n25910 );
    or g3525 ( n8232 , n10612 , n27502 );
    or g3526 ( n6494 , n32095 , n14987 );
    or g3527 ( n16277 , n17744 , n5252 );
    and g3528 ( n27525 , n26954 , n17555 );
    or g3529 ( n7203 , n27226 , n12586 );
    or g3530 ( n8896 , n16288 , n12953 );
    not g3531 ( n28806 , n2685 );
    or g3532 ( n5810 , n3205 , n29006 );
    nor g3533 ( n23150 , n16857 , n30137 );
    xnor g3534 ( n14917 , n22837 , n27426 );
    or g3535 ( n7781 , n24310 , n3165 );
    not g3536 ( n16257 , n30840 );
    xnor g3537 ( n19693 , n32485 , n12357 );
    or g3538 ( n24255 , n18136 , n26002 );
    xnor g3539 ( n31407 , n26211 , n8805 );
    or g3540 ( n21400 , n33127 , n30732 );
    or g3541 ( n15366 , n9658 , n14327 );
    and g3542 ( n35732 , n23313 , n11545 );
    or g3543 ( n3253 , n24043 , n2502 );
    or g3544 ( n35463 , n14121 , n30287 );
    or g3545 ( n17533 , n13740 , n6340 );
    and g3546 ( n687 , n28280 , n31360 );
    not g3547 ( n13935 , n22471 );
    or g3548 ( n34368 , n18424 , n34248 );
    xnor g3549 ( n30805 , n20626 , n31289 );
    or g3550 ( n34309 , n9005 , n30380 );
    nor g3551 ( n32931 , n10894 , n785 );
    or g3552 ( n2355 , n1455 , n30654 );
    or g3553 ( n32245 , n19456 , n19173 );
    or g3554 ( n18319 , n28659 , n4318 );
    or g3555 ( n35044 , n22300 , n31055 );
    nor g3556 ( n27367 , n9658 , n18837 );
    or g3557 ( n17154 , n175 , n23402 );
    or g3558 ( n16157 , n4288 , n31284 );
    or g3559 ( n11183 , n5335 , n21321 );
    or g3560 ( n17366 , n26208 , n29592 );
    or g3561 ( n7179 , n237 , n16077 );
    or g3562 ( n16921 , n27766 , n3958 );
    or g3563 ( n35698 , n23208 , n16326 );
    and g3564 ( n13863 , n12770 , n12271 );
    nor g3565 ( n31442 , n25602 , n29433 );
    nor g3566 ( n784 , n15745 , n20457 );
    or g3567 ( n670 , n10217 , n32923 );
    and g3568 ( n5186 , n1002 , n12505 );
    xnor g3569 ( n14773 , n4813 , n18200 );
    or g3570 ( n32169 , n4962 , n9016 );
    and g3571 ( n2429 , n29747 , n7753 );
    and g3572 ( n11248 , n31706 , n11138 );
    nor g3573 ( n5419 , n30742 , n24930 );
    nor g3574 ( n35484 , n30742 , n12257 );
    and g3575 ( n31651 , n17569 , n17107 );
    and g3576 ( n35770 , n17109 , n34310 );
    or g3577 ( n27531 , n6558 , n7763 );
    or g3578 ( n18666 , n19897 , n3842 );
    xnor g3579 ( n4162 , n17896 , n21675 );
    or g3580 ( n21007 , n32711 , n12165 );
    and g3581 ( n14778 , n29314 , n34601 );
    not g3582 ( n26019 , n6775 );
    not g3583 ( n1091 , n23667 );
    and g3584 ( n26675 , n21807 , n33 );
    or g3585 ( n1789 , n21069 , n6965 );
    and g3586 ( n330 , n15533 , n26252 );
    and g3587 ( n20780 , n17453 , n10136 );
    and g3588 ( n6606 , n7338 , n26841 );
    not g3589 ( n26406 , n28814 );
    xnor g3590 ( n7967 , n34082 , n32740 );
    or g3591 ( n33051 , n27021 , n32329 );
    not g3592 ( n24329 , n3205 );
    or g3593 ( n26059 , n18837 , n29592 );
    or g3594 ( n13151 , n2027 , n35792 );
    and g3595 ( n12864 , n2755 , n4461 );
    and g3596 ( n33251 , n7782 , n21740 );
    and g3597 ( n11071 , n13847 , n25635 );
    or g3598 ( n33667 , n20439 , n6441 );
    or g3599 ( n5365 , n13300 , n30292 );
    or g3600 ( n35469 , n30742 , n16169 );
    or g3601 ( n17762 , n18681 , n584 );
    and g3602 ( n8362 , n21710 , n9098 );
    or g3603 ( n23199 , n24371 , n33648 );
    and g3604 ( n1867 , n23074 , n31639 );
    not g3605 ( n3599 , n7759 );
    or g3606 ( n4626 , n12790 , n4328 );
    xnor g3607 ( n5640 , n24380 , n11605 );
    or g3608 ( n16774 , n2570 , n33737 );
    or g3609 ( n28128 , n31272 , n23759 );
    or g3610 ( n35730 , n28489 , n23626 );
    not g3611 ( n18642 , n31559 );
    and g3612 ( n35017 , n4137 , n5444 );
    not g3613 ( n15158 , n7697 );
    or g3614 ( n25769 , n4616 , n24330 );
    or g3615 ( n31007 , n12289 , n34467 );
    and g3616 ( n31387 , n14542 , n8906 );
    xnor g3617 ( n14330 , n28224 , n28190 );
    not g3618 ( n26095 , n787 );
    and g3619 ( n12431 , n156 , n28138 );
    or g3620 ( n26433 , n12489 , n10762 );
    xnor g3621 ( n3732 , n16004 , n14399 );
    or g3622 ( n20532 , n5335 , n20963 );
    and g3623 ( n3893 , n20594 , n6792 );
    xnor g3624 ( n9261 , n5402 , n16922 );
    xnor g3625 ( n4041 , n30801 , n11212 );
    and g3626 ( n8959 , n26462 , n21182 );
    or g3627 ( n1539 , n26456 , n5618 );
    and g3628 ( n3307 , n25630 , n17274 );
    or g3629 ( n23011 , n4853 , n16005 );
    or g3630 ( n29423 , n6311 , n15145 );
    or g3631 ( n13403 , n25129 , n28668 );
    nor g3632 ( n31855 , n32095 , n24853 );
    or g3633 ( n11102 , n16937 , n24710 );
    or g3634 ( n35254 , n31289 , n34491 );
    xor g3635 ( n28572 , n2317 , n32226 );
    or g3636 ( n870 , n23019 , n32793 );
    and g3637 ( n15210 , n21872 , n10575 );
    or g3638 ( n13827 , n32953 , n18143 );
    or g3639 ( n8694 , n32715 , n20305 );
    and g3640 ( n14719 , n25824 , n16810 );
    nor g3641 ( n25763 , n30479 , n19843 );
    or g3642 ( n3695 , n23661 , n1824 );
    and g3643 ( n31552 , n2598 , n27335 );
    xnor g3644 ( n15380 , n805 , n34937 );
    or g3645 ( n19610 , n32660 , n15145 );
    or g3646 ( n8925 , n23322 , n11312 );
    and g3647 ( n3041 , n19564 , n29012 );
    and g3648 ( n31332 , n32474 , n8383 );
    or g3649 ( n24263 , n15179 , n4907 );
    or g3650 ( n19176 , n695 , n4130 );
    not g3651 ( n18991 , n35173 );
    or g3652 ( n27859 , n20203 , n34375 );
    or g3653 ( n18620 , n6025 , n4847 );
    or g3654 ( n21899 , n9396 , n18173 );
    or g3655 ( n23232 , n14253 , n4363 );
    not g3656 ( n16348 , n20558 );
    and g3657 ( n24833 , n3275 , n9664 );
    and g3658 ( n3485 , n32399 , n21136 );
    and g3659 ( n4604 , n28663 , n31076 );
    and g3660 ( n29767 , n19805 , n28530 );
    or g3661 ( n28464 , n4288 , n32160 );
    and g3662 ( n20272 , n27048 , n21530 );
    or g3663 ( n36054 , n25609 , n20773 );
    and g3664 ( n23322 , n5680 , n11962 );
    and g3665 ( n13149 , n23528 , n22764 );
    or g3666 ( n13825 , n5287 , n7442 );
    nor g3667 ( n30427 , n31864 , n28062 );
    or g3668 ( n18657 , n3222 , n28342 );
    or g3669 ( n32310 , n18092 , n11211 );
    or g3670 ( n3862 , n32715 , n17677 );
    xnor g3671 ( n18861 , n4405 , n25602 );
    not g3672 ( n10424 , n3222 );
    or g3673 ( n14122 , n12236 , n3239 );
    or g3674 ( n11809 , n23420 , n3437 );
    and g3675 ( n2546 , n14548 , n24784 );
    or g3676 ( n13378 , n23519 , n10380 );
    and g3677 ( n10176 , n7995 , n20077 );
    or g3678 ( n25375 , n24890 , n6857 );
    xnor g3679 ( n25217 , n26158 , n21560 );
    or g3680 ( n12793 , n5062 , n28191 );
    and g3681 ( n26100 , n33313 , n10384 );
    and g3682 ( n21248 , n10592 , n22995 );
    xnor g3683 ( n24857 , n24468 , n11455 );
    nor g3684 ( n28250 , n5335 , n21371 );
    or g3685 ( n9987 , n34109 , n35913 );
    or g3686 ( n2789 , n5303 , n34639 );
    or g3687 ( n27780 , n4960 , n16691 );
    nor g3688 ( n20004 , n6524 , n20573 );
    or g3689 ( n22786 , n2641 , n15653 );
    or g3690 ( n32721 , n6767 , n33906 );
    or g3691 ( n12004 , n31289 , n14158 );
    and g3692 ( n286 , n17200 , n24079 );
    or g3693 ( n26734 , n18820 , n17872 );
    or g3694 ( n7244 , n25115 , n2712 );
    or g3695 ( n8765 , n28935 , n28456 );
    or g3696 ( n23881 , n36034 , n19814 );
    xnor g3697 ( n28243 , n34908 , n16496 );
    xnor g3698 ( n7319 , n9900 , n17364 );
    and g3699 ( n6052 , n35165 , n33150 );
    and g3700 ( n29373 , n20779 , n24911 );
    xnor g3701 ( n18719 , n11621 , n4878 );
    xnor g3702 ( n20192 , n15985 , n15255 );
    and g3703 ( n18633 , n3853 , n25961 );
    and g3704 ( n15064 , n28466 , n22867 );
    xnor g3705 ( n27123 , n9583 , n24643 );
    xnor g3706 ( n34510 , n28073 , n32289 );
    and g3707 ( n16216 , n17519 , n18701 );
    or g3708 ( n20034 , n25817 , n3437 );
    xnor g3709 ( n1699 , n18066 , n36072 );
    or g3710 ( n6327 , n29274 , n14242 );
    or g3711 ( n9651 , n4960 , n11671 );
    xnor g3712 ( n11992 , n35916 , n5287 );
    nor g3713 ( n18772 , n30742 , n11041 );
    or g3714 ( n23592 , n6626 , n7748 );
    not g3715 ( n5821 , n7357 );
    or g3716 ( n2797 , n24211 , n12201 );
    and g3717 ( n3295 , n9749 , n34904 );
    or g3718 ( n22698 , n14740 , n19887 );
    nor g3719 ( n17763 , n1950 , n4030 );
    xnor g3720 ( n926 , n3520 , n4743 );
    xnor g3721 ( n22579 , n11309 , n6415 );
    or g3722 ( n35861 , n33772 , n19105 );
    not g3723 ( n11115 , n33168 );
    nor g3724 ( n4333 , n35950 , n31058 );
    or g3725 ( n25251 , n23292 , n30708 );
    or g3726 ( n31678 , n17482 , n188 );
    nor g3727 ( n15349 , n31559 , n19319 );
    xnor g3728 ( n33787 , n8286 , n24371 );
    xnor g3729 ( n31091 , n16595 , n9789 );
    or g3730 ( n29312 , n34244 , n9867 );
    or g3731 ( n20307 , n23255 , n14298 );
    xnor g3732 ( n33037 , n33697 , n4962 );
    xnor g3733 ( n19587 , n6125 , n30577 );
    and g3734 ( n12886 , n19911 , n14896 );
    or g3735 ( n19289 , n19827 , n1511 );
    nor g3736 ( n32006 , n35112 , n33933 );
    and g3737 ( n32958 , n31428 , n275 );
    xnor g3738 ( n27939 , n7155 , n31632 );
    xnor g3739 ( n831 , n17193 , n12564 );
    or g3740 ( n1242 , n32584 , n26258 );
    not g3741 ( n24260 , n18649 );
    not g3742 ( n29430 , n7028 );
    xnor g3743 ( n27839 , n32017 , n19194 );
    or g3744 ( n23293 , n30742 , n6206 );
    xnor g3745 ( n35856 , n26039 , n17140 );
    or g3746 ( n12070 , n24419 , n13480 );
    or g3747 ( n17667 , n22260 , n20840 );
    xnor g3748 ( n28863 , n12502 , n24371 );
    xnor g3749 ( n21762 , n28819 , n30608 );
    xnor g3750 ( n19510 , n5883 , n14979 );
    not g3751 ( n17621 , n27291 );
    or g3752 ( n7260 , n35927 , n23760 );
    xnor g3753 ( n12360 , n3005 , n4962 );
    and g3754 ( n21271 , n19063 , n11397 );
    and g3755 ( n24864 , n28936 , n35594 );
    or g3756 ( n14853 , n8277 , n31773 );
    not g3757 ( n24711 , n4758 );
    xnor g3758 ( n26579 , n7302 , n25602 );
    or g3759 ( n12233 , n10287 , n21644 );
    xnor g3760 ( n25045 , n21738 , n25127 );
    and g3761 ( n17726 , n11642 , n12008 );
    or g3762 ( n28919 , n23020 , n14706 );
    xnor g3763 ( n29836 , n24251 , n21625 );
    or g3764 ( n619 , n32419 , n2117 );
    or g3765 ( n6244 , n5763 , n32505 );
    or g3766 ( n14838 , n9663 , n8353 );
    or g3767 ( n29463 , n25054 , n17612 );
    or g3768 ( n5957 , n33053 , n10140 );
    xnor g3769 ( n26669 , n14848 , n25867 );
    and g3770 ( n9193 , n24988 , n2372 );
    or g3771 ( n26361 , n28609 , n19939 );
    or g3772 ( n35270 , n19057 , n11850 );
    or g3773 ( n16681 , n22437 , n1715 );
    or g3774 ( n14527 , n26049 , n9915 );
    or g3775 ( n33359 , n28178 , n16919 );
    or g3776 ( n5572 , n30742 , n17806 );
    not g3777 ( n26329 , n35938 );
    not g3778 ( n11238 , n21320 );
    nor g3779 ( n23750 , n22929 , n8832 );
    nor g3780 ( n35749 , n1027 , n5088 );
    or g3781 ( n8603 , n10894 , n29103 );
    not g3782 ( n8524 , n25602 );
    or g3783 ( n17832 , n24458 , n19421 );
    or g3784 ( n33696 , n5024 , n3514 );
    xnor g3785 ( n5472 , n26362 , n25340 );
    and g3786 ( n31149 , n14013 , n493 );
    or g3787 ( n13098 , n15825 , n5537 );
    xnor g3788 ( n19926 , n11058 , n32857 );
    or g3789 ( n31839 , n5901 , n21976 );
    xnor g3790 ( n13771 , n7188 , n20603 );
    or g3791 ( n1030 , n23612 , n18542 );
    or g3792 ( n3366 , n3222 , n15272 );
    or g3793 ( n12463 , n10702 , n7726 );
    or g3794 ( n11069 , n26267 , n19336 );
    and g3795 ( n17788 , n765 , n13733 );
    xnor g3796 ( n17836 , n5770 , n31227 );
    xnor g3797 ( n9019 , n11446 , n8398 );
    and g3798 ( n27551 , n12903 , n25259 );
    and g3799 ( n17298 , n191 , n23062 );
    or g3800 ( n25188 , n18583 , n12465 );
    xnor g3801 ( n25561 , n19998 , n5738 );
    or g3802 ( n1569 , n4834 , n28643 );
    or g3803 ( n25787 , n30742 , n22050 );
    or g3804 ( n3866 , n5910 , n578 );
    nor g3805 ( n30195 , n26861 , n32801 );
    or g3806 ( n22143 , n5964 , n35043 );
    or g3807 ( n9646 , n24024 , n13015 );
    and g3808 ( n15345 , n27958 , n26723 );
    or g3809 ( n7675 , n2943 , n22858 );
    xnor g3810 ( n561 , n10418 , n8432 );
    or g3811 ( n1335 , n3222 , n29248 );
    or g3812 ( n31159 , n32863 , n30234 );
    or g3813 ( n9587 , n1918 , n22464 );
    nor g3814 ( n12526 , n31559 , n32590 );
    or g3815 ( n13503 , n25389 , n9663 );
    or g3816 ( n34071 , n26669 , n30519 );
    xnor g3817 ( n19740 , n6982 , n24185 );
    or g3818 ( n9823 , n26053 , n17153 );
    or g3819 ( n35628 , n25342 , n30708 );
    nor g3820 ( n8463 , n19632 , n8919 );
    or g3821 ( n18712 , n11513 , n842 );
    or g3822 ( n17201 , n11544 , n28668 );
    and g3823 ( n3469 , n35438 , n15790 );
    xnor g3824 ( n33929 , n26386 , n35927 );
    or g3825 ( n3061 , n13411 , n5222 );
    xnor g3826 ( n14597 , n22955 , n29884 );
    not g3827 ( n3294 , n25130 );
    or g3828 ( n6236 , n30050 , n5671 );
    nor g3829 ( n13167 , n27226 , n4491 );
    nor g3830 ( n31691 , n22347 , n18115 );
    or g3831 ( n2652 , n17600 , n10973 );
    buf g3832 ( n31627 , n17372 );
    and g3833 ( n11709 , n23780 , n35503 );
    not g3834 ( n24338 , n5952 );
    nor g3835 ( n26894 , n28907 , n6715 );
    or g3836 ( n26905 , n1845 , n32697 );
    not g3837 ( n16259 , n11996 );
    or g3838 ( n14185 , n22163 , n20440 );
    xnor g3839 ( n26235 , n29520 , n28740 );
    or g3840 ( n17005 , n12285 , n14171 );
    and g3841 ( n31812 , n8868 , n25049 );
    or g3842 ( n15302 , n10688 , n30431 );
    xnor g3843 ( n18034 , n7458 , n17931 );
    xnor g3844 ( n29324 , n25828 , n28887 );
    and g3845 ( n15663 , n17822 , n1975 );
    xnor g3846 ( n22552 , n28624 , n1864 );
    or g3847 ( n8116 , n28306 , n4450 );
    or g3848 ( n13590 , n12167 , n33482 );
    and g3849 ( n34350 , n11054 , n2853 );
    xnor g3850 ( n9326 , n1643 , n1950 );
    or g3851 ( n8769 , n14990 , n18477 );
    and g3852 ( n14161 , n11279 , n35183 );
    xnor g3853 ( n25932 , n27269 , n14564 );
    or g3854 ( n4376 , n5280 , n25952 );
    not g3855 ( n3958 , n2092 );
    nor g3856 ( n10248 , n16620 , n2358 );
    or g3857 ( n34137 , n6647 , n26023 );
    or g3858 ( n29846 , n5554 , n14064 );
    xnor g3859 ( n4805 , n17958 , n10885 );
    xnor g3860 ( n26201 , n19133 , n21944 );
    xnor g3861 ( n35897 , n24216 , n29514 );
    and g3862 ( n20960 , n23230 , n3505 );
    and g3863 ( n859 , n35975 , n531 );
    nor g3864 ( n18606 , n4960 , n1447 );
    or g3865 ( n29261 , n15088 , n30280 );
    and g3866 ( n12442 , n27818 , n12211 );
    or g3867 ( n13288 , n35927 , n12830 );
    nor g3868 ( n16337 , n4288 , n14654 );
    or g3869 ( n22563 , n8816 , n4482 );
    and g3870 ( n22014 , n12963 , n6249 );
    xnor g3871 ( n31402 , n9853 , n31289 );
    and g3872 ( n28952 , n29642 , n34187 );
    or g3873 ( n25737 , n8215 , n32329 );
    or g3874 ( n1620 , n15982 , n1942 );
    xnor g3875 ( n32648 , n20095 , n19158 );
    or g3876 ( n18384 , n20336 , n25306 );
    or g3877 ( n16978 , n5765 , n17337 );
    or g3878 ( n3040 , n10894 , n12015 );
    not g3879 ( n4687 , n29713 );
    and g3880 ( n26555 , n31376 , n20606 );
    nor g3881 ( n6365 , n2190 , n20879 );
    or g3882 ( n1325 , n35927 , n3696 );
    or g3883 ( n10196 , n3594 , n16326 );
    xnor g3884 ( n31748 , n17565 , n35151 );
    or g3885 ( n33816 , n2690 , n8295 );
    or g3886 ( n9087 , n28954 , n33098 );
    or g3887 ( n14431 , n15841 , n15290 );
    or g3888 ( n32540 , n36068 , n27812 );
    and g3889 ( n21034 , n6118 , n33777 );
    and g3890 ( n20590 , n21566 , n36060 );
    or g3891 ( n22326 , n22274 , n4426 );
    or g3892 ( n26202 , n34207 , n7726 );
    or g3893 ( n33336 , n29433 , n24710 );
    and g3894 ( n27268 , n24888 , n20706 );
    and g3895 ( n15952 , n17252 , n9972 );
    and g3896 ( n24302 , n1964 , n12940 );
    xnor g3897 ( n3547 , n11201 , n35901 );
    or g3898 ( n19062 , n16527 , n20352 );
    or g3899 ( n30642 , n32584 , n1119 );
    not g3900 ( n28100 , n33450 );
    xnor g3901 ( n25177 , n15979 , n11428 );
    or g3902 ( n19633 , n422 , n33461 );
    or g3903 ( n14895 , n33643 , n8022 );
    nor g3904 ( n33562 , n7253 , n3516 );
    xnor g3905 ( n19809 , n34743 , n31633 );
    nor g3906 ( n6961 , n34855 , n10490 );
    not g3907 ( n22809 , n31951 );
    xnor g3908 ( n25687 , n10207 , n31289 );
    and g3909 ( n6504 , n3413 , n18766 );
    or g3910 ( n23595 , n3178 , n25355 );
    xnor g3911 ( n34878 , n26731 , n9989 );
    xnor g3912 ( n17835 , n26928 , n15086 );
    not g3913 ( n9538 , n19277 );
    or g3914 ( n3526 , n23208 , n23028 );
    or g3915 ( n22203 , n19590 , n22206 );
    and g3916 ( n10678 , n8441 , n19778 );
    and g3917 ( n19800 , n28071 , n33240 );
    xnor g3918 ( n33304 , n16384 , n8750 );
    xnor g3919 ( n30123 , n20329 , n19263 );
    or g3920 ( n34010 , n25346 , n11703 );
    and g3921 ( n23368 , n14933 , n10940 );
    nor g3922 ( n2182 , n32857 , n32080 );
    and g3923 ( n9605 , n28238 , n25356 );
    xnor g3924 ( n32127 , n14910 , n3205 );
    or g3925 ( n32208 , n25894 , n27580 );
    nor g3926 ( n30812 , n13613 , n8000 );
    or g3927 ( n24639 , n9367 , n11703 );
    xnor g3928 ( n34941 , n15844 , n9920 );
    xnor g3929 ( n12493 , n17299 , n19666 );
    and g3930 ( n29942 , n2669 , n8732 );
    and g3931 ( n623 , n28059 , n19292 );
    not g3932 ( n22026 , n34807 );
    and g3933 ( n21456 , n3797 , n936 );
    or g3934 ( n1271 , n30129 , n28324 );
    buf g3935 ( n30826 , n9003 );
    or g3936 ( n88 , n25383 , n18364 );
    xnor g3937 ( n18563 , n345 , n17816 );
    xnor g3938 ( n35446 , n31996 , n26896 );
    nor g3939 ( n976 , n1950 , n29298 );
    or g3940 ( n9705 , n5452 , n33017 );
    or g3941 ( n6926 , n33213 , n2211 );
    nor g3942 ( n20719 , n17568 , n26926 );
    or g3943 ( n30935 , n102 , n16919 );
    xnor g3944 ( n28518 , n26029 , n31768 );
    or g3945 ( n16725 , n5738 , n28780 );
    and g3946 ( n21714 , n27101 , n17489 );
    not g3947 ( n19722 , n27437 );
    nor g3948 ( n16254 , n3946 , n23352 );
    or g3949 ( n26016 , n16212 , n1642 );
    nor g3950 ( n3539 , n4878 , n19287 );
    nor g3951 ( n27015 , n15886 , n34691 );
    or g3952 ( n34682 , n23178 , n23538 );
    or g3953 ( n13772 , n15537 , n2712 );
    or g3954 ( n10100 , n5335 , n12218 );
    and g3955 ( n35265 , n32010 , n15404 );
    and g3956 ( n14327 , n18322 , n19193 );
    or g3957 ( n34678 , n16646 , n12622 );
    xnor g3958 ( n14802 , n31099 , n10894 );
    or g3959 ( n25364 , n8432 , n21700 );
    and g3960 ( n17681 , n3727 , n450 );
    and g3961 ( n30688 , n35050 , n12696 );
    xnor g3962 ( n16842 , n22173 , n729 );
    xnor g3963 ( n12645 , n10433 , n4960 );
    and g3964 ( n22717 , n22325 , n30197 );
    and g3965 ( n24716 , n13945 , n17387 );
    or g3966 ( n16313 , n23781 , n21042 );
    or g3967 ( n4458 , n9793 , n6643 );
    and g3968 ( n31038 , n18545 , n12496 );
    xnor g3969 ( n413 , n29150 , n11357 );
    xnor g3970 ( n34082 , n22791 , n30742 );
    or g3971 ( n5291 , n32532 , n27652 );
    or g3972 ( n9751 , n6757 , n28837 );
    not g3973 ( n16077 , n17316 );
    and g3974 ( n35004 , n3582 , n23340 );
    xnor g3975 ( n1131 , n6230 , n8112 );
    xnor g3976 ( n33705 , n18195 , n7540 );
    and g3977 ( n2438 , n9148 , n15588 );
    xnor g3978 ( n18429 , n31294 , n3261 );
    or g3979 ( n3373 , n30516 , n15805 );
    xnor g3980 ( n13903 , n4276 , n4744 );
    or g3981 ( n17706 , n24371 , n6959 );
    or g3982 ( n5004 , n791 , n3738 );
    and g3983 ( n9768 , n8571 , n14909 );
    or g3984 ( n20298 , n24817 , n8364 );
    and g3985 ( n27811 , n18793 , n29724 );
    xnor g3986 ( n11639 , n32531 , n830 );
    or g3987 ( n9274 , n12645 , n26018 );
    or g3988 ( n16807 , n6528 , n30646 );
    not g3989 ( n10042 , n5382 );
    xnor g3990 ( n3127 , n32139 , n2044 );
    or g3991 ( n7356 , n25275 , n1763 );
    or g3992 ( n31088 , n20092 , n4507 );
    or g3993 ( n6784 , n3136 , n7293 );
    and g3994 ( n30156 , n22875 , n19588 );
    xnor g3995 ( n32241 , n10075 , n11046 );
    and g3996 ( n24953 , n31585 , n3248 );
    or g3997 ( n8251 , n14085 , n19490 );
    or g3998 ( n24828 , n26912 , n10289 );
    or g3999 ( n29755 , n11611 , n23921 );
    not g4000 ( n3004 , n35927 );
    or g4001 ( n23397 , n5995 , n1557 );
    or g4002 ( n35956 , n770 , n10417 );
    or g4003 ( n7551 , n27465 , n24710 );
    and g4004 ( n33764 , n19739 , n34291 );
    or g4005 ( n26793 , n9789 , n8632 );
    or g4006 ( n15723 , n9102 , n25268 );
    not g4007 ( n13963 , n14202 );
    or g4008 ( n35428 , n4962 , n31307 );
    and g4009 ( n549 , n29889 , n10538 );
    or g4010 ( n26402 , n8559 , n17155 );
    or g4011 ( n9645 , n29399 , n26504 );
    and g4012 ( n23471 , n4836 , n21425 );
    xnor g4013 ( n321 , n11955 , n31272 );
    or g4014 ( n35032 , n6812 , n28064 );
    xnor g4015 ( n23063 , n14039 , n31272 );
    nor g4016 ( n9217 , n7885 , n13935 );
    xnor g4017 ( n11935 , n12819 , n9629 );
    and g4018 ( n32446 , n13554 , n21137 );
    nor g4019 ( n12972 , n830 , n26521 );
    or g4020 ( n4298 , n1338 , n32697 );
    not g4021 ( n28586 , n25761 );
    xnor g4022 ( n24814 , n20196 , n27449 );
    or g4023 ( n5799 , n9789 , n1122 );
    xnor g4024 ( n5958 , n24947 , n6417 );
    not g4025 ( n573 , n11046 );
    or g4026 ( n14 , n19532 , n22858 );
    or g4027 ( n21960 , n29713 , n30838 );
    or g4028 ( n17435 , n19197 , n29540 );
    and g4029 ( n8802 , n24 , n33153 );
    or g4030 ( n30430 , n35556 , n28064 );
    or g4031 ( n3580 , n31289 , n20176 );
    and g4032 ( n25896 , n10399 , n10165 );
    not g4033 ( n6441 , n11389 );
    or g4034 ( n3999 , n14832 , n21370 );
    not g4035 ( n23545 , n35481 );
    and g4036 ( n31811 , n5014 , n15035 );
    or g4037 ( n24914 , n21384 , n22783 );
    xnor g4038 ( n28990 , n25454 , n31811 );
    or g4039 ( n3665 , n20071 , n20310 );
    or g4040 ( n28976 , n32906 , n11295 );
    and g4041 ( n9947 , n13317 , n28896 );
    or g4042 ( n6601 , n12532 , n23748 );
    xnor g4043 ( n27823 , n22155 , n32043 );
    xnor g4044 ( n28414 , n14194 , n18189 );
    xnor g4045 ( n21492 , n34434 , n5547 );
    and g4046 ( n26609 , n5328 , n19747 );
    xnor g4047 ( n30396 , n27120 , n23325 );
    xnor g4048 ( n29238 , n14023 , n5620 );
    and g4049 ( n18258 , n10080 , n31281 );
    or g4050 ( n12186 , n16310 , n14699 );
    and g4051 ( n27715 , n21348 , n33818 );
    xnor g4052 ( n1027 , n21781 , n9708 );
    or g4053 ( n24395 , n11530 , n29650 );
    or g4054 ( n15140 , n6376 , n24672 );
    and g4055 ( n11326 , n25944 , n9335 );
    not g4056 ( n6406 , n30714 );
    xnor g4057 ( n15414 , n23350 , n16620 );
    or g4058 ( n7189 , n1757 , n20601 );
    xnor g4059 ( n31398 , n25043 , n20354 );
    xnor g4060 ( n31676 , n14584 , n6279 );
    and g4061 ( n14737 , n20313 , n24576 );
    or g4062 ( n27972 , n19783 , n21673 );
    xnor g4063 ( n14459 , n12556 , n34552 );
    xnor g4064 ( n1503 , n23459 , n19551 );
    xnor g4065 ( n23987 , n5506 , n30178 );
    and g4066 ( n3129 , n20103 , n22404 );
    xnor g4067 ( n24228 , n29600 , n20650 );
    and g4068 ( n639 , n25406 , n34831 );
    or g4069 ( n20472 , n33058 , n1856 );
    or g4070 ( n34966 , n17747 , n3215 );
    or g4071 ( n28602 , n3205 , n28114 );
    and g4072 ( n26921 , n9152 , n14061 );
    and g4073 ( n30434 , n12688 , n20809 );
    xnor g4074 ( n31958 , n8277 , n4962 );
    buf g4075 ( n6950 , n22783 );
    or g4076 ( n2180 , n12617 , n8153 );
    not g4077 ( n18283 , n35927 );
    or g4078 ( n29039 , n24085 , n11204 );
    xnor g4079 ( n24111 , n1 , n32256 );
    not g4080 ( n22851 , n16716 );
    and g4081 ( n3416 , n9563 , n5399 );
    not g4082 ( n10973 , n33711 );
    or g4083 ( n3798 , n14751 , n34542 );
    nor g4084 ( n22397 , n32584 , n34999 );
    or g4085 ( n7592 , n24539 , n17354 );
    not g4086 ( n2105 , n22471 );
    not g4087 ( n23991 , n5892 );
    not g4088 ( n15736 , n36041 );
    or g4089 ( n16844 , n4140 , n23462 );
    or g4090 ( n35357 , n17802 , n22501 );
    or g4091 ( n35512 , n17273 , n34794 );
    or g4092 ( n16960 , n3222 , n14655 );
    or g4093 ( n22472 , n32938 , n25735 );
    not g4094 ( n9106 , n23978 );
    or g4095 ( n30518 , n31960 , n17974 );
    nor g4096 ( n2534 , n830 , n16087 );
    or g4097 ( n28525 , n9800 , n24356 );
    not g4098 ( n23543 , n26724 );
    not g4099 ( n34493 , n33435 );
    or g4100 ( n27023 , n29081 , n10336 );
    and g4101 ( n3128 , n36001 , n5757 );
    buf g4102 ( n12326 , n3477 );
    xnor g4103 ( n21304 , n23840 , n25174 );
    xnor g4104 ( n23154 , n27271 , n6191 );
    or g4105 ( n11556 , n22182 , n23099 );
    or g4106 ( n4424 , n29839 , n6504 );
    or g4107 ( n34418 , n26406 , n23452 );
    xnor g4108 ( n16657 , n11041 , n889 );
    and g4109 ( n20873 , n8127 , n26518 );
    and g4110 ( n23612 , n12937 , n14011 );
    xnor g4111 ( n12017 , n26165 , n524 );
    xnor g4112 ( n7566 , n13913 , n33821 );
    and g4113 ( n7916 , n11950 , n6350 );
    buf g4114 ( n17337 , n29718 );
    or g4115 ( n15200 , n7651 , n34537 );
    xnor g4116 ( n19557 , n32863 , n30234 );
    nor g4117 ( n34835 , n1274 , n10007 );
    or g4118 ( n13137 , n23912 , n5779 );
    not g4119 ( n20813 , n20850 );
    xnor g4120 ( n16167 , n24822 , n30742 );
    and g4121 ( n16445 , n7179 , n16425 );
    xnor g4122 ( n10742 , n13615 , n26647 );
    or g4123 ( n24913 , n34283 , n2955 );
    not g4124 ( n18845 , n32608 );
    or g4125 ( n16429 , n5287 , n1978 );
    xnor g4126 ( n5098 , n31212 , n8888 );
    or g4127 ( n10666 , n23604 , n17127 );
    and g4128 ( n22996 , n27450 , n2375 );
    or g4129 ( n16440 , n25982 , n25831 );
    and g4130 ( n11578 , n5371 , n20914 );
    and g4131 ( n32944 , n3011 , n6688 );
    and g4132 ( n9817 , n35040 , n16626 );
    and g4133 ( n24102 , n4862 , n1527 );
    or g4134 ( n20054 , n3205 , n26693 );
    or g4135 ( n5947 , n2721 , n15256 );
    or g4136 ( n3589 , n25440 , n34862 );
    nor g4137 ( n24564 , n24879 , n8835 );
    xnor g4138 ( n13894 , n8627 , n24371 );
    xnor g4139 ( n22371 , n29353 , n6132 );
    nor g4140 ( n8919 , n14646 , n15849 );
    or g4141 ( n17473 , n28686 , n3756 );
    or g4142 ( n35709 , n21235 , n30423 );
    or g4143 ( n21416 , n28968 , n12899 );
    or g4144 ( n4925 , n23660 , n12897 );
    and g4145 ( n20642 , n13405 , n5659 );
    nor g4146 ( n6962 , n19551 , n17986 );
    xnor g4147 ( n34681 , n30704 , n25174 );
    buf g4148 ( n949 , n14956 );
    or g4149 ( n15993 , n7095 , n31231 );
    not g4150 ( n18603 , n24371 );
    or g4151 ( n8570 , n22174 , n33447 );
    or g4152 ( n23272 , n34322 , n34600 );
    xnor g4153 ( n11201 , n29692 , n23524 );
    or g4154 ( n14537 , n15614 , n9813 );
    or g4155 ( n11853 , n4833 , n24176 );
    xnor g4156 ( n27493 , n13998 , n16436 );
    or g4157 ( n24039 , n9699 , n19649 );
    xnor g4158 ( n21499 , n11181 , n27390 );
    nor g4159 ( n31264 , n9658 , n30675 );
    or g4160 ( n33819 , n1507 , n17068 );
    or g4161 ( n14216 , n2906 , n5972 );
    and g4162 ( n30659 , n2234 , n23247 );
    or g4163 ( n12888 , n16959 , n9194 );
    or g4164 ( n7552 , n9658 , n30701 );
    or g4165 ( n26372 , n8432 , n983 );
    xnor g4166 ( n7898 , n25928 , n32889 );
    not g4167 ( n21993 , n1874 );
    or g4168 ( n10440 , n21433 , n20806 );
    or g4169 ( n18896 , n8227 , n16649 );
    and g4170 ( n33269 , n27137 , n25875 );
    or g4171 ( n24189 , n10894 , n838 );
    and g4172 ( n35216 , n34733 , n30330 );
    and g4173 ( n1832 , n20429 , n25310 );
    xnor g4174 ( n36013 , n28187 , n8432 );
    nor g4175 ( n24844 , n11309 , n20037 );
    not g4176 ( n31700 , n15886 );
    or g4177 ( n31978 , n32074 , n4363 );
    or g4178 ( n22368 , n3205 , n10410 );
    or g4179 ( n2307 , n24786 , n32808 );
    or g4180 ( n30880 , n10143 , n32808 );
    xnor g4181 ( n1940 , n30417 , n32715 );
    or g4182 ( n23747 , n15886 , n32674 );
    not g4183 ( n13608 , n25602 );
    xnor g4184 ( n19380 , n16945 , n1693 );
    or g4185 ( n26281 , n19551 , n6384 );
    nor g4186 ( n24949 , n1950 , n9075 );
    xnor g4187 ( n25816 , n34208 , n10498 );
    and g4188 ( n7903 , n22438 , n13014 );
    or g4189 ( n6881 , n8432 , n20072 );
    or g4190 ( n18713 , n7802 , n11568 );
    xnor g4191 ( n20602 , n31120 , n26265 );
    xnor g4192 ( n31659 , n3371 , n19551 );
    or g4193 ( n23803 , n15820 , n27053 );
    not g4194 ( n15971 , n24304 );
    or g4195 ( n20874 , n21394 , n32589 );
    nor g4196 ( n13122 , n3205 , n33927 );
    or g4197 ( n26620 , n32820 , n5618 );
    or g4198 ( n31154 , n4962 , n22621 );
    and g4199 ( n34627 , n8721 , n12106 );
    nor g4200 ( n7719 , n30742 , n18381 );
    and g4201 ( n15572 , n18237 , n19426 );
    nor g4202 ( n1865 , n9793 , n26055 );
    or g4203 ( n20591 , n20076 , n31984 );
    and g4204 ( n30665 , n16704 , n33465 );
    not g4205 ( n5824 , n17448 );
    xnor g4206 ( n35853 , n16858 , n1950 );
    nor g4207 ( n22692 , n4288 , n26183 );
    not g4208 ( n13254 , n3205 );
    or g4209 ( n14942 , n23018 , n14973 );
    or g4210 ( n23326 , n16975 , n5779 );
    xnor g4211 ( n22500 , n28781 , n32359 );
    xnor g4212 ( n32543 , n20042 , n8036 );
    and g4213 ( n19710 , n33841 , n10934 );
    not g4214 ( n4361 , n28758 );
    or g4215 ( n9594 , n7597 , n28789 );
    nor g4216 ( n18482 , n10639 , n20340 );
    nor g4217 ( n22730 , n24732 , n24505 );
    or g4218 ( n6410 , n11248 , n21002 );
    or g4219 ( n17997 , n8056 , n27625 );
    or g4220 ( n3173 , n14252 , n9030 );
    xnor g4221 ( n16450 , n11533 , n26927 );
    not g4222 ( n34456 , n22518 );
    or g4223 ( n24033 , n1911 , n12913 );
    or g4224 ( n17589 , n31289 , n30975 );
    or g4225 ( n20735 , n36069 , n35630 );
    nor g4226 ( n5570 , n18538 , n16272 );
    and g4227 ( n12340 , n16281 , n12418 );
    xnor g4228 ( n9017 , n11020 , n8749 );
    xnor g4229 ( n11448 , n9517 , n5335 );
    and g4230 ( n1133 , n3398 , n25009 );
    xnor g4231 ( n27078 , n692 , n32095 );
    or g4232 ( n7331 , n9658 , n1172 );
    not g4233 ( n30904 , n22200 );
    and g4234 ( n5041 , n31888 , n23747 );
    or g4235 ( n12068 , n6062 , n4081 );
    xnor g4236 ( n7774 , n10281 , n4878 );
    or g4237 ( n20204 , n17587 , n26465 );
    nor g4238 ( n33591 , n9793 , n12131 );
    or g4239 ( n10361 , n31799 , n13595 );
    xnor g4240 ( n12713 , n33284 , n18379 );
    xnor g4241 ( n11508 , n2841 , n15886 );
    xnor g4242 ( n5235 , n34668 , n29459 );
    and g4243 ( n21608 , n25152 , n3190 );
    nor g4244 ( n9181 , n3205 , n14536 );
    xnor g4245 ( n5564 , n33633 , n11046 );
    or g4246 ( n16785 , n18524 , n13213 );
    and g4247 ( n22798 , n32296 , n31081 );
    or g4248 ( n34088 , n6777 , n18933 );
    and g4249 ( n35205 , n31271 , n19294 );
    xnor g4250 ( n31898 , n9824 , n36070 );
    and g4251 ( n26265 , n15776 , n35439 );
    or g4252 ( n32024 , n29801 , n8831 );
    buf g4253 ( n33098 , n33464 );
    or g4254 ( n8728 , n10459 , n3052 );
    xnor g4255 ( n5420 , n25257 , n35755 );
    and g4256 ( n18201 , n26990 , n24536 );
    or g4257 ( n31311 , n11247 , n5721 );
    not g4258 ( n25899 , n8447 );
    or g4259 ( n12710 , n8396 , n9855 );
    not g4260 ( n16213 , n18121 );
    or g4261 ( n33991 , n9793 , n25115 );
    or g4262 ( n35485 , n4724 , n32408 );
    xnor g4263 ( n20882 , n6360 , n30742 );
    not g4264 ( n14618 , n35650 );
    or g4265 ( n19847 , n28058 , n2798 );
    or g4266 ( n26203 , n9789 , n6332 );
    and g4267 ( n33125 , n12828 , n30404 );
    or g4268 ( n32954 , n20183 , n15319 );
    xnor g4269 ( n19859 , n12822 , n14501 );
    xnor g4270 ( n32051 , n19878 , n34367 );
    xnor g4271 ( n25454 , n21159 , n3222 );
    or g4272 ( n33612 , n4717 , n24829 );
    or g4273 ( n8403 , n3946 , n34041 );
    or g4274 ( n34565 , n25602 , n25249 );
    and g4275 ( n19387 , n13833 , n24443 );
    not g4276 ( n6487 , n15772 );
    nor g4277 ( n19654 , n16922 , n13127 );
    or g4278 ( n11273 , n24595 , n32091 );
    xnor g4279 ( n21875 , n24243 , n23604 );
    xnor g4280 ( n28007 , n658 , n7540 );
    or g4281 ( n9378 , n28312 , n25710 );
    nor g4282 ( n20489 , n29037 , n16411 );
    or g4283 ( n6840 , n7661 , n31104 );
    or g4284 ( n19899 , n27138 , n29071 );
    and g4285 ( n8804 , n4084 , n30970 );
    xnor g4286 ( n32340 , n27587 , n8432 );
    or g4287 ( n20108 , n32101 , n27501 );
    nor g4288 ( n18723 , n18650 , n14748 );
    and g4289 ( n5625 , n465 , n32212 );
    or g4290 ( n10483 , n22014 , n6683 );
    and g4291 ( n2543 , n7264 , n16418 );
    and g4292 ( n19851 , n17160 , n35145 );
    nor g4293 ( n20774 , n29595 , n32329 );
    buf g4294 ( n12332 , n5339 );
    xnor g4295 ( n6610 , n2690 , n26698 );
    or g4296 ( n34462 , n12450 , n6328 );
    xnor g4297 ( n25702 , n35497 , n274 );
    and g4298 ( n18374 , n34332 , n30863 );
    nor g4299 ( n20377 , n13619 , n27963 );
    or g4300 ( n2430 , n14897 , n23879 );
    nor g4301 ( n14839 , n22831 , n7089 );
    not g4302 ( n19767 , n30732 );
    or g4303 ( n14237 , n27955 , n20595 );
    xor g4304 ( n24509 , n15029 , n16845 );
    and g4305 ( n7096 , n17333 , n28491 );
    or g4306 ( n13851 , n17568 , n35712 );
    or g4307 ( n25600 , n3002 , n34634 );
    nor g4308 ( n28685 , n3938 , n1142 );
    or g4309 ( n32586 , n23896 , n10464 );
    or g4310 ( n22907 , n33988 , n8617 );
    or g4311 ( n23389 , n11818 , n32073 );
    and g4312 ( n7208 , n12400 , n23604 );
    xnor g4313 ( n27217 , n32656 , n31539 );
    or g4314 ( n19326 , n13491 , n3634 );
    and g4315 ( n29322 , n16618 , n11073 );
    not g4316 ( n35728 , n2893 );
    and g4317 ( n23579 , n29777 , n12070 );
    or g4318 ( n9470 , n27005 , n7061 );
    xnor g4319 ( n32098 , n32992 , n29241 );
    and g4320 ( n28070 , n9770 , n15180 );
    or g4321 ( n11384 , n5379 , n35111 );
    or g4322 ( n12518 , n33143 , n12465 );
    and g4323 ( n20952 , n16624 , n21474 );
    or g4324 ( n33644 , n27226 , n31229 );
    nor g4325 ( n2851 , n4574 , n35804 );
    xnor g4326 ( n19002 , n3966 , n4962 );
    and g4327 ( n19395 , n5268 , n18853 );
    or g4328 ( n29924 , n6569 , n12254 );
    or g4329 ( n3049 , n19551 , n9543 );
    or g4330 ( n8497 , n6906 , n25831 );
    or g4331 ( n18105 , n3629 , n1642 );
    and g4332 ( n17078 , n27002 , n19060 );
    not g4333 ( n15517 , n3842 );
    buf g4334 ( n10289 , n17068 );
    or g4335 ( n3886 , n16391 , n5618 );
    xnor g4336 ( n4640 , n6652 , n33689 );
    or g4337 ( n8987 , n20912 , n9915 );
    xnor g4338 ( n19136 , n5940 , n26219 );
    or g4339 ( n18506 , n13489 , n3356 );
    nor g4340 ( n1683 , n5287 , n1764 );
    not g4341 ( n10477 , n5793 );
    xnor g4342 ( n13781 , n17783 , n35072 );
    and g4343 ( n30218 , n15487 , n20736 );
    or g4344 ( n31328 , n20065 , n15444 );
    xnor g4345 ( n3522 , n5022 , n15403 );
    xnor g4346 ( n1925 , n1413 , n1438 );
    or g4347 ( n20276 , n15886 , n12315 );
    or g4348 ( n2365 , n22110 , n15369 );
    and g4349 ( n918 , n31547 , n32254 );
    or g4350 ( n29927 , n16669 , n17111 );
    xnor g4351 ( n24908 , n29265 , n21248 );
    and g4352 ( n20082 , n8854 , n13825 );
    or g4353 ( n29181 , n19809 , n14076 );
    not g4354 ( n26979 , n30742 );
    and g4355 ( n2473 , n33217 , n28061 );
    and g4356 ( n29604 , n13699 , n8243 );
    and g4357 ( n13148 , n19980 , n32317 );
    or g4358 ( n10685 , n18927 , n26659 );
    xnor g4359 ( n17338 , n15884 , n5335 );
    and g4360 ( n36030 , n23673 , n20810 );
    or g4361 ( n3528 , n1378 , n25786 );
    or g4362 ( n28925 , n23604 , n28633 );
    and g4363 ( n5613 , n27194 , n17374 );
    or g4364 ( n30850 , n27457 , n5245 );
    or g4365 ( n29182 , n32600 , n9702 );
    or g4366 ( n31350 , n3946 , n2735 );
    not g4367 ( n19373 , n21884 );
    xnor g4368 ( n1690 , n8080 , n36072 );
    nor g4369 ( n17776 , n30229 , n20148 );
    xnor g4370 ( n25512 , n7200 , n3222 );
    or g4371 ( n32384 , n2329 , n30732 );
    and g4372 ( n4186 , n938 , n21241 );
    or g4373 ( n6549 , n34271 , n28734 );
    xnor g4374 ( n18327 , n11648 , n30553 );
    or g4375 ( n17733 , n3972 , n17133 );
    or g4376 ( n3849 , n31098 , n15109 );
    or g4377 ( n34536 , n7161 , n32959 );
    not g4378 ( n33023 , n4805 );
    or g4379 ( n10373 , n10723 , n27623 );
    xnor g4380 ( n33597 , n18327 , n6370 );
    and g4381 ( n2503 , n13723 , n195 );
    or g4382 ( n11168 , n5178 , n8392 );
    or g4383 ( n847 , n636 , n24259 );
    or g4384 ( n17426 , n30025 , n4254 );
    not g4385 ( n32039 , n34865 );
    and g4386 ( n18574 , n7386 , n7226 );
    or g4387 ( n30794 , n11190 , n33076 );
    not g4388 ( n12223 , n18826 );
    and g4389 ( n3822 , n6245 , n12497 );
    and g4390 ( n282 , n10359 , n32623 );
    and g4391 ( n24091 , n24874 , n25700 );
    xnor g4392 ( n33665 , n26596 , n5781 );
    or g4393 ( n35702 , n22446 , n20576 );
    or g4394 ( n20624 , n19500 , n32634 );
    not g4395 ( n10519 , n12266 );
    xnor g4396 ( n16731 , n28888 , n35927 );
    or g4397 ( n21483 , n7472 , n4318 );
    and g4398 ( n2748 , n10431 , n26178 );
    and g4399 ( n22530 , n4432 , n28913 );
    xnor g4400 ( n25250 , n23535 , n9658 );
    and g4401 ( n11770 , n11421 , n25380 );
    or g4402 ( n35758 , n32095 , n23937 );
    xnor g4403 ( n25750 , n27318 , n35891 );
    xnor g4404 ( n19225 , n27436 , n34967 );
    or g4405 ( n15489 , n19551 , n6528 );
    or g4406 ( n27221 , n1276 , n31627 );
    nor g4407 ( n15045 , n17568 , n4475 );
    and g4408 ( n28867 , n7622 , n13593 );
    or g4409 ( n21925 , n21299 , n8153 );
    xnor g4410 ( n34533 , n34175 , n15060 );
    xnor g4411 ( n7130 , n22447 , n34183 );
    not g4412 ( n8885 , n9658 );
    xnor g4413 ( n14477 , n4720 , n20266 );
    or g4414 ( n16560 , n21213 , n5168 );
    and g4415 ( n1689 , n27789 , n21046 );
    and g4416 ( n8771 , n18628 , n18449 );
    xnor g4417 ( n3650 , n569 , n33014 );
    and g4418 ( n30672 , n7976 , n26859 );
    and g4419 ( n34437 , n10605 , n4676 );
    not g4420 ( n17665 , n19225 );
    xnor g4421 ( n27240 , n34473 , n7966 );
    not g4422 ( n2448 , n30418 );
    or g4423 ( n21856 , n24863 , n5456 );
    or g4424 ( n31035 , n5565 , n3437 );
    xnor g4425 ( n34083 , n19948 , n23352 );
    and g4426 ( n10693 , n26682 , n10255 );
    or g4427 ( n19670 , n4878 , n32348 );
    and g4428 ( n17478 , n18916 , n33736 );
    and g4429 ( n22123 , n8497 , n13621 );
    or g4430 ( n22443 , n21104 , n3188 );
    or g4431 ( n6304 , n3249 , n28191 );
    or g4432 ( n30723 , n9132 , n32958 );
    not g4433 ( n27096 , n7588 );
    or g4434 ( n12733 , n19583 , n30993 );
    and g4435 ( n505 , n13323 , n2670 );
    and g4436 ( n7762 , n6552 , n10436 );
    xnor g4437 ( n18356 , n34791 , n33972 );
    nor g4438 ( n31057 , n5335 , n28417 );
    nor g4439 ( n31020 , n19305 , n1666 );
    and g4440 ( n9690 , n26378 , n16576 );
    and g4441 ( n25904 , n24066 , n29426 );
    buf g4442 ( n20318 , n648 );
    xnor g4443 ( n13790 , n18923 , n830 );
    nor g4444 ( n4817 , n19761 , n24505 );
    buf g4445 ( n26480 , n32572 );
    or g4446 ( n22775 , n35401 , n1402 );
    or g4447 ( n5175 , n7322 , n21977 );
    xnor g4448 ( n30745 , n25978 , n11801 );
    or g4449 ( n9737 , n11334 , n27171 );
    or g4450 ( n7554 , n4771 , n34472 );
    or g4451 ( n20259 , n25473 , n2005 );
    xnor g4452 ( n4038 , n22982 , n24864 );
    xnor g4453 ( n741 , n5942 , n27929 );
    or g4454 ( n26828 , n14730 , n16797 );
    xnor g4455 ( n10201 , n35104 , n4695 );
    xnor g4456 ( n12881 , n6231 , n3774 );
    xnor g4457 ( n28849 , n15906 , n18638 );
    and g4458 ( n17907 , n20868 , n31480 );
    xnor g4459 ( n23849 , n23010 , n35927 );
    or g4460 ( n12347 , n30581 , n6689 );
    or g4461 ( n30900 , n6516 , n20300 );
    nor g4462 ( n5228 , n29713 , n31947 );
    or g4463 ( n4408 , n10894 , n29010 );
    not g4464 ( n10531 , n32424 );
    or g4465 ( n8512 , n6731 , n9240 );
    xnor g4466 ( n12729 , n27227 , n17799 );
    not g4467 ( n4983 , n16620 );
    xnor g4468 ( n6125 , n6735 , n7540 );
    and g4469 ( n15394 , n23395 , n11262 );
    not g4470 ( n12107 , n12460 );
    nor g4471 ( n16116 , n22291 , n29287 );
    xor g4472 ( n19565 , n73 , n21323 );
    xnor g4473 ( n1758 , n29778 , n25673 );
    or g4474 ( n10111 , n30729 , n8203 );
    xnor g4475 ( n5568 , n16657 , n35838 );
    or g4476 ( n15146 , n19485 , n9601 );
    or g4477 ( n26085 , n29920 , n23225 );
    and g4478 ( n4668 , n9444 , n11729 );
    or g4479 ( n8029 , n6885 , n2119 );
    or g4480 ( n11101 , n26280 , n8276 );
    or g4481 ( n7908 , n10894 , n23959 );
    xnor g4482 ( n33780 , n15565 , n15886 );
    or g4483 ( n10576 , n26161 , n34687 );
    or g4484 ( n14750 , n3222 , n15987 );
    or g4485 ( n27712 , n24981 , n17004 );
    or g4486 ( n27313 , n32715 , n3284 );
    and g4487 ( n21884 , n32150 , n5471 );
    not g4488 ( n8511 , n13612 );
    not g4489 ( n1641 , n33041 );
    or g4490 ( n19030 , n10369 , n8259 );
    nor g4491 ( n12983 , n11023 , n32356 );
    or g4492 ( n4275 , n26391 , n23278 );
    and g4493 ( n12912 , n15582 , n12303 );
    nor g4494 ( n23249 , n12696 , n19373 );
    or g4495 ( n1668 , n22798 , n20812 );
    xnor g4496 ( n29791 , n34728 , n32335 );
    xnor g4497 ( n3033 , n20688 , n31784 );
    and g4498 ( n21223 , n25615 , n32548 );
    nor g4499 ( n2505 , n3205 , n34434 );
    and g4500 ( n12201 , n34167 , n19301 );
    and g4501 ( n34985 , n11860 , n8146 );
    xnor g4502 ( n29719 , n12947 , n15464 );
    xnor g4503 ( n5977 , n17353 , n22291 );
    or g4504 ( n21340 , n23241 , n30708 );
    and g4505 ( n10418 , n22902 , n14413 );
    or g4506 ( n2464 , n29557 , n8392 );
    xnor g4507 ( n18442 , n27943 , n4758 );
    or g4508 ( n20134 , n31806 , n4172 );
    and g4509 ( n12389 , n35215 , n2558 );
    not g4510 ( n16293 , n35927 );
    or g4511 ( n16322 , n27070 , n5252 );
    nor g4512 ( n30235 , n9658 , n9523 );
    and g4513 ( n7113 , n5528 , n9012 );
    xnor g4514 ( n5464 , n33652 , n32095 );
    or g4515 ( n27364 , n4288 , n15962 );
    and g4516 ( n32239 , n22000 , n3297 );
    or g4517 ( n4963 , n19984 , n10001 );
    and g4518 ( n14798 , n34799 , n21586 );
    nor g4519 ( n11066 , n25174 , n19590 );
    and g4520 ( n31261 , n2411 , n25124 );
    and g4521 ( n4416 , n13579 , n12687 );
    or g4522 ( n30171 , n18297 , n11712 );
    and g4523 ( n4639 , n21767 , n15687 );
    and g4524 ( n10862 , n27744 , n4252 );
    not g4525 ( n14666 , n2292 );
    xnor g4526 ( n3385 , n2089 , n12973 );
    and g4527 ( n12447 , n17760 , n20538 );
    xnor g4528 ( n7496 , n33056 , n22291 );
    or g4529 ( n32980 , n6440 , n27113 );
    or g4530 ( n32548 , n32857 , n35727 );
    and g4531 ( n8277 , n31818 , n1544 );
    or g4532 ( n14398 , n23608 , n25392 );
    or g4533 ( n24888 , n17591 , n10823 );
    or g4534 ( n35906 , n10008 , n18477 );
    and g4535 ( n29810 , n35742 , n15661 );
    and g4536 ( n7847 , n6450 , n35147 );
    or g4537 ( n5569 , n6861 , n8924 );
    and g4538 ( n22003 , n23167 , n6575 );
    and g4539 ( n34214 , n32048 , n15244 );
    xnor g4540 ( n21930 , n31875 , n21490 );
    and g4541 ( n14119 , n5725 , n34377 );
    or g4542 ( n7109 , n3205 , n6864 );
    nor g4543 ( n35492 , n33279 , n13883 );
    or g4544 ( n17688 , n17713 , n28675 );
    or g4545 ( n24449 , n13663 , n10229 );
    nor g4546 ( n1972 , n5335 , n36019 );
    and g4547 ( n27043 , n35957 , n34726 );
    or g4548 ( n13993 , n917 , n22224 );
    xnor g4549 ( n9683 , n22944 , n31289 );
    xnor g4550 ( n30546 , n17562 , n8432 );
    and g4551 ( n16690 , n13468 , n31323 );
    or g4552 ( n17165 , n296 , n10400 );
    not g4553 ( n33224 , n9435 );
    or g4554 ( n29435 , n24221 , n11295 );
    nor g4555 ( n8181 , n12647 , n10533 );
    not g4556 ( n26728 , n14420 );
    or g4557 ( n28732 , n11046 , n16641 );
    and g4558 ( n29818 , n21284 , n3147 );
    or g4559 ( n27019 , n4396 , n9091 );
    and g4560 ( n1264 , n19342 , n29817 );
    and g4561 ( n29418 , n27900 , n28131 );
    nor g4562 ( n20932 , n21 , n19904 );
    not g4563 ( n3685 , n9361 );
    and g4564 ( n35164 , n33860 , n15516 );
    or g4565 ( n28949 , n17422 , n32329 );
    and g4566 ( n15157 , n18089 , n13369 );
    or g4567 ( n32754 , n19136 , n26002 );
    xnor g4568 ( n19709 , n18181 , n5289 );
    or g4569 ( n19673 , n15767 , n16086 );
    or g4570 ( n21471 , n10401 , n8913 );
    xnor g4571 ( n21132 , n14958 , n25602 );
    or g4572 ( n5059 , n15887 , n34869 );
    and g4573 ( n13130 , n16727 , n10494 );
    xnor g4574 ( n2656 , n4682 , n27177 );
    or g4575 ( n16334 , n21981 , n8392 );
    xnor g4576 ( n25218 , n6915 , n3222 );
    and g4577 ( n24941 , n32784 , n11582 );
    nor g4578 ( n34695 , n6518 , n6104 );
    and g4579 ( n2462 , n6969 , n17420 );
    and g4580 ( n20869 , n5500 , n25703 );
    not g4581 ( n7569 , n26731 );
    xnor g4582 ( n22697 , n9664 , n3275 );
    not g4583 ( n5965 , n26756 );
    or g4584 ( n20135 , n20258 , n20690 );
    not g4585 ( n29941 , n14132 );
    and g4586 ( n16124 , n28754 , n3203 );
    xnor g4587 ( n6375 , n4002 , n32278 );
    xnor g4588 ( n21205 , n32940 , n7861 );
    xnor g4589 ( n27532 , n34965 , n4960 );
    and g4590 ( n5263 , n5196 , n14392 );
    or g4591 ( n34645 , n7396 , n5941 );
    or g4592 ( n29227 , n28180 , n26974 );
    xnor g4593 ( n15142 , n22457 , n30553 );
    and g4594 ( n15278 , n34877 , n7403 );
    and g4595 ( n11569 , n1431 , n16126 );
    or g4596 ( n20365 , n27202 , n14145 );
    or g4597 ( n19727 , n35529 , n23492 );
    not g4598 ( n22646 , n8923 );
    xnor g4599 ( n31267 , n32160 , n4288 );
    and g4600 ( n9024 , n25437 , n35462 );
    and g4601 ( n19451 , n2243 , n10495 );
    nor g4602 ( n18443 , n1786 , n10913 );
    or g4603 ( n2349 , n6137 , n31514 );
    xnor g4604 ( n11535 , n22056 , n28934 );
    not g4605 ( n19010 , n13421 );
    or g4606 ( n33243 , n25870 , n12434 );
    or g4607 ( n30387 , n32857 , n22154 );
    xnor g4608 ( n17437 , n1584 , n35223 );
    and g4609 ( n1295 , n30403 , n2135 );
    and g4610 ( n8418 , n22108 , n15485 );
    and g4611 ( n34955 , n6709 , n9656 );
    not g4612 ( n51 , n6288 );
    not g4613 ( n1873 , n13358 );
    and g4614 ( n5786 , n7478 , n32395 );
    or g4615 ( n20949 , n28123 , n14791 );
    or g4616 ( n9272 , n17716 , n25392 );
    or g4617 ( n11672 , n22067 , n287 );
    or g4618 ( n30547 , n23098 , n3738 );
    and g4619 ( n11001 , n24256 , n29017 );
    xnor g4620 ( n20804 , n19494 , n35099 );
    xnor g4621 ( n958 , n416 , n31687 );
    nor g4622 ( n26189 , n22990 , n1121 );
    and g4623 ( n24539 , n32142 , n12113 );
    or g4624 ( n22805 , n32857 , n13275 );
    or g4625 ( n11687 , n10784 , n12879 );
    xnor g4626 ( n11284 , n8131 , n27536 );
    xnor g4627 ( n34175 , n3141 , n4962 );
    nor g4628 ( n0 , n15886 , n18270 );
    xnor g4629 ( n2803 , n4905 , n22291 );
    xnor g4630 ( n9640 , n22406 , n35509 );
    or g4631 ( n26858 , n830 , n32531 );
    or g4632 ( n20860 , n1639 , n10417 );
    and g4633 ( n20827 , n3261 , n31294 );
    or g4634 ( n25685 , n3421 , n6340 );
    and g4635 ( n23846 , n7451 , n30601 );
    xnor g4636 ( n18020 , n15412 , n13768 );
    xor g4637 ( n28879 , n29331 , n34403 );
    nor g4638 ( n8682 , n16370 , n17829 );
    xnor g4639 ( n29034 , n23749 , n15464 );
    nor g4640 ( n1617 , n11046 , n18238 );
    and g4641 ( n14489 , n20144 , n13108 );
    not g4642 ( n5332 , n27156 );
    or g4643 ( n29621 , n33455 , n15568 );
    and g4644 ( n7876 , n5870 , n14679 );
    xnor g4645 ( n16384 , n2876 , n11455 );
    or g4646 ( n29025 , n35955 , n10630 );
    and g4647 ( n29998 , n13964 , n3077 );
    not g4648 ( n12652 , n11455 );
    or g4649 ( n35887 , n31272 , n17500 );
    and g4650 ( n725 , n28395 , n14346 );
    xnor g4651 ( n20907 , n6290 , n16500 );
    buf g4652 ( n1796 , n16649 );
    nor g4653 ( n16305 , n10072 , n24566 );
    xnor g4654 ( n22412 , n17390 , n7540 );
    not g4655 ( n27998 , n18278 );
    or g4656 ( n26017 , n27196 , n32576 );
    xnor g4657 ( n28022 , n11501 , n4960 );
    or g4658 ( n20410 , n35927 , n9576 );
    nor g4659 ( n29356 , n35666 , n1176 );
    xnor g4660 ( n293 , n25041 , n19551 );
    not g4661 ( n33962 , n19602 );
    nor g4662 ( n8254 , n10981 , n31964 );
    not g4663 ( n12547 , n1552 );
    or g4664 ( n9677 , n32935 , n17974 );
    and g4665 ( n17827 , n21390 , n17973 );
    xnor g4666 ( n6403 , n33927 , n2727 );
    nor g4667 ( n2508 , n4896 , n34015 );
    not g4668 ( n5820 , n24957 );
    nor g4669 ( n24362 , n32611 , n29366 );
    nor g4670 ( n15648 , n25602 , n1625 );
    xnor g4671 ( n30342 , n26849 , n32095 );
    and g4672 ( n28066 , n9573 , n20740 );
    and g4673 ( n24415 , n4459 , n10661 );
    or g4674 ( n4862 , n25828 , n28887 );
    and g4675 ( n7170 , n30612 , n5484 );
    and g4676 ( n20492 , n23100 , n11365 );
    xnor g4677 ( n2329 , n17457 , n9958 );
    or g4678 ( n27335 , n3205 , n18063 );
    or g4679 ( n14493 , n6348 , n33761 );
    xnor g4680 ( n27120 , n9204 , n35927 );
    or g4681 ( n15199 , n3081 , n35402 );
    not g4682 ( n19422 , n1127 );
    or g4683 ( n33035 , n14840 , n21002 );
    xnor g4684 ( n2240 , n29732 , n29555 );
    or g4685 ( n24850 , n28354 , n1474 );
    or g4686 ( n2059 , n5912 , n34038 );
    or g4687 ( n2885 , n5676 , n12149 );
    or g4688 ( n29186 , n19984 , n5190 );
    or g4689 ( n29473 , n4177 , n11850 );
    or g4690 ( n25935 , n14578 , n1557 );
    xnor g4691 ( n19346 , n21798 , n15886 );
    and g4692 ( n4285 , n7334 , n10927 );
    xnor g4693 ( n14280 , n2192 , n24130 );
    not g4694 ( n8683 , n27176 );
    nor g4695 ( n16824 , n5214 , n35518 );
    not g4696 ( n13374 , n3243 );
    or g4697 ( n13066 , n8425 , n27253 );
    and g4698 ( n1435 , n26071 , n20117 );
    xnor g4699 ( n12162 , n16081 , n16620 );
    and g4700 ( n5161 , n17960 , n7593 );
    xnor g4701 ( n33094 , n26956 , n27960 );
    and g4702 ( n15649 , n29423 , n24014 );
    and g4703 ( n10739 , n25971 , n18108 );
    xnor g4704 ( n12932 , n611 , n9253 );
    xnor g4705 ( n30862 , n7284 , n14427 );
    or g4706 ( n15927 , n20213 , n35111 );
    or g4707 ( n28201 , n15074 , n5337 );
    or g4708 ( n34146 , n8672 , n2823 );
    not g4709 ( n17674 , n22871 );
    or g4710 ( n33477 , n9735 , n4895 );
    or g4711 ( n5934 , n1365 , n13217 );
    or g4712 ( n10687 , n16670 , n28668 );
    or g4713 ( n26034 , n9220 , n27963 );
    and g4714 ( n35507 , n21736 , n15708 );
    or g4715 ( n19517 , n8712 , n21486 );
    xnor g4716 ( n4825 , n12354 , n7540 );
    or g4717 ( n11988 , n10102 , n17695 );
    and g4718 ( n30774 , n18900 , n19320 );
    not g4719 ( n11874 , n8378 );
    xnor g4720 ( n15771 , n35495 , n20045 );
    xnor g4721 ( n19621 , n4826 , n24371 );
    and g4722 ( n19077 , n23955 , n18854 );
    or g4723 ( n12303 , n32715 , n10999 );
    xnor g4724 ( n5374 , n9820 , n25602 );
    xnor g4725 ( n31954 , n473 , n32388 );
    xnor g4726 ( n29558 , n1378 , n32095 );
    and g4727 ( n8354 , n29645 , n2129 );
    not g4728 ( n2718 , n27422 );
    or g4729 ( n4119 , n26505 , n6133 );
    or g4730 ( n15661 , n11046 , n27710 );
    or g4731 ( n14825 , n16222 , n11977 );
    not g4732 ( n18635 , n14597 );
    not g4733 ( n17592 , n23953 );
    nor g4734 ( n12080 , n30742 , n10514 );
    or g4735 ( n10541 , n33121 , n22339 );
    xnor g4736 ( n24251 , n4938 , n29713 );
    xnor g4737 ( n16487 , n11018 , n19260 );
    or g4738 ( n14524 , n24332 , n3443 );
    and g4739 ( n11980 , n8785 , n26552 );
    or g4740 ( n12383 , n23250 , n24254 );
    or g4741 ( n32131 , n25602 , n8775 );
    not g4742 ( n34853 , n2650 );
    or g4743 ( n26943 , n15299 , n23678 );
    or g4744 ( n25152 , n10636 , n33642 );
    and g4745 ( n31558 , n29927 , n33834 );
    or g4746 ( n8507 , n20209 , n35451 );
    or g4747 ( n8036 , n11008 , n8877 );
    xnor g4748 ( n16215 , n23245 , n7540 );
    or g4749 ( n17507 , n10894 , n7195 );
    xnor g4750 ( n22075 , n20071 , n20310 );
    or g4751 ( n843 , n19908 , n35313 );
    and g4752 ( n27870 , n35092 , n19226 );
    nor g4753 ( n34287 , n8232 , n27947 );
    and g4754 ( n35516 , n9769 , n18557 );
    not g4755 ( n15001 , n7101 );
    xnor g4756 ( n22877 , n28938 , n22291 );
    xnor g4757 ( n22302 , n14816 , n16620 );
    or g4758 ( n11198 , n12565 , n17974 );
    or g4759 ( n23152 , n8606 , n11977 );
    xnor g4760 ( n30254 , n35052 , n14286 );
    not g4761 ( n26951 , n19033 );
    or g4762 ( n28672 , n18338 , n27056 );
    nor g4763 ( n12034 , n8777 , n28072 );
    and g4764 ( n3628 , n20861 , n17260 );
    and g4765 ( n33757 , n30971 , n9508 );
    xnor g4766 ( n16699 , n6598 , n24500 );
    xnor g4767 ( n22277 , n16842 , n24846 );
    xnor g4768 ( n18875 , n505 , n4960 );
    not g4769 ( n27396 , n16217 );
    and g4770 ( n28106 , n27316 , n14928 );
    xnor g4771 ( n9722 , n28345 , n33901 );
    or g4772 ( n10985 , n33974 , n28191 );
    or g4773 ( n12534 , n3974 , n669 );
    not g4774 ( n95 , n4878 );
    and g4775 ( n19319 , n28459 , n25823 );
    and g4776 ( n20048 , n23097 , n28359 );
    xnor g4777 ( n5553 , n7881 , n32095 );
    or g4778 ( n27666 , n24530 , n2479 );
    or g4779 ( n14181 , n34595 , n22519 );
    or g4780 ( n31115 , n10138 , n14146 );
    and g4781 ( n4858 , n1044 , n13417 );
    xnor g4782 ( n32478 , n14943 , n17751 );
    or g4783 ( n12501 , n31127 , n35992 );
    and g4784 ( n34491 , n3402 , n22034 );
    or g4785 ( n25876 , n19457 , n4490 );
    nor g4786 ( n24187 , n25602 , n33670 );
    or g4787 ( n22748 , n9658 , n28713 );
    and g4788 ( n15985 , n12691 , n6863 );
    nor g4789 ( n14651 , n30020 , n13943 );
    or g4790 ( n26288 , n31972 , n2749 );
    or g4791 ( n15954 , n25602 , n32382 );
    or g4792 ( n3538 , n32232 , n10341 );
    or g4793 ( n17552 , n7826 , n35148 );
    not g4794 ( n23147 , n15886 );
    or g4795 ( n15390 , n1321 , n31182 );
    and g4796 ( n19401 , n32920 , n34910 );
    nor g4797 ( n8338 , n4960 , n29617 );
    or g4798 ( n6249 , n16582 , n27447 );
    not g4799 ( n23 , n14530 );
    xnor g4800 ( n9397 , n30097 , n21351 );
    not g4801 ( n28045 , n5446 );
    nor g4802 ( n16561 , n7540 , n14354 );
    or g4803 ( n34589 , n26272 , n34084 );
    or g4804 ( n12176 , n27125 , n1642 );
    and g4805 ( n15150 , n32578 , n23693 );
    xnor g4806 ( n30032 , n15926 , n17308 );
    or g4807 ( n16524 , n31025 , n23170 );
    or g4808 ( n19853 , n25176 , n5457 );
    and g4809 ( n564 , n17511 , n26739 );
    not g4810 ( n19435 , n714 );
    or g4811 ( n14175 , n16620 , n29031 );
    or g4812 ( n16630 , n3222 , n26175 );
    or g4813 ( n31213 , n14882 , n5501 );
    or g4814 ( n2566 , n25779 , n1796 );
    and g4815 ( n3458 , n29282 , n30101 );
    or g4816 ( n7694 , n15973 , n23450 );
    or g4817 ( n23141 , n16671 , n27625 );
    not g4818 ( n28141 , n2686 );
    not g4819 ( n26110 , n93 );
    nor g4820 ( n7123 , n28942 , n22124 );
    or g4821 ( n17424 , n9793 , n29614 );
    nor g4822 ( n34344 , n12024 , n33157 );
    and g4823 ( n14727 , n4368 , n3148 );
    xnor g4824 ( n18561 , n20870 , n25174 );
    xnor g4825 ( n33847 , n5977 , n29132 );
    or g4826 ( n28079 , n30613 , n16600 );
    or g4827 ( n20167 , n16114 , n10417 );
    xnor g4828 ( n28180 , n33911 , n23604 );
    and g4829 ( n3931 , n16099 , n326 );
    nor g4830 ( n8355 , n4878 , n2468 );
    and g4831 ( n27116 , n31088 , n33253 );
    or g4832 ( n22660 , n17558 , n3352 );
    nor g4833 ( n5754 , n4962 , n13244 );
    or g4834 ( n170 , n17751 , n1072 );
    xnor g4835 ( n25208 , n17606 , n32624 );
    or g4836 ( n34833 , n18750 , n17742 );
    nor g4837 ( n23217 , n25070 , n27753 );
    nor g4838 ( n2374 , n30792 , n799 );
    xnor g4839 ( n12509 , n24020 , n5492 );
    or g4840 ( n35225 , n3573 , n24893 );
    and g4841 ( n8167 , n22469 , n7017 );
    or g4842 ( n33315 , n13162 , n21873 );
    or g4843 ( n14474 , n20816 , n1511 );
    xnor g4844 ( n25893 , n11567 , n4960 );
    and g4845 ( n21338 , n27888 , n21362 );
    not g4846 ( n12796 , n24212 );
    or g4847 ( n4593 , n32095 , n12850 );
    not g4848 ( n33989 , n26502 );
    not g4849 ( n3438 , n28866 );
    and g4850 ( n32546 , n11843 , n25504 );
    not g4851 ( n6584 , n18414 );
    nor g4852 ( n10299 , n2527 , n17687 );
    or g4853 ( n24915 , n11144 , n24333 );
    or g4854 ( n22410 , n26314 , n10762 );
    xnor g4855 ( n31191 , n31394 , n4590 );
    or g4856 ( n22629 , n30742 , n3278 );
    and g4857 ( n35746 , n28338 , n16890 );
    xnor g4858 ( n2345 , n32229 , n5738 );
    and g4859 ( n28713 , n9839 , n27142 );
    or g4860 ( n6517 , n18508 , n19652 );
    xnor g4861 ( n13291 , n26449 , n4288 );
    and g4862 ( n17785 , n25796 , n9456 );
    and g4863 ( n6435 , n5790 , n2582 );
    xnor g4864 ( n12392 , n3157 , n16620 );
    nor g4865 ( n33298 , n19551 , n7282 );
    or g4866 ( n30271 , n15464 , n1591 );
    or g4867 ( n8762 , n32584 , n27125 );
    or g4868 ( n26739 , n4288 , n29559 );
    xnor g4869 ( n29183 , n23992 , n32197 );
    or g4870 ( n27469 , n22633 , n15952 );
    or g4871 ( n28077 , n22755 , n16622 );
    xnor g4872 ( n11490 , n12628 , n11493 );
    or g4873 ( n22662 , n3975 , n3019 );
    or g4874 ( n23682 , n21232 , n2524 );
    or g4875 ( n32554 , n25804 , n12622 );
    or g4876 ( n1346 , n32748 , n26106 );
    or g4877 ( n32576 , n13088 , n10701 );
    xnor g4878 ( n28796 , n5931 , n11194 );
    nor g4879 ( n20064 , n9789 , n28106 );
    or g4880 ( n31443 , n4962 , n9923 );
    and g4881 ( n15894 , n15425 , n14134 );
    and g4882 ( n23729 , n13151 , n14028 );
    xnor g4883 ( n6861 , n16886 , n29020 );
    and g4884 ( n15969 , n6227 , n25182 );
    not g4885 ( n23990 , n27857 );
    not g4886 ( n23379 , n32411 );
    and g4887 ( n10718 , n29863 , n11076 );
    and g4888 ( n27763 , n12139 , n18714 );
    and g4889 ( n29873 , n10368 , n1794 );
    xnor g4890 ( n11829 , n29400 , n4297 );
    buf g4891 ( n18255 , n14611 );
    or g4892 ( n12219 , n28092 , n4043 );
    xnor g4893 ( n28052 , n16243 , n21237 );
    and g4894 ( n6821 , n15370 , n35818 );
    or g4895 ( n22588 , n31332 , n3437 );
    or g4896 ( n14828 , n16922 , n22571 );
    not g4897 ( n9410 , n25761 );
    or g4898 ( n29858 , n6375 , n9555 );
    or g4899 ( n33307 , n26941 , n18761 );
    or g4900 ( n31910 , n31068 , n19421 );
    or g4901 ( n11297 , n11634 , n8366 );
    and g4902 ( n17839 , n14867 , n1807 );
    and g4903 ( n21453 , n9144 , n17097 );
    or g4904 ( n2944 , n6694 , n8090 );
    not g4905 ( n17336 , n408 );
    xnor g4906 ( n11363 , n31955 , n9789 );
    xnor g4907 ( n10321 , n18597 , n1682 );
    or g4908 ( n19325 , n5490 , n10336 );
    and g4909 ( n7706 , n4119 , n10262 );
    and g4910 ( n5765 , n10763 , n16323 );
    and g4911 ( n23264 , n5597 , n11455 );
    xnor g4912 ( n34907 , n6807 , n11046 );
    or g4913 ( n20063 , n35008 , n32634 );
    or g4914 ( n31681 , n31295 , n15036 );
    or g4915 ( n22520 , n2259 , n16556 );
    or g4916 ( n18489 , n7559 , n10107 );
    and g4917 ( n25888 , n29051 , n7805 );
    and g4918 ( n15477 , n35387 , n18587 );
    and g4919 ( n35271 , n8646 , n15268 );
    nor g4920 ( n26205 , n26070 , n22061 );
    and g4921 ( n13361 , n21824 , n7078 );
    or g4922 ( n20896 , n33397 , n12332 );
    xnor g4923 ( n17206 , n29816 , n16331 );
    or g4924 ( n18539 , n19551 , n10021 );
    or g4925 ( n7341 , n23604 , n610 );
    or g4926 ( n30991 , n13007 , n29643 );
    xnor g4927 ( n34646 , n4209 , n9135 );
    and g4928 ( n28643 , n12020 , n9100 );
    xnor g4929 ( n19794 , n21083 , n32178 );
    not g4930 ( n31403 , n8471 );
    xnor g4931 ( n32832 , n6627 , n10587 );
    and g4932 ( n22814 , n19681 , n13448 );
    or g4933 ( n24293 , n5376 , n5868 );
    or g4934 ( n11457 , n23665 , n35141 );
    xnor g4935 ( n17433 , n26706 , n29839 );
    or g4936 ( n22058 , n30594 , n28710 );
    or g4937 ( n20815 , n10182 , n5317 );
    or g4938 ( n2213 , n9937 , n15290 );
    or g4939 ( n5134 , n12012 , n19490 );
    or g4940 ( n2929 , n25368 , n5168 );
    nor g4941 ( n17417 , n25602 , n30293 );
    or g4942 ( n3051 , n31679 , n16995 );
    or g4943 ( n30872 , n30716 , n13664 );
    and g4944 ( n16570 , n33221 , n23570 );
    or g4945 ( n35142 , n33573 , n4175 );
    or g4946 ( n22867 , n6140 , n32634 );
    or g4947 ( n34197 , n32412 , n26000 );
    xnor g4948 ( n19661 , n28509 , n15501 );
    or g4949 ( n26426 , n35814 , n19653 );
    or g4950 ( n9353 , n19956 , n3634 );
    or g4951 ( n4509 , n6437 , n25306 );
    xnor g4952 ( n342 , n14785 , n18379 );
    and g4953 ( n24963 , n3107 , n27967 );
    or g4954 ( n24152 , n1446 , n28574 );
    or g4955 ( n17317 , n8820 , n3386 );
    or g4956 ( n29386 , n15886 , n17750 );
    not g4957 ( n6347 , n653 );
    or g4958 ( n14937 , n21072 , n21880 );
    and g4959 ( n28696 , n32025 , n9234 );
    and g4960 ( n18203 , n13378 , n2737 );
    or g4961 ( n14339 , n14097 , n28526 );
    xnor g4962 ( n18848 , n15734 , n24163 );
    xnor g4963 ( n1555 , n32061 , n27912 );
    not g4964 ( n4760 , n16262 );
    xor g4965 ( n482 , n3404 , n31478 );
    and g4966 ( n27174 , n26964 , n31450 );
    or g4967 ( n27382 , n19740 , n25019 );
    xnor g4968 ( n17923 , n425 , n24371 );
    and g4969 ( n26966 , n11230 , n28823 );
    xor g4970 ( n5963 , n3545 , n22302 );
    xnor g4971 ( n6647 , n19926 , n30983 );
    or g4972 ( n24470 , n35947 , n15538 );
    or g4973 ( n21211 , n19551 , n27739 );
    or g4974 ( n31016 , n22449 , n850 );
    or g4975 ( n10781 , n17510 , n26483 );
    and g4976 ( n22626 , n5889 , n35828 );
    and g4977 ( n4113 , n9843 , n16032 );
    xnor g4978 ( n23768 , n32295 , n1950 );
    xnor g4979 ( n2795 , n30393 , n9793 );
    not g4980 ( n10573 , n30742 );
    xnor g4981 ( n30452 , n22308 , n28396 );
    and g4982 ( n10292 , n5349 , n27035 );
    xnor g4983 ( n10143 , n25627 , n11980 );
    or g4984 ( n27881 , n18618 , n5972 );
    not g4985 ( n3236 , n17751 );
    and g4986 ( n30313 , n12536 , n22392 );
    nor g4987 ( n23830 , n10894 , n4785 );
    or g4988 ( n1064 , n17896 , n21675 );
    or g4989 ( n31667 , n3590 , n9999 );
    and g4990 ( n16538 , n2855 , n28775 );
    xnor g4991 ( n34444 , n35853 , n15025 );
    xnor g4992 ( n30961 , n30373 , n13433 );
    and g4993 ( n3647 , n5827 , n2809 );
    and g4994 ( n35665 , n28511 , n22821 );
    nor g4995 ( n33905 , n7540 , n25699 );
    or g4996 ( n9393 , n27416 , n1474 );
    nor g4997 ( n1750 , n26056 , n19834 );
    or g4998 ( n27184 , n768 , n9672 );
    xnor g4999 ( n19494 , n35369 , n36049 );
    not g5000 ( n12516 , n4878 );
    or g5001 ( n26554 , n5313 , n31554 );
    not g5002 ( n34161 , n9793 );
    xnor g5003 ( n24237 , n33648 , n24371 );
    or g5004 ( n20612 , n21852 , n13077 );
    xnor g5005 ( n1612 , n18262 , n4329 );
    or g5006 ( n30640 , n7925 , n35644 );
    or g5007 ( n4586 , n17568 , n3128 );
    or g5008 ( n26092 , n24021 , n31282 );
    or g5009 ( n22557 , n22346 , n35132 );
    nor g5010 ( n5023 , n26587 , n189 );
    or g5011 ( n21749 , n11455 , n2876 );
    and g5012 ( n12252 , n5130 , n1043 );
    and g5013 ( n6502 , n29403 , n16189 );
    xnor g5014 ( n33066 , n838 , n10894 );
    or g5015 ( n21475 , n11111 , n29229 );
    or g5016 ( n1977 , n9565 , n34923 );
    and g5017 ( n21200 , n16732 , n26297 );
    xnor g5018 ( n5021 , n13154 , n12340 );
    or g5019 ( n32175 , n3946 , n11760 );
    or g5020 ( n4402 , n26760 , n26931 );
    xnor g5021 ( n23093 , n11634 , n30253 );
    or g5022 ( n33230 , n25602 , n15235 );
    xnor g5023 ( n1152 , n14294 , n8240 );
    or g5024 ( n8591 , n19949 , n4772 );
    xnor g5025 ( n11555 , n13513 , n9024 );
    and g5026 ( n6796 , n24910 , n4786 );
    or g5027 ( n34422 , n31289 , n17139 );
    nor g5028 ( n20417 , n17751 , n34717 );
    not g5029 ( n31590 , n3226 );
    xnor g5030 ( n30180 , n14744 , n23604 );
    or g5031 ( n24734 , n16860 , n22783 );
    or g5032 ( n28078 , n28700 , n6682 );
    xnor g5033 ( n26500 , n32341 , n16875 );
    or g5034 ( n32161 , n11396 , n9069 );
    or g5035 ( n28699 , n11933 , n1314 );
    and g5036 ( n4707 , n10291 , n5407 );
    xnor g5037 ( n21228 , n3650 , n18630 );
    not g5038 ( n25792 , n23407 );
    or g5039 ( n15948 , n19466 , n35402 );
    xnor g5040 ( n9247 , n28308 , n10894 );
    and g5041 ( n34119 , n24668 , n28057 );
    nor g5042 ( n27024 , n29713 , n7140 );
    or g5043 ( n24492 , n32823 , n24672 );
    and g5044 ( n7733 , n322 , n16012 );
    xnor g5045 ( n17445 , n27353 , n31289 );
    or g5046 ( n19869 , n15540 , n34036 );
    and g5047 ( n16382 , n18678 , n28196 );
    nor g5048 ( n29940 , n3205 , n33752 );
    and g5049 ( n35148 , n3083 , n9471 );
    nor g5050 ( n7873 , n15464 , n2024 );
    xnor g5051 ( n20246 , n9179 , n11578 );
    or g5052 ( n19016 , n13575 , n6936 );
    not g5053 ( n1762 , n328 );
    nor g5054 ( n32766 , n9984 , n21964 );
    not g5055 ( n21873 , n25761 );
    and g5056 ( n24940 , n13100 , n16815 );
    not g5057 ( n10183 , n6024 );
    xnor g5058 ( n11084 , n20787 , n28513 );
    or g5059 ( n3987 , n33990 , n393 );
    xnor g5060 ( n8230 , n10454 , n174 );
    and g5061 ( n3088 , n27904 , n125 );
    not g5062 ( n2540 , n25472 );
    xnor g5063 ( n23091 , n22370 , n5335 );
    xnor g5064 ( n28614 , n17585 , n21419 );
    or g5065 ( n28681 , n29508 , n2712 );
    xnor g5066 ( n3078 , n6427 , n4878 );
    and g5067 ( n24679 , n34042 , n29190 );
    or g5068 ( n16400 , n21485 , n30978 );
    not g5069 ( n22124 , n29560 );
    or g5070 ( n14195 , n25745 , n23090 );
    or g5071 ( n28714 , n9918 , n27447 );
    or g5072 ( n18888 , n19984 , n12136 );
    not g5073 ( n14258 , n8628 );
    or g5074 ( n13293 , n2379 , n5905 );
    xnor g5075 ( n1665 , n9627 , n33892 );
    not g5076 ( n3810 , n7941 );
    or g5077 ( n25031 , n7259 , n3310 );
    and g5078 ( n33649 , n17053 , n7570 );
    xnor g5079 ( n3097 , n8935 , n8144 );
    xnor g5080 ( n25170 , n12192 , n32034 );
    and g5081 ( n24820 , n23042 , n13932 );
    or g5082 ( n11500 , n11415 , n25447 );
    or g5083 ( n25724 , n26029 , n31768 );
    not g5084 ( n14486 , n20558 );
    and g5085 ( n6958 , n24667 , n20497 );
    or g5086 ( n34652 , n34331 , n20812 );
    or g5087 ( n5641 , n36055 , n21977 );
    and g5088 ( n5428 , n7497 , n3874 );
    not g5089 ( n2527 , n31125 );
    xnor g5090 ( n18847 , n32538 , n11455 );
    and g5091 ( n34014 , n123 , n147 );
    or g5092 ( n11436 , n18403 , n2712 );
    not g5093 ( n7089 , n24341 );
    or g5094 ( n6250 , n22291 , n21234 );
    and g5095 ( n11901 , n5406 , n24428 );
    or g5096 ( n523 , n25174 , n31492 );
    nor g5097 ( n3658 , n25602 , n34061 );
    and g5098 ( n35605 , n28328 , n6222 );
    and g5099 ( n30992 , n27569 , n25820 );
    or g5100 ( n34446 , n17751 , n636 );
    and g5101 ( n24160 , n31574 , n31305 );
    xnor g5102 ( n30835 , n34879 , n31024 );
    or g5103 ( n10053 , n31146 , n17111 );
    and g5104 ( n25466 , n15241 , n5643 );
    or g5105 ( n13434 , n17293 , n23462 );
    and g5106 ( n23128 , n3161 , n17846 );
    and g5107 ( n8674 , n18128 , n32791 );
    or g5108 ( n18042 , n14553 , n3979 );
    or g5109 ( n21637 , n10101 , n2501 );
    or g5110 ( n17527 , n31953 , n17354 );
    or g5111 ( n7193 , n1950 , n15157 );
    or g5112 ( n8947 , n35808 , n13480 );
    or g5113 ( n1879 , n32715 , n30659 );
    xnor g5114 ( n19761 , n24314 , n25751 );
    and g5115 ( n26960 , n27720 , n20008 );
    nor g5116 ( n21708 , n8432 , n30207 );
    or g5117 ( n26367 , n29918 , n10331 );
    xnor g5118 ( n21660 , n13158 , n31799 );
    or g5119 ( n14395 , n19820 , n18542 );
    or g5120 ( n16531 , n13167 , n22553 );
    or g5121 ( n4632 , n28250 , n24491 );
    and g5122 ( n29448 , n12368 , n24405 );
    xnor g5123 ( n35880 , n8613 , n19551 );
    and g5124 ( n478 , n10774 , n22078 );
    or g5125 ( n1890 , n31497 , n14877 );
    buf g5126 ( n3251 , n1761 );
    or g5127 ( n17891 , n8225 , n15889 );
    not g5128 ( n1250 , n3842 );
    or g5129 ( n29530 , n971 , n26569 );
    or g5130 ( n2279 , n26226 , n17978 );
    nor g5131 ( n55 , n24371 , n27811 );
    or g5132 ( n19006 , n9161 , n14903 );
    not g5133 ( n26296 , n8267 );
    xnor g5134 ( n7183 , n35995 , n5701 );
    xnor g5135 ( n35075 , n12127 , n3205 );
    and g5136 ( n18152 , n6326 , n23727 );
    or g5137 ( n26803 , n20955 , n34707 );
    or g5138 ( n19428 , n3316 , n34472 );
    or g5139 ( n28650 , n15691 , n32634 );
    xnor g5140 ( n12169 , n24131 , n26344 );
    xnor g5141 ( n23044 , n29728 , n33033 );
    or g5142 ( n10368 , n18580 , n11115 );
    or g5143 ( n17947 , n4709 , n11258 );
    or g5144 ( n30842 , n14340 , n30431 );
    or g5145 ( n5110 , n8164 , n11520 );
    or g5146 ( n35863 , n28309 , n578 );
    and g5147 ( n18433 , n10354 , n2768 );
    or g5148 ( n35129 , n22474 , n8416 );
    or g5149 ( n26975 , n9200 , n34045 );
    and g5150 ( n30207 , n13080 , n34120 );
    xnor g5151 ( n1358 , n35152 , n27243 );
    or g5152 ( n18206 , n3541 , n2005 );
    or g5153 ( n5380 , n10785 , n28191 );
    nor g5154 ( n23242 , n16571 , n25993 );
    or g5155 ( n22667 , n9847 , n34022 );
    or g5156 ( n326 , n29162 , n25940 );
    or g5157 ( n7749 , n31417 , n8490 );
    and g5158 ( n4314 , n24984 , n32488 );
    not g5159 ( n33542 , n16620 );
    and g5160 ( n28004 , n33330 , n35821 );
    or g5161 ( n35218 , n4369 , n17962 );
    or g5162 ( n18911 , n29839 , n12142 );
    xnor g5163 ( n20455 , n19424 , n7676 );
    xnor g5164 ( n20042 , n12581 , n19070 );
    xnor g5165 ( n32879 , n6528 , n19551 );
    xnor g5166 ( n26029 , n12653 , n31799 );
    not g5167 ( n26485 , n5635 );
    xnor g5168 ( n12441 , n3909 , n7706 );
    not g5169 ( n17408 , n10894 );
    not g5170 ( n22267 , n25442 );
    and g5171 ( n16539 , n20943 , n16289 );
    or g5172 ( n5357 , n20206 , n1715 );
    or g5173 ( n21912 , n10894 , n25342 );
    and g5174 ( n32294 , n22610 , n4288 );
    and g5175 ( n20173 , n2766 , n35678 );
    and g5176 ( n32883 , n32352 , n17840 );
    or g5177 ( n21607 , n11150 , n25594 );
    or g5178 ( n17053 , n29389 , n23757 );
    and g5179 ( n29395 , n31485 , n5893 );
    xnor g5180 ( n1439 , n14084 , n14331 );
    not g5181 ( n4769 , n17939 );
    not g5182 ( n30470 , n2533 );
    or g5183 ( n32524 , n16403 , n14918 );
    or g5184 ( n5057 , n24222 , n27447 );
    xnor g5185 ( n20311 , n15456 , n15464 );
    or g5186 ( n7581 , n34578 , n2524 );
    not g5187 ( n6349 , n4288 );
    or g5188 ( n17110 , n1377 , n24025 );
    xnor g5189 ( n29597 , n11550 , n24099 );
    or g5190 ( n28046 , n11963 , n14434 );
    and g5191 ( n29438 , n7060 , n22673 );
    xnor g5192 ( n30806 , n7238 , n28756 );
    and g5193 ( n4871 , n23263 , n5810 );
    xnor g5194 ( n28878 , n9516 , n27418 );
    xnor g5195 ( n2420 , n26671 , n5336 );
    or g5196 ( n4481 , n4183 , n1796 );
    not g5197 ( n4500 , n27275 );
    and g5198 ( n2834 , n3905 , n17850 );
    or g5199 ( n22085 , n14541 , n18588 );
    xnor g5200 ( n26168 , n17156 , n8649 );
    or g5201 ( n5479 , n4296 , n31134 );
    or g5202 ( n31129 , n28833 , n27172 );
    and g5203 ( n31075 , n13293 , n9372 );
    or g5204 ( n34449 , n20044 , n15144 );
    and g5205 ( n12500 , n2037 , n1950 );
    or g5206 ( n28947 , n1016 , n28842 );
    xnor g5207 ( n11335 , n2721 , n34781 );
    or g5208 ( n21530 , n9793 , n20937 );
    and g5209 ( n1785 , n21443 , n16597 );
    and g5210 ( n26930 , n18169 , n17659 );
    or g5211 ( n28573 , n926 , n20576 );
    or g5212 ( n2015 , n18606 , n35449 );
    xnor g5213 ( n25148 , n12083 , n25545 );
    or g5214 ( n10090 , n32715 , n24963 );
    or g5215 ( n16147 , n8432 , n11538 );
    xnor g5216 ( n10917 , n33507 , n5717 );
    nor g5217 ( n16503 , n7827 , n18264 );
    or g5218 ( n9307 , n11034 , n25831 );
    or g5219 ( n3459 , n12803 , n11312 );
    or g5220 ( n36057 , n10581 , n19125 );
    or g5221 ( n5686 , n15503 , n9731 );
    xnor g5222 ( n9062 , n3503 , n7373 );
    xnor g5223 ( n25798 , n18569 , n22432 );
    or g5224 ( n19964 , n27716 , n23090 );
    nor g5225 ( n33201 , n17406 , n14146 );
    or g5226 ( n4932 , n15311 , n19402 );
    or g5227 ( n23753 , n17677 , n27501 );
    and g5228 ( n10514 , n14015 , n30583 );
    or g5229 ( n30469 , n34320 , n4525 );
    xnor g5230 ( n34390 , n27346 , n10871 );
    xnor g5231 ( n20713 , n14174 , n31375 );
    xnor g5232 ( n2013 , n5214 , n35518 );
    or g5233 ( n34512 , n29649 , n1911 );
    nor g5234 ( n15188 , n11378 , n27635 );
    and g5235 ( n5546 , n565 , n28847 );
    or g5236 ( n33452 , n31617 , n2814 );
    not g5237 ( n17313 , n20840 );
    or g5238 ( n27368 , n7708 , n15538 );
    or g5239 ( n9368 , n14916 , n16115 );
    or g5240 ( n35221 , n11066 , n22789 );
    xnor g5241 ( n17563 , n8642 , n5149 );
    and g5242 ( n25435 , n32467 , n32594 );
    and g5243 ( n24004 , n1401 , n10024 );
    and g5244 ( n13287 , n32659 , n4703 );
    or g5245 ( n8883 , n25076 , n8153 );
    and g5246 ( n8953 , n13487 , n30977 );
    and g5247 ( n16272 , n28433 , n21467 );
    xnor g5248 ( n26665 , n33114 , n28398 );
    not g5249 ( n7327 , n9117 );
    or g5250 ( n758 , n32037 , n30519 );
    or g5251 ( n27837 , n29139 , n31902 );
    and g5252 ( n22869 , n6517 , n1559 );
    or g5253 ( n15770 , n15167 , n13482 );
    or g5254 ( n6284 , n22529 , n17111 );
    and g5255 ( n15800 , n12571 , n4810 );
    or g5256 ( n17917 , n32997 , n3716 );
    or g5257 ( n36076 , n4597 , n529 );
    or g5258 ( n29737 , n11469 , n13307 );
    or g5259 ( n13659 , n19182 , n28123 );
    or g5260 ( n27333 , n35447 , n26404 );
    or g5261 ( n9250 , n1149 , n28455 );
    or g5262 ( n24614 , n5478 , n25831 );
    or g5263 ( n33782 , n1418 , n14316 );
    and g5264 ( n5304 , n15765 , n18071 );
    or g5265 ( n25211 , n10955 , n2157 );
    and g5266 ( n33099 , n13778 , n4434 );
    not g5267 ( n24823 , n3205 );
    and g5268 ( n5327 , n34309 , n31121 );
    nor g5269 ( n23795 , n7058 , n29203 );
    and g5270 ( n12927 , n32757 , n2145 );
    xnor g5271 ( n28137 , n10965 , n10894 );
    buf g5272 ( n9975 , n31372 );
    and g5273 ( n668 , n30981 , n15466 );
    and g5274 ( n33533 , n21595 , n1615 );
    xnor g5275 ( n8978 , n15360 , n27356 );
    or g5276 ( n33111 , n29839 , n31750 );
    and g5277 ( n9349 , n26746 , n11504 );
    or g5278 ( n20499 , n5416 , n3979 );
    and g5279 ( n1764 , n11783 , n20135 );
    nor g5280 ( n25095 , n15731 , n33956 );
    xnor g5281 ( n16555 , n4263 , n26884 );
    and g5282 ( n12602 , n29601 , n577 );
    xnor g5283 ( n7418 , n35227 , n29884 );
    or g5284 ( n476 , n1808 , n19939 );
    or g5285 ( n2843 , n24896 , n5457 );
    or g5286 ( n9776 , n30158 , n19297 );
    and g5287 ( n25794 , n27105 , n2662 );
    and g5288 ( n3888 , n794 , n2649 );
    nor g5289 ( n29569 , n9145 , n5720 );
    xnor g5290 ( n15973 , n28261 , n9658 );
    or g5291 ( n11076 , n19984 , n3565 );
    and g5292 ( n9501 , n35528 , n30719 );
    or g5293 ( n27079 , n16886 , n29020 );
    not g5294 ( n8253 , n16223 );
    or g5295 ( n19342 , n12083 , n25545 );
    xnor g5296 ( n11854 , n36016 , n33161 );
    or g5297 ( n8519 , n9734 , n9930 );
    nor g5298 ( n4906 , n17568 , n19645 );
    xnor g5299 ( n25820 , n35923 , n24329 );
    xnor g5300 ( n13753 , n33405 , n17881 );
    or g5301 ( n33607 , n31044 , n9848 );
    xnor g5302 ( n1406 , n13802 , n4416 );
    or g5303 ( n21472 , n20461 , n17204 );
    and g5304 ( n26748 , n8806 , n17503 );
    and g5305 ( n26175 , n10053 , n11840 );
    xnor g5306 ( n22982 , n8045 , n15464 );
    or g5307 ( n20493 , n6053 , n1856 );
    and g5308 ( n9812 , n29394 , n5792 );
    or g5309 ( n26006 , n8686 , n12950 );
    or g5310 ( n26965 , n24924 , n33105 );
    and g5311 ( n1969 , n8287 , n22304 );
    xnor g5312 ( n16654 , n32772 , n4962 );
    or g5313 ( n34733 , n13521 , n3490 );
    not g5314 ( n10007 , n26485 );
    nor g5315 ( n13901 , n4500 , n22036 );
    or g5316 ( n34783 , n3997 , n21268 );
    or g5317 ( n15777 , n32857 , n27950 );
    not g5318 ( n21459 , n29713 );
    and g5319 ( n189 , n30111 , n2153 );
    and g5320 ( n17150 , n1077 , n2914 );
    not g5321 ( n29794 , n26722 );
    xnor g5322 ( n20820 , n23551 , n8704 );
    and g5323 ( n10749 , n18506 , n1205 );
    not g5324 ( n32089 , n27144 );
    or g5325 ( n31485 , n14401 , n27728 );
    and g5326 ( n27166 , n10037 , n21542 );
    nor g5327 ( n4789 , n32299 , n16649 );
    not g5328 ( n16770 , n34353 );
    nor g5329 ( n3901 , n23604 , n3813 );
    or g5330 ( n6657 , n1939 , n4871 );
    or g5331 ( n1508 , n6624 , n15256 );
    or g5332 ( n16484 , n5353 , n6336 );
    or g5333 ( n23610 , n2300 , n9832 );
    not g5334 ( n12953 , n25648 );
    or g5335 ( n5042 , n23604 , n27031 );
    and g5336 ( n35354 , n35352 , n16098 );
    or g5337 ( n19330 , n31771 , n13307 );
    or g5338 ( n17732 , n21277 , n29643 );
    not g5339 ( n8157 , n376 );
    or g5340 ( n1692 , n35927 , n9819 );
    or g5341 ( n12106 , n8432 , n20185 );
    or g5342 ( n4729 , n30866 , n4175 );
    nor g5343 ( n10990 , n4288 , n31843 );
    xnor g5344 ( n31808 , n20205 , n5455 );
    xnor g5345 ( n8625 , n5275 , n25602 );
    or g5346 ( n11298 , n1478 , n17223 );
    or g5347 ( n14037 , n16965 , n17286 );
    and g5348 ( n29549 , n27608 , n19492 );
    and g5349 ( n10767 , n31849 , n16201 );
    xnor g5350 ( n31506 , n34081 , n23071 );
    or g5351 ( n32467 , n13781 , n1474 );
    and g5352 ( n17725 , n3454 , n8693 );
    or g5353 ( n31325 , n17655 , n3239 );
    or g5354 ( n6862 , n24371 , n16834 );
    or g5355 ( n27634 , n20543 , n6075 );
    or g5356 ( n21041 , n30530 , n4490 );
    or g5357 ( n27971 , n32856 , n22946 );
    or g5358 ( n1354 , n7273 , n31773 );
    or g5359 ( n29479 , n29882 , n11312 );
    and g5360 ( n25317 , n15510 , n4251 );
    xnor g5361 ( n8384 , n27496 , n13463 );
    nor g5362 ( n21202 , n9870 , n21481 );
    or g5363 ( n3077 , n4288 , n18667 );
    nor g5364 ( n5926 , n12599 , n7601 );
    or g5365 ( n11641 , n18709 , n21732 );
    xnor g5366 ( n14763 , n29381 , n17568 );
    or g5367 ( n29057 , n32587 , n7962 );
    or g5368 ( n35201 , n16143 , n12179 );
    not g5369 ( n31502 , n35714 );
    and g5370 ( n31388 , n30392 , n231 );
    and g5371 ( n6966 , n2328 , n26564 );
    and g5372 ( n6660 , n1881 , n26657 );
    nor g5373 ( n13890 , n4960 , n17123 );
    and g5374 ( n18111 , n4397 , n29030 );
    and g5375 ( n21321 , n14852 , n15847 );
    and g5376 ( n35388 , n26193 , n3714 );
    or g5377 ( n12056 , n31799 , n8434 );
    or g5378 ( n25554 , n25602 , n19574 );
    xnor g5379 ( n1316 , n28051 , n4288 );
    not g5380 ( n11782 , n32857 );
    and g5381 ( n32217 , n17217 , n6428 );
    not g5382 ( n27756 , n28866 );
    or g5383 ( n5445 , n24824 , n33382 );
    and g5384 ( n23360 , n33194 , n9185 );
    or g5385 ( n4150 , n29884 , n32558 );
    xnor g5386 ( n8838 , n3137 , n1599 );
    and g5387 ( n30200 , n18320 , n25624 );
    xnor g5388 ( n27550 , n7172 , n31215 );
    and g5389 ( n3806 , n27307 , n4265 );
    xnor g5390 ( n23770 , n20211 , n15403 );
    or g5391 ( n27964 , n4991 , n34039 );
    and g5392 ( n27473 , n17358 , n23224 );
    or g5393 ( n19980 , n35455 , n16797 );
    not g5394 ( n19257 , n19551 );
    and g5395 ( n11372 , n21546 , n33690 );
    and g5396 ( n2563 , n5907 , n30811 );
    buf g5397 ( n31514 , n25648 );
    and g5398 ( n9112 , n27132 , n3300 );
    and g5399 ( n11663 , n11988 , n26963 );
    or g5400 ( n29370 , n7460 , n407 );
    and g5401 ( n9183 , n17732 , n15323 );
    and g5402 ( n5941 , n22183 , n2740 );
    xnor g5403 ( n486 , n27122 , n25174 );
    or g5404 ( n18250 , n9793 , n10528 );
    or g5405 ( n28413 , n33959 , n23462 );
    not g5406 ( n19918 , n30316 );
    xnor g5407 ( n23431 , n1567 , n13976 );
    xnor g5408 ( n8443 , n3244 , n33722 );
    or g5409 ( n29706 , n3205 , n10099 );
    or g5410 ( n12909 , n36015 , n34016 );
    xnor g5411 ( n30728 , n10197 , n11967 );
    or g5412 ( n20819 , n16505 , n24289 );
    nor g5413 ( n31186 , n34698 , n33562 );
    and g5414 ( n20829 , n6914 , n12759 );
    or g5415 ( n17551 , n17642 , n2712 );
    or g5416 ( n32905 , n16049 , n21042 );
    and g5417 ( n12715 , n6179 , n3569 );
    or g5418 ( n6993 , n31559 , n12073 );
    or g5419 ( n20950 , n14910 , n30708 );
    or g5420 ( n588 , n360 , n3756 );
    and g5421 ( n31626 , n26278 , n21051 );
    xnor g5422 ( n28931 , n27258 , n32579 );
    xnor g5423 ( n18009 , n35505 , n4960 );
    xnor g5424 ( n9251 , n16573 , n4288 );
    xnor g5425 ( n20031 , n6751 , n4272 );
    and g5426 ( n35324 , n11366 , n16581 );
    and g5427 ( n9642 , n33002 , n7465 );
    and g5428 ( n18525 , n22109 , n22911 );
    and g5429 ( n4957 , n4665 , n9963 );
    and g5430 ( n3950 , n29455 , n20967 );
    or g5431 ( n10231 , n26748 , n4772 );
    and g5432 ( n25982 , n18764 , n4819 );
    xnor g5433 ( n29222 , n15432 , n26121 );
    or g5434 ( n8076 , n14743 , n23869 );
    xnor g5435 ( n9199 , n13837 , n20141 );
    or g5436 ( n23129 , n234 , n19649 );
    xnor g5437 ( n35882 , n20506 , n4758 );
    not g5438 ( n27969 , n27628 );
    or g5439 ( n14347 , n32781 , n12622 );
    xnor g5440 ( n14127 , n17854 , n17316 );
    and g5441 ( n31656 , n27333 , n33426 );
    not g5442 ( n26369 , n22471 );
    or g5443 ( n1703 , n11488 , n23626 );
    or g5444 ( n11962 , n27911 , n21977 );
    or g5445 ( n16993 , n23604 , n4013 );
    and g5446 ( n7945 , n13590 , n35378 );
    or g5447 ( n12688 , n17699 , n12950 );
    xnor g5448 ( n32509 , n27039 , n6151 );
    nor g5449 ( n19922 , n9789 , n7472 );
    not g5450 ( n3884 , n6596 );
    xnor g5451 ( n28289 , n30840 , n265 );
    or g5452 ( n31648 , n9706 , n2267 );
    xnor g5453 ( n15747 , n25013 , n25174 );
    or g5454 ( n27222 , n87 , n23921 );
    or g5455 ( n22580 , n11880 , n35623 );
    xnor g5456 ( n17564 , n7742 , n4960 );
    xnor g5457 ( n24898 , n28633 , n23604 );
    or g5458 ( n11262 , n32095 , n11248 );
    or g5459 ( n21356 , n19551 , n18838 );
    or g5460 ( n21498 , n11455 , n14006 );
    or g5461 ( n16873 , n12986 , n28455 );
    or g5462 ( n17011 , n23346 , n11833 );
    and g5463 ( n30490 , n18306 , n12939 );
    nor g5464 ( n32728 , n4878 , n17041 );
    xnor g5465 ( n8270 , n20416 , n4285 );
    nor g5466 ( n29486 , n26117 , n8004 );
    and g5467 ( n12205 , n21400 , n10614 );
    and g5468 ( n32020 , n24402 , n1777 );
    or g5469 ( n33841 , n17691 , n27782 );
    or g5470 ( n7135 , n3066 , n35422 );
    xnor g5471 ( n35175 , n28997 , n24371 );
    nor g5472 ( n8108 , n30854 , n542 );
    not g5473 ( n527 , n30586 );
    not g5474 ( n26800 , n27090 );
    not g5475 ( n18649 , n19939 );
    and g5476 ( n23001 , n1773 , n23949 );
    or g5477 ( n25112 , n26755 , n34219 );
    and g5478 ( n22641 , n33184 , n85 );
    or g5479 ( n35342 , n25174 , n33346 );
    and g5480 ( n28463 , n5504 , n21549 );
    or g5481 ( n34916 , n35150 , n21080 );
    and g5482 ( n35866 , n3827 , n23058 );
    or g5483 ( n11584 , n19542 , n16014 );
    or g5484 ( n12422 , n33148 , n29626 );
    not g5485 ( n13620 , n24834 );
    nor g5486 ( n1344 , n33524 , n29018 );
    or g5487 ( n2529 , n3543 , n4912 );
    or g5488 ( n28850 , n12015 , n6683 );
    and g5489 ( n26521 , n30872 , n4663 );
    and g5490 ( n24312 , n1147 , n6078 );
    or g5491 ( n34293 , n29421 , n35858 );
    and g5492 ( n17399 , n20112 , n24214 );
    and g5493 ( n208 , n11136 , n2567 );
    or g5494 ( n22510 , n7822 , n7961 );
    or g5495 ( n14463 , n25174 , n5166 );
    and g5496 ( n15079 , n11175 , n29016 );
    buf g5497 ( n2814 , n32194 );
    and g5498 ( n18676 , n5567 , n10890 );
    or g5499 ( n33852 , n30742 , n35404 );
    or g5500 ( n22606 , n18835 , n17730 );
    xnor g5501 ( n31364 , n1500 , n31559 );
    or g5502 ( n16712 , n15595 , n35630 );
    or g5503 ( n5264 , n19551 , n25041 );
    or g5504 ( n31723 , n33016 , n25896 );
    not g5505 ( n24502 , n26851 );
    or g5506 ( n23669 , n31109 , n11703 );
    and g5507 ( n957 , n13359 , n31289 );
    nor g5508 ( n14032 , n24362 , n13591 );
    and g5509 ( n2746 , n6298 , n6083 );
    xnor g5510 ( n21889 , n25931 , n14160 );
    or g5511 ( n33814 , n35927 , n8586 );
    and g5512 ( n31109 , n974 , n4471 );
    xnor g5513 ( n32066 , n20724 , n5323 );
    or g5514 ( n4731 , n32416 , n31134 );
    and g5515 ( n7564 , n34024 , n7384 );
    xnor g5516 ( n18405 , n20106 , n27866 );
    and g5517 ( n32878 , n15436 , n33623 );
    not g5518 ( n9016 , n2962 );
    xnor g5519 ( n15469 , n3178 , n32857 );
    or g5520 ( n12292 , n4592 , n3805 );
    and g5521 ( n16184 , n12134 , n21122 );
    nor g5522 ( n35754 , n32095 , n27833 );
    not g5523 ( n27511 , n16223 );
    xnor g5524 ( n18784 , n16552 , n18944 );
    xnor g5525 ( n7321 , n16881 , n3348 );
    or g5526 ( n4048 , n17641 , n28404 );
    or g5527 ( n34577 , n20697 , n2168 );
    xnor g5528 ( n19204 , n18158 , n17560 );
    xnor g5529 ( n1007 , n21397 , n17505 );
    and g5530 ( n1383 , n32661 , n17615 );
    or g5531 ( n8252 , n8994 , n19288 );
    or g5532 ( n14027 , n34800 , n13203 );
    and g5533 ( n30335 , n23180 , n22041 );
    or g5534 ( n28905 , n28416 , n29643 );
    and g5535 ( n30739 , n7798 , n10648 );
    or g5536 ( n19039 , n1156 , n2117 );
    or g5537 ( n19744 , n13332 , n27447 );
    and g5538 ( n34066 , n27389 , n30410 );
    nor g5539 ( n28111 , n31056 , n8298 );
    or g5540 ( n11117 , n4758 , n19450 );
    xnor g5541 ( n4803 , n16119 , n28295 );
    and g5542 ( n29760 , n20939 , n30845 );
    xnor g5543 ( n6182 , n4314 , n31799 );
    or g5544 ( n18330 , n6500 , n31006 );
    xnor g5545 ( n7108 , n28772 , n25513 );
    and g5546 ( n10301 , n12097 , n33835 );
    xnor g5547 ( n15419 , n3731 , n4059 );
    nor g5548 ( n881 , n30553 , n11810 );
    xnor g5549 ( n8661 , n23062 , n191 );
    xnor g5550 ( n10034 , n15747 , n13478 );
    or g5551 ( n3335 , n19280 , n35355 );
    or g5552 ( n35309 , n27568 , n26633 );
    and g5553 ( n11428 , n32773 , n11845 );
    and g5554 ( n31869 , n20661 , n5483 );
    xnor g5555 ( n32246 , n24852 , n5343 );
    xnor g5556 ( n34538 , n3720 , n20669 );
    xnor g5557 ( n20485 , n25016 , n5517 );
    and g5558 ( n5178 , n8989 , n29192 );
    xnor g5559 ( n20383 , n6156 , n31065 );
    xnor g5560 ( n12173 , n2909 , n5428 );
    or g5561 ( n10426 , n27892 , n33658 );
    xnor g5562 ( n19841 , n214 , n29839 );
    and g5563 ( n24930 , n14050 , n9158 );
    xnor g5564 ( n12611 , n17095 , n15623 );
    and g5565 ( n32734 , n3614 , n16656 );
    or g5566 ( n24423 , n27066 , n17962 );
    or g5567 ( n5498 , n31911 , n33157 );
    and g5568 ( n4915 , n11016 , n14796 );
    or g5569 ( n34017 , n22029 , n23715 );
    not g5570 ( n3523 , n6236 );
    or g5571 ( n20968 , n20875 , n33656 );
    or g5572 ( n4138 , n24164 , n23792 );
    or g5573 ( n7689 , n23269 , n26931 );
    and g5574 ( n5118 , n21878 , n10116 );
    not g5575 ( n32851 , n8432 );
    or g5576 ( n10308 , n24371 , n1652 );
    or g5577 ( n3965 , n34691 , n13015 );
    not g5578 ( n402 , n20316 );
    or g5579 ( n3010 , n20090 , n22858 );
    or g5580 ( n20274 , n11046 , n25301 );
    or g5581 ( n27155 , n35927 , n15509 );
    or g5582 ( n12847 , n9658 , n12093 );
    not g5583 ( n28299 , n6793 );
    or g5584 ( n16745 , n2784 , n5779 );
    not g5585 ( n3863 , n558 );
    or g5586 ( n20359 , n33326 , n16457 );
    or g5587 ( n5369 , n30655 , n19571 );
    or g5588 ( n24219 , n335 , n5752 );
    and g5589 ( n22312 , n29678 , n26983 );
    or g5590 ( n14624 , n19458 , n5424 );
    xnor g5591 ( n15208 , n14354 , n13976 );
    xnor g5592 ( n19172 , n32452 , n25602 );
    or g5593 ( n13415 , n13798 , n2611 );
    and g5594 ( n30695 , n11503 , n13124 );
    nor g5595 ( n23606 , n22366 , n32379 );
    or g5596 ( n7980 , n5584 , n19767 );
    or g5597 ( n3672 , n7853 , n28675 );
    and g5598 ( n34673 , n19981 , n33671 );
    or g5599 ( n12717 , n12972 , n7903 );
    or g5600 ( n35178 , n13789 , n23655 );
    or g5601 ( n15551 , n6780 , n949 );
    xnor g5602 ( n18699 , n27538 , n5598 );
    or g5603 ( n30344 , n3960 , n4545 );
    or g5604 ( n9304 , n11557 , n27973 );
    or g5605 ( n8732 , n27567 , n27973 );
    xnor g5606 ( n20554 , n30345 , n34635 );
    nor g5607 ( n34314 , n22291 , n26267 );
    nor g5608 ( n12052 , n23915 , n23921 );
    or g5609 ( n10365 , n18982 , n24479 );
    or g5610 ( n27595 , n5335 , n34098 );
    or g5611 ( n5962 , n9658 , n34096 );
    and g5612 ( n640 , n31975 , n3418 );
    and g5613 ( n24829 , n2377 , n514 );
    or g5614 ( n17268 , n30251 , n34084 );
    or g5615 ( n25077 , n27386 , n28036 );
    or g5616 ( n11007 , n18791 , n5900 );
    xnor g5617 ( n2143 , n19995 , n9909 );
    xnor g5618 ( n18408 , n8579 , n4016 );
    and g5619 ( n15921 , n3748 , n32884 );
    xnor g5620 ( n26259 , n25351 , n24267 );
    or g5621 ( n26334 , n17568 , n20872 );
    xnor g5622 ( n9187 , n9538 , n16922 );
    and g5623 ( n1968 , n19704 , n7004 );
    and g5624 ( n17434 , n31615 , n14768 );
    nor g5625 ( n19993 , n350 , n7653 );
    xnor g5626 ( n2248 , n10454 , n33025 );
    or g5627 ( n6640 , n5876 , n34229 );
    or g5628 ( n1622 , n4484 , n31055 );
    xnor g5629 ( n31438 , n12319 , n15886 );
    or g5630 ( n26996 , n31289 , n21679 );
    or g5631 ( n34963 , n19931 , n28060 );
    or g5632 ( n2869 , n35927 , n11048 );
    and g5633 ( n33417 , n10541 , n13179 );
    or g5634 ( n22740 , n17474 , n24336 );
    or g5635 ( n9762 , n5608 , n13307 );
    xnor g5636 ( n337 , n16715 , n9658 );
    or g5637 ( n26444 , n5654 , n16553 );
    and g5638 ( n25372 , n2229 , n30728 );
    or g5639 ( n24870 , n28265 , n5771 );
    nor g5640 ( n1535 , n20696 , n21251 );
    not g5641 ( n26958 , n28699 );
    xnor g5642 ( n2644 , n11684 , n32715 );
    or g5643 ( n18452 , n7540 , n5226 );
    xnor g5644 ( n27540 , n12991 , n830 );
    xnor g5645 ( n30209 , n10845 , n21220 );
    and g5646 ( n11308 , n19296 , n2071 );
    and g5647 ( n4316 , n11196 , n25979 );
    or g5648 ( n18821 , n5235 , n20300 );
    and g5649 ( n7998 , n4256 , n14663 );
    and g5650 ( n10745 , n2403 , n20476 );
    not g5651 ( n7892 , n20427 );
    or g5652 ( n31901 , n20995 , n83 );
    or g5653 ( n23810 , n4878 , n2986 );
    xnor g5654 ( n29480 , n16475 , n19633 );
    and g5655 ( n29787 , n28095 , n10454 );
    xnor g5656 ( n19924 , n9623 , n4288 );
    and g5657 ( n17869 , n3031 , n20745 );
    or g5658 ( n12369 , n34080 , n31464 );
    and g5659 ( n12197 , n23716 , n26991 );
    or g5660 ( n5328 , n941 , n15144 );
    nor g5661 ( n4307 , n17568 , n33114 );
    or g5662 ( n19662 , n26441 , n908 );
    and g5663 ( n25066 , n16850 , n15133 );
    nor g5664 ( n17281 , n6111 , n21673 );
    xnor g5665 ( n11780 , n29031 , n27760 );
    or g5666 ( n21046 , n9793 , n9265 );
    not g5667 ( n19594 , n8066 );
    or g5668 ( n23862 , n32095 , n11001 );
    xnor g5669 ( n29297 , n18700 , n28012 );
    or g5670 ( n8162 , n2624 , n16797 );
    or g5671 ( n16808 , n11455 , n29919 );
    and g5672 ( n18181 , n625 , n25840 );
    and g5673 ( n5368 , n22125 , n1971 );
    or g5674 ( n1258 , n3291 , n25786 );
    xnor g5675 ( n36043 , n26253 , n32851 );
    or g5676 ( n24079 , n1950 , n14464 );
    and g5677 ( n21486 , n22903 , n34056 );
    and g5678 ( n33284 , n2681 , n19266 );
    or g5679 ( n32177 , n16922 , n19949 );
    or g5680 ( n5574 , n23877 , n3756 );
    or g5681 ( n4601 , n7005 , n10400 );
    not g5682 ( n20037 , n14585 );
    nor g5683 ( n1863 , n32857 , n27783 );
    or g5684 ( n33080 , n32314 , n29872 );
    or g5685 ( n5728 , n19001 , n11712 );
    and g5686 ( n30146 , n27110 , n26788 );
    or g5687 ( n24201 , n18354 , n31071 );
    or g5688 ( n34984 , n24681 , n21210 );
    and g5689 ( n26834 , n35901 , n11201 );
    and g5690 ( n14938 , n33191 , n33849 );
    xnor g5691 ( n29546 , n31461 , n16922 );
    and g5692 ( n1222 , n33282 , n31122 );
    or g5693 ( n29331 , n25137 , n9034 );
    xnor g5694 ( n17273 , n15376 , n10894 );
    xnor g5695 ( n9939 , n23026 , n7055 );
    or g5696 ( n29727 , n13283 , n35762 );
    xnor g5697 ( n4255 , n9962 , n12724 );
    or g5698 ( n3457 , n16228 , n31554 );
    xnor g5699 ( n34770 , n9401 , n29990 );
    or g5700 ( n15385 , n15528 , n28324 );
    xnor g5701 ( n3259 , n17285 , n12437 );
    or g5702 ( n21624 , n1240 , n31589 );
    or g5703 ( n5983 , n4758 , n6124 );
    and g5704 ( n29754 , n2059 , n24155 );
    or g5705 ( n34407 , n29839 , n6817 );
    and g5706 ( n15056 , n8862 , n20796 );
    or g5707 ( n12978 , n28720 , n4772 );
    or g5708 ( n11725 , n33460 , n20762 );
    and g5709 ( n31633 , n20000 , n14422 );
    or g5710 ( n13392 , n19465 , n16305 );
    or g5711 ( n19377 , n18680 , n25500 );
    xnor g5712 ( n10571 , n30212 , n17301 );
    xnor g5713 ( n8931 , n5286 , n32857 );
    or g5714 ( n16472 , n9793 , n31467 );
    xnor g5715 ( n21991 , n24689 , n16480 );
    and g5716 ( n31232 , n35083 , n1984 );
    or g5717 ( n28054 , n28520 , n1142 );
    or g5718 ( n8200 , n4972 , n13664 );
    or g5719 ( n9606 , n32095 , n4749 );
    and g5720 ( n19391 , n1985 , n11199 );
    and g5721 ( n11390 , n16093 , n10883 );
    or g5722 ( n17291 , n900 , n19058 );
    xnor g5723 ( n21610 , n17701 , n29713 );
    xnor g5724 ( n13298 , n32360 , n8949 );
    and g5725 ( n79 , n24031 , n9468 );
    xnor g5726 ( n22586 , n23269 , n31287 );
    nor g5727 ( n6085 , n318 , n32329 );
    xnor g5728 ( n12542 , n14665 , n33251 );
    and g5729 ( n23399 , n16269 , n14417 );
    or g5730 ( n29339 , n3599 , n22886 );
    or g5731 ( n35705 , n1950 , n11010 );
    not g5732 ( n12367 , n8353 );
    not g5733 ( n22281 , n30742 );
    or g5734 ( n24846 , n1863 , n19909 );
    xnor g5735 ( n1885 , n10228 , n12951 );
    and g5736 ( n16145 , n10588 , n1037 );
    xnor g5737 ( n9824 , n21142 , n25889 );
    xnor g5738 ( n8551 , n31762 , n32095 );
    not g5739 ( n34939 , n35775 );
    and g5740 ( n34667 , n25143 , n16070 );
    nor g5741 ( n817 , n1248 , n6017 );
    or g5742 ( n10020 , n11337 , n30519 );
    xnor g5743 ( n22283 , n20955 , n34707 );
    xnor g5744 ( n7011 , n32604 , n20836 );
    xnor g5745 ( n4247 , n27868 , n3205 );
    nor g5746 ( n4732 , n30306 , n18913 );
    not g5747 ( n3344 , n22501 );
    xnor g5748 ( n11114 , n11139 , n33894 );
    nor g5749 ( n20944 , n10894 , n33887 );
    and g5750 ( n20301 , n19514 , n31199 );
    and g5751 ( n11029 , n14348 , n16686 );
    and g5752 ( n15319 , n35664 , n14463 );
    xnor g5753 ( n21114 , n2429 , n11455 );
    xnor g5754 ( n23781 , n1749 , n32570 );
    xnor g5755 ( n6848 , n27102 , n25602 );
    not g5756 ( n24695 , n19551 );
    or g5757 ( n9857 , n8432 , n16953 );
    not g5758 ( n7125 , n3222 );
    not g5759 ( n22926 , n16620 );
    xnor g5760 ( n17896 , n8317 , n1950 );
    and g5761 ( n14126 , n35770 , n6263 );
    and g5762 ( n12897 , n3691 , n18973 );
    xnor g5763 ( n11557 , n34706 , n5800 );
    or g5764 ( n2003 , n9614 , n19166 );
    and g5765 ( n27164 , n24914 , n19199 );
    or g5766 ( n28362 , n8263 , n27143 );
    and g5767 ( n27085 , n21905 , n7491 );
    or g5768 ( n35528 , n22488 , n12596 );
    or g5769 ( n13815 , n23404 , n7340 );
    or g5770 ( n12379 , n4758 , n27943 );
    xnor g5771 ( n1495 , n9218 , n29624 );
    not g5772 ( n36049 , n10894 );
    and g5773 ( n34117 , n26340 , n30380 );
    xnor g5774 ( n11964 , n26390 , n31559 );
    or g5775 ( n3612 , n14780 , n17162 );
    or g5776 ( n33909 , n19425 , n13015 );
    xnor g5777 ( n17114 , n17755 , n31559 );
    nor g5778 ( n33740 , n16620 , n2451 );
    nor g5779 ( n1372 , n15695 , n19432 );
    and g5780 ( n22572 , n3435 , n10633 );
    or g5781 ( n18975 , n14693 , n34609 );
    or g5782 ( n7042 , n22218 , n21681 );
    nor g5783 ( n11433 , n31799 , n23068 );
    nor g5784 ( n25424 , n14848 , n25867 );
    xnor g5785 ( n7963 , n7713 , n2090 );
    or g5786 ( n32202 , n32847 , n23567 );
    or g5787 ( n33495 , n12836 , n16464 );
    not g5788 ( n4788 , n18121 );
    not g5789 ( n35306 , n8366 );
    or g5790 ( n5069 , n4204 , n20762 );
    or g5791 ( n33828 , n7144 , n15497 );
    and g5792 ( n3349 , n14032 , n12154 );
    or g5793 ( n485 , n12251 , n16019 );
    and g5794 ( n4970 , n10781 , n7996 );
    and g5795 ( n27276 , n28994 , n15848 );
    not g5796 ( n21478 , n7912 );
    not g5797 ( n30140 , n32857 );
    or g5798 ( n33305 , n31297 , n22010 );
    xnor g5799 ( n10589 , n9980 , n8008 );
    xnor g5800 ( n28731 , n4955 , n13096 );
    or g5801 ( n25738 , n32080 , n22858 );
    or g5802 ( n18256 , n29583 , n34404 );
    xor g5803 ( n23960 , n6218 , n16911 );
    or g5804 ( n6248 , n23963 , n33578 );
    not g5805 ( n23887 , n11931 );
    and g5806 ( n255 , n9716 , n15314 );
    and g5807 ( n16749 , n31491 , n34083 );
    xnor g5808 ( n32137 , n1900 , n4962 );
    or g5809 ( n24392 , n28390 , n22081 );
    or g5810 ( n18587 , n30506 , n3979 );
    or g5811 ( n12980 , n34599 , n27625 );
    or g5812 ( n30789 , n34002 , n2524 );
    or g5813 ( n985 , n4288 , n33604 );
    xnor g5814 ( n5908 , n7901 , n9789 );
    xnor g5815 ( n34632 , n32055 , n21328 );
    or g5816 ( n9495 , n13093 , n24937 );
    or g5817 ( n1912 , n12498 , n3858 );
    and g5818 ( n20181 , n278 , n1325 );
    and g5819 ( n18527 , n5432 , n33876 );
    and g5820 ( n26146 , n952 , n29085 );
    xnor g5821 ( n8930 , n27125 , n32584 );
    not g5822 ( n17161 , n1091 );
    nor g5823 ( n29813 , n4607 , n20127 );
    nor g5824 ( n14670 , n527 , n18807 );
    not g5825 ( n27564 , n368 );
    and g5826 ( n35292 , n11689 , n11723 );
    not g5827 ( n27402 , n23604 );
    or g5828 ( n14543 , n2644 , n8288 );
    or g5829 ( n33029 , n33060 , n22858 );
    xnor g5830 ( n27896 , n15609 , n3205 );
    or g5831 ( n6428 , n26379 , n26220 );
    or g5832 ( n12439 , n13548 , n27625 );
    or g5833 ( n31613 , n10303 , n6568 );
    or g5834 ( n30101 , n4878 , n4898 );
    xnor g5835 ( n16004 , n9380 , n16922 );
    or g5836 ( n21589 , n3068 , n16456 );
    and g5837 ( n1768 , n9252 , n16054 );
    and g5838 ( n19812 , n26902 , n20520 );
    xnor g5839 ( n27133 , n4991 , n34039 );
    or g5840 ( n26104 , n792 , n16006 );
    and g5841 ( n24520 , n30058 , n16383 );
    xnor g5842 ( n10293 , n35088 , n27225 );
    and g5843 ( n32693 , n2520 , n19358 );
    or g5844 ( n26145 , n31438 , n14077 );
    and g5845 ( n31302 , n5211 , n14123 );
    or g5846 ( n21390 , n11134 , n1846 );
    xnor g5847 ( n4726 , n17517 , n26885 );
    or g5848 ( n32651 , n12135 , n11703 );
    nor g5849 ( n8772 , n19998 , n27501 );
    xnor g5850 ( n16810 , n12696 , n15003 );
    nor g5851 ( n10804 , n35856 , n2494 );
    xnor g5852 ( n24050 , n18756 , n35258 );
    xnor g5853 ( n15673 , n35680 , n4868 );
    or g5854 ( n6602 , n29661 , n34537 );
    or g5855 ( n33097 , n33639 , n5230 );
    or g5856 ( n6001 , n33044 , n13912 );
    or g5857 ( n23745 , n3093 , n15290 );
    and g5858 ( n23677 , n31251 , n34535 );
    nor g5859 ( n28420 , n32407 , n18115 );
    or g5860 ( n7307 , n8418 , n21673 );
    or g5861 ( n26065 , n19738 , n14295 );
    nor g5862 ( n21208 , n10454 , n23495 );
    buf g5863 ( n6683 , n34923 );
    xnor g5864 ( n31106 , n4157 , n4878 );
    or g5865 ( n20020 , n11455 , n3093 );
    or g5866 ( n3996 , n30953 , n2524 );
    xnor g5867 ( n27761 , n9467 , n9789 );
    or g5868 ( n13899 , n9789 , n7901 );
    or g5869 ( n9769 , n18149 , n25914 );
    and g5870 ( n8103 , n14771 , n19801 );
    or g5871 ( n20609 , n31298 , n21579 );
    xnor g5872 ( n20666 , n16016 , n31289 );
    or g5873 ( n13811 , n34203 , n24356 );
    nor g5874 ( n35400 , n34567 , n6017 );
    or g5875 ( n18129 , n32857 , n14662 );
    nor g5876 ( n21961 , n12637 , n9921 );
    xnor g5877 ( n4913 , n14883 , n4878 );
    or g5878 ( n20876 , n24371 , n19216 );
    and g5879 ( n2523 , n4799 , n28294 );
    nor g5880 ( n28579 , n11455 , n25015 );
    and g5881 ( n20541 , n32344 , n23084 );
    and g5882 ( n21701 , n32099 , n18773 );
    or g5883 ( n12134 , n36048 , n19487 );
    and g5884 ( n31099 , n2715 , n4385 );
    xnor g5885 ( n13381 , n18636 , n30397 );
    or g5886 ( n6079 , n11171 , n20589 );
    or g5887 ( n15994 , n10562 , n19213 );
    and g5888 ( n21890 , n22454 , n11102 );
    not g5889 ( n33530 , n32857 );
    not g5890 ( n35472 , n7699 );
    or g5891 ( n26881 , n4077 , n23921 );
    or g5892 ( n14240 , n30502 , n8139 );
    or g5893 ( n34875 , n7704 , n13924 );
    xnor g5894 ( n605 , n242 , n2085 );
    and g5895 ( n14148 , n7007 , n10875 );
    xnor g5896 ( n11546 , n24552 , n32584 );
    xnor g5897 ( n23618 , n747 , n35709 );
    or g5898 ( n32078 , n7350 , n34865 );
    nor g5899 ( n12011 , n25602 , n35521 );
    or g5900 ( n11748 , n20981 , n15518 );
    or g5901 ( n32865 , n29807 , n19391 );
    or g5902 ( n26414 , n16620 , n13142 );
    or g5903 ( n13183 , n19482 , n33157 );
    or g5904 ( n31688 , n10378 , n22967 );
    xnor g5905 ( n18876 , n32568 , n10982 );
    or g5906 ( n23167 , n21924 , n6779 );
    and g5907 ( n3308 , n4070 , n1242 );
    xnor g5908 ( n16030 , n16242 , n4878 );
    or g5909 ( n24301 , n24810 , n22316 );
    nor g5910 ( n8399 , n23766 , n33287 );
    xnor g5911 ( n7498 , n1819 , n7240 );
    and g5912 ( n3357 , n28387 , n25101 );
    or g5913 ( n30662 , n34840 , n27694 );
    or g5914 ( n9624 , n242 , n19058 );
    or g5915 ( n19784 , n28915 , n2798 );
    xnor g5916 ( n20198 , n30798 , n30742 );
    or g5917 ( n2120 , n11623 , n26689 );
    or g5918 ( n11207 , n59 , n9030 );
    and g5919 ( n35005 , n35061 , n28542 );
    nor g5920 ( n29805 , n26449 , n18115 );
    and g5921 ( n28554 , n23596 , n22731 );
    or g5922 ( n9159 , n3009 , n1511 );
    and g5923 ( n6684 , n35184 , n29524 );
    and g5924 ( n24643 , n14996 , n1270 );
    xnor g5925 ( n7951 , n31750 , n29871 );
    or g5926 ( n16309 , n4878 , n26256 );
    or g5927 ( n26399 , n764 , n27232 );
    not g5928 ( n19708 , n10894 );
    or g5929 ( n30564 , n14561 , n31134 );
    or g5930 ( n2025 , n35136 , n31549 );
    or g5931 ( n17344 , n10322 , n1322 );
    or g5932 ( n4143 , n8466 , n14055 );
    or g5933 ( n18188 , n33291 , n31484 );
    xnor g5934 ( n17228 , n29271 , n22736 );
    or g5935 ( n4643 , n1339 , n10872 );
    xnor g5936 ( n20106 , n6741 , n24371 );
    and g5937 ( n32964 , n18373 , n14177 );
    xnor g5938 ( n30108 , n7282 , n1225 );
    or g5939 ( n31979 , n1295 , n35935 );
    or g5940 ( n4384 , n10948 , n30179 );
    xnor g5941 ( n35008 , n32832 , n14994 );
    and g5942 ( n9550 , n3509 , n20034 );
    or g5943 ( n36089 , n23991 , n13931 );
    not g5944 ( n16698 , n2029 );
    xnor g5945 ( n34960 , n1694 , n35295 );
    or g5946 ( n3152 , n20738 , n3026 );
    nor g5947 ( n12225 , n16620 , n28947 );
    nor g5948 ( n23715 , n25926 , n16548 );
    or g5949 ( n7524 , n2863 , n34865 );
    or g5950 ( n6639 , n12678 , n19767 );
    or g5951 ( n31263 , n29911 , n1511 );
    xnor g5952 ( n6123 , n15234 , n29713 );
    and g5953 ( n19736 , n12976 , n3775 );
    or g5954 ( n2006 , n25420 , n15102 );
    and g5955 ( n28365 , n29691 , n31064 );
    or g5956 ( n28762 , n14231 , n30461 );
    not g5957 ( n5290 , n8547 );
    xnor g5958 ( n8183 , n23483 , n24839 );
    or g5959 ( n24912 , n27179 , n34484 );
    or g5960 ( n17059 , n12877 , n22682 );
    and g5961 ( n26910 , n21326 , n4107 );
    or g5962 ( n24146 , n10208 , n8090 );
    xnor g5963 ( n3384 , n6189 , n11849 );
    or g5964 ( n336 , n31284 , n949 );
    or g5965 ( n35471 , n9556 , n31606 );
    or g5966 ( n20430 , n1706 , n15742 );
    or g5967 ( n30609 , n16113 , n22501 );
    or g5968 ( n10782 , n34329 , n12326 );
    or g5969 ( n5294 , n13845 , n20579 );
    or g5970 ( n1056 , n20242 , n32268 );
    not g5971 ( n13096 , n24371 );
    xnor g5972 ( n1883 , n27212 , n32095 );
    or g5973 ( n17719 , n17195 , n35630 );
    or g5974 ( n32696 , n17568 , n20155 );
    not g5975 ( n35943 , n25135 );
    or g5976 ( n3404 , n18552 , n26264 );
    or g5977 ( n14546 , n1364 , n14681 );
    not g5978 ( n10133 , n22873 );
    and g5979 ( n18195 , n7638 , n15833 );
    and g5980 ( n1480 , n26171 , n21879 );
    or g5981 ( n27930 , n9693 , n20812 );
    or g5982 ( n8261 , n23604 , n25847 );
    and g5983 ( n15037 , n28056 , n10190 );
    and g5984 ( n2705 , n33595 , n7696 );
    or g5985 ( n2507 , n16174 , n16345 );
    or g5986 ( n35077 , n5098 , n31464 );
    not g5987 ( n32484 , n18296 );
    and g5988 ( n6205 , n35844 , n5814 );
    not g5989 ( n955 , n7713 );
    or g5990 ( n3408 , n3846 , n15791 );
    or g5991 ( n26639 , n31559 , n22942 );
    xnor g5992 ( n34611 , n15380 , n31712 );
    or g5993 ( n13844 , n30670 , n6683 );
    or g5994 ( n8690 , n17375 , n19153 );
    xnor g5995 ( n11382 , n19824 , n30804 );
    or g5996 ( n24992 , n21930 , n2798 );
    xnor g5997 ( n31969 , n28733 , n16801 );
    and g5998 ( n23773 , n6614 , n24182 );
    or g5999 ( n3734 , n4962 , n21026 );
    or g6000 ( n8751 , n18622 , n13307 );
    not g6001 ( n8461 , n27627 );
    nor g6002 ( n6543 , n29874 , n15145 );
    or g6003 ( n28535 , n11455 , n13689 );
    and g6004 ( n21488 , n20006 , n7186 );
    or g6005 ( n25578 , n10298 , n9773 );
    or g6006 ( n32790 , n15403 , n19810 );
    and g6007 ( n13161 , n7641 , n12177 );
    or g6008 ( n1137 , n35307 , n30646 );
    and g6009 ( n22834 , n14974 , n20663 );
    or g6010 ( n10797 , n15403 , n14578 );
    xnor g6011 ( n1220 , n3570 , n16922 );
    xnor g6012 ( n33348 , n18742 , n15896 );
    nor g6013 ( n35629 , n11835 , n28605 );
    or g6014 ( n32163 , n17835 , n35402 );
    xnor g6015 ( n20171 , n3041 , n5067 );
    xnor g6016 ( n34913 , n24460 , n2454 );
    or g6017 ( n8272 , n26643 , n12578 );
    nor g6018 ( n3290 , n31289 , n5765 );
    xnor g6019 ( n13181 , n4693 , n20401 );
    xnor g6020 ( n30422 , n10252 , n28088 );
    or g6021 ( n18003 , n10856 , n13397 );
    nor g6022 ( n31303 , n4962 , n30865 );
    or g6023 ( n19207 , n20031 , n14746 );
    and g6024 ( n21521 , n34153 , n35632 );
    and g6025 ( n35518 , n29303 , n25921 );
    xnor g6026 ( n11064 , n17086 , n32866 );
    or g6027 ( n13588 , n30320 , n32505 );
    or g6028 ( n35014 , n35505 , n17233 );
    or g6029 ( n18662 , n34213 , n27769 );
    or g6030 ( n34598 , n21021 , n6981 );
    xnor g6031 ( n35162 , n34259 , n18363 );
    nor g6032 ( n19688 , n35927 , n18158 );
    xnor g6033 ( n7336 , n30425 , n4288 );
    xnor g6034 ( n28690 , n27379 , n26752 );
    or g6035 ( n5525 , n9658 , n28139 );
    not g6036 ( n8495 , n9658 );
    or g6037 ( n19885 , n29839 , n933 );
    or g6038 ( n20169 , n34949 , n20189 );
    or g6039 ( n24668 , n17398 , n4363 );
    nor g6040 ( n9327 , n32584 , n33765 );
    or g6041 ( n26107 , n9676 , n16919 );
    or g6042 ( n20538 , n849 , n949 );
    or g6043 ( n69 , n6315 , n4478 );
    and g6044 ( n5045 , n11795 , n1562 );
    and g6045 ( n5150 , n21501 , n26592 );
    and g6046 ( n23757 , n13959 , n12241 );
    xnor g6047 ( n14222 , n14873 , n19317 );
    or g6048 ( n13251 , n31839 , n12658 );
    and g6049 ( n613 , n17167 , n18094 );
    and g6050 ( n19 , n32440 , n26530 );
    or g6051 ( n5551 , n10281 , n17337 );
    xnor g6052 ( n1626 , n28043 , n20486 );
    or g6053 ( n9602 , n24942 , n9983 );
    or g6054 ( n14033 , n8966 , n27728 );
    nor g6055 ( n14256 , n9793 , n19752 );
    not g6056 ( n2817 , n3239 );
    or g6057 ( n9572 , n35716 , n25773 );
    or g6058 ( n1285 , n5335 , n21998 );
    xnor g6059 ( n34195 , n30276 , n33440 );
    or g6060 ( n17255 , n9658 , n27722 );
    and g6061 ( n20727 , n28452 , n2427 );
    or g6062 ( n7517 , n8945 , n19952 );
    or g6063 ( n14604 , n13911 , n32572 );
    or g6064 ( n4190 , n19822 , n7553 );
    and g6065 ( n25366 , n30915 , n16967 );
    and g6066 ( n18694 , n25628 , n29834 );
    xnor g6067 ( n21067 , n27783 , n6791 );
    and g6068 ( n32298 , n21024 , n33603 );
    or g6069 ( n4031 , n24134 , n13390 );
    not g6070 ( n22870 , n25648 );
    xnor g6071 ( n33838 , n20768 , n31289 );
    and g6072 ( n20853 , n19625 , n32319 );
    or g6073 ( n28461 , n32860 , n8905 );
    or g6074 ( n32942 , n21116 , n13145 );
    xnor g6075 ( n13135 , n20937 , n9793 );
    or g6076 ( n2196 , n19871 , n30826 );
    or g6077 ( n12795 , n4878 , n11621 );
    not g6078 ( n8027 , n12822 );
    nor g6079 ( n23076 , n35927 , n1297 );
    nor g6080 ( n9256 , n3222 , n29418 );
    xnor g6081 ( n33735 , n3707 , n15299 );
    xnor g6082 ( n7021 , n34178 , n30558 );
    or g6083 ( n33638 , n9543 , n16457 );
    not g6084 ( n28864 , n11807 );
    xnor g6085 ( n17274 , n25633 , n31919 );
    or g6086 ( n3359 , n8154 , n26486 );
    xnor g6087 ( n14646 , n8182 , n27912 );
    and g6088 ( n18427 , n28824 , n27586 );
    not g6089 ( n13396 , n19602 );
    or g6090 ( n21848 , n632 , n12563 );
    xnor g6091 ( n15017 , n2462 , n22291 );
    and g6092 ( n15378 , n12609 , n23467 );
    or g6093 ( n24083 , n14734 , n7584 );
    xnor g6094 ( n19900 , n18677 , n29445 );
    xnor g6095 ( n32976 , n18781 , n29372 );
    or g6096 ( n13774 , n26286 , n3552 );
    or g6097 ( n4961 , n4288 , n4915 );
    xnor g6098 ( n35684 , n29831 , n25778 );
    or g6099 ( n32151 , n9944 , n25447 );
    not g6100 ( n31050 , n14532 );
    or g6101 ( n25388 , n25174 , n4186 );
    and g6102 ( n27778 , n13986 , n5135 );
    or g6103 ( n28660 , n16941 , n31850 );
    or g6104 ( n24601 , n22538 , n35757 );
    or g6105 ( n14488 , n13920 , n8878 );
    and g6106 ( n3052 , n898 , n22432 );
    or g6107 ( n34843 , n18781 , n29372 );
    buf g6108 ( n8865 , n13343 );
    or g6109 ( n29199 , n16257 , n34378 );
    nor g6110 ( n9679 , n6534 , n26672 );
    and g6111 ( n6591 , n35450 , n30376 );
    or g6112 ( n25050 , n23853 , n25761 );
    or g6113 ( n21468 , n15431 , n27075 );
    xnor g6114 ( n11652 , n12300 , n5929 );
    or g6115 ( n28526 , n4267 , n35209 );
    xnor g6116 ( n18867 , n15163 , n9789 );
    xnor g6117 ( n33255 , n31180 , n9789 );
    or g6118 ( n12960 , n19888 , n30826 );
    and g6119 ( n14464 , n24871 , n12788 );
    and g6120 ( n32297 , n34949 , n12460 );
    xnor g6121 ( n22077 , n18271 , n16620 );
    xnor g6122 ( n8706 , n12133 , n19551 );
    buf g6123 ( n7588 , n18441 );
    xnor g6124 ( n2915 , n30987 , n4962 );
    or g6125 ( n1310 , n35383 , n33435 );
    xnor g6126 ( n27713 , n15157 , n1950 );
    or g6127 ( n5904 , n24972 , n19732 );
    or g6128 ( n1290 , n31056 , n681 );
    and g6129 ( n11786 , n26478 , n3885 );
    xnor g6130 ( n2635 , n5695 , n29713 );
    and g6131 ( n28631 , n10327 , n24067 );
    or g6132 ( n35531 , n21196 , n30826 );
    xnor g6133 ( n20899 , n2952 , n15281 );
    or g6134 ( n2856 , n24633 , n6553 );
    xnor g6135 ( n10401 , n23959 , n10894 );
    or g6136 ( n11746 , n6730 , n10417 );
    nor g6137 ( n31611 , n21068 , n10335 );
    or g6138 ( n25393 , n12164 , n17354 );
    and g6139 ( n19213 , n22898 , n7502 );
    or g6140 ( n28424 , n6316 , n13305 );
    or g6141 ( n33202 , n26649 , n5440 );
    and g6142 ( n12482 , n35222 , n23468 );
    and g6143 ( n29488 , n29503 , n25308 );
    and g6144 ( n32997 , n31646 , n25188 );
    xnor g6145 ( n26154 , n19064 , n8324 );
    xnor g6146 ( n15597 , n33621 , n7540 );
    or g6147 ( n15312 , n19551 , n17713 );
    or g6148 ( n2220 , n13601 , n10432 );
    or g6149 ( n5485 , n10375 , n3345 );
    not g6150 ( n26448 , n19984 );
    xnor g6151 ( n16336 , n18114 , n21441 );
    or g6152 ( n15370 , n16062 , n24551 );
    or g6153 ( n22164 , n27280 , n23323 );
    and g6154 ( n10999 , n12784 , n21908 );
    and g6155 ( n26312 , n7979 , n33532 );
    xnor g6156 ( n23754 , n1565 , n31289 );
    or g6157 ( n3001 , n1950 , n5263 );
    and g6158 ( n3420 , n13780 , n35448 );
    xnor g6159 ( n20764 , n12661 , n23327 );
    xnor g6160 ( n12735 , n32143 , n29713 );
    and g6161 ( n36019 , n9211 , n25467 );
    and g6162 ( n35822 , n27576 , n11768 );
    or g6163 ( n28970 , n2952 , n15281 );
    and g6164 ( n35540 , n2160 , n6925 );
    or g6165 ( n9909 , n12311 , n16059 );
    not g6166 ( n3148 , n16620 );
    or g6167 ( n32698 , n29895 , n5779 );
    and g6168 ( n22096 , n28277 , n2178 );
    and g6169 ( n12456 , n24049 , n15427 );
    or g6170 ( n8114 , n34517 , n31643 );
    or g6171 ( n34483 , n35853 , n15025 );
    and g6172 ( n20251 , n14829 , n31604 );
    nor g6173 ( n11661 , n19551 , n3543 );
    xnor g6174 ( n8554 , n3202 , n32135 );
    and g6175 ( n23492 , n11778 , n27149 );
    not g6176 ( n16728 , n12326 );
    xnor g6177 ( n9039 , n27283 , n6665 );
    xnor g6178 ( n29648 , n9038 , n3950 );
    xnor g6179 ( n6472 , n16025 , n33605 );
    nor g6180 ( n31961 , n19551 , n6685 );
    or g6181 ( n17145 , n13372 , n7422 );
    or g6182 ( n27068 , n19145 , n29854 );
    xnor g6183 ( n25238 , n4901 , n9789 );
    or g6184 ( n16201 , n9273 , n22858 );
    not g6185 ( n4132 , n17108 );
    and g6186 ( n12188 , n8339 , n7985 );
    and g6187 ( n11128 , n2677 , n18077 );
    or g6188 ( n4006 , n3138 , n25306 );
    and g6189 ( n22663 , n21070 , n19680 );
    or g6190 ( n24787 , n5190 , n15538 );
    or g6191 ( n10618 , n9658 , n35042 );
    not g6192 ( n15548 , n9789 );
    or g6193 ( n28715 , n4960 , n21089 );
    or g6194 ( n13406 , n5958 , n2798 );
    xnor g6195 ( n6173 , n3584 , n6720 );
    xnor g6196 ( n8544 , n29364 , n6088 );
    nor g6197 ( n606 , n27328 , n19834 );
    or g6198 ( n2682 , n14079 , n2119 );
    not g6199 ( n533 , n15886 );
    and g6200 ( n25710 , n19737 , n32165 );
    xnor g6201 ( n9614 , n12490 , n29713 );
    buf g6202 ( n16464 , n20749 );
    and g6203 ( n20902 , n29335 , n21662 );
    not g6204 ( n31268 , n10351 );
    or g6205 ( n27162 , n4513 , n10142 );
    nor g6206 ( n29980 , n391 , n24505 );
    not g6207 ( n13362 , n19076 );
    nor g6208 ( n2820 , n11125 , n28993 );
    or g6209 ( n21934 , n29994 , n24333 );
    xnor g6210 ( n31098 , n33985 , n1013 );
    or g6211 ( n7103 , n20937 , n13015 );
    or g6212 ( n7631 , n3693 , n10379 );
    or g6213 ( n26283 , n6658 , n20681 );
    or g6214 ( n29371 , n17580 , n26480 );
    or g6215 ( n15118 , n14138 , n26112 );
    xnor g6216 ( n25329 , n12413 , n30141 );
    xnor g6217 ( n31000 , n2443 , n22376 );
    xnor g6218 ( n27819 , n18641 , n32339 );
    xnor g6219 ( n12424 , n14081 , n18598 );
    and g6220 ( n26865 , n3266 , n31352 );
    and g6221 ( n22102 , n16714 , n6957 );
    buf g6222 ( n1942 , n11184 );
    and g6223 ( n35784 , n19062 , n20989 );
    xnor g6224 ( n12877 , n4926 , n384 );
    xnor g6225 ( n9738 , n17756 , n11046 );
    buf g6226 ( n11518 , n34643 );
    nor g6227 ( n2364 , n24371 , n32336 );
    or g6228 ( n29002 , n29881 , n24333 );
    or g6229 ( n19399 , n18491 , n25652 );
    nor g6230 ( n475 , n24853 , n16803 );
    or g6231 ( n36060 , n4962 , n27596 );
    or g6232 ( n31640 , n14704 , n32608 );
    and g6233 ( n22080 , n18928 , n33423 );
    buf g6234 ( n15497 , n21624 );
    or g6235 ( n10436 , n28165 , n8203 );
    not g6236 ( n33933 , n29203 );
    or g6237 ( n11658 , n12775 , n12996 );
    and g6238 ( n22456 , n20384 , n22249 );
    and g6239 ( n14844 , n13549 , n9914 );
    and g6240 ( n17246 , n35270 , n11923 );
    xnor g6241 ( n2453 , n31089 , n5197 );
    and g6242 ( n20830 , n32966 , n31151 );
    or g6243 ( n21605 , n8334 , n33558 );
    not g6244 ( n26513 , n5067 );
    or g6245 ( n13930 , n8817 , n32634 );
    or g6246 ( n34628 , n4030 , n27574 );
    or g6247 ( n15817 , n14485 , n1557 );
    or g6248 ( n19768 , n4761 , n22934 );
    nor g6249 ( n17515 , n27436 , n3292 );
    buf g6250 ( n19952 , n15573 );
    or g6251 ( n9750 , n11813 , n12913 );
    xnor g6252 ( n30042 , n9140 , n4962 );
    and g6253 ( n2841 , n9231 , n17323 );
    not g6254 ( n26199 , n28811 );
    nor g6255 ( n6717 , n15464 , n7115 );
    or g6256 ( n21655 , n33941 , n19403 );
    or g6257 ( n29658 , n8206 , n22997 );
    or g6258 ( n35361 , n16936 , n7578 );
    not g6259 ( n32395 , n9793 );
    xnor g6260 ( n14609 , n10833 , n4554 );
    and g6261 ( n21322 , n26520 , n1333 );
    and g6262 ( n17475 , n5498 , n35160 );
    nor g6263 ( n10760 , n34054 , n12088 );
    xnor g6264 ( n2447 , n34938 , n24371 );
    xnor g6265 ( n26137 , n18581 , n31968 );
    or g6266 ( n14519 , n31449 , n35422 );
    not g6267 ( n32658 , n4878 );
    xnor g6268 ( n32660 , n31506 , n9254 );
    and g6269 ( n17722 , n29925 , n22601 );
    or g6270 ( n1871 , n29900 , n29411 );
    xnor g6271 ( n27504 , n28142 , n21782 );
    or g6272 ( n12593 , n33220 , n22858 );
    and g6273 ( n15585 , n6032 , n32402 );
    not g6274 ( n12228 , n3222 );
    not g6275 ( n14167 , n20287 );
    xnor g6276 ( n7769 , n11166 , n946 );
    xnor g6277 ( n18469 , n26207 , n35445 );
    and g6278 ( n9104 , n22266 , n744 );
    xnor g6279 ( n2822 , n19028 , n31056 );
    nor g6280 ( n26847 , n31799 , n15531 );
    or g6281 ( n5125 , n22057 , n5008 );
    and g6282 ( n30117 , n5439 , n15867 );
    not g6283 ( n15704 , n32857 );
    or g6284 ( n34115 , n12624 , n31198 );
    and g6285 ( n33725 , n33972 , n34791 );
    and g6286 ( n19038 , n22729 , n30781 );
    not g6287 ( n33353 , n4962 );
    nor g6288 ( n5953 , n22421 , n9921 );
    not g6289 ( n2528 , n23788 );
    or g6290 ( n5308 , n19988 , n29917 );
    and g6291 ( n12840 , n29074 , n7804 );
    not g6292 ( n33925 , n22980 );
    or g6293 ( n8213 , n10456 , n20690 );
    or g6294 ( n7850 , n9789 , n22637 );
    not g6295 ( n1793 , n32572 );
    xor g6296 ( n30404 , n6880 , n19551 );
    or g6297 ( n27439 , n30512 , n15496 );
    or g6298 ( n26076 , n20907 , n20576 );
    or g6299 ( n10342 , n18832 , n31134 );
    xnor g6300 ( n28616 , n31956 , n19999 );
    or g6301 ( n5006 , n28026 , n31626 );
    or g6302 ( n15130 , n30175 , n10336 );
    not g6303 ( n14411 , n25602 );
    nor g6304 ( n19252 , n4960 , n17603 );
    xnor g6305 ( n25534 , n18886 , n13035 );
    or g6306 ( n35634 , n22861 , n12474 );
    xnor g6307 ( n14401 , n11623 , n26689 );
    xnor g6308 ( n35823 , n27095 , n18097 );
    xnor g6309 ( n20615 , n23455 , n11455 );
    nor g6310 ( n2601 , n5287 , n16536 );
    xnor g6311 ( n19995 , n31966 , n2056 );
    or g6312 ( n22705 , n35950 , n25897 );
    or g6313 ( n22756 , n3786 , n8152 );
    or g6314 ( n15379 , n23190 , n23790 );
    and g6315 ( n8486 , n5938 , n28524 );
    and g6316 ( n26360 , n10390 , n23146 );
    and g6317 ( n16107 , n30310 , n22407 );
    not g6318 ( n2698 , n3858 );
    and g6319 ( n26955 , n26947 , n729 );
    and g6320 ( n16716 , n1711 , n1398 );
    nor g6321 ( n9034 , n20525 , n22077 );
    or g6322 ( n426 , n11699 , n256 );
    or g6323 ( n24182 , n27291 , n2222 );
    or g6324 ( n642 , n21810 , n31001 );
    xnor g6325 ( n28055 , n24945 , n29537 );
    nor g6326 ( n10394 , n8696 , n8657 );
    and g6327 ( n33447 , n11627 , n11036 );
    xnor g6328 ( n11306 , n14991 , n9165 );
    or g6329 ( n25408 , n10988 , n9443 );
    or g6330 ( n34712 , n28752 , n28939 );
    xnor g6331 ( n5901 , n2254 , n16620 );
    xnor g6332 ( n12018 , n33454 , n4962 );
    and g6333 ( n1317 , n24523 , n32635 );
    or g6334 ( n9559 , n10016 , n12612 );
    xnor g6335 ( n1349 , n2148 , n15886 );
    or g6336 ( n19068 , n28133 , n11741 );
    not g6337 ( n31854 , n32608 );
    xnor g6338 ( n10462 , n13505 , n5260 );
    or g6339 ( n34114 , n18039 , n51 );
    not g6340 ( n35340 , n7950 );
    or g6341 ( n19644 , n35882 , n32351 );
    or g6342 ( n23818 , n34073 , n32608 );
    not g6343 ( n31608 , n10184 );
    and g6344 ( n19311 , n30814 , n34461 );
    or g6345 ( n6843 , n29458 , n11518 );
    or g6346 ( n4537 , n10542 , n27952 );
    or g6347 ( n23273 , n16922 , n19277 );
    not g6348 ( n30911 , n19182 );
    xnor g6349 ( n24387 , n17794 , n8855 );
    or g6350 ( n10330 , n9789 , n20393 );
    or g6351 ( n19627 , n29520 , n28740 );
    and g6352 ( n23030 , n6496 , n25640 );
    xnor g6353 ( n17083 , n32825 , n32857 );
    or g6354 ( n17113 , n34511 , n25411 );
    xnor g6355 ( n20729 , n8975 , n25402 );
    and g6356 ( n23319 , n34107 , n21444 );
    or g6357 ( n10713 , n14354 , n5168 );
    nor g6358 ( n3343 , n15464 , n16582 );
    and g6359 ( n26321 , n12738 , n7390 );
    xnor g6360 ( n2893 , n34649 , n31559 );
    or g6361 ( n20763 , n11928 , n5900 );
    or g6362 ( n1854 , n30097 , n11977 );
    or g6363 ( n18108 , n1950 , n24950 );
    xnor g6364 ( n2758 , n4749 , n32095 );
    or g6365 ( n16951 , n12396 , n32321 );
    or g6366 ( n22875 , n10252 , n28088 );
    not g6367 ( n26701 , n7523 );
    or g6368 ( n13030 , n33245 , n25567 );
    or g6369 ( n10831 , n8742 , n15756 );
    or g6370 ( n10190 , n22638 , n28248 );
    or g6371 ( n21487 , n30951 , n13646 );
    and g6372 ( n8026 , n1822 , n35032 );
    xnor g6373 ( n24531 , n2899 , n35230 );
    or g6374 ( n23220 , n33891 , n26002 );
    or g6375 ( n10124 , n30553 , n35879 );
    or g6376 ( n9143 , n28151 , n29899 );
    or g6377 ( n15400 , n18096 , n21042 );
    or g6378 ( n5674 , n3350 , n14924 );
    or g6379 ( n7020 , n19810 , n24653 );
    buf g6380 ( n25786 , n33368 );
    or g6381 ( n29041 , n1015 , n9488 );
    buf g6382 ( n14746 , n32434 );
    not g6383 ( n23678 , n25839 );
    buf g6384 ( n17111 , n22761 );
    xnor g6385 ( n27496 , n350 , n34792 );
    xnor g6386 ( n25542 , n35753 , n35696 );
    nor g6387 ( n25205 , n4960 , n13770 );
    and g6388 ( n16389 , n35527 , n22830 );
    or g6389 ( n23023 , n11901 , n20318 );
    buf g6390 ( n4952 , n15871 );
    or g6391 ( n8850 , n20566 , n9672 );
    or g6392 ( n4349 , n3773 , n10872 );
    not g6393 ( n27428 , n16475 );
    xnor g6394 ( n10325 , n16591 , n29565 );
    and g6395 ( n5707 , n24135 , n34550 );
    and g6396 ( n13213 , n2015 , n31223 );
    nor g6397 ( n1196 , n9689 , n1218 );
    or g6398 ( n26558 , n20215 , n6950 );
    and g6399 ( n23069 , n16982 , n2493 );
    or g6400 ( n20509 , n10894 , n17208 );
    or g6401 ( n12784 , n18827 , n15145 );
    xnor g6402 ( n12140 , n17423 , n10915 );
    xnor g6403 ( n20962 , n2635 , n8663 );
    or g6404 ( n20745 , n13520 , n27053 );
    or g6405 ( n15181 , n24371 , n5894 );
    and g6406 ( n31582 , n5518 , n13665 );
    and g6407 ( n26239 , n20283 , n30693 );
    and g6408 ( n9926 , n16544 , n6357 );
    or g6409 ( n27316 , n9820 , n26737 );
    xnor g6410 ( n23134 , n15558 , n22746 );
    or g6411 ( n25433 , n31195 , n15012 );
    and g6412 ( n35801 , n28427 , n2165 );
    and g6413 ( n17565 , n29654 , n11762 );
    xnor g6414 ( n32064 , n3429 , n13059 );
    or g6415 ( n5838 , n18379 , n2539 );
    or g6416 ( n20409 , n25314 , n35721 );
    not g6417 ( n26366 , n34620 );
    or g6418 ( n33427 , n29733 , n4956 );
    xnor g6419 ( n22797 , n35150 , n3940 );
    or g6420 ( n10956 , n21497 , n2104 );
    and g6421 ( n24331 , n1029 , n5573 );
    or g6422 ( n28777 , n15316 , n25567 );
    xnor g6423 ( n27683 , n890 , n12272 );
    xnor g6424 ( n7188 , n25717 , n4878 );
    nor g6425 ( n17389 , n3205 , n3291 );
    and g6426 ( n35187 , n27440 , n8643 );
    and g6427 ( n34361 , n32702 , n13367 );
    or g6428 ( n30392 , n9490 , n22105 );
    and g6429 ( n13010 , n25955 , n1927 );
    and g6430 ( n7118 , n29606 , n4660 );
    not g6431 ( n8364 , n30292 );
    or g6432 ( n35885 , n10393 , n6749 );
    or g6433 ( n13369 , n35727 , n2524 );
    or g6434 ( n509 , n12603 , n19496 );
    or g6435 ( n17310 , n27432 , n28591 );
    not g6436 ( n16125 , n4960 );
    or g6437 ( n23364 , n2622 , n24489 );
    xnor g6438 ( n1510 , n32518 , n5287 );
    or g6439 ( n18732 , n33415 , n25648 );
    or g6440 ( n9843 , n33047 , n3756 );
    not g6441 ( n26486 , n6288 );
    and g6442 ( n7169 , n31785 , n15312 );
    and g6443 ( n2122 , n12891 , n11339 );
    or g6444 ( n31162 , n15779 , n25592 );
    xnor g6445 ( n1082 , n10568 , n30553 );
    or g6446 ( n33297 , n8432 , n25814 );
    or g6447 ( n184 , n18875 , n27453 );
    or g6448 ( n24658 , n16705 , n16797 );
    and g6449 ( n1097 , n34282 , n21574 );
    and g6450 ( n35786 , n12386 , n12981 );
    xnor g6451 ( n9687 , n21533 , n4960 );
    and g6452 ( n16086 , n13938 , n20534 );
    and g6453 ( n28295 , n2365 , n17456 );
    xnor g6454 ( n17602 , n35666 , n30742 );
    and g6455 ( n14648 , n21310 , n4313 );
    xnor g6456 ( n21748 , n5584 , n4962 );
    xnor g6457 ( n31157 , n7144 , n35113 );
    or g6458 ( n23021 , n19309 , n23462 );
    and g6459 ( n20448 , n28800 , n10270 );
    or g6460 ( n15408 , n5287 , n9435 );
    and g6461 ( n120 , n17913 , n27466 );
    and g6462 ( n32618 , n26511 , n28259 );
    xnor g6463 ( n4381 , n31531 , n35151 );
    nor g6464 ( n2125 , n597 , n20689 );
    or g6465 ( n6237 , n21668 , n25019 );
    not g6466 ( n21315 , n10946 );
    or g6467 ( n35147 , n25013 , n1715 );
    or g6468 ( n15589 , n17749 , n12128 );
    xnor g6469 ( n17910 , n16827 , n16285 );
    nor g6470 ( n14877 , n35958 , n33933 );
    and g6471 ( n35355 , n20097 , n16877 );
    and g6472 ( n30809 , n23679 , n15557 );
    or g6473 ( n31719 , n30742 , n4044 );
    and g6474 ( n27813 , n18302 , n29474 );
    not g6475 ( n31641 , n6890 );
    not g6476 ( n5060 , n23910 );
    xnor g6477 ( n7057 , n18000 , n18521 );
    or g6478 ( n23463 , n7119 , n4175 );
    and g6479 ( n12955 , n33315 , n323 );
    or g6480 ( n21331 , n24687 , n15109 );
    or g6481 ( n12889 , n5067 , n19830 );
    or g6482 ( n21807 , n24007 , n15625 );
    and g6483 ( n19820 , n28029 , n23145 );
    xnor g6484 ( n32040 , n5677 , n3205 );
    or g6485 ( n33820 , n57 , n1832 );
    or g6486 ( n14234 , n525 , n3634 );
    not g6487 ( n21735 , n11455 );
    xnor g6488 ( n22260 , n31439 , n33931 );
    xnor g6489 ( n29903 , n32972 , n29839 );
    and g6490 ( n27370 , n34925 , n2290 );
    or g6491 ( n26809 , n26619 , n3680 );
    and g6492 ( n7861 , n30211 , n12870 );
    nor g6493 ( n5692 , n29238 , n6424 );
    xnor g6494 ( n6822 , n8658 , n4430 );
    or g6495 ( n9043 , n7157 , n27756 );
    or g6496 ( n26984 , n35177 , n33730 );
    and g6497 ( n27218 , n5269 , n18461 );
    or g6498 ( n12139 , n637 , n19105 );
    xnor g6499 ( n34480 , n32230 , n16943 );
    or g6500 ( n6019 , n17753 , n26352 );
    and g6501 ( n14140 , n13997 , n3487 );
    xnor g6502 ( n17361 , n33487 , n3968 );
    not g6503 ( n25524 , n10894 );
    or g6504 ( n34720 , n20477 , n19338 );
    or g6505 ( n12121 , n18232 , n32572 );
    or g6506 ( n21431 , n19551 , n22202 );
    or g6507 ( n31965 , n26875 , n31134 );
    or g6508 ( n21821 , n4962 , n22713 );
    or g6509 ( n29584 , n24798 , n7167 );
    or g6510 ( n32149 , n20294 , n4508 );
    or g6511 ( n12050 , n3865 , n24696 );
    and g6512 ( n32671 , n19691 , n28168 );
    or g6513 ( n23207 , n24520 , n4912 );
    and g6514 ( n14747 , n17674 , n11599 );
    xnor g6515 ( n17529 , n2770 , n3946 );
    xnor g6516 ( n9474 , n27135 , n26103 );
    and g6517 ( n1730 , n16787 , n7117 );
    not g6518 ( n20997 , n30948 );
    and g6519 ( n29666 , n16507 , n15374 );
    or g6520 ( n5377 , n16397 , n19659 );
    or g6521 ( n33153 , n29713 , n8238 );
    and g6522 ( n18300 , n6129 , n68 );
    and g6523 ( n17126 , n23166 , n16375 );
    and g6524 ( n27426 , n26445 , n30029 );
    or g6525 ( n4750 , n21186 , n16133 );
    xnor g6526 ( n3183 , n17578 , n28696 );
    or g6527 ( n31355 , n35372 , n22548 );
    or g6528 ( n8226 , n20962 , n35630 );
    nor g6529 ( n10816 , n31289 , n7029 );
    and g6530 ( n5412 , n13552 , n2007 );
    xnor g6531 ( n19323 , n27925 , n7540 );
    or g6532 ( n20831 , n15116 , n11850 );
    and g6533 ( n11085 , n23844 , n2020 );
    or g6534 ( n6407 , n3205 , n24161 );
    or g6535 ( n33600 , n17075 , n9194 );
    not g6536 ( n559 , n35422 );
    and g6537 ( n22700 , n34629 , n8502 );
    or g6538 ( n28448 , n5282 , n3188 );
    or g6539 ( n11936 , n31264 , n6210 );
    not g6540 ( n26190 , n3614 );
    or g6541 ( n9743 , n13734 , n6259 );
    or g6542 ( n22630 , n11014 , n15497 );
    nor g6543 ( n1582 , n35994 , n33287 );
    xnor g6544 ( n32545 , n12748 , n20360 );
    or g6545 ( n10216 , n27445 , n7337 );
    and g6546 ( n15022 , n30912 , n3155 );
    xnor g6547 ( n32858 , n20504 , n25602 );
    or g6548 ( n16369 , n6508 , n12913 );
    or g6549 ( n12492 , n32378 , n15781 );
    not g6550 ( n35224 , n11294 );
    or g6551 ( n22683 , n8819 , n31718 );
    nor g6552 ( n27528 , n4962 , n25088 );
    and g6553 ( n30975 , n33552 , n34964 );
    and g6554 ( n15599 , n15177 , n2862 );
    xnor g6555 ( n31682 , n13718 , n31477 );
    or g6556 ( n15492 , n7035 , n11996 );
    or g6557 ( n33123 , n32731 , n35179 );
    or g6558 ( n11886 , n26830 , n28438 );
    xnor g6559 ( n4400 , n20794 , n8674 );
    or g6560 ( n29450 , n22327 , n12622 );
    and g6561 ( n17257 , n5185 , n32024 );
    or g6562 ( n22093 , n31215 , n25435 );
    not g6563 ( n1824 , n33435 );
    or g6564 ( n1065 , n3946 , n22222 );
    or g6565 ( n31380 , n7876 , n16543 );
    or g6566 ( n5997 , n12696 , n21313 );
    xnor g6567 ( n26408 , n11188 , n7540 );
    or g6568 ( n6154 , n14656 , n4014 );
    and g6569 ( n27596 , n13219 , n7687 );
    or g6570 ( n1509 , n23855 , n10762 );
    xnor g6571 ( n29094 , n14166 , n30037 );
    nor g6572 ( n22458 , n18655 , n30595 );
    or g6573 ( n18522 , n31212 , n8888 );
    or g6574 ( n10738 , n5604 , n8292 );
    and g6575 ( n11041 , n28829 , n34628 );
    or g6576 ( n20778 , n113 , n2745 );
    xnor g6577 ( n35071 , n31913 , n25135 );
    and g6578 ( n16775 , n18485 , n30430 );
    and g6579 ( n33812 , n33175 , n24219 );
    and g6580 ( n23602 , n32787 , n17014 );
    and g6581 ( n29508 , n1053 , n13410 );
    nor g6582 ( n2905 , n25602 , n31400 );
    xnor g6583 ( n223 , n16113 , n31215 );
    or g6584 ( n13888 , n4756 , n19734 );
    and g6585 ( n913 , n13972 , n15411 );
    not g6586 ( n30381 , n31411 );
    and g6587 ( n1076 , n24297 , n28147 );
    nor g6588 ( n3841 , n17568 , n11522 );
    or g6589 ( n7520 , n14654 , n22316 );
    and g6590 ( n19135 , n10865 , n20886 );
    or g6591 ( n2245 , n31802 , n29383 );
    or g6592 ( n24133 , n31478 , n29909 );
    or g6593 ( n12592 , n31976 , n1069 );
    or g6594 ( n16846 , n22409 , n1934 );
    or g6595 ( n2833 , n31781 , n29592 );
    and g6596 ( n9295 , n23383 , n15773 );
    xnor g6597 ( n15693 , n8140 , n17409 );
    xnor g6598 ( n21225 , n12656 , n25488 );
    or g6599 ( n23656 , n129 , n21771 );
    and g6600 ( n4662 , n1954 , n5845 );
    or g6601 ( n4156 , n25002 , n21691 );
    nor g6602 ( n30679 , n18293 , n24505 );
    nor g6603 ( n30541 , n31382 , n34360 );
    xnor g6604 ( n33734 , n12647 , n36040 );
    nor g6605 ( n7398 , n32857 , n10450 );
    xnor g6606 ( n26614 , n12911 , n33007 );
    or g6607 ( n10359 , n17923 , n27218 );
    nor g6608 ( n3624 , n31799 , n16244 );
    or g6609 ( n26506 , n5700 , n6288 );
    xnor g6610 ( n27448 , n25478 , n15464 );
    or g6611 ( n7039 , n19856 , n19939 );
    or g6612 ( n8106 , n7546 , n35935 );
    nor g6613 ( n16290 , n1950 , n11148 );
    not g6614 ( n889 , n30742 );
    and g6615 ( n27907 , n34417 , n9243 );
    or g6616 ( n28134 , n27474 , n1586 );
    and g6617 ( n10027 , n26767 , n20845 );
    not g6618 ( n11594 , n6919 );
    xnor g6619 ( n26637 , n7998 , n35927 );
    not g6620 ( n18233 , n4960 );
    or g6621 ( n35477 , n10411 , n30431 );
    or g6622 ( n989 , n18597 , n1682 );
    and g6623 ( n5397 , n25759 , n19533 );
    or g6624 ( n18391 , n13153 , n4952 );
    or g6625 ( n18727 , n6817 , n1176 );
    buf g6626 ( n12622 , n6037 );
    xnor g6627 ( n25923 , n1736 , n17568 );
    xnor g6628 ( n18463 , n27292 , n773 );
    and g6629 ( n35420 , n22385 , n19969 );
    or g6630 ( n5817 , n1389 , n28404 );
    not g6631 ( n3380 , n15539 );
    xnor g6632 ( n719 , n21116 , n13145 );
    or g6633 ( n31545 , n4077 , n7671 );
    or g6634 ( n33771 , n1638 , n585 );
    nor g6635 ( n33693 , n15403 , n14617 );
    and g6636 ( n29278 , n29112 , n33575 );
    and g6637 ( n17041 , n11272 , n26992 );
    or g6638 ( n26012 , n10957 , n28248 );
    or g6639 ( n17741 , n4634 , n23544 );
    or g6640 ( n6590 , n32545 , n21210 );
    or g6641 ( n35040 , n33610 , n33707 );
    or g6642 ( n11412 , n20405 , n2918 );
    not g6643 ( n23717 , n12622 );
    or g6644 ( n32439 , n13702 , n15538 );
    or g6645 ( n5362 , n24818 , n1345 );
    and g6646 ( n33897 , n25202 , n7715 );
    or g6647 ( n1530 , n26597 , n16919 );
    and g6648 ( n212 , n15893 , n2109 );
    nor g6649 ( n25570 , n9568 , n3671 );
    and g6650 ( n24959 , n31263 , n20315 );
    or g6651 ( n29073 , n14765 , n8366 );
    not g6652 ( n32148 , n17480 );
    and g6653 ( n5064 , n8522 , n22267 );
    xnor g6654 ( n11870 , n615 , n32095 );
    and g6655 ( n7745 , n13725 , n29613 );
    or g6656 ( n21745 , n3867 , n26480 );
    or g6657 ( n3297 , n5039 , n6181 );
    or g6658 ( n28084 , n30720 , n32071 );
    or g6659 ( n35248 , n17175 , n24294 );
    not g6660 ( n21587 , n32857 );
    or g6661 ( n24471 , n29531 , n2104 );
    or g6662 ( n27847 , n8813 , n9951 );
    or g6663 ( n20641 , n29995 , n17233 );
    or g6664 ( n6179 , n11597 , n23043 );
    or g6665 ( n4633 , n18374 , n27574 );
    or g6666 ( n32409 , n3584 , n10336 );
    or g6667 ( n21938 , n26900 , n945 );
    and g6668 ( n25999 , n5415 , n32544 );
    or g6669 ( n14133 , n2795 , n34801 );
    or g6670 ( n22232 , n29839 , n21269 );
    or g6671 ( n15461 , n34296 , n34084 );
    or g6672 ( n12066 , n15235 , n2384 );
    xnor g6673 ( n5585 , n19294 , n31271 );
    and g6674 ( n4629 , n1146 , n22433 );
    xnor g6675 ( n712 , n13296 , n13257 );
    and g6676 ( n6094 , n24977 , n1471 );
    xnor g6677 ( n33601 , n8356 , n18248 );
    xnor g6678 ( n24606 , n4863 , n24868 );
    or g6679 ( n18688 , n19717 , n32808 );
    nor g6680 ( n3341 , n13281 , n25390 );
    xnor g6681 ( n30228 , n12218 , n5335 );
    or g6682 ( n31846 , n1439 , n10952 );
    or g6683 ( n29086 , n7577 , n19084 );
    and g6684 ( n34558 , n29120 , n12696 );
    or g6685 ( n19081 , n29983 , n24356 );
    or g6686 ( n34129 , n10894 , n15959 );
    and g6687 ( n4213 , n8013 , n6547 );
    not g6688 ( n33142 , n17475 );
    and g6689 ( n20175 , n3213 , n24618 );
    xnor g6690 ( n25382 , n21108 , n24371 );
    xnor g6691 ( n16954 , n12830 , n35927 );
    xnor g6692 ( n35980 , n14489 , n24332 );
    or g6693 ( n20287 , n35033 , n30992 );
    xnor g6694 ( n11882 , n10102 , n17695 );
    and g6695 ( n14354 , n6337 , n3564 );
    and g6696 ( n3906 , n32609 , n21580 );
    nor g6697 ( n13920 , n21846 , n31411 );
    and g6698 ( n3917 , n24379 , n17001 );
    xnor g6699 ( n119 , n7985 , n8339 );
    or g6700 ( n30263 , n18107 , n1796 );
    or g6701 ( n7798 , n29361 , n10432 );
    xnor g6702 ( n246 , n27036 , n25459 );
    xnor g6703 ( n32037 , n1632 , n24582 );
    xnor g6704 ( n30603 , n20226 , n35216 );
    xnor g6705 ( n8038 , n24760 , n29713 );
    or g6706 ( n31779 , n14851 , n19952 );
    not g6707 ( n21186 , n20249 );
    or g6708 ( n30891 , n28051 , n25625 );
    nor g6709 ( n22647 , n31382 , n30770 );
    and g6710 ( n20664 , n24678 , n33930 );
    nor g6711 ( n20312 , n31289 , n13359 );
    and g6712 ( n32624 , n28694 , n9713 );
    or g6713 ( n9514 , n2883 , n31514 );
    and g6714 ( n24566 , n7747 , n28563 );
    or g6715 ( n20782 , n33880 , n20762 );
    xnor g6716 ( n22119 , n34502 , n17751 );
    xnor g6717 ( n23516 , n13812 , n19575 );
    nor g6718 ( n7164 , n31799 , n3812 );
    or g6719 ( n23385 , n20417 , n28198 );
    or g6720 ( n30258 , n14025 , n30292 );
    not g6721 ( n23689 , n17939 );
    or g6722 ( n1976 , n24371 , n18343 );
    or g6723 ( n14562 , n4908 , n6825 );
    and g6724 ( n18287 , n25158 , n19144 );
    and g6725 ( n2506 , n22184 , n30437 );
    and g6726 ( n33185 , n27668 , n35110 );
    nor g6727 ( n20628 , n31610 , n2629 );
    xnor g6728 ( n26326 , n8418 , n281 );
    or g6729 ( n2009 , n11046 , n16314 );
    and g6730 ( n13326 , n17639 , n32181 );
    or g6731 ( n20809 , n32392 , n25940 );
    and g6732 ( n12334 , n801 , n24809 );
    not g6733 ( n117 , n4878 );
    nor g6734 ( n21882 , n11190 , n18353 );
    and g6735 ( n25123 , n23782 , n24077 );
    or g6736 ( n30174 , n22799 , n10634 );
    or g6737 ( n24577 , n177 , n31337 );
    or g6738 ( n31235 , n31038 , n9731 );
    xnor g6739 ( n25838 , n14063 , n13170 );
    xnor g6740 ( n23699 , n35183 , n11279 );
    and g6741 ( n20789 , n574 , n8093 );
    or g6742 ( n15666 , n22681 , n14963 );
    and g6743 ( n20090 , n24146 , n26889 );
    nor g6744 ( n20115 , n29839 , n19925 );
    buf g6745 ( n11712 , n11770 );
    and g6746 ( n19206 , n3701 , n27492 );
    or g6747 ( n15562 , n25699 , n30646 );
    or g6748 ( n26684 , n10623 , n28574 );
    not g6749 ( n28544 , n17939 );
    xnor g6750 ( n10362 , n11606 , n35078 );
    or g6751 ( n34949 , n33856 , n1014 );
    xnor g6752 ( n33226 , n23737 , n4288 );
    xnor g6753 ( n32936 , n20132 , n22992 );
    or g6754 ( n7058 , n27482 , n1372 );
    not g6755 ( n19285 , n32324 );
    or g6756 ( n19396 , n29083 , n33310 );
    or g6757 ( n9185 , n30742 , n16230 );
    or g6758 ( n9714 , n124 , n12958 );
    nor g6759 ( n20568 , n11455 , n23221 );
    or g6760 ( n22184 , n19444 , n11977 );
    nor g6761 ( n17608 , n30742 , n32569 );
    or g6762 ( n3544 , n22549 , n139 );
    and g6763 ( n3387 , n28346 , n24418 );
    or g6764 ( n33032 , n10293 , n8203 );
    xnor g6765 ( n16061 , n24624 , n9789 );
    not g6766 ( n29855 , n16620 );
    and g6767 ( n11993 , n303 , n34060 );
    or g6768 ( n2882 , n32715 , n27485 );
    and g6769 ( n31638 , n7837 , n20656 );
    not g6770 ( n20358 , n20427 );
    and g6771 ( n19475 , n10205 , n34037 );
    or g6772 ( n8393 , n6093 , n26747 );
    and g6773 ( n33430 , n16170 , n31628 );
    or g6774 ( n5642 , n12947 , n5168 );
    or g6775 ( n1275 , n8779 , n8399 );
    nor g6776 ( n9648 , n33037 , n35720 );
    or g6777 ( n887 , n15886 , n12319 );
    or g6778 ( n22848 , n24807 , n12791 );
    or g6779 ( n13103 , n23675 , n31514 );
    and g6780 ( n10383 , n16355 , n11443 );
    xnor g6781 ( n22134 , n31109 , n22291 );
    and g6782 ( n19827 , n21541 , n8883 );
    nor g6783 ( n35559 , n8911 , n23921 );
    or g6784 ( n21482 , n15299 , n19736 );
    or g6785 ( n17428 , n9502 , n139 );
    not g6786 ( n538 , n25300 );
    or g6787 ( n24514 , n8695 , n16153 );
    xnor g6788 ( n27038 , n18208 , n29839 );
    and g6789 ( n32943 , n32927 , n29605 );
    or g6790 ( n19920 , n983 , n1942 );
    and g6791 ( n3532 , n15352 , n19298 );
    or g6792 ( n20156 , n18492 , n35422 );
    and g6793 ( n1948 , n15441 , n2301 );
    and g6794 ( n7220 , n21141 , n18153 );
    or g6795 ( n8050 , n16987 , n19584 );
    not g6796 ( n11473 , n14427 );
    or g6797 ( n14891 , n7540 , n17390 );
    or g6798 ( n30882 , n4611 , n32505 );
    and g6799 ( n33320 , n25470 , n30352 );
    or g6800 ( n3086 , n2051 , n19125 );
    or g6801 ( n26983 , n19551 , n28996 );
    and g6802 ( n24856 , n26417 , n27835 );
    xnor g6803 ( n4154 , n4147 , n24928 );
    nor g6804 ( n28439 , n25602 , n1383 );
    and g6805 ( n1306 , n35864 , n13069 );
    or g6806 ( n34485 , n6412 , n11258 );
    xnor g6807 ( n25122 , n8129 , n35290 );
    or g6808 ( n4372 , n33962 , n28811 );
    xnor g6809 ( n2942 , n5172 , n24129 );
    or g6810 ( n11388 , n5040 , n17204 );
    and g6811 ( n35555 , n25733 , n26913 );
    not g6812 ( n19942 , n22241 );
    and g6813 ( n7758 , n31778 , n15104 );
    and g6814 ( n14545 , n16131 , n27403 );
    not g6815 ( n7787 , n4354 );
    or g6816 ( n23994 , n6572 , n26659 );
    or g6817 ( n14894 , n11455 , n28865 );
    or g6818 ( n13787 , n8417 , n20922 );
    or g6819 ( n28764 , n10185 , n15519 );
    nor g6820 ( n24038 , n8683 , n29203 );
    and g6821 ( n4436 , n30341 , n22889 );
    and g6822 ( n23611 , n12717 , n28049 );
    or g6823 ( n804 , n19551 , n23459 );
    and g6824 ( n2770 , n30371 , n31614 );
    xnor g6825 ( n33334 , n28798 , n9793 );
    or g6826 ( n20117 , n3205 , n13632 );
    xnor g6827 ( n29837 , n30105 , n10911 );
    and g6828 ( n5403 , n9470 , n25754 );
    xnor g6829 ( n35308 , n19590 , n23027 );
    and g6830 ( n4826 , n1772 , n19240 );
    and g6831 ( n32518 , n32998 , n6356 );
    xnor g6832 ( n33501 , n21865 , n34598 );
    xnor g6833 ( n25544 , n27461 , n19433 );
    xnor g6834 ( n6310 , n27503 , n28330 );
    xnor g6835 ( n1086 , n3394 , n6987 );
    or g6836 ( n9004 , n5287 , n24589 );
    or g6837 ( n7833 , n23394 , n14076 );
    or g6838 ( n15711 , n31777 , n6288 );
    or g6839 ( n11979 , n32857 , n32272 );
    and g6840 ( n15291 , n18939 , n23510 );
    or g6841 ( n12865 , n14200 , n10139 );
    xnor g6842 ( n22965 , n8797 , n12431 );
    or g6843 ( n28282 , n954 , n12966 );
    and g6844 ( n3291 , n23964 , n28832 );
    or g6845 ( n4794 , n9717 , n6554 );
    or g6846 ( n6039 , n11120 , n24653 );
    or g6847 ( n35818 , n3222 , n9588 );
    or g6848 ( n29455 , n27399 , n32930 );
    not g6849 ( n8879 , n9658 );
    and g6850 ( n23026 , n33619 , n29275 );
    xnor g6851 ( n5489 , n18748 , n20664 );
    not g6852 ( n1041 , n3480 );
    or g6853 ( n30240 , n1359 , n18811 );
    xnor g6854 ( n7756 , n7654 , n8432 );
    or g6855 ( n25029 , n21715 , n17046 );
    or g6856 ( n31454 , n33436 , n20840 );
    and g6857 ( n25684 , n25655 , n20551 );
    or g6858 ( n30535 , n9658 , n14445 );
    or g6859 ( n24443 , n15403 , n21832 );
    not g6860 ( n7748 , n18296 );
    xnor g6861 ( n1466 , n10887 , n9658 );
    or g6862 ( n23520 , n30790 , n20318 );
    or g6863 ( n27415 , n12643 , n33227 );
    xnor g6864 ( n35344 , n35404 , n30742 );
    xnor g6865 ( n12708 , n4381 , n5975 );
    or g6866 ( n26990 , n12938 , n17974 );
    or g6867 ( n33196 , n12380 , n11163 );
    or g6868 ( n13382 , n31966 , n12996 );
    or g6869 ( n29032 , n27956 , n21923 );
    or g6870 ( n3190 , n24371 , n8438 );
    xnor g6871 ( n22599 , n14025 , n4928 );
    or g6872 ( n3698 , n29839 , n10112 );
    nor g6873 ( n2282 , n879 , n15566 );
    and g6874 ( n35608 , n19798 , n34255 );
    nor g6875 ( n14290 , n4288 , n19524 );
    or g6876 ( n27586 , n11041 , n8723 );
    xnor g6877 ( n30573 , n34258 , n16922 );
    or g6878 ( n24987 , n27062 , n5972 );
    and g6879 ( n12281 , n18961 , n35489 );
    and g6880 ( n18938 , n9423 , n2857 );
    and g6881 ( n4930 , n7613 , n7069 );
    xnor g6882 ( n11368 , n3532 , n4962 );
    and g6883 ( n10855 , n18940 , n24197 );
    xor g6884 ( n14826 , n6567 , n33960 );
    or g6885 ( n3130 , n7365 , n20308 );
    xnor g6886 ( n2318 , n32953 , n18143 );
    xnor g6887 ( n15759 , n24646 , n17898 );
    xnor g6888 ( n14653 , n26275 , n8432 );
    or g6889 ( n33266 , n3668 , n30305 );
    xnor g6890 ( n10174 , n17729 , n9789 );
    or g6891 ( n16181 , n20030 , n11977 );
    or g6892 ( n18145 , n30144 , n3858 );
    or g6893 ( n592 , n31215 , n34623 );
    and g6894 ( n791 , n4479 , n35626 );
    and g6895 ( n33880 , n13488 , n10569 );
    xnor g6896 ( n5766 , n15807 , n4047 );
    and g6897 ( n20732 , n11065 , n1426 );
    or g6898 ( n8082 , n25793 , n29266 );
    nor g6899 ( n19443 , n29713 , n31087 );
    or g6900 ( n27296 , n4131 , n25255 );
    xnor g6901 ( n10360 , n1304 , n508 );
    not g6902 ( n28398 , n17568 );
    xnor g6903 ( n13064 , n22586 , n17092 );
    xnor g6904 ( n17195 , n17919 , n32738 );
    or g6905 ( n12759 , n27290 , n22682 );
    and g6906 ( n33192 , n9061 , n25056 );
    or g6907 ( n15636 , n20888 , n32071 );
    or g6908 ( n10853 , n3222 , n5917 );
    or g6909 ( n34881 , n30911 , n8328 );
    or g6910 ( n11098 , n22277 , n23790 );
    xnor g6911 ( n12266 , n10454 , n18710 );
    and g6912 ( n21061 , n10672 , n23417 );
    xnor g6913 ( n35118 , n7646 , n10894 );
    or g6914 ( n15275 , n22292 , n3352 );
    and g6915 ( n6159 , n3273 , n13472 );
    or g6916 ( n24373 , n6063 , n20515 );
    and g6917 ( n8341 , n1513 , n9350 );
    or g6918 ( n7563 , n24332 , n20267 );
    or g6919 ( n30676 , n832 , n27728 );
    xnor g6920 ( n22810 , n33569 , n31799 );
    and g6921 ( n9301 , n18124 , n18735 );
    or g6922 ( n9634 , n29839 , n29802 );
    or g6923 ( n31609 , n25414 , n15538 );
    or g6924 ( n12690 , n23604 , n33716 );
    xnor g6925 ( n5257 , n19886 , n23201 );
    or g6926 ( n5986 , n12802 , n16456 );
    or g6927 ( n31754 , n35060 , n12876 );
    or g6928 ( n18389 , n1343 , n3736 );
    xnor g6929 ( n7766 , n4427 , n10583 );
    and g6930 ( n18383 , n17490 , n3836 );
    nor g6931 ( n20563 , n3205 , n12590 );
    or g6932 ( n16255 , n6828 , n27574 );
    nor g6933 ( n21723 , n12732 , n13302 );
    or g6934 ( n13754 , n5794 , n22858 );
    or g6935 ( n13836 , n7540 , n30282 );
    and g6936 ( n21330 , n14305 , n19239 );
    xnor g6937 ( n26379 , n31364 , n19690 );
    or g6938 ( n26412 , n19668 , n33310 );
    or g6939 ( n31868 , n30517 , n18052 );
    or g6940 ( n10493 , n7411 , n32507 );
    or g6941 ( n15885 , n21951 , n26480 );
    xnor g6942 ( n14565 , n5606 , n6930 );
    or g6943 ( n6162 , n27604 , n20553 );
    nor g6944 ( n7727 , n34976 , n30431 );
    or g6945 ( n32144 , n18839 , n183 );
    buf g6946 ( n28675 , n13216 );
    and g6947 ( n20148 , n23137 , n19495 );
    and g6948 ( n4366 , n9491 , n31979 );
    not g6949 ( n14582 , n12301 );
    and g6950 ( n34761 , n30477 , n16335 );
    nor g6951 ( n27614 , n19551 , n2232 );
    or g6952 ( n3377 , n9900 , n17364 );
    or g6953 ( n11860 , n28760 , n4363 );
    xnor g6954 ( n9222 , n8948 , n9658 );
    or g6955 ( n19279 , n30816 , n12622 );
    or g6956 ( n22787 , n17206 , n34084 );
    or g6957 ( n609 , n3946 , n34 );
    nor g6958 ( n3257 , n35718 , n24634 );
    or g6959 ( n14870 , n22031 , n5457 );
    or g6960 ( n23000 , n18326 , n655 );
    xnor g6961 ( n27452 , n5253 , n2672 );
    and g6962 ( n849 , n12065 , n28253 );
    or g6963 ( n507 , n32508 , n18127 );
    and g6964 ( n11233 , n25296 , n31344 );
    and g6965 ( n17991 , n33393 , n12762 );
    xnor g6966 ( n17292 , n30955 , n18161 );
    or g6967 ( n27733 , n21896 , n19732 );
    and g6968 ( n13338 , n32542 , n12060 );
    nor g6969 ( n27617 , n15299 , n29647 );
    or g6970 ( n22374 , n9818 , n20827 );
    and g6971 ( n11959 , n26277 , n24918 );
    nor g6972 ( n11165 , n4288 , n32404 );
    or g6973 ( n1367 , n20598 , n33723 );
    xnor g6974 ( n21214 , n5995 , n27226 );
    and g6975 ( n26238 , n31246 , n7554 );
    xnor g6976 ( n2018 , n4690 , n9604 );
    xnor g6977 ( n10393 , n9549 , n4878 );
    or g6978 ( n20524 , n15464 , n10027 );
    or g6979 ( n27810 , n28181 , n33034 );
    or g6980 ( n16447 , n3503 , n7373 );
    or g6981 ( n28270 , n12257 , n9317 );
    not g6982 ( n14963 , n13784 );
    xnor g6983 ( n14811 , n856 , n24547 );
    nor g6984 ( n25510 , n7857 , n17368 );
    not g6985 ( n9115 , n4210 );
    and g6986 ( n18486 , n65 , n22908 );
    or g6987 ( n10969 , n9052 , n24479 );
    or g6988 ( n34506 , n12351 , n13015 );
    or g6989 ( n31893 , n32095 , n26676 );
    xnor g6990 ( n22344 , n5049 , n4715 );
    or g6991 ( n6264 , n623 , n5395 );
    nor g6992 ( n3504 , n16620 , n17470 );
    or g6993 ( n19408 , n7540 , n17532 );
    and g6994 ( n3838 , n29179 , n32012 );
    or g6995 ( n16437 , n28417 , n11833 );
    nor g6996 ( n9460 , n5335 , n15191 );
    or g6997 ( n20795 , n8059 , n23741 );
    xnor g6998 ( n20825 , n17875 , n13000 );
    xnor g6999 ( n14109 , n180 , n34218 );
    xnor g7000 ( n7155 , n26568 , n31289 );
    and g7001 ( n8663 , n18154 , n16266 );
    and g7002 ( n33138 , n23745 , n9620 );
    xnor g7003 ( n9416 , n11333 , n14563 );
    or g7004 ( n21295 , n22289 , n20576 );
    or g7005 ( n15323 , n33652 , n7293 );
    or g7006 ( n10851 , n22291 , n22437 );
    not g7007 ( n8139 , n30204 );
    or g7008 ( n21087 , n22426 , n9899 );
    or g7009 ( n20221 , n19906 , n4175 );
    not g7010 ( n15581 , n6987 );
    or g7011 ( n17328 , n13299 , n11712 );
    xnor g7012 ( n24107 , n12458 , n8432 );
    and g7013 ( n6748 , n8946 , n29832 );
    xnor g7014 ( n9895 , n12565 , n9658 );
    not g7015 ( n10264 , n16326 );
    xnor g7016 ( n7528 , n13142 , n16620 );
    or g7017 ( n33768 , n11414 , n31739 );
    and g7018 ( n14728 , n14502 , n11256 );
    xnor g7019 ( n1192 , n10404 , n3730 );
    xnor g7020 ( n26021 , n1015 , n3946 );
    and g7021 ( n9253 , n33768 , n1664 );
    not g7022 ( n22624 , n30295 );
    xnor g7023 ( n33016 , n24810 , n31799 );
    xnor g7024 ( n9964 , n22614 , n24371 );
    xnor g7025 ( n4984 , n18849 , n30077 );
    xnor g7026 ( n6363 , n19272 , n12222 );
    xnor g7027 ( n16225 , n19347 , n8273 );
    or g7028 ( n4465 , n31799 , n13158 );
    or g7029 ( n35578 , n11190 , n29194 );
    not g7030 ( n23549 , n16620 );
    not g7031 ( n19542 , n16575 );
    or g7032 ( n31647 , n30348 , n33379 );
    or g7033 ( n33527 , n5949 , n25786 );
    and g7034 ( n9072 , n13327 , n10180 );
    xnor g7035 ( n16971 , n24968 , n3946 );
    and g7036 ( n10463 , n12184 , n27684 );
    or g7037 ( n16498 , n15930 , n12057 );
    or g7038 ( n32188 , n15081 , n27251 );
    or g7039 ( n32345 , n28289 , n35630 );
    or g7040 ( n25229 , n16620 , n16279 );
    or g7041 ( n28162 , n2961 , n29643 );
    xnor g7042 ( n15779 , n10742 , n17848 );
    and g7043 ( n9631 , n15958 , n19073 );
    and g7044 ( n23737 , n7135 , n23957 );
    and g7045 ( n5094 , n19491 , n1123 );
    or g7046 ( n27112 , n30746 , n27518 );
    and g7047 ( n32335 , n24734 , n15845 );
    or g7048 ( n2679 , n25478 , n15517 );
    and g7049 ( n24286 , n5859 , n2461 );
    nor g7050 ( n12438 , n17303 , n10690 );
    or g7051 ( n17388 , n11046 , n21396 );
    or g7052 ( n21174 , n16922 , n11338 );
    xnor g7053 ( n32939 , n13527 , n11077 );
    and g7054 ( n23438 , n24137 , n35809 );
    and g7055 ( n31906 , n27103 , n19842 );
    and g7056 ( n32769 , n13072 , n12597 );
    not g7057 ( n26117 , n17066 );
    or g7058 ( n25875 , n26719 , n17125 );
    xnor g7059 ( n20566 , n12161 , n21468 );
    xnor g7060 ( n6009 , n19530 , n17751 );
    nor g7061 ( n34571 , n16652 , n30463 );
    not g7062 ( n28323 , n3842 );
    and g7063 ( n2325 , n33771 , n17720 );
    or g7064 ( n4665 , n1197 , n2384 );
    or g7065 ( n26394 , n14415 , n2798 );
    or g7066 ( n26301 , n11344 , n26002 );
    nor g7067 ( n30222 , n33732 , n14672 );
    or g7068 ( n20796 , n14662 , n16961 );
    or g7069 ( n2804 , n21165 , n26589 );
    or g7070 ( n2777 , n8382 , n15547 );
    or g7071 ( n2306 , n3669 , n16345 );
    or g7072 ( n34581 , n31957 , n9832 );
    xnor g7073 ( n33497 , n31242 , n19657 );
    or g7074 ( n501 , n9568 , n24141 );
    xnor g7075 ( n25159 , n20366 , n4675 );
    and g7076 ( n10908 , n16295 , n15777 );
    xnor g7077 ( n28911 , n28307 , n9782 );
    or g7078 ( n24393 , n10894 , n19768 );
    or g7079 ( n16136 , n6067 , n544 );
    xnor g7080 ( n9457 , n31569 , n30513 );
    xnor g7081 ( n32436 , n24863 , n5456 );
    and g7082 ( n7555 , n9489 , n14277 );
    xnor g7083 ( n25048 , n33657 , n27997 );
    or g7084 ( n29925 , n21040 , n17829 );
    or g7085 ( n11657 , n5839 , n8766 );
    or g7086 ( n20507 , n23760 , n31554 );
    and g7087 ( n17027 , n11310 , n10043 );
    not g7088 ( n11705 , n2827 );
    and g7089 ( n11055 , n5851 , n26169 );
    xnor g7090 ( n8382 , n14327 , n9658 );
    not g7091 ( n17881 , n16922 );
    and g7092 ( n13869 , n14442 , n26738 );
    nor g7093 ( n28605 , n25037 , n35954 );
    or g7094 ( n299 , n16620 , n19018 );
    and g7095 ( n25139 , n30043 , n9799 );
    or g7096 ( n15524 , n11046 , n32304 );
    and g7097 ( n33668 , n29392 , n5986 );
    or g7098 ( n5851 , n2657 , n26032 );
    and g7099 ( n13094 , n21256 , n42 );
    or g7100 ( n22094 , n13149 , n17354 );
    or g7101 ( n15888 , n26048 , n1942 );
    or g7102 ( n11662 , n25174 , n25764 );
    and g7103 ( n13948 , n11864 , n5667 );
    or g7104 ( n1894 , n16415 , n21673 );
    nor g7105 ( n11943 , n23604 , n31387 );
    or g7106 ( n22903 , n3720 , n20669 );
    and g7107 ( n14246 , n29207 , n18410 );
    and g7108 ( n22865 , n15151 , n1880 );
    nor g7109 ( n35787 , n26701 , n33157 );
    or g7110 ( n16321 , n21432 , n19579 );
    and g7111 ( n11698 , n24480 , n32000 );
    and g7112 ( n1757 , n6174 , n14234 );
    and g7113 ( n6912 , n8599 , n1101 );
    or g7114 ( n25981 , n27822 , n18477 );
    xnor g7115 ( n16886 , n31999 , n1950 );
    and g7116 ( n11673 , n27412 , n28298 );
    xnor g7117 ( n26030 , n9980 , n21372 );
    or g7118 ( n18140 , n3994 , n12128 );
    or g7119 ( n16850 , n7616 , n6075 );
    or g7120 ( n22769 , n8432 , n4170 );
    or g7121 ( n15783 , n4288 , n15037 );
    or g7122 ( n4046 , n33454 , n24356 );
    or g7123 ( n35845 , n14079 , n18811 );
    xnor g7124 ( n31305 , n25715 , n11782 );
    and g7125 ( n13601 , n26593 , n26661 );
    nor g7126 ( n12030 , n12160 , n16770 );
    and g7127 ( n34691 , n21316 , n25184 );
    or g7128 ( n23354 , n32382 , n30292 );
    or g7129 ( n2736 , n27367 , n21019 );
    or g7130 ( n12280 , n26973 , n22206 );
    or g7131 ( n13357 , n18087 , n24489 );
    buf g7132 ( n10140 , n12869 );
    xnor g7133 ( n15972 , n34023 , n5295 );
    and g7134 ( n11472 , n16303 , n793 );
    or g7135 ( n26373 , n2397 , n8937 );
    or g7136 ( n1298 , n25102 , n28438 );
    or g7137 ( n10344 , n13033 , n32425 );
    xnor g7138 ( n33837 , n3814 , n14800 );
    or g7139 ( n29962 , n27544 , n8254 );
    xnor g7140 ( n10030 , n27885 , n15299 );
    or g7141 ( n15485 , n14336 , n20318 );
    or g7142 ( n16226 , n16105 , n21873 );
    xnor g7143 ( n35672 , n1316 , n3115 );
    or g7144 ( n23012 , n21457 , n25773 );
    xnor g7145 ( n26743 , n10941 , n27512 );
    and g7146 ( n9517 , n28872 , n24584 );
    or g7147 ( n27918 , n34955 , n10417 );
    xnor g7148 ( n26330 , n11745 , n19154 );
    or g7149 ( n15575 , n35855 , n16543 );
    or g7150 ( n10937 , n29387 , n14844 );
    and g7151 ( n22947 , n34652 , n5072 );
    not g7152 ( n616 , n21359 );
    and g7153 ( n3 , n3896 , n17693 );
    nor g7154 ( n15431 , n24371 , n996 );
    and g7155 ( n34696 , n25916 , n23571 );
    or g7156 ( n14952 , n20180 , n29953 );
    or g7157 ( n21398 , n34040 , n12001 );
    or g7158 ( n21958 , n31215 , n781 );
    xnor g7159 ( n15032 , n34613 , n16301 );
    or g7160 ( n21319 , n29010 , n33416 );
    or g7161 ( n8548 , n22531 , n24489 );
    not g7162 ( n24627 , n9383 );
    not g7163 ( n13840 , n4520 );
    and g7164 ( n10166 , n30138 , n25064 );
    not g7165 ( n23027 , n25174 );
    or g7166 ( n24901 , n11991 , n3842 );
    xnor g7167 ( n26941 , n33311 , n3205 );
    or g7168 ( n26020 , n14477 , n33098 );
    and g7169 ( n6210 , n5188 , n25199 );
    xnor g7170 ( n11997 , n35786 , n1950 );
    or g7171 ( n8069 , n14288 , n24317 );
    or g7172 ( n15237 , n20531 , n19173 );
    and g7173 ( n32740 , n18789 , n19196 );
    or g7174 ( n29646 , n23310 , n26292 );
    or g7175 ( n21904 , n29839 , n18208 );
    or g7176 ( n8633 , n12999 , n20690 );
    or g7177 ( n7938 , n30053 , n23462 );
    or g7178 ( n22862 , n20746 , n7931 );
    or g7179 ( n30743 , n21273 , n8833 );
    and g7180 ( n35235 , n7915 , n9793 );
    or g7181 ( n35066 , n33569 , n559 );
    and g7182 ( n23118 , n7145 , n1209 );
    xnor g7183 ( n28922 , n4801 , n32857 );
    or g7184 ( n10726 , n16922 , n639 );
    xnor g7185 ( n34719 , n30442 , n24560 );
    and g7186 ( n27420 , n7839 , n8370 );
    or g7187 ( n23188 , n1950 , n31311 );
    and g7188 ( n7823 , n35435 , n16443 );
    or g7189 ( n27916 , n35089 , n20762 );
    nor g7190 ( n14762 , n4960 , n17307 );
    or g7191 ( n35474 , n8455 , n15344 );
    xnor g7192 ( n6430 , n28901 , n5335 );
    or g7193 ( n1579 , n29719 , n5103 );
    xnor g7194 ( n4599 , n12212 , n7773 );
    or g7195 ( n13152 , n6092 , n28404 );
    or g7196 ( n868 , n4322 , n556 );
    or g7197 ( n18350 , n5243 , n2104 );
    or g7198 ( n11913 , n17996 , n6340 );
    and g7199 ( n13117 , n8291 , n12889 );
    not g7200 ( n11776 , n7769 );
    and g7201 ( n4231 , n35440 , n32957 );
    xor g7202 ( n26867 , n34627 , n26033 );
    not g7203 ( n12744 , n19828 );
    and g7204 ( n18253 , n13919 , n1085 );
    xnor g7205 ( n17619 , n35537 , n33192 );
    xnor g7206 ( n20659 , n11625 , n10081 );
    and g7207 ( n35916 , n10049 , n15504 );
    or g7208 ( n5836 , n20411 , n11218 );
    xnor g7209 ( n19873 , n10623 , n26577 );
    or g7210 ( n30957 , n5013 , n808 );
    or g7211 ( n32204 , n6275 , n21644 );
    or g7212 ( n34564 , n32766 , n14361 );
    nor g7213 ( n33265 , n29600 , n26467 );
    nor g7214 ( n28225 , n21907 , n1176 );
    and g7215 ( n20486 , n11301 , n26182 );
    or g7216 ( n9644 , n19591 , n21977 );
    buf g7217 ( n11593 , n11833 );
    and g7218 ( n5960 , n1469 , n5583 );
    xnor g7219 ( n18669 , n10366 , n32666 );
    or g7220 ( n14863 , n23351 , n3188 );
    or g7221 ( n7258 , n1676 , n17306 );
    or g7222 ( n33278 , n32725 , n25447 );
    not g7223 ( n3252 , n17628 );
    and g7224 ( n2590 , n34695 , n12148 );
    or g7225 ( n16195 , n14109 , n27801 );
    and g7226 ( n20768 , n22073 , n8475 );
    or g7227 ( n4850 , n31052 , n26480 );
    xnor g7228 ( n6595 , n13714 , n32715 );
    xnor g7229 ( n14541 , n12433 , n7540 );
    or g7230 ( n10238 , n7063 , n29366 );
    xnor g7231 ( n26053 , n35907 , n9793 );
    not g7232 ( n10195 , n15917 );
    not g7233 ( n28286 , n4878 );
    or g7234 ( n31036 , n8481 , n2814 );
    xnor g7235 ( n6477 , n22069 , n2543 );
    xnor g7236 ( n9978 , n31165 , n19440 );
    or g7237 ( n32252 , n13583 , n542 );
    or g7238 ( n6695 , n31578 , n11892 );
    or g7239 ( n11493 , n11038 , n33396 );
    or g7240 ( n2316 , n16750 , n24653 );
    and g7241 ( n5791 , n34980 , n21187 );
    or g7242 ( n15093 , n1135 , n3437 );
    or g7243 ( n35829 , n35988 , n12596 );
    or g7244 ( n1729 , n4288 , n24363 );
    not g7245 ( n22276 , n26683 );
    or g7246 ( n4371 , n11046 , n16209 );
    nor g7247 ( n32309 , n31187 , n4161 );
    or g7248 ( n31866 , n19760 , n5779 );
    nor g7249 ( n10283 , n32095 , n5096 );
    or g7250 ( n8961 , n15376 , n28064 );
    and g7251 ( n4076 , n11869 , n21871 );
    and g7252 ( n15539 , n21817 , n22980 );
    xnor g7253 ( n16638 , n32170 , n5171 );
    or g7254 ( n8411 , n10910 , n7673 );
    not g7255 ( n35545 , n2327 );
    xnor g7256 ( n23636 , n12916 , n15299 );
    and g7257 ( n34270 , n206 , n18133 );
    or g7258 ( n27076 , n19886 , n23201 );
    and g7259 ( n2216 , n4274 , n26016 );
    and g7260 ( n17042 , n24797 , n14524 );
    xnor g7261 ( n25084 , n7564 , n4288 );
    nor g7262 ( n5578 , n16620 , n23350 );
    or g7263 ( n9433 , n32174 , n34600 );
    or g7264 ( n26898 , n9493 , n19544 );
    or g7265 ( n16546 , n521 , n5208 );
    or g7266 ( n4503 , n4962 , n3966 );
    or g7267 ( n22770 , n11927 , n35935 );
    or g7268 ( n28471 , n11442 , n8366 );
    or g7269 ( n18799 , n21193 , n949 );
    or g7270 ( n20297 , n2305 , n1856 );
    or g7271 ( n36056 , n34842 , n34971 );
    xnor g7272 ( n11031 , n22892 , n20732 );
    and g7273 ( n27505 , n22015 , n21640 );
    or g7274 ( n5321 , n29559 , n29052 );
    and g7275 ( n9480 , n1233 , n6971 );
    nor g7276 ( n26151 , n17568 , n25346 );
    nor g7277 ( n18382 , n16922 , n14682 );
    or g7278 ( n6737 , n4321 , n23891 );
    buf g7279 ( n25019 , n4175 );
    and g7280 ( n14709 , n12337 , n21997 );
    and g7281 ( n7649 , n34217 , n22232 );
    or g7282 ( n22898 , n28087 , n12353 );
    or g7283 ( n3007 , n14941 , n9104 );
    or g7284 ( n1614 , n21391 , n11459 );
    and g7285 ( n11002 , n14027 , n32511 );
    not g7286 ( n11460 , n15546 );
    nor g7287 ( n16438 , n33413 , n29366 );
    or g7288 ( n31093 , n4116 , n5741 );
    or g7289 ( n32514 , n32864 , n36000 );
    and g7290 ( n3317 , n32662 , n22980 );
    xnor g7291 ( n723 , n28927 , n11455 );
    or g7292 ( n31776 , n2187 , n8379 );
    and g7293 ( n31815 , n26454 , n15354 );
    and g7294 ( n26927 , n8678 , n14518 );
    or g7295 ( n35919 , n4630 , n12332 );
    and g7296 ( n24140 , n25022 , n8889 );
    buf g7297 ( n5900 , n4361 );
    or g7298 ( n24965 , n33539 , n363 );
    or g7299 ( n29046 , n17745 , n31285 );
    xnor g7300 ( n21591 , n30231 , n29970 );
    xnor g7301 ( n14031 , n18518 , n18379 );
    xnor g7302 ( n28735 , n26823 , n35927 );
    or g7303 ( n5827 , n22337 , n1970 );
    xnor g7304 ( n2193 , n32402 , n6032 );
    nor g7305 ( n17941 , n28463 , n6548 );
    and g7306 ( n2771 , n15612 , n25816 );
    not g7307 ( n25924 , n34396 );
    and g7308 ( n17633 , n12766 , n12559 );
    not g7309 ( n6651 , n1950 );
    and g7310 ( n27539 , n21309 , n25361 );
    xnor g7311 ( n2678 , n566 , n30742 );
    xnor g7312 ( n13957 , n31703 , n7113 );
    not g7313 ( n22457 , n32067 );
    and g7314 ( n3780 , n29472 , n29641 );
    xnor g7315 ( n2965 , n3895 , n33398 );
    or g7316 ( n15758 , n10894 , n14688 );
    or g7317 ( n12607 , n10920 , n34089 );
    or g7318 ( n31315 , n7321 , n18264 );
    and g7319 ( n6559 , n7574 , n27829 );
    and g7320 ( n7177 , n16441 , n8009 );
    and g7321 ( n26429 , n20591 , n3767 );
    xnor g7322 ( n31610 , n29089 , n33948 );
    or g7323 ( n35635 , n21450 , n2117 );
    xnor g7324 ( n17946 , n29968 , n12005 );
    xnor g7325 ( n3496 , n10594 , n3388 );
    and g7326 ( n21294 , n13342 , n1571 );
    and g7327 ( n21739 , n8139 , n18770 );
    and g7328 ( n4645 , n29129 , n14692 );
    xnor g7329 ( n30942 , n58 , n24878 );
    or g7330 ( n31447 , n32584 , n3892 );
    xnor g7331 ( n27546 , n10798 , n7345 );
    not g7332 ( n30654 , n28969 );
    nor g7333 ( n19675 , n4878 , n15502 );
    and g7334 ( n33440 , n989 , n30275 );
    xnor g7335 ( n17423 , n26070 , n29713 );
    nor g7336 ( n21094 , n28958 , n15184 );
    or g7337 ( n32521 , n3222 , n11713 );
    and g7338 ( n25647 , n12325 , n25516 );
    xnor g7339 ( n19278 , n8514 , n32090 );
    or g7340 ( n21262 , n28345 , n33901 );
    or g7341 ( n19538 , n5655 , n1796 );
    or g7342 ( n977 , n22363 , n29953 );
    nor g7343 ( n11765 , n4960 , n16534 );
    xnor g7344 ( n27130 , n20981 , n15518 );
    or g7345 ( n22250 , n10878 , n17125 );
    and g7346 ( n17469 , n35099 , n19494 );
    xnor g7347 ( n4011 , n2118 , n830 );
    not g7348 ( n2727 , n3205 );
    or g7349 ( n10538 , n18165 , n35143 );
    or g7350 ( n3309 , n27452 , n18017 );
    xnor g7351 ( n17965 , n6421 , n15552 );
    and g7352 ( n11774 , n1047 , n26236 );
    xnor g7353 ( n12999 , n13941 , n14570 );
    and g7354 ( n18164 , n31880 , n3285 );
    and g7355 ( n16228 , n12861 , n19039 );
    and g7356 ( n14075 , n13264 , n6045 );
    and g7357 ( n5881 , n23228 , n13803 );
    xnor g7358 ( n18750 , n16925 , n22291 );
    or g7359 ( n22905 , n25698 , n15439 );
    and g7360 ( n25845 , n27703 , n17144 );
    not g7361 ( n19137 , n28273 );
    and g7362 ( n27603 , n24674 , n34714 );
    or g7363 ( n23839 , n34987 , n16797 );
    buf g7364 ( n22961 , n544 );
    or g7365 ( n26592 , n16922 , n29083 );
    not g7366 ( n6712 , n27786 );
    and g7367 ( n405 , n24980 , n7552 );
    or g7368 ( n15137 , n13636 , n30519 );
    or g7369 ( n15500 , n22765 , n22946 );
    or g7370 ( n20355 , n5110 , n17162 );
    xnor g7371 ( n9715 , n22818 , n24389 );
    and g7372 ( n19376 , n23441 , n11857 );
    or g7373 ( n22249 , n4962 , n6591 );
    not g7374 ( n24723 , n34677 );
    or g7375 ( n35650 , n3572 , n6107 );
    or g7376 ( n1731 , n18576 , n23396 );
    or g7377 ( n8306 , n25602 , n14043 );
    and g7378 ( n6829 , n8415 , n33032 );
    xnor g7379 ( n28486 , n15767 , n16086 );
    or g7380 ( n2676 , n17941 , n31674 );
    or g7381 ( n2670 , n33354 , n16961 );
    xnor g7382 ( n14629 , n17038 , n24486 );
    not g7383 ( n34011 , n29713 );
    xnor g7384 ( n27953 , n18745 , n19257 );
    or g7385 ( n12386 , n25788 , n34484 );
    or g7386 ( n6597 , n32230 , n16943 );
    and g7387 ( n30216 , n16094 , n29690 );
    or g7388 ( n27330 , n23076 , n19493 );
    nor g7389 ( n1375 , n21664 , n22847 );
    or g7390 ( n33059 , n20387 , n22316 );
    not g7391 ( n30478 , n2780 );
    or g7392 ( n26073 , n9793 , n30393 );
    xnor g7393 ( n12300 , n22082 , n16135 );
    xnor g7394 ( n13475 , n23764 , n15403 );
    or g7395 ( n7497 , n8407 , n3756 );
    or g7396 ( n19092 , n24371 , n4826 );
    xnor g7397 ( n11228 , n12989 , n23360 );
    xnor g7398 ( n2936 , n6907 , n9658 );
    and g7399 ( n18569 , n25574 , n9469 );
    xnor g7400 ( n35024 , n19429 , n10607 );
    or g7401 ( n8281 , n25991 , n26296 );
    xnor g7402 ( n30004 , n31216 , n23735 );
    and g7403 ( n9386 , n10652 , n3555 );
    not g7404 ( n4426 , n11996 );
    or g7405 ( n7405 , n34274 , n9951 );
    xnor g7406 ( n12167 , n11164 , n4962 );
    and g7407 ( n11749 , n2900 , n33363 );
    and g7408 ( n7918 , n25546 , n24186 );
    xnor g7409 ( n14415 , n6667 , n10028 );
    or g7410 ( n6724 , n12102 , n9947 );
    or g7411 ( n17383 , n1978 , n24653 );
    or g7412 ( n16127 , n21551 , n14554 );
    and g7413 ( n27758 , n7757 , n1684 );
    or g7414 ( n16913 , n2949 , n30732 );
    xnor g7415 ( n9125 , n34681 , n32049 );
    or g7416 ( n12037 , n7172 , n23209 );
    nor g7417 ( n29092 , n24775 , n24556 );
    xnor g7418 ( n4816 , n26389 , n30091 );
    not g7419 ( n23910 , n7555 );
    or g7420 ( n26749 , n24662 , n35141 );
    and g7421 ( n9592 , n29305 , n6797 );
    and g7422 ( n28051 , n10863 , n36025 );
    xnor g7423 ( n5056 , n17672 , n21162 );
    or g7424 ( n20759 , n5489 , n3805 );
    nor g7425 ( n23751 , n23604 , n15985 );
    or g7426 ( n6362 , n7540 , n26472 );
    or g7427 ( n32383 , n10027 , n17125 );
    or g7428 ( n18511 , n4962 , n30987 );
    or g7429 ( n25100 , n20961 , n12332 );
    or g7430 ( n34299 , n17161 , n34693 );
    and g7431 ( n11522 , n5974 , n28408 );
    xnor g7432 ( n26044 , n9821 , n26756 );
    nor g7433 ( n9818 , n4960 , n8372 );
    or g7434 ( n30178 , n3721 , n14794 );
    or g7435 ( n34167 , n7416 , n35937 );
    nor g7436 ( n30268 , n9116 , n7448 );
    xnor g7437 ( n31420 , n21497 , n30742 );
    xnor g7438 ( n33554 , n3099 , n30742 );
    xnor g7439 ( n3406 , n36087 , n11455 );
    and g7440 ( n12209 , n11430 , n7045 );
    and g7441 ( n26477 , n34502 , n895 );
    not g7442 ( n7814 , n22980 );
    or g7443 ( n16325 , n34666 , n9670 );
    or g7444 ( n17796 , n11046 , n16711 );
    or g7445 ( n5831 , n11046 , n29984 );
    or g7446 ( n1545 , n4710 , n17233 );
    or g7447 ( n11736 , n35927 , n30334 );
    xnor g7448 ( n33333 , n3540 , n31056 );
    not g7449 ( n30365 , n28273 );
    and g7450 ( n4059 , n6497 , n28025 );
    and g7451 ( n12470 , n18693 , n15746 );
    and g7452 ( n14683 , n4006 , n33445 );
    nor g7453 ( n17509 , n22135 , n18115 );
    xnor g7454 ( n28965 , n28318 , n19551 );
    and g7455 ( n18801 , n10991 , n14608 );
    or g7456 ( n21966 , n32857 , n14387 );
    and g7457 ( n34135 , n4207 , n24805 );
    xnor g7458 ( n29162 , n31425 , n28135 );
    and g7459 ( n35891 , n10757 , n2704 );
    xnor g7460 ( n19276 , n28709 , n8738 );
    or g7461 ( n18457 , n14435 , n21456 );
    or g7462 ( n4479 , n4409 , n19105 );
    nor g7463 ( n11635 , n9111 , n33956 );
    and g7464 ( n5139 , n17508 , n6610 );
    nor g7465 ( n32871 , n26695 , n35498 );
    nor g7466 ( n30897 , n10894 , n7495 );
    or g7467 ( n16784 , n24371 , n20572 );
    or g7468 ( n33835 , n35927 , n20875 );
    xnor g7469 ( n11304 , n19948 , n5476 );
    xnor g7470 ( n9339 , n2509 , n27186 );
    xnor g7471 ( n32747 , n13763 , n25052 );
    nor g7472 ( n16033 , n18988 , n31232 );
    and g7473 ( n14605 , n31860 , n32700 );
    or g7474 ( n11564 , n7033 , n21691 );
    xnor g7475 ( n18261 , n33875 , n29713 );
    and g7476 ( n12494 , n11325 , n7476 );
    or g7477 ( n3953 , n15403 , n9325 );
    and g7478 ( n5278 , n4883 , n18347 );
    xnor g7479 ( n21201 , n31084 , n31147 );
    or g7480 ( n29099 , n23455 , n11593 );
    and g7481 ( n21055 , n12598 , n32183 );
    xnor g7482 ( n30638 , n13445 , n23801 );
    and g7483 ( n15531 , n2043 , n24951 );
    and g7484 ( n31687 , n14333 , n20876 );
    or g7485 ( n28029 , n11603 , n4363 );
    or g7486 ( n19227 , n17767 , n1796 );
    or g7487 ( n3230 , n34767 , n16543 );
    and g7488 ( n23504 , n23437 , n27906 );
    nor g7489 ( n22382 , n4758 , n14739 );
    xnor g7490 ( n22518 , n25118 , n34002 );
    and g7491 ( n2984 , n28937 , n5229 );
    xnor g7492 ( n13867 , n12346 , n3308 );
    xnor g7493 ( n34074 , n25520 , n34315 );
    xnor g7494 ( n23306 , n6634 , n11841 );
    or g7495 ( n16480 , n2601 , n35603 );
    or g7496 ( n25215 , n12680 , n15112 );
    not g7497 ( n17801 , n11046 );
    xnor g7498 ( n7809 , n24458 , n29713 );
    or g7499 ( n18684 , n7318 , n11312 );
    or g7500 ( n23331 , n21927 , n35093 );
    not g7501 ( n25958 , n30742 );
    or g7502 ( n31671 , n17158 , n20427 );
    or g7503 ( n35092 , n23541 , n28668 );
    or g7504 ( n12314 , n7346 , n17337 );
    and g7505 ( n636 , n11388 , n1670 );
    and g7506 ( n7987 , n11815 , n23728 );
    xnor g7507 ( n9566 , n9980 , n4284 );
    and g7508 ( n945 , n20280 , n27378 );
    or g7509 ( n25590 , n35776 , n25761 );
    or g7510 ( n15525 , n15299 , n3707 );
    or g7511 ( n11507 , n9658 , n22470 );
    xnor g7512 ( n23746 , n28695 , n25713 );
    nor g7513 ( n8159 , n31165 , n19440 );
    and g7514 ( n10142 , n14724 , n17460 );
    xnor g7515 ( n3816 , n4641 , n5335 );
    or g7516 ( n29236 , n14821 , n12016 );
    xor g7517 ( n15637 , n23784 , n3003 );
    or g7518 ( n17200 , n21344 , n21974 );
    or g7519 ( n23944 , n8258 , n4363 );
    or g7520 ( n30958 , n1282 , n29592 );
    xnor g7521 ( n13812 , n3128 , n17568 );
    nor g7522 ( n35084 , n24371 , n10623 );
    and g7523 ( n28933 , n19758 , n8499 );
    or g7524 ( n27306 , n28242 , n33416 );
    and g7525 ( n27381 , n9745 , n9180 );
    nor g7526 ( n19293 , n30578 , n25293 );
    or g7527 ( n7513 , n11829 , n26480 );
    nor g7528 ( n10348 , n2459 , n11663 );
    or g7529 ( n8061 , n298 , n33951 );
    and g7530 ( n35371 , n17367 , n6869 );
    xnor g7531 ( n34244 , n20816 , n4878 );
    or g7532 ( n27092 , n32066 , n9955 );
    or g7533 ( n23345 , n18379 , n32058 );
    or g7534 ( n2852 , n830 , n18710 );
    xnor g7535 ( n641 , n2942 , n10715 );
    and g7536 ( n11159 , n29746 , n1820 );
    or g7537 ( n19658 , n23271 , n33098 );
    or g7538 ( n4559 , n24979 , n908 );
    or g7539 ( n17826 , n27622 , n26220 );
    nor g7540 ( n34365 , n32857 , n19878 );
    and g7541 ( n26706 , n23370 , n2929 );
    or g7542 ( n9505 , n5894 , n25255 );
    xnor g7543 ( n6500 , n14978 , n29713 );
    or g7544 ( n8848 , n4960 , n25373 );
    or g7545 ( n32594 , n35318 , n26112 );
    or g7546 ( n35768 , n25174 , n1377 );
    xnor g7547 ( n22186 , n28130 , n13613 );
    or g7548 ( n17168 , n24569 , n7918 );
    or g7549 ( n16346 , n24867 , n33435 );
    or g7550 ( n31600 , n5236 , n6972 );
    and g7551 ( n35913 , n29105 , n136 );
    and g7552 ( n9961 , n31405 , n4615 );
    not g7553 ( n6609 , n30519 );
    and g7554 ( n11179 , n21690 , n30794 );
    or g7555 ( n25734 , n28066 , n21862 );
    or g7556 ( n10834 , n29980 , n13383 );
    and g7557 ( n83 , n35076 , n158 );
    and g7558 ( n3696 , n23835 , n15868 );
    xnor g7559 ( n8992 , n29387 , n14844 );
    and g7560 ( n10099 , n5914 , n14936 );
    or g7561 ( n6636 , n749 , n24785 );
    or g7562 ( n6484 , n31268 , n11035 );
    xnor g7563 ( n13259 , n5939 , n26873 );
    and g7564 ( n13121 , n27930 , n10204 );
    or g7565 ( n22461 , n18379 , n13319 );
    nor g7566 ( n16397 , n4878 , n35947 );
    or g7567 ( n21905 , n6122 , n34270 );
    xnor g7568 ( n23884 , n1328 , n30504 );
    or g7569 ( n16427 , n3579 , n20762 );
    xnor g7570 ( n16062 , n9588 , n3222 );
    and g7571 ( n7127 , n21274 , n22306 );
    and g7572 ( n8109 , n7534 , n30325 );
    and g7573 ( n32838 , n9433 , n33640 );
    not g7574 ( n31967 , n16321 );
    not g7575 ( n263 , n9789 );
    or g7576 ( n25386 , n25854 , n31487 );
    not g7577 ( n16444 , n4960 );
    and g7578 ( n3415 , n428 , n14005 );
    or g7579 ( n32937 , n14254 , n14746 );
    and g7580 ( n13393 , n15196 , n10458 );
    nor g7581 ( n34128 , n30742 , n7110 );
    not g7582 ( n33952 , n31799 );
    and g7583 ( n31362 , n33873 , n20718 );
    xnor g7584 ( n24590 , n19972 , n25174 );
    or g7585 ( n19024 , n5396 , n2955 );
    or g7586 ( n23936 , n31013 , n24704 );
    not g7587 ( n26091 , n19182 );
    or g7588 ( n6342 , n13913 , n33821 );
    or g7589 ( n22853 , n32804 , n35111 );
    xor g7590 ( n13260 , n20030 , n35927 );
    and g7591 ( n26010 , n35896 , n35426 );
    or g7592 ( n3402 , n19586 , n31067 );
    nor g7593 ( n24961 , n3887 , n10709 );
    xnor g7594 ( n15038 , n35598 , n15942 );
    nor g7595 ( n1219 , n2527 , n33243 );
    and g7596 ( n12669 , n33126 , n280 );
    xnor g7597 ( n32585 , n26632 , n17568 );
    and g7598 ( n35451 , n11984 , n29580 );
    or g7599 ( n17684 , n29121 , n32379 );
    or g7600 ( n10121 , n10776 , n8203 );
    and g7601 ( n6726 , n4657 , n27508 );
    or g7602 ( n26343 , n30742 , n33136 );
    xnor g7603 ( n22259 , n6829 , n32857 );
    not g7604 ( n5592 , n311 );
    xnor g7605 ( n17820 , n6400 , n22027 );
    and g7606 ( n5850 , n4688 , n11515 );
    xnor g7607 ( n353 , n6463 , n9793 );
    xnor g7608 ( n10404 , n26055 , n9793 );
    or g7609 ( n27028 , n35701 , n12465 );
    xnor g7610 ( n25721 , n29385 , n13241 );
    xnor g7611 ( n4568 , n292 , n25241 );
    or g7612 ( n30717 , n9658 , n6907 );
    not g7613 ( n16896 , n1528 );
    or g7614 ( n31 , n27228 , n3188 );
    or g7615 ( n4173 , n6761 , n4254 );
    xnor g7616 ( n19273 , n2915 , n17675 );
    or g7617 ( n23969 , n28126 , n19125 );
    or g7618 ( n8916 , n22344 , n3344 );
    and g7619 ( n10402 , n923 , n31752 );
    xnor g7620 ( n2051 , n20715 , n27531 );
    nor g7621 ( n13556 , n17412 , n11511 );
    xnor g7622 ( n14466 , n28622 , n10243 );
    not g7623 ( n27407 , n32857 );
    and g7624 ( n12925 , n22310 , n26776 );
    not g7625 ( n752 , n9793 );
    or g7626 ( n30903 , n22877 , n18858 );
    and g7627 ( n16065 , n19839 , n23750 );
    or g7628 ( n457 , n20229 , n29562 );
    or g7629 ( n23947 , n14885 , n9601 );
    xnor g7630 ( n656 , n13364 , n9793 );
    or g7631 ( n4354 , n28121 , n29290 );
    and g7632 ( n10777 , n5199 , n11649 );
    or g7633 ( n10993 , n3205 , n21488 );
    xnor g7634 ( n31210 , n18601 , n35927 );
    xnor g7635 ( n15808 , n17558 , n12296 );
    or g7636 ( n11542 , n12655 , n29804 );
    or g7637 ( n11700 , n30705 , n13393 );
    not g7638 ( n346 , n17179 );
    and g7639 ( n29887 , n6073 , n6014 );
    xnor g7640 ( n22324 , n3063 , n21077 );
    and g7641 ( n5129 , n15850 , n21828 );
    or g7642 ( n8979 , n32064 , n26023 );
    nor g7643 ( n34430 , n14531 , n32379 );
    not g7644 ( n33399 , n3842 );
    and g7645 ( n20851 , n6021 , n7858 );
    or g7646 ( n21841 , n13387 , n4172 );
    not g7647 ( n19120 , n4769 );
    or g7648 ( n13444 , n11510 , n27564 );
    and g7649 ( n8489 , n29154 , n5641 );
    xnor g7650 ( n1185 , n21596 , n36007 );
    and g7651 ( n20849 , n11558 , n15161 );
    or g7652 ( n32578 , n15191 , n1511 );
    xnor g7653 ( n28030 , n24237 , n32031 );
    or g7654 ( n14199 , n4878 , n34761 );
    not g7655 ( n10902 , n20169 );
    xnor g7656 ( n27757 , n11944 , n17549 );
    and g7657 ( n838 , n13927 , n25720 );
    not g7658 ( n12606 , n15290 );
    or g7659 ( n8734 , n35673 , n32808 );
    buf g7660 ( n13217 , n4036 );
    and g7661 ( n14071 , n27726 , n26097 );
    or g7662 ( n17654 , n9793 , n5412 );
    xnor g7663 ( n3602 , n35443 , n19771 );
    and g7664 ( n11079 , n7771 , n25078 );
    or g7665 ( n2033 , n31799 , n19509 );
    or g7666 ( n1081 , n15881 , n27973 );
    or g7667 ( n22235 , n33632 , n19173 );
    and g7668 ( n3166 , n27798 , n22827 );
    or g7669 ( n3233 , n14057 , n22241 );
    or g7670 ( n7176 , n10110 , n8269 );
    or g7671 ( n14159 , n32584 , n5160 );
    or g7672 ( n5099 , n4962 , n23270 );
    and g7673 ( n33039 , n20612 , n7298 );
    or g7674 ( n17224 , n11993 , n13286 );
    and g7675 ( n16297 , n26344 , n24131 );
    xnor g7676 ( n9281 , n19915 , n7540 );
    nor g7677 ( n19348 , n16315 , n13646 );
    xnor g7678 ( n143 , n19485 , n9789 );
    and g7679 ( n277 , n31434 , n2166 );
    and g7680 ( n32391 , n5043 , n6827 );
    or g7681 ( n28567 , n22526 , n16569 );
    or g7682 ( n20026 , n26159 , n26002 );
    xnor g7683 ( n34149 , n33968 , n3059 );
    and g7684 ( n29843 , n7376 , n33048 );
    or g7685 ( n18186 , n8005 , n19084 );
    nor g7686 ( n3370 , n25602 , n4131 );
    buf g7687 ( n3738 , n21862 );
    or g7688 ( n3991 , n16087 , n25355 );
    xnor g7689 ( n28445 , n4636 , n725 );
    or g7690 ( n24747 , n34414 , n22316 );
    nor g7691 ( n33978 , n30742 , n35719 );
    or g7692 ( n19969 , n32095 , n7881 );
    and g7693 ( n32825 , n22600 , n28450 );
    or g7694 ( n17970 , n28276 , n27305 );
    and g7695 ( n12250 , n24133 , n35194 );
    xnor g7696 ( n13358 , n21706 , n29884 );
    or g7697 ( n7249 , n21602 , n31195 );
    and g7698 ( n1218 , n10259 , n8091 );
    not g7699 ( n28783 , n15638 );
    or g7700 ( n1388 , n31620 , n20068 );
    and g7701 ( n23599 , n17073 , n19067 );
    not g7702 ( n20138 , n3205 );
    and g7703 ( n30290 , n30495 , n9982 );
    or g7704 ( n8065 , n25794 , n8392 );
    or g7705 ( n11539 , n3545 , n15344 );
    or g7706 ( n17032 , n2354 , n28191 );
    not g7707 ( n12437 , n23604 );
    or g7708 ( n13428 , n20465 , n27053 );
    and g7709 ( n13703 , n29814 , n17958 );
    xor g7710 ( n6334 , n5529 , n6331 );
    or g7711 ( n35275 , n29417 , n22051 );
    and g7712 ( n4328 , n22112 , n18959 );
    or g7713 ( n28458 , n23347 , n25107 );
    xnor g7714 ( n35876 , n31793 , n12787 );
    xnor g7715 ( n23833 , n2822 , n33615 );
    or g7716 ( n10650 , n3616 , n2005 );
    xnor g7717 ( n5582 , n20712 , n25174 );
    xnor g7718 ( n32060 , n30944 , n24371 );
    or g7719 ( n27033 , n2248 , n32086 );
    xnor g7720 ( n35395 , n19516 , n34474 );
    or g7721 ( n15630 , n3977 , n19084 );
    xnor g7722 ( n24404 , n22335 , n19892 );
    xnor g7723 ( n24702 , n18029 , n31795 );
    or g7724 ( n9093 , n22291 , n6572 );
    xnor g7725 ( n10260 , n9612 , n2800 );
    nor g7726 ( n31391 , n30973 , n13261 );
    and g7727 ( n10064 , n30787 , n9434 );
    xnor g7728 ( n31620 , n22991 , n24371 );
    and g7729 ( n28011 , n19541 , n9931 );
    nor g7730 ( n27692 , n3205 , n13732 );
    and g7731 ( n1069 , n15583 , n609 );
    or g7732 ( n16130 , n18913 , n19939 );
    not g7733 ( n18095 , n16223 );
    xnor g7734 ( n27637 , n13683 , n9067 );
    or g7735 ( n2298 , n11157 , n29626 );
    or g7736 ( n25985 , n29839 , n28431 );
    xnor g7737 ( n16684 , n28860 , n21301 );
    and g7738 ( n24826 , n32755 , n18394 );
    or g7739 ( n29797 , n30648 , n1168 );
    or g7740 ( n27791 , n9351 , n19755 );
    and g7741 ( n22914 , n13450 , n9110 );
    or g7742 ( n2401 , n23195 , n5779 );
    or g7743 ( n3337 , n9789 , n15163 );
    or g7744 ( n13972 , n17288 , n1511 );
    or g7745 ( n16094 , n19883 , n35317 );
    and g7746 ( n10758 , n23353 , n71 );
    and g7747 ( n4684 , n2060 , n16653 );
    or g7748 ( n2173 , n21504 , n19448 );
    nor g7749 ( n33870 , n4701 , n32379 );
    or g7750 ( n31708 , n4878 , n19603 );
    and g7751 ( n11752 , n18590 , n3214 );
    or g7752 ( n25168 , n19984 , n1725 );
    and g7753 ( n866 , n22103 , n1532 );
    and g7754 ( n14308 , n4195 , n23267 );
    or g7755 ( n10282 , n18084 , n6553 );
    xnor g7756 ( n16398 , n30774 , n34440 );
    and g7757 ( n19593 , n10699 , n14830 );
    or g7758 ( n9927 , n10477 , n2585 );
    or g7759 ( n32207 , n15886 , n20511 );
    xnor g7760 ( n8156 , n8219 , n28103 );
    xnor g7761 ( n12137 , n30185 , n32584 );
    or g7762 ( n5882 , n11208 , n5457 );
    nor g7763 ( n14102 , n383 , n1480 );
    and g7764 ( n6447 , n13542 , n10347 );
    and g7765 ( n30362 , n13045 , n29011 );
    and g7766 ( n19604 , n10687 , n5672 );
    or g7767 ( n22454 , n5420 , n30519 );
    and g7768 ( n30238 , n18363 , n34259 );
    or g7769 ( n10172 , n28388 , n7215 );
    xnor g7770 ( n32864 , n4063 , n26 );
    not g7771 ( n9088 , n5287 );
    or g7772 ( n35231 , n25196 , n15090 );
    xnor g7773 ( n168 , n13501 , n16781 );
    and g7774 ( n8371 , n17443 , n1206 );
    and g7775 ( n8613 , n32184 , n2307 );
    xnor g7776 ( n22725 , n8365 , n4856 );
    nor g7777 ( n20670 , n31799 , n16114 );
    or g7778 ( n2615 , n13951 , n15667 );
    xnor g7779 ( n15665 , n15293 , n3659 );
    not g7780 ( n29594 , n31711 );
    xnor g7781 ( n9407 , n23940 , n22130 );
    or g7782 ( n16242 , n22730 , n6510 );
    xnor g7783 ( n32363 , n15142 , n9295 );
    or g7784 ( n10296 , n2263 , n29873 );
    or g7785 ( n18445 , n22132 , n10793 );
    or g7786 ( n8998 , n32857 , n31481 );
    or g7787 ( n15268 , n35927 , n4551 );
    or g7788 ( n22141 , n20838 , n22316 );
    and g7789 ( n3224 , n29634 , n19140 );
    not g7790 ( n28638 , n20689 );
    xnor g7791 ( n27457 , n30600 , n4878 );
    or g7792 ( n27425 , n8543 , n5752 );
    nor g7793 ( n9293 , n23102 , n29062 );
    or g7794 ( n30784 , n31289 , n10714 );
    xnor g7795 ( n9333 , n12696 , n12494 );
    not g7796 ( n6859 , n24081 );
    or g7797 ( n1112 , n23604 , n28143 );
    and g7798 ( n24955 , n20036 , n46 );
    not g7799 ( n31022 , n22677 );
    or g7800 ( n5268 , n22690 , n24356 );
    and g7801 ( n3508 , n709 , n13163 );
    not g7802 ( n9981 , n32584 );
    or g7803 ( n31795 , n32461 , n21753 );
    or g7804 ( n31369 , n9564 , n23707 );
    xnor g7805 ( n6299 , n19860 , n17568 );
    xnor g7806 ( n32587 , n29166 , n12392 );
    xnor g7807 ( n34987 , n3590 , n9999 );
    and g7808 ( n35494 , n18184 , n30294 );
    xnor g7809 ( n30962 , n469 , n3222 );
    not g7810 ( n1931 , n9208 );
    or g7811 ( n18079 , n33657 , n27997 );
    xnor g7812 ( n26501 , n21781 , n1663 );
    xnor g7813 ( n21796 , n2400 , n35766 );
    xnor g7814 ( n7616 , n14329 , n30813 );
    or g7815 ( n4068 , n25015 , n25306 );
    and g7816 ( n23442 , n22699 , n4341 );
    or g7817 ( n3948 , n12261 , n31004 );
    or g7818 ( n6245 , n3677 , n3756 );
    nor g7819 ( n33661 , n35437 , n28778 );
    xnor g7820 ( n34207 , n12969 , n1442 );
    buf g7821 ( n763 , n33368 );
    or g7822 ( n21473 , n31827 , n11295 );
    not g7823 ( n34342 , n2092 );
    and g7824 ( n11789 , n5829 , n18971 );
    xnor g7825 ( n10119 , n29661 , n1260 );
    or g7826 ( n17107 , n121 , n7726 );
    xnor g7827 ( n13333 , n20176 , n31289 );
    not g7828 ( n33017 , n2095 );
    and g7829 ( n18955 , n23477 , n34147 );
    or g7830 ( n19832 , n2646 , n19464 );
    not g7831 ( n19968 , n28273 );
    and g7832 ( n7931 , n34857 , n3293 );
    or g7833 ( n18545 , n7209 , n20601 );
    xnor g7834 ( n12524 , n33735 , n2757 );
    not g7835 ( n22819 , n10894 );
    and g7836 ( n24866 , n2722 , n24306 );
    or g7837 ( n979 , n15399 , n27268 );
    or g7838 ( n23799 , n32446 , n30708 );
    xnor g7839 ( n17851 , n36043 , n13950 );
    or g7840 ( n8976 , n8432 , n32284 );
    nor g7841 ( n35189 , n27662 , n29203 );
    or g7842 ( n31555 , n31225 , n268 );
    not g7843 ( n12538 , n12428 );
    or g7844 ( n13092 , n6359 , n19732 );
    xnor g7845 ( n33520 , n8662 , n15266 );
    or g7846 ( n6429 , n7316 , n5278 );
    xnor g7847 ( n23057 , n1296 , n7540 );
    or g7848 ( n18229 , n14623 , n2384 );
    or g7849 ( n24257 , n15886 , n11401 );
    buf g7850 ( n32634 , n544 );
    and g7851 ( n11225 , n30979 , n5744 );
    or g7852 ( n25169 , n17568 , n11709 );
    or g7853 ( n27119 , n7343 , n34084 );
    and g7854 ( n4542 , n31994 , n18708 );
    or g7855 ( n10250 , n1633 , n351 );
    or g7856 ( n2993 , n13796 , n35748 );
    xnor g7857 ( n27442 , n6297 , n21553 );
    and g7858 ( n6586 , n16333 , n29610 );
    xnor g7859 ( n3937 , n13528 , n31056 );
    xnor g7860 ( n1148 , n31899 , n10739 );
    or g7861 ( n1817 , n20880 , n6742 );
    or g7862 ( n11441 , n18743 , n20576 );
    nor g7863 ( n28615 , n9793 , n12544 );
    and g7864 ( n27720 , n13576 , n27780 );
    or g7865 ( n34820 , n5210 , n6618 );
    or g7866 ( n31941 , n5335 , n30670 );
    xnor g7867 ( n15426 , n10351 , n4240 );
    or g7868 ( n19638 , n21869 , n24489 );
    not g7869 ( n6965 , n25553 );
    and g7870 ( n28798 , n9677 , n29590 );
    nor g7871 ( n26908 , n3205 , n27385 );
    and g7872 ( n22570 , n35098 , n25305 );
    and g7873 ( n29926 , n11650 , n31341 );
    or g7874 ( n12589 , n22637 , n14918 );
    buf g7875 ( n1176 , n2436 );
    or g7876 ( n28793 , n35220 , n5457 );
    or g7877 ( n23223 , n31307 , n25831 );
    or g7878 ( n16374 , n24998 , n13788 );
    or g7879 ( n22230 , n21293 , n32572 );
    and g7880 ( n11048 , n6515 , n26570 );
    or g7881 ( n1469 , n23815 , n12596 );
    and g7882 ( n19113 , n28762 , n13079 );
    xnor g7883 ( n32187 , n32476 , n15464 );
    and g7884 ( n20399 , n374 , n3534 );
    or g7885 ( n16224 , n32715 , n34599 );
    or g7886 ( n29931 , n33066 , n23060 );
    xnor g7887 ( n1738 , n2248 , n15936 );
    not g7888 ( n20526 , n22980 );
    not g7889 ( n15075 , n33274 );
    or g7890 ( n10406 , n5172 , n10140 );
    not g7891 ( n24220 , n13463 );
    or g7892 ( n35805 , n19319 , n1942 );
    buf g7893 ( n30586 , n3396 );
    or g7894 ( n25890 , n34641 , n6913 );
    nor g7895 ( n24511 , n34959 , n19834 );
    xnor g7896 ( n19439 , n321 , n19387 );
    or g7897 ( n6808 , n13436 , n29516 );
    or g7898 ( n32165 , n4288 , n23315 );
    and g7899 ( n20832 , n24100 , n35198 );
    nor g7900 ( n62 , n14317 , n32324 );
    xnor g7901 ( n10286 , n28556 , n10246 );
    xnor g7902 ( n19489 , n16280 , n27257 );
    and g7903 ( n17436 , n11899 , n13655 );
    nor g7904 ( n13598 , n4878 , n11042 );
    or g7905 ( n8144 , n2561 , n27573 );
    not g7906 ( n13452 , n31289 );
    or g7907 ( n6228 , n16738 , n14918 );
    xnor g7908 ( n26566 , n15883 , n10216 );
    xnor g7909 ( n20699 , n9187 , n27759 );
    not g7910 ( n1849 , n34943 );
    or g7911 ( n15911 , n8468 , n33388 );
    or g7912 ( n30757 , n2512 , n33098 );
    xnor g7913 ( n3770 , n19837 , n10424 );
    and g7914 ( n32178 , n12633 , n4730 );
    not g7915 ( n18936 , n12622 );
    or g7916 ( n24205 , n15464 , n24528 );
    xnor g7917 ( n30599 , n32663 , n29769 );
    xnor g7918 ( n6699 , n33037 , n35720 );
    and g7919 ( n24061 , n29679 , n12997 );
    xnor g7920 ( n2048 , n9354 , n16648 );
    and g7921 ( n24450 , n12998 , n24391 );
    or g7922 ( n5845 , n1553 , n26292 );
    or g7923 ( n22976 , n15464 , n27657 );
    nor g7924 ( n7253 , n3186 , n12913 );
    and g7925 ( n20872 , n5433 , n17849 );
    xnor g7926 ( n10227 , n6684 , n4288 );
    and g7927 ( n32110 , n21458 , n33602 );
    and g7928 ( n19255 , n34125 , n15382 );
    or g7929 ( n29369 , n25313 , n1763 );
    and g7930 ( n23299 , n14895 , n375 );
    nor g7931 ( n2660 , n27738 , n9591 );
    or g7932 ( n32025 , n24098 , n31283 );
    or g7933 ( n4219 , n31899 , n10739 );
    or g7934 ( n25437 , n23106 , n12442 );
    and g7935 ( n10415 , n6770 , n14408 );
    and g7936 ( n3837 , n15491 , n34928 );
    or g7937 ( n6138 , n31289 , n24194 );
    or g7938 ( n10226 , n4878 , n20816 );
    not g7939 ( n8638 , n2487 );
    or g7940 ( n18352 , n29839 , n8481 );
    not g7941 ( n27245 , n22595 );
    and g7942 ( n4491 , n19592 , n33003 );
    and g7943 ( n35826 , n4114 , n20083 );
    and g7944 ( n12973 , n15751 , n7438 );
    and g7945 ( n4239 , n21812 , n3040 );
    or g7946 ( n2273 , n22590 , n15117 );
    and g7947 ( n858 , n12578 , n23261 );
    or g7948 ( n14815 , n5341 , n32330 );
    or g7949 ( n27034 , n32694 , n16961 );
    or g7950 ( n10912 , n12315 , n11833 );
    and g7951 ( n8476 , n8952 , n27913 );
    and g7952 ( n6753 , n19289 , n30120 );
    and g7953 ( n25015 , n6849 , n22481 );
    xnor g7954 ( n198 , n34358 , n21919 );
    or g7955 ( n21501 , n686 , n33757 );
    not g7956 ( n24051 , n9789 );
    not g7957 ( n14717 , n17539 );
    or g7958 ( n35675 , n10050 , n4508 );
    or g7959 ( n25004 , n3946 , n8881 );
    xnor g7960 ( n3076 , n28180 , n26974 );
    or g7961 ( n33281 , n21022 , n11977 );
    or g7962 ( n2259 , n19984 , n3981 );
    or g7963 ( n21573 , n21323 , n73 );
    or g7964 ( n31079 , n10798 , n7345 );
    or g7965 ( n14338 , n32584 , n22689 );
    or g7966 ( n7710 , n9568 , n24267 );
    xnor g7967 ( n8933 , n19975 , n19551 );
    or g7968 ( n15451 , n23681 , n1812 );
    or g7969 ( n35039 , n1799 , n16488 );
    not g7970 ( n21282 , n9789 );
    xnor g7971 ( n12819 , n6569 , n7540 );
    nor g7972 ( n14858 , n20526 , n21811 );
    xnor g7973 ( n10249 , n17474 , n24336 );
    and g7974 ( n35827 , n29233 , n27061 );
    xnor g7975 ( n1850 , n3162 , n22291 );
    not g7976 ( n7730 , n4769 );
    and g7977 ( n23847 , n5276 , n12814 );
    nor g7978 ( n17810 , n12264 , n11594 );
    xnor g7979 ( n9331 , n9510 , n12674 );
    or g7980 ( n33131 , n23604 , n4979 );
    not g7981 ( n23149 , n7588 );
    xnor g7982 ( n26098 , n6347 , n16135 );
    or g7983 ( n5288 , n17967 , n25133 );
    not g7984 ( n22245 , n5411 );
    or g7985 ( n25156 , n3707 , n23805 );
    or g7986 ( n5205 , n24898 , n6338 );
    xnor g7987 ( n6567 , n14639 , n8781 );
    or g7988 ( n23206 , n8467 , n12596 );
    or g7989 ( n33711 , n20848 , n217 );
    xnor g7990 ( n28984 , n11697 , n4818 );
    or g7991 ( n24495 , n12544 , n30708 );
    and g7992 ( n34273 , n26715 , n10608 );
    xnor g7993 ( n15325 , n35782 , n16017 );
    xnor g7994 ( n6495 , n3729 , n5738 );
    nor g7995 ( n15416 , n16319 , n24091 );
    buf g7996 ( n18542 , n12956 );
    and g7997 ( n17978 , n3159 , n30500 );
    or g7998 ( n13916 , n17505 , n29366 );
    or g7999 ( n11166 , n20489 , n27730 );
    not g8000 ( n26919 , n28969 );
    and g8001 ( n24592 , n30699 , n9339 );
    and g8002 ( n19976 , n4579 , n35406 );
    or g8003 ( n30155 , n15207 , n13991 );
    or g8004 ( n4144 , n33958 , n12791 );
    or g8005 ( n9423 , n5942 , n27929 );
    not g8006 ( n32186 , n2029 );
    or g8007 ( n35137 , n24371 , n21799 );
    or g8008 ( n34569 , n20434 , n15109 );
    buf g8009 ( n8090 , n11755 );
    and g8010 ( n20253 , n31221 , n33852 );
    or g8011 ( n17130 , n13769 , n3736 );
    xnor g8012 ( n31199 , n17345 , n7081 );
    xor g8013 ( n34186 , n17646 , n18279 );
    and g8014 ( n15310 , n19337 , n9939 );
    xnor g8015 ( n31900 , n2102 , n8218 );
    or g8016 ( n34141 , n17955 , n14076 );
    or g8017 ( n31279 , n28105 , n19952 );
    or g8018 ( n20978 , n29276 , n5168 );
    and g8019 ( n27283 , n2014 , n9701 );
    and g8020 ( n24168 , n15679 , n13989 );
    or g8021 ( n34698 , n15963 , n34298 );
    or g8022 ( n23409 , n20106 , n27866 );
    and g8023 ( n32569 , n26355 , n29809 );
    and g8024 ( n34447 , n10626 , n19202 );
    or g8025 ( n14932 , n14299 , n8392 );
    and g8026 ( n9190 , n8669 , n7134 );
    xnor g8027 ( n35776 , n21520 , n12294 );
    or g8028 ( n18011 , n14655 , n3736 );
    xnor g8029 ( n15528 , n26772 , n23605 );
    and g8030 ( n4664 , n4958 , n3182 );
    nor g8031 ( n20271 , n32393 , n26346 );
    or g8032 ( n22000 , n17946 , n15439 );
    or g8033 ( n10068 , n8431 , n8242 );
    not g8034 ( n5452 , n11195 );
    or g8035 ( n15367 , n35846 , n15383 );
    and g8036 ( n7221 , n17620 , n23555 );
    nor g8037 ( n16153 , n19348 , n18264 );
    xnor g8038 ( n5841 , n34694 , n995 );
    or g8039 ( n28763 , n2376 , n31549 );
    or g8040 ( n15440 , n28924 , n6266 );
    not g8041 ( n8755 , n33786 );
    or g8042 ( n28817 , n15190 , n21977 );
    xnor g8043 ( n25665 , n8481 , n29839 );
    or g8044 ( n23563 , n14366 , n22946 );
    or g8045 ( n12997 , n22291 , n320 );
    nor g8046 ( n10058 , n3205 , n3584 );
    or g8047 ( n21050 , n918 , n28064 );
    or g8048 ( n17870 , n35123 , n24860 );
    not g8049 ( n21097 , n4962 );
    and g8050 ( n22590 , n4658 , n12812 );
    not g8051 ( n18652 , n6205 );
    or g8052 ( n18939 , n8435 , n5868 );
    not g8053 ( n22861 , n18438 );
    xnor g8054 ( n18293 , n4553 , n31388 );
    or g8055 ( n20491 , n11300 , n27631 );
    and g8056 ( n13862 , n35905 , n5934 );
    xnor g8057 ( n20565 , n12142 , n29839 );
    and g8058 ( n35947 , n28886 , n30598 );
    or g8059 ( n5269 , n23361 , n29535 );
    not g8060 ( n16296 , n4791 );
    not g8061 ( n21602 , n31233 );
    not g8062 ( n24635 , n30732 );
    or g8063 ( n14086 , n5512 , n22707 );
    xnor g8064 ( n28774 , n34278 , n205 );
    or g8065 ( n4094 , n9793 , n19750 );
    or g8066 ( n28068 , n25602 , n15298 );
    and g8067 ( n32338 , n19658 , n30474 );
    and g8068 ( n9827 , n32862 , n14711 );
    not g8069 ( n15942 , n7540 );
    not g8070 ( n17480 , n14766 );
    xnor g8071 ( n32050 , n8634 , n33680 );
    xnor g8072 ( n17897 , n34044 , n27355 );
    or g8073 ( n11792 , n7355 , n25567 );
    and g8074 ( n8437 , n15080 , n33252 );
    and g8075 ( n32220 , n24575 , n20581 );
    xnor g8076 ( n2192 , n313 , n30742 );
    or g8077 ( n25593 , n13209 , n28136 );
    nor g8078 ( n8737 , n16620 , n18594 );
    xnor g8079 ( n28107 , n18927 , n30742 );
    not g8080 ( n34458 , n30292 );
    or g8081 ( n13432 , n696 , n24696 );
    and g8082 ( n10197 , n15400 , n24612 );
    or g8083 ( n5768 , n17099 , n5752 );
    and g8084 ( n11702 , n10795 , n312 );
    xnor g8085 ( n9682 , n33868 , n1350 );
    nor g8086 ( n6866 , n8432 , n15800 );
    or g8087 ( n29424 , n28340 , n26517 );
    and g8088 ( n24549 , n15428 , n21259 );
    not g8089 ( n10976 , n10405 );
    nor g8090 ( n15070 , n21635 , n3763 );
    or g8091 ( n17217 , n1500 , n31606 );
    or g8092 ( n2958 , n24280 , n5924 );
    or g8093 ( n7843 , n31191 , n31514 );
    nor g8094 ( n11894 , n17568 , n683 );
    or g8095 ( n26511 , n11155 , n13459 );
    and g8096 ( n11401 , n14173 , n6445 );
    or g8097 ( n4787 , n15021 , n20584 );
    nor g8098 ( n5184 , n7814 , n22628 );
    xnor g8099 ( n4765 , n15340 , n21803 );
    or g8100 ( n303 , n19474 , n16934 );
    or g8101 ( n159 , n25463 , n35748 );
    or g8102 ( n14909 , n26464 , n20579 );
    or g8103 ( n32903 , n24371 , n12845 );
    and g8104 ( n11575 , n27681 , n13852 );
    nor g8105 ( n33935 , n3222 , n449 );
    xnor g8106 ( n23704 , n30546 , n16423 );
    and g8107 ( n36007 , n7333 , n35065 );
    or g8108 ( n8760 , n31929 , n35978 );
    and g8109 ( n25107 , n20630 , n32132 );
    and g8110 ( n30036 , n35044 , n9438 );
    or g8111 ( n18505 , n31651 , n10336 );
    and g8112 ( n15657 , n13092 , n27299 );
    and g8113 ( n9513 , n32540 , n7206 );
    xnor g8114 ( n6136 , n26353 , n15994 );
    or g8115 ( n29308 , n19333 , n26365 );
    or g8116 ( n33587 , n30742 , n33099 );
    or g8117 ( n29472 , n13557 , n30732 );
    not g8118 ( n21760 , n22200 );
    and g8119 ( n26612 , n13687 , n10753 );
    and g8120 ( n27985 , n28353 , n3980 );
    xnor g8121 ( n35088 , n13956 , n35927 );
    xnor g8122 ( n12382 , n31324 , n23128 );
    and g8123 ( n30832 , n24169 , n14176 );
    and g8124 ( n15055 , n21185 , n11210 );
    or g8125 ( n1138 , n10519 , n14618 );
    or g8126 ( n12418 , n1950 , n34356 );
    and g8127 ( n320 , n5192 , n34006 );
    or g8128 ( n17269 , n33038 , n19490 );
    and g8129 ( n15498 , n15127 , n31935 );
    not g8130 ( n26341 , n8087 );
    and g8131 ( n10082 , n27334 , n9526 );
    and g8132 ( n8450 , n20890 , n12240 );
    and g8133 ( n29983 , n6555 , n33926 );
    nor g8134 ( n3657 , n17568 , n29306 );
    not g8135 ( n24719 , n28438 );
    or g8136 ( n23719 , n3195 , n19244 );
    or g8137 ( n15950 , n30553 , n12550 );
    not g8138 ( n17008 , n8123 );
    or g8139 ( n3262 , n23547 , n25424 );
    or g8140 ( n17596 , n28684 , n25392 );
    or g8141 ( n4232 , n26977 , n23882 );
    and g8142 ( n15422 , n26557 , n24409 );
    xnor g8143 ( n2555 , n26758 , n18968 );
    nor g8144 ( n13896 , n16620 , n20057 );
    or g8145 ( n33584 , n16672 , n18007 );
    and g8146 ( n33969 , n28505 , n3781 );
    nor g8147 ( n27180 , n32857 , n11802 );
    or g8148 ( n2223 , n16663 , n7312 );
    and g8149 ( n19283 , n23317 , n20896 );
    xnor g8150 ( n34073 , n3078 , n9241 );
    or g8151 ( n21667 , n27637 , n17964 );
    and g8152 ( n22257 , n26439 , n510 );
    xnor g8153 ( n12278 , n20682 , n24538 );
    nor g8154 ( n19351 , n23630 , n25390 );
    or g8155 ( n22800 , n28906 , n33956 );
    nor g8156 ( n3809 , n29713 , n284 );
    or g8157 ( n29415 , n35927 , n6780 );
    or g8158 ( n25356 , n28701 , n24696 );
    not g8159 ( n20716 , n2395 );
    and g8160 ( n25312 , n15430 , n15391 );
    or g8161 ( n5639 , n1821 , n35422 );
    xnor g8162 ( n15149 , n34796 , n22294 );
    or g8163 ( n14518 , n24371 , n16583 );
    xnor g8164 ( n34294 , n21834 , n29544 );
    xnor g8165 ( n21460 , n5937 , n18379 );
    or g8166 ( n14534 , n26944 , n15805 );
    and g8167 ( n22574 , n27296 , n18069 );
    not g8168 ( n2340 , n27437 );
    or g8169 ( n1291 , n20832 , n21644 );
    not g8170 ( n35209 , n14126 );
    and g8171 ( n18921 , n5632 , n18284 );
    and g8172 ( n19145 , n25885 , n21377 );
    or g8173 ( n6545 , n32095 , n33652 );
    xnor g8174 ( n36023 , n34085 , n6966 );
    or g8175 ( n34823 , n9793 , n28163 );
    or g8176 ( n32200 , n27291 , n22353 );
    xnor g8177 ( n33280 , n4377 , n30742 );
    or g8178 ( n31459 , n31591 , n28702 );
    and g8179 ( n33515 , n34803 , n17263 );
    and g8180 ( n28318 , n7520 , n5383 );
    and g8181 ( n33285 , n1536 , n504 );
    buf g8182 ( n4318 , n21853 );
    or g8183 ( n22329 , n31580 , n10960 );
    or g8184 ( n25212 , n16825 , n6950 );
    xnor g8185 ( n17647 , n15305 , n3946 );
    nor g8186 ( n10892 , n30873 , n9921 );
    or g8187 ( n11753 , n29064 , n16462 );
    and g8188 ( n23205 , n16871 , n4944 );
    or g8189 ( n12523 , n14981 , n21307 );
    xnor g8190 ( n9465 , n7572 , n29205 );
    xnor g8191 ( n2628 , n23594 , n9793 );
    buf g8192 ( n2168 , n33590 );
    or g8193 ( n1713 , n26519 , n15714 );
    or g8194 ( n23437 , n9432 , n31780 );
    or g8195 ( n24125 , n16616 , n24025 );
    or g8196 ( n6916 , n6452 , n25712 );
    and g8197 ( n1909 , n27475 , n15276 );
    buf g8198 ( n9832 , n9731 );
    xnor g8199 ( n14921 , n10636 , n33642 );
    or g8200 ( n22609 , n6559 , n20797 );
    nor g8201 ( n24499 , n33166 , n9811 );
    and g8202 ( n4744 , n30875 , n29313 );
    and g8203 ( n4058 , n13571 , n32734 );
    xnor g8204 ( n19586 , n36080 , n1132 );
    xnor g8205 ( n7932 , n9697 , n21899 );
    or g8206 ( n22912 , n26335 , n25567 );
    or g8207 ( n29447 , n29000 , n31794 );
    and g8208 ( n19071 , n30887 , n10202 );
    and g8209 ( n5122 , n35807 , n28377 );
    or g8210 ( n10095 , n18379 , n14785 );
    xnor g8211 ( n30115 , n17433 , n29323 );
    or g8212 ( n200 , n16832 , n4172 );
    and g8213 ( n30462 , n33508 , n14539 );
    or g8214 ( n16128 , n25948 , n31773 );
    and g8215 ( n707 , n16587 , n9245 );
    or g8216 ( n3883 , n31954 , n26468 );
    xnor g8217 ( n8852 , n14510 , n14580 );
    or g8218 ( n22411 , n17750 , n23209 );
    xnor g8219 ( n14982 , n12683 , n10894 );
    or g8220 ( n35685 , n31153 , n2600 );
    not g8221 ( n33144 , n32451 );
    not g8222 ( n25193 , n18003 );
    and g8223 ( n30600 , n34055 , n23837 );
    xnor g8224 ( n4212 , n21371 , n33910 );
    xnor g8225 ( n5803 , n29030 , n4397 );
    nor g8226 ( n10094 , n9414 , n27091 );
    xnor g8227 ( n17332 , n10620 , n3946 );
    and g8228 ( n11852 , n25741 , n9170 );
    nor g8229 ( n31200 , n21224 , n32720 );
    not g8230 ( n1946 , n28124 );
    or g8231 ( n12846 , n30742 , n22791 );
    and g8232 ( n19617 , n30408 , n31383 );
    or g8233 ( n18227 , n6373 , n3647 );
    nor g8234 ( n30517 , n4962 , n11683 );
    not g8235 ( n35174 , n32002 );
    and g8236 ( n16294 , n2930 , n4139 );
    or g8237 ( n25601 , n34057 , n17964 );
    not g8238 ( n27351 , n33744 );
    or g8239 ( n9364 , n31289 , n16479 );
    or g8240 ( n15472 , n13274 , n18878 );
    or g8241 ( n2740 , n4962 , n8277 );
    or g8242 ( n5217 , n11190 , n1890 );
    or g8243 ( n31103 , n16347 , n27728 );
    not g8244 ( n2585 , n5674 );
    not g8245 ( n89 , n4143 );
    or g8246 ( n4227 , n24508 , n11238 );
    xnor g8247 ( n28851 , n27370 , n29713 );
    or g8248 ( n26542 , n2786 , n14745 );
    or g8249 ( n32117 , n4962 , n33454 );
    xnor g8250 ( n8940 , n4987 , n28311 );
    and g8251 ( n24035 , n3441 , n13025 );
    xnor g8252 ( n15483 , n9768 , n23219 );
    xnor g8253 ( n27107 , n6512 , n19551 );
    or g8254 ( n12916 , n24285 , n24622 );
    xnor g8255 ( n30729 , n23092 , n16837 );
    nor g8256 ( n17790 , n12636 , n34556 );
    not g8257 ( n5713 , n22793 );
    or g8258 ( n32100 , n25977 , n31134 );
    xnor g8259 ( n14421 , n1421 , n8432 );
    xnor g8260 ( n22282 , n6241 , n17317 );
    xnor g8261 ( n1269 , n16026 , n19442 );
    and g8262 ( n9121 , n4462 , n20119 );
    or g8263 ( n25042 , n19880 , n33593 );
    or g8264 ( n7247 , n7000 , n4635 );
    and g8265 ( n32719 , n18459 , n3062 );
    or g8266 ( n3336 , n28278 , n12428 );
    xnor g8267 ( n5886 , n17747 , n3215 );
    xnor g8268 ( n7597 , n14350 , n30742 );
    not g8269 ( n35046 , n8977 );
    xnor g8270 ( n2907 , n32981 , n17568 );
    xnor g8271 ( n16481 , n14631 , n35657 );
    not g8272 ( n16468 , n35291 );
    xnor g8273 ( n15454 , n22524 , n30674 );
    nor g8274 ( n9615 , n25602 , n7005 );
    or g8275 ( n227 , n23644 , n26023 );
    or g8276 ( n14453 , n5678 , n16152 );
    or g8277 ( n33263 , n3063 , n21077 );
    and g8278 ( n25043 , n18447 , n32845 );
    or g8279 ( n19165 , n24371 , n17395 );
    or g8280 ( n18376 , n24897 , n1642 );
    nor g8281 ( n2098 , n24865 , n3550 );
    xnor g8282 ( n26314 , n7811 , n15004 );
    or g8283 ( n8033 , n10647 , n12950 );
    and g8284 ( n22301 , n30691 , n13251 );
    xnor g8285 ( n25698 , n7316 , n5278 );
    and g8286 ( n33683 , n1095 , n757 );
    or g8287 ( n16120 , n32127 , n20066 );
    and g8288 ( n18047 , n32564 , n11107 );
    or g8289 ( n12190 , n1999 , n14746 );
    or g8290 ( n16568 , n23150 , n11418 );
    or g8291 ( n1661 , n30046 , n29953 );
    not g8292 ( n1603 , n22471 );
    xnor g8293 ( n34439 , n22798 , n6279 );
    xnor g8294 ( n21729 , n4004 , n23627 );
    or g8295 ( n29682 , n10894 , n9387 );
    and g8296 ( n2986 , n1315 , n20754 );
    or g8297 ( n19775 , n846 , n5150 );
    or g8298 ( n25190 , n34527 , n25831 );
    or g8299 ( n2292 , n13666 , n9648 );
    or g8300 ( n29347 , n23721 , n26686 );
    nor g8301 ( n28895 , n7690 , n13426 );
    and g8302 ( n19519 , n27285 , n5018 );
    and g8303 ( n22091 , n8968 , n34228 );
    buf g8304 ( n12879 , n30732 );
    xnor g8305 ( n28110 , n17278 , n29134 );
    or g8306 ( n3039 , n9509 , n29411 );
    or g8307 ( n3910 , n15978 , n20817 );
    or g8308 ( n14881 , n35980 , n31175 );
    xnor g8309 ( n6072 , n9850 , n23604 );
    or g8310 ( n32282 , n19606 , n5168 );
    not g8311 ( n30773 , n14045 );
    nor g8312 ( n10615 , n22291 , n23269 );
    and g8313 ( n23566 , n10520 , n18213 );
    or g8314 ( n14598 , n11110 , n585 );
    or g8315 ( n14455 , n28465 , n21956 );
    xnor g8316 ( n17186 , n29882 , n35927 );
    not g8317 ( n16307 , n22291 );
    or g8318 ( n11386 , n34448 , n15980 );
    xnor g8319 ( n2169 , n5379 , n8495 );
    or g8320 ( n15664 , n24531 , n7726 );
    xnor g8321 ( n1877 , n26753 , n25714 );
    and g8322 ( n1576 , n25566 , n1798 );
    xnor g8323 ( n4091 , n17274 , n25630 );
    or g8324 ( n31714 , n20115 , n19475 );
    nor g8325 ( n13782 , n16996 , n11826 );
    or g8326 ( n34402 , n6451 , n20690 );
    and g8327 ( n22013 , n11457 , n6228 );
    or g8328 ( n16721 , n12704 , n25648 );
    and g8329 ( n14566 , n7729 , n8222 );
    and g8330 ( n941 , n21020 , n27848 );
    and g8331 ( n27682 , n21233 , n32686 );
    and g8332 ( n14196 , n10373 , n3924 );
    nor g8333 ( n27041 , n13396 , n6406 );
    or g8334 ( n795 , n21603 , n16961 );
    or g8335 ( n14480 , n14792 , n21747 );
    or g8336 ( n5814 , n23621 , n8253 );
    xnor g8337 ( n14712 , n29975 , n19551 );
    nor g8338 ( n2164 , n31289 , n10134 );
    and g8339 ( n14677 , n15324 , n1841 );
    xnor g8340 ( n29348 , n25988 , n9812 );
    or g8341 ( n18541 , n15163 , n24025 );
    or g8342 ( n15410 , n9048 , n12457 );
    or g8343 ( n30996 , n20574 , n17068 );
    or g8344 ( n22220 , n23676 , n1414 );
    xnor g8345 ( n1819 , n3093 , n11455 );
    xnor g8346 ( n26944 , n30938 , n21056 );
    xnor g8347 ( n2379 , n1852 , n9793 );
    and g8348 ( n35202 , n35662 , n159 );
    and g8349 ( n18878 , n24680 , n27981 );
    xnor g8350 ( n23487 , n24834 , n17711 );
    xnor g8351 ( n24327 , n6173 , n26402 );
    and g8352 ( n21870 , n10120 , n1876 );
    xnor g8353 ( n17912 , n31332 , n13021 );
    xnor g8354 ( n13879 , n15108 , n14637 );
    nor g8355 ( n13522 , n9793 , n29782 );
    or g8356 ( n18898 , n10318 , n32806 );
    or g8357 ( n18961 , n16755 , n22024 );
    xnor g8358 ( n20682 , n9265 , n9793 );
    xnor g8359 ( n31802 , n24963 , n32715 );
    or g8360 ( n14457 , n23694 , n29502 );
    not g8361 ( n5216 , n6815 );
    or g8362 ( n13171 , n4881 , n17046 );
    or g8363 ( n4518 , n16135 , n5644 );
    not g8364 ( n2313 , n6363 );
    or g8365 ( n19806 , n26568 , n13900 );
    or g8366 ( n29213 , n4962 , n9140 );
    nor g8367 ( n6020 , n10930 , n4508 );
    xnor g8368 ( n7098 , n9901 , n30127 );
    nor g8369 ( n19180 , n21602 , n289 );
    or g8370 ( n15668 , n1787 , n9504 );
    xnor g8371 ( n16051 , n25058 , n17227 );
    or g8372 ( n2202 , n19924 , n7869 );
    or g8373 ( n11986 , n16805 , n32842 );
    xnor g8374 ( n24896 , n16735 , n22016 );
    and g8375 ( n12093 , n26491 , n25225 );
    and g8376 ( n32441 , n23416 , n32117 );
    or g8377 ( n1875 , n25602 , n29603 );
    or g8378 ( n12788 , n32092 , n6018 );
    or g8379 ( n31246 , n5250 , n2005 );
    xnor g8380 ( n11110 , n15587 , n21110 );
    or g8381 ( n728 , n409 , n19336 );
    not g8382 ( n13691 , n6252 );
    or g8383 ( n16413 , n26477 , n9747 );
    and g8384 ( n4178 , n19503 , n25846 );
    and g8385 ( n8903 , n12292 , n18241 );
    and g8386 ( n35660 , n7556 , n24396 );
    or g8387 ( n11270 , n19506 , n31627 );
    and g8388 ( n35663 , n27019 , n23371 );
    xnor g8389 ( n17156 , n21397 , n26921 );
    not g8390 ( n22909 , n30652 );
    xnor g8391 ( n9269 , n7880 , n25705 );
    nor g8392 ( n9562 , n12399 , n17582 );
    not g8393 ( n14748 , n8637 );
    xnor g8394 ( n5382 , n9881 , n14106 );
    and g8395 ( n11644 , n6946 , n16983 );
    or g8396 ( n21720 , n33822 , n5976 );
    or g8397 ( n18940 , n10093 , n10762 );
    not g8398 ( n18654 , n18296 );
    nor g8399 ( n5461 , n33041 , n35894 );
    xnor g8400 ( n22182 , n23608 , n9658 );
    or g8401 ( n29772 , n22569 , n33435 );
    xnor g8402 ( n3066 , n21863 , n1606 );
    or g8403 ( n19018 , n1344 , n15262 );
    or g8404 ( n12411 , n10249 , n27580 );
    or g8405 ( n34020 , n32840 , n35604 );
    xnor g8406 ( n12253 , n14571 , n7698 );
    or g8407 ( n7194 , n10894 , n33189 );
    nor g8408 ( n317 , n13947 , n1067 );
    or g8409 ( n24059 , n9191 , n32808 );
    and g8410 ( n14315 , n2789 , n33089 );
    or g8411 ( n9329 , n9658 , n5960 );
    or g8412 ( n20210 , n14287 , n11711 );
    xnor g8413 ( n18744 , n20926 , n28453 );
    or g8414 ( n1160 , n35312 , n1919 );
    xnor g8415 ( n21168 , n32627 , n19753 );
    and g8416 ( n19530 , n15140 , n11847 );
    or g8417 ( n15618 , n5739 , n10901 );
    and g8418 ( n5533 , n25433 , n18929 );
    or g8419 ( n3306 , n2933 , n29065 );
    xnor g8420 ( n25425 , n19478 , n25174 );
    or g8421 ( n12600 , n2133 , n11613 );
    or g8422 ( n8021 , n741 , n17046 );
    xnor g8423 ( n10716 , n17339 , n1950 );
    or g8424 ( n28916 , n1118 , n26818 );
    and g8425 ( n11995 , n9159 , n7841 );
    xnor g8426 ( n31981 , n20698 , n13724 );
    or g8427 ( n8590 , n28307 , n9782 );
    xnor g8428 ( n20924 , n20293 , n33338 );
    or g8429 ( n11370 , n6100 , n4645 );
    xnor g8430 ( n28224 , n7853 , n17568 );
    nor g8431 ( n15869 , n16620 , n12318 );
    nor g8432 ( n23713 , n12140 , n6017 );
    or g8433 ( n6600 , n34999 , n27447 );
    and g8434 ( n28489 , n18637 , n19916 );
    and g8435 ( n12377 , n6840 , n1908 );
    xnor g8436 ( n27260 , n21424 , n13074 );
    xnor g8437 ( n18244 , n29338 , n29368 );
    not g8438 ( n19322 , n30589 );
    not g8439 ( n25023 , n20840 );
    and g8440 ( n17082 , n16601 , n4633 );
    or g8441 ( n35405 , n15926 , n17308 );
    and g8442 ( n15813 , n33045 , n24876 );
    and g8443 ( n12384 , n3492 , n22980 );
    and g8444 ( n12653 , n3697 , n10337 );
    or g8445 ( n6450 , n10034 , n25594 );
    and g8446 ( n21621 , n18998 , n5391 );
    and g8447 ( n21261 , n6345 , n5775 );
    or g8448 ( n678 , n4765 , n28668 );
    xnor g8449 ( n19615 , n5345 , n16620 );
    and g8450 ( n24950 , n8048 , n6768 );
    or g8451 ( n34703 , n12944 , n9194 );
    nor g8452 ( n15253 , n1950 , n17907 );
    or g8453 ( n14172 , n11190 , n3751 );
    or g8454 ( n16011 , n16508 , n8871 );
    or g8455 ( n35223 , n14256 , n31572 );
    or g8456 ( n28611 , n4921 , n4172 );
    or g8457 ( n22642 , n34538 , n8924 );
    nor g8458 ( n33178 , n4288 , n30715 );
    and g8459 ( n15768 , n33800 , n32062 );
    xnor g8460 ( n34005 , n33997 , n19313 );
    or g8461 ( n12193 , n7563 , n25447 );
    or g8462 ( n24960 , n11253 , n26360 );
    or g8463 ( n6659 , n3097 , n1090 );
    and g8464 ( n13320 , n29039 , n5241 );
    or g8465 ( n16267 , n32160 , n25255 );
    or g8466 ( n5407 , n19106 , n6678 );
    xnor g8467 ( n30764 , n17091 , n15073 );
    nor g8468 ( n12047 , n1950 , n7242 );
    buf g8469 ( n25773 , n2979 );
    and g8470 ( n22356 , n5251 , n15600 );
    xnor g8471 ( n3623 , n15874 , n5335 );
    and g8472 ( n33311 , n6385 , n17212 );
    and g8473 ( n26039 , n2772 , n30750 );
    or g8474 ( n6166 , n7204 , n4564 );
    or g8475 ( n3035 , n24700 , n18857 );
    not g8476 ( n31071 , n17685 );
    xnor g8477 ( n27521 , n32361 , n4960 );
    xnor g8478 ( n5392 , n11330 , n33036 );
    and g8479 ( n11010 , n16454 , n2180 );
    or g8480 ( n1501 , n27291 , n33460 );
    or g8481 ( n31145 , n348 , n34484 );
    or g8482 ( n20153 , n16950 , n1474 );
    or g8483 ( n17225 , n32857 , n30957 );
    xnor g8484 ( n24999 , n10255 , n26682 );
    nor g8485 ( n21931 , n7480 , n25185 );
    nor g8486 ( n6082 , n3909 , n7706 );
    xnor g8487 ( n33941 , n16265 , n15172 );
    xnor g8488 ( n16049 , n19148 , n35516 );
    nor g8489 ( n14428 , n1950 , n34350 );
    nor g8490 ( n11348 , n3205 , n21121 );
    and g8491 ( n1980 , n27415 , n6453 );
    nor g8492 ( n7051 , n5335 , n6973 );
    xnor g8493 ( n16793 , n11683 , n16175 );
    xnor g8494 ( n28443 , n23311 , n34249 );
    xnor g8495 ( n16833 , n33945 , n31577 );
    and g8496 ( n24676 , n27781 , n25134 );
    or g8497 ( n3993 , n27992 , n8071 );
    and g8498 ( n33257 , n15741 , n17823 );
    or g8499 ( n35338 , n21112 , n17962 );
    and g8500 ( n5163 , n22744 , n19224 );
    xnor g8501 ( n18073 , n10734 , n18437 );
    xnor g8502 ( n31077 , n15263 , n4758 );
    or g8503 ( n27014 , n2674 , n23414 );
    or g8504 ( n7970 , n32478 , n33158 );
    or g8505 ( n2012 , n31523 , n13215 );
    nor g8506 ( n6689 , n18742 , n15896 );
    not g8507 ( n24394 , n9789 );
    xnor g8508 ( n12836 , n8931 , n10593 );
    or g8509 ( n10295 , n12006 , n6340 );
    xnor g8510 ( n23985 , n26201 , n17870 );
    and g8511 ( n32736 , n5003 , n29070 );
    nor g8512 ( n14558 , n5344 , n6017 );
    nor g8513 ( n11879 , n17568 , n26177 );
    or g8514 ( n11199 , n24371 , n17249 );
    and g8515 ( n23201 , n24475 , n35263 );
    or g8516 ( n33363 , n25174 , n35327 );
    xnor g8517 ( n26250 , n213 , n15390 );
    or g8518 ( n24143 , n8753 , n1090 );
    xnor g8519 ( n27622 , n25609 , n20773 );
    xnor g8520 ( n15587 , n2387 , n19090 );
    or g8521 ( n33478 , n10894 , n3652 );
    or g8522 ( n6252 , n27489 , n11969 );
    and g8523 ( n28406 , n13888 , n32394 );
    or g8524 ( n9613 , n4010 , n11354 );
    xnor g8525 ( n32827 , n15617 , n9072 );
    nor g8526 ( n8617 , n2544 , n50 );
    xnor g8527 ( n9094 , n23850 , n4288 );
    xnor g8528 ( n12904 , n3236 , n29408 );
    and g8529 ( n27086 , n22016 , n16735 );
    and g8530 ( n15179 , n30629 , n29224 );
    or g8531 ( n1101 , n31406 , n4478 );
    nor g8532 ( n22990 , n19565 , n6017 );
    xnor g8533 ( n30343 , n14259 , n31277 );
    or g8534 ( n21697 , n27585 , n7965 );
    xnor g8535 ( n30073 , n31027 , n22916 );
    or g8536 ( n33849 , n22291 , n18403 );
    or g8537 ( n28487 , n4962 , n30114 );
    xnor g8538 ( n27422 , n32275 , n15707 );
    and g8539 ( n8871 , n19674 , n13954 );
    nor g8540 ( n5610 , n29149 , n23149 );
    xnor g8541 ( n31090 , n5564 , n6711 );
    or g8542 ( n20119 , n32715 , n5376 );
    or g8543 ( n34863 , n29859 , n6537 );
    or g8544 ( n1640 , n33633 , n9675 );
    or g8545 ( n5438 , n16156 , n11922 );
    or g8546 ( n17979 , n18463 , n585 );
    xnor g8547 ( n32796 , n19880 , n33593 );
    xnor g8548 ( n8717 , n27164 , n8432 );
    or g8549 ( n2004 , n377 , n11850 );
    not g8550 ( n24816 , n11929 );
    or g8551 ( n10757 , n16880 , n23532 );
    or g8552 ( n34686 , n18706 , n28574 );
    and g8553 ( n8337 , n34996 , n34789 );
    and g8554 ( n4271 , n21086 , n15212 );
    or g8555 ( n14151 , n32715 , n13149 );
    xnor g8556 ( n25094 , n9524 , n24758 );
    or g8557 ( n17821 , n4050 , n34865 );
    or g8558 ( n25726 , n23604 , n6796 );
    xnor g8559 ( n30498 , n1591 , n15464 );
    and g8560 ( n35238 , n3163 , n29720 );
    or g8561 ( n33213 , n16438 , n8108 );
    xnor g8562 ( n6830 , n11509 , n2492 );
    or g8563 ( n26807 , n11391 , n33310 );
    or g8564 ( n2916 , n13133 , n10872 );
    and g8565 ( n29232 , n21500 , n30240 );
    xnor g8566 ( n8334 , n12586 , n27226 );
    and g8567 ( n9163 , n19746 , n7830 );
    or g8568 ( n34206 , n16834 , n24356 );
    not g8569 ( n22841 , n17568 );
    xnor g8570 ( n7691 , n33446 , n6546 );
    or g8571 ( n28745 , n674 , n35141 );
    or g8572 ( n20480 , n9658 , n34359 );
    and g8573 ( n25397 , n4770 , n12610 );
    or g8574 ( n20151 , n8608 , n10762 );
    xnor g8575 ( n11268 , n8994 , n19288 );
    xnor g8576 ( n13802 , n6753 , n4288 );
    or g8577 ( n30627 , n11824 , n17302 );
    and g8578 ( n5978 , n8652 , n5824 );
    and g8579 ( n32682 , n18777 , n30609 );
    or g8580 ( n25308 , n32531 , n31554 );
    and g8581 ( n9529 , n18898 , n32470 );
    and g8582 ( n12112 , n10172 , n11836 );
    and g8583 ( n1413 , n11441 , n5352 );
    xnor g8584 ( n2034 , n668 , n3205 );
    xnor g8585 ( n17404 , n31617 , n31289 );
    buf g8586 ( n1474 , n20140 );
    not g8587 ( n15073 , n16620 );
    or g8588 ( n18292 , n17800 , n16919 );
    or g8589 ( n4867 , n31219 , n19105 );
    and g8590 ( n16073 , n2049 , n10344 );
    xnor g8591 ( n5872 , n13315 , n17568 );
    or g8592 ( n10390 , n12796 , n14070 );
    or g8593 ( n2183 , n10894 , n12683 );
    or g8594 ( n30060 , n19379 , n11866 );
    xnor g8595 ( n23661 , n3468 , n28422 );
    or g8596 ( n273 , n26763 , n7673 );
    xnor g8597 ( n9139 , n32879 , n19989 );
    or g8598 ( n26144 , n29670 , n1856 );
    or g8599 ( n14417 , n17568 , n33701 );
    or g8600 ( n10069 , n8486 , n10417 );
    xnor g8601 ( n8708 , n34955 , n32095 );
    or g8602 ( n28382 , n3506 , n14554 );
    xnor g8603 ( n28651 , n12091 , n18045 );
    xnor g8604 ( n10532 , n16641 , n11046 );
    or g8605 ( n27311 , n15641 , n26737 );
    and g8606 ( n26627 , n28483 , n21960 );
    and g8607 ( n32504 , n18170 , n25128 );
    nor g8608 ( n34298 , n3222 , n24009 );
    not g8609 ( n9798 , n17071 );
    or g8610 ( n34003 , n23037 , n25191 );
    xnor g8611 ( n6710 , n2735 , n3946 );
    not g8612 ( n2331 , n14068 );
    or g8613 ( n24788 , n10516 , n14691 );
    xnor g8614 ( n34364 , n35789 , n24371 );
    not g8615 ( n21801 , n5453 );
    and g8616 ( n284 , n23283 , n7854 );
    and g8617 ( n24243 , n15794 , n2115 );
    or g8618 ( n663 , n30073 , n18811 );
    xnor g8619 ( n9049 , n35788 , n3843 );
    or g8620 ( n5386 , n12090 , n25761 );
    and g8621 ( n32157 , n896 , n29511 );
    not g8622 ( n25415 , n22980 );
    and g8623 ( n31284 , n20843 , n33975 );
    xnor g8624 ( n8982 , n2024 , n15464 );
    or g8625 ( n5532 , n32498 , n16824 );
    xnor g8626 ( n15832 , n19874 , n4962 );
    not g8627 ( n31731 , n13243 );
    nor g8628 ( n30489 , n18849 , n3312 );
    and g8629 ( n25541 , n15362 , n7493 );
    and g8630 ( n22227 , n32298 , n24752 );
    or g8631 ( n10278 , n22782 , n24148 );
    or g8632 ( n22459 , n9793 , n13971 );
    and g8633 ( n669 , n5563 , n9755 );
    or g8634 ( n24802 , n25602 , n3780 );
    and g8635 ( n2342 , n29532 , n5212 );
    or g8636 ( n24938 , n11604 , n28799 );
    buf g8637 ( n9555 , n1796 );
    nor g8638 ( n25662 , n15299 , n18567 );
    xnor g8639 ( n30471 , n16000 , n5335 );
    or g8640 ( n16217 , n20680 , n8175 );
    and g8641 ( n32889 , n7360 , n10178 );
    and g8642 ( n3840 , n33806 , n33355 );
    xnor g8643 ( n35000 , n22650 , n33628 );
    or g8644 ( n14189 , n20626 , n28675 );
    or g8645 ( n29291 , n1950 , n9673 );
    nor g8646 ( n29044 , n9793 , n3784 );
    or g8647 ( n8315 , n11454 , n12412 );
    or g8648 ( n22828 , n2898 , n18488 );
    or g8649 ( n35713 , n31799 , n7050 );
    and g8650 ( n17500 , n18647 , n32283 );
    xnor g8651 ( n24114 , n28594 , n17568 );
    xnor g8652 ( n4524 , n22296 , n18887 );
    not g8653 ( n17067 , n22471 );
    or g8654 ( n8502 , n28174 , n1642 );
    xnor g8655 ( n12129 , n24212 , n27148 );
    or g8656 ( n25470 , n22037 , n24525 );
    or g8657 ( n34285 , n31386 , n16835 );
    or g8658 ( n10840 , n4793 , n10225 );
    or g8659 ( n7383 , n18013 , n29096 );
    not g8660 ( n2082 , n11455 );
    xnor g8661 ( n15553 , n21479 , n1969 );
    xnor g8662 ( n28686 , n1657 , n23015 );
    or g8663 ( n16838 , n34590 , n19421 );
    not g8664 ( n6678 , n12326 );
    and g8665 ( n22238 , n28950 , n9946 );
    and g8666 ( n30384 , n6355 , n7047 );
    or g8667 ( n4663 , n8188 , n27963 );
    xnor g8668 ( n8929 , n29001 , n19135 );
    or g8669 ( n11153 , n31799 , n19694 );
    and g8670 ( n14905 , n2423 , n18543 );
    and g8671 ( n18112 , n29814 , n7872 );
    nor g8672 ( n27393 , n13335 , n34391 );
    or g8673 ( n35924 , n29805 , n9498 );
    and g8674 ( n16554 , n3264 , n2442 );
    xnor g8675 ( n17121 , n4979 , n23604 );
    xnor g8676 ( n15457 , n13351 , n34263 );
    xnor g8677 ( n28178 , n30331 , n19637 );
    and g8678 ( n25394 , n16363 , n30868 );
    or g8679 ( n11075 , n7969 , n4646 );
    or g8680 ( n29978 , n27226 , n5995 );
    or g8681 ( n10989 , n1679 , n14717 );
    not g8682 ( n7844 , n6257 );
    not g8683 ( n5389 , n272 );
    nor g8684 ( n15793 , n17751 , n26921 );
    and g8685 ( n8266 , n9645 , n35289 );
    or g8686 ( n5542 , n18195 , n7647 );
    or g8687 ( n27323 , n9357 , n14699 );
    or g8688 ( n1301 , n16632 , n11703 );
    and g8689 ( n4939 , n8126 , n23229 );
    or g8690 ( n4672 , n28911 , n6075 );
    or g8691 ( n35021 , n31801 , n1856 );
    xnor g8692 ( n2250 , n27254 , n4758 );
    xor g8693 ( n27554 , n32692 , n12570 );
    not g8694 ( n29201 , n29029 );
    or g8695 ( n1672 , n12968 , n35748 );
    and g8696 ( n16585 , n8014 , n14188 );
    or g8697 ( n35082 , n13291 , n6764 );
    or g8698 ( n3355 , n19551 , n12797 );
    xnor g8699 ( n9255 , n33554 , n32257 );
    nor g8700 ( n4189 , n27493 , n25185 );
    not g8701 ( n18198 , n8695 );
    or g8702 ( n23955 , n2217 , n29592 );
    xnor g8703 ( n3320 , n22135 , n24371 );
    and g8704 ( n29023 , n5425 , n10724 );
    or g8705 ( n32743 , n24371 , n29497 );
    and g8706 ( n10818 , n9533 , n13507 );
    or g8707 ( n33779 , n28875 , n3188 );
    or g8708 ( n18717 , n19509 , n9601 );
    or g8709 ( n21101 , n1626 , n29562 );
    or g8710 ( n13984 , n5481 , n9030 );
    and g8711 ( n26256 , n2775 , n30890 );
    and g8712 ( n5770 , n24492 , n14395 );
    nor g8713 ( n11520 , n24265 , n2083 );
    or g8714 ( n7804 , n27849 , n14706 );
    and g8715 ( n34130 , n3057 , n32177 );
    or g8716 ( n28590 , n8432 , n36014 );
    or g8717 ( n24094 , n4906 , n28656 );
    or g8718 ( n24591 , n12307 , n16464 );
    or g8719 ( n20482 , n35671 , n25019 );
    and g8720 ( n11229 , n33987 , n10655 );
    and g8721 ( n19341 , n13658 , n17465 );
    or g8722 ( n4516 , n8176 , n2798 );
    or g8723 ( n28524 , n12073 , n26931 );
    xnor g8724 ( n15505 , n25793 , n4962 );
    not g8725 ( n21080 , n22241 );
    nor g8726 ( n30466 , n1950 , n20961 );
    xnor g8727 ( n12445 , n32332 , n20747 );
    or g8728 ( n29838 , n15878 , n30204 );
    xnor g8729 ( n25073 , n31911 , n4288 );
    not g8730 ( n28512 , n30742 );
    nor g8731 ( n34716 , n4960 , n1076 );
    or g8732 ( n13311 , n24371 , n8627 );
    nor g8733 ( n19379 , n3205 , n21995 );
    xnor g8734 ( n5801 , n10452 , n32584 );
    or g8735 ( n2868 , n34406 , n35845 );
    nor g8736 ( n7124 , n21336 , n29365 );
    not g8737 ( n30871 , n28273 );
    or g8738 ( n20479 , n9141 , n23626 );
    or g8739 ( n17717 , n25602 , n14958 );
    or g8740 ( n32800 , n5351 , n9930 );
    xnor g8741 ( n33773 , n14685 , n34323 );
    xnor g8742 ( n20226 , n4324 , n4962 );
    not g8743 ( n560 , n16102 );
    or g8744 ( n21535 , n33962 , n30714 );
    or g8745 ( n11192 , n7540 , n27994 );
    or g8746 ( n36 , n873 , n6026 );
    or g8747 ( n23856 , n29713 , n17701 );
    not g8748 ( n25941 , n11833 );
    or g8749 ( n1542 , n9687 , n29438 );
    and g8750 ( n16757 , n9594 , n2052 );
    and g8751 ( n28467 , n33344 , n25109 );
    xnor g8752 ( n7291 , n17351 , n9478 );
    xnor g8753 ( n34100 , n20647 , n31215 );
    or g8754 ( n15347 , n13654 , n17790 );
    or g8755 ( n12562 , n34821 , n959 );
    not g8756 ( n16156 , n5923 );
    or g8757 ( n28050 , n15863 , n9555 );
    nor g8758 ( n12227 , n23604 , n28393 );
    and g8759 ( n24836 , n3491 , n31346 );
    and g8760 ( n26354 , n9613 , n15836 );
    and g8761 ( n28661 , n24850 , n21006 );
    or g8762 ( n4528 , n6787 , n9030 );
    or g8763 ( n10927 , n5335 , n6469 );
    and g8764 ( n5020 , n10891 , n7596 );
    and g8765 ( n21525 , n1824 , n14998 );
    xnor g8766 ( n19015 , n27761 , n20104 );
    and g8767 ( n6945 , n22332 , n23029 );
    or g8768 ( n19268 , n9558 , n13822 );
    or g8769 ( n19648 , n21984 , n30389 );
    xnor g8770 ( n3103 , n8150 , n21903 );
    nor g8771 ( n24969 , n9980 , n12662 );
    nor g8772 ( n15925 , n31612 , n7700 );
    or g8773 ( n22760 , n5789 , n19125 );
    xnor g8774 ( n4141 , n35587 , n10894 );
    and g8775 ( n29748 , n26392 , n23465 );
    or g8776 ( n871 , n10571 , n5972 );
    or g8777 ( n11353 , n32857 , n27309 );
    xnor g8778 ( n10132 , n75 , n29713 );
    xnor g8779 ( n28943 , n24114 , n11823 );
    xnor g8780 ( n9220 , n25328 , n35561 );
    and g8781 ( n16905 , n6295 , n16165 );
    or g8782 ( n28775 , n27212 , n28866 );
    and g8783 ( n25478 , n15433 , n13460 );
    or g8784 ( n1443 , n6141 , n32808 );
    or g8785 ( n13016 , n26262 , n14076 );
    or g8786 ( n24605 , n25445 , n21644 );
    xnor g8787 ( n1272 , n23937 , n32095 );
    xnor g8788 ( n3029 , n6581 , n33471 );
    and g8789 ( n20109 , n16181 , n7852 );
    and g8790 ( n27759 , n27856 , n15227 );
    or g8791 ( n13157 , n9793 , n196 );
    or g8792 ( n6709 , n27805 , n30419 );
    or g8793 ( n18985 , n4924 , n7313 );
    not g8794 ( n31672 , n29801 );
    xnor g8795 ( n34403 , n31363 , n4878 );
    and g8796 ( n32875 , n30264 , n2606 );
    or g8797 ( n8532 , n6514 , n28455 );
    and g8798 ( n14990 , n7806 , n2463 );
    or g8799 ( n27703 , n19984 , n34300 );
    xnor g8800 ( n23444 , n26025 , n29178 );
    xnor g8801 ( n34432 , n22877 , n18858 );
    or g8802 ( n9854 , n30862 , n22783 );
    not g8803 ( n4659 , n17215 );
    xnor g8804 ( n4558 , n7068 , n15886 );
    xnor g8805 ( n23706 , n4196 , n5287 );
    or g8806 ( n4600 , n11285 , n29352 );
    or g8807 ( n5467 , n34883 , n10417 );
    and g8808 ( n35458 , n6436 , n1111 );
    and g8809 ( n22991 , n19020 , n11022 );
    nor g8810 ( n11597 , n4962 , n35128 );
    not g8811 ( n12024 , n10003 );
    or g8812 ( n22248 , n1658 , n19876 );
    and g8813 ( n33136 , n27618 , n28448 );
    nor g8814 ( n25755 , n4878 , n24539 );
    or g8815 ( n33834 , n2047 , n34888 );
    and g8816 ( n4624 , n12121 , n22523 );
    or g8817 ( n15019 , n19813 , n32808 );
    and g8818 ( n23307 , n21008 , n27204 );
    not g8819 ( n4739 , n16064 );
    buf g8820 ( n24489 , n3325 );
    nor g8821 ( n35736 , n4962 , n24349 );
    and g8822 ( n8223 , n11579 , n9056 );
    or g8823 ( n17770 , n7540 , n19915 );
    or g8824 ( n13142 , n14357 , n8665 );
    or g8825 ( n23645 , n21521 , n949 );
    or g8826 ( n136 , n15464 , n29995 );
    and g8827 ( n22222 , n11108 , n35560 );
    nor g8828 ( n28582 , n17568 , n1505 );
    xnor g8829 ( n21570 , n19768 , n10894 );
    not g8830 ( n33000 , n16223 );
    and g8831 ( n33043 , n4569 , n29095 );
    not g8832 ( n22243 , n6822 );
    or g8833 ( n20828 , n10197 , n4318 );
    or g8834 ( n10729 , n24371 , n20126 );
    or g8835 ( n26036 , n31215 , n30218 );
    or g8836 ( n32616 , n32476 , n16961 );
    or g8837 ( n13752 , n5559 , n19867 );
    and g8838 ( n34199 , n27566 , n10260 );
    nor g8839 ( n34834 , n4263 , n19942 );
    or g8840 ( n16701 , n7223 , n19971 );
    and g8841 ( n30256 , n26094 , n20828 );
    or g8842 ( n30678 , n30742 , n2061 );
    or g8843 ( n35571 , n1169 , n28668 );
    and g8844 ( n34891 , n34515 , n3825 );
    xnor g8845 ( n34156 , n28903 , n4546 );
    or g8846 ( n19839 , n21524 , n34995 );
    and g8847 ( n13796 , n21393 , n16873 );
    xnor g8848 ( n28779 , n36090 , n24371 );
    and g8849 ( n15148 , n21331 , n16211 );
    or g8850 ( n20100 , n26559 , n31464 );
    and g8851 ( n29391 , n7550 , n3499 );
    and g8852 ( n35170 , n727 , n23125 );
    not g8853 ( n20197 , n19551 );
    or g8854 ( n840 , n3946 , n14592 );
    xnor g8855 ( n2921 , n14445 , n9658 );
    or g8856 ( n14783 , n26671 , n5336 );
    not g8857 ( n22831 , n25174 );
    and g8858 ( n12155 , n29572 , n26981 );
    xnor g8859 ( n9664 , n12696 , n35292 );
    or g8860 ( n30424 , n18405 , n7673 );
    nor g8861 ( n35615 , n32715 , n7388 );
    or g8862 ( n24166 , n12890 , n2823 );
    or g8863 ( n310 , n26909 , n21691 );
    or g8864 ( n6109 , n15375 , n3352 );
    and g8865 ( n18269 , n20508 , n26845 );
    or g8866 ( n25969 , n11825 , n25306 );
    xnor g8867 ( n3375 , n13783 , n8851 );
    or g8868 ( n11065 , n24617 , n436 );
    or g8869 ( n24878 , n27180 , n10151 );
    and g8870 ( n33781 , n21291 , n32264 );
    and g8871 ( n26584 , n4339 , n20507 );
    not g8872 ( n18303 , n31977 );
    not g8873 ( n6081 , n2029 );
    or g8874 ( n25547 , n25319 , n7102 );
    or g8875 ( n2742 , n35691 , n21042 );
    or g8876 ( n20118 , n5685 , n33519 );
    or g8877 ( n10307 , n1950 , n27820 );
    not g8878 ( n35616 , n19455 );
    nor g8879 ( n20918 , n29839 , n14269 );
    and g8880 ( n13837 , n27058 , n35600 );
    or g8881 ( n22813 , n30921 , n18171 );
    and g8882 ( n33113 , n23734 , n7374 );
    and g8883 ( n239 , n15961 , n24891 );
    xnor g8884 ( n28027 , n31556 , n27476 );
    and g8885 ( n7365 , n20493 , n7581 );
    nor g8886 ( n25096 , n19984 , n21450 );
    xnor g8887 ( n4513 , n19333 , n8432 );
    or g8888 ( n27529 , n14533 , n25036 );
    or g8889 ( n33800 , n7470 , n11977 );
    or g8890 ( n27495 , n2357 , n15333 );
    and g8891 ( n5704 , n30783 , n34948 );
    and g8892 ( n14197 , n21842 , n8035 );
    xnor g8893 ( n5631 , n19977 , n24332 );
    xnor g8894 ( n34690 , n3885 , n26478 );
    or g8895 ( n23868 , n13544 , n8723 );
    xnor g8896 ( n8422 , n23333 , n24371 );
    nor g8897 ( n21179 , n3628 , n6548 );
    xnor g8898 ( n18625 , n17918 , n27643 );
    xnor g8899 ( n124 , n20838 , n4960 );
    xnor g8900 ( n8119 , n21231 , n28461 );
    not g8901 ( n28095 , n17335 );
    and g8902 ( n21056 , n8598 , n21858 );
    or g8903 ( n27183 , n32095 , n16989 );
    and g8904 ( n28941 , n12936 , n34592 );
    and g8905 ( n34081 , n1347 , n35298 );
    or g8906 ( n11723 , n34604 , n1715 );
    or g8907 ( n16142 , n16884 , n34971 );
    not g8908 ( n36072 , n1950 );
    or g8909 ( n8143 , n30417 , n26486 );
    not g8910 ( n27237 , n27226 );
    not g8911 ( n26600 , n25110 );
    and g8912 ( n14407 , n30580 , n10590 );
    or g8913 ( n20561 , n11567 , n25355 );
    or g8914 ( n20322 , n10437 , n7293 );
    or g8915 ( n9945 , n33989 , n15084 );
    or g8916 ( n3791 , n19551 , n10317 );
    or g8917 ( n8754 , n25997 , n27574 );
    or g8918 ( n29801 , n4519 , n28123 );
    and g8919 ( n13315 , n30548 , n29482 );
    or g8920 ( n33404 , n17607 , n30732 );
    nor g8921 ( n29581 , n1160 , n14677 );
    and g8922 ( n30054 , n9781 , n19806 );
    xnor g8923 ( n18299 , n24940 , n32857 );
    or g8924 ( n2738 , n27811 , n27625 );
    or g8925 ( n16474 , n11296 , n26705 );
    xnor g8926 ( n17606 , n18689 , n32715 );
    or g8927 ( n18584 , n28389 , n6020 );
    and g8928 ( n5626 , n16214 , n33794 );
    or g8929 ( n3789 , n34545 , n530 );
    xnor g8930 ( n22390 , n22413 , n24371 );
    xnor g8931 ( n18988 , n4857 , n32715 );
    or g8932 ( n15227 , n5335 , n27337 );
    or g8933 ( n4849 , n4186 , n9731 );
    and g8934 ( n17441 , n24649 , n7977 );
    or g8935 ( n30463 , n4878 , n32169 );
    or g8936 ( n14622 , n22705 , n12163 );
    xnor g8937 ( n21116 , n18891 , n9793 );
    xnor g8938 ( n30374 , n24713 , n27226 );
    or g8939 ( n21423 , n11010 , n3858 );
    xnor g8940 ( n12549 , n10589 , n23895 );
    xnor g8941 ( n15388 , n13691 , n3312 );
    xnor g8942 ( n12346 , n14849 , n32715 );
    and g8943 ( n25149 , n34603 , n2969 );
    or g8944 ( n31033 , n30399 , n27574 );
    nor g8945 ( n32896 , n16620 , n21941 );
    or g8946 ( n20309 , n12881 , n6340 );
    or g8947 ( n19119 , n10604 , n29754 );
    and g8948 ( n25657 , n33516 , n34788 );
    nor g8949 ( n9298 , n29202 , n753 );
    and g8950 ( n3348 , n22207 , n18586 );
    or g8951 ( n30001 , n8231 , n6478 );
    not g8952 ( n10452 , n7775 );
    not g8953 ( n4442 , n969 );
    not g8954 ( n21950 , n24731 );
    and g8955 ( n20603 , n25034 , n26414 );
    xnor g8956 ( n23800 , n7577 , n4288 );
    xnor g8957 ( n12866 , n11709 , n17568 );
    or g8958 ( n16047 , n31799 , n4314 );
    or g8959 ( n31905 , n16966 , n18406 );
    xnor g8960 ( n30506 , n8902 , n8077 );
    xnor g8961 ( n21296 , n35803 , n870 );
    nor g8962 ( n26087 , n16620 , n20205 );
    and g8963 ( n23811 , n31066 , n9001 );
    or g8964 ( n15725 , n29184 , n19490 );
    and g8965 ( n23221 , n22509 , n1017 );
    xnor g8966 ( n15114 , n4220 , n30481 );
    and g8967 ( n6437 , n2070 , n12513 );
    not g8968 ( n15351 , n18002 );
    xnor g8969 ( n18072 , n16508 , n8871 );
    or g8970 ( n9972 , n15886 , n2841 );
    not g8971 ( n2799 , n25174 );
    and g8972 ( n31507 , n23904 , n32383 );
    xnor g8973 ( n10805 , n32080 , n34367 );
    or g8974 ( n28753 , n32857 , n14817 );
    or g8975 ( n7409 , n16620 , n16081 );
    or g8976 ( n2100 , n23824 , n34816 );
    and g8977 ( n14766 , n4542 , n27961 );
    xnor g8978 ( n10798 , n17633 , n19551 );
    xnor g8979 ( n27941 , n10940 , n14933 );
    or g8980 ( n25877 , n33429 , n24375 );
    or g8981 ( n6797 , n24371 , n9760 );
    or g8982 ( n8102 , n31602 , n13952 );
    or g8983 ( n23873 , n18270 , n26659 );
    xnor g8984 ( n19682 , n21138 , n28282 );
    xnor g8985 ( n12928 , n11964 , n34381 );
    or g8986 ( n31444 , n12902 , n10397 );
    or g8987 ( n20162 , n22291 , n2462 );
    or g8988 ( n34163 , n1425 , n28438 );
    not g8989 ( n8876 , n19577 );
    or g8990 ( n26992 , n5963 , n14746 );
    nor g8991 ( n20859 , n32857 , n20109 );
    or g8992 ( n23197 , n32778 , n26737 );
    nor g8993 ( n28169 , n16620 , n6116 );
    nor g8994 ( n10627 , n27226 , n18301 );
    or g8995 ( n35272 , n23666 , n4081 );
    or g8996 ( n25287 , n30228 , n29288 );
    or g8997 ( n323 , n19047 , n27801 );
    xnor g8998 ( n18531 , n5627 , n17751 );
    or g8999 ( n4052 , n20269 , n16797 );
    or g9000 ( n14869 , n12926 , n3044 );
    and g9001 ( n15906 , n19081 , n17949 );
    xnor g9002 ( n8901 , n25118 , n781 );
    or g9003 ( n26403 , n28308 , n18358 );
    or g9004 ( n28977 , n19048 , n34084 );
    or g9005 ( n10970 , n17568 , n1222 );
    and g9006 ( n7385 , n20839 , n35127 );
    not g9007 ( n11028 , n18198 );
    or g9008 ( n4942 , n22842 , n12596 );
    buf g9009 ( n12696 , n9088 );
    xnor g9010 ( n7713 , n32601 , n16135 );
    and g9011 ( n13290 , n23005 , n14222 );
    not g9012 ( n1635 , n31054 );
    xnor g9013 ( n27992 , n22050 , n30742 );
    or g9014 ( n21031 , n7108 , n18264 );
    xnor g9015 ( n12656 , n8609 , n35927 );
    or g9016 ( n25132 , n15022 , n34971 );
    not g9017 ( n19512 , n31460 );
    xnor g9018 ( n6038 , n7452 , n26092 );
    or g9019 ( n4688 , n12832 , n18877 );
    and g9020 ( n14700 , n28282 , n21138 );
    xnor g9021 ( n6004 , n4948 , n8538 );
    or g9022 ( n4968 , n6872 , n1744 );
    not g9023 ( n35644 , n10423 );
    xnor g9024 ( n9442 , n28863 , n19267 );
    xnor g9025 ( n4855 , n32060 , n4185 );
    xnor g9026 ( n24764 , n35914 , n9793 );
    and g9027 ( n17539 , n34674 , n26740 );
    and g9028 ( n23133 , n857 , n15680 );
    not g9029 ( n17009 , n30732 );
    not g9030 ( n27391 , n3205 );
    or g9031 ( n32432 , n8260 , n26595 );
    xnor g9032 ( n21032 , n8229 , n24061 );
    nor g9033 ( n17164 , n16703 , n31411 );
    nor g9034 ( n30925 , n22291 , n26950 );
    and g9035 ( n24120 , n24799 , n17350 );
    xnor g9036 ( n13575 , n29194 , n11190 );
    and g9037 ( n33060 , n28768 , n30959 );
    or g9038 ( n8003 , n32060 , n4185 );
    and g9039 ( n30687 , n6167 , n18751 );
    and g9040 ( n14357 , n20865 , n22980 );
    and g9041 ( n5152 , n14872 , n28112 );
    or g9042 ( n7070 , n21496 , n30431 );
    or g9043 ( n15136 , n5335 , n25492 );
    or g9044 ( n4680 , n24107 , n7709 );
    or g9045 ( n17064 , n13501 , n16781 );
    or g9046 ( n33020 , n29056 , n8575 );
    or g9047 ( n8757 , n4165 , n19125 );
    xnor g9048 ( n9943 , n21275 , n19113 );
    and g9049 ( n13952 , n2150 , n11082 );
    or g9050 ( n11462 , n14957 , n2119 );
    or g9051 ( n31340 , n13101 , n32505 );
    and g9052 ( n2621 , n7986 , n16208 );
    or g9053 ( n1004 , n31215 , n12669 );
    not g9054 ( n28780 , n16045 );
    or g9055 ( n21427 , n1003 , n28252 );
    xnor g9056 ( n2510 , n30368 , n5335 );
    xnor g9057 ( n13515 , n34580 , n23927 );
    or g9058 ( n34858 , n20554 , n22961 );
    not g9059 ( n26317 , n25847 );
    nor g9060 ( n24772 , n4860 , n26292 );
    or g9061 ( n30916 , n13266 , n32959 );
    xnor g9062 ( n30955 , n30328 , n9793 );
    and g9063 ( n6314 , n16572 , n13371 );
    or g9064 ( n17999 , n3542 , n19107 );
    xnor g9065 ( n7799 , n8121 , n16897 );
    or g9066 ( n17669 , n18574 , n25306 );
    nor g9067 ( n28202 , n26376 , n15185 );
    xnor g9068 ( n25081 , n897 , n3222 );
    or g9069 ( n12141 , n16808 , n7306 );
    or g9070 ( n19716 , n26041 , n13255 );
    or g9071 ( n22605 , n33222 , n9951 );
    or g9072 ( n33292 , n5691 , n10313 );
    or g9073 ( n27048 , n13135 , n8539 );
    xnor g9074 ( n14641 , n24445 , n11455 );
    and g9075 ( n4742 , n24149 , n28473 );
    or g9076 ( n27768 , n23380 , n14308 );
    and g9077 ( n7711 , n29826 , n6389 );
    and g9078 ( n4635 , n31795 , n18029 );
    or g9079 ( n33603 , n35995 , n26653 );
    and g9080 ( n25373 , n2101 , n29128 );
    or g9081 ( n15830 , n11706 , n11261 );
    xnor g9082 ( n15824 , n24703 , n7784 );
    or g9083 ( n30612 , n2420 , n31464 );
    xnor g9084 ( n25931 , n14179 , n5114 );
    or g9085 ( n32342 , n17028 , n15210 );
    xnor g9086 ( n23632 , n32885 , n8446 );
    nor g9087 ( n15251 , n29177 , n3806 );
    or g9088 ( n4625 , n31056 , n22483 );
    xnor g9089 ( n2400 , n7014 , n25602 );
    or g9090 ( n16916 , n16135 , n6205 );
    or g9091 ( n13494 , n12867 , n31606 );
    xnor g9092 ( n3008 , n23768 , n21223 );
    xnor g9093 ( n8356 , n16953 , n8432 );
    or g9094 ( n6112 , n30094 , n1856 );
    and g9095 ( n17744 , n16308 , n4182 );
    xnor g9096 ( n6751 , n19948 , n21630 );
    xnor g9097 ( n32156 , n449 , n7125 );
    xnor g9098 ( n35424 , n16891 , n28255 );
    or g9099 ( n26845 , n11046 , n19741 );
    xnor g9100 ( n17573 , n11546 , n13642 );
    or g9101 ( n16658 , n4475 , n21862 );
    or g9102 ( n16093 , n13897 , n4187 );
    nor g9103 ( n175 , n23604 , n20821 );
    or g9104 ( n12706 , n25331 , n13058 );
    not g9105 ( n16577 , n28336 );
    xnor g9106 ( n5844 , n16906 , n6201 );
    xnor g9107 ( n20834 , n7043 , n27226 );
    xnor g9108 ( n26875 , n8083 , n4639 );
    or g9109 ( n29100 , n10239 , n33117 );
    and g9110 ( n21477 , n3065 , n31915 );
    or g9111 ( n35836 , n23213 , n14706 );
    and g9112 ( n28104 , n18010 , n11920 );
    or g9113 ( n34562 , n12692 , n32495 );
    xnor g9114 ( n16173 , n22808 , n26008 );
    or g9115 ( n36047 , n3205 , n33311 );
    or g9116 ( n25843 , n3946 , n13796 );
    or g9117 ( n1167 , n20694 , n28455 );
    or g9118 ( n17333 , n3332 , n15459 );
    xnor g9119 ( n3574 , n2176 , n11190 );
    xnor g9120 ( n19757 , n750 , n30680 );
    and g9121 ( n29514 , n23000 , n3407 );
    or g9122 ( n11583 , n21381 , n4478 );
    nor g9123 ( n14471 , n32095 , n12677 );
    and g9124 ( n28743 , n27579 , n3366 );
    xor g9125 ( n26056 , n6093 , n26747 );
    and g9126 ( n16390 , n11169 , n30 );
    and g9127 ( n1010 , n30379 , n4392 );
    and g9128 ( n8063 , n25756 , n27677 );
    xnor g9129 ( n24847 , n9379 , n32658 );
    or g9130 ( n20185 , n9574 , n1424 );
    nor g9131 ( n6328 , n32574 , n25795 );
    or g9132 ( n5651 , n28802 , n33924 );
    nor g9133 ( n21887 , n2647 , n35429 );
    not g9134 ( n8098 , n22241 );
    or g9135 ( n11100 , n10041 , n23266 );
    or g9136 ( n27200 , n27098 , n5146 );
    xnor g9137 ( n6877 , n1496 , n35815 );
    not g9138 ( n5138 , n20558 );
    nor g9139 ( n19304 , n3205 , n948 );
    or g9140 ( n19003 , n16034 , n35043 );
    nor g9141 ( n30613 , n30742 , n15697 );
    nor g9142 ( n20824 , n24816 , n16698 );
    nor g9143 ( n27921 , n12062 , n28503 );
    and g9144 ( n11471 , n2687 , n16359 );
    xnor g9145 ( n1726 , n19210 , n4288 );
    not g9146 ( n25629 , n22980 );
    and g9147 ( n7428 , n24661 , n15761 );
    and g9148 ( n13537 , n8769 , n18732 );
    nor g9149 ( n19438 , n32584 , n682 );
    buf g9150 ( n16649 , n27816 );
    or g9151 ( n32015 , n25883 , n16338 );
    and g9152 ( n34994 , n24676 , n25517 );
    xnor g9153 ( n28968 , n28981 , n30742 );
    or g9154 ( n32115 , n30768 , n4203 );
    and g9155 ( n23435 , n5105 , n11861 );
    xnor g9156 ( n6440 , n27824 , n32857 );
    or g9157 ( n9866 , n22082 , n474 );
    or g9158 ( n21751 , n26703 , n20318 );
    or g9159 ( n26605 , n34327 , n5779 );
    not g9160 ( n4367 , n28893 );
    or g9161 ( n4535 , n16988 , n13949 );
    and g9162 ( n32603 , n547 , n20388 );
    or g9163 ( n16714 , n5350 , n640 );
    buf g9164 ( n29953 , n14292 );
    xnor g9165 ( n12185 , n6864 , n3205 );
    xnor g9166 ( n6765 , n11456 , n4288 );
    or g9167 ( n14644 , n19323 , n9933 );
    and g9168 ( n16534 , n13653 , n30420 );
    not g9169 ( n30636 , n24332 );
    or g9170 ( n3801 , n16286 , n14841 );
    xnor g9171 ( n17542 , n7847 , n31559 );
    or g9172 ( n2858 , n32622 , n27580 );
    and g9173 ( n15213 , n34581 , n18476 );
    xnor g9174 ( n7233 , n27899 , n13056 );
    nor g9175 ( n23342 , n5287 , n15621 );
    not g9176 ( n9661 , n2029 );
    xnor g9177 ( n28173 , n25943 , n5337 );
    not g9178 ( n34724 , n24847 );
    xnor g9179 ( n18247 , n28549 , n32095 );
    and g9180 ( n19338 , n24706 , n23548 );
    not g9181 ( n7101 , n27738 );
    or g9182 ( n4943 , n31531 , n17829 );
    and g9183 ( n35457 , n8741 , n7558 );
    or g9184 ( n19222 , n16620 , n23478 );
    xnor g9185 ( n30649 , n9552 , n24836 );
    xnor g9186 ( n16234 , n24766 , n3222 );
    and g9187 ( n113 , n31213 , n6404 );
    and g9188 ( n13284 , n32384 , n5935 );
    xnor g9189 ( n22538 , n10575 , n21872 );
    not g9190 ( n17758 , n2664 );
    or g9191 ( n9152 , n10498 , n9832 );
    or g9192 ( n21246 , n20395 , n20812 );
    and g9193 ( n20717 , n31162 , n32805 );
    xnor g9194 ( n27358 , n1538 , n35927 );
    or g9195 ( n34266 , n6796 , n19942 );
    xnor g9196 ( n1575 , n20995 , n83 );
    xnor g9197 ( n36086 , n2587 , n31310 );
    or g9198 ( n5715 , n4878 , n29515 );
    or g9199 ( n17834 , n6895 , n11996 );
    xor g9200 ( n16650 , n33450 , n15473 );
    and g9201 ( n21396 , n6491 , n9908 );
    not g9202 ( n14174 , n31272 );
    or g9203 ( n3435 , n28892 , n30752 );
    and g9204 ( n569 , n23207 , n13354 );
    and g9205 ( n11274 , n14203 , n20320 );
    nor g9206 ( n4086 , n830 , n32597 );
    xnor g9207 ( n4539 , n5503 , n11067 );
    or g9208 ( n12716 , n8358 , n4490 );
    or g9209 ( n24507 , n13732 , n7293 );
    not g9210 ( n19245 , n23786 );
    or g9211 ( n30163 , n31415 , n18930 );
    and g9212 ( n32688 , n29405 , n7946 );
    xnor g9213 ( n11966 , n22126 , n12523 );
    or g9214 ( n22315 , n10893 , n18995 );
    or g9215 ( n18928 , n20677 , n6950 );
    xnor g9216 ( n33490 , n29699 , n23604 );
    or g9217 ( n23016 , n7336 , n17879 );
    xnor g9218 ( n8525 , n16366 , n34285 );
    or g9219 ( n18031 , n6556 , n24259 );
    or g9220 ( n3661 , n15204 , n27973 );
    or g9221 ( n1651 , n32436 , n27392 );
    xnor g9222 ( n2045 , n33611 , n15299 );
    or g9223 ( n35135 , n14344 , n26308 );
    nor g9224 ( n14089 , n21171 , n29847 );
    or g9225 ( n34194 , n1429 , n30039 );
    xnor g9226 ( n20184 , n31591 , n28702 );
    and g9227 ( n32549 , n16901 , n22593 );
    or g9228 ( n14913 , n18196 , n3298 );
    xnor g9229 ( n29964 , n7631 , n15403 );
    or g9230 ( n8424 , n4232 , n11226 );
    xnor g9231 ( n32900 , n11111 , n29229 );
    or g9232 ( n9056 , n22101 , n20701 );
    or g9233 ( n7141 , n7909 , n15265 );
    or g9234 ( n10136 , n22291 , n26287 );
    and g9235 ( n2509 , n1668 , n31021 );
    and g9236 ( n22689 , n17997 , n12960 );
    nor g9237 ( n27673 , n25174 , n21778 );
    or g9238 ( n25666 , n11190 , n5690 );
    and g9239 ( n12678 , n30118 , n30900 );
    or g9240 ( n11664 , n6114 , n957 );
    or g9241 ( n14779 , n5402 , n17962 );
    xnor g9242 ( n34411 , n1702 , n1318 );
    or g9243 ( n22714 , n27295 , n27447 );
    xnor g9244 ( n10916 , n3992 , n14563 );
    or g9245 ( n9654 , n12886 , n17354 );
    or g9246 ( n33237 , n16491 , n8090 );
    xnor g9247 ( n24990 , n2342 , n29277 );
    xnor g9248 ( n21629 , n34497 , n26770 );
    nor g9249 ( n2460 , n26317 , n20379 );
    or g9250 ( n27273 , n21045 , n13480 );
    not g9251 ( n34850 , n16467 );
    and g9252 ( n29156 , n11099 , n19350 );
    and g9253 ( n31804 , n26722 , n31604 );
    xnor g9254 ( n1556 , n27038 , n32391 );
    xnor g9255 ( n4021 , n19476 , n26877 );
    and g9256 ( n20303 , n32547 , n22128 );
    or g9257 ( n26932 , n35769 , n8924 );
    not g9258 ( n18580 , n33024 );
    nor g9259 ( n13654 , n19551 , n17322 );
    and g9260 ( n8387 , n24490 , n21770 );
    or g9261 ( n17283 , n15464 , n5015 );
    nor g9262 ( n24375 , n29130 , n5457 );
    and g9263 ( n11538 , n14155 , n3039 );
    xnor g9264 ( n3258 , n21786 , n29995 );
    or g9265 ( n22179 , n34819 , n3979 );
    xnor g9266 ( n7129 , n28 , n13254 );
    nor g9267 ( n17006 , n34677 , n27641 );
    or g9268 ( n4238 , n18300 , n11703 );
    or g9269 ( n22078 , n31559 , n17725 );
    or g9270 ( n14036 , n32857 , n5286 );
    or g9271 ( n14509 , n4962 , n23064 );
    and g9272 ( n28549 , n22897 , n21772 );
    or g9273 ( n11931 , n26695 , n28123 );
    or g9274 ( n20145 , n1950 , n21707 );
    and g9275 ( n27960 , n8055 , n27591 );
    or g9276 ( n25007 , n22090 , n19403 );
    not g9277 ( n12409 , n9506 );
    xnor g9278 ( n4257 , n1541 , n4758 );
    xnor g9279 ( n13041 , n8124 , n13933 );
    or g9280 ( n24977 , n29802 , n2955 );
    or g9281 ( n28366 , n13831 , n20690 );
    and g9282 ( n26428 , n36028 , n15633 );
    or g9283 ( n22721 , n8025 , n35714 );
    or g9284 ( n16853 , n3222 , n12286 );
    or g9285 ( n13891 , n26255 , n9966 );
    and g9286 ( n29273 , n1184 , n14403 );
    or g9287 ( n23771 , n23604 , n30530 );
    and g9288 ( n2651 , n1720 , n4133 );
    or g9289 ( n26516 , n28247 , n21644 );
    or g9290 ( n3085 , n29681 , n20817 );
    and g9291 ( n4868 , n23802 , n22 );
    or g9292 ( n14521 , n6732 , n24672 );
    xnor g9293 ( n2344 , n14320 , n32689 );
    or g9294 ( n3122 , n16052 , n29761 );
    and g9295 ( n33578 , n23331 , n33934 );
    xnor g9296 ( n13566 , n6127 , n1950 );
    xnor g9297 ( n11481 , n27585 , n7965 );
    xnor g9298 ( n11143 , n8625 , n7883 );
    and g9299 ( n5587 , n16902 , n16393 );
    and g9300 ( n28789 , n33820 , n20116 );
    and g9301 ( n35584 , n26766 , n33235 );
    or g9302 ( n32162 , n7658 , n9030 );
    xnor g9303 ( n22025 , n11253 , n26360 );
    and g9304 ( n32083 , n32211 , n34589 );
    xnor g9305 ( n21165 , n28143 , n23604 );
    or g9306 ( n35018 , n31742 , n29643 );
    or g9307 ( n30841 , n13736 , n12128 );
    or g9308 ( n34522 , n5356 , n16668 );
    xnor g9309 ( n7917 , n21679 , n31289 );
    and g9310 ( n21410 , n25864 , n20454 );
    or g9311 ( n28991 , n30164 , n18203 );
    or g9312 ( n31126 , n17407 , n23537 );
    xnor g9313 ( n23171 , n30799 , n32857 );
    or g9314 ( n13441 , n29662 , n35422 );
    or g9315 ( n16198 , n29009 , n1250 );
    and g9316 ( n13786 , n238 , n5496 );
    xnor g9317 ( n22401 , n8351 , n2716 );
    or g9318 ( n21442 , n11455 , n33485 );
    and g9319 ( n9379 , n20004 , n22721 );
    and g9320 ( n17401 , n32893 , n1956 );
    or g9321 ( n21449 , n28342 , n3858 );
    xnor g9322 ( n11349 , n16794 , n11455 );
    and g9323 ( n33733 , n404 , n33408 );
    nor g9324 ( n5135 , n15475 , n16564 );
    or g9325 ( n19735 , n1950 , n24550 );
    or g9326 ( n10092 , n4288 , n2639 );
    or g9327 ( n9305 , n25760 , n24356 );
    or g9328 ( n15859 , n28073 , n4751 );
    or g9329 ( n7992 , n18074 , n29852 );
    and g9330 ( n33633 , n13873 , n10006 );
    buf g9331 ( n29393 , n6521 );
    or g9332 ( n7045 , n31289 , n5066 );
    or g9333 ( n29035 , n34876 , n25240 );
    and g9334 ( n3864 , n4453 , n12919 );
    and g9335 ( n15752 , n13309 , n6188 );
    or g9336 ( n34643 , n16156 , n32366 );
    xnor g9337 ( n15480 , n30006 , n19984 );
    xor g9338 ( n26271 , n20933 , n29558 );
    or g9339 ( n25880 , n31215 , n7172 );
    or g9340 ( n30977 , n30742 , n17312 );
    xor g9341 ( n24972 , n19811 , n14547 );
    and g9342 ( n10128 , n21306 , n11087 );
    and g9343 ( n14959 , n18684 , n13206 );
    or g9344 ( n1834 , n3780 , n35111 );
    or g9345 ( n15511 , n3271 , n23790 );
    or g9346 ( n15612 , n3484 , n29439 );
    not g9347 ( n2064 , n16620 );
    or g9348 ( n16351 , n23221 , n26112 );
    xnor g9349 ( n6769 , n1867 , n16135 );
    and g9350 ( n508 , n9143 , n7890 );
    nor g9351 ( n9008 , n32857 , n21420 );
    or g9352 ( n20835 , n11326 , n5252 );
    and g9353 ( n7363 , n23364 , n7862 );
    or g9354 ( n34838 , n22291 , n11254 );
    or g9355 ( n20149 , n11004 , n10463 );
    or g9356 ( n404 , n31214 , n12058 );
    xnor g9357 ( n34553 , n18266 , n31799 );
    nor g9358 ( n6240 , n30636 , n27858 );
    xnor g9359 ( n12095 , n3136 , n17568 );
    xnor g9360 ( n1054 , n35241 , n32857 );
    and g9361 ( n22610 , n8133 , n9750 );
    and g9362 ( n7674 , n29406 , n24792 );
    or g9363 ( n31689 , n5075 , n19952 );
    xnor g9364 ( n651 , n34562 , n11046 );
    or g9365 ( n13669 , n35915 , n30569 );
    xnor g9366 ( n7420 , n15300 , n2177 );
    or g9367 ( n28263 , n15156 , n23512 );
    xnor g9368 ( n4547 , n3353 , n2472 );
    not g9369 ( n31919 , n4878 );
    or g9370 ( n25929 , n16986 , n5752 );
    and g9371 ( n23334 , n2530 , n13584 );
    xnor g9372 ( n11838 , n22846 , n29510 );
    and g9373 ( n20295 , n17768 , n16857 );
    xnor g9374 ( n5036 , n34586 , n8910 );
    or g9375 ( n8906 , n29831 , n4318 );
    xnor g9376 ( n6854 , n13497 , n18850 );
    xnor g9377 ( n18067 , n26625 , n31918 );
    and g9378 ( n14306 , n24516 , n2062 );
    xnor g9379 ( n23983 , n23106 , n12442 );
    or g9380 ( n30131 , n21857 , n35294 );
    or g9381 ( n35159 , n34512 , n25761 );
    and g9382 ( n34297 , n3117 , n35300 );
    not g9383 ( n19927 , n252 );
    and g9384 ( n28314 , n17574 , n24540 );
    or g9385 ( n13070 , n3520 , n4743 );
    nor g9386 ( n33944 , n32584 , n30049 );
    or g9387 ( n1002 , n30664 , n25548 );
    nor g9388 ( n6782 , n11046 , n30070 );
    nor g9389 ( n5998 , n8432 , n15669 );
    buf g9390 ( n27053 , n1793 );
    xnor g9391 ( n15201 , n15918 , n478 );
    and g9392 ( n13123 , n7107 , n30842 );
    or g9393 ( n8873 , n27941 , n28404 );
    or g9394 ( n34490 , n29839 , n2276 );
    or g9395 ( n4870 , n4796 , n21926 );
    and g9396 ( n15547 , n13289 , n34838 );
    or g9397 ( n627 , n32774 , n25255 );
    or g9398 ( n35139 , n9625 , n28248 );
    and g9399 ( n8881 , n6744 , n29689 );
    xnor g9400 ( n22888 , n16879 , n30883 );
    or g9401 ( n11946 , n18724 , n19783 );
    not g9402 ( n9232 , n14017 );
    or g9403 ( n31132 , n27548 , n5900 );
    or g9404 ( n21437 , n34390 , n22682 );
    or g9405 ( n9372 , n9793 , n1852 );
    or g9406 ( n22112 , n15336 , n28553 );
    or g9407 ( n7725 , n16336 , n5779 );
    nor g9408 ( n9986 , n31559 , n25690 );
    nor g9409 ( n27729 , n20212 , n31411 );
    xnor g9410 ( n30090 , n29011 , n8298 );
    or g9411 ( n22387 , n7239 , n18264 );
    or g9412 ( n8912 , n11595 , n36000 );
    or g9413 ( n3065 , n20190 , n2513 );
    or g9414 ( n18690 , n3103 , n27728 );
    and g9415 ( n35719 , n12551 , n32247 );
    not g9416 ( n28541 , n33596 );
    xnor g9417 ( n34798 , n6098 , n14550 );
    or g9418 ( n7806 , n23980 , n11850 );
    xnor g9419 ( n20183 , n31112 , n31559 );
    and g9420 ( n12328 , n12460 , n17621 );
    or g9421 ( n19072 , n24371 , n22991 );
    or g9422 ( n29893 , n14458 , n28866 );
    nor g9423 ( n10303 , n31799 , n27803 );
    or g9424 ( n25885 , n13282 , n6075 );
    not g9425 ( n9447 , n33381 );
    or g9426 ( n7741 , n32473 , n11638 );
    and g9427 ( n25475 , n30044 , n12946 );
    or g9428 ( n26530 , n32095 , n28212 );
    and g9429 ( n18918 , n14919 , n14900 );
    or g9430 ( n2643 , n3222 , n8564 );
    or g9431 ( n30275 , n15886 , n26010 );
    not g9432 ( n7940 , n14126 );
    and g9433 ( n12834 , n2652 , n19343 );
    and g9434 ( n33475 , n22969 , n22012 );
    or g9435 ( n32355 , n22595 , n9847 );
    or g9436 ( n11668 , n30488 , n28064 );
    or g9437 ( n17956 , n13701 , n19866 );
    xnor g9438 ( n32102 , n10860 , n18379 );
    or g9439 ( n32737 , n22539 , n29231 );
    and g9440 ( n8882 , n14331 , n14084 );
    and g9441 ( n8487 , n8029 , n1075 );
    nor g9442 ( n19917 , n31559 , n32157 );
    and g9443 ( n489 , n14052 , n14125 );
    not g9444 ( n18478 , n10072 );
    and g9445 ( n10887 , n30991 , n35843 );
    nor g9446 ( n31155 , n32952 , n9555 );
    nor g9447 ( n10562 , n27226 , n26048 );
    xnor g9448 ( n5660 , n29151 , n16717 );
    xnor g9449 ( n8543 , n5604 , n8292 );
    or g9450 ( n10468 , n8655 , n30292 );
    xnor g9451 ( n24778 , n32325 , n29855 );
    not g9452 ( n24700 , n10068 );
    and g9453 ( n35328 , n12471 , n34935 );
    or g9454 ( n34768 , n13910 , n30708 );
    or g9455 ( n19480 , n28014 , n25306 );
    and g9456 ( n29640 , n19238 , n853 );
    or g9457 ( n23623 , n3326 , n28438 );
    or g9458 ( n25777 , n7693 , n14161 );
    or g9459 ( n21584 , n20246 , n6553 );
    and g9460 ( n30658 , n18251 , n2858 );
    buf g9461 ( n5752 , n31990 );
    and g9462 ( n26866 , n32954 , n2347 );
    xnor g9463 ( n30360 , n13791 , n8701 );
    and g9464 ( n29148 , n15046 , n8216 );
    or g9465 ( n20046 , n1593 , n34363 );
    and g9466 ( n6742 , n13066 , n12426 );
    buf g9467 ( n1557 , n22753 );
    or g9468 ( n22913 , n12935 , n4348 );
    or g9469 ( n13170 , n11576 , n26374 );
    buf g9470 ( n8366 , n14579 );
    xnor g9471 ( n20981 , n19509 , n31799 );
    nor g9472 ( n15067 , n35075 , n7184 );
    and g9473 ( n18381 , n16513 , n10546 );
    or g9474 ( n34584 , n19088 , n11261 );
    xnor g9475 ( n28401 , n14980 , n3016 );
    or g9476 ( n12891 , n7991 , n11940 );
    xnor g9477 ( n30630 , n26146 , n7540 );
    not g9478 ( n1066 , n14068 );
    or g9479 ( n1073 , n10754 , n24929 );
    xnor g9480 ( n1332 , n20785 , n10894 );
    or g9481 ( n33402 , n30976 , n16566 );
    or g9482 ( n26564 , n3222 , n4050 );
    not g9483 ( n15515 , n29839 );
    and g9484 ( n10905 , n18948 , n25766 );
    and g9485 ( n15534 , n11493 , n12628 );
    and g9486 ( n23455 , n10438 , n8020 );
    and g9487 ( n13565 , n4588 , n12777 );
    xnor g9488 ( n16967 , n699 , n24053 );
    xnor g9489 ( n9775 , n7245 , n15757 );
    buf g9490 ( n3805 , n30441 );
    or g9491 ( n6268 , n1883 , n16060 );
    not g9492 ( n10607 , n4960 );
    nor g9493 ( n10217 , n17568 , n10660 );
    or g9494 ( n8280 , n32857 , n21611 );
    and g9495 ( n32114 , n25974 , n15325 );
    or g9496 ( n4240 , n19362 , n9796 );
    or g9497 ( n27409 , n35668 , n12606 );
    or g9498 ( n33895 , n24640 , n12465 );
    not g9499 ( n21792 , n29203 );
    xnor g9500 ( n14944 , n16547 , n31056 );
    or g9501 ( n24352 , n6685 , n23805 );
    not g9502 ( n24699 , n18310 );
    or g9503 ( n8763 , n32857 , n17436 );
    or g9504 ( n3242 , n9463 , n16555 );
    or g9505 ( n15992 , n22080 , n6678 );
    not g9506 ( n9848 , n6489 );
    and g9507 ( n35227 , n3130 , n12195 );
    or g9508 ( n23236 , n5548 , n25597 );
    and g9509 ( n8044 , n470 , n34901 );
    nor g9510 ( n11458 , n6028 , n12658 );
    or g9511 ( n29293 , n9658 , n623 );
    and g9512 ( n5995 , n10782 , n3967 );
    or g9513 ( n25009 , n31056 , n3540 );
    xnor g9514 ( n17854 , n12838 , n26128 );
    and g9515 ( n14732 , n8477 , n31748 );
    or g9516 ( n31396 , n5441 , n4912 );
    or g9517 ( n18725 , n11943 , n2957 );
    and g9518 ( n27675 , n4215 , n19870 );
    and g9519 ( n9549 , n25586 , n4199 );
    or g9520 ( n7234 , n4878 , n10281 );
    or g9521 ( n29795 , n2684 , n16659 );
    and g9522 ( n33694 , n6897 , n2752 );
    or g9523 ( n322 , n5472 , n12128 );
    or g9524 ( n13034 , n8432 , n21465 );
    or g9525 ( n32223 , n34053 , n19451 );
    or g9526 ( n23158 , n3455 , n9601 );
    and g9527 ( n21232 , n28321 , n34684 );
    not g9528 ( n13908 , n20621 );
    nor g9529 ( n2895 , n16620 , n11790 );
    nor g9530 ( n20513 , n1950 , n8418 );
    or g9531 ( n14627 , n1779 , n865 );
    not g9532 ( n25870 , n4896 );
    or g9533 ( n18984 , n31289 , n26568 );
    or g9534 ( n17254 , n29269 , n10900 );
    or g9535 ( n32563 , n22397 , n18357 );
    and g9536 ( n23930 , n2847 , n3648 );
    and g9537 ( n32930 , n29026 , n16412 );
    and g9538 ( n17713 , n9610 , n1114 );
    and g9539 ( n12230 , n17552 , n30552 );
    or g9540 ( n30168 , n35940 , n29872 );
    or g9541 ( n16218 , n2099 , n1397 );
    and g9542 ( n9437 , n15053 , n22831 );
    xnor g9543 ( n8611 , n25923 , n25219 );
    or g9544 ( n9526 , n22291 , n31558 );
    or g9545 ( n13871 , n31559 , n29278 );
    xnor g9546 ( n20556 , n27675 , n9793 );
    xnor g9547 ( n31178 , n9586 , n11681 );
    or g9548 ( n21682 , n7001 , n29633 );
    and g9549 ( n24435 , n951 , n15488 );
    or g9550 ( n11343 , n22291 , n24819 );
    or g9551 ( n10482 , n7880 , n25705 );
    or g9552 ( n25344 , n3813 , n10140 );
    or g9553 ( n5643 , n32857 , n29232 );
    xnor g9554 ( n22042 , n10164 , n25778 );
    and g9555 ( n24626 , n11198 , n31299 );
    xnor g9556 ( n24306 , n29253 , n822 );
    buf g9557 ( n27196 , n26610 );
    or g9558 ( n26536 , n32989 , n9930 );
    not g9559 ( n25078 , n25492 );
    or g9560 ( n10294 , n28148 , n9911 );
    or g9561 ( n13738 , n34455 , n15144 );
    or g9562 ( n16278 , n27995 , n20812 );
    and g9563 ( n19123 , n28567 , n13067 );
    xnor g9564 ( n21635 , n30559 , n11455 );
    and g9565 ( n6979 , n16124 , n2868 );
    or g9566 ( n20886 , n9793 , n33285 );
    xnor g9567 ( n10955 , n32304 , n11046 );
    xnor g9568 ( n20910 , n20592 , n31559 );
    and g9569 ( n8175 , n7247 , n16638 );
    and g9570 ( n1792 , n3262 , n30188 );
    and g9571 ( n20211 , n34384 , n20782 );
    or g9572 ( n26957 , n30152 , n14841 );
    and g9573 ( n31595 , n29043 , n33991 );
    or g9574 ( n23709 , n9463 , n11407 );
    or g9575 ( n1917 , n34716 , n25732 );
    or g9576 ( n14596 , n1358 , n13307 );
    or g9577 ( n23562 , n12490 , n9832 );
    nor g9578 ( n14601 , n33882 , n19128 );
    xnor g9579 ( n27498 , n25543 , n9658 );
    nor g9580 ( n20058 , n34728 , n4896 );
    nor g9581 ( n28813 , n11046 , n13097 );
    or g9582 ( n23321 , n21759 , n34484 );
    buf g9583 ( n4172 , n29872 );
    xnor g9584 ( n1702 , n24530 , n1341 );
    or g9585 ( n13295 , n15819 , n22783 );
    nor g9586 ( n19671 , n27431 , n10314 );
    xnor g9587 ( n28229 , n15860 , n15321 );
    xnor g9588 ( n25173 , n33190 , n27072 );
    and g9589 ( n14000 , n32506 , n26507 );
    or g9590 ( n31657 , n29884 , n918 );
    or g9591 ( n22214 , n29336 , n32152 );
    xnor g9592 ( n34710 , n18988 , n31232 );
    or g9593 ( n35341 , n4960 , n52 );
    or g9594 ( n4302 , n20166 , n18488 );
    or g9595 ( n23977 , n30521 , n8503 );
    or g9596 ( n1874 , n30707 , n2405 );
    or g9597 ( n28886 , n31629 , n7673 );
    xnor g9598 ( n26236 , n15143 , n5547 );
    or g9599 ( n23251 , n25244 , n24672 );
    and g9600 ( n28192 , n333 , n35606 );
    or g9601 ( n7867 , n5953 , n5509 );
    not g9602 ( n21413 , n10895 );
    or g9603 ( n14872 , n20325 , n12879 );
    xnor g9604 ( n10998 , n1890 , n11190 );
    xnor g9605 ( n3638 , n34747 , n13988 );
    xnor g9606 ( n26928 , n27863 , n10894 );
    or g9607 ( n10170 , n9139 , n10762 );
    or g9608 ( n32615 , n21845 , n18803 );
    or g9609 ( n23317 , n19489 , n5821 );
    or g9610 ( n20386 , n15299 , n33220 );
    not g9611 ( n13433 , n29713 );
    and g9612 ( n34975 , n14384 , n31113 );
    or g9613 ( n7539 , n9793 , n28798 );
    xnor g9614 ( n546 , n25711 , n33515 );
    and g9615 ( n14113 , n27259 , n17751 );
    xnor g9616 ( n8142 , n18734 , n29839 );
    or g9617 ( n25406 , n24978 , n32071 );
    xnor g9618 ( n30556 , n26501 , n13958 );
    xnor g9619 ( n34921 , n20656 , n7837 );
    or g9620 ( n4628 , n12231 , n17612 );
    nor g9621 ( n6452 , n17751 , n30467 );
    xnor g9622 ( n19398 , n1699 , n20502 );
    xnor g9623 ( n27319 , n19718 , n9793 );
    xnor g9624 ( n13729 , n19621 , n33889 );
    and g9625 ( n25061 , n11100 , n21415 );
    xnor g9626 ( n23430 , n9870 , n21481 );
    not g9627 ( n30039 , n21043 );
    nor g9628 ( n10309 , n14150 , n8827 );
    xnor g9629 ( n13502 , n11537 , n29839 );
    and g9630 ( n26106 , n26213 , n3013 );
    and g9631 ( n16831 , n20414 , n26298 );
    and g9632 ( n34168 , n9598 , n24987 );
    or g9633 ( n21455 , n27863 , n20812 );
    and g9634 ( n15363 , n31766 , n11189 );
    xnor g9635 ( n22489 , n11478 , n19984 );
    xnor g9636 ( n7976 , n2358 , n35541 );
    xnor g9637 ( n26667 , n14885 , n29839 );
    or g9638 ( n6948 , n30375 , n9951 );
    or g9639 ( n802 , n3021 , n29317 );
    and g9640 ( n15604 , n2343 , n22938 );
    and g9641 ( n5929 , n23668 , n31366 );
    nor g9642 ( n35529 , n11455 , n22159 );
    or g9643 ( n35636 , n4839 , n31134 );
    not g9644 ( n13421 , n28649 );
    and g9645 ( n28934 , n15532 , n6494 );
    xnor g9646 ( n22233 , n10260 , n27566 );
    and g9647 ( n23033 , n2003 , n21849 );
    not g9648 ( n26382 , n29522 );
    or g9649 ( n23318 , n28633 , n20601 );
    or g9650 ( n16653 , n22968 , n22858 );
    or g9651 ( n13510 , n19976 , n34865 );
    and g9652 ( n26423 , n18952 , n9227 );
    xnor g9653 ( n4783 , n33130 , n3871 );
    and g9654 ( n26458 , n4136 , n21491 );
    or g9655 ( n6919 , n28746 , n3756 );
    nor g9656 ( n2581 , n2838 , n4838 );
    or g9657 ( n25410 , n13083 , n19490 );
    or g9658 ( n12896 , n11855 , n24356 );
    and g9659 ( n5358 , n32365 , n18888 );
    or g9660 ( n2301 , n7171 , n34084 );
    and g9661 ( n30675 , n20578 , n25251 );
    or g9662 ( n1108 , n4288 , n9623 );
    and g9663 ( n1338 , n23595 , n9151 );
    xnor g9664 ( n27787 , n17869 , n25174 );
    or g9665 ( n25491 , n11802 , n34472 );
    and g9666 ( n32305 , n24498 , n2208 );
    nor g9667 ( n19243 , n7555 , n30610 );
    or g9668 ( n10859 , n11724 , n17964 );
    not g9669 ( n3940 , n29713 );
    or g9670 ( n14015 , n17495 , n31055 );
    xnor g9671 ( n7004 , n32404 , n18554 );
    and g9672 ( n32215 , n35651 , n12094 );
    or g9673 ( n9889 , n2281 , n31062 );
    and g9674 ( n15831 , n13347 , n14624 );
    xnor g9675 ( n34057 , n29969 , n32198 );
    and g9676 ( n19975 , n10036 , n18530 );
    or g9677 ( n9801 , n30070 , n24489 );
    or g9678 ( n22949 , n13457 , n12950 );
    xnor g9679 ( n27933 , n5582 , n31656 );
    or g9680 ( n29605 , n32095 , n1745 );
    nor g9681 ( n26060 , n35927 , n33582 );
    and g9682 ( n4170 , n300 , n7152 );
    and g9683 ( n19755 , n31763 , n18617 );
    or g9684 ( n7493 , n8236 , n11996 );
    or g9685 ( n24297 , n14630 , n12428 );
    and g9686 ( n16219 , n30378 , n7459 );
    or g9687 ( n22688 , n24086 , n20579 );
    or g9688 ( n11057 , n22234 , n11258 );
    and g9689 ( n25172 , n2350 , n17494 );
    or g9690 ( n25093 , n33645 , n24172 );
    or g9691 ( n11526 , n27130 , n10289 );
    not g9692 ( n27582 , n3357 );
    nor g9693 ( n5968 , n32500 , n13245 );
    or g9694 ( n25056 , n24371 , n26321 );
    or g9695 ( n26102 , n24371 , n22413 );
    or g9696 ( n31669 , n6475 , n31464 );
    and g9697 ( n21611 , n28538 , n18960 );
    or g9698 ( n18721 , n4882 , n513 );
    and g9699 ( n35591 , n1621 , n28006 );
    and g9700 ( n29248 , n25689 , n1137 );
    or g9701 ( n30590 , n31461 , n30708 );
    nor g9702 ( n27936 , n3676 , n9921 );
    and g9703 ( n17270 , n24558 , n19222 );
    or g9704 ( n28300 , n3914 , n32959 );
    or g9705 ( n33798 , n24332 , n35190 );
    buf g9706 ( n14918 , n19385 );
    not g9707 ( n29417 , n11529 );
    or g9708 ( n32768 , n7320 , n33850 );
    or g9709 ( n9406 , n26631 , n8153 );
    not g9710 ( n1753 , n34926 );
    or g9711 ( n18894 , n13745 , n35143 );
    nor g9712 ( n27533 , n17568 , n11747 );
    or g9713 ( n24110 , n27532 , n25863 );
    or g9714 ( n12063 , n18102 , n18512 );
    and g9715 ( n33220 , n4794 , n28576 );
    and g9716 ( n34289 , n30426 , n29507 );
    or g9717 ( n2481 , n4962 , n25066 );
    nor g9718 ( n10379 , n13029 , n26282 );
    or g9719 ( n16574 , n21297 , n4595 );
    and g9720 ( n9108 , n34870 , n32596 );
    or g9721 ( n23679 , n14718 , n25255 );
    or g9722 ( n32566 , n1740 , n18255 );
    xnor g9723 ( n21722 , n19284 , n24371 );
    and g9724 ( n4264 , n5205 , n28925 );
    xnor g9725 ( n34668 , n4662 , n29713 );
    or g9726 ( n12099 , n25746 , n16409 );
    or g9727 ( n15643 , n27800 , n21042 );
    and g9728 ( n34660 , n7066 , n26854 );
    xnor g9729 ( n22400 , n30146 , n32857 );
    xnor g9730 ( n29756 , n18012 , n15663 );
    or g9731 ( n21649 , n26521 , n2241 );
    and g9732 ( n34604 , n19638 , n9803 );
    xnor g9733 ( n35219 , n16495 , n1605 );
    or g9734 ( n15087 , n29395 , n22501 );
    or g9735 ( n4866 , n12735 , n30780 );
    and g9736 ( n4956 , n14546 , n2605 );
    xnor g9737 ( n16206 , n19694 , n31799 );
    or g9738 ( n27045 , n21709 , n23323 );
    xnor g9739 ( n16446 , n11885 , n8815 );
    nor g9740 ( n32938 , n1950 , n7702 );
    nor g9741 ( n18338 , n4960 , n22798 );
    or g9742 ( n14936 , n8125 , n26220 );
    or g9743 ( n18138 , n6911 , n7038 );
    or g9744 ( n35011 , n24478 , n10960 );
    and g9745 ( n20747 , n19719 , n27654 );
    and g9746 ( n26393 , n7626 , n10305 );
    or g9747 ( n11754 , n9183 , n22946 );
    and g9748 ( n27305 , n19799 , n12372 );
    xnor g9749 ( n31219 , n18870 , n19441 );
    or g9750 ( n3145 , n32604 , n20836 );
    and g9751 ( n4446 , n28764 , n31470 );
    and g9752 ( n12621 , n28038 , n3531 );
    or g9753 ( n8322 , n19045 , n8956 );
    or g9754 ( n18645 , n6763 , n6216 );
    or g9755 ( n3776 , n30829 , n33720 );
    or g9756 ( n23609 , n15419 , n6374 );
    or g9757 ( n28339 , n6719 , n4057 );
    and g9758 ( n22328 , n26950 , n22291 );
    not g9759 ( n5521 , n35422 );
    or g9760 ( n21412 , n25174 , n16915 );
    or g9761 ( n35240 , n33932 , n18676 );
    xor g9762 ( n24478 , n14420 , n10210 );
    or g9763 ( n31607 , n35732 , n28240 );
    xnor g9764 ( n19906 , n161 , n31243 );
    or g9765 ( n4615 , n7654 , n11593 );
    nor g9766 ( n8541 , n19214 , n2119 );
    not g9767 ( n19297 , n4467 );
    not g9768 ( n30932 , n14468 );
    not g9769 ( n22502 , n35256 );
    xnor g9770 ( n20356 , n27662 , n33014 );
    or g9771 ( n4441 , n5287 , n31356 );
    or g9772 ( n20617 , n30385 , n22215 );
    xnor g9773 ( n35652 , n16432 , n774 );
    or g9774 ( n30997 , n21815 , n35422 );
    nor g9775 ( n30549 , n20567 , n1574 );
    xnor g9776 ( n3372 , n11911 , n677 );
    and g9777 ( n2998 , n30245 , n24227 );
    or g9778 ( n23865 , n32715 , n12217 );
    or g9779 ( n4473 , n11455 , n34842 );
    or g9780 ( n23561 , n18030 , n32505 );
    and g9781 ( n11074 , n35512 , n22104 );
    xnor g9782 ( n15606 , n10155 , n20292 );
    xnor g9783 ( n35260 , n18149 , n25914 );
    or g9784 ( n32757 , n4310 , n23825 );
    or g9785 ( n18783 , n16827 , n16285 );
    or g9786 ( n20483 , n16381 , n14699 );
    and g9787 ( n27943 , n24803 , n22733 );
    xnor g9788 ( n28752 , n17127 , n23604 );
    or g9789 ( n652 , n16689 , n5482 );
    or g9790 ( n17381 , n23857 , n20375 );
    or g9791 ( n21250 , n16186 , n16659 );
    not g9792 ( n24287 , n22471 );
    nor g9793 ( n23968 , n23604 , n24082 );
    or g9794 ( n27857 , n4974 , n5891 );
    and g9795 ( n9036 , n23533 , n2545 );
    not g9796 ( n24247 , n25354 );
    xnor g9797 ( n25973 , n5520 , n28933 );
    or g9798 ( n7849 , n3837 , n15117 );
    or g9799 ( n7609 , n3923 , n18477 );
    or g9800 ( n27986 , n30554 , n30826 );
    and g9801 ( n9999 , n2231 , n18035 );
    xnor g9802 ( n8151 , n15183 , n7163 );
    or g9803 ( n13962 , n9793 , n11617 );
    or g9804 ( n35678 , n29273 , n763 );
    xnor g9805 ( n6787 , n22539 , n29231 );
    or g9806 ( n30137 , n22217 , n12344 );
    not g9807 ( n27159 , n1543 );
    or g9808 ( n32779 , n31114 , n19084 );
    or g9809 ( n6485 , n19040 , n35665 );
    and g9810 ( n2511 , n16063 , n20522 );
    not g9811 ( n7474 , n15886 );
    or g9812 ( n27877 , n10714 , n21002 );
    not g9813 ( n12764 , n32857 );
    or g9814 ( n27732 , n19993 , n27551 );
    and g9815 ( n19166 , n30455 , n886 );
    and g9816 ( n12133 , n28028 , n315 );
    or g9817 ( n18 , n1503 , n2303 );
    not g9818 ( n20734 , n7857 );
    nor g9819 ( n920 , n21645 , n16762 );
    nor g9820 ( n29056 , n31215 , n29800 );
    nor g9821 ( n18573 , n32715 , n1117 );
    and g9822 ( n30650 , n35708 , n9789 );
    or g9823 ( n18553 , n17416 , n18264 );
    or g9824 ( n11976 , n16840 , n35393 );
    xnor g9825 ( n16882 , n22540 , n11499 );
    or g9826 ( n27449 , n34488 , n1407 );
    or g9827 ( n25653 , n32857 , n26615 );
    or g9828 ( n11024 , n19322 , n19125 );
    and g9829 ( n29459 , n33700 , n14657 );
    not g9830 ( n1171 , n12428 );
    or g9831 ( n14227 , n15273 , n36003 );
    and g9832 ( n25603 , n10582 , n29671 );
    or g9833 ( n24738 , n14864 , n20300 );
    or g9834 ( n31890 , n29475 , n20559 );
    nor g9835 ( n33296 , n22291 , n13544 );
    and g9836 ( n12203 , n13424 , n3089 );
    and g9837 ( n12910 , n7724 , n12620 );
    and g9838 ( n5800 , n25906 , n17397 );
    or g9839 ( n7226 , n14484 , n30826 );
    nor g9840 ( n34982 , n25602 , n31651 );
    xnor g9841 ( n12440 , n1503 , n2303 );
    xnor g9842 ( n22527 , n2216 , n11046 );
    and g9843 ( n24383 , n14952 , n27672 );
    xnor g9844 ( n18076 , n25992 , n9496 );
    or g9845 ( n16743 , n7836 , n26002 );
    and g9846 ( n11570 , n14104 , n14738 );
    xnor g9847 ( n33879 , n19278 , n24028 );
    xnor g9848 ( n20376 , n298 , n33951 );
    buf g9849 ( n19421 , n19385 );
    or g9850 ( n29840 , n23591 , n139 );
    nor g9851 ( n23486 , n21663 , n31411 );
    or g9852 ( n32454 , n15740 , n26112 );
    xnor g9853 ( n13803 , n12696 , n15621 );
    and g9854 ( n22027 , n18570 , n13874 );
    not g9855 ( n18660 , n12173 );
    or g9856 ( n13855 , n16103 , n35535 );
    not g9857 ( n729 , n1950 );
    and g9858 ( n194 , n15694 , n29688 );
    xnor g9859 ( n35803 , n35936 , n8885 );
    or g9860 ( n27818 , n31210 , n31048 );
    not g9861 ( n3681 , n6075 );
    not g9862 ( n27126 , n13408 );
    or g9863 ( n31653 , n31548 , n2270 );
    and g9864 ( n23546 , n31262 , n6443 );
    xnor g9865 ( n7378 , n29306 , n18267 );
    and g9866 ( n4914 , n19101 , n23388 );
    or g9867 ( n4126 , n3654 , n3906 );
    or g9868 ( n9569 , n15480 , n4742 );
    and g9869 ( n14703 , n23103 , n4053 );
    xnor g9870 ( n20158 , n15820 , n27226 );
    and g9871 ( n5733 , n32128 , n17475 );
    or g9872 ( n26831 , n13710 , n21937 );
    not g9873 ( n21819 , n25602 );
    and g9874 ( n33808 , n15668 , n16190 );
    and g9875 ( n1118 , n9646 , n1724 );
    or g9876 ( n34780 , n17702 , n28123 );
    and g9877 ( n27158 , n2944 , n16908 );
    and g9878 ( n27997 , n10719 , n31111 );
    or g9879 ( n21694 , n4962 , n34205 );
    not g9880 ( n31996 , n31236 );
    not g9881 ( n9847 , n29378 );
    xnor g9882 ( n25975 , n1440 , n24789 );
    and g9883 ( n6183 , n34442 , n14454 );
    and g9884 ( n14708 , n17334 , n24736 );
    xnor g9885 ( n5218 , n16288 , n29713 );
    not g9886 ( n30162 , n26482 );
    and g9887 ( n20126 , n31476 , n15446 );
    and g9888 ( n27288 , n24448 , n12444 );
    and g9889 ( n1256 , n28749 , n10835 );
    xnor g9890 ( n1939 , n18633 , n25602 );
    not g9891 ( n16262 , n6592 );
    or g9892 ( n27440 , n13467 , n1105 );
    xnor g9893 ( n10981 , n5488 , n9789 );
    or g9894 ( n13249 , n35927 , n4911 );
    nor g9895 ( n10524 , n17702 , n5216 );
    xnor g9896 ( n19611 , n29782 , n26736 );
    not g9897 ( n16709 , n6199 );
    xnor g9898 ( n2911 , n1338 , n1950 );
    or g9899 ( n7165 , n361 , n28668 );
    or g9900 ( n25134 , n5095 , n13305 );
    not g9901 ( n23769 , n32095 );
    and g9902 ( n23972 , n19008 , n30137 );
    and g9903 ( n14043 , n32602 , n33008 );
    or g9904 ( n8506 , n14325 , n2168 );
    or g9905 ( n30121 , n34049 , n25648 );
    xnor g9906 ( n12574 , n30084 , n23604 );
    or g9907 ( n4109 , n17934 , n22550 );
    or g9908 ( n12180 , n24948 , n35693 );
    nor g9909 ( n29355 , n3205 , n18718 );
    or g9910 ( n31119 , n9347 , n17111 );
    xnor g9911 ( n13 , n32500 , n15886 );
    not g9912 ( n8357 , n1091 );
    nor g9913 ( n25683 , n35523 , n16501 );
    or g9914 ( n21043 , n14747 , n20070 );
    or g9915 ( n3797 , n20863 , n18385 );
    xnor g9916 ( n21275 , n4213 , n9789 );
    not g9917 ( n20738 , n9163 );
    or g9918 ( n16513 , n29518 , n19125 );
    xnor g9919 ( n16891 , n33902 , n4962 );
    or g9920 ( n35352 , n33734 , n25592 );
    xnor g9921 ( n1089 , n14767 , n27794 );
    nor g9922 ( n32726 , n17568 , n5877 );
    or g9923 ( n5016 , n28415 , n11850 );
    and g9924 ( n25575 , n9216 , n14026 );
    xnor g9925 ( n28348 , n22503 , n14845 );
    xnor g9926 ( n27605 , n13575 , n6936 );
    and g9927 ( n785 , n33721 , n22329 );
    or g9928 ( n19746 , n29436 , n25247 );
    and g9929 ( n31333 , n34257 , n17377 );
    and g9930 ( n23040 , n20635 , n25485 );
    or g9931 ( n11154 , n24332 , n20462 );
    or g9932 ( n33225 , n18738 , n21691 );
    not g9933 ( n5637 , n21658 );
    or g9934 ( n19365 , n19624 , n28324 );
    and g9935 ( n26969 , n35159 , n16374 );
    or g9936 ( n700 , n12502 , n4912 );
    and g9937 ( n12262 , n9263 , n28682 );
    and g9938 ( n15025 , n19481 , n25620 );
    not g9939 ( n30372 , n14079 );
    and g9940 ( n22051 , n23785 , n11945 );
    or g9941 ( n22059 , n4878 , n1088 );
    or g9942 ( n9635 , n31481 , n23209 );
    not g9943 ( n9278 , n16620 );
    xnor g9944 ( n5606 , n20050 , n1815 );
    or g9945 ( n29412 , n33947 , n34484 );
    xnor g9946 ( n20818 , n2222 , n27291 );
    and g9947 ( n19977 , n12420 , n21283 );
    and g9948 ( n20406 , n20390 , n3482 );
    or g9949 ( n7154 , n31215 , n4604 );
    or g9950 ( n18176 , n10364 , n7090 );
    and g9951 ( n9385 , n12552 , n24456 );
    and g9952 ( n32538 , n20151 , n9299 );
    or g9953 ( n6227 , n30588 , n13760 );
    nor g9954 ( n17070 , n27755 , n13193 );
    nor g9955 ( n18098 , n31799 , n30337 );
    and g9956 ( n15727 , n14825 , n13996 );
    xnor g9957 ( n21874 , n24534 , n11046 );
    or g9958 ( n19008 , n26802 , n3274 );
    or g9959 ( n6432 , n2986 , n4595 );
    or g9960 ( n3361 , n31420 , n26865 );
    or g9961 ( n34825 , n28445 , n34727 );
    or g9962 ( n21967 , n18893 , n28613 );
    xnor g9963 ( n33115 , n13392 , n16620 );
    not g9964 ( n18286 , n23108 );
    or g9965 ( n17903 , n30435 , n3842 );
    or g9966 ( n3022 , n25862 , n14441 );
    or g9967 ( n12761 , n21159 , n9731 );
    not g9968 ( n16064 , n4874 );
    or g9969 ( n428 , n27109 , n1371 );
    or g9970 ( n26796 , n11889 , n4363 );
    not g9971 ( n29378 , n16611 );
    or g9972 ( n22265 , n4962 , n16632 );
    xnor g9973 ( n35144 , n35446 , n5320 );
    and g9974 ( n26770 , n19030 , n30606 );
    not g9975 ( n8377 , n16620 );
    or g9976 ( n5136 , n6735 , n27447 );
    xnor g9977 ( n26359 , n34514 , n1826 );
    not g9978 ( n15153 , n6690 );
    not g9979 ( n3020 , n9894 );
    xnor g9980 ( n768 , n25900 , n14100 );
    nor g9981 ( n7314 , n19551 , n7342 );
    xnor g9982 ( n28354 , n29173 , n30083 );
    xnor g9983 ( n10888 , n33195 , n23852 );
    or g9984 ( n25796 , n34900 , n32505 );
    or g9985 ( n6270 , n7091 , n33649 );
    or g9986 ( n29042 , n32418 , n4488 );
    and g9987 ( n152 , n15089 , n14309 );
    nor g9988 ( n4560 , n16620 , n31436 );
    xnor g9989 ( n19415 , n4634 , n23544 );
    or g9990 ( n1589 , n27195 , n25773 );
    not g9991 ( n3627 , n35927 );
    or g9992 ( n16787 , n16836 , n19933 );
    or g9993 ( n28459 , n25045 , n16762 );
    xnor g9994 ( n35921 , n20336 , n25174 );
    xnor g9995 ( n22057 , n7973 , n32929 );
    xnor g9996 ( n9720 , n35398 , n13648 );
    nor g9997 ( n15099 , n16664 , n13898 );
    or g9998 ( n14760 , n6254 , n35393 );
    and g9999 ( n18964 , n21427 , n17904 );
    xnor g10000 ( n31821 , n22702 , n29107 );
    or g10001 ( n20903 , n17986 , n20579 );
    and g10002 ( n32531 , n1036 , n24174 );
    or g10003 ( n10677 , n25543 , n25355 );
    and g10004 ( n33063 , n2871 , n27946 );
    or g10005 ( n15797 , n24430 , n25594 );
    or g10006 ( n22404 , n10894 , n14379 );
    or g10007 ( n12862 , n27602 , n9672 );
    or g10008 ( n3559 , n27742 , n19421 );
    or g10009 ( n13529 , n27921 , n5184 );
    not g10010 ( n27172 , n30459 );
    and g10011 ( n9449 , n16635 , n2419 );
    xnor g10012 ( n20837 , n19106 , n33622 );
    xnor g10013 ( n10506 , n18430 , n30413 );
    and g10014 ( n34756 , n9167 , n4964 );
    or g10015 ( n28514 , n24862 , n14839 );
    or g10016 ( n25001 , n14978 , n2524 );
    and g10017 ( n528 , n15810 , n4602 );
    or g10018 ( n8942 , n14696 , n14918 );
    or g10019 ( n26370 , n14019 , n28548 );
    xnor g10020 ( n6230 , n24361 , n2492 );
    xnor g10021 ( n34545 , n14990 , n9793 );
    or g10022 ( n18800 , n16284 , n7673 );
    or g10023 ( n33900 , n10285 , n17125 );
    and g10024 ( n7003 , n24232 , n32996 );
    or g10025 ( n15010 , n1596 , n9092 );
    or g10026 ( n30532 , n7714 , n6479 );
    xnor g10027 ( n102 , n9383 , n17108 );
    and g10028 ( n24095 , n28870 , n12064 );
    not g10029 ( n32371 , n5096 );
    not g10030 ( n34025 , n15886 );
    xnor g10031 ( n33309 , n4365 , n22823 );
    xnor g10032 ( n12573 , n18973 , n3691 );
    xor g10033 ( n24342 , n8447 , n10256 );
    and g10034 ( n2854 , n32946 , n3661 );
    xnor g10035 ( n33598 , n7733 , n4758 );
    or g10036 ( n10735 , n31986 , n25594 );
    and g10037 ( n33875 , n6335 , n15443 );
    xnor g10038 ( n26819 , n5052 , n4288 );
    or g10039 ( n25743 , n5048 , n30204 );
    not g10040 ( n33328 , n1950 );
    xnor g10041 ( n2886 , n19099 , n25381 );
    or g10042 ( n14317 , n17652 , n8831 );
    and g10043 ( n24582 , n31365 , n30170 );
    or g10044 ( n6887 , n28096 , n14699 );
    nor g10045 ( n21145 , n9401 , n19218 );
    and g10046 ( n27203 , n7781 , n23277 );
    not g10047 ( n35151 , n11046 );
    or g10048 ( n30249 , n13446 , n23921 );
    or g10049 ( n34730 , n16620 , n8182 );
    xnor g10050 ( n20372 , n8930 , n36021 );
    or g10051 ( n18916 , n28173 , n32379 );
    nor g10052 ( n22634 , n26550 , n30456 );
    xnor g10053 ( n28709 , n2931 , n3627 );
    nor g10054 ( n26664 , n2865 , n16649 );
    or g10055 ( n35838 , n14236 , n12693 );
    and g10056 ( n21703 , n33078 , n663 );
    not g10057 ( n13926 , n14143 );
    or g10058 ( n3664 , n4817 , n9998 );
    or g10059 ( n5083 , n4962 , n14728 );
    xnor g10060 ( n17026 , n14688 , n10894 );
    and g10061 ( n8719 , n9314 , n25576 );
    and g10062 ( n20785 , n28084 , n18799 );
    or g10063 ( n33987 , n1806 , n6945 );
    and g10064 ( n6936 , n18351 , n3175 );
    or g10065 ( n20265 , n29790 , n2701 );
    or g10066 ( n7106 , n29736 , n21332 );
    or g10067 ( n757 , n31799 , n24920 );
    or g10068 ( n6223 , n4973 , n10749 );
    and g10069 ( n34243 , n29460 , n26513 );
    and g10070 ( n14414 , n28845 , n8228 );
    and g10071 ( n20773 , n2388 , n29950 );
    and g10072 ( n15959 , n33306 , n12720 );
    and g10073 ( n7881 , n31791 , n31567 );
    and g10074 ( n26862 , n3472 , n16857 );
    buf g10075 ( n26292 , n11518 );
    nor g10076 ( n23652 , n32857 , n16805 );
    or g10077 ( n19626 , n13971 , n25255 );
    or g10078 ( n24835 , n28224 , n28190 );
    xnor g10079 ( n6247 , n23369 , n15886 );
    nor g10080 ( n30279 , n3205 , n14959 );
    or g10081 ( n16358 , n23276 , n27574 );
    or g10082 ( n20544 , n32275 , n2712 );
    and g10083 ( n4305 , n2588 , n14260 );
    nor g10084 ( n5980 , n7300 , n5780 );
    nor g10085 ( n2744 , n3222 , n12816 );
    not g10086 ( n16636 , n9793 );
    or g10087 ( n12880 , n27844 , n10336 );
    or g10088 ( n1716 , n25602 , n14786 );
    xnor g10089 ( n1855 , n3316 , n35927 );
    and g10090 ( n2077 , n12730 , n15203 );
    not g10091 ( n10382 , n26209 );
    xnor g10092 ( n13527 , n7342 , n19551 );
    or g10093 ( n1395 , n33945 , n31577 );
    or g10094 ( n23765 , n4878 , n5533 );
    not g10095 ( n1596 , n1052 );
    buf g10096 ( n14706 , n2092 );
    or g10097 ( n25230 , n20084 , n34865 );
    xnor g10098 ( n25151 , n16258 , n30028 );
    nor g10099 ( n15207 , n31800 , n9921 );
    or g10100 ( n10815 , n8841 , n17068 );
    or g10101 ( n34102 , n24104 , n21862 );
    nor g10102 ( n11722 , n15886 , n29363 );
    nor g10103 ( n2198 , n25811 , n22738 );
    or g10104 ( n15762 , n21844 , n1386 );
    and g10105 ( n7651 , n14062 , n32886 );
    or g10106 ( n7638 , n12331 , n25447 );
    xnor g10107 ( n8462 , n9902 , n26395 );
    not g10108 ( n11263 , n1217 );
    or g10109 ( n1078 , n2637 , n22359 );
    and g10110 ( n25735 , n2491 , n30186 );
    or g10111 ( n21100 , n31447 , n17120 );
    or g10112 ( n7735 , n4685 , n19722 );
    and g10113 ( n12358 , n31408 , n14162 );
    or g10114 ( n7949 , n8577 , n628 );
    xnor g10115 ( n29242 , n34795 , n23847 );
    xnor g10116 ( n6885 , n35120 , n29388 );
    or g10117 ( n7083 , n21892 , n10066 );
    or g10118 ( n601 , n19359 , n27266 );
    or g10119 ( n11596 , n11598 , n21742 );
    xnor g10120 ( n28744 , n5687 , n1158 );
    not g10121 ( n10587 , n19551 );
    and g10122 ( n18534 , n33477 , n27423 );
    and g10123 ( n20147 , n28625 , n766 );
    not g10124 ( n27917 , n31056 );
    nor g10125 ( n29588 , n26656 , n29907 );
    buf g10126 ( n4595 , n29176 );
    or g10127 ( n9262 , n22243 , n20055 );
    not g10128 ( n33767 , n15886 );
    and g10129 ( n24170 , n26534 , n22812 );
    or g10130 ( n17493 , n22923 , n18593 );
    or g10131 ( n6049 , n11870 , n3517 );
    not g10132 ( n34679 , n17804 );
    not g10133 ( n20330 , n33948 );
    and g10134 ( n31307 , n26874 , n27519 );
    nor g10135 ( n28498 , n16620 , n5110 );
    and g10136 ( n6191 , n18817 , n29566 );
    not g10137 ( n34015 , n12434 );
    xnor g10138 ( n29844 , n6595 , n1048 );
    or g10139 ( n21131 , n1819 , n7240 );
    xnor g10140 ( n27020 , n33770 , n7656 );
    xnor g10141 ( n33324 , n30629 , n34744 );
    and g10142 ( n35519 , n4489 , n32420 );
    or g10143 ( n26893 , n9688 , n21042 );
    or g10144 ( n29582 , n1514 , n10872 );
    xnor g10145 ( n30566 , n4316 , n25602 );
    and g10146 ( n15321 , n34106 , n9988 );
    xnor g10147 ( n9421 , n11257 , n32917 );
    not g10148 ( n25686 , n9793 );
    or g10149 ( n3509 , n24754 , n15805 );
    and g10150 ( n25264 , n27128 , n17414 );
    and g10151 ( n29497 , n3811 , n35956 );
    or g10152 ( n31889 , n3978 , n1402 );
    and g10153 ( n813 , n27076 , n6391 );
    and g10154 ( n7306 , n17678 , n8326 );
    and g10155 ( n7399 , n34206 , n10254 );
    xnor g10156 ( n32027 , n27717 , n35540 );
    xnor g10157 ( n3739 , n10010 , n35927 );
    xnor g10158 ( n10093 , n30385 , n22215 );
    xnor g10159 ( n16737 , n34398 , n5287 );
    nor g10160 ( n22299 , n17568 , n32190 );
    or g10161 ( n15564 , n27575 , n32517 );
    or g10162 ( n2568 , n9568 , n18808 );
    xnor g10163 ( n15111 , n18403 , n22291 );
    and g10164 ( n22293 , n36004 , n28618 );
    or g10165 ( n25635 , n27291 , n18935 );
    and g10166 ( n21880 , n6429 , n23588 );
    not g10167 ( n35417 , n16223 );
    or g10168 ( n17147 , n22881 , n27201 );
    or g10169 ( n22424 , n1353 , n3756 );
    and g10170 ( n32917 , n21534 , n14707 );
    not g10171 ( n33990 , n4519 );
    and g10172 ( n19720 , n15193 , n13766 );
    and g10173 ( n10583 , n20121 , n20276 );
    or g10174 ( n5842 , n2750 , n13023 );
    xnor g10175 ( n30786 , n3927 , n3518 );
    xnor g10176 ( n33550 , n28397 , n3205 );
    or g10177 ( n471 , n30221 , n2422 );
    and g10178 ( n5516 , n28177 , n18657 );
    or g10179 ( n2229 , n30302 , n13099 );
    nor g10180 ( n9101 , n30133 , n18115 );
    or g10181 ( n33425 , n9793 , n2794 );
    xnor g10182 ( n16798 , n4258 , n32857 );
    nor g10183 ( n28120 , n10387 , n23921 );
    xnor g10184 ( n16852 , n35773 , n4364 );
    or g10185 ( n1772 , n30343 , n544 );
    xnor g10186 ( n26762 , n23241 , n29713 );
    and g10187 ( n19860 , n10686 , n16614 );
    or g10188 ( n20648 , n30835 , n20690 );
    or g10189 ( n534 , n26323 , n24204 );
    and g10190 ( n2622 , n331 , n6214 );
    or g10191 ( n27861 , n3946 , n30485 );
    or g10192 ( n10049 , n24963 , n22316 );
    or g10193 ( n14346 , n31559 , n6703 );
    or g10194 ( n2145 , n31799 , n9161 );
    xnor g10195 ( n23108 , n2878 , n11046 );
    or g10196 ( n34253 , n12535 , n1079 );
    nor g10197 ( n15438 , n11182 , n10265 );
    or g10198 ( n20315 , n30727 , n35757 );
    nor g10199 ( n12194 , n33068 , n35643 );
    xnor g10200 ( n30848 , n17151 , n28510 );
    or g10201 ( n35807 , n1087 , n25355 );
    not g10202 ( n22548 , n22980 );
    xnor g10203 ( n11675 , n32069 , n6079 );
    not g10204 ( n28748 , n26259 );
    xnor g10205 ( n14753 , n29730 , n34717 );
    or g10206 ( n6587 , n9718 , n18855 );
    xnor g10207 ( n10984 , n3522 , n35164 );
    or g10208 ( n32320 , n20666 , n27592 );
    and g10209 ( n32912 , n12156 , n22461 );
    xnor g10210 ( n15527 , n6999 , n27715 );
    or g10211 ( n32631 , n14797 , n20091 );
    or g10212 ( n24718 , n30492 , n32425 );
    xnor g10213 ( n21389 , n4122 , n7692 );
    or g10214 ( n20893 , n17592 , n2851 );
    nor g10215 ( n22398 , n16922 , n5493 );
    nor g10216 ( n8330 , n30366 , n16649 );
    or g10217 ( n11682 , n12249 , n12428 );
    or g10218 ( n4846 , n3014 , n5546 );
    or g10219 ( n13551 , n23307 , n20074 );
    xnor g10220 ( n30594 , n23020 , n11190 );
    xnor g10221 ( n7612 , n18321 , n15403 );
    or g10222 ( n2317 , n13413 , n9352 );
    or g10223 ( n29521 , n1453 , n10383 );
    xnor g10224 ( n15926 , n17356 , n11046 );
    nor g10225 ( n26611 , n10894 , n8313 );
    xnor g10226 ( n942 , n24550 , n1950 );
    and g10227 ( n4013 , n26536 , n27119 );
    or g10228 ( n68 , n25642 , n23462 );
    xnor g10229 ( n18756 , n5917 , n3222 );
    or g10230 ( n34330 , n35398 , n13648 );
    and g10231 ( n23010 , n17275 , n25391 );
    and g10232 ( n11728 , n29757 , n13742 );
    or g10233 ( n1246 , n25238 , n32362 );
    nor g10234 ( n22977 , n26038 , n30989 );
    or g10235 ( n28149 , n12971 , n16464 );
    or g10236 ( n8812 , n23834 , n36000 );
    or g10237 ( n24428 , n5533 , n15497 );
    and g10238 ( n34463 , n18440 , n14034 );
    or g10239 ( n9263 , n20265 , n35629 );
    or g10240 ( n6957 , n19551 , n4807 );
    and g10241 ( n26008 , n21416 , n35073 );
    or g10242 ( n32598 , n31120 , n26265 );
    not g10243 ( n31557 , n8278 );
    xnor g10244 ( n18870 , n31453 , n8432 );
    xnor g10245 ( n27653 , n1427 , n1922 );
    buf g10246 ( n24505 , n16649 );
    not g10247 ( n27650 , n30151 );
    xnor g10248 ( n8927 , n1698 , n15828 );
    or g10249 ( n4617 , n15565 , n16961 );
    or g10250 ( n6 , n7100 , n11295 );
    not g10251 ( n6554 , n26112 );
    and g10252 ( n29617 , n3576 , n15555 );
    and g10253 ( n1538 , n19724 , n3268 );
    or g10254 ( n6838 , n33787 , n18665 );
    or g10255 ( n6214 , n22007 , n4448 );
    or g10256 ( n2239 , n17902 , n27501 );
    or g10257 ( n5809 , n18561 , n3241 );
    xnor g10258 ( n8085 , n23151 , n3611 );
    xnor g10259 ( n33528 , n30434 , n16922 );
    or g10260 ( n16675 , n9738 , n18938 );
    or g10261 ( n26599 , n27596 , n2745 );
    or g10262 ( n25225 , n30004 , n23462 );
    or g10263 ( n4448 , n17454 , n12596 );
    and g10264 ( n10809 , n960 , n10584 );
    or g10265 ( n29785 , n25544 , n27704 );
    nor g10266 ( n29635 , n31799 , n5625 );
    and g10267 ( n17878 , n17963 , n7456 );
    and g10268 ( n23402 , n9602 , n10173 );
    or g10269 ( n10554 , n28820 , n22996 );
    not g10270 ( n21671 , n22797 );
    buf g10271 ( n31055 , n19939 );
    or g10272 ( n13711 , n1421 , n21956 );
    or g10273 ( n27556 , n2713 , n17068 );
    not g10274 ( n22361 , n25687 );
    or g10275 ( n10906 , n25460 , n9113 );
    xnor g10276 ( n11693 , n12678 , n16922 );
    or g10277 ( n32659 , n496 , n30732 );
    or g10278 ( n28179 , n7586 , n32634 );
    xnor g10279 ( n34924 , n1633 , n351 );
    xnor g10280 ( n21430 , n23068 , n31799 );
    buf g10281 ( n20427 , n33204 );
    not g10282 ( n5411 , n19754 );
    and g10283 ( n4637 , n3329 , n8699 );
    or g10284 ( n35873 , n13322 , n9036 );
    xnor g10285 ( n5562 , n7559 , n10107 );
    xnor g10286 ( n7219 , n7704 , n13924 );
    and g10287 ( n3340 , n20673 , n34446 );
    or g10288 ( n5329 , n22766 , n22946 );
    or g10289 ( n3967 , n2222 , n17354 );
    xnor g10290 ( n32192 , n17324 , n9789 );
    or g10291 ( n1283 , n20146 , n8090 );
    or g10292 ( n11260 , n24946 , n3314 );
    and g10293 ( n9118 , n5375 , n3792 );
    nor g10294 ( n14679 , n33738 , n34782 );
    xnor g10295 ( n27594 , n35089 , n3222 );
    nor g10296 ( n25334 , n33041 , n24899 );
    not g10297 ( n3101 , n12245 );
    or g10298 ( n26683 , n12638 , n14517 );
    and g10299 ( n2225 , n20193 , n4655 );
    and g10300 ( n4715 , n29289 , n24825 );
    not g10301 ( n32649 , n3205 );
    xor g10302 ( n9834 , n25451 , n1883 );
    or g10303 ( n12998 , n7564 , n21002 );
    or g10304 ( n2084 , n14209 , n2479 );
    and g10305 ( n28834 , n11112 , n23778 );
    and g10306 ( n19659 , n1499 , n11585 );
    or g10307 ( n22915 , n27940 , n3508 );
    or g10308 ( n12854 , n19975 , n27053 );
    xor g10309 ( n1680 , n12811 , n3255 );
    not g10310 ( n33629 , n31559 );
    or g10311 ( n13585 , n30040 , n35402 );
    or g10312 ( n33624 , n15976 , n12596 );
    and g10313 ( n9367 , n31410 , n21724 );
    or g10314 ( n35817 , n28123 , n22583 );
    xnor g10315 ( n3590 , n23843 , n31799 );
    nor g10316 ( n7608 , n31289 , n26474 );
    xnor g10317 ( n31925 , n13229 , n23219 );
    buf g10318 ( n5208 , n6288 );
    or g10319 ( n13380 , n10227 , n35420 );
    and g10320 ( n27822 , n22573 , n34685 );
    and g10321 ( n29630 , n24849 , n8687 );
    or g10322 ( n13458 , n13312 , n28544 );
    xnor g10323 ( n12048 , n17961 , n1950 );
    and g10324 ( n2090 , n26260 , n24386 );
    or g10325 ( n7770 , n22771 , n7758 );
    and g10326 ( n8955 , n26039 , n3059 );
    or g10327 ( n15389 , n29713 , n10285 );
    xnor g10328 ( n19516 , n6812 , n33328 );
    or g10329 ( n15555 , n5017 , n23462 );
    or g10330 ( n789 , n31500 , n23090 );
    xnor g10331 ( n27193 , n27341 , n1549 );
    and g10332 ( n13074 , n25285 , n30730 );
    nor g10333 ( n34873 , n16421 , n6081 );
    nor g10334 ( n12902 , n1950 , n27066 );
    xnor g10335 ( n3753 , n2936 , n22824 );
    and g10336 ( n3631 , n23927 , n34580 );
    or g10337 ( n17400 , n5166 , n21862 );
    and g10338 ( n3046 , n7812 , n8432 );
    not g10339 ( n26759 , n16631 );
    xnor g10340 ( n21148 , n4558 , n6956 );
    and g10341 ( n5556 , n21011 , n19094 );
    nor g10342 ( n28304 , n25602 , n33197 );
    not g10343 ( n27432 , n1220 );
    and g10344 ( n16854 , n30860 , n24773 );
    xnor g10345 ( n26638 , n10469 , n13817 );
    nor g10346 ( n5509 , n34260 , n16698 );
    or g10347 ( n2763 , n1950 , n3387 );
    xnor g10348 ( n1963 , n26989 , n29884 );
    xnor g10349 ( n3445 , n36009 , n29835 );
    or g10350 ( n484 , n28221 , n15439 );
    or g10351 ( n29710 , n12930 , n29643 );
    xnor g10352 ( n7316 , n9758 , n24371 );
    and g10353 ( n22394 , n4832 , n8639 );
    or g10354 ( n3124 , n26871 , n8153 );
    and g10355 ( n29899 , n15608 , n5255 );
    or g10356 ( n10084 , n12768 , n8636 );
    and g10357 ( n20866 , n5698 , n33472 );
    xnor g10358 ( n3471 , n27005 , n7061 );
    and g10359 ( n9105 , n30436 , n27409 );
    or g10360 ( n26917 , n1950 , n7907 );
    or g10361 ( n1199 , n5158 , n23090 );
    and g10362 ( n4026 , n2569 , n5767 );
    xnor g10363 ( n21669 , n9409 , n14056 );
    xnor g10364 ( n23309 , n27552 , n5335 );
    nor g10365 ( n21177 , n28965 , n28728 );
    or g10366 ( n1449 , n18417 , n23264 );
    not g10367 ( n4382 , n6830 );
    nor g10368 ( n2641 , n15206 , n9555 );
    xnor g10369 ( n13175 , n30848 , n1202 );
    xnor g10370 ( n8553 , n24453 , n10489 );
    and g10371 ( n29976 , n18967 , n3042 );
    or g10372 ( n32196 , n5460 , n9832 );
    and g10373 ( n18521 , n17239 , n4424 );
    not g10374 ( n3725 , n22291 );
    xnor g10375 ( n23815 , n26396 , n20500 );
    or g10376 ( n35954 , n11731 , n28737 );
    or g10377 ( n24250 , n22283 , n4172 );
    and g10378 ( n8514 , n23274 , n458 );
    xnor g10379 ( n23198 , n4396 , n9091 );
    or g10380 ( n8235 , n23494 , n24259 );
    or g10381 ( n2266 , n26217 , n5208 );
    xnor g10382 ( n3551 , n30736 , n16922 );
    or g10383 ( n13954 , n29713 , n35985 );
    nor g10384 ( n26545 , n11046 , n11995 );
    or g10385 ( n11417 , n19211 , n8107 );
    nor g10386 ( n11498 , n22670 , n33157 );
    or g10387 ( n447 , n7430 , n5900 );
    or g10388 ( n4087 , n9658 , n23535 );
    xnor g10389 ( n6525 , n2442 , n3264 );
    and g10390 ( n1021 , n5862 , n13709 );
    not g10391 ( n5833 , n8865 );
    or g10392 ( n23575 , n5738 , n26428 );
    xnor g10393 ( n20705 , n32785 , n4960 );
    nor g10394 ( n14326 , n25602 , n18027 );
    or g10395 ( n7737 , n29713 , n34555 );
    xnor g10396 ( n3520 , n21990 , n15403 );
    or g10397 ( n3500 , n23087 , n16606 );
    or g10398 ( n12335 , n19546 , n30292 );
    or g10399 ( n28726 , n14970 , n27728 );
    or g10400 ( n31349 , n35276 , n32691 );
    or g10401 ( n13762 , n29884 , n1785 );
    or g10402 ( n4820 , n7594 , n10557 );
    xnor g10403 ( n10255 , n14964 , n14278 );
    or g10404 ( n19161 , n31559 , n26916 );
    nor g10405 ( n18963 , n19730 , n31825 );
    and g10406 ( n32257 , n30361 , n10307 );
    and g10407 ( n30127 , n22622 , n8887 );
    xnor g10408 ( n20357 , n32009 , n6747 );
    not g10409 ( n13235 , n29327 );
    and g10410 ( n26335 , n34995 , n24224 );
    xnor g10411 ( n9578 , n30149 , n22291 );
    not g10412 ( n23697 , n27009 );
    xnor g10413 ( n9946 , n24349 , n18495 );
    and g10414 ( n17695 , n3999 , n16122 );
    xnor g10415 ( n33517 , n583 , n5180 );
    and g10416 ( n3997 , n20847 , n16857 );
    or g10417 ( n21335 , n32857 , n28693 );
    xnor g10418 ( n31082 , n10873 , n11190 );
    xnor g10419 ( n3660 , n15997 , n14069 );
    or g10420 ( n13639 , n32673 , n23559 );
    or g10421 ( n24321 , n29487 , n6459 );
    or g10422 ( n5906 , n26508 , n27501 );
    and g10423 ( n33713 , n30906 , n23161 );
    not g10424 ( n7015 , n22517 );
    or g10425 ( n27373 , n34411 , n19946 );
    or g10426 ( n19350 , n4758 , n19001 );
    or g10427 ( n31192 , n31178 , n35402 );
    and g10428 ( n17447 , n5322 , n21431 );
    and g10429 ( n34159 , n26163 , n15701 );
    or g10430 ( n5458 , n28429 , n9194 );
    xnor g10431 ( n22068 , n28727 , n7859 );
    or g10432 ( n18362 , n6309 , n35143 );
    not g10433 ( n2903 , n10336 );
    xnor g10434 ( n30322 , n35249 , n8432 );
    or g10435 ( n28057 , n27587 , n15538 );
    xnor g10436 ( n1234 , n3955 , n17657 );
    nor g10437 ( n10397 , n20363 , n13076 );
    and g10438 ( n23792 , n9877 , n35596 );
    and g10439 ( n217 , n29447 , n17132 );
    and g10440 ( n31853 , n31774 , n4758 );
    or g10441 ( n10262 , n9793 , n9937 );
    xnor g10442 ( n14510 , n19991 , n27325 );
    xnor g10443 ( n7956 , n7197 , n1950 );
    and g10444 ( n6629 , n35178 , n10026 );
    and g10445 ( n35177 , n23378 , n12741 );
    or g10446 ( n14568 , n10300 , n31773 );
    xnor g10447 ( n25957 , n10184 , n18003 );
    xnor g10448 ( n6772 , n7159 , n14512 );
    xnor g10449 ( n9237 , n26287 , n22291 );
    and g10450 ( n29945 , n11976 , n14863 );
    xnor g10451 ( n10958 , n7505 , n23246 );
    xnor g10452 ( n31193 , n14495 , n12663 );
    or g10453 ( n24678 , n1355 , n29848 );
    or g10454 ( n20217 , n27746 , n25036 );
    or g10455 ( n4195 , n7560 , n28533 );
    xnor g10456 ( n8792 , n24725 , n4460 );
    xnor g10457 ( n13849 , n735 , n13081 );
    or g10458 ( n18091 , n4734 , n10402 );
    and g10459 ( n7442 , n32947 , n29680 );
    or g10460 ( n20788 , n7797 , n16264 );
    or g10461 ( n4393 , n24339 , n25831 );
    xnor g10462 ( n6076 , n4869 , n31354 );
    or g10463 ( n3270 , n7540 , n30660 );
    or g10464 ( n15241 , n6180 , n12774 );
    not g10465 ( n12578 , n16326 );
    or g10466 ( n14206 , n32095 , n26849 );
    or g10467 ( n8509 , n4878 , n6979 );
    xnor g10468 ( n8278 , n27571 , n30253 );
    or g10469 ( n22792 , n31289 , n19462 );
    and g10470 ( n15846 , n8548 , n5982 );
    xnor g10471 ( n7035 , n4824 , n29100 );
    or g10472 ( n3988 , n3347 , n35402 );
    and g10473 ( n18043 , n5878 , n28008 );
    or g10474 ( n3796 , n32715 , n11684 );
    xnor g10475 ( n4833 , n33880 , n31056 );
    and g10476 ( n3383 , n21559 , n12170 );
    and g10477 ( n3653 , n5427 , n6458 );
    xnor g10478 ( n7049 , n10916 , n15685 );
    xnor g10479 ( n31603 , n17379 , n16135 );
    or g10480 ( n21278 , n15037 , n20797 );
    xnor g10481 ( n23687 , n32840 , n35604 );
    and g10482 ( n6046 , n2503 , n31799 );
    or g10483 ( n18010 , n21874 , n8630 );
    xnor g10484 ( n20016 , n28641 , n18857 );
    or g10485 ( n19749 , n28585 , n10736 );
    or g10486 ( n6578 , n27291 , n19914 );
    or g10487 ( n2796 , n4960 , n34965 );
    or g10488 ( n16132 , n18456 , n924 );
    nor g10489 ( n10935 , n25533 , n11050 );
    or g10490 ( n28435 , n34907 , n15814 );
    and g10491 ( n13791 , n23457 , n10448 );
    or g10492 ( n19454 , n22619 , n18752 );
    or g10493 ( n18836 , n33346 , n16710 );
    or g10494 ( n21779 , n36087 , n25773 );
    nor g10495 ( n33299 , n35057 , n6548 );
    xnor g10496 ( n34900 , n27616 , n5615 );
    or g10497 ( n21244 , n1537 , n12128 );
    or g10498 ( n26417 , n22069 , n2543 );
    not g10499 ( n24289 , n25648 );
    not g10500 ( n24685 , n7527 );
    nor g10501 ( n24319 , n30167 , n35358 );
    xnor g10502 ( n11611 , n17647 , n17543 );
    or g10503 ( n28370 , n14557 , n12791 );
    or g10504 ( n21908 , n1801 , n23209 );
    or g10505 ( n22367 , n18790 , n27166 );
    not g10506 ( n30047 , n35481 );
    not g10507 ( n8295 , n12428 );
    xnor g10508 ( n26351 , n23250 , n24254 );
    xnor g10509 ( n738 , n23218 , n27226 );
    and g10510 ( n16344 , n28281 , n7194 );
    or g10511 ( n1409 , n30795 , n10717 );
    xnor g10512 ( n7158 , n26584 , n33530 );
    xnor g10513 ( n15360 , n21410 , n4960 );
    or g10514 ( n13435 , n35613 , n32634 );
    and g10515 ( n18877 , n34460 , n26138 );
    or g10516 ( n29898 , n28365 , n12996 );
    or g10517 ( n21385 , n29839 , n3210 );
    or g10518 ( n3724 , n28007 , n25419 );
    or g10519 ( n3495 , n23604 , n1723 );
    and g10520 ( n9504 , n13914 , n4146 );
    and g10521 ( n35603 , n14086 , n32219 );
    not g10522 ( n4989 , n25018 );
    and g10523 ( n5010 , n3605 , n13759 );
    or g10524 ( n7207 , n35154 , n7664 );
    not g10525 ( n13656 , n24879 );
    and g10526 ( n14006 , n31296 , n6876 );
    or g10527 ( n125 , n31272 , n4603 );
    nor g10528 ( n35824 , n18032 , n4952 );
    or g10529 ( n16948 , n15299 , n16777 );
    xnor g10530 ( n17545 , n9566 , n2485 );
    and g10531 ( n2457 , n5485 , n20822 );
    not g10532 ( n6540 , n20393 );
    and g10533 ( n13076 , n30269 , n15939 );
    or g10534 ( n2130 , n2188 , n23790 );
    and g10535 ( n5703 , n25585 , n3946 );
    not g10536 ( n13821 , n3444 );
    and g10537 ( n30076 , n10135 , n15998 );
    not g10538 ( n36064 , n7284 );
    not g10539 ( n34038 , n11101 );
    or g10540 ( n23280 , n19702 , n26549 );
    or g10541 ( n24886 , n32841 , n31554 );
    or g10542 ( n3168 , n25674 , n4042 );
    or g10543 ( n20594 , n10228 , n12951 );
    and g10544 ( n29952 , n18085 , n11439 );
    or g10545 ( n16402 , n3758 , n26052 );
    xnor g10546 ( n6814 , n18006 , n6502 );
    or g10547 ( n11136 , n33540 , n32507 );
    xnor g10548 ( n4410 , n8985 , n28989 );
    and g10549 ( n18471 , n2839 , n15790 );
    xnor g10550 ( n32508 , n16812 , n1950 );
    xnor g10551 ( n10155 , n27401 , n32095 );
    or g10552 ( n30210 , n2568 , n12843 );
    or g10553 ( n25655 , n13537 , n34865 );
    or g10554 ( n16188 , n8818 , n5208 );
    or g10555 ( n13829 , n32857 , n14363 );
    xnor g10556 ( n16527 , n14291 , n25602 );
    not g10557 ( n30877 , n25031 );
    and g10558 ( n26806 , n6657 , n6235 );
    and g10559 ( n15814 , n29025 , n7531 );
    xnor g10560 ( n26567 , n33255 , n3144 );
    xnor g10561 ( n33770 , n15079 , n34369 );
    or g10562 ( n27519 , n8001 , n29953 );
    and g10563 ( n28292 , n2130 , n11305 );
    or g10564 ( n1765 , n22626 , n17337 );
    xnor g10565 ( n17831 , n31672 , n31945 );
    and g10566 ( n6033 , n1907 , n34003 );
    or g10567 ( n2310 , n9200 , n1701 );
    or g10568 ( n26155 , n9793 , n24867 );
    or g10569 ( n1205 , n27291 , n5613 );
    or g10570 ( n13535 , n18000 , n18521 );
    or g10571 ( n27481 , n12223 , n22624 );
    or g10572 ( n25906 , n28137 , n24740 );
    and g10573 ( n19025 , n13685 , n18100 );
    xnor g10574 ( n25207 , n10813 , n16141 );
    xnor g10575 ( n23542 , n19550 , n9789 );
    or g10576 ( n939 , n4366 , n3694 );
    or g10577 ( n3157 , n32871 , n35492 );
    or g10578 ( n9348 , n27552 , n29366 );
    not g10579 ( n31044 , n26817 );
    xnor g10580 ( n35180 , n31012 , n23604 );
    or g10581 ( n29275 , n12129 , n8153 );
    or g10582 ( n21283 , n16565 , n30870 );
    or g10583 ( n22852 , n11404 , n25761 );
    or g10584 ( n18387 , n24697 , n15144 );
    xnor g10585 ( n3063 , n8890 , n3946 );
    or g10586 ( n18473 , n10075 , n15290 );
    or g10587 ( n11022 , n30987 , n28969 );
    or g10588 ( n17365 , n5085 , n15700 );
    and g10589 ( n13850 , n29970 , n30231 );
    nor g10590 ( n19763 , n32857 , n20474 );
    not g10591 ( n14956 , n32071 );
    or g10592 ( n8136 , n4897 , n30519 );
    or g10593 ( n7060 , n3731 , n4059 );
    or g10594 ( n4477 , n26460 , n8972 );
    or g10595 ( n31151 , n27291 , n3715 );
    or g10596 ( n5621 , n20646 , n12055 );
    and g10597 ( n11488 , n6244 , n30924 );
    and g10598 ( n34212 , n2725 , n12583 );
    or g10599 ( n30579 , n30468 , n19173 );
    nor g10600 ( n14313 , n22790 , n14171 );
    nor g10601 ( n19023 , n3205 , n19235 );
    xnor g10602 ( n15620 , n19209 , n16620 );
    or g10603 ( n4655 , n1187 , n3988 );
    buf g10604 ( n35141 , n22783 );
    not g10605 ( n24115 , n34865 );
    and g10606 ( n4784 , n29534 , n16784 );
    xnor g10607 ( n28599 , n15808 , n16795 );
    xnor g10608 ( n16693 , n9281 , n14184 );
    or g10609 ( n5140 , n20934 , n3694 );
    or g10610 ( n15965 , n11455 , n11872 );
    or g10611 ( n26345 , n15886 , n12466 );
    or g10612 ( n13584 , n17806 , n11833 );
    nor g10613 ( n27825 , n8432 , n26253 );
    or g10614 ( n13539 , n4288 , n9360 );
    or g10615 ( n23094 , n25130 , n16763 );
    and g10616 ( n7457 , n35838 , n16657 );
    and g10617 ( n25444 , n13670 , n31125 );
    and g10618 ( n5835 , n11698 , n24711 );
    and g10619 ( n16486 , n26920 , n33769 );
    or g10620 ( n21298 , n26436 , n29760 );
    xnor g10621 ( n15448 , n9205 , n31273 );
    and g10622 ( n16736 , n24178 , n15950 );
    not g10623 ( n9350 , n17568 );
    or g10624 ( n28583 , n12708 , n14076 );
    xnor g10625 ( n3048 , n20092 , n4507 );
    not g10626 ( n9960 , n16620 );
    and g10627 ( n22723 , n9548 , n29738 );
    or g10628 ( n20018 , n18009 , n3512 );
    or g10629 ( n18236 , n6314 , n4318 );
    or g10630 ( n6621 , n27871 , n3224 );
    or g10631 ( n16748 , n3552 , n6815 );
    and g10632 ( n7361 , n26170 , n30243 );
    and g10633 ( n18993 , n6752 , n11629 );
    or g10634 ( n28538 , n30334 , n23626 );
    or g10635 ( n31042 , n26396 , n20500 );
    buf g10636 ( n27501 , n6548 );
    or g10637 ( n6949 , n17441 , n12996 );
    or g10638 ( n15271 , n14329 , n30813 );
    xnor g10639 ( n12189 , n32614 , n24371 );
    not g10640 ( n5469 , n31215 );
    or g10641 ( n13806 , n34681 , n32049 );
    or g10642 ( n24309 , n5227 , n8924 );
    or g10643 ( n571 , n25581 , n6340 );
    not g10644 ( n26962 , n26365 );
    or g10645 ( n13833 , n21219 , n2705 );
    xnor g10646 ( n11416 , n19948 , n13677 );
    or g10647 ( n6860 , n20501 , n34756 );
    or g10648 ( n25413 , n23604 , n35724 );
    or g10649 ( n10451 , n31131 , n20318 );
    or g10650 ( n15306 , n16620 , n32325 );
    and g10651 ( n23499 , n24083 , n7889 );
    or g10652 ( n30793 , n33708 , n34862 );
    or g10653 ( n30071 , n24629 , n13795 );
    or g10654 ( n22484 , n23604 , n12813 );
    or g10655 ( n6032 , n9597 , n9938 );
    and g10656 ( n7929 , n233 , n20480 );
    and g10657 ( n27122 , n21449 , n23984 );
    nor g10658 ( n4706 , n3670 , n7453 );
    or g10659 ( n26430 , n19065 , n15826 );
    not g10660 ( n7698 , n16922 );
    xnor g10661 ( n16367 , n9891 , n7598 );
    nor g10662 ( n13591 , n1540 , n26881 );
    xnor g10663 ( n28701 , n10724 , n5425 );
    or g10664 ( n28378 , n20885 , n35402 );
    nor g10665 ( n20842 , n18353 , n29366 );
    and g10666 ( n6947 , n29965 , n17507 );
    or g10667 ( n31728 , n28368 , n4739 );
    or g10668 ( n6946 , n27653 , n29562 );
    or g10669 ( n34818 , n13364 , n13215 );
    xnor g10670 ( n32403 , n28430 , n30248 );
    and g10671 ( n5937 , n12002 , n17579 );
    nor g10672 ( n14236 , n1950 , n27473 );
    or g10673 ( n6303 , n14269 , n1511 );
    and g10674 ( n31229 , n10803 , n11725 );
    xnor g10675 ( n16491 , n10471 , n8710 );
    or g10676 ( n2579 , n24611 , n26251 );
    or g10677 ( n29766 , n9926 , n24710 );
    or g10678 ( n29938 , n26258 , n25447 );
    or g10679 ( n28207 , n22340 , n25392 );
    or g10680 ( n7660 , n9154 , n9951 );
    or g10681 ( n3781 , n4962 , n1900 );
    or g10682 ( n22584 , n6557 , n8924 );
    xnor g10683 ( n2956 , n20920 , n27226 );
    not g10684 ( n23696 , n15029 );
    and g10685 ( n10603 , n31274 , n11411 );
    or g10686 ( n28468 , n16446 , n11601 );
    not g10687 ( n5806 , n4960 );
    or g10688 ( n10254 , n32011 , n27973 );
    and g10689 ( n25471 , n16229 , n35635 );
    nor g10690 ( n16970 , n9204 , n4496 );
    xnor g10691 ( n33891 , n19122 , n10775 );
    and g10692 ( n18668 , n15130 , n28552 );
    not g10693 ( n2626 , n10521 );
    or g10694 ( n27029 , n14555 , n16797 );
    or g10695 ( n23301 , n29358 , n17872 );
    and g10696 ( n14849 , n26797 , n9475 );
    nor g10697 ( n29053 , n3946 , n22859 );
    or g10698 ( n8141 , n28654 , n27704 );
    xnor g10699 ( n3244 , n31829 , n17182 );
    and g10700 ( n3769 , n15514 , n31837 );
    xnor g10701 ( n5157 , n15619 , n4784 );
    not g10702 ( n20548 , n18478 );
    xnor g10703 ( n17791 , n27345 , n18860 );
    not g10704 ( n27497 , n937 );
    xnor g10705 ( n6917 , n30217 , n31215 );
    or g10706 ( n1460 , n24237 , n32031 );
    or g10707 ( n23724 , n9703 , n15290 );
    and g10708 ( n22318 , n34418 , n16309 );
    or g10709 ( n23125 , n830 , n5112 );
    and g10710 ( n33362 , n19648 , n32051 );
    xnor g10711 ( n894 , n27050 , n8087 );
    and g10712 ( n12894 , n28158 , n24881 );
    or g10713 ( n32201 , n34349 , n15256 );
    not g10714 ( n10823 , n1580 );
    not g10715 ( n31337 , n22501 );
    xnor g10716 ( n14396 , n16154 , n23604 );
    nor g10717 ( n7521 , n29713 , n4642 );
    and g10718 ( n26589 , n10129 , n14191 );
    and g10719 ( n17525 , n28595 , n2897 );
    and g10720 ( n20748 , n16648 , n9354 );
    and g10721 ( n7105 , n6921 , n29951 );
    or g10722 ( n32247 , n9049 , n29411 );
    and g10723 ( n16230 , n17486 , n19846 );
    or g10724 ( n9148 , n10162 , n26019 );
    and g10725 ( n28533 , n3789 , n13146 );
    or g10726 ( n27708 , n657 , n17337 );
    or g10727 ( n1194 , n11452 , n11850 );
    xnor g10728 ( n4611 , n23255 , n14298 );
    and g10729 ( n13880 , n18882 , n17571 );
    or g10730 ( n29877 , n2143 , n21210 );
    or g10731 ( n21564 , n25320 , n25067 );
    or g10732 ( n24568 , n18668 , n33435 );
    and g10733 ( n21129 , n30927 , n29774 );
    or g10734 ( n21511 , n17980 , n29562 );
    xnor g10735 ( n2035 , n20395 , n4288 );
    nor g10736 ( n12120 , n16620 , n21243 );
    not g10737 ( n19957 , n22200 );
    xnor g10738 ( n12962 , n18144 , n30421 );
    and g10739 ( n16812 , n15797 , n17461 );
    and g10740 ( n13343 , n5519 , n26526 );
    xnor g10741 ( n16495 , n34742 , n32857 );
    xnor g10742 ( n13870 , n12866 , n30725 );
    and g10743 ( n6474 , n23994 , n19437 );
    xnor g10744 ( n30311 , n5451 , n4960 );
    or g10745 ( n8256 , n12349 , n28332 );
    not g10746 ( n19748 , n32563 );
    and g10747 ( n15870 , n4870 , n155 );
    xnor g10748 ( n19237 , n13331 , n30567 );
    nor g10749 ( n8164 , n13159 , n31683 );
    and g10750 ( n30737 , n19321 , n17837 );
    nor g10751 ( n16847 , n29484 , n18026 );
    xnor g10752 ( n12152 , n13863 , n11455 );
    and g10753 ( n7845 , n7627 , n5261 );
    or g10754 ( n19453 , n27291 , n324 );
    and g10755 ( n17928 , n4514 , n1574 );
    xnor g10756 ( n4387 , n2027 , n35792 );
    or g10757 ( n35331 , n31799 , n17802 );
    or g10758 ( n35795 , n8438 , n30204 );
    or g10759 ( n8172 , n3222 , n21606 );
    not g10760 ( n3649 , n3292 );
    or g10761 ( n15494 , n5530 , n24259 );
    xnor g10762 ( n7950 , n21941 , n26337 );
    nor g10763 ( n17871 , n16620 , n9851 );
    or g10764 ( n17367 , n18769 , n3858 );
    xnor g10765 ( n13734 , n28014 , n17568 );
    or g10766 ( n21123 , n4962 , n15727 );
    xnor g10767 ( n4344 , n2022 , n36030 );
    or g10768 ( n25553 , n30466 , n11229 );
    and g10769 ( n24551 , n34303 , n30307 );
    or g10770 ( n15307 , n14629 , n19939 );
    and g10771 ( n31180 , n33823 , n15019 );
    and g10772 ( n28962 , n33278 , n17597 );
    nor g10773 ( n21791 , n3222 , n9952 );
    and g10774 ( n19892 , n21298 , n9634 );
    or g10775 ( n7469 , n11765 , n10808 );
    xnor g10776 ( n34044 , n31229 , n27226 );
    or g10777 ( n27000 , n5076 , n19421 );
    not g10778 ( n26736 , n9793 );
    xnor g10779 ( n20196 , n6730 , n18638 );
    or g10780 ( n21994 , n35176 , n32505 );
    or g10781 ( n2732 , n12062 , n10074 );
    or g10782 ( n33722 , n5429 , n19940 );
    or g10783 ( n24988 , n12284 , n23790 );
    and g10784 ( n8948 , n31664 , n35942 );
    and g10785 ( n22690 , n33509 , n1681 );
    and g10786 ( n8446 , n18624 , n3337 );
    or g10787 ( n8482 , n14676 , n11518 );
    buf g10788 ( n29411 , n266 );
    or g10789 ( n31488 , n20636 , n28586 );
    or g10790 ( n4885 , n30219 , n1582 );
    and g10791 ( n30988 , n18926 , n7752 );
    xnor g10792 ( n26757 , n27532 , n25863 );
    not g10793 ( n8312 , n2092 );
    not g10794 ( n20640 , n19310 );
    or g10795 ( n29328 , n20652 , n7169 );
    or g10796 ( n7603 , n18758 , n35329 );
    or g10797 ( n33795 , n10403 , n35400 );
    xnor g10798 ( n7765 , n33060 , n31056 );
    xnor g10799 ( n11893 , n13253 , n2874 );
    not g10800 ( n1880 , n5738 );
    not g10801 ( n33592 , n2590 );
    nor g10802 ( n18499 , n4962 , n32220 );
    and g10803 ( n8977 , n16586 , n35859 );
    or g10804 ( n16081 , n17966 , n30520 );
    nor g10805 ( n25568 , n23277 , n3165 );
    xnor g10806 ( n17104 , n11254 , n22291 );
    and g10807 ( n1846 , n16816 , n1237 );
    not g10808 ( n32722 , n7759 );
    or g10809 ( n28972 , n22257 , n33001 );
    or g10810 ( n15287 , n32939 , n11295 );
    or g10811 ( n33564 , n35494 , n3858 );
    or g10812 ( n26163 , n2439 , n12428 );
    or g10813 ( n6816 , n35827 , n21862 );
    or g10814 ( n26790 , n1045 , n18851 );
    xnor g10815 ( n19390 , n3291 , n13477 );
    or g10816 ( n29374 , n33728 , n24356 );
    nor g10817 ( n11133 , n13586 , n10327 );
    and g10818 ( n32557 , n7512 , n20729 );
    and g10819 ( n15185 , n12909 , n32974 );
    or g10820 ( n32159 , n35246 , n10663 );
    xnor g10821 ( n2346 , n1741 , n29884 );
    or g10822 ( n15058 , n22402 , n23209 );
    or g10823 ( n4581 , n34786 , n19515 );
    or g10824 ( n28433 , n30710 , n34001 );
    or g10825 ( n32173 , n30473 , n5355 );
    xor g10826 ( n94 , n1825 , n10044 );
    or g10827 ( n19902 , n9789 , n35708 );
    or g10828 ( n33423 , n17027 , n14918 );
    or g10829 ( n276 , n17577 , n25786 );
    or g10830 ( n17185 , n34837 , n10061 );
    or g10831 ( n8383 , n24422 , n24710 );
    and g10832 ( n6399 , n32637 , n7478 );
    and g10833 ( n28717 , n6887 , n3831 );
    or g10834 ( n17857 , n13326 , n6683 );
    buf g10835 ( n19464 , n13523 );
    xnor g10836 ( n2421 , n5396 , n16922 );
    or g10837 ( n10648 , n35255 , n3188 );
    or g10838 ( n7827 , n31641 , n29153 );
    xnor g10839 ( n462 , n22797 , n34380 );
    xnor g10840 ( n20936 , n23662 , n26555 );
    xnor g10841 ( n30693 , n13244 , n23071 );
    and g10842 ( n6397 , n15091 , n15662 );
    xnor g10843 ( n3197 , n19574 , n25602 );
    or g10844 ( n17511 , n29955 , n9450 );
    and g10845 ( n18706 , n9149 , n4319 );
    and g10846 ( n29125 , n13982 , n2002 );
    or g10847 ( n31660 , n16620 , n21733 );
    or g10848 ( n4137 , n27831 , n31606 );
    and g10849 ( n21700 , n35077 , n9319 );
    nor g10850 ( n35330 , n27489 , n26774 );
    not g10851 ( n12705 , n32857 );
    or g10852 ( n14368 , n4524 , n35757 );
    buf g10853 ( n9921 , n19834 );
    not g10854 ( n7477 , n651 );
    or g10855 ( n34715 , n498 , n13217 );
    or g10856 ( n14663 , n23118 , n27447 );
    and g10857 ( n14786 , n13060 , n10295 );
    or g10858 ( n7533 , n10728 , n31627 );
    or g10859 ( n2450 , n10005 , n12128 );
    or g10860 ( n26307 , n15665 , n34600 );
    or g10861 ( n7311 , n8461 , n7960 );
    and g10862 ( n34556 , n21327 , n2452 );
    or g10863 ( n10188 , n14418 , n17337 );
    and g10864 ( n32288 , n23338 , n23384 );
    xnor g10865 ( n9786 , n31862 , n6756 );
    and g10866 ( n9079 , n19831 , n14526 );
    not g10867 ( n10954 , n14831 );
    and g10868 ( n19940 , n26965 , n16761 );
    or g10869 ( n22593 , n25357 , n9832 );
    buf g10870 ( n25447 , n28783 );
    not g10871 ( n21705 , n34558 );
    or g10872 ( n10271 , n1381 , n15784 );
    or g10873 ( n4101 , n2389 , n21851 );
    xnor g10874 ( n30720 , n18758 , n35329 );
    or g10875 ( n34773 , n8432 , n25858 );
    or g10876 ( n33571 , n19443 , n4529 );
    or g10877 ( n15018 , n8212 , n23729 );
    nor g10878 ( n30319 , n5287 , n9734 );
    xnor g10879 ( n21099 , n10635 , n7032 );
    and g10880 ( n16209 , n32196 , n8979 );
    and g10881 ( n23658 , n30427 , n20639 );
    or g10882 ( n12449 , n18801 , n35244 );
    xnor g10883 ( n30442 , n20244 , n31799 );
    or g10884 ( n19548 , n16050 , n23323 );
    and g10885 ( n35737 , n23318 , n18688 );
    or g10886 ( n2881 , n4308 , n2814 );
    or g10887 ( n20207 , n31874 , n3640 );
    or g10888 ( n8868 , n14466 , n6075 );
    not g10889 ( n9506 , n4440 );
    xnor g10890 ( n16939 , n19695 , n34702 );
    xnor g10891 ( n11322 , n28855 , n15877 );
    xnor g10892 ( n764 , n17265 , n17568 );
    xnor g10893 ( n127 , n6009 , n20562 );
    or g10894 ( n30359 , n34960 , n30519 );
    or g10895 ( n17455 , n31017 , n10171 );
    or g10896 ( n27410 , n6973 , n15290 );
    and g10897 ( n1955 , n34483 , n21835 );
    xnor g10898 ( n32448 , n20615 , n19617 );
    xnor g10899 ( n22008 , n18064 , n16392 );
    or g10900 ( n26062 , n639 , n24259 );
    and g10901 ( n14512 , n18058 , n28948 );
    and g10902 ( n10290 , n32045 , n31521 );
    xor g10903 ( n6434 , n32699 , n15620 );
    xnor g10904 ( n18149 , n33170 , n32095 );
    not g10905 ( n29657 , n18919 );
    xnor g10906 ( n29918 , n27739 , n19551 );
    nor g10907 ( n6938 , n8745 , n31770 );
    and g10908 ( n26121 , n14859 , n6320 );
    or g10909 ( n2859 , n535 , n4952 );
    or g10910 ( n13126 , n26600 , n14202 );
    and g10911 ( n17622 , n5731 , n12176 );
    or g10912 ( n9340 , n22291 , n33056 );
    xnor g10913 ( n10864 , n22801 , n6077 );
    or g10914 ( n22582 , n17751 , n22968 );
    and g10915 ( n19829 , n14474 , n7492 );
    xnor g10916 ( n28349 , n14222 , n23005 );
    xnor g10917 ( n23252 , n9271 , n20623 );
    and g10918 ( n31621 , n17455 , n4567 );
    and g10919 ( n13528 , n33510 , n5992 );
    xnor g10920 ( n29001 , n13537 , n22291 );
    xnor g10921 ( n5165 , n12801 , n31289 );
    and g10922 ( n12938 , n15913 , n2517 );
    or g10923 ( n21013 , n4979 , n34888 );
    nor g10924 ( n28283 , n16617 , n6017 );
    xnor g10925 ( n13176 , n208 , n11190 );
    or g10926 ( n2343 , n7811 , n15004 );
    or g10927 ( n16856 , n23574 , n16961 );
    not g10928 ( n1090 , n30459 );
    buf g10929 ( n35630 , n3188 );
    or g10930 ( n12327 , n23613 , n24013 );
    not g10931 ( n21894 , n5298 );
    xnor g10932 ( n24727 , n29603 , n25602 );
    and g10933 ( n6348 , n25806 , n3844 );
    and g10934 ( n34398 , n13668 , n48 );
    not g10935 ( n7650 , n12436 );
    xnor g10936 ( n21867 , n19172 , n7636 );
    and g10937 ( n30062 , n27032 , n35839 );
    or g10938 ( n22659 , n23422 , n30656 );
    or g10939 ( n14880 , n4344 , n32507 );
    or g10940 ( n12976 , n8554 , n31464 );
    or g10941 ( n22269 , n22020 , n481 );
    or g10942 ( n9130 , n14059 , n2104 );
    and g10943 ( n28360 , n26987 , n31729 );
    or g10944 ( n7168 , n830 , n20535 );
    xnor g10945 ( n8656 , n11339 , n12891 );
    not g10946 ( n34744 , n9789 );
    or g10947 ( n5181 , n1950 , n34029 );
    or g10948 ( n22108 , n26499 , n2823 );
    xnor g10949 ( n30905 , n21322 , n17384 );
    not g10950 ( n17271 , n7191 );
    or g10951 ( n17014 , n15693 , n3634 );
    or g10952 ( n22145 , n16922 , n23558 );
    or g10953 ( n888 , n31955 , n30646 );
    or g10954 ( n27365 , n17304 , n35748 );
    xnor g10955 ( n8984 , n4257 , n5495 );
    not g10956 ( n6360 , n1046 );
    or g10957 ( n12336 , n32719 , n4772 );
    xnor g10958 ( n20527 , n4911 , n35927 );
    or g10959 ( n18308 , n17568 , n32981 );
    nor g10960 ( n9389 , n16620 , n33372 );
    and g10961 ( n1826 , n11584 , n19022 );
    or g10962 ( n21415 , n29839 , n33112 );
    and g10963 ( n16666 , n8555 , n33980 );
    and g10964 ( n35865 , n35730 , n34336 );
    or g10965 ( n33763 , n20050 , n19058 );
    or g10966 ( n22704 , n10465 , n27447 );
    or g10967 ( n32344 , n9451 , n26480 );
    or g10968 ( n22393 , n14103 , n19732 );
    and g10969 ( n27774 , n32001 , n9390 );
    not g10970 ( n26465 , n19939 );
    and g10971 ( n4529 , n8815 , n11885 );
    or g10972 ( n10633 , n10894 , n4540 );
    or g10973 ( n35953 , n8612 , n35388 );
    and g10974 ( n4718 , n25771 , n18785 );
    and g10975 ( n16512 , n4990 , n15864 );
    or g10976 ( n26816 , n18379 , n6573 );
    or g10977 ( n8222 , n9066 , n12996 );
    and g10978 ( n21029 , n10525 , n21191 );
    or g10979 ( n6175 , n5421 , n29626 );
    or g10980 ( n4848 , n35538 , n13900 );
    or g10981 ( n17738 , n27948 , n17046 );
    and g10982 ( n17576 , n20938 , n11026 );
    or g10983 ( n17502 , n7990 , n31554 );
    xnor g10984 ( n33511 , n19390 , n34479 );
    or g10985 ( n28697 , n13252 , n28329 );
    and g10986 ( n2217 , n7278 , n17735 );
    or g10987 ( n20710 , n9094 , n29988 );
    xnor g10988 ( n25256 , n35972 , n9957 );
    or g10989 ( n25085 , n2954 , n17554 );
    xnor g10990 ( n9370 , n21748 , n18219 );
    and g10991 ( n6089 , n4738 , n27581 );
    not g10992 ( n33218 , n9789 );
    xnor g10993 ( n3795 , n21425 , n4836 );
    or g10994 ( n23224 , n3995 , n19058 );
    or g10995 ( n7236 , n34798 , n21977 );
    xnor g10996 ( n5502 , n2648 , n1580 );
    nor g10997 ( n10717 , n25131 , n29707 );
    and g10998 ( n3546 , n31733 , n12108 );
    not g10999 ( n1179 , n6538 );
    xnor g11000 ( n34286 , n25073 , n25605 );
    and g11001 ( n14342 , n34809 , n22568 );
    or g11002 ( n27555 , n25602 , n1370 );
    xnor g11003 ( n2263 , n22713 , n4962 );
    or g11004 ( n33736 , n30998 , n27770 );
    or g11005 ( n30363 , n24315 , n28574 );
    and g11006 ( n26101 , n33359 , n34412 );
    not g11007 ( n31544 , n19551 );
    not g11008 ( n22931 , n6086 );
    and g11009 ( n20875 , n10018 , n26324 );
    xnor g11010 ( n25930 , n35557 , n27226 );
    and g11011 ( n770 , n23821 , n18396 );
    or g11012 ( n22857 , n7540 , n26037 );
    xnor g11013 ( n25105 , n10999 , n32715 );
    xnor g11014 ( n19152 , n35808 , n7540 );
    xnor g11015 ( n30933 , n26315 , n27085 );
    xnor g11016 ( n15720 , n26047 , n15886 );
    and g11017 ( n15170 , n21325 , n24052 );
    or g11018 ( n12967 , n8988 , n19173 );
    not g11019 ( n9153 , n20532 );
    xnor g11020 ( n229 , n16159 , n441 );
    or g11021 ( n10780 , n16620 , n11166 );
    or g11022 ( n81 , n15006 , n18542 );
    and g11023 ( n19374 , n23451 , n3449 );
    or g11024 ( n25865 , n29778 , n25673 );
    and g11025 ( n746 , n5783 , n10013 );
    or g11026 ( n17973 , n31289 , n10676 );
    not g11027 ( n14310 , n23007 );
    xnor g11028 ( n29320 , n12514 , n34440 );
    or g11029 ( n30508 , n19951 , n6459 );
    or g11030 ( n9732 , n19049 , n31049 );
    or g11031 ( n17199 , n8356 , n18248 );
    and g11032 ( n15565 , n5001 , n12589 );
    or g11033 ( n31458 , n4288 , n30025 );
    or g11034 ( n11660 , n13712 , n25763 );
    or g11035 ( n16144 , n30239 , n31514 );
    or g11036 ( n11917 , n31194 , n28675 );
    xnor g11037 ( n24403 , n32973 , n282 );
    xnor g11038 ( n26499 , n19290 , n7433 );
    nor g11039 ( n32860 , n27291 , n27295 );
    or g11040 ( n20131 , n14954 , n15774 );
    or g11041 ( n34107 , n18120 , n7481 );
    and g11042 ( n8778 , n34031 , n33580 );
    or g11043 ( n8991 , n33753 , n33956 );
    and g11044 ( n10808 , n14550 , n6098 );
    xnor g11045 ( n19513 , n3284 , n32715 );
    nor g11046 ( n12931 , n31215 , n30492 );
    or g11047 ( n9342 , n3303 , n7046 );
    xnor g11048 ( n9814 , n27465 , n29884 );
    and g11049 ( n13526 , n34112 , n32560 );
    and g11050 ( n14570 , n33817 , n21367 );
    and g11051 ( n3995 , n8736 , n12119 );
    or g11052 ( n30864 , n2819 , n1143 );
    or g11053 ( n24655 , n19772 , n29393 );
    not g11054 ( n14689 , n9361 );
    xnor g11055 ( n15535 , n12044 , n3205 );
    or g11056 ( n23515 , n13082 , n28866 );
    or g11057 ( n35015 , n31361 , n28248 );
    nor g11058 ( n26295 , n10894 , n18569 );
    and g11059 ( n15060 , n28589 , n14199 );
    and g11060 ( n7074 , n21593 , n975 );
    and g11061 ( n27769 , n3192 , n27953 );
    or g11062 ( n23246 , n27825 , n22338 );
    or g11063 ( n22556 , n31819 , n8366 );
    and g11064 ( n3824 , n33097 , n12258 );
    buf g11065 ( n3239 , n13758 );
    xnor g11066 ( n32818 , n8042 , n7065 );
    and g11067 ( n31275 , n29198 , n19902 );
    or g11068 ( n15632 , n34554 , n21691 );
    xnor g11069 ( n5483 , n23196 , n15745 );
    xnor g11070 ( n19211 , n6698 , n23604 );
    nor g11071 ( n24611 , n30141 , n8807 );
    and g11072 ( n32785 , n31950 , n19745 );
    nor g11073 ( n27114 , n13020 , n4719 );
    and g11074 ( n34434 , n9912 , n33832 );
    or g11075 ( n35049 , n1950 , n7645 );
    and g11076 ( n4954 , n13191 , n8591 );
    or g11077 ( n18259 , n18978 , n29830 );
    or g11078 ( n25125 , n25995 , n423 );
    xnor g11079 ( n28630 , n24669 , n9941 );
    or g11080 ( n18640 , n28721 , n12913 );
    and g11081 ( n13805 , n25868 , n35549 );
    or g11082 ( n15910 , n15924 , n25447 );
    xnor g11083 ( n1396 , n14960 , n33936 );
    not g11084 ( n4128 , n26007 );
    or g11085 ( n28341 , n27226 , n26966 );
    or g11086 ( n29849 , n23604 , n4972 );
    or g11087 ( n18586 , n27291 , n24104 );
    not g11088 ( n8285 , n15883 );
    and g11089 ( n6755 , n23474 , n5468 );
    and g11090 ( n32685 , n28041 , n28516 );
    or g11091 ( n24958 , n32584 , n29391 );
    and g11092 ( n34162 , n16682 , n11434 );
    and g11093 ( n18061 , n7406 , n27220 );
    not g11094 ( n31745 , n6535 );
    or g11095 ( n23927 , n15648 , n16562 );
    xnor g11096 ( n24213 , n27599 , n16620 );
    and g11097 ( n1207 , n32512 , n8620 );
    xnor g11098 ( n9724 , n2357 , n15333 );
    or g11099 ( n3179 , n19170 , n17354 );
    xnor g11100 ( n11070 , n25141 , n21540 );
    or g11101 ( n30920 , n12441 , n578 );
    or g11102 ( n21306 , n35188 , n28940 );
    buf g11103 ( n585 , n27728 );
    and g11104 ( n27868 , n13357 , n33054 );
    nor g11105 ( n14193 , n20678 , n31411 );
    or g11106 ( n19046 , n32246 , n3188 );
    or g11107 ( n15405 , n3222 , n469 );
    xnor g11108 ( n2442 , n8487 , n22017 );
    xnor g11109 ( n26522 , n28882 , n25381 );
    and g11110 ( n30393 , n15629 , n30941 );
    or g11111 ( n2775 , n11239 , n23344 );
    or g11112 ( n8736 , n23500 , n3738 );
    or g11113 ( n25487 , n24371 , n16831 );
    nor g11114 ( n33979 , n1698 , n15828 );
    or g11115 ( n24558 , n402 , n11239 );
    not g11116 ( n13449 , n17204 );
    not g11117 ( n19402 , n8366 );
    or g11118 ( n4020 , n154 , n16192 );
    and g11119 ( n1244 , n31074 , n19066 );
    or g11120 ( n34026 , n28022 , n30109 );
    or g11121 ( n16354 , n32614 , n4661 );
    nor g11122 ( n1016 , n4461 , n1511 );
    and g11123 ( n15638 , n28912 , n5256 );
    or g11124 ( n4752 , n4624 , n20762 );
    not g11125 ( n28711 , n17568 );
    or g11126 ( n11685 , n16894 , n6436 );
    and g11127 ( n10416 , n9046 , n27291 );
    or g11128 ( n12746 , n30526 , n23762 );
    or g11129 ( n5132 , n22655 , n29061 );
    or g11130 ( n31490 , n32639 , n12622 );
    buf g11131 ( n34923 , n35080 );
    or g11132 ( n4714 , n25602 , n15148 );
    or g11133 ( n17685 , n10175 , n5980 );
    and g11134 ( n18621 , n29962 , n15634 );
    or g11135 ( n8146 , n10164 , n20762 );
    xnor g11136 ( n24264 , n4638 , n16579 );
    or g11137 ( n1017 , n34119 , n4254 );
    nor g11138 ( n22040 , n4758 , n20169 );
    not g11139 ( n1386 , n20029 );
    xnor g11140 ( n29543 , n34751 , n17970 );
    nor g11141 ( n4761 , n23339 , n33956 );
    or g11142 ( n9710 , n1576 , n24333 );
    or g11143 ( n13597 , n9853 , n15743 );
    or g11144 ( n10836 , n2413 , n7673 );
    xnor g11145 ( n26166 , n28972 , n16620 );
    not g11146 ( n12092 , n16225 );
    nor g11147 ( n16755 , n7540 , n20717 );
    and g11148 ( n12798 , n13119 , n12975 );
    xnor g11149 ( n24057 , n31972 , n2749 );
    not g11150 ( n30908 , n10967 );
    and g11151 ( n16729 , n3507 , n16256 );
    xnor g11152 ( n25894 , n19406 , n25497 );
    and g11153 ( n34467 , n21203 , n8603 );
    not g11154 ( n24996 , n7619 );
    and g11155 ( n24165 , n26150 , n26793 );
    and g11156 ( n34792 , n25261 , n27034 );
    or g11157 ( n18685 , n1657 , n23015 );
    and g11158 ( n24967 , n6147 , n11423 );
    or g11159 ( n28663 , n6051 , n1511 );
    or g11160 ( n35233 , n19715 , n3961 );
    or g11161 ( n34000 , n10965 , n24356 );
    or g11162 ( n35001 , n9409 , n18407 );
    xnor g11163 ( n10228 , n2076 , n11046 );
    xnor g11164 ( n34400 , n1768 , n4878 );
    or g11165 ( n32303 , n19331 , n15778 );
    or g11166 ( n24500 , n109 , n29841 );
    xnor g11167 ( n3771 , n2493 , n16982 );
    or g11168 ( n19803 , n26210 , n20840 );
    and g11169 ( n24791 , n11374 , n19175 );
    nor g11170 ( n33498 , n8634 , n33680 );
    or g11171 ( n4521 , n33517 , n29953 );
    and g11172 ( n16609 , n6126 , n22152 );
    and g11173 ( n35820 , n11061 , n18528 );
    xnor g11174 ( n27175 , n25324 , n22198 );
    xnor g11175 ( n14553 , n18222 , n33521 );
    xnor g11176 ( n28565 , n23634 , n24837 );
    xnor g11177 ( n9902 , n19630 , n33767 );
    xnor g11178 ( n24245 , n32393 , n27291 );
    not g11179 ( n27954 , n29579 );
    or g11180 ( n26191 , n22614 , n17829 );
    and g11181 ( n7926 , n816 , n17563 );
    or g11182 ( n4339 , n19201 , n28668 );
    buf g11183 ( n2798 , n7446 );
    nor g11184 ( n2649 , n12751 , n34165 );
    or g11185 ( n24691 , n8355 , n15977 );
    or g11186 ( n12974 , n28203 , n19994 );
    xnor g11187 ( n5158 , n10508 , n16139 );
    or g11188 ( n23388 , n24371 , n35356 );
    xnor g11189 ( n31513 , n24442 , n22281 );
    xnor g11190 ( n5422 , n18935 , n27291 );
    or g11191 ( n1190 , n13502 , n34130 );
    or g11192 ( n18496 , n30742 , n29631 );
    and g11193 ( n12272 , n19539 , n19361 );
    and g11194 ( n20937 , n2146 , n19929 );
    xnor g11195 ( n15412 , n29515 , n4878 );
    xnor g11196 ( n20164 , n30192 , n20177 );
    or g11197 ( n19725 , n35750 , n19732 );
    nor g11198 ( n15778 , n23940 , n22130 );
    nor g11199 ( n24562 , n15886 , n14073 );
    or g11200 ( n27706 , n32857 , n28678 );
    or g11201 ( n15955 , n12845 , n4595 );
    and g11202 ( n9411 , n34191 , n22980 );
    or g11203 ( n5418 , n25602 , n5351 );
    or g11204 ( n35952 , n27741 , n1715 );
    or g11205 ( n8228 , n27226 , n23218 );
    or g11206 ( n8 , n21369 , n18240 );
    not g11207 ( n1404 , n30732 );
    or g11208 ( n5859 , n8564 , n4490 );
    xnor g11209 ( n378 , n35737 , n9793 );
    and g11210 ( n34224 , n9537 , n15749 );
    or g11211 ( n25063 , n8440 , n19421 );
    or g11212 ( n12528 , n4673 , n16213 );
    or g11213 ( n28671 , n35927 , n26833 );
    or g11214 ( n9996 , n35002 , n5618 );
    or g11215 ( n10427 , n17982 , n28123 );
    and g11216 ( n23312 , n34102 , n56 );
    and g11217 ( n22578 , n1241 , n10909 );
    or g11218 ( n6893 , n11551 , n3553 );
    and g11219 ( n13943 , n26241 , n2414 );
    or g11220 ( n34230 , n1616 , n13215 );
    or g11221 ( n12393 , n28501 , n16510 );
    nor g11222 ( n17743 , n29713 , n29831 );
    nor g11223 ( n12244 , n19736 , n11161 );
    or g11224 ( n24370 , n21243 , n13909 );
    xnor g11225 ( n18641 , n11575 , n31581 );
    and g11226 ( n7793 , n34672 , n24451 );
    or g11227 ( n11610 , n11862 , n20498 );
    or g11228 ( n116 , n29031 , n7293 );
    or g11229 ( n9797 , n19054 , n22749 );
    and g11230 ( n54 , n16785 , n8697 );
    or g11231 ( n8111 , n10748 , n23990 );
    not g11232 ( n16817 , n30732 );
    xnor g11233 ( n6093 , n6207 , n30451 );
    or g11234 ( n10032 , n35791 , n19464 );
    or g11235 ( n1214 , n25435 , n26365 );
    nor g11236 ( n5487 , n16620 , n19272 );
    or g11237 ( n26487 , n31289 , n14718 );
    xnor g11238 ( n34915 , n16857 , n29949 );
    xnor g11239 ( n6180 , n29232 , n32857 );
    nor g11240 ( n33382 , n20416 , n4285 );
    xnor g11241 ( n15660 , n28157 , n24528 );
    xnor g11242 ( n23727 , n28571 , n21553 );
    xnor g11243 ( n16332 , n12480 , n31559 );
    or g11244 ( n20394 , n23067 , n9317 );
    or g11245 ( n16349 , n11956 , n7254 );
    or g11246 ( n6969 , n35737 , n9731 );
    or g11247 ( n15411 , n2632 , n35757 );
    xnor g11248 ( n10821 , n9814 , n25350 );
    nor g11249 ( n8016 , n32095 , n7925 );
    or g11250 ( n5265 , n35811 , n35998 );
    or g11251 ( n12810 , n4208 , n3756 );
    not g11252 ( n10067 , n30742 );
    and g11253 ( n23324 , n6737 , n30108 );
    and g11254 ( n4273 , n13500 , n2990 );
    or g11255 ( n14334 , n17445 , n30354 );
    and g11256 ( n13046 , n16994 , n29526 );
    or g11257 ( n30868 , n11455 , n30386 );
    and g11258 ( n17321 , n26076 , n25353 );
    or g11259 ( n30247 , n5394 , n13008 );
    not g11260 ( n15383 , n2433 );
    and g11261 ( n18204 , n7160 , n24313 );
    xnor g11262 ( n6199 , n9980 , n7587 );
    and g11263 ( n1712 , n30336 , n30849 );
    not g11264 ( n26672 , n2029 );
    nor g11265 ( n12895 , n13998 , n30624 );
    not g11266 ( n15094 , n4962 );
    not g11267 ( n30299 , n28438 );
    or g11268 ( n25039 , n33380 , n1946 );
    and g11269 ( n14800 , n31313 , n11402 );
    or g11270 ( n3743 , n32095 , n28549 );
    and g11271 ( n23939 , n19563 , n22795 );
    xnor g11272 ( n12122 , n899 , n3222 );
    and g11273 ( n3461 , n14094 , n8529 );
    and g11274 ( n14295 , n13724 , n20698 );
    or g11275 ( n26880 , n32095 , n11193 );
    and g11276 ( n8201 , n21909 , n369 );
    or g11277 ( n12113 , n5009 , n19421 );
    and g11278 ( n18403 , n13882 , n24604 );
    xnor g11279 ( n26481 , n27949 , n703 );
    or g11280 ( n12551 , n30994 , n3738 );
    or g11281 ( n16171 , n21049 , n2119 );
    or g11282 ( n24487 , n31900 , n26480 );
    xnor g11283 ( n2354 , n3467 , n26514 );
    xnor g11284 ( n27429 , n1393 , n34025 );
    xnor g11285 ( n19591 , n23443 , n17116 );
    not g11286 ( n31896 , n20009 );
    xnor g11287 ( n4755 , n12630 , n9882 );
    nor g11288 ( n23138 , n11190 , n28211 );
    and g11289 ( n32331 , n32125 , n33714 );
    or g11290 ( n10480 , n3635 , n25592 );
    or g11291 ( n19696 , n14396 , n15611 );
    and g11292 ( n18778 , n7329 , n32454 );
    and g11293 ( n14516 , n11095 , n9122 );
    xnor g11294 ( n27629 , n14381 , n29370 );
    nor g11295 ( n6120 , n12942 , n12879 );
    or g11296 ( n17625 , n15669 , n17162 );
    and g11297 ( n34997 , n5856 , n11358 );
    and g11298 ( n4405 , n26572 , n10123 );
    and g11299 ( n1019 , n32364 , n22463 );
    or g11300 ( n6158 , n3205 , n24279 );
    or g11301 ( n36073 , n34434 , n11977 );
    and g11302 ( n29821 , n14596 , n14153 );
    buf g11303 ( n26220 , n29533 );
    or g11304 ( n12305 , n30276 , n33440 );
    and g11305 ( n34867 , n32610 , n21600 );
    nor g11306 ( n10182 , n23953 , n6984 );
    nor g11307 ( n9315 , n20774 , n2098 );
    or g11308 ( n17712 , n27613 , n26002 );
    or g11309 ( n6542 , n2694 , n15925 );
    or g11310 ( n28543 , n35927 , n32685 );
    and g11311 ( n25907 , n2017 , n5409 );
    or g11312 ( n1896 , n22837 , n27426 );
    and g11313 ( n15296 , n7205 , n4083 );
    or g11314 ( n31316 , n25094 , n32634 );
    or g11315 ( n15077 , n9658 , n27275 );
    and g11316 ( n5677 , n3625 , n23117 );
    xnor g11317 ( n8797 , n23621 , n24332 );
    or g11318 ( n23330 , n28358 , n14232 );
    xnor g11319 ( n1847 , n26502 , n15084 );
    and g11320 ( n11866 , n4934 , n24715 );
    xnor g11321 ( n12921 , n5740 , n13857 );
    or g11322 ( n13044 , n22291 , n3162 );
    and g11323 ( n34132 , n22156 , n4576 );
    and g11324 ( n1718 , n33203 , n13981 );
    and g11325 ( n13923 , n929 , n18436 );
    or g11326 ( n13017 , n8388 , n544 );
    and g11327 ( n27011 , n26221 , n14583 );
    and g11328 ( n27643 , n7764 , n22629 );
    xnor g11329 ( n25327 , n19346 , n16660 );
    xnor g11330 ( n15716 , n13794 , n26089 );
    or g11331 ( n14479 , n7540 , n1296 );
    xnor g11332 ( n3194 , n24210 , n19044 );
    and g11333 ( n657 , n6164 , n2255 );
    or g11334 ( n11214 , n29864 , n23489 );
    or g11335 ( n2114 , n31570 , n17068 );
    or g11336 ( n35499 , n14021 , n16457 );
    or g11337 ( n19004 , n8294 , n18542 );
    xnor g11338 ( n35925 , n146 , n1145 );
    not g11339 ( n1529 , n26229 );
    xnor g11340 ( n34374 , n22750 , n35927 );
    xnor g11341 ( n33374 , n4379 , n1950 );
    and g11342 ( n32270 , n908 , n35037 );
    or g11343 ( n11191 , n24413 , n27588 );
    not g11344 ( n24508 , n4920 );
    and g11345 ( n32284 , n33345 , n3700 );
    xnor g11346 ( n8198 , n18061 , n29839 );
    or g11347 ( n28959 , n9289 , n12086 );
    not g11348 ( n35269 , n344 );
    or g11349 ( n3608 , n24930 , n34484 );
    and g11350 ( n6582 , n4054 , n15245 );
    or g11351 ( n19082 , n11797 , n5556 );
    and g11352 ( n17304 , n32201 , n327 );
    or g11353 ( n12337 , n26356 , n15290 );
    and g11354 ( n33139 , n20617 , n27081 );
    xnor g11355 ( n6192 , n21846 , n5067 );
    or g11356 ( n31499 , n3222 , n17998 );
    and g11357 ( n5309 , n16474 , n28662 );
    not g11358 ( n15068 , n3904 );
    or g11359 ( n2272 , n12885 , n30462 );
    nor g11360 ( n34778 , n5335 , n17558 );
    or g11361 ( n31628 , n4878 , n4157 );
    and g11362 ( n28882 , n20575 , n24436 );
    or g11363 ( n18314 , n3128 , n34865 );
    or g11364 ( n2477 , n33299 , n12052 );
    nor g11365 ( n30741 , n26851 , n13312 );
    and g11366 ( n25914 , n21764 , n32743 );
    buf g11367 ( n8723 , n10083 );
    and g11368 ( n13426 , n13379 , n7400 );
    or g11369 ( n17714 , n12 , n24479 );
    or g11370 ( n11726 , n11068 , n5779 );
    not g11371 ( n10617 , n32105 );
    nor g11372 ( n1593 , n16620 , n26969 );
    xnor g11373 ( n12989 , n3653 , n17568 );
    or g11374 ( n13484 , n32095 , n32950 );
    not g11375 ( n31563 , n30732 );
    or g11376 ( n20388 , n32274 , n13016 );
    or g11377 ( n9531 , n30080 , n11756 );
    xnor g11378 ( n21647 , n4336 , n16760 );
    and g11379 ( n23459 , n9632 , n2988 );
    and g11380 ( n17756 , n23563 , n4375 );
    or g11381 ( n7904 , n33511 , n19105 );
    and g11382 ( n29078 , n20579 , n1456 );
    or g11383 ( n5276 , n33276 , n17698 );
    or g11384 ( n16605 , n20349 , n28248 );
    or g11385 ( n14002 , n2913 , n529 );
    or g11386 ( n31568 , n22308 , n28396 );
    xnor g11387 ( n30099 , n28315 , n5287 );
    xnor g11388 ( n26998 , n14944 , n6414 );
    xnor g11389 ( n16722 , n31516 , n9422 );
    and g11390 ( n3747 , n14002 , n17832 );
    and g11391 ( n13540 , n460 , n17222 );
    or g11392 ( n24090 , n32625 , n4450 );
    or g11393 ( n11651 , n24806 , n1414 );
    not g11394 ( n13255 , n5390 );
    xnor g11395 ( n30129 , n31751 , n4718 );
    xnor g11396 ( n35870 , n24791 , n29884 );
    and g11397 ( n11060 , n8069 , n20208 );
    xnor g11398 ( n22652 , n32192 , n20 );
    nor g11399 ( n24147 , n4962 , n9703 );
    or g11400 ( n35569 , n19420 , n8366 );
    or g11401 ( n25974 , n14326 , n24277 );
    or g11402 ( n28002 , n24580 , n12879 );
    or g11403 ( n23119 , n11745 , n34484 );
    and g11404 ( n14991 , n18387 , n28392 );
    or g11405 ( n29668 , n33670 , n31773 );
    and g11406 ( n1739 , n9888 , n21957 );
    and g11407 ( n29229 , n31670 , n3667 );
    and g11408 ( n32874 , n14111 , n32405 );
    or g11409 ( n30560 , n7228 , n7803 );
    or g11410 ( n74 , n18795 , n22946 );
    and g11411 ( n15164 , n9941 , n24669 );
    or g11412 ( n20607 , n1172 , n21862 );
    or g11413 ( n16416 , n10500 , n6340 );
    and g11414 ( n17775 , n14337 , n35850 );
    nor g11415 ( n25438 , n4878 , n19291 );
    or g11416 ( n13868 , n4960 , n15755 );
    or g11417 ( n29210 , n32796 , n16762 );
    nor g11418 ( n28363 , n27717 , n35540 );
    and g11419 ( n11750 , n10642 , n20299 );
    xnor g11420 ( n35964 , n25400 , n17447 );
    not g11421 ( n33791 , n3545 );
    or g11422 ( n35984 , n4414 , n10603 );
    xor g11423 ( n25277 , n26840 , n29304 );
    xnor g11424 ( n11534 , n33407 , n4288 );
    or g11425 ( n33512 , n20926 , n28453 );
    and g11426 ( n7404 , n22092 , n28840 );
    or g11427 ( n21581 , n21184 , n32634 );
    xnor g11428 ( n32536 , n32636 , n28168 );
    or g11429 ( n6461 , n13515 , n28843 );
    nor g11430 ( n15568 , n28003 , n17120 );
    or g11431 ( n12287 , n25980 , n16802 );
    xnor g11432 ( n35596 , n29136 , n9858 );
    buf g11433 ( n19939 , n32586 );
    and g11434 ( n1345 , n2816 , n33715 );
    or g11435 ( n19308 , n29839 , n17246 );
    xnor g11436 ( n19580 , n21806 , n10345 );
    xnor g11437 ( n3054 , n19534 , n4702 );
    xnor g11438 ( n20260 , n26846 , n16820 );
    and g11439 ( n14397 , n17549 , n11944 );
    or g11440 ( n26011 , n24290 , n19945 );
    and g11441 ( n23906 , n35333 , n29827 );
    or g11442 ( n1906 , n23080 , n3352 );
    or g11443 ( n35910 , n15403 , n18321 );
    nor g11444 ( n31466 , n16620 , n27599 );
    and g11445 ( n30417 , n11564 , n19815 );
    not g11446 ( n6793 , n20227 );
    and g11447 ( n25228 , n19840 , n20903 );
    xnor g11448 ( n7224 , n15057 , n148 );
    and g11449 ( n12929 , n27304 , n18148 );
    or g11450 ( n20741 , n18744 , n26002 );
    or g11451 ( n23841 , n8286 , n26112 );
    or g11452 ( n12842 , n5844 , n28544 );
    or g11453 ( n16270 , n25474 , n23399 );
    or g11454 ( n33329 , n2506 , n13305 );
    and g11455 ( n1051 , n10746 , n34797 );
    not g11456 ( n916 , n20558 );
    and g11457 ( n7734 , n33147 , n34692 );
    or g11458 ( n4111 , n1936 , n585 );
    xnor g11459 ( n26072 , n9883 , n19317 );
    and g11460 ( n30205 , n16772 , n5463 );
    not g11461 ( n33590 , n34865 );
    or g11462 ( n1237 , n7540 , n6755 );
    or g11463 ( n30673 , n10108 , n1856 );
    and g11464 ( n34965 , n24301 , n21952 );
    xor g11465 ( n35414 , n9686 , n10192 );
    or g11466 ( n18070 , n35927 , n20934 );
    and g11467 ( n33331 , n30071 , n16997 );
    not g11468 ( n7962 , n30204 );
    xnor g11469 ( n31503 , n9980 , n5648 );
    xnor g11470 ( n18468 , n21711 , n31496 );
    or g11471 ( n35718 , n12520 , n21800 );
    or g11472 ( n1722 , n9658 , n6906 );
    nor g11473 ( n14551 , n11190 , n35017 );
    or g11474 ( n33383 , n16199 , n22682 );
    xnor g11475 ( n5688 , n29009 , n8677 );
    and g11476 ( n27356 , n31123 , n10361 );
    buf g11477 ( n24333 , n3681 );
    xnor g11478 ( n3014 , n11424 , n9793 );
    and g11479 ( n6302 , n18728 , n20550 );
    or g11480 ( n2926 , n11916 , n2275 );
    xnor g11481 ( n23997 , n7484 , n3222 );
    and g11482 ( n29611 , n21312 , n5386 );
    and g11483 ( n18915 , n31325 , n35620 );
    or g11484 ( n4502 , n10167 , n8153 );
    or g11485 ( n16976 , n14734 , n14076 );
    xnor g11486 ( n20697 , n35175 , n14003 );
    not g11487 ( n28853 , n5990 );
    nor g11488 ( n3440 , n27291 , n23008 );
    and g11489 ( n26390 , n23135 , n20011 );
    or g11490 ( n32985 , n30207 , n2104 );
    xnor g11491 ( n18026 , n19881 , n16620 );
    and g11492 ( n20518 , n11207 , n18894 );
    and g11493 ( n21699 , n32483 , n20974 );
    or g11494 ( n8644 , n32316 , n13923 );
    and g11495 ( n29531 , n20298 , n28109 );
    or g11496 ( n16704 , n6206 , n24489 );
    nor g11497 ( n32263 , n23427 , n18115 );
    nor g11498 ( n1497 , n3664 , n33956 );
    xnor g11499 ( n12251 , n1524 , n32095 );
    or g11500 ( n17 , n1567 , n18542 );
    and g11501 ( n25332 , n3709 , n4714 );
    nor g11502 ( n7610 , n24445 , n31411 );
    or g11503 ( n24273 , n7691 , n31464 );
    or g11504 ( n17593 , n5628 , n11601 );
    xnor g11505 ( n28975 , n28862 , n29148 );
    or g11506 ( n35226 , n27352 , n10634 );
    xnor g11507 ( n14532 , n21507 , n19984 );
    or g11508 ( n19021 , n18470 , n26457 );
    not g11509 ( n22811 , n303 );
    or g11510 ( n13970 , n19168 , n5900 );
    and g11511 ( n3368 , n27029 , n25053 );
    or g11512 ( n6255 , n2702 , n6868 );
    or g11513 ( n22711 , n31804 , n27539 );
    xnor g11514 ( n35706 , n18120 , n7481 );
    xnor g11515 ( n30529 , n15975 , n18267 );
    not g11516 ( n20765 , n24778 );
    and g11517 ( n29276 , n28645 , n31592 );
    or g11518 ( n21676 , n14621 , n11274 );
    or g11519 ( n26640 , n9454 , n23890 );
    xnor g11520 ( n21394 , n1282 , n1950 );
    and g11521 ( n26132 , n6260 , n22748 );
    or g11522 ( n22891 , n27936 , n20201 );
    and g11523 ( n10882 , n23073 , n25639 );
    or g11524 ( n3787 , n15101 , n1957 );
    xnor g11525 ( n17134 , n11416 , n9903 );
    nor g11526 ( n13961 , n4878 , n25633 );
    or g11527 ( n21443 , n18518 , n32329 );
    xnor g11528 ( n32069 , n1115 , n30126 );
    xnor g11529 ( n23362 , n11639 , n16137 );
    or g11530 ( n27136 , n33490 , n23300 );
    or g11531 ( n31152 , n11621 , n4772 );
    and g11532 ( n24530 , n13105 , n28379 );
    or g11533 ( n16572 , n5689 , n2005 );
    xnor g11534 ( n7969 , n5565 , n24332 );
    xnor g11535 ( n27252 , n33214 , n8034 );
    and g11536 ( n28308 , n7468 , n8990 );
    and g11537 ( n11148 , n26149 , n23220 );
    or g11538 ( n33391 , n14450 , n35402 );
    or g11539 ( n15362 , n18651 , n32961 );
    nor g11540 ( n12671 , n8445 , n23499 );
    xnor g11541 ( n14388 , n33555 , n13902 );
    or g11542 ( n9233 , n29713 , n1740 );
    nor g11543 ( n13437 , n5335 , n17321 );
    or g11544 ( n2231 , n14763 , n28592 );
    nor g11545 ( n30766 , n4878 , n4682 );
    xnor g11546 ( n19477 , n31676 , n11998 );
    nor g11547 ( n26778 , n30742 , n16381 );
    xnor g11548 ( n9600 , n13375 , n31053 );
    nor g11549 ( n6524 , n5883 , n19084 );
    or g11550 ( n30356 , n4684 , n28064 );
    xnor g11551 ( n26303 , n14897 , n23879 );
    or g11552 ( n4452 , n12821 , n9706 );
    and g11553 ( n423 , n11580 , n17680 );
    or g11554 ( n35864 , n12047 , n23529 );
    and g11555 ( n26472 , n26976 , n1860 );
    xnor g11556 ( n34441 , n25218 , n23981 );
    and g11557 ( n1049 , n20850 , n21119 );
    and g11558 ( n14447 , n6006 , n4548 );
    buf g11559 ( n17872 , n33200 );
    or g11560 ( n5596 , n26237 , n30708 );
    nor g11561 ( n3351 , n12914 , n11877 );
    nor g11562 ( n21044 , n32924 , n20040 );
    xnor g11563 ( n13736 , n8816 , n4482 );
    or g11564 ( n33754 , n7466 , n17872 );
    and g11565 ( n35307 , n19365 , n964 );
    and g11566 ( n8298 , n33193 , n5661 );
    and g11567 ( n6589 , n1517 , n1994 );
    or g11568 ( n4114 , n880 , n13246 );
    not g11569 ( n7359 , n8050 );
    or g11570 ( n26708 , n19551 , n29975 );
    or g11571 ( n10972 , n23604 , n34168 );
    and g11572 ( n5260 , n8095 , n732 );
    and g11573 ( n3310 , n8694 , n1201 );
    or g11574 ( n24557 , n26638 , n10872 );
    not g11575 ( n16079 , n25602 );
    or g11576 ( n4886 , n14154 , n30177 );
    or g11577 ( n24144 , n4120 , n35935 );
    or g11578 ( n7402 , n34839 , n3239 );
    xnor g11579 ( n28142 , n19118 , n4288 );
    xnor g11580 ( n4890 , n18760 , n947 );
    not g11581 ( n11350 , n29928 );
    or g11582 ( n17112 , n27375 , n9672 );
    xnor g11583 ( n16655 , n27979 , n439 );
    not g11584 ( n8269 , n3480 );
    or g11585 ( n9486 , n8528 , n489 );
    xnor g11586 ( n11645 , n17577 , n21358 );
    or g11587 ( n22128 , n35927 , n5421 );
    nor g11588 ( n10819 , n4288 , n14983 );
    nor g11589 ( n20901 , n8431 , n3015 );
    xnor g11590 ( n7811 , n31069 , n15886 );
    not g11591 ( n15737 , n35783 );
    or g11592 ( n23962 , n34424 , n13062 );
    or g11593 ( n6974 , n35867 , n33581 );
    or g11594 ( n36061 , n9721 , n32959 );
    or g11595 ( n2627 , n4962 , n24613 );
    nor g11596 ( n31269 , n32857 , n24455 );
    and g11597 ( n27619 , n29894 , n15489 );
    nor g11598 ( n32068 , n27291 , n32393 );
    and g11599 ( n12073 , n31810 , n22493 );
    and g11600 ( n4725 , n13908 , n25078 );
    or g11601 ( n31353 , n10922 , n29562 );
    or g11602 ( n1973 , n2469 , n29562 );
    and g11603 ( n1018 , n13559 , n9932 );
    xnor g11604 ( n680 , n31311 , n1950 );
    or g11605 ( n6625 , n19802 , n8473 );
    or g11606 ( n1471 , n25902 , n1763 );
    or g11607 ( n6174 , n14744 , n25355 );
    xnor g11608 ( n23156 , n1076 , n16125 );
    or g11609 ( n29567 , n987 , n6459 );
    and g11610 ( n3759 , n15911 , n25374 );
    or g11611 ( n15873 , n11784 , n18307 );
    xnor g11612 ( n25995 , n20212 , n13553 );
    or g11613 ( n14859 , n28945 , n27758 );
    or g11614 ( n14559 , n35888 , n22097 );
    or g11615 ( n17341 , n10974 , n19970 );
    and g11616 ( n3178 , n17797 , n13164 );
    or g11617 ( n9252 , n27671 , n27790 );
    xnor g11618 ( n32056 , n33928 , n15422 );
    and g11619 ( n12218 , n16754 , n7607 );
    and g11620 ( n52 , n20471 , n5586 );
    and g11621 ( n30045 , n16458 , n15147 );
    or g11622 ( n32556 , n32361 , n2524 );
    nor g11623 ( n873 , n20983 , n22200 );
    or g11624 ( n25114 , n25932 , n27801 );
    or g11625 ( n13687 , n5419 , n34251 );
    and g11626 ( n18007 , n34410 , n11875 );
    nor g11627 ( n16161 , n32715 , n16038 );
    or g11628 ( n18957 , n8432 , n27587 );
    or g11629 ( n33625 , n26673 , n23332 );
    or g11630 ( n35539 , n21671 , n29256 );
    nor g11631 ( n9287 , n32588 , n8761 );
    or g11632 ( n23204 , n6013 , n33655 );
    or g11633 ( n19332 , n1556 , n3756 );
    nor g11634 ( n23475 , n4878 , n10008 );
    or g11635 ( n31096 , n5625 , n16594 );
    and g11636 ( n14183 , n6187 , n4944 );
    and g11637 ( n11810 , n30539 , n34308 );
    or g11638 ( n12965 , n7767 , n17872 );
    xnor g11639 ( n31421 , n25118 , n30218 );
    xnor g11640 ( n23132 , n30838 , n29713 );
    or g11641 ( n27101 , n2592 , n3090 );
    nor g11642 ( n11758 , n10894 , n18318 );
    or g11643 ( n13258 , n997 , n32071 );
    nor g11644 ( n18932 , n13517 , n34945 );
    or g11645 ( n13950 , n1280 , n3561 );
    xnor g11646 ( n11608 , n2719 , n3807 );
    not g11647 ( n7584 , n26268 );
    not g11648 ( n17893 , n14890 );
    or g11649 ( n10431 , n28779 , n31704 );
    xnor g11650 ( n14202 , n27179 , n9960 );
    and g11651 ( n27724 , n10203 , n30666 );
    not g11652 ( n691 , n25803 );
    nor g11653 ( n3848 , n19347 , n35935 );
    or g11654 ( n31078 , n9123 , n9979 );
    nor g11655 ( n31301 , n34051 , n4508 );
    xnor g11656 ( n21924 , n18525 , n5067 );
    or g11657 ( n14499 , n25731 , n24716 );
    xnor g11658 ( n18832 , n17938 , n13747 );
    nor g11659 ( n16039 , n24728 , n11113 );
    xnor g11660 ( n7142 , n29081 , n1950 );
    or g11661 ( n306 , n11318 , n12221 );
    or g11662 ( n32553 , n10918 , n8392 );
    or g11663 ( n13958 , n28111 , n6565 );
    and g11664 ( n8985 , n18186 , n22640 );
    or g11665 ( n17693 , n4288 , n33407 );
    or g11666 ( n4764 , n4540 , n23748 );
    or g11667 ( n14868 , n19203 , n19939 );
    or g11668 ( n20345 , n6513 , n6401 );
    buf g11669 ( n15496 , n7650 );
    and g11670 ( n3026 , n33427 , n18215 );
    and g11671 ( n25793 , n5971 , n10552 );
    or g11672 ( n9158 , n20610 , n16345 );
    or g11673 ( n24667 , n23231 , n31991 );
    and g11674 ( n1026 , n34523 , n1387 );
    xnor g11675 ( n24956 , n14817 , n32857 );
    or g11676 ( n31452 , n18050 , n5752 );
    not g11677 ( n25194 , n32857 );
    or g11678 ( n15710 , n10 , n21977 );
    xnor g11679 ( n13278 , n23461 , n33950 );
    and g11680 ( n31128 , n28310 , n17959 );
    or g11681 ( n9424 , n18431 , n17964 );
    or g11682 ( n34067 , n19276 , n26962 );
    or g11683 ( n595 , n9789 , n4901 );
    or g11684 ( n23578 , n1495 , n10872 );
    or g11685 ( n1059 , n23604 , n27288 );
    nor g11686 ( n22029 , n9658 , n28174 );
    xnor g11687 ( n29410 , n31792 , n7540 );
    or g11688 ( n25505 , n1643 , n33416 );
    or g11689 ( n25886 , n20447 , n19848 );
    or g11690 ( n35602 , n14945 , n301 );
    or g11691 ( n3082 , n2711 , n1200 );
    or g11692 ( n4432 , n20199 , n15099 );
    and g11693 ( n19450 , n23397 , n15711 );
    or g11694 ( n6232 , n4878 , n6468 );
    nor g11695 ( n17968 , n10678 , n23377 );
    or g11696 ( n1571 , n11455 , n15055 );
    or g11697 ( n22779 , n1784 , n13307 );
    or g11698 ( n279 , n30742 , n498 );
    not g11699 ( n8282 , n30459 );
    and g11700 ( n7240 , n9595 , n15027 );
    or g11701 ( n31277 , n32728 , n807 );
    and g11702 ( n5884 , n3886 , n31520 );
    xnor g11703 ( n16095 , n21666 , n29866 );
    or g11704 ( n1947 , n3769 , n29393 );
    not g11705 ( n12781 , n35927 );
    or g11706 ( n27371 , n5936 , n2384 );
    or g11707 ( n33181 , n24737 , n10082 );
    nor g11708 ( n5174 , n35927 , n2931 );
    nor g11709 ( n35109 , n10233 , n5699 );
    buf g11710 ( n18488 , n32209 );
    nor g11711 ( n19742 , n19551 , n19975 );
    nor g11712 ( n27689 , n3749 , n9767 );
    or g11713 ( n2884 , n25602 , n19934 );
    buf g11714 ( n9601 , n34048 );
    or g11715 ( n5647 , n6710 , n30448 );
    or g11716 ( n9400 , n15285 , n32505 );
    or g11717 ( n3300 , n32584 , n14485 );
    or g11718 ( n6455 , n8432 , n27164 );
    and g11719 ( n23574 , n24815 , n35041 );
    or g11720 ( n26302 , n29163 , n16896 );
    and g11721 ( n24602 , n3173 , n22504 );
    or g11722 ( n34217 , n22817 , n18974 );
    or g11723 ( n27951 , n4962 , n12883 );
    or g11724 ( n15335 , n9355 , n28240 );
    xnor g11725 ( n35680 , n15128 , n19984 );
    or g11726 ( n34318 , n23095 , n14874 );
    not g11727 ( n31727 , n10894 );
    xnor g11728 ( n8563 , n11335 , n21181 );
    or g11729 ( n24367 , n14311 , n5993 );
    or g11730 ( n24190 , n14105 , n28248 );
    and g11731 ( n33301 , n15589 , n35836 );
    or g11732 ( n31142 , n15882 , n5161 );
    not g11733 ( n18103 , n15886 );
    xnor g11734 ( n5144 , n5690 , n11190 );
    or g11735 ( n35456 , n31272 , n16980 );
    xnor g11736 ( n9045 , n3036 , n4716 );
    not g11737 ( n9670 , n28167 );
    not g11738 ( n12473 , n2732 );
    or g11739 ( n31001 , n8206 , n14289 );
    nor g11740 ( n13283 , n31056 , n16547 );
    xnor g11741 ( n4296 , n4766 , n20001 );
    or g11742 ( n7276 , n16250 , n25773 );
    or g11743 ( n17074 , n660 , n29630 );
    xnor g11744 ( n26978 , n21124 , n32857 );
    or g11745 ( n465 , n19395 , n20812 );
    or g11746 ( n20081 , n1094 , n20540 );
    and g11747 ( n22279 , n25960 , n28474 );
    or g11748 ( n19463 , n9627 , n33892 );
    or g11749 ( n8173 , n22068 , n32572 );
    not g11750 ( n19385 , n26860 );
    or g11751 ( n3201 , n11535 , n20427 );
    and g11752 ( n3637 , n24526 , n13391 );
    or g11753 ( n19221 , n10873 , n27574 );
    xnor g11754 ( n25991 , n16666 , n4878 );
    not g11755 ( n20913 , n33256 );
    or g11756 ( n5486 , n25058 , n17227 );
    or g11757 ( n26840 , n23859 , n12174 );
    xnor g11758 ( n20299 , n10287 , n14024 );
    not g11759 ( n33621 , n5226 );
    or g11760 ( n10343 , n30692 , n15145 );
    xnor g11761 ( n29579 , n20411 , n26337 );
    xnor g11762 ( n17586 , n410 , n10894 );
    nor g11763 ( n18535 , n22291 , n23292 );
    or g11764 ( n30571 , n25454 , n31811 );
    and g11765 ( n31794 , n480 , n6287 );
    and g11766 ( n20277 , n30458 , n4087 );
    or g11767 ( n15557 , n30599 , n29953 );
    or g11768 ( n26482 , n31799 , n29464 );
    xnor g11769 ( n31986 , n57 , n1832 );
    xnor g11770 ( n13355 , n25189 , n30553 );
    or g11771 ( n33128 , n17454 , n4175 );
    nor g11772 ( n10772 , n17043 , n5087 );
    or g11773 ( n6552 , n29208 , n33435 );
    or g11774 ( n35926 , n8432 , n31453 );
    and g11775 ( n32707 , n30220 , n5381 );
    xnor g11776 ( n24519 , n31420 , n26865 );
    and g11777 ( n27794 , n16020 , n33587 );
    xnor g11778 ( n31394 , n7987 , n19984 );
    nor g11779 ( n17385 , n15479 , n24672 );
    or g11780 ( n8314 , n15886 , n11157 );
    xnor g11781 ( n20331 , n19216 , n24371 );
    or g11782 ( n20267 , n25637 , n26017 );
    or g11783 ( n32609 , n1726 , n19979 );
    not g11784 ( n14158 , n6534 );
    xnor g11785 ( n11087 , n19395 , n11967 );
    or g11786 ( n31585 , n31190 , n5868 );
    xnor g11787 ( n7801 , n12883 , n31744 );
    xnor g11788 ( n32745 , n26098 , n33118 );
    or g11789 ( n31764 , n1496 , n35815 );
    and g11790 ( n2157 , n28729 , n35926 );
    xnor g11791 ( n13561 , n24082 , n27402 );
    xnor g11792 ( n5356 , n2113 , n21453 );
    or g11793 ( n13778 , n22268 , n28240 );
    or g11794 ( n19442 , n32068 , n26437 );
    xnor g11795 ( n22892 , n12867 , n7540 );
    xnor g11796 ( n30876 , n378 , n3815 );
    or g11797 ( n12694 , n25090 , n10762 );
    not g11798 ( n28094 , n11600 );
    or g11799 ( n23391 , n2864 , n14196 );
    xnor g11800 ( n34926 , n17557 , n970 );
    not g11801 ( n23452 , n7535 );
    and g11802 ( n35858 , n29285 , n18980 );
    not g11803 ( n3673 , n35379 );
    or g11804 ( n160 , n4878 , n4179 );
    xnor g11805 ( n4538 , n3889 , n29125 );
    not g11806 ( n10422 , n3258 );
    xnor g11807 ( n23142 , n22489 , n3340 );
    or g11808 ( n27856 , n19422 , n15834 );
    xnor g11809 ( n18815 , n19235 , n5837 );
    xnor g11810 ( n23718 , n2258 , n3199 );
    nor g11811 ( n16328 , n5631 , n7571 );
    or g11812 ( n25557 , n14233 , n32959 );
    xnor g11813 ( n29946 , n29583 , n34404 );
    and g11814 ( n29361 , n12884 , n25490 );
    or g11815 ( n24597 , n17315 , n17111 );
    xnor g11816 ( n35497 , n29108 , n34937 );
    and g11817 ( n14284 , n1915 , n33845 );
    xnor g11818 ( n35534 , n27804 , n19551 );
    or g11819 ( n27197 , n18694 , n13305 );
    or g11820 ( n32910 , n30821 , n25594 );
    or g11821 ( n4459 , n11164 , n19084 );
    not g11822 ( n31257 , n25398 );
    and g11823 ( n13949 , n21422 , n17654 );
    or g11824 ( n1043 , n30742 , n2271 );
    or g11825 ( n21495 , n10609 , n31163 );
    and g11826 ( n35854 , n25479 , n17826 );
    or g11827 ( n11707 , n19172 , n7636 );
    xnor g11828 ( n33868 , n23507 , n25602 );
    or g11829 ( n4198 , n30742 , n23924 );
    and g11830 ( n19019 , n11631 , n20195 );
    or g11831 ( n13554 , n33492 , n13307 );
    or g11832 ( n24451 , n28978 , n18488 );
    or g11833 ( n33907 , n35175 , n14003 );
    and g11834 ( n3897 , n26828 , n15922 );
    and g11835 ( n24088 , n10551 , n7625 );
    or g11836 ( n31642 , n5335 , n12172 );
    or g11837 ( n11515 , n5335 , n15040 );
    or g11838 ( n21182 , n16620 , n35368 );
    or g11839 ( n250 , n20956 , n7553 );
    xnor g11840 ( n20092 , n18201 , n17568 );
    and g11841 ( n29633 , n5364 , n27312 );
    and g11842 ( n8776 , n35829 , n33385 );
    xnor g11843 ( n4863 , n21297 , n5335 );
    xnor g11844 ( n18959 , n14855 , n35832 );
    and g11845 ( n13478 , n32490 , n29429 );
    and g11846 ( n7230 , n16962 , n19116 );
    or g11847 ( n16627 , n910 , n19403 );
    or g11848 ( n18451 , n25775 , n18255 );
    xnor g11849 ( n3322 , n31743 , n29434 );
    or g11850 ( n21503 , n24371 , n3821 );
    xnor g11851 ( n25033 , n12122 , n10656 );
    xnor g11852 ( n13634 , n8038 , n23257 );
    and g11853 ( n18819 , n207 , n26808 );
    and g11854 ( n6780 , n31645 , n35566 );
    and g11855 ( n29363 , n8873 , n5069 );
    xnor g11856 ( n5687 , n11538 , n8432 );
    or g11857 ( n15176 , n13572 , n20830 );
    not g11858 ( n21550 , n5786 );
    not g11859 ( n29645 , n16930 );
    xnor g11860 ( n1139 , n12696 , n1764 );
    nor g11861 ( n2412 , n31289 , n2521 );
    or g11862 ( n8746 , n32337 , n3546 );
    or g11863 ( n5629 , n30907 , n29562 );
    xnor g11864 ( n11202 , n31051 , n11589 );
    and g11865 ( n5313 , n30338 , n23530 );
    xnor g11866 ( n11742 , n16967 , n30915 );
    nor g11867 ( n34626 , n18831 , n8724 );
    nor g11868 ( n24926 , n22891 , n28987 );
    not g11869 ( n134 , n35168 );
    xnor g11870 ( n27461 , n34482 , n19551 );
    xnor g11871 ( n35183 , n32774 , n7081 );
    xnor g11872 ( n28869 , n8534 , n31550 );
    nor g11873 ( n33162 , n4960 , n4948 );
    and g11874 ( n19878 , n15885 , n21672 );
    nor g11875 ( n26476 , n24774 , n29932 );
    not g11876 ( n33275 , n32608 );
    and g11877 ( n24583 , n1162 , n22980 );
    or g11878 ( n9314 , n29253 , n13305 );
    and g11879 ( n8154 , n25936 , n29498 );
    not g11880 ( n3619 , n30575 );
    xnor g11881 ( n24607 , n20403 , n4288 );
    nor g11882 ( n287 , n35144 , n26369 );
    or g11883 ( n33234 , n9793 , n26581 );
    xnor g11884 ( n19996 , n19127 , n35971 );
    xnor g11885 ( n9589 , n7432 , n12857 );
    nor g11886 ( n472 , n16620 , n13392 );
    and g11887 ( n33977 , n29047 , n21677 );
    xnor g11888 ( n2782 , n23478 , n11013 );
    and g11889 ( n12833 , n26774 , n172 );
    not g11890 ( n7122 , n23604 );
    or g11891 ( n1851 , n5695 , n5252 );
    and g11892 ( n3419 , n6163 , n35884 );
    and g11893 ( n31768 , n981 , n5046 );
    or g11894 ( n23135 , n20530 , n17111 );
    xnor g11895 ( n33129 , n30236 , n30284 );
    or g11896 ( n8558 , n34802 , n5208 );
    or g11897 ( n25253 , n26325 , n28438 );
    or g11898 ( n7936 , n12558 , n12540 );
    or g11899 ( n35755 , n11019 , n4627 );
    xnor g11900 ( n2269 , n22341 , n8735 );
    or g11901 ( n18540 , n25602 , n20032 );
    or g11902 ( n14304 , n24161 , n24653 );
    xnor g11903 ( n20232 , n22157 , n16767 );
    and g11904 ( n13717 , n35851 , n20122 );
    xnor g11905 ( n34595 , n25814 , n8432 );
    and g11906 ( n22871 , n27384 , n22980 );
    or g11907 ( n35278 , n31289 , n1565 );
    xnor g11908 ( n29357 , n1767 , n26626 );
    or g11909 ( n33303 , n14589 , n27053 );
    and g11910 ( n27573 , n934 , n8715 );
    or g11911 ( n10023 , n23653 , n28668 );
    not g11912 ( n16586 , n30335 );
    or g11913 ( n27340 , n31582 , n22946 );
    nor g11914 ( n25296 , n9472 , n4875 );
    xnor g11915 ( n7826 , n296 , n32857 );
    xnor g11916 ( n3521 , n27377 , n3915 );
    not g11917 ( n4102 , n12084 );
    or g11918 ( n35654 , n25602 , n7589 );
    not g11919 ( n31599 , n22001 );
    and g11920 ( n228 , n17911 , n33481 );
    or g11921 ( n15750 , n16501 , n10273 );
    or g11922 ( n8442 , n5617 , n30853 );
    or g11923 ( n32665 , n20991 , n3733 );
    nor g11924 ( n13951 , n11455 , n10767 );
    nor g11925 ( n35568 , n16620 , n22511 );
    or g11926 ( n26338 , n7978 , n1511 );
    xnor g11927 ( n26871 , n12914 , n11877 );
    or g11928 ( n7607 , n10691 , n30870 );
    not g11929 ( n22881 , n9808 );
    or g11930 ( n32819 , n8432 , n34829 );
    or g11931 ( n8010 , n6870 , n6278 );
    or g11932 ( n15769 , n30182 , n13887 );
    or g11933 ( n30691 , n23564 , n4443 );
    and g11934 ( n980 , n18720 , n30110 );
    and g11935 ( n13234 , n16231 , n34686 );
    xnor g11936 ( n33789 , n4918 , n19708 );
    or g11937 ( n24831 , n339 , n12791 );
    or g11938 ( n24313 , n10885 , n22858 );
    buf g11939 ( n24672 , n30519 );
    and g11940 ( n26184 , n4309 , n10618 );
    or g11941 ( n23788 , n395 , n30561 );
    xnor g11942 ( n34758 , n19789 , n31799 );
    or g11943 ( n3417 , n24141 , n35315 );
    or g11944 ( n30203 , n8895 , n10960 );
    xnor g11945 ( n16034 , n483 , n10889 );
    or g11946 ( n4571 , n4089 , n34493 );
    or g11947 ( n5558 , n7766 , n33098 );
    or g11948 ( n9491 , n5640 , n16797 );
    or g11949 ( n9560 , n4960 , n15846 );
    xnor g11950 ( n4208 , n8230 , n27792 );
    and g11951 ( n25597 , n8904 , n27442 );
    not g11952 ( n25167 , n31977 );
    or g11953 ( n12754 , n20184 , n19952 );
    xnor g11954 ( n11817 , n28851 , n18829 );
    xnor g11955 ( n11604 , n5076 , n16922 );
    or g11956 ( n11828 , n29218 , n35757 );
    or g11957 ( n21070 , n17038 , n24486 );
    or g11958 ( n6635 , n23428 , n7673 );
    not g11959 ( n29545 , n23784 );
    or g11960 ( n15391 , n16404 , n29872 );
    or g11961 ( n20411 , n44 , n20711 );
    nor g11962 ( n13053 , n2254 , n8018 );
    or g11963 ( n5007 , n23604 , n34737 );
    or g11964 ( n25706 , n12726 , n30732 );
    or g11965 ( n32839 , n24258 , n6339 );
    or g11966 ( n35686 , n32538 , n12996 );
    not g11967 ( n29315 , n29830 );
    xnor g11968 ( n30511 , n17707 , n28184 );
    or g11969 ( n13206 , n11242 , n12465 );
    and g11970 ( n991 , n24348 , n19522 );
    or g11971 ( n16300 , n27161 , n17111 );
    or g11972 ( n33241 , n5354 , n19732 );
    xnor g11973 ( n14107 , n32478 , n33158 );
    xnor g11974 ( n25141 , n20025 , n5335 );
    or g11975 ( n19282 , n12382 , n20300 );
    not g11976 ( n7162 , n8262 );
    nor g11977 ( n2488 , n5679 , n2211 );
    or g11978 ( n13009 , n5684 , n8723 );
    and g11979 ( n3633 , n23739 , n6934 );
    xnor g11980 ( n9218 , n21603 , n24371 );
    xnor g11981 ( n35349 , n21089 , n4960 );
    or g11982 ( n25509 , n6022 , n33174 );
    or g11983 ( n2398 , n1950 , n1057 );
    xnor g11984 ( n11404 , n353 , n11690 );
    xnor g11985 ( n4814 , n29079 , n8262 );
    or g11986 ( n22987 , n13690 , n21210 );
    and g11987 ( n9879 , n15543 , n5895 );
    not g11988 ( n33380 , n21337 );
    or g11989 ( n20165 , n30742 , n35854 );
    or g11990 ( n11449 , n15545 , n28438 );
    or g11991 ( n35003 , n18379 , n16944 );
    xnor g11992 ( n11559 , n22174 , n33447 );
    or g11993 ( n33484 , n34052 , n21386 );
    or g11994 ( n11130 , n29713 , n7272 );
    xnor g11995 ( n9384 , n7756 , n1245 );
    or g11996 ( n15327 , n24371 , n1228 );
    or g11997 ( n17874 , n12095 , n11896 );
    or g11998 ( n8788 , n22099 , n32071 );
    or g11999 ( n9167 , n35167 , n21081 );
    xnor g12000 ( n31051 , n8778 , n32095 );
    and g12001 ( n20806 , n15455 , n23006 );
    xnor g12002 ( n13266 , n5987 , n9668 );
    and g12003 ( n7200 , n30570 , n33563 );
    xnor g12004 ( n15300 , n1135 , n6720 );
    nor g12005 ( n8671 , n223 , n2774 );
    or g12006 ( n15129 , n22291 , n24840 );
    or g12007 ( n16758 , n23924 , n3736 );
    or g12008 ( n28682 , n35927 , n18584 );
    xnor g12009 ( n26222 , n19577 , n5707 );
    or g12010 ( n10205 , n3092 , n33854 );
    not g12011 ( n25533 , n22980 );
    and g12012 ( n31150 , n25782 , n31597 );
    xnor g12013 ( n453 , n3833 , n10752 );
    xnor g12014 ( n13253 , n16365 , n9858 );
    or g12015 ( n34539 , n11020 , n8749 );
    or g12016 ( n2373 , n25602 , n10647 );
    or g12017 ( n17496 , n4878 , n17441 );
    and g12018 ( n23633 , n14833 , n8309 );
    or g12019 ( n22121 , n4962 , n8703 );
    or g12020 ( n11210 , n8304 , n17046 );
    xnor g12021 ( n6022 , n31467 , n9793 );
    and g12022 ( n20426 , n9874 , n21493 );
    xnor g12023 ( n28126 , n27723 , n6099 );
    nor g12024 ( n7538 , n23027 , n34764 );
    or g12025 ( n31026 , n6291 , n27704 );
    or g12026 ( n34454 , n10747 , n30287 );
    and g12027 ( n9790 , n27686 , n24125 );
    xnor g12028 ( n2654 , n15903 , n18565 );
    or g12029 ( n5484 , n26238 , n31554 );
    nor g12030 ( n34543 , n33629 , n22758 );
    xnor g12031 ( n13007 , n17104 , n8109 );
    or g12032 ( n23861 , n3532 , n35111 );
    or g12033 ( n1953 , n35071 , n31549 );
    xnor g12034 ( n12110 , n8488 , n29771 );
    and g12035 ( n12758 , n8448 , n15049 );
    or g12036 ( n3606 , n4811 , n19258 );
    and g12037 ( n21497 , n28944 , n26855 );
    or g12038 ( n7721 , n26687 , n908 );
    and g12039 ( n12851 , n15994 , n26353 );
    or g12040 ( n8691 , n27009 , n10159 );
    xnor g12041 ( n29027 , n14912 , n29510 );
    xnor g12042 ( n11280 , n7195 , n10894 );
    xnor g12043 ( n22247 , n11919 , n29102 );
    or g12044 ( n26153 , n34174 , n35749 );
    or g12045 ( n11549 , n342 , n8237 );
    or g12046 ( n7128 , n482 , n12128 );
    not g12047 ( n10449 , n4758 );
    or g12048 ( n29155 , n19460 , n842 );
    not g12049 ( n34408 , n19551 );
    or g12050 ( n9755 , n15886 , n15477 );
    xnor g12051 ( n30792 , n14653 , n15781 );
    nor g12052 ( n775 , n3946 , n330 );
    or g12053 ( n114 , n10192 , n23279 );
    or g12054 ( n6612 , n31879 , n16797 );
    or g12055 ( n2584 , n3662 , n11126 );
    or g12056 ( n33217 , n28214 , n28407 );
    not g12057 ( n9297 , n6257 );
    not g12058 ( n22546 , n26745 );
    xnor g12059 ( n30154 , n12401 , n11360 );
    not g12060 ( n20905 , n28273 );
    or g12061 ( n6611 , n9789 , n34665 );
    xnor g12062 ( n21366 , n9837 , n25508 );
    not g12063 ( n30167 , n27699 );
    and g12064 ( n7288 , n8315 , n9313 );
    not g12065 ( n22294 , n8432 );
    not g12066 ( n16110 , n5335 );
    or g12067 ( n671 , n26479 , n34889 );
    xnor g12068 ( n26903 , n27636 , n713 );
    or g12069 ( n6135 , n35009 , n5389 );
    or g12070 ( n24683 , n32020 , n14745 );
    or g12071 ( n9399 , n17041 , n17125 );
    or g12072 ( n4403 , n26295 , n5747 );
    and g12073 ( n6976 , n6874 , n32698 );
    or g12074 ( n16433 , n11455 , n4842 );
    and g12075 ( n28720 , n25190 , n23624 );
    or g12076 ( n12613 , n19757 , n5208 );
    xnor g12077 ( n28932 , n34 , n3946 );
    or g12078 ( n33450 , n23674 , n34284 );
    and g12079 ( n23698 , n16640 , n29320 );
    buf g12080 ( n32608 , n34076 );
    xnor g12081 ( n35788 , n30994 , n21351 );
    or g12082 ( n29714 , n4960 , n22723 );
    xor g12083 ( n35682 , n2547 , n16620 );
    not g12084 ( n17177 , n34448 );
    xnor g12085 ( n6462 , n26819 , n8349 );
    not g12086 ( n21189 , n4962 );
    or g12087 ( n30038 , n25324 , n22198 );
    nor g12088 ( n15854 , n3450 , n19244 );
    nor g12089 ( n766 , n20567 , n21657 );
    and g12090 ( n23333 , n1509 , n2482 );
    not g12091 ( n34378 , n265 );
    or g12092 ( n27598 , n3946 , n17178 );
    and g12093 ( n28288 , n24645 , n30717 );
    or g12094 ( n27055 , n4558 , n6956 );
    xnor g12095 ( n7701 , n8860 , n11412 );
    and g12096 ( n21091 , n11245 , n29713 );
    or g12097 ( n33811 , n23111 , n6692 );
    or g12098 ( n19117 , n4878 , n7876 );
    or g12099 ( n25680 , n9190 , n3736 );
    or g12100 ( n11573 , n19499 , n30708 );
    xnor g12101 ( n10466 , n6119 , n31596 );
    or g12102 ( n17697 , n17186 , n22158 );
    xnor g12103 ( n22054 , n49 , n18713 );
    or g12104 ( n21578 , n16275 , n18407 );
    xnor g12105 ( n23127 , n20383 , n26153 );
    or g12106 ( n6795 , n27879 , n29643 );
    and g12107 ( n29988 , n2830 , n30225 );
    nor g12108 ( n5852 , n19551 , n28318 );
    or g12109 ( n15059 , n32095 , n1244 );
    or g12110 ( n3601 , n30645 , n30419 );
    or g12111 ( n3047 , n11455 , n10145 );
    xor g12112 ( n14769 , n24455 , n32857 );
    xnor g12113 ( n8012 , n19948 , n11760 );
    or g12114 ( n19103 , n19251 , n4437 );
    and g12115 ( n5324 , n34449 , n16067 );
    or g12116 ( n2441 , n10894 , n31239 );
    or g12117 ( n26113 , n30922 , n3842 );
    or g12118 ( n15089 , n15609 , n28240 );
    or g12119 ( n30738 , n30224 , n10616 );
    not g12120 ( n18481 , n2597 );
    xnor g12121 ( n11888 , n23703 , n15024 );
    or g12122 ( n31179 , n33550 , n13965 );
    nor g12123 ( n7525 , n27448 , n22940 );
    not g12124 ( n31329 , n16725 );
    xnor g12125 ( n29353 , n25118 , n32694 );
    nor g12126 ( n29656 , n29456 , n33430 );
    or g12127 ( n32951 , n15886 , n28564 );
    xnor g12128 ( n6352 , n3225 , n3633 );
    or g12129 ( n1870 , n4960 , n35505 );
    xnor g12130 ( n16909 , n14616 , n19115 );
    or g12131 ( n19027 , n29185 , n1250 );
    or g12132 ( n29235 , n15317 , n17125 );
    or g12133 ( n29537 , n17868 , n25603 );
    xnor g12134 ( n15836 , n13462 , n24053 );
    not g12135 ( n18282 , n1299 );
    or g12136 ( n8847 , n17751 , n19530 );
    or g12137 ( n9508 , n5335 , n28560 );
    not g12138 ( n11000 , n22980 );
    or g12139 ( n18494 , n2765 , n35043 );
    or g12140 ( n11439 , n31981 , n28455 );
    xnor g12141 ( n87 , n34758 , n34452 );
    and g12142 ( n7488 , n8200 , n13625 );
    nor g12143 ( n29852 , n17602 , n33468 );
    nor g12144 ( n11615 , n13782 , n6069 );
    or g12145 ( n35862 , n31743 , n4058 );
    or g12146 ( n2844 , n4336 , n16760 );
    not g12147 ( n7371 , n31289 );
    xnor g12148 ( n29197 , n34187 , n29642 );
    or g12149 ( n21945 , n4677 , n4175 );
    xnor g12150 ( n8860 , n5490 , n33952 );
    or g12151 ( n19340 , n9789 , n22578 );
    xnor g12152 ( n5763 , n10328 , n2473 );
    not g12153 ( n26859 , n34856 );
    or g12154 ( n5474 , n35927 , n36033 );
    and g12155 ( n7350 , n20819 , n29812 );
    or g12156 ( n12405 , n32170 , n8366 );
    xnor g12157 ( n14301 , n35823 , n33984 );
    or g12158 ( n26982 , n15616 , n32669 );
    or g12159 ( n1742 , n20037 , n20762 );
    xnor g12160 ( n22175 , n9388 , n34806 );
    and g12161 ( n7339 , n27272 , n31241 );
    or g12162 ( n19825 , n5677 , n35609 );
    and g12163 ( n29547 , n32123 , n28470 );
    and g12164 ( n676 , n35221 , n32705 );
    buf g12165 ( n128 , n12626 );
    xnor g12166 ( n26772 , n8914 , n4962 );
    not g12167 ( n28757 , n7588 );
    or g12168 ( n9284 , n25534 , n3979 );
    xnor g12169 ( n5017 , n14482 , n5624 );
    not g12170 ( n25311 , n9077 );
    not g12171 ( n16112 , n14143 );
    or g12172 ( n11951 , n29133 , n3738 );
    or g12173 ( n8915 , n29839 , n7523 );
    and g12174 ( n25298 , n18168 , n23878 );
    xnor g12175 ( n7048 , n23550 , n10031 );
    or g12176 ( n9522 , n30054 , n10634 );
    or g12177 ( n26713 , n2729 , n5868 );
    not g12178 ( n35832 , n35927 );
    not g12179 ( n31014 , n15564 );
    or g12180 ( n32104 , n14281 , n32697 );
    or g12181 ( n2806 , n19100 , n30826 );
    xnor g12182 ( n17650 , n20198 , n14632 );
    nor g12183 ( n26255 , n3497 , n10065 );
    or g12184 ( n3117 , n14245 , n13394 );
    xnor g12185 ( n679 , n11787 , n12302 );
    and g12186 ( n12565 , n11531 , n21910 );
    xnor g12187 ( n23993 , n23602 , n10894 );
    or g12188 ( n28232 , n29741 , n12715 );
    xnor g12189 ( n4724 , n6316 , n24371 );
    xnor g12190 ( n32113 , n17441 , n4878 );
    nor g12191 ( n28076 , n5287 , n15003 );
    or g12192 ( n21127 , n6935 , n25592 );
    or g12193 ( n9830 , n32095 , n35869 );
    buf g12194 ( n6548 , n11227 );
    xnor g12195 ( n28350 , n19054 , n22749 );
    or g12196 ( n7121 , n34597 , n20817 );
    xnor g12197 ( n7030 , n13502 , n34130 );
    and g12198 ( n17050 , n29811 , n820 );
    xnor g12199 ( n31884 , n3942 , n16922 );
    and g12200 ( n35356 , n3473 , n7475 );
    buf g12201 ( n25392 , n23909 );
    and g12202 ( n4679 , n2011 , n32415 );
    not g12203 ( n32289 , n5335 );
    or g12204 ( n26071 , n20256 , n18643 );
    xnor g12205 ( n3859 , n32590 , n31559 );
    or g12206 ( n7948 , n26475 , n18264 );
    xnor g12207 ( n27771 , n33341 , n16396 );
    xnor g12208 ( n10968 , n6674 , n4470 );
    not g12209 ( n35429 , n16223 );
    and g12210 ( n35124 , n19872 , n32326 );
    and g12211 ( n16222 , n11027 , n26173 );
    or g12212 ( n31931 , n24631 , n673 );
    nor g12213 ( n23567 , n27582 , n34615 );
    nor g12214 ( n11880 , n31799 , n9768 );
    xnor g12215 ( n7452 , n29730 , n18204 );
    xnor g12216 ( n23271 , n28922 , n25397 );
    and g12217 ( n30183 , n6097 , n14509 );
    or g12218 ( n2423 , n21168 , n30419 );
    nor g12219 ( n32753 , n18114 , n21441 );
    not g12220 ( n25293 , n33128 );
    or g12221 ( n19781 , n26768 , n32447 );
    nor g12222 ( n25037 , n10070 , n12913 );
    xnor g12223 ( n604 , n9518 , n10479 );
    xnor g12224 ( n28978 , n4527 , n2981 );
    and g12225 ( n1343 , n30564 , n9114 );
    or g12226 ( n33246 , n10486 , n24112 );
    or g12227 ( n14442 , n7997 , n29050 );
    or g12228 ( n8843 , n16922 , n19170 );
    or g12229 ( n31692 , n15097 , n26594 );
    or g12230 ( n35738 , n7645 , n949 );
    or g12231 ( n24877 , n28622 , n10243 );
    and g12232 ( n12124 , n31136 , n10124 );
    and g12233 ( n28163 , n3970 , n29770 );
    xnor g12234 ( n1423 , n11907 , n29916 );
    xnor g12235 ( n35796 , n2665 , n17037 );
    or g12236 ( n1203 , n12932 , n9030 );
    and g12237 ( n24923 , n4491 , n27226 );
    xnor g12238 ( n4480 , n1978 , n5287 );
    and g12239 ( n6817 , n24901 , n14779 );
    or g12240 ( n29538 , n830 , n12991 );
    or g12241 ( n2383 , n4746 , n11844 );
    or g12242 ( n24620 , n22043 , n10952 );
    and g12243 ( n15827 , n12888 , n33531 );
    or g12244 ( n16814 , n34534 , n3806 );
    or g12245 ( n9991 , n33405 , n34537 );
    or g12246 ( n29610 , n16915 , n23072 );
    nor g12247 ( n34832 , n15299 , n318 );
    or g12248 ( n14795 , n2700 , n9930 );
    and g12249 ( n25672 , n3044 , n22964 );
    or g12250 ( n8794 , n26773 , n2814 );
    or g12251 ( n30041 , n36051 , n20817 );
    nor g12252 ( n6209 , n2314 , n4508 );
    not g12253 ( n21286 , n2045 );
    and g12254 ( n1311 , n31465 , n32776 );
    and g12255 ( n824 , n16123 , n11822 );
    and g12256 ( n8380 , n24742 , n30121 );
    xnor g12257 ( n21369 , n6314 , n31289 );
    xnor g12258 ( n28654 , n16664 , n13898 );
    or g12259 ( n30110 , n4984 , n11996 );
    xnor g12260 ( n9259 , n25811 , n22738 );
    or g12261 ( n2917 , n17751 , n2837 );
    xnor g12262 ( n6044 , n25104 , n35631 );
    or g12263 ( n4332 , n1148 , n11518 );
    buf g12264 ( n22682 , n16502 );
    and g12265 ( n17524 , n451 , n34896 );
    not g12266 ( n5952 , n603 );
    or g12267 ( n6943 , n11190 , n22292 );
    or g12268 ( n14822 , n35598 , n33310 );
    or g12269 ( n458 , n2214 , n13235 );
    xnor g12270 ( n6344 , n9980 , n20402 );
    nor g12271 ( n26280 , n16922 , n33405 );
    nor g12272 ( n22802 , n1950 , n25445 );
    or g12273 ( n13749 , n397 , n2384 );
    or g12274 ( n23454 , n7702 , n20762 );
    or g12275 ( n11920 , n11046 , n24534 );
    or g12276 ( n18211 , n9789 , n31180 );
    not g12277 ( n32502 , n15527 );
    and g12278 ( n27887 , n14942 , n3246 );
    xnor g12279 ( n25473 , n30243 , n26170 );
    or g12280 ( n22623 , n34480 , n25594 );
    not g12281 ( n33358 , n714 );
    nor g12282 ( n35348 , n9789 , n146 );
    buf g12283 ( n3858 , n27433 );
    and g12284 ( n30698 , n31018 , n30407 );
    and g12285 ( n29390 , n22141 , n34774 );
    or g12286 ( n24527 , n28988 , n16919 );
    or g12287 ( n8904 , n11216 , n14089 );
    xnor g12288 ( n31080 , n10932 , n20722 );
    or g12289 ( n24656 , n5550 , n6061 );
    or g12290 ( n24755 , n21478 , n16179 );
    or g12291 ( n26416 , n10247 , n16797 );
    nor g12292 ( n26431 , n8920 , n34615 );
    or g12293 ( n31436 , n34892 , n15135 );
    or g12294 ( n5907 , n16945 , n1693 );
    or g12295 ( n2097 , n4962 , n32811 );
    or g12296 ( n17828 , n21089 , n19421 );
    or g12297 ( n25815 , n26183 , n13900 );
    nor g12298 ( n32647 , n9658 , n255 );
    xnor g12299 ( n25313 , n20419 , n32878 );
    and g12300 ( n28710 , n24609 , n21843 );
    and g12301 ( n35078 , n34127 , n18885 );
    xnor g12302 ( n9536 , n2271 , n30742 );
    nor g12303 ( n3378 , n27074 , n25757 );
    or g12304 ( n12651 , n1551 , n1980 );
    or g12305 ( n16791 , n17764 , n27192 );
    xnor g12306 ( n21384 , n22962 , n27996 );
    xnor g12307 ( n4897 , n31206 , n20969 );
    and g12308 ( n19630 , n1782 , n20725 );
    and g12309 ( n26253 , n10020 , n9128 );
    or g12310 ( n16679 , n15768 , n13305 );
    xnor g12311 ( n24216 , n28640 , n1950 );
    or g12312 ( n34204 , n35897 , n20817 );
    xnor g12313 ( n9725 , n6156 , n19604 );
    or g12314 ( n25399 , n7224 , n23921 );
    nor g12315 ( n33539 , n30742 , n8026 );
    or g12316 ( n952 , n5960 , n24489 );
    and g12317 ( n26219 , n2245 , n10090 );
    or g12318 ( n26409 , n33188 , n34862 );
    or g12319 ( n6925 , n4878 , n3888 );
    and g12320 ( n9478 , n26940 , n5499 );
    or g12321 ( n26808 , n25602 , n20504 );
    or g12322 ( n35610 , n30537 , n23323 );
    or g12323 ( n22049 , n6136 , n14554 );
    xnor g12324 ( n11469 , n33528 , n1920 );
    and g12325 ( n35724 , n6590 , n16080 );
    nor g12326 ( n29259 , n9538 , n29203 );
    not g12327 ( n19128 , n28273 );
    or g12328 ( n33204 , n6566 , n27603 );
    and g12329 ( n21659 , n19349 , n35653 );
    nor g12330 ( n2767 , n13770 , n29045 );
    xnor g12331 ( n23511 , n26356 , n25602 );
    xnor g12332 ( n13624 , n17744 , n16922 );
    or g12333 ( n19066 , n3821 , n33034 );
    and g12334 ( n31253 , n31280 , n19384 );
    xnor g12335 ( n532 , n17500 , n31272 );
    or g12336 ( n6676 , n30498 , n26453 );
    not g12337 ( n33630 , n16922 );
    or g12338 ( n7201 , n4816 , n27392 );
    or g12339 ( n34056 , n35927 , n30960 );
    not g12340 ( n26740 , n11455 );
    not g12341 ( n12647 , n21650 );
    or g12342 ( n35293 , n2560 , n27973 );
    or g12343 ( n22428 , n28692 , n16904 );
    and g12344 ( n23032 , n16940 , n6250 );
    xnor g12345 ( n13472 , n16857 , n32225 );
    nor g12346 ( n15482 , n15886 , n10052 );
    or g12347 ( n1631 , n262 , n1474 );
    and g12348 ( n27243 , n21856 , n18540 );
    and g12349 ( n73 , n5054 , n24278 );
    or g12350 ( n10025 , n15000 , n25940 );
    or g12351 ( n2713 , n14540 , n23078 );
    xnor g12352 ( n4746 , n3448 , n22291 );
    and g12353 ( n12782 , n18473 , n21626 );
    or g12354 ( n11291 , n7227 , n26468 );
    or g12355 ( n33005 , n28769 , n14472 );
    not g12356 ( n30703 , n15886 );
    or g12357 ( n3920 , n9499 , n34537 );
    or g12358 ( n5499 , n4288 , n23737 );
    not g12359 ( n20141 , n23604 );
    or g12360 ( n17093 , n35131 , n22475 );
    or g12361 ( n23596 , n27979 , n14699 );
    xnor g12362 ( n10703 , n27620 , n7632 );
    not g12363 ( n6207 , n21102 );
    not g12364 ( n18724 , n3205 );
    not g12365 ( n4241 , n3742 );
    or g12366 ( n5126 , n26758 , n18968 );
    xnor g12367 ( n33089 , n33878 , n19090 );
    and g12368 ( n26608 , n12033 , n4959 );
    or g12369 ( n4103 , n5335 , n22693 );
    and g12370 ( n16403 , n1239 , n11158 );
    xnor g12371 ( n15270 , n33780 , n12026 );
    or g12372 ( n21527 , n5866 , n30150 );
    and g12373 ( n10246 , n33181 , n19905 );
    or g12374 ( n23054 , n9323 , n6950 );
    xnor g12375 ( n20656 , n9980 , n34604 );
    and g12376 ( n12434 , n10857 , n27942 );
    nor g12377 ( n4321 , n4288 , n16275 );
    or g12378 ( n24761 , n11592 , n35422 );
    and g12379 ( n10134 , n14178 , n7467 );
    or g12380 ( n34929 , n13823 , n33128 );
    or g12381 ( n34935 , n31534 , n20690 );
    or g12382 ( n33797 , n4169 , n11996 );
    and g12383 ( n34 , n2504 , n27708 );
    or g12384 ( n18602 , n28335 , n8872 );
    or g12385 ( n18440 , n6606 , n25255 );
    or g12386 ( n23007 , n11968 , n20982 );
    and g12387 ( n29451 , n27057 , n29476 );
    and g12388 ( n2127 , n35656 , n6273 );
    or g12389 ( n25618 , n28770 , n908 );
    or g12390 ( n13932 , n33170 , n10140 );
    and g12391 ( n30753 , n29780 , n13174 );
    or g12392 ( n22380 , n611 , n9253 );
    or g12393 ( n2934 , n13065 , n12465 );
    and g12394 ( n13619 , n19297 , n27917 );
    or g12395 ( n8427 , n12077 , n11850 );
    xnor g12396 ( n7248 , n17703 , n14141 );
    and g12397 ( n865 , n23007 , n34370 );
    or g12398 ( n29303 , n20807 , n13840 );
    or g12399 ( n3446 , n4960 , n28489 );
    or g12400 ( n2971 , n34128 , n33474 );
    and g12401 ( n17558 , n14604 , n24390 );
    xnor g12402 ( n16975 , n29808 , n30822 );
    xnor g12403 ( n18508 , n34844 , n7540 );
    or g12404 ( n22585 , n18301 , n32425 );
    or g12405 ( n1759 , n34482 , n11703 );
    xnor g12406 ( n26293 , n15678 , n31215 );
    or g12407 ( n10002 , n22190 , n21042 );
    and g12408 ( n18180 , n31732 , n6758 );
    or g12409 ( n23554 , n22534 , n20528 );
    nor g12410 ( n17407 , n4997 , n6548 );
    or g12411 ( n24396 , n1950 , n32295 );
    or g12412 ( n34887 , n21115 , n10872 );
    or g12413 ( n10795 , n35079 , n5618 );
    or g12414 ( n13182 , n6662 , n32634 );
    or g12415 ( n13814 , n22291 , n31863 );
    and g12416 ( n20540 , n24103 , n2474 );
    not g12417 ( n28641 , n10068 );
    or g12418 ( n28245 , n22906 , n34236 );
    or g12419 ( n27524 , n32095 , n33947 );
    nor g12420 ( n34860 , n4960 , n30096 );
    or g12421 ( n14610 , n31215 , n18620 );
    xnor g12422 ( n26666 , n5915 , n20911 );
    or g12423 ( n32450 , n19608 , n3188 );
    xnor g12424 ( n26234 , n5530 , n4962 );
    or g12425 ( n15833 , n17605 , n1763 );
    xnor g12426 ( n9967 , n30905 , n16589 );
    or g12427 ( n5027 , n8419 , n20427 );
    and g12428 ( n27454 , n14875 , n18539 );
    or g12429 ( n2280 , n24735 , n35402 );
    xnor g12430 ( n4778 , n3846 , n15791 );
    and g12431 ( n14628 , n33942 , n11514 );
    and g12432 ( n26211 , n476 , n276 );
    or g12433 ( n31903 , n32017 , n1307 );
    or g12434 ( n19153 , n34718 , n13880 );
    xnor g12435 ( n32360 , n23906 , n22357 );
    or g12436 ( n17514 , n6634 , n11841 );
    not g12437 ( n31625 , n19781 );
    or g12438 ( n11293 , n26398 , n1511 );
    or g12439 ( n25145 , n31289 , n31617 );
    or g12440 ( n32999 , n9658 , n5696 );
    or g12441 ( n13102 , n33635 , n34084 );
    and g12442 ( n11391 , n27523 , n2614 );
    and g12443 ( n26879 , n26618 , n21649 );
    xnor g12444 ( n31917 , n13708 , n28186 );
    and g12445 ( n16747 , n25062 , n28715 );
    or g12446 ( n8669 , n8647 , n6075 );
    or g12447 ( n17676 , n19878 , n3352 );
    buf g12448 ( n29872 , n8675 );
    or g12449 ( n24742 , n21998 , n24289 );
    and g12450 ( n1446 , n15511 , n29505 );
    nor g12451 ( n1492 , n9658 , n13462 );
    nor g12452 ( n20110 , n19551 , n18706 );
    not g12453 ( n19470 , n32601 );
    or g12454 ( n3301 , n33046 , n5850 );
    or g12455 ( n20583 , n25144 , n18033 );
    xnor g12456 ( n6141 , n17564 , n23410 );
    xnor g12457 ( n1009 , n27917 , n2753 );
    and g12458 ( n25837 , n2283 , n26432 );
    not g12459 ( n24128 , n13553 );
    or g12460 ( n35844 , n22965 , n24505 );
    or g12461 ( n21448 , n12989 , n23360 );
    or g12462 ( n12479 , n27049 , n16311 );
    xnor g12463 ( n18537 , n5382 , n32411 );
    xnor g12464 ( n13633 , n6680 , n4962 );
    or g12465 ( n30631 , n18370 , n5145 );
    and g12466 ( n15444 , n9927 , n20319 );
    xnor g12467 ( n6282 , n31722 , n17045 );
    and g12468 ( n14756 , n10251 , n27146 );
    and g12469 ( n15154 , n31093 , n29329 );
    or g12470 ( n28914 , n13553 , n34529 );
    or g12471 ( n38 , n19551 , n19444 );
    and g12472 ( n14328 , n24055 , n31767 );
    and g12473 ( n22215 , n17656 , n24644 );
    and g12474 ( n7422 , n19558 , n14891 );
    xnor g12475 ( n1289 , n4355 , n15345 );
    xnor g12476 ( n1662 , n4740 , n30742 );
    and g12477 ( n23241 , n19330 , n35890 );
    and g12478 ( n20203 , n29280 , n982 );
    not g12479 ( n9229 , n2254 );
    or g12480 ( n28957 , n15529 , n7015 );
    and g12481 ( n33327 , n16900 , n32605 );
    xnor g12482 ( n32357 , n33093 , n2799 );
    xnor g12483 ( n8401 , n3305 , n31515 );
    or g12484 ( n8941 , n2760 , n5170 );
    xnor g12485 ( n26753 , n14277 , n19286 );
    and g12486 ( n21576 , n29799 , n19948 );
    nor g12487 ( n32691 , n11000 , n22487 );
    xnor g12488 ( n1752 , n32729 , n8128 );
    and g12489 ( n6456 , n7249 , n710 );
    or g12490 ( n15122 , n21679 , n23187 );
    buf g12491 ( n23748 , n13221 );
    buf g12492 ( n12128 , n30940 );
    not g12493 ( n22017 , n29713 );
    and g12494 ( n25292 , n17124 , n22960 );
    or g12495 ( n35387 , n19328 , n10336 );
    xnor g12496 ( n7807 , n9366 , n15169 );
    and g12497 ( n18567 , n5854 , n9922 );
    or g12498 ( n4096 , n18054 , n15145 );
    or g12499 ( n14100 , n33503 , n166 );
    or g12500 ( n19423 , n16922 , n35694 );
    xnor g12501 ( n14038 , n12894 , n31056 );
    and g12502 ( n7019 , n27446 , n985 );
    or g12503 ( n4588 , n11684 , n14699 );
    xnor g12504 ( n32315 , n31209 , n33827 );
    xnor g12505 ( n8494 , n17957 , n27291 );
    and g12506 ( n20346 , n28134 , n1925 );
    and g12507 ( n27968 , n2703 , n11759 );
    xnor g12508 ( n13018 , n10064 , n31799 );
    or g12509 ( n2945 , n31808 , n30770 );
    or g12510 ( n32464 , n16939 , n18264 );
    or g12511 ( n18333 , n11403 , n24833 );
    nor g12512 ( n21891 , n17568 , n9831 );
    and g12513 ( n25760 , n21128 , n25280 );
    and g12514 ( n29049 , n4417 , n35552 );
    and g12515 ( n7914 , n9694 , n23082 );
    xnor g12516 ( n19302 , n35847 , n25174 );
    or g12517 ( n4922 , n24415 , n34484 );
    or g12518 ( n9859 , n7277 , n19241 );
    or g12519 ( n35127 , n6864 , n11833 );
    or g12520 ( n22339 , n32169 , n23396 );
    and g12521 ( n11359 , n29667 , n32741 );
    and g12522 ( n5505 , n17116 , n23443 );
    or g12523 ( n30928 , n31169 , n11850 );
    and g12524 ( n6705 , n22388 , n14902 );
    and g12525 ( n1428 , n27877 , n7988 );
    xnor g12526 ( n33143 , n34544 , n9529 );
    and g12527 ( n6649 , n23204 , n18125 );
    or g12528 ( n5885 , n34352 , n35141 );
    xnor g12529 ( n9494 , n5920 , n22989 );
    and g12530 ( n32797 , n12534 , n17847 );
    nor g12531 ( n30400 , n5716 , n11715 );
    and g12532 ( n17931 , n24420 , n4000 );
    xnor g12533 ( n23116 , n25457 , n3331 );
    xnor g12534 ( n16489 , n29006 , n3205 );
    or g12535 ( n32702 , n33296 , n9028 );
    and g12536 ( n22544 , n10238 , n32291 );
    and g12537 ( n23495 , n28095 , n22482 );
    or g12538 ( n34412 , n32255 , n10417 );
    or g12539 ( n23383 , n20475 , n13618 );
    or g12540 ( n3206 , n8881 , n1511 );
    or g12541 ( n20391 , n31977 , n24400 );
    or g12542 ( n4736 , n35690 , n31381 );
    not g12543 ( n18682 , n26720 );
    xnor g12544 ( n3875 , n35506 , n4288 );
    nor g12545 ( n6398 , n25568 , n11850 );
    and g12546 ( n28593 , n31456 , n32949 );
    or g12547 ( n35976 , n32857 , n4801 );
    not g12548 ( n5088 , n30602 );
    or g12549 ( n35648 , n18220 , n25752 );
    or g12550 ( n27670 , n24920 , n30708 );
    xnor g12551 ( n10594 , n3956 , n32095 );
    or g12552 ( n12608 , n35074 , n18264 );
    xnor g12553 ( n35229 , n12105 , n4446 );
    nor g12554 ( n12166 , n3205 , n15143 );
    or g12555 ( n5661 , n33467 , n31554 );
    and g12556 ( n8886 , n1896 , n32456 );
    not g12557 ( n6900 , n6640 );
    or g12558 ( n16541 , n9062 , n5900 );
    xnor g12559 ( n5435 , n34810 , n9658 );
    xnor g12560 ( n10930 , n19828 , n12112 );
    not g12561 ( n29703 , n14190 );
    and g12562 ( n15755 , n20482 , n17051 );
    or g12563 ( n26933 , n30742 , n8274 );
    or g12564 ( n32978 , n9793 , n7915 );
    xnor g12565 ( n24117 , n8062 , n4962 );
    not g12566 ( n19726 , n5801 );
    and g12567 ( n4044 , n22680 , n2476 );
    not g12568 ( n23066 , n4960 );
    xnor g12569 ( n14394 , n14987 , n27145 );
    or g12570 ( n14742 , n11938 , n261 );
    or g12571 ( n17049 , n6462 , n35141 );
    or g12572 ( n32700 , n28550 , n16961 );
    or g12573 ( n35409 , n9077 , n22293 );
    xnor g12574 ( n20929 , n28713 , n9658 );
    or g12575 ( n4738 , n30322 , n1207 );
    nor g12576 ( n10645 , n31799 , n11745 );
    or g12577 ( n28575 , n24792 , n29406 );
    and g12578 ( n31861 , n5370 , n20374 );
    or g12579 ( n3155 , n32682 , n34923 );
    and g12580 ( n10221 , n1635 , n22980 );
    and g12581 ( n26732 , n21059 , n21216 );
    xnor g12582 ( n29900 , n29297 , n26065 );
    and g12583 ( n27782 , n2514 , n16109 );
    or g12584 ( n25615 , n783 , n20285 );
    nor g12585 ( n25747 , n1950 , n6812 );
    xnor g12586 ( n5 , n28731 , n12469 );
    and g12587 ( n29159 , n17551 , n24832 );
    xnor g12588 ( n13197 , n15240 , n25174 );
    xnor g12589 ( n23834 , n10805 , n11045 );
    and g12590 ( n34232 , n22670 , n27327 );
    or g12591 ( n33747 , n4847 , n33915 );
    xnor g12592 ( n25058 , n8215 , n15403 );
    or g12593 ( n12279 , n5111 , n26931 );
    and g12594 ( n11800 , n6894 , n23191 );
    or g12595 ( n35366 , n1598 , n9642 );
    xnor g12596 ( n2370 , n21703 , n1950 );
    xnor g12597 ( n10369 , n17081 , n30742 );
    or g12598 ( n15113 , n10461 , n35633 );
    and g12599 ( n12171 , n21642 , n1257 );
    nor g12600 ( n1278 , n26063 , n24905 );
    or g12601 ( n17630 , n10044 , n21134 );
    and g12602 ( n23287 , n25270 , n26085 );
    and g12603 ( n24497 , n25884 , n12366 );
    nor g12604 ( n11135 , n25889 , n33069 );
    or g12605 ( n10481 , n3100 , n21002 );
    or g12606 ( n26874 , n17526 , n25255 );
    not g12607 ( n21754 , n3222 );
    and g12608 ( n2702 , n21417 , n8209 );
    and g12609 ( n28479 , n20304 , n17807 );
    and g12610 ( n34623 , n21719 , n9965 );
    or g12611 ( n8408 , n2018 , n6950 );
    not g12612 ( n3468 , n23622 );
    or g12613 ( n12805 , n21392 , n25447 );
    xnor g12614 ( n1362 , n15699 , n10662 );
    or g12615 ( n34464 , n5087 , n24207 );
    and g12616 ( n23139 , n5107 , n35726 );
    nor g12617 ( n16035 , n31625 , n20172 );
    xnor g12618 ( n7455 , n20046 , n9242 );
    or g12619 ( n19177 , n23604 , n13284 );
    or g12620 ( n33532 , n14090 , n29872 );
    or g12621 ( n30755 , n17481 , n14985 );
    or g12622 ( n9749 , n3496 , n1414 );
    and g12623 ( n27508 , n22800 , n8316 );
    or g12624 ( n15892 , n35967 , n27501 );
    or g12625 ( n15212 , n25174 , n17618 );
    xnor g12626 ( n16619 , n11873 , n32799 );
    not g12627 ( n32005 , n35677 );
    and g12628 ( n25115 , n16318 , n13607 );
    or g12629 ( n17860 , n10001 , n19421 );
    nor g12630 ( n30980 , n14380 , n1796 );
    or g12631 ( n33496 , n27339 , n17964 );
    xnor g12632 ( n11444 , n12269 , n23421 );
    or g12633 ( n25879 , n22252 , n5752 );
    xnor g12634 ( n26461 , n14444 , n31289 );
    or g12635 ( n25315 , n30278 , n15215 );
    or g12636 ( n35695 , n18144 , n32842 );
    xnor g12637 ( n31760 , n29262 , n4758 );
    or g12638 ( n5426 , n324 , n17974 );
    xnor g12639 ( n187 , n20873 , n15886 );
    xnor g12640 ( n13031 , n13572 , n20830 );
    or g12641 ( n9142 , n15724 , n34084 );
    and g12642 ( n35914 , n4767 , n19706 );
    or g12643 ( n27674 , n17123 , n6459 );
    or g12644 ( n12444 , n27817 , n8702 );
    nor g12645 ( n10549 , n15886 , n2943 );
    xor g12646 ( n12207 , n33571 , n11346 );
    not g12647 ( n20049 , n33691 );
    or g12648 ( n27485 , n5287 , n5413 );
    nor g12649 ( n24971 , n25124 , n18884 );
    or g12650 ( n24884 , n24119 , n13301 );
    xnor g12651 ( n31508 , n28463 , n15299 );
    or g12652 ( n1482 , n29578 , n24300 );
    or g12653 ( n26495 , n24371 , n27734 );
    or g12654 ( n21076 , n3946 , n20216 );
    or g12655 ( n2634 , n23604 , n17002 );
    or g12656 ( n3169 , n22157 , n16767 );
    or g12657 ( n11044 , n26408 , n3167 );
    nor g12658 ( n11905 , n32715 , n900 );
    not g12659 ( n23103 , n28305 );
    or g12660 ( n6413 , n4429 , n32507 );
    or g12661 ( n35421 , n30742 , n21497 );
    and g12662 ( n27181 , n248 , n34382 );
    and g12663 ( n9840 , n7750 , n13034 );
    or g12664 ( n13942 , n29713 , n3357 );
    xnor g12665 ( n97 , n34793 , n32259 );
    or g12666 ( n28725 , n31546 , n1176 );
    or g12667 ( n10700 , n30003 , n35868 );
    xnor g12668 ( n33 , n7472 , n26782 );
    or g12669 ( n5875 , n9789 , n34585 );
    nor g12670 ( n7313 , n26762 , n14808 );
    or g12671 ( n10245 , n29006 , n25773 );
    and g12672 ( n29258 , n22806 , n28998 );
    and g12673 ( n25104 , n2046 , n7846 );
    or g12674 ( n35155 , n25542 , n24672 );
    and g12675 ( n32780 , n15012 , n17501 );
    or g12676 ( n23353 , n9042 , n17872 );
    not g12677 ( n18113 , n16223 );
    not g12678 ( n5981 , n1181 );
    or g12679 ( n28395 , n15844 , n9920 );
    or g12680 ( n31390 , n24050 , n1796 );
    and g12681 ( n13275 , n32607 , n24578 );
    nor g12682 ( n4266 , n13553 , n27656 );
    and g12683 ( n12852 , n12465 , n24283 );
    nor g12684 ( n8225 , n17568 , n30790 );
    not g12685 ( n24789 , n22291 );
    and g12686 ( n16019 , n33402 , n7305 );
    xnor g12687 ( n24936 , n15007 , n21989 );
    xnor g12688 ( n28047 , n8965 , n11455 );
    not g12689 ( n33874 , n34563 );
    xnor g12690 ( n11544 , n6364 , n25647 );
    xnor g12691 ( n4277 , n20586 , n5234 );
    xnor g12692 ( n31101 , n682 , n32584 );
    xnor g12693 ( n31052 , n9426 , n33149 );
    or g12694 ( n25200 , n13546 , n9951 );
    xnor g12695 ( n33104 , n6392 , n31799 );
    or g12696 ( n379 , n26707 , n27801 );
    xor g12697 ( n21317 , n28044 , n28568 );
    or g12698 ( n19366 , n31363 , n20318 );
    and g12699 ( n18272 , n355 , n23123 );
    xnor g12700 ( n15162 , n17186 , n22158 );
    and g12701 ( n15899 , n19021 , n8023 );
    or g12702 ( n19514 , n35715 , n7232 );
    buf g12703 ( n30459 , n9449 );
    or g12704 ( n11883 , n30735 , n22961 );
    and g12705 ( n31775 , n35471 , n33904 );
    or g12706 ( n10584 , n18500 , n26468 );
    or g12707 ( n25759 , n10635 , n7032 );
    or g12708 ( n30811 , n31559 , n19271 );
    or g12709 ( n14079 , n835 , n2235 );
    nor g12710 ( n34091 , n17568 , n12809 );
    nor g12711 ( n9289 , n22291 , n24608 );
    and g12712 ( n33277 , n29347 , n24401 );
    nor g12713 ( n33884 , n25602 , n18651 );
    xnor g12714 ( n16537 , n12949 , n17751 );
    or g12715 ( n25187 , n2665 , n17037 );
    or g12716 ( n2731 , n1990 , n5618 );
    or g12717 ( n27855 , n17985 , n2680 );
    xnor g12718 ( n10691 , n33838 , n8465 );
    or g12719 ( n22509 , n15426 , n30519 );
    and g12720 ( n26126 , n15556 , n3526 );
    or g12721 ( n34445 , n33249 , n5346 );
    and g12722 ( n31161 , n33514 , n21913 );
    and g12723 ( n14584 , n13738 , n24916 );
    xnor g12724 ( n19488 , n18318 , n22819 );
    or g12725 ( n14008 , n11341 , n36000 );
    and g12726 ( n5396 , n2450 , n32894 );
    or g12727 ( n18604 , n31731 , n2237 );
    and g12728 ( n21349 , n2100 , n8709 );
    not g12729 ( n35756 , n19551 );
    buf g12730 ( n27625 , n2712 );
    xnor g12731 ( n18493 , n29188 , n4758 );
    xnor g12732 ( n796 , n6004 , n29236 );
    or g12733 ( n30572 , n25172 , n13305 );
    or g12734 ( n28019 , n24148 , n17065 );
    or g12735 ( n4795 , n21650 , n4550 );
    xnor g12736 ( n16685 , n25933 , n17553 );
    or g12737 ( n4697 , n23603 , n1252 );
    or g12738 ( n29466 , n16775 , n10140 );
    or g12739 ( n32523 , n31799 , n11034 );
    and g12740 ( n21990 , n22230 , n13009 );
    or g12741 ( n22155 , n7800 , n9174 );
    xnor g12742 ( n23644 , n5394 , n13008 );
    xnor g12743 ( n8081 , n15156 , n23512 );
    or g12744 ( n5037 , n35929 , n24102 );
    or g12745 ( n20523 , n8211 , n14523 );
    buf g12746 ( n35244 , n24338 );
    or g12747 ( n20144 , n34301 , n10872 );
    xnor g12748 ( n3773 , n30374 , n23773 );
    and g12749 ( n3584 , n29004 , n35997 );
    xnor g12750 ( n517 , n24872 , n29897 );
    or g12751 ( n709 , n7796 , n17976 );
    or g12752 ( n17362 , n948 , n908 );
    or g12753 ( n12619 , n4960 , n18087 );
    or g12754 ( n25345 , n3363 , n23249 );
    xnor g12755 ( n25245 , n32997 , n9164 );
    or g12756 ( n22133 , n5830 , n20812 );
    xnor g12757 ( n7972 , n77 , n20805 );
    or g12758 ( n23941 , n2546 , n21956 );
    or g12759 ( n46 , n4288 , n24086 );
    xnor g12760 ( n29187 , n16955 , n19261 );
    nor g12761 ( n31883 , n3251 , n3417 );
    or g12762 ( n26873 , n17648 , n18490 );
    and g12763 ( n9933 , n26935 , n13111 );
    xnor g12764 ( n5793 , n20426 , n95 );
    xnor g12765 ( n32286 , n13799 , n25744 );
    and g12766 ( n12683 , n25279 , n16188 );
    or g12767 ( n24072 , n16206 , n15507 );
    not g12768 ( n34450 , n3259 );
    not g12769 ( n28989 , n25602 );
    or g12770 ( n27314 , n28045 , n15506 );
    or g12771 ( n35689 , n20368 , n20762 );
    not g12772 ( n17944 , n23509 );
    or g12773 ( n20623 , n35806 , n10978 );
    or g12774 ( n21773 , n5287 , n4196 );
    or g12775 ( n9035 , n19835 , n4203 );
    xnor g12776 ( n32770 , n4604 , n31215 );
    or g12777 ( n25641 , n10362 , n24479 );
    and g12778 ( n32417 , n14868 , n13279 );
    buf g12779 ( n35935 , n15033 );
    xnor g12780 ( n19856 , n34262 , n9316 );
    or g12781 ( n27900 , n30739 , n24555 );
    xnor g12782 ( n16988 , n13745 , n22291 );
    or g12783 ( n31885 , n18160 , n2960 );
    xnor g12784 ( n28117 , n23439 , n32457 );
    xnor g12785 ( n21551 , n17157 , n21192 );
    and g12786 ( n11351 , n23227 , n14491 );
    not g12787 ( n28444 , n3394 );
    or g12788 ( n17263 , n5428 , n9675 );
    and g12789 ( n24534 , n35480 , n32891 );
    and g12790 ( n16583 , n15571 , n30508 );
    not g12791 ( n22782 , n34521 );
    and g12792 ( n30070 , n12750 , n32985 );
    not g12793 ( n21149 , n30333 );
    or g12794 ( n18942 , n1391 , n19105 );
    or g12795 ( n4584 , n27875 , n7072 );
    and g12796 ( n15828 , n3007 , n19372 );
    not g12797 ( n32191 , n3205 );
    and g12798 ( n8405 , n8573 , n8726 );
    or g12799 ( n2987 , n28562 , n35630 );
    or g12800 ( n17617 , n13414 , n33098 );
    or g12801 ( n25180 , n19922 , n26675 );
    or g12802 ( n31825 , n21466 , n18767 );
    or g12803 ( n24767 , n364 , n6950 );
    xnor g12804 ( n4677 , n13753 , n6625 );
    not g12805 ( n9021 , n17568 );
    and g12806 ( n3144 , n15932 , n21557 );
    xnor g12807 ( n24206 , n16857 , n34999 );
    and g12808 ( n3800 , n4806 , n9343 );
    nor g12809 ( n8165 , n22953 , n33155 );
    xnor g12810 ( n24909 , n1551 , n1980 );
    and g12811 ( n22944 , n2026 , n80 );
    and g12812 ( n13595 , n14460 , n19138 );
    and g12813 ( n22213 , n13994 , n20223 );
    not g12814 ( n15074 , n25943 );
    or g12815 ( n35418 , n7540 , n10761 );
    or g12816 ( n15729 , n20638 , n12510 );
    or g12817 ( n20622 , n12582 , n11827 );
    and g12818 ( n19462 , n29725 , n29663 );
    or g12819 ( n2853 , n28292 , n28574 );
    nor g12820 ( n29127 , n13705 , n23325 );
    xnor g12821 ( n34914 , n25441 , n25638 );
    xnor g12822 ( n4262 , n14340 , n3222 );
    and g12823 ( n15305 , n25876 , n12204 );
    xnor g12824 ( n21072 , n18426 , n32095 );
    and g12825 ( n5172 , n3544 , n24188 );
    and g12826 ( n17265 , n13474 , n25484 );
    and g12827 ( n16858 , n5142 , n21860 );
    xnor g12828 ( n32916 , n25813 , n25307 );
    xnor g12829 ( n12267 , n6937 , n1950 );
    or g12830 ( n14502 , n16650 , n4895 );
    and g12831 ( n9448 , n2848 , n18166 );
    xnor g12832 ( n23694 , n5696 , n9658 );
    or g12833 ( n13983 , n13704 , n7525 );
    and g12834 ( n3895 , n5068 , n33971 );
    and g12835 ( n32031 , n1800 , n22121 );
    or g12836 ( n20218 , n10894 , n4608 );
    and g12837 ( n32276 , n34340 , n11304 );
    or g12838 ( n23897 , n12542 , n6950 );
    and g12839 ( n4536 , n8718 , n25050 );
    not g12840 ( n27559 , n25110 );
    nor g12841 ( n9404 , n30189 , n13222 );
    or g12842 ( n13022 , n169 , n32697 );
    or g12843 ( n11052 , n6145 , n3188 );
    and g12844 ( n1983 , n24642 , n11480 );
    or g12845 ( n27478 , n7098 , n23921 );
    and g12846 ( n11077 , n963 , n9948 );
    not g12847 ( n20957 , n17568 );
    or g12848 ( n9561 , n5917 , n1176 );
    or g12849 ( n35908 , n19789 , n27501 );
    xnor g12850 ( n33439 , n20223 , n13994 );
    or g12851 ( n14508 , n4288 , n16841 );
    xor g12852 ( n12935 , n25553 , n21069 );
    and g12853 ( n5493 , n35126 , n16437 );
    and g12854 ( n35186 , n12974 , n47 );
    or g12855 ( n25323 , n7719 , n22634 );
    xnor g12856 ( n11485 , n19628 , n35927 );
    xnor g12857 ( n26812 , n22815 , n22377 );
    or g12858 ( n5846 , n20413 , n3188 );
    buf g12859 ( n23921 , n2658 );
    or g12860 ( n32798 , n21705 , n4311 );
    or g12861 ( n23075 , n23731 , n29411 );
    or g12862 ( n6260 , n20929 , n19335 );
    or g12863 ( n26427 , n3702 , n6075 );
    nor g12864 ( n1878 , n32967 , n19968 );
    or g12865 ( n11043 , n4962 , n4981 );
    or g12866 ( n31845 , n15148 , n20579 );
    or g12867 ( n17348 , n18610 , n30708 );
    or g12868 ( n28994 , n5706 , n11570 );
    or g12869 ( n12665 , n942 , n31116 );
    and g12870 ( n33799 , n35984 , n34407 );
    and g12871 ( n23269 , n9285 , n11809 );
    or g12872 ( n2219 , n23968 , n20552 );
    or g12873 ( n16126 , n11338 , n2117 );
    or g12874 ( n17023 , n31559 , n4893 );
    and g12875 ( n15917 , n31479 , n25118 );
    buf g12876 ( n18115 , n31411 );
    xnor g12877 ( n3669 , n27549 , n34682 );
    or g12878 ( n17144 , n35224 , n31833 );
    or g12879 ( n34986 , n4732 , n26381 );
    xnor g12880 ( n32226 , n34697 , n16620 );
    and g12881 ( n15376 , n35122 , n4902 );
    or g12882 ( n32677 , n9321 , n21962 );
    xnor g12883 ( n20941 , n20331 , n16417 );
    and g12884 ( n19476 , n26059 , n19865 );
    and g12885 ( n30944 , n13116 , n14257 );
    xnor g12886 ( n22491 , n29942 , n19551 );
    and g12887 ( n23277 , n32070 , n22107 );
    or g12888 ( n577 , n24371 , n22135 );
    and g12889 ( n22381 , n25942 , n31831 );
    and g12890 ( n4938 , n6329 , n28812 );
    or g12891 ( n33769 , n9789 , n6402 );
    and g12892 ( n18795 , n27790 , n10879 );
    xnor g12893 ( n30244 , n7661 , n31104 );
    and g12894 ( n14146 , n7083 , n28326 );
    or g12895 ( n23548 , n22291 , n17353 );
    xnor g12896 ( n18779 , n10660 , n34749 );
    not g12897 ( n5338 , n30459 );
    or g12898 ( n33392 , n18013 , n17102 );
    or g12899 ( n6546 , n1380 , n24811 );
    or g12900 ( n28983 , n5359 , n16525 );
    or g12901 ( n18025 , n9010 , n35935 );
    or g12902 ( n6983 , n3141 , n106 );
    xnor g12903 ( n20051 , n27843 , n19141 );
    and g12904 ( n18665 , n16695 , n20373 );
    nor g12905 ( n22966 , n1836 , n12731 );
    and g12906 ( n2706 , n10332 , n1059 );
    and g12907 ( n12269 , n18093 , n35001 );
    nor g12908 ( n22707 , n14616 , n19115 );
    and g12909 ( n20292 , n24252 , n3204 );
    or g12910 ( n24543 , n9793 , n20101 );
    or g12911 ( n2520 , n27258 , n32579 );
    and g12912 ( n9883 , n10215 , n25206 );
    xnor g12913 ( n2688 , n2421 , n15110 );
    or g12914 ( n34753 , n31799 , n23065 );
    or g12915 ( n30377 , n17751 , n33027 );
    and g12916 ( n1377 , n10925 , n31510 );
    xnor g12917 ( n5029 , n15928 , n25174 );
    or g12918 ( n26026 , n24249 , n9709 );
    not g12919 ( n35481 , n34476 );
    and g12920 ( n31948 , n11863 , n14030 );
    or g12921 ( n13131 , n19477 , n12428 );
    and g12922 ( n3784 , n34307 , n21085 );
    not g12923 ( n27146 , n21657 );
    xnor g12924 ( n4534 , n20435 , n20654 );
    or g12925 ( n26655 , n13893 , n21210 );
    or g12926 ( n14705 , n15403 , n13862 );
    or g12927 ( n13095 , n17353 , n24489 );
    or g12928 ( n14369 , n4517 , n28438 );
    xnor g12929 ( n13133 , n28924 , n6266 );
    not g12930 ( n16668 , n30586 );
    and g12931 ( n11741 , n20307 , n26400 );
    or g12932 ( n22625 , n17568 , n27060 );
    or g12933 ( n17066 , n33367 , n25183 );
    or g12934 ( n16359 , n9789 , n32834 );
    xnor g12935 ( n12410 , n23067 , n20959 );
    or g12936 ( n32429 , n25878 , n29854 );
    or g12937 ( n19242 , n10894 , n8974 );
    or g12938 ( n3000 , n35927 , n16310 );
    nor g12939 ( n23429 , n16620 , n24218 );
    xnor g12940 ( n13281 , n20356 , n7141 );
    and g12941 ( n16000 , n35055 , n26863 );
    not g12942 ( n33677 , n12622 );
    and g12943 ( n30233 , n11560 , n9970 );
    and g12944 ( n19259 , n23944 , n23454 );
    xnor g12945 ( n26649 , n555 , n9793 );
    or g12946 ( n1024 , n28154 , n2798 );
    xnor g12947 ( n29122 , n16857 , n20847 );
    xnor g12948 ( n20477 , n5960 , n9658 );
    xnor g12949 ( n27224 , n7139 , n29884 );
    xnor g12950 ( n11251 , n10333 , n16893 );
    or g12951 ( n32085 , n19462 , n18255 );
    nor g12952 ( n20252 , n24376 , n26369 );
    and g12953 ( n1340 , n24614 , n27982 );
    and g12954 ( n22657 , n32631 , n29820 );
    or g12955 ( n23476 , n17539 , n26172 );
    xnor g12956 ( n31800 , n13358 , n21554 );
    or g12957 ( n34233 , n33837 , n7673 );
    nor g12958 ( n2262 , n24016 , n27359 );
    and g12959 ( n14640 , n20969 , n31206 );
    and g12960 ( n7147 , n18079 , n592 );
    or g12961 ( n19541 , n19163 , n30507 );
    or g12962 ( n3714 , n15403 , n23764 );
    or g12963 ( n19226 , n18918 , n31554 );
    and g12964 ( n21301 , n25660 , n29958 );
    and g12965 ( n32476 , n23009 , n12760 );
    or g12966 ( n5828 , n22914 , n26931 );
    and g12967 ( n22777 , n4601 , n5405 );
    xnor g12968 ( n27817 , n3675 , n24226 );
    and g12969 ( n6741 , n661 , n1672 );
    xnor g12970 ( n29895 , n12338 , n27527 );
    or g12971 ( n10600 , n22320 , n25752 );
    or g12972 ( n28872 , n12801 , n25831 );
    or g12973 ( n26262 , n1836 , n30884 );
    and g12974 ( n21680 , n7513 , n29567 );
    and g12975 ( n5590 , n26305 , n34220 );
    or g12976 ( n29642 , n1774 , n3279 );
    xnor g12977 ( n7294 , n10454 , n6714 );
    xnor g12978 ( n7119 , n9481 , n14283 );
    xnor g12979 ( n34606 , n22747 , n29839 );
    and g12980 ( n23211 , n30593 , n9651 );
    xnor g12981 ( n32915 , n31619 , n17568 );
    xnor g12982 ( n23958 , n13544 , n6321 );
    nor g12983 ( n23776 , n19085 , n25322 );
    or g12984 ( n26300 , n9658 , n27362 );
    not g12985 ( n20425 , n30879 );
    and g12986 ( n16566 , n25077 , n21445 );
    or g12987 ( n156 , n1963 , n29963 );
    and g12988 ( n2276 , n12754 , n11037 );
    not g12989 ( n31887 , n25392 );
    or g12990 ( n23984 , n2708 , n35757 );
    and g12991 ( n1072 , n6928 , n5897 );
    not g12992 ( n33622 , n4962 );
    not g12993 ( n7863 , n15842 );
    or g12994 ( n10273 , n22001 , n24672 );
    not g12995 ( n1462 , n27792 );
    or g12996 ( n31766 , n12707 , n30762 );
    or g12997 ( n1809 , n22177 , n27053 );
    or g12998 ( n7974 , n1269 , n1796 );
    nor g12999 ( n15460 , n10894 , n23026 );
    xnor g13000 ( n32792 , n2992 , n3222 );
    or g13001 ( n26027 , n31799 , n4123 );
    xnor g13002 ( n21247 , n15973 , n23450 );
    or g13003 ( n27709 , n31881 , n9601 );
    or g13004 ( n33500 , n1131 , n12879 );
    not g13005 ( n2600 , n16659 );
    and g13006 ( n18102 , n29479 , n8169 );
    or g13007 ( n12420 , n35227 , n34865 );
    or g13008 ( n951 , n17278 , n25255 );
    not g13009 ( n27588 , n8644 );
    or g13010 ( n24045 , n23252 , n7673 );
    and g13011 ( n14973 , n13184 , n6862 );
    or g13012 ( n5624 , n20719 , n8024 );
    or g13013 ( n18153 , n18258 , n24710 );
    xnor g13014 ( n6405 , n1477 , n34481 );
    not g13015 ( n11633 , n11307 );
    and g13016 ( n22224 , n13599 , n33644 );
    and g13017 ( n27824 , n30172 , n8822 );
    and g13018 ( n23185 , n18314 , n13091 );
    not g13019 ( n16411 , n34022 );
    not g13020 ( n3497 , n20185 );
    not g13021 ( n26949 , n34319 );
    nor g13022 ( n14517 , n5374 , n734 );
    xnor g13023 ( n29957 , n7912 , n28032 );
    and g13024 ( n1119 , n17538 , n22936 );
    xnor g13025 ( n3202 , n17267 , n16135 );
    or g13026 ( n6630 , n4288 , n13562 );
    xnor g13027 ( n1062 , n15006 , n16307 );
    buf g13028 ( n915 , n11379 );
    or g13029 ( n31073 , n14223 , n17906 );
    or g13030 ( n32960 , n5408 , n3882 );
    and g13031 ( n8191 , n10224 , n16574 );
    nor g13032 ( n4395 , n19984 , n33467 );
    or g13033 ( n23145 , n16539 , n15538 );
    xnor g13034 ( n14063 , n2639 , n24651 );
    and g13035 ( n6469 , n21260 , n14189 );
    or g13036 ( n31320 , n24332 , n22914 );
    xnor g13037 ( n15206 , n24932 , n29759 );
    or g13038 ( n10202 , n7319 , n4203 );
    nor g13039 ( n10334 , n3222 , n28546 );
    xnor g13040 ( n34320 , n20387 , n16922 );
    nor g13041 ( n7788 , n22503 , n14845 );
    and g13042 ( n14623 , n8410 , n29435 );
    and g13043 ( n2667 , n24003 , n35743 );
    xnor g13044 ( n2902 , n15941 , n21684 );
    nor g13045 ( n34281 , n29839 , n23906 );
    or g13046 ( n4000 , n17568 , n24121 );
    nor g13047 ( n35483 , n27226 , n9550 );
    or g13048 ( n1300 , n28981 , n34971 );
    xnor g13049 ( n7930 , n15752 , n4960 );
    nor g13050 ( n2187 , n830 , n24024 );
    or g13051 ( n14911 , n22201 , n6052 );
    or g13052 ( n7841 , n13024 , n6306 );
    xnor g13053 ( n34705 , n27919 , n32857 );
    xnor g13054 ( n9100 , n2393 , n21531 );
    xnor g13055 ( n12161 , n10149 , n24382 );
    xnor g13056 ( n18257 , n34244 , n9867 );
    or g13057 ( n1804 , n14225 , n10651 );
    not g13058 ( n14812 , n1528 );
    xnor g13059 ( n18835 , n27089 , n25174 );
    or g13060 ( n26469 , n12780 , n32507 );
    not g13061 ( n21240 , n26725 );
    buf g13062 ( n31067 , n17111 );
    or g13063 ( n14914 , n31289 , n10003 );
    or g13064 ( n18271 , n6617 , n32185 );
    xnor g13065 ( n33090 , n1256 , n31289 );
    nor g13066 ( n29003 , n21775 , n20642 );
    and g13067 ( n1087 , n34435 , n4383 );
    and g13068 ( n1922 , n14092 , n2793 );
    and g13069 ( n23608 , n5225 , n24982 );
    and g13070 ( n32593 , n27776 , n31061 );
    and g13071 ( n6837 , n22711 , n4071 );
    or g13072 ( n249 , n3946 , n31812 );
    or g13073 ( n6747 , n16111 , n17815 );
    not g13074 ( n4683 , n33171 );
    nor g13075 ( n30230 , n830 , n16716 );
    nor g13076 ( n17248 , n20247 , n6017 );
    xnor g13077 ( n32168 , n15731 , n17751 );
    or g13078 ( n19194 , n18722 , n7514 );
    or g13079 ( n9770 , n33136 , n19464 );
    or g13080 ( n29345 , n24332 , n21271 );
    or g13081 ( n20522 , n28560 , n33310 );
    and g13082 ( n14436 , n21592 , n29726 );
    or g13083 ( n19944 , n608 , n24505 );
    or g13084 ( n21269 , n16283 , n16903 );
    xnor g13085 ( n15856 , n33373 , n18379 );
    or g13086 ( n24226 , n12032 , n8474 );
    nor g13087 ( n15686 , n9789 , n6980 );
    and g13088 ( n27587 , n8411 , n1159 );
    or g13089 ( n18187 , n2688 , n21579 );
    not g13090 ( n9344 , n30117 );
    xnor g13091 ( n8697 , n18651 , n8524 );
    xnor g13092 ( n12276 , n28564 , n15886 );
    and g13093 ( n17024 , n22161 , n9913 );
    or g13094 ( n10835 , n16693 , n34852 );
    or g13095 ( n14050 , n26732 , n19084 );
    or g13096 ( n6967 , n31559 , n12844 );
    and g13097 ( n12883 , n30072 , n8964 );
    xnor g13098 ( n31086 , n32735 , n16922 );
    or g13099 ( n24307 , n2508 , n19793 );
    or g13100 ( n23105 , n27397 , n22501 );
    and g13101 ( n1048 , n19701 , n24958 );
    or g13102 ( n12293 , n16481 , n34727 );
    and g13103 ( n19496 , n21308 , n6262 );
    and g13104 ( n15889 , n25323 , n7688 );
    and g13105 ( n2753 , n13606 , n30356 );
    and g13106 ( n10918 , n1310 , n30303 );
    not g13107 ( n32481 , n29331 );
    and g13108 ( n23169 , n19279 , n7922 );
    or g13109 ( n29244 , n174 , n24025 );
    nor g13110 ( n12032 , n15886 , n26441 );
    xnor g13111 ( n15356 , n17026 , n17405 );
    and g13112 ( n10407 , n18178 , n2021 );
    buf g13113 ( n24259 , n14706 );
    or g13114 ( n8309 , n4758 , n7733 );
    buf g13115 ( n31549 , n16919 );
    nor g13116 ( n19493 , n19142 , n12702 );
    not g13117 ( n15002 , n2029 );
    and g13118 ( n19901 , n12733 , n31343 );
    xnor g13119 ( n21359 , n3125 , n2548 );
    and g13120 ( n3111 , n1949 , n15971 );
    or g13121 ( n9182 , n6297 , n20797 );
    or g13122 ( n11531 , n7745 , n20308 );
    or g13123 ( n12270 , n9667 , n8362 );
    and g13124 ( n32590 , n32381 , n28428 );
    and g13125 ( n21073 , n20093 , n25118 );
    or g13126 ( n19616 , n20790 , n16659 );
    or g13127 ( n29996 , n27605 , n22961 );
    and g13128 ( n23393 , n7548 , n2129 );
    or g13129 ( n32787 , n32370 , n1942 );
    nor g13130 ( n18092 , n9658 , n35936 );
    and g13131 ( n18672 , n6099 , n27723 );
    not g13132 ( n25711 , n15403 );
    xnor g13133 ( n14090 , n25269 , n33706 );
    or g13134 ( n7890 , n32095 , n3917 );
    or g13135 ( n22758 , n10678 , n12298 );
    and g13136 ( n24455 , n34067 , n9778 );
    xnor g13137 ( n5557 , n13716 , n15393 );
    or g13138 ( n33472 , n29713 , n30373 );
    xnor g13139 ( n7285 , n33529 , n830 );
    and g13140 ( n18309 , n30547 , n27131 );
    or g13141 ( n32850 , n4604 , n2712 );
    or g13142 ( n34215 , n19530 , n9317 );
    not g13143 ( n3492 , n19418 );
    and g13144 ( n1015 , n33225 , n18228 );
    not g13145 ( n19090 , n31559 );
    or g13146 ( n30585 , n5089 , n17125 );
    nor g13147 ( n17934 , n12507 , n30871 );
    and g13148 ( n3921 , n19381 , n25939 );
    not g13149 ( n5729 , n8966 );
    nor g13150 ( n24579 , n27383 , n19834 );
    or g13151 ( n34787 , n25679 , n25036 );
    nor g13152 ( n1839 , n11955 , n2535 );
    and g13153 ( n16212 , n906 , n13582 );
    or g13154 ( n7257 , n19551 , n18106 );
    or g13155 ( n20261 , n29839 , n550 );
    or g13156 ( n15175 , n4447 , n10319 );
    and g13157 ( n4449 , n9315 , n28019 );
    or g13158 ( n31338 , n19129 , n12668 );
    or g13159 ( n15236 , n29839 , n8988 );
    not g13160 ( n5989 , n3417 );
    and g13161 ( n5190 , n6562 , n28375 );
    xnor g13162 ( n4300 , n17696 , n1516 );
    or g13163 ( n26718 , n16161 , n21339 );
    or g13164 ( n18417 , n16035 , n28606 );
    or g13165 ( n7132 , n11046 , n7250 );
    and g13166 ( n29176 , n34470 , n35438 );
    or g13167 ( n32568 , n24156 , n8619 );
    nor g13168 ( n21634 , n29501 , n28113 );
    and g13169 ( n32366 , n18842 , n34477 );
    or g13170 ( n33563 , n30386 , n30708 );
    or g13171 ( n29613 , n23594 , n3694 );
    or g13172 ( n33807 , n9120 , n2728 );
    not g13173 ( n17007 , n12098 );
    or g13174 ( n25443 , n28830 , n24653 );
    and g13175 ( n32816 , n22452 , n21836 );
    nor g13176 ( n25915 , n7048 , n4657 );
    nor g13177 ( n26479 , n5287 , n5089 );
    or g13178 ( n20270 , n8198 , n6975 );
    or g13179 ( n26889 , n29306 , n9317 );
    nor g13180 ( n8517 , n7779 , n18115 );
    or g13181 ( n27129 , n4035 , n16797 );
    nor g13182 ( n13992 , n31799 , n13229 );
    or g13183 ( n16376 , n18599 , n15154 );
    not g13184 ( n4439 , n22241 );
    or g13185 ( n15647 , n9057 , n23323 );
    and g13186 ( n18874 , n10440 , n9525 );
    buf g13187 ( n4175 , n25031 );
    xnor g13188 ( n12443 , n32535 , n17751 );
    nor g13189 ( n24347 , n9793 , n2342 );
    and g13190 ( n16387 , n12694 , n26131 );
    or g13191 ( n13530 , n27736 , n19490 );
    or g13192 ( n6849 , n11995 , n27625 );
    and g13193 ( n22734 , n26893 , n35103 );
    xnor g13194 ( n2208 , n19097 , n35800 );
    and g13195 ( n7112 , n1674 , n18042 );
    xnor g13196 ( n31594 , n33346 , n25174 );
    or g13197 ( n29684 , n30282 , n4318 );
    or g13198 ( n16483 , n9789 , n19328 );
    or g13199 ( n22180 , n16172 , n1924 );
    xnor g13200 ( n7509 , n302 , n24088 );
    xnor g13201 ( n18436 , n34992 , n26698 );
    xnor g13202 ( n30820 , n5374 , n734 );
    or g13203 ( n10129 , n4427 , n10583 );
    or g13204 ( n23937 , n35250 , n4244 );
    xnor g13205 ( n13048 , n13456 , n16922 );
    and g13206 ( n1852 , n34775 , n23629 );
    or g13207 ( n7656 , n28698 , n19410 );
    and g13208 ( n13770 , n3851 , n5712 );
    or g13209 ( n14935 , n4286 , n17872 );
    xnor g13210 ( n9228 , n32202 , n23604 );
    or g13211 ( n5251 , n33090 , n12203 );
    xnor g13212 ( n15276 , n22479 , n8855 );
    and g13213 ( n33545 , n12933 , n23647 );
    xnor g13214 ( n23912 , n19041 , n4664 );
    or g13215 ( n1397 , n15728 , n20147 );
    and g13216 ( n3553 , n30153 , n21406 );
    nor g13217 ( n32933 , n15886 , n14643 );
    xnor g13218 ( n15409 , n22483 , n31056 );
    or g13219 ( n6213 , n4288 , n26449 );
    nor g13220 ( n10962 , n16531 , n6204 );
    or g13221 ( n16085 , n19551 , n9386 );
    or g13222 ( n24522 , n18748 , n20664 );
    and g13223 ( n24842 , n22219 , n26684 );
    or g13224 ( n3011 , n10371 , n31143 );
    or g13225 ( n13431 , n32187 , n26929 );
    and g13226 ( n1682 , n35602 , n20951 );
    and g13227 ( n12743 , n11098 , n2268 );
    xnor g13228 ( n9885 , n11743 , n19551 );
    or g13229 ( n30441 , n27196 , n27203 );
    or g13230 ( n15072 , n17729 , n3736 );
    or g13231 ( n11767 , n31392 , n25255 );
    or g13232 ( n12766 , n13112 , n12879 );
    not g13233 ( n24299 , n15290 );
    xnor g13234 ( n15406 , n7978 , n3205 );
    xnor g13235 ( n29326 , n26004 , n27226 );
    nor g13236 ( n28170 , n1578 , n33956 );
    and g13237 ( n12448 , n19716 , n33912 );
    not g13238 ( n21018 , n22980 );
    or g13239 ( n26661 , n30665 , n1715 );
    or g13240 ( n35085 , n35983 , n29356 );
    and g13241 ( n8088 , n33710 , n4780 );
    or g13242 ( n30388 , n20688 , n31784 );
    or g13243 ( n20006 , n32224 , n15290 );
    not g13244 ( n29350 , n1843 );
    or g13245 ( n30570 , n14343 , n28438 );
    and g13246 ( n16631 , n30165 , n17599 );
    xor g13247 ( n33390 , n21287 , n18412 );
    xnor g13248 ( n23439 , n27742 , n3946 );
    xnor g13249 ( n29742 , n3551 , n33923 );
    or g13250 ( n12633 , n23970 , n23593 );
    not g13251 ( n35401 , n22980 );
    nor g13252 ( n11670 , n9789 , n11787 );
    xnor g13253 ( n66 , n5218 , n31587 );
    xnor g13254 ( n29865 , n23017 , n5404 );
    xnor g13255 ( n23055 , n1891 , n18097 );
    and g13256 ( n36046 , n29563 , n24541 );
    or g13257 ( n28805 , n21279 , n9394 );
    not g13258 ( n237 , n17854 );
    xnor g13259 ( n13586 , n27738 , n10235 );
    nor g13260 ( n24937 , n9795 , n19215 );
    xnor g13261 ( n18125 , n34334 , n3725 );
    xnor g13262 ( n28736 , n17175 , n24294 );
    or g13263 ( n24386 , n24332 , n3177 );
    nor g13264 ( n31564 , n1611 , n15599 );
    or g13265 ( n17541 , n2197 , n35043 );
    or g13266 ( n2289 , n5115 , n29626 );
    or g13267 ( n197 , n14605 , n29393 );
    or g13268 ( n5914 , n14788 , n9832 );
    nor g13269 ( n28389 , n31765 , n4496 );
    and g13270 ( n9556 , n12454 , n34636 );
    nor g13271 ( n32182 , n29856 , n27199 );
    or g13272 ( n7008 , n3290 , n12679 );
    and g13273 ( n15914 , n20317 , n28268 );
    or g13274 ( n31379 , n25871 , n23090 );
    and g13275 ( n15371 , n35996 , n18250 );
    not g13276 ( n1956 , n19615 );
    not g13277 ( n4996 , n5147 );
    or g13278 ( n2403 , n4262 , n17050 );
    not g13279 ( n11142 , n21832 );
    or g13280 ( n15392 , n24840 , n763 );
    nor g13281 ( n10950 , n20392 , n20917 );
    or g13282 ( n18595 , n26021 , n26443 );
    or g13283 ( n6350 , n10112 , n28787 );
    xnor g13284 ( n28929 , n23270 , n4962 );
    or g13285 ( n31288 , n2304 , n20690 );
    or g13286 ( n5347 , n11590 , n25306 );
    and g13287 ( n935 , n15229 , n23868 );
    and g13288 ( n26332 , n3110 , n26571 );
    or g13289 ( n34877 , n31895 , n29640 );
    and g13290 ( n24048 , n21023 , n20735 );
    xnor g13291 ( n26041 , n10529 , n4878 );
    not g13292 ( n14473 , n29609 );
    not g13293 ( n17140 , n31799 );
    or g13294 ( n726 , n1718 , n11977 );
    nor g13295 ( n31424 , n1950 , n32239 );
    and g13296 ( n7937 , n25598 , n28382 );
    or g13297 ( n27932 , n31216 , n23735 );
    and g13298 ( n36045 , n789 , n27972 );
    xnor g13299 ( n13112 , n129 , n21771 );
    xnor g13300 ( n32445 , n647 , n24371 );
    or g13301 ( n7604 , n14031 , n3088 );
    or g13302 ( n22507 , n22291 , n4957 );
    or g13303 ( n15386 , n990 , n3708 );
    or g13304 ( n3983 , n24550 , n11703 );
    or g13305 ( n27285 , n29283 , n33694 );
    not g13306 ( n34254 , n25602 );
    and g13307 ( n7621 , n31721 , n10103 );
    or g13308 ( n15016 , n8432 , n5117 );
    xnor g13309 ( n4856 , n35697 , n16620 );
    or g13310 ( n4958 , n4809 , n24220 );
    or g13311 ( n36063 , n23550 , n10031 );
    nor g13312 ( n14625 , n16938 , n16976 );
    xnor g13313 ( n2404 , n8374 , n26306 );
    or g13314 ( n2000 , n15473 , n28100 );
    and g13315 ( n35815 , n25865 , n5927 );
    xnor g13316 ( n28265 , n23979 , n16739 );
    and g13317 ( n28939 , n32815 , n25175 );
    nor g13318 ( n21188 , n31829 , n25153 );
    nor g13319 ( n33117 , n6225 , n32982 );
    xnor g13320 ( n23386 , n27224 , n20441 );
    or g13321 ( n9230 , n4007 , n19241 );
    or g13322 ( n20423 , n29270 , n8567 );
    or g13323 ( n32761 , n29839 , n29139 );
    and g13324 ( n33529 , n10684 , n14701 );
    or g13325 ( n17937 , n9793 , n11424 );
    or g13326 ( n30443 , n12138 , n15109 );
    or g13327 ( n31463 , n25218 , n23981 );
    xnor g13328 ( n21118 , n24136 , n31823 );
    xnor g13329 ( n34178 , n10454 , n23804 );
    nor g13330 ( n954 , n3205 , n34203 );
    xnor g13331 ( n31212 , n11569 , n29839 );
    or g13332 ( n18729 , n4962 , n5584 );
    or g13333 ( n16604 , n10767 , n5168 );
    and g13334 ( n6051 , n15335 , n20019 );
    nor g13335 ( n26699 , n11455 , n6527 );
    or g13336 ( n17700 , n2489 , n11104 );
    and g13337 ( n30611 , n34088 , n2656 );
    or g13338 ( n31522 , n751 , n10670 );
    or g13339 ( n20754 , n11776 , n33401 );
    and g13340 ( n2124 , n16739 , n23979 );
    or g13341 ( n28000 , n18994 , n32557 );
    or g13342 ( n31663 , n19112 , n31696 );
    or g13343 ( n20473 , n5920 , n22989 );
    and g13344 ( n2419 , n33815 , n34461 );
    or g13345 ( n12154 , n7671 , n10598 );
    not g13346 ( n28266 , n28099 );
    or g13347 ( n32352 , n10696 , n13307 );
    or g13348 ( n22795 , n30742 , n16324 );
    and g13349 ( n2683 , n6144 , n22389 );
    and g13350 ( n9288 , n4543 , n28010 );
    or g13351 ( n3879 , n7115 , n13480 );
    or g13352 ( n13644 , n15057 , n148 );
    or g13353 ( n12235 , n29839 , n22811 );
    not g13354 ( n25980 , n3171 );
    and g13355 ( n10822 , n12200 , n35063 );
    nor g13356 ( n32532 , n4960 , n22347 );
    xnor g13357 ( n26025 , n32811 , n4962 );
    or g13358 ( n21156 , n27291 , n16228 );
    or g13359 ( n24982 , n16925 , n18358 );
    nor g13360 ( n1124 , n1950 , n30097 );
    and g13361 ( n20692 , n29328 , n20509 );
    or g13362 ( n35638 , n32065 , n27801 );
    or g13363 ( n17209 , n31215 , n10758 );
    or g13364 ( n22804 , n3342 , n32572 );
    xnor g13365 ( n13107 , n19709 , n8941 );
    or g13366 ( n26149 , n6480 , n17162 );
    xnor g13367 ( n27399 , n21510 , n27291 );
    or g13368 ( n28589 , n7267 , n22807 );
    or g13369 ( n28097 , n33285 , n17974 );
    nor g13370 ( n23095 , n3205 , n13845 );
    or g13371 ( n31990 , n24400 , n35804 );
    or g13372 ( n32802 , n230 , n35402 );
    or g13373 ( n20304 , n17246 , n12953 );
    xnor g13374 ( n2079 , n27025 , n7993 );
    nor g13375 ( n26437 , n24245 , n19087 );
    xnor g13376 ( n28416 , n12247 , n35763 );
    xnor g13377 ( n29561 , n19524 , n4288 );
    or g13378 ( n211 , n21142 , n28866 );
    buf g13379 ( n29203 , n34588 );
    or g13380 ( n17460 , n29839 , n26760 );
    or g13381 ( n16957 , n4539 , n14746 );
    nor g13382 ( n11540 , n10813 , n33157 );
    xnor g13383 ( n3622 , n18498 , n5335 );
    xnor g13384 ( n5678 , n14387 , n32857 );
    and g13385 ( n11487 , n9766 , n7414 );
    or g13386 ( n26742 , n16922 , n8932 );
    xnor g13387 ( n32781 , n5194 , n17060 );
    or g13388 ( n15718 , n14921 , n22682 );
    xnor g13389 ( n9242 , n23658 , n18873 );
    and g13390 ( n1907 , n22659 , n8054 );
    or g13391 ( n10036 , n17609 , n34600 );
    and g13392 ( n15509 , n1620 , n17148 );
    xnor g13393 ( n2469 , n12643 , n33227 );
    and g13394 ( n4078 , n16011 , n1966 );
    buf g13395 ( n35143 , n29718 );
    not g13396 ( n2979 , n15344 );
    or g13397 ( n25283 , n34516 , n29592 );
    or g13398 ( n774 , n6604 , n27041 );
    or g13399 ( n28297 , n9277 , n31134 );
    or g13400 ( n24488 , n5703 , n23192 );
    and g13401 ( n34590 , n13212 , n34577 );
    or g13402 ( n16997 , n32857 , n9657 );
    and g13403 ( n22569 , n1945 , n5342 );
    or g13404 ( n28483 , n23132 , n29015 );
    xnor g13405 ( n18413 , n24326 , n23939 );
    or g13406 ( n29827 , n5493 , n5521 );
    or g13407 ( n20661 , n11670 , n27563 );
    or g13408 ( n29240 , n20198 , n14632 );
    and g13409 ( n11859 , n440 , n16605 );
    and g13410 ( n27094 , n20502 , n1699 );
    or g13411 ( n5202 , n29614 , n1642 );
    xnor g13412 ( n26325 , n16001 , n17827 );
    or g13413 ( n9286 , n8940 , n12428 );
    or g13414 ( n11275 , n2404 , n35141 );
    and g13415 ( n18297 , n20220 , n18116 );
    buf g13416 ( n24653 , n24022 );
    and g13417 ( n3961 , n14562 , n31813 );
    and g13418 ( n762 , n4777 , n21751 );
    xnor g13419 ( n12969 , n31906 , n5795 );
    or g13420 ( n23842 , n5388 , n8364 );
    or g13421 ( n26031 , n7195 , n16457 );
    and g13422 ( n21554 , n8864 , n12948 );
    or g13423 ( n1029 , n28827 , n31606 );
    or g13424 ( n30227 , n30092 , n4892 );
    xnor g13425 ( n26364 , n19001 , n4758 );
    nor g13426 ( n1653 , n11455 , n27979 );
    or g13427 ( n13342 , n27718 , n20120 );
    nor g13428 ( n11216 , n4960 , n6559 );
    and g13429 ( n17382 , n8360 , n20731 );
    nor g13430 ( n18979 , n19450 , n6548 );
    or g13431 ( n29541 , n1277 , n31334 );
    or g13432 ( n17122 , n31559 , n28004 );
    not g13433 ( n16849 , n30250 );
    and g13434 ( n3640 , n6492 , n3682 );
    xnor g13435 ( n16665 , n999 , n10721 );
    xnor g13436 ( n24324 , n25385 , n8076 );
    and g13437 ( n1565 , n13631 , n29170 );
    or g13438 ( n13371 , n1296 , n2117 );
    and g13439 ( n17409 , n25161 , n9570 );
    xnor g13440 ( n21098 , n31417 , n35326 );
    or g13441 ( n20551 , n8929 , n11258 );
    xnor g13442 ( n27807 , n18246 , n1097 );
    xnor g13443 ( n7424 , n30467 , n17751 );
    or g13444 ( n13780 , n1873 , n21554 );
    nor g13445 ( n6835 , n6596 , n33115 );
    and g13446 ( n33107 , n33196 , n15818 );
    or g13447 ( n2424 , n11368 , n22496 );
    or g13448 ( n26616 , n14565 , n32507 );
    and g13449 ( n16180 , n31965 , n20012 );
    and g13450 ( n1619 , n34683 , n14733 );
    or g13451 ( n23774 , n4753 , n13015 );
    or g13452 ( n16380 , n30553 , n16775 );
    nor g13453 ( n15644 , n10894 , n30902 );
    and g13454 ( n26833 , n598 , n1661 );
    xnor g13455 ( n23907 , n4973 , n10749 );
    xnor g13456 ( n10011 , n8938 , n4523 );
    and g13457 ( n27152 , n35857 , n28607 );
    xnor g13458 ( n27869 , n28119 , n21071 );
    or g13459 ( n17238 , n23439 , n32457 );
    or g13460 ( n17520 , n14905 , n5168 );
    or g13461 ( n26636 , n8798 , n13495 );
    or g13462 ( n30376 , n32348 , n8723 );
    xnor g13463 ( n16353 , n29956 , n35928 );
    xnor g13464 ( n22106 , n8445 , n23499 );
    or g13465 ( n17752 , n14536 , n18936 );
    not g13466 ( n15052 , n35295 );
    or g13467 ( n7870 , n33501 , n9955 );
    or g13468 ( n21797 , n23833 , n31055 );
    xnor g13469 ( n28309 , n33259 , n29196 );
    or g13470 ( n20779 , n14793 , n25394 );
    not g13471 ( n4691 , n33827 );
    xnor g13472 ( n12196 , n1447 , n30397 );
    and g13473 ( n13359 , n12568 , n5082 );
    xnor g13474 ( n2573 , n444 , n13498 );
    nor g13475 ( n34657 , n13144 , n14258 );
    xnor g13476 ( n285 , n17012 , n5326 );
    or g13477 ( n10744 , n28813 , n1630 );
    nor g13478 ( n33493 , n14208 , n6209 );
    or g13479 ( n14989 , n35927 , n22750 );
    or g13480 ( n21968 , n3645 , n20690 );
    or g13481 ( n9377 , n17794 , n11977 );
    and g13482 ( n8435 , n21793 , n30119 );
    xnor g13483 ( n31013 , n12217 , n32715 );
    and g13484 ( n10168 , n6277 , n35474 );
    buf g13485 ( n1528 , n16778 );
    xnor g13486 ( n19852 , n20518 , n9658 );
    or g13487 ( n27494 , n1656 , n14918 );
    or g13488 ( n11267 , n33673 , n27947 );
    and g13489 ( n5296 , n31188 , n6196 );
    or g13490 ( n368 , n34226 , n18152 );
    or g13491 ( n26691 , n21205 , n25594 );
    or g13492 ( n23398 , n27599 , n28866 );
    and g13493 ( n29829 , n32237 , n16681 );
    xnor g13494 ( n16237 , n24737 , n10082 );
    not g13495 ( n15738 , n24247 );
    or g13496 ( n29526 , n34132 , n2479 );
    and g13497 ( n27322 , n22775 , n33650 );
    xnor g13498 ( n2818 , n4805 , n19310 );
    or g13499 ( n35653 , n17568 , n31133 );
    xnor g13500 ( n33070 , n1083 , n5067 );
    or g13501 ( n1128 , n19551 , n34527 );
    xnor g13502 ( n15578 , n2948 , n35541 );
    and g13503 ( n6394 , n9040 , n18560 );
    nor g13504 ( n8555 , n3848 , n5601 );
    and g13505 ( n5566 , n1058 , n6444 );
    and g13506 ( n11952 , n22984 , n16869 );
    xnor g13507 ( n23758 , n16771 , n16444 );
    and g13508 ( n34016 , n11677 , n8670 );
    or g13509 ( n24986 , n4878 , n2225 );
    and g13510 ( n12640 , n19662 , n26370 );
    xnor g13511 ( n23721 , n35392 , n4960 );
    xnor g13512 ( n29979 , n6469 , n5335 );
    nor g13513 ( n25963 , n18259 , n27057 );
    xnor g13514 ( n28902 , n31481 , n32857 );
    or g13515 ( n34951 , n35911 , n4172 );
    or g13516 ( n26063 , n24954 , n867 );
    and g13517 ( n19631 , n19383 , n32007 );
    or g13518 ( n34325 , n15886 , n2148 );
    or g13519 ( n18579 , n4281 , n29853 );
    or g13520 ( n5913 , n11713 , n24489 );
    xnor g13521 ( n19191 , n12334 , n29839 );
    or g13522 ( n24 , n12401 , n11360 );
    not g13523 ( n12275 , n3239 );
    and g13524 ( n25276 , n7642 , n16504 );
    or g13525 ( n32142 , n17831 , n6950 );
    xnor g13526 ( n29360 , n29060 , n2563 );
    xnor g13527 ( n12920 , n7916 , n8432 );
    or g13528 ( n19660 , n9235 , n10762 );
    xnor g13529 ( n29456 , n20044 , n4962 );
    nor g13530 ( n8779 , n23485 , n31411 );
    not g13531 ( n19154 , n31799 );
    and g13532 ( n30896 , n25802 , n15594 );
    or g13533 ( n12605 , n691 , n6229 );
    and g13534 ( n15658 , n12343 , n15082 );
    or g13535 ( n26872 , n23034 , n3893 );
    or g13536 ( n31524 , n27226 , n21227 );
    and g13537 ( n25500 , n33141 , n31993 );
    and g13538 ( n1549 , n32015 , n5491 );
    not g13539 ( n4438 , n32922 );
    not g13540 ( n12222 , n16620 );
    and g13541 ( n12827 , n30413 , n18430 );
    not g13542 ( n4899 , n22200 );
    xnor g13543 ( n10764 , n17261 , n4421 );
    or g13544 ( n15802 , n31215 , n19456 );
    and g13545 ( n18947 , n1737 , n35963 );
    nor g13546 ( n8275 , n32095 , n9409 );
    nor g13547 ( n24556 , n3317 , n19600 );
    or g13548 ( n23555 , n9789 , n27849 );
    not g13549 ( n11389 , n14756 );
    not g13550 ( n35618 , n9975 );
    not g13551 ( n18354 , n8901 );
    or g13552 ( n29142 , n30313 , n17962 );
    and g13553 ( n8910 , n11657 , n10198 );
    or g13554 ( n2372 , n22829 , n15742 );
    or g13555 ( n7185 , n3533 , n585 );
    xnor g13556 ( n20688 , n34414 , n27291 );
    xnor g13557 ( n26783 , n8932 , n16922 );
    and g13558 ( n19910 , n7656 , n33770 );
    or g13559 ( n1077 , n19152 , n32676 );
    not g13560 ( n20567 , n26947 );
    not g13561 ( n7392 , n12698 );
    not g13562 ( n2484 , n27111 );
    not g13563 ( n26815 , n19771 );
    xnor g13564 ( n16092 , n15429 , n25402 );
    or g13565 ( n17456 , n4878 , n7779 );
    xnor g13566 ( n11259 , n31819 , n35927 );
    or g13567 ( n26766 , n12809 , n31773 );
    not g13568 ( n30364 , n2495 );
    or g13569 ( n33004 , n17509 , n34765 );
    xnor g13570 ( n31469 , n18456 , n924 );
    and g13571 ( n5026 , n20808 , n20704 );
    or g13572 ( n7953 , n19414 , n22961 );
    or g13573 ( n3151 , n9884 , n1414 );
    and g13574 ( n27251 , n2430 , n25905 );
    xnor g13575 ( n4268 , n11671 , n4960 );
    or g13576 ( n32901 , n32164 , n8203 );
    or g13577 ( n20702 , n35927 , n12482 );
    xnor g13578 ( n11068 , n29068 , n33403 );
    and g13579 ( n19951 , n26616 , n33763 );
    and g13580 ( n3651 , n2640 , n21749 );
    or g13581 ( n22325 , n34612 , n9022 );
    and g13582 ( n21978 , n21206 , n32459 );
    not g13583 ( n24751 , n670 );
    xnor g13584 ( n11706 , n33090 , n12203 );
    xnor g13585 ( n30587 , n32250 , n4288 );
    and g13586 ( n18075 , n35309 , n3804 );
    xnor g13587 ( n8217 , n10786 , n4129 );
    and g13588 ( n4369 , n7402 , n15908 );
    xnor g13589 ( n33166 , n35521 , n25602 );
    or g13590 ( n7206 , n9793 , n2047 );
    or g13591 ( n15031 , n28647 , n33435 );
    nor g13592 ( n13516 , n180 , n34218 );
    or g13593 ( n16504 , n11455 , n23494 );
    xnor g13594 ( n18001 , n35057 , n3222 );
    or g13595 ( n16624 , n8893 , n19732 );
    and g13596 ( n23067 , n26711 , n1030 );
    xnor g13597 ( n5394 , n19720 , n4288 );
    xnor g13598 ( n28945 , n27021 , n29839 );
    and g13599 ( n29139 , n29737 , n15561 );
    buf g13600 ( n4081 , n28438 );
    not g13601 ( n34991 , n11539 );
    and g13602 ( n13509 , n25027 , n32849 );
    or g13603 ( n6036 , n24371 , n19875 );
    nor g13604 ( n32052 , n2522 , n15496 );
    or g13605 ( n27731 , n20132 , n12996 );
    and g13606 ( n16794 , n35210 , n14004 );
    not g13607 ( n7648 , n7588 );
    or g13608 ( n17179 , n27393 , n24454 );
    or g13609 ( n18647 , n15282 , n15805 );
    or g13610 ( n10977 , n9862 , n8366 );
    and g13611 ( n30177 , n4040 , n31878 );
    or g13612 ( n15749 , n610 , n949 );
    nor g13613 ( n16941 , n9793 , n24721 );
    or g13614 ( n5718 , n18670 , n28837 );
    or g13615 ( n30694 , n31799 , n2503 );
    xnor g13616 ( n33487 , n24194 , n31289 );
    or g13617 ( n31327 , n7868 , n1474 );
    or g13618 ( n598 , n20829 , n25255 );
    or g13619 ( n30595 , n30470 , n4172 );
    xnor g13620 ( n29389 , n15841 , n31799 );
    nor g13621 ( n10386 , n21737 , n20762 );
    nor g13622 ( n30067 , n4960 , n22668 );
    or g13623 ( n33688 , n16487 , n9030 );
    or g13624 ( n34164 , n8533 , n29823 );
    or g13625 ( n12318 , n15780 , n19863 );
    or g13626 ( n5798 , n31855 , n13466 );
    and g13627 ( n33569 , n343 , n1188 );
    or g13628 ( n6118 , n27692 , n18705 );
    or g13629 ( n1270 , n23604 , n35667 );
    and g13630 ( n13457 , n14093 , n15530 );
    xnor g13631 ( n3193 , n9360 , n4288 );
    xnor g13632 ( n18757 , n2644 , n8288 );
    not g13633 ( n30432 , n23604 );
    or g13634 ( n8457 , n27226 , n18955 );
    xnor g13635 ( n2892 , n31038 , n27291 );
    or g13636 ( n14606 , n4960 , n30173 );
    or g13637 ( n19384 , n5335 , n28827 );
    and g13638 ( n8007 , n30908 , n19948 );
    or g13639 ( n5266 , n33879 , n628 );
    or g13640 ( n27830 , n9500 , n12950 );
    and g13641 ( n33968 , n27282 , n28793 );
    and g13642 ( n33400 , n16364 , n9557 );
    or g13643 ( n27312 , n24371 , n3837 );
    xnor g13644 ( n20302 , n468 , n19997 );
    or g13645 ( n1141 , n29839 , n18734 );
    not g13646 ( n1452 , n28172 );
    and g13647 ( n1093 , n17900 , n30041 );
    nor g13648 ( n12344 , n10967 , n21956 );
    and g13649 ( n7857 , n19764 , n32809 );
    or g13650 ( n6096 , n32911 , n4254 );
    and g13651 ( n30224 , n10077 , n2542 );
    or g13652 ( n2978 , n4379 , n2712 );
    not g13653 ( n4029 , n9793 );
    or g13654 ( n10715 , n2096 , n11447 );
    not g13655 ( n33244 , n33013 );
    xnor g13656 ( n35687 , n31781 , n19551 );
    and g13657 ( n10611 , n35277 , n11369 );
    xnor g13658 ( n25627 , n27195 , n31799 );
    and g13659 ( n6643 , n2139 , n1107 );
    xnor g13660 ( n13907 , n12048 , n10340 );
    and g13661 ( n33940 , n26104 , n26331 );
    and g13662 ( n24486 , n31463 , n4754 );
    buf g13663 ( n16797 , n6075 );
    and g13664 ( n22066 , n27439 , n30002 );
    not g13665 ( n21081 , n16413 );
    xnor g13666 ( n32390 , n13089 , n33674 );
    xnor g13667 ( n21038 , n15650 , n21007 );
    and g13668 ( n30389 , n28000 , n28529 );
    and g13669 ( n19261 , n25538 , n13334 );
    xnor g13670 ( n7683 , n7419 , n1459 );
    and g13671 ( n21084 , n35982 , n29708 );
    xnor g13672 ( n18123 , n7078 , n21824 );
    xnor g13673 ( n9249 , n13566 , n25887 );
    nor g13674 ( n18491 , n30742 , n762 );
    xnor g13675 ( n2913 , n7809 , n17183 );
    or g13676 ( n11212 , n26611 , n7516 );
    and g13677 ( n12601 , n8463 , n14838 );
    or g13678 ( n18863 , n26677 , n9108 );
    or g13679 ( n6620 , n26447 , n26737 );
    or g13680 ( n2392 , n33483 , n18949 );
    or g13681 ( n1005 , n21817 , n11800 );
    not g13682 ( n5413 , n34027 );
    and g13683 ( n21192 , n4851 , n16043 );
    or g13684 ( n18281 , n12407 , n28222 );
    or g13685 ( n33865 , n30742 , n31190 );
    xnor g13686 ( n20437 , n19085 , n25322 );
    or g13687 ( n32904 , n5627 , n10634 );
    or g13688 ( n16766 , n1088 , n32425 );
    xnor g13689 ( n28016 , n32515 , n11587 );
    or g13690 ( n6778 , n8930 , n36021 );
    and g13691 ( n29445 , n24459 , n16134 );
    not g13692 ( n3716 , n7726 );
    xnor g13693 ( n29420 , n21601 , n593 );
    xnor g13694 ( n12375 , n8147 , n16905 );
    not g13695 ( n14979 , n16620 );
    or g13696 ( n16454 , n33011 , n28240 );
    xnor g13697 ( n14740 , n23435 , n19551 );
    nor g13698 ( n25964 , n8431 , n35677 );
    xnor g13699 ( n1045 , n5884 , n4960 );
    or g13700 ( n1431 , n30059 , n2005 );
    or g13701 ( n31136 , n19990 , n9730 );
    nor g13702 ( n8981 , n25375 , n2479 );
    or g13703 ( n23779 , n23604 , n11727 );
    and g13704 ( n31675 , n20221 , n12800 );
    not g13705 ( n10689 , n33275 );
    xnor g13706 ( n24732 , n29121 , n7565 );
    or g13707 ( n26711 , n1410 , n30519 );
    nor g13708 ( n24208 , n18892 , n17895 );
    xnor g13709 ( n24542 , n18561 , n3241 );
    or g13710 ( n16231 , n30538 , n15496 );
    and g13711 ( n32559 , n17710 , n34148 );
    nor g13712 ( n10628 , n24371 , n22115 );
    not g13713 ( n879 , n22980 );
    or g13714 ( n17975 , n22942 , n35748 );
    or g13715 ( n33699 , n16821 , n18264 );
    or g13716 ( n27842 , n32883 , n30708 );
    or g13717 ( n9189 , n9789 , n21532 );
    buf g13718 ( n18811 , n21579 );
    or g13719 ( n26082 , n14456 , n13307 );
    xor g13720 ( n9502 , n2615 , n13308 );
    nor g13721 ( n3043 , n10894 , n1706 );
    and g13722 ( n19814 , n17514 , n30007 );
    or g13723 ( n19388 , n10163 , n35692 );
    and g13724 ( n30697 , n5966 , n13202 );
    or g13725 ( n27901 , n16164 , n23504 );
    xnor g13726 ( n35974 , n32642 , n30250 );
    or g13727 ( n8989 , n26472 , n10400 );
    not g13728 ( n17652 , n22980 );
    and g13729 ( n32806 , n26160 , n22565 );
    and g13730 ( n3321 , n31911 , n21674 );
    or g13731 ( n30972 , n14108 , n4595 );
    xnor g13732 ( n33130 , n4017 , n29434 );
    and g13733 ( n25469 , n2223 , n14047 );
    or g13734 ( n34436 , n16922 , n9267 );
    or g13735 ( n29109 , n255 , n23626 );
    nor g13736 ( n22165 , n18963 , n2999 );
    not g13737 ( n2502 , n31073 );
    and g13738 ( n5417 , n1651 , n23304 );
    or g13739 ( n11365 , n35522 , n21579 );
    xnor g13740 ( n23996 , n26637 , n4239 );
    or g13741 ( n9219 , n10097 , n11850 );
    or g13742 ( n1468 , n7540 , n658 );
    xnor g13743 ( n611 , n20651 , n23604 );
    xnor g13744 ( n9846 , n4013 , n23604 );
    or g13745 ( n35273 , n517 , n12128 );
    xnor g13746 ( n32139 , n4957 , n22291 );
    not g13747 ( n20595 , n8366 );
    xnor g13748 ( n4032 , n18343 , n24371 );
    xnor g13749 ( n8943 , n31895 , n29640 );
    or g13750 ( n22109 , n22552 , n22783 );
    xnor g13751 ( n7751 , n31867 , n7344 );
    xnor g13752 ( n30879 , n19948 , n29117 );
    and g13753 ( n692 , n30843 , n14282 );
    xnor g13754 ( n31686 , n29139 , n29839 );
    nor g13755 ( n11081 , n23604 , n5830 );
    or g13756 ( n13264 , n27099 , n13261 );
    nor g13757 ( n13383 , n7479 , n24431 );
    xnor g13758 ( n25440 , n25367 , n17259 );
    not g13759 ( n13312 , n22980 );
    or g13760 ( n30671 , n8516 , n4175 );
    or g13761 ( n11868 , n28706 , n32071 );
    or g13762 ( n31168 , n12468 , n34532 );
    or g13763 ( n18600 , n21058 , n2939 );
    or g13764 ( n29024 , n25602 , n18039 );
    or g13765 ( n24927 , n34151 , n4175 );
    xnor g13766 ( n24380 , n1295 , n32095 );
    or g13767 ( n22724 , n782 , n1689 );
    or g13768 ( n25722 , n3949 , n28675 );
    nor g13769 ( n32389 , n24371 , n1155 );
    xnor g13770 ( n34934 , n20823 , n19643 );
    xnor g13771 ( n9962 , n25775 , n29839 );
    xnor g13772 ( n22742 , n2385 , n4246 );
    or g13773 ( n1387 , n24371 , n22614 );
    nor g13774 ( n26662 , n25021 , n1928 );
    not g13775 ( n14674 , n28625 );
    xnor g13776 ( n35284 , n5830 , n30432 );
    xnor g13777 ( n5250 , n14678 , n17226 );
    and g13778 ( n21371 , n33349 , n34465 );
    not g13779 ( n34615 , n2029 );
    or g13780 ( n7579 , n3385 , n16797 );
    not g13781 ( n29277 , n9793 );
    and g13782 ( n33931 , n29711 , n22507 );
    xnor g13783 ( n19506 , n10664 , n23643 );
    or g13784 ( n3207 , n8955 , n10804 );
    or g13785 ( n18147 , n32981 , n9915 );
    and g13786 ( n12058 , n22472 , n28016 );
    nor g13787 ( n19354 , n31799 , n14071 );
    xnor g13788 ( n7277 , n16702 , n5041 );
    or g13789 ( n26776 , n24328 , n8153 );
    and g13790 ( n20038 , n16647 , n14888 );
    not g13791 ( n20262 , n25931 );
    xnor g13792 ( n10392 , n19323 , n9933 );
    or g13793 ( n5633 , n29839 , n7828 );
    xnor g13794 ( n12739 , n8422 , n23736 );
    or g13795 ( n17236 , n17457 , n9958 );
    and g13796 ( n2330 , n12262 , n32857 );
    xnor g13797 ( n14980 , n18780 , n31289 );
    nor g13798 ( n16185 , n4962 , n18209 );
    or g13799 ( n2115 , n17701 , n24025 );
    or g13800 ( n4404 , n22291 , n2284 );
    or g13801 ( n23433 , n30018 , n14708 );
    not g13802 ( n21674 , n4288 );
    or g13803 ( n26860 , n8831 , n32324 );
    nor g13804 ( n13704 , n15464 , n25478 );
    xnor g13805 ( n12376 , n30100 , n7808 );
    or g13806 ( n15083 , n18402 , n9601 );
    xnor g13807 ( n34290 , n14737 , n31215 );
    xnor g13808 ( n26821 , n14740 , n19887 );
    and g13809 ( n32262 , n12100 , n24034 );
    xnor g13810 ( n15139 , n8037 , n8921 );
    xnor g13811 ( n24314 , n3687 , n21983 );
    buf g13812 ( n2433 , n13098 );
    xnor g13813 ( n17098 , n34443 , n32260 );
    xnor g13814 ( n29427 , n16197 , n32857 );
    nor g13815 ( n15030 , n22150 , n7105 );
    or g13816 ( n20342 , n9136 , n11312 );
    xnor g13817 ( n23929 , n29519 , n17568 );
    and g13818 ( n14179 , n11221 , n34507 );
    and g13819 ( n34967 , n2319 , n7725 );
    xnor g13820 ( n2686 , n21604 , n12516 );
    xnor g13821 ( n2133 , n34767 , n29713 );
    and g13822 ( n23308 , n3644 , n18903 );
    or g13823 ( n1202 , n3790 , n32919 );
    nor g13824 ( n16100 , n11142 , n35168 );
    or g13825 ( n21158 , n15 , n6950 );
    or g13826 ( n31695 , n10444 , n13361 );
    and g13827 ( n6915 , n9794 , n22221 );
    or g13828 ( n30030 , n29839 , n13457 );
    or g13829 ( n2123 , n25174 , n13123 );
    or g13830 ( n10733 , n4962 , n31601 );
    and g13831 ( n4711 , n14273 , n34160 );
    xnor g13832 ( n3587 , n7939 , n10683 );
    xnor g13833 ( n32011 , n12684 , n32441 );
    nor g13834 ( n31509 , n31215 , n29622 );
    and g13835 ( n18240 , n30663 , n13836 );
    xnor g13836 ( n2708 , n29146 , n12834 );
    xnor g13837 ( n2879 , n2911 , n11372 );
    xnor g13838 ( n9607 , n6991 , n15886 );
    or g13839 ( n11131 , n16620 , n18937 );
    or g13840 ( n21133 , n4962 , n8062 );
    or g13841 ( n30055 , n4962 , n30313 );
    and g13842 ( n15235 , n18023 , n22131 );
    or g13843 ( n10013 , n4878 , n20038 );
    or g13844 ( n15120 , n18038 , n7831 );
    xnor g13845 ( n14530 , n14379 , n22819 );
    or g13846 ( n34605 , n15258 , n4930 );
    xor g13847 ( n5359 , n19727 , n30962 );
    or g13848 ( n14475 , n6622 , n28324 );
    or g13849 ( n30719 , n2335 , n2104 );
    or g13850 ( n3712 , n35927 , n8609 );
    or g13851 ( n3505 , n7488 , n25786 );
    xnor g13852 ( n13911 , n438 , n7225 );
    not g13853 ( n9155 , n19551 );
    or g13854 ( n24490 , n29333 , n8090 );
    and g13855 ( n15202 , n16520 , n34256 );
    xnor g13856 ( n26985 , n13275 , n32857 );
    or g13857 ( n467 , n16580 , n290 );
    xnor g13858 ( n13042 , n26751 , n14265 );
    not g13859 ( n3059 , n31799 );
    xnor g13860 ( n28784 , n22494 , n4758 );
    or g13861 ( n7859 , n23460 , n36029 );
    xnor g13862 ( n8960 , n13548 , n23604 );
    not g13863 ( n2629 , n18481 );
    or g13864 ( n24871 , n13661 , n25592 );
    or g13865 ( n12248 , n1950 , n7197 );
    and g13866 ( n13023 , n34288 , n6545 );
    or g13867 ( n16862 , n7368 , n8585 );
    and g13868 ( n33648 , n5758 , n2754 );
    or g13869 ( n21229 , n21060 , n29953 );
    xnor g13870 ( n27948 , n13561 , n4163 );
    and g13871 ( n28665 , n31195 , n15738 );
    or g13872 ( n10439 , n19551 , n14009 );
    not g13873 ( n6763 , n22980 );
    xnor g13874 ( n28924 , n19170 , n16922 );
    or g13875 ( n13442 , n12189 , n19786 );
    and g13876 ( n20387 , n4509 , n82 );
    xor g13877 ( n17158 , n14394 , n13350 );
    or g13878 ( n9133 , n6820 , n32329 );
    xnor g13879 ( n20494 , n12374 , n21851 );
    xnor g13880 ( n21523 , n25699 , n7540 );
    not g13881 ( n20807 , n6541 );
    or g13882 ( n30901 , n31247 , n30925 );
    xnor g13883 ( n1109 , n7336 , n17879 );
    xnor g13884 ( n12911 , n28114 , n3205 );
    or g13885 ( n2514 , n29786 , n11987 );
    or g13886 ( n33687 , n4960 , n15878 );
    or g13887 ( n18872 , n14350 , n16457 );
    or g13888 ( n9674 , n20643 , n33476 );
    xnor g13889 ( n10579 , n12621 , n30742 );
    and g13890 ( n16154 , n19857 , n32494 );
    and g13891 ( n7601 , n19318 , n4106 );
    or g13892 ( n31207 , n18802 , n28574 );
    and g13893 ( n15733 , n4237 , n2967 );
    and g13894 ( n25295 , n31868 , n17803 );
    or g13895 ( n31456 , n18020 , n28668 );
    xnor g13896 ( n16243 , n396 , n4878 );
    or g13897 ( n18177 , n8556 , n24479 );
    xnor g13898 ( n3607 , n13268 , n18047 );
    or g13899 ( n25280 , n12104 , n17612 );
    xnor g13900 ( n26631 , n30531 , n25866 );
    xnor g13901 ( n6551 , n11702 , n7540 );
    or g13902 ( n18331 , n31559 , n17016 );
    xnor g13903 ( n535 , n18719 , n26179 );
    xnor g13904 ( n21865 , n11406 , n21189 );
    or g13905 ( n9469 , n18745 , n24851 );
    or g13906 ( n1039 , n3371 , n3738 );
    xnor g13907 ( n4733 , n5081 , n23024 );
    xnor g13908 ( n16591 , n25664 , n30742 );
    and g13909 ( n31198 , n30827 , n6108 );
    or g13910 ( n12994 , n7197 , n15383 );
    or g13911 ( n9871 , n3448 , n3736 );
    or g13912 ( n8246 , n24533 , n12913 );
    and g13913 ( n17307 , n28763 , n20167 );
    nor g13914 ( n16734 , n12137 , n8041 );
    or g13915 ( n9395 , n34553 , n4557 );
    xnor g13916 ( n5788 , n22412 , n28288 );
    or g13917 ( n8900 , n2167 , n12332 );
    or g13918 ( n28569 , n3054 , n5779 );
    xnor g13919 ( n32021 , n26926 , n27300 );
    not g13920 ( n17115 , n1950 );
    and g13921 ( n8775 , n21158 , n8289 );
    or g13922 ( n15730 , n9792 , n23122 );
    xnor g13923 ( n8484 , n12732 , n13302 );
    or g13924 ( n15374 , n10408 , n10140 );
    not g13925 ( n7615 , n4494 );
    or g13926 ( n35655 , n2639 , n15256 );
    or g13927 ( n20898 , n16989 , n17233 );
    and g13928 ( n16261 , n21295 , n8758 );
    or g13929 ( n13881 , n34709 , n21078 );
    or g13930 ( n5002 , n9789 , n31955 );
    nor g13931 ( n35930 , n9789 , n28855 );
    xnor g13932 ( n16031 , n23970 , n23593 );
    xnor g13933 ( n19608 , n24956 , n16854 );
    or g13934 ( n23695 , n739 , n15145 );
    and g13935 ( n23544 , n4020 , n23771 );
    xnor g13936 ( n14023 , n24721 , n752 );
    or g13937 ( n32646 , n17000 , n17256 );
    buf g13938 ( n4254 , n6609 );
    or g13939 ( n21770 , n7173 , n3437 );
    and g13940 ( n6677 , n23948 , n29734 );
    xnor g13941 ( n13347 , n21243 , n2549 );
    or g13942 ( n17106 , n23305 , n34234 );
    or g13943 ( n31445 , n943 , n9030 );
    or g13944 ( n7330 , n21510 , n11712 );
    and g13945 ( n29896 , n31987 , n19392 );
    xnor g13946 ( n25363 , n1519 , n17173 );
    or g13947 ( n34636 , n14388 , n28837 );
    and g13948 ( n373 , n13422 , n12472 );
    xnor g13949 ( n24131 , n15531 , n14386 );
    or g13950 ( n24215 , n35927 , n19401 );
    and g13951 ( n32738 , n14377 , n31933 );
    nor g13952 ( n11763 , n3205 , n33269 );
    xnor g13953 ( n3094 , n23314 , n24559 );
    xnor g13954 ( n11653 , n6263 , n14098 );
    or g13955 ( n14069 , n26980 , n23484 );
    and g13956 ( n3560 , n23256 , n35438 );
    xnor g13957 ( n13710 , n19444 , n19551 );
    or g13958 ( n11586 , n17603 , n4254 );
    nor g13959 ( n18109 , n29713 , n11377 );
    or g13960 ( n30528 , n23604 , n3747 );
    not g13961 ( n18348 , n16980 );
    xnor g13962 ( n34346 , n27515 , n24473 );
    and g13963 ( n34763 , n29685 , n10447 );
    xnor g13964 ( n31202 , n1889 , n16162 );
    and g13965 ( n16673 , n32677 , n11788 );
    or g13966 ( n13568 , n11496 , n12159 );
    xnor g13967 ( n14364 , n6215 , n10894 );
    xnor g13968 ( n29681 , n25697 , n5445 );
    xnor g13969 ( n12489 , n18513 , n813 );
    xnor g13970 ( n24437 , n21359 , n8378 );
    or g13971 ( n28115 , n9373 , n25831 );
    nor g13972 ( n3187 , n31289 , n15398 );
    and g13973 ( n28623 , n28185 , n6918 );
    or g13974 ( n27259 , n2877 , n35359 );
    xnor g13975 ( n5416 , n1054 , n28314 );
    xnor g13976 ( n18973 , n15540 , n25524 );
    or g13977 ( n26450 , n9936 , n29393 );
    or g13978 ( n22648 , n12739 , n21210 );
    not g13979 ( n25897 , n22980 );
    nor g13980 ( n18752 , n27133 , n7175 );
    and g13981 ( n12873 , n8347 , n20686 );
    xnor g13982 ( n30965 , n23275 , n2834 );
    xnor g13983 ( n27669 , n33982 , n22576 );
    and g13984 ( n7380 , n25737 , n10597 );
    buf g13985 ( n24356 , n30033 );
    not g13986 ( n33154 , n33753 );
    or g13987 ( n24784 , n5117 , n33034 );
    and g13988 ( n9500 , n818 , n5380 );
    or g13989 ( n14011 , n30293 , n20762 );
    or g13990 ( n25748 , n3943 , n1474 );
    and g13991 ( n34248 , n26832 , n2612 );
    or g13992 ( n7449 , n33428 , n23287 );
    or g13993 ( n929 , n31840 , n28467 );
    or g13994 ( n9456 , n15962 , n23187 );
    or g13995 ( n18078 , n334 , n3703 );
    and g13996 ( n8997 , n31179 , n28537 );
    or g13997 ( n29340 , n34268 , n18841 );
    and g13998 ( n8928 , n20270 , n24709 );
    xnor g13999 ( n5964 , n15038 , n7778 );
    or g14000 ( n7246 , n9658 , n23213 );
    or g14001 ( n1189 , n11091 , n19421 );
    and g14002 ( n31601 , n8897 , n26700 );
    xnor g14003 ( n28441 , n990 , n3708 );
    or g14004 ( n8679 , n7793 , n16457 );
    and g14005 ( n3812 , n16273 , n5848 );
    xnor g14006 ( n2697 , n5872 , n5223 );
    and g14007 ( n32197 , n2559 , n33865 );
    or g14008 ( n15103 , n9510 , n12674 );
    or g14009 ( n25822 , n35028 , n34537 );
    or g14010 ( n24473 , n19345 , n19555 );
    xnor g14011 ( n20071 , n17575 , n16922 );
    or g14012 ( n15328 , n1983 , n17354 );
    or g14013 ( n12871 , n20803 , n4078 );
    or g14014 ( n8475 , n11465 , n34862 );
    and g14015 ( n21452 , n4859 , n6280 );
    xnor g14016 ( n34795 , n1948 , n16922 );
    or g14017 ( n35622 , n7324 , n21055 );
    not g14018 ( n13533 , n15036 );
    not g14019 ( n7271 , n3480 );
    or g14020 ( n21767 , n35680 , n4868 );
    xnor g14021 ( n35411 , n33027 , n17751 );
    nor g14022 ( n21235 , n9789 , n17794 );
    not g14023 ( n6263 , n18379 );
    or g14024 ( n10204 , n24064 , n35402 );
    buf g14025 ( n32379 , n19834 );
    or g14026 ( n28338 , n15230 , n25306 );
    or g14027 ( n24402 , n120 , n10867 );
    xnor g14028 ( n26799 , n22645 , n27016 );
    or g14029 ( n16917 , n12727 , n2384 );
    not g14030 ( n19448 , n26112 );
    and g14031 ( n30173 , n25494 , n33608 );
    and g14032 ( n17301 , n35135 , n9876 );
    nor g14033 ( n12380 , n11455 , n23455 );
    or g14034 ( n8087 , n19779 , n4090 );
    not g14035 ( n3276 , n1326 );
    and g14036 ( n28716 , n15010 , n3102 );
    not g14037 ( n29437 , n311 );
    or g14038 ( n7323 , n17202 , n12929 );
    xnor g14039 ( n22767 , n20057 , n9278 );
    nor g14040 ( n7095 , n25174 , n10465 );
    and g14041 ( n14476 , n6088 , n29364 );
    or g14042 ( n13128 , n21330 , n26931 );
    not g14043 ( n14813 , n27538 );
    xnor g14044 ( n25519 , n31107 , n4960 );
    or g14045 ( n32132 , n9789 , n12054 );
    or g14046 ( n28037 , n4288 , n5048 );
    or g14047 ( n2966 , n13287 , n35111 );
    xnor g14048 ( n13231 , n12771 , n30395 );
    xnor g14049 ( n24687 , n25820 , n27569 );
    or g14050 ( n1919 , n11046 , n9479 );
    nor g14051 ( n7975 , n11046 , n16539 );
    and g14052 ( n35900 , n27557 , n9364 );
    xnor g14053 ( n28856 , n16708 , n3415 );
    not g14054 ( n19158 , n35927 );
    or g14055 ( n26786 , n32340 , n22417 );
    or g14056 ( n17909 , n18015 , n6459 );
    and g14057 ( n32101 , n34114 , n28569 );
    nor g14058 ( n35814 , n1096 , n34949 );
    or g14059 ( n5295 , n8770 , n33733 );
    or g14060 ( n32899 , n1948 , n13480 );
    not g14061 ( n10266 , n21146 );
    not g14062 ( n14976 , n4878 );
    or g14063 ( n1216 , n21374 , n30287 );
    nor g14064 ( n25857 , n9789 , n34268 );
    xnor g14065 ( n14673 , n15398 , n7371 );
    and g14066 ( n12172 , n14814 , n7954 );
    and g14067 ( n4131 , n11400 , n29584 );
    not g14068 ( n12296 , n5335 );
    not g14069 ( n24364 , n2540 );
    nor g14070 ( n13223 , n23942 , n24564 );
    or g14071 ( n30497 , n4876 , n16456 );
    nor g14072 ( n25179 , n2331 , n24685 );
    or g14073 ( n23160 , n21304 , n28275 );
    or g14074 ( n32880 , n23604 , n16154 );
    or g14075 ( n1587 , n21321 , n21002 );
    xnor g14076 ( n35300 , n32569 , n14612 );
    or g14077 ( n28344 , n10664 , n23643 );
    and g14078 ( n11787 , n4039 , n11476 );
    and g14079 ( n25514 , n31380 , n19958 );
    or g14080 ( n24743 , n1312 , n30204 );
    nor g14081 ( n18692 , n9290 , n4508 );
    or g14082 ( n4520 , n2534 , n7934 );
    or g14083 ( n18843 , n4962 , n10125 );
    or g14084 ( n25806 , n19874 , n31606 );
    or g14085 ( n3443 , n24038 , n9404 );
    nor g14086 ( n33483 , n17568 , n3353 );
    xnor g14087 ( n23375 , n7281 , n33826 );
    xnor g14088 ( n209 , n27070 , n30742 );
    and g14089 ( n9507 , n23733 , n24931 );
    not g14090 ( n2800 , n11046 );
    and g14091 ( n28904 , n18157 , n34915 );
    or g14092 ( n21586 , n32715 , n14575 );
    not g14093 ( n24129 , n25602 );
    xnor g14094 ( n13830 , n31503 , n32022 );
    not g14095 ( n799 , n22471 );
    not g14096 ( n17905 , n1528 );
    not g14097 ( n14311 , n26688 );
    or g14098 ( n30379 , n3287 , n11527 );
    xnor g14099 ( n22540 , n8387 , n4962 );
    or g14100 ( n24076 , n20463 , n3858 );
    and g14101 ( n26950 , n26333 , n32978 );
    nor g14102 ( n3235 , n33916 , n478 );
    not g14103 ( n10946 , n33116 );
    and g14104 ( n17990 , n24755 , n2896 );
    or g14105 ( n25409 , n19374 , n17125 );
    and g14106 ( n20982 , n5975 , n4381 );
    or g14107 ( n4168 , n23604 , n29699 );
    and g14108 ( n10324 , n31709 , n17593 );
    nor g14109 ( n6510 , n12318 , n18095 );
    and g14110 ( n11294 , n35849 , n7485 );
    or g14111 ( n32626 , n4287 , n17775 );
    nor g14112 ( n26015 , n9789 , n14873 );
    and g14113 ( n21481 , n18425 , n20142 );
    xnor g14114 ( n17040 , n13662 , n18388 );
    and g14115 ( n30808 , n4164 , n26366 );
    or g14116 ( n31409 , n2412 , n24961 );
    not g14117 ( n17256 , n8501 );
    xnor g14118 ( n19959 , n26177 , n22841 );
    or g14119 ( n2060 , n7149 , n30419 );
    and g14120 ( n28680 , n14096 , n5207 );
    buf g14121 ( n3736 , n30406 );
    and g14122 ( n22496 , n17276 , n10779 );
    and g14123 ( n1365 , n29717 , n19315 );
    or g14124 ( n12415 , n10832 , n23001 );
    and g14125 ( n31496 , n5823 , n35968 );
    not g14126 ( n12268 , n10137 );
    or g14127 ( n34420 , n10256 , n25899 );
    or g14128 ( n11863 , n17575 , n128 );
    nor g14129 ( n901 , n19762 , n6705 );
    or g14130 ( n344 , n25214 , n8163 );
    or g14131 ( n21308 , n33935 , n14659 );
    not g14132 ( n28620 , n21545 );
    or g14133 ( n27182 , n15860 , n15321 );
    nor g14134 ( n6042 , n23880 , n35429 );
    xnor g14135 ( n5283 , n6918 , n28185 );
    and g14136 ( n14350 , n29494 , n34204 );
    or g14137 ( n1031 , n17568 , n33433 );
    xnor g14138 ( n21082 , n13149 , n32715 );
    or g14139 ( n4613 , n17839 , n10499 );
    xnor g14140 ( n28809 , n21808 , n11190 );
    or g14141 ( n14022 , n7987 , n27872 );
    and g14142 ( n9113 , n34366 , n26385 );
    or g14143 ( n32210 , n7900 , n12209 );
    and g14144 ( n30670 , n25681 , n1363 );
    and g14145 ( n11157 , n19156 , n5857 );
    nor g14146 ( n27214 , n2242 , n15497 );
    or g14147 ( n10126 , n1117 , n20601 );
    or g14148 ( n28428 , n21778 , n26931 );
    nor g14149 ( n34328 , n23604 , n29133 );
    or g14150 ( n9445 , n1174 , n5868 );
    xnor g14151 ( n16 , n23581 , n5668 );
    and g14152 ( n22303 , n10245 , n24059 );
    or g14153 ( n2593 , n23393 , n32297 );
    or g14154 ( n13807 , n14709 , n34537 );
    and g14155 ( n10319 , n19134 , n7710 );
    or g14156 ( n21936 , n13592 , n23442 );
    or g14157 ( n5982 , n27869 , n18488 );
    xnor g14158 ( n19883 , n13348 , n22291 );
    xnor g14159 ( n15915 , n8052 , n12501 );
    xnor g14160 ( n10184 , n25794 , n29644 );
    or g14161 ( n21388 , n5144 , n23633 );
    nor g14162 ( n19052 , n30587 , n20458 );
    xnor g14163 ( n28766 , n32529 , n5335 );
    not g14164 ( n1225 , n19551 );
    or g14165 ( n28122 , n32857 , n32567 );
    or g14166 ( n2294 , n30559 , n2814 );
    or g14167 ( n7117 , n19551 , n28610 );
    and g14168 ( n17300 , n28271 , n17491 );
    or g14169 ( n15751 , n5888 , n14192 );
    xnor g14170 ( n34351 , n10609 , n31163 );
    and g14171 ( n26995 , n21661 , n635 );
    or g14172 ( n5196 , n21124 , n12950 );
    nor g14173 ( n10085 , n15452 , n22086 );
    or g14174 ( n2914 , n7540 , n35808 );
    not g14175 ( n266 , n30999 );
    xnor g14176 ( n8576 , n686 , n33757 );
    or g14177 ( n9653 , n7540 , n11702 );
    and g14178 ( n9065 , n13110 , n1906 );
    xor g14179 ( n1572 , n26007 , n21949 );
    or g14180 ( n33548 , n21254 , n35170 );
    nor g14181 ( n27575 , n4960 , n16365 );
    xnor g14182 ( n10555 , n21660 , n29310 );
    and g14183 ( n202 , n1831 , n23746 );
    or g14184 ( n34395 , n4550 , n24488 );
    nor g14185 ( n20180 , n844 , n914 );
    or g14186 ( n12059 , n20541 , n3352 );
    and g14187 ( n33707 , n1555 , n11078 );
    xnor g14188 ( n15289 , n9846 , n15304 );
    nor g14189 ( n17242 , n4440 , n31774 );
    xnor g14190 ( n31945 , n5009 , n16620 );
    nor g14191 ( n8714 , n16620 , n2948 );
    not g14192 ( n6018 , n25592 );
    or g14193 ( n34766 , n29651 , n5296 );
    and g14194 ( n2137 , n19377 , n17094 );
    and g14195 ( n34041 , n5922 , n24202 );
    and g14196 ( n21258 , n29721 , n34188 );
    or g14197 ( n14337 , n8131 , n27536 );
    or g14198 ( n29653 , n1591 , n13449 );
    or g14199 ( n11961 , n17164 , n32503 );
    not g14200 ( n1455 , n32814 );
    or g14201 ( n30859 , n19307 , n7726 );
    and g14202 ( n15625 , n18122 , n17546 );
    xnor g14203 ( n30345 , n11747 , n17568 );
    nor g14204 ( n2808 , n30742 , n345 );
    xnor g14205 ( n24344 , n20596 , n34025 );
    buf g14206 ( n21862 , n18682 );
    xnor g14207 ( n23253 , n26375 , n4861 );
    or g14208 ( n28161 , n30682 , n35748 );
    and g14209 ( n18143 , n17030 , n7109 );
    and g14210 ( n10915 , n23330 , n15931 );
    not g14211 ( n27124 , n1950 );
    nor g14212 ( n2586 , n15299 , n9828 );
    or g14213 ( n1989 , n2732 , n3239 );
    xnor g14214 ( n1487 , n15474 , n32584 );
    or g14215 ( n25848 , n22991 , n7892 );
    buf g14216 ( n20797 , n17224 );
    or g14217 ( n35054 , n32584 , n7220 );
    and g14218 ( n17127 , n16870 , n35380 );
    not g14219 ( n22847 , n20035 );
    xnor g14220 ( n3017 , n32187 , n26929 );
    and g14221 ( n26773 , n10209 , n31005 );
    or g14222 ( n21429 , n29742 , n15344 );
    nor g14223 ( n15088 , n6573 , n22200 );
    xnor g14224 ( n15254 , n21669 , n534 );
    xnor g14225 ( n3506 , n14225 , n10651 );
    xnor g14226 ( n23411 , n8243 , n13699 );
    or g14227 ( n28432 , n19504 , n35757 );
    not g14228 ( n16361 , n4288 );
    xnor g14229 ( n36009 , n12938 , n30742 );
    or g14230 ( n33191 , n15111 , n31595 );
    or g14231 ( n25874 , n10958 , n15805 );
    or g14232 ( n30657 , n7310 , n24489 );
    or g14233 ( n17631 , n7540 , n19568 );
    or g14234 ( n4992 , n4960 , n21533 );
    and g14235 ( n31617 , n27927 , n33609 );
    not g14236 ( n19190 , n6773 );
    or g14237 ( n28999 , n13849 , n16464 );
    xnor g14238 ( n5628 , n10371 , n31143 );
    and g14239 ( n8550 , n21507 , n15904 );
    and g14240 ( n3956 , n25291 , n579 );
    xnor g14241 ( n22188 , n409 , n18603 );
    and g14242 ( n12947 , n24097 , n1214 );
    not g14243 ( n23148 , n3101 );
    or g14244 ( n28138 , n29884 , n26989 );
    and g14245 ( n34349 , n2577 , n26310 );
    xnor g14246 ( n21721 , n4915 , n4288 );
    xnor g14247 ( n5550 , n14405 , n17568 );
    or g14248 ( n3234 , n32857 , n27824 );
    xnor g14249 ( n6364 , n29666 , n15299 );
    and g14250 ( n23173 , n10665 , n14318 );
    or g14251 ( n5883 , n29054 , n14183 );
    and g14252 ( n33146 , n28874 , n11347 );
    or g14253 ( n31015 , n21721 , n34154 );
    xnor g14254 ( n13701 , n19401 , n35927 );
    not g14255 ( n22703 , n583 );
    or g14256 ( n15435 , n31265 , n17884 );
    xnor g14257 ( n10472 , n3397 , n15278 );
    or g14258 ( n11375 , n10833 , n4554 );
    nor g14259 ( n13666 , n4962 , n33697 );
    or g14260 ( n28578 , n2510 , n32688 );
    or g14261 ( n32453 , n29246 , n3188 );
    xnor g14262 ( n3833 , n17052 , n9793 );
    or g14263 ( n26413 , n22814 , n10634 );
    xnor g14264 ( n12986 , n20183 , n15319 );
    not g14265 ( n3405 , n8531 );
    and g14266 ( n25867 , n28237 , n31458 );
    and g14267 ( n7685 , n30662 , n19785 );
    xnor g14268 ( n11907 , n12131 , n16636 );
    and g14269 ( n25911 , n3641 , n6599 );
    or g14270 ( n10022 , n21555 , n9163 );
    xnor g14271 ( n35154 , n19374 , n16922 );
    xnor g14272 ( n32908 , n22167 , n3075 );
    nor g14273 ( n30686 , n10894 , n35369 );
    or g14274 ( n10642 , n33178 , n5183 );
    and g14275 ( n4176 , n25212 , n27000 );
    or g14276 ( n33074 , n13464 , n13664 );
    and g14277 ( n5280 , n12646 , n13985 );
    and g14278 ( n15757 , n3642 , n20707 );
    or g14279 ( n11681 , n2171 , n24769 );
    xnor g14280 ( n2385 , n7546 , n22291 );
    or g14281 ( n1735 , n15272 , n25447 );
    and g14282 ( n21089 , n23899 , n6530 );
    or g14283 ( n6655 , n9658 , n6474 );
    or g14284 ( n22887 , n18719 , n26179 );
    or g14285 ( n29556 , n24677 , n12791 );
    or g14286 ( n26654 , n34152 , n3694 );
    or g14287 ( n26277 , n32322 , n25306 );
    xnor g14288 ( n12698 , n34260 , n830 );
    or g14289 ( n29688 , n15403 , n2575 );
    not g14290 ( n2224 , n17423 );
    or g14291 ( n631 , n10048 , n3577 );
    and g14292 ( n31705 , n17296 , n29914 );
    not g14293 ( n32075 , n24371 );
    or g14294 ( n29860 , n16874 , n13015 );
    xnor g14295 ( n13944 , n35719 , n28512 );
    or g14296 ( n21183 , n19984 , n18411 );
    or g14297 ( n788 , n9065 , n24710 );
    and g14298 ( n240 , n33957 , n34494 );
    nor g14299 ( n2261 , n7769 , n15566 );
    nor g14300 ( n1067 , n16395 , n12438 );
    nor g14301 ( n11643 , n30771 , n6017 );
    not g14302 ( n10867 , n6257 );
    or g14303 ( n4083 , n6717 , n13490 );
    and g14304 ( n22154 , n16010 , n1899 );
    and g14305 ( n23883 , n3232 , n27398 );
    or g14306 ( n27838 , n30962 , n930 );
    and g14307 ( n24525 , n23895 , n10589 );
    or g14308 ( n32032 , n30742 , n27444 );
    or g14309 ( n32122 , n17863 , n21042 );
    or g14310 ( n33830 , n25755 , n720 );
    or g14311 ( n32155 , n30032 , n21042 );
    xnor g14312 ( n28165 , n23654 , n1042 );
    and g14313 ( n28089 , n35709 , n747 );
    nor g14314 ( n35500 , n31215 , n1564 );
    xnor g14315 ( n8125 , n14694 , n6064 );
    or g14316 ( n14896 , n18780 , n14918 );
    xnor g14317 ( n29146 , n28342 , n3222 );
    not g14318 ( n35960 , n5529 );
    nor g14319 ( n29309 , n14339 , n14075 );
    and g14320 ( n26568 , n23197 , n35501 );
    or g14321 ( n9741 , n572 , n20817 );
    or g14322 ( n27349 , n23253 , n34727 );
    xnor g14323 ( n12238 , n12696 , n34530 );
    xnor g14324 ( n28642 , n30018 , n14708 );
    and g14325 ( n25732 , n33209 , n23156 );
    or g14326 ( n8402 , n15621 , n27574 );
    and g14327 ( n14637 , n33809 , n5099 );
    or g14328 ( n8013 , n17098 , n4175 );
    or g14329 ( n7778 , n23826 , n11237 );
    or g14330 ( n21215 , n10054 , n27663 );
    or g14331 ( n21744 , n35927 , n27655 );
    or g14332 ( n29725 , n25266 , n4081 );
    xnor g14333 ( n35384 , n35690 , n31381 );
    or g14334 ( n857 , n21509 , n19939 );
    xnor g14335 ( n8635 , n3613 , n28636 );
    or g14336 ( n10868 , n22291 , n21354 );
    not g14337 ( n16246 , n14069 );
    or g14338 ( n29937 , n16279 , n5868 );
    xnor g14339 ( n33024 , n31624 , n12516 );
    or g14340 ( n10814 , n32349 , n12259 );
    xnor g14341 ( n31324 , n5855 , n10894 );
    or g14342 ( n12641 , n23142 , n15809 );
    xnor g14343 ( n8229 , n15317 , n9658 );
    or g14344 ( n9111 , n9628 , n22147 );
    xnor g14345 ( n1094 , n1057 , n1950 );
    or g14346 ( n32072 , n12286 , n24653 );
    or g14347 ( n11778 , n22896 , n29569 );
    and g14348 ( n30701 , n31047 , n24142 );
    or g14349 ( n4292 , n16327 , n31514 );
    or g14350 ( n11196 , n3615 , n31067 );
    nor g14351 ( n31500 , n33973 , n31014 );
    and g14352 ( n1143 , n26885 , n17517 );
    or g14353 ( n4224 , n32715 , n29159 );
    xnor g14354 ( n8846 , n23993 , n11205 );
    or g14355 ( n17911 , n11859 , n20797 );
    or g14356 ( n22352 , n7233 , n20576 );
    and g14357 ( n11089 , n3145 , n15802 );
    or g14358 ( n16430 , n830 , n20636 );
    nor g14359 ( n18552 , n16620 , n7387 );
    xnor g14360 ( n33012 , n31843 , n35909 );
    xnor g14361 ( n13546 , n34050 , n23565 );
    and g14362 ( n18220 , n27184 , n15730 );
    and g14363 ( n29298 , n12789 , n6932 );
    xnor g14364 ( n2618 , n3121 , n4878 );
    or g14365 ( n12452 , n28423 , n11258 );
    and g14366 ( n5676 , n21315 , n11133 );
    xnor g14367 ( n15978 , n14712 , n4454 );
    xnor g14368 ( n25374 , n21420 , n6791 );
    xnor g14369 ( n27983 , n17784 , n8802 );
    or g14370 ( n29779 , n681 , n28064 );
    or g14371 ( n11340 , n25318 , n7417 );
    or g14372 ( n31434 , n34795 , n23847 );
    or g14373 ( n31729 , n35927 , n26386 );
    or g14374 ( n4360 , n16135 , n21699 );
    xnor g14375 ( n41 , n32792 , n25276 );
    or g14376 ( n35266 , n27226 , n4468 );
    or g14377 ( n34354 , n27226 , n12447 );
    or g14378 ( n20454 , n10555 , n9951 );
    and g14379 ( n31331 , n25180 , n24344 );
    and g14380 ( n7883 , n16120 , n29481 );
    or g14381 ( n33003 , n21451 , n7448 );
    xnor g14382 ( n10279 , n29326 , n27185 );
    xnor g14383 ( n32299 , n24245 , n19087 );
    or g14384 ( n34042 , n1982 , n20852 );
    or g14385 ( n17883 , n32294 , n317 );
    xnor g14386 ( n18375 , n15696 , n6995 );
    or g14387 ( n6697 , n9852 , n2524 );
    and g14388 ( n7703 , n18783 , n10898 );
    or g14389 ( n33233 , n36091 , n32572 );
    or g14390 ( n12504 , n27943 , n3736 );
    or g14391 ( n2002 , n11046 , n2216 );
    or g14392 ( n32815 , n16702 , n5041 );
    or g14393 ( n21326 , n13181 , n19952 );
    or g14394 ( n11374 , n11249 , n35141 );
    or g14395 ( n3292 , n2586 , n11615 );
    or g14396 ( n31335 , n12949 , n18542 );
    or g14397 ( n26767 , n34623 , n11703 );
    nor g14398 ( n34223 , n9658 , n699 );
    not g14399 ( n26105 , n11996 );
    or g14400 ( n14647 , n27721 , n6340 );
    nor g14401 ( n8196 , n8885 , n19507 );
    buf g14402 ( n25355 , n1942 );
    or g14403 ( n13668 , n29844 , n16797 );
    nor g14404 ( n1418 , n13608 , n14351 );
    and g14405 ( n22142 , n17916 , n35688 );
    and g14406 ( n10061 , n15811 , n34316 );
    xnor g14407 ( n13367 , n9523 , n26896 );
    or g14408 ( n21393 , n31112 , n21862 );
    not g14409 ( n14903 , n35938 );
    xnor g14410 ( n13740 , n28820 , n22996 );
    xnor g14411 ( n24631 , n24840 , n22291 );
    or g14412 ( n9680 , n12355 , n33683 );
    or g14413 ( n31616 , n10512 , n17181 );
    or g14414 ( n24983 , n28108 , n25625 );
    buf g14415 ( n23089 , n10316 );
    not g14416 ( n12362 , n28563 );
    and g14417 ( n35847 , n61 , n9406 );
    xnor g14418 ( n2883 , n22337 , n1970 );
    or g14419 ( n1114 , n23737 , n12996 );
    xnor g14420 ( n8190 , n29722 , n35775 );
    and g14421 ( n8292 , n16291 , n14080 );
    or g14422 ( n9716 , n17437 , n4952 );
    or g14423 ( n18310 , n9789 , n25602 );
    xnor g14424 ( n26327 , n10832 , n23001 );
    or g14425 ( n7351 , n4962 , n31413 );
    xnor g14426 ( n17798 , n34364 , n9879 );
    and g14427 ( n23900 , n32081 , n1568 );
    xnor g14428 ( n32617 , n18424 , n34248 );
    and g14429 ( n9067 , n4903 , n10880 );
    and g14430 ( n28996 , n15214 , n25682 );
    or g14431 ( n2041 , n35914 , n20797 );
    or g14432 ( n12792 , n25602 , n21404 );
    xnor g14433 ( n30775 , n11620 , n27821 );
    or g14434 ( n32862 , n24936 , n19448 );
    not g14435 ( n1465 , n16620 );
    xnor g14436 ( n30840 , n25764 , n17887 );
    xnor g14437 ( n8131 , n120 , n31289 );
    or g14438 ( n31240 , n32780 , n15497 );
    xnor g14439 ( n32219 , n12696 , n16536 );
    or g14440 ( n5261 , n10894 , n31099 );
    or g14441 ( n19185 , n5102 , n5779 );
    and g14442 ( n25605 , n30856 , n16251 );
    or g14443 ( n2319 , n29647 , n33785 );
    xnor g14444 ( n690 , n35023 , n13741 );
    and g14445 ( n33027 , n23974 , n29002 );
    or g14446 ( n24951 , n33114 , n24851 );
    and g14447 ( n753 , n3035 , n629 );
    nor g14448 ( n23908 , n23937 , n31411 );
    or g14449 ( n1499 , n472 , n6835 );
    xnor g14450 ( n26922 , n16238 , n19079 );
    and g14451 ( n25953 , n17741 , n4094 );
    and g14452 ( n10230 , n11936 , n35576 );
    and g14453 ( n479 , n10814 , n30465 );
    or g14454 ( n10682 , n21543 , n1522 );
    or g14455 ( n20241 , n52 , n25255 );
    or g14456 ( n13498 , n13598 , n2126 );
    or g14457 ( n10291 , n3470 , n21691 );
    xnor g14458 ( n9179 , n5566 , n1950 );
    or g14459 ( n11524 , n29713 , n36084 );
    or g14460 ( n16782 , n13696 , n19105 );
    and g14461 ( n12532 , n35700 , n6432 );
    or g14462 ( n1577 , n29046 , n28031 );
    or g14463 ( n25955 , n7328 , n14841 );
    and g14464 ( n5230 , n7778 , n15038 );
    or g14465 ( n32558 , n19642 , n26431 );
    or g14466 ( n28618 , n29839 , n21311 );
    or g14467 ( n17350 , n23604 , n28545 );
    xnor g14468 ( n4007 , n3021 , n29317 );
    not g14469 ( n29270 , n24947 );
    nor g14470 ( n26531 , n9789 , n23880 );
    and g14471 ( n6686 , n35053 , n23989 );
    xnor g14472 ( n12580 , n3622 , n35585 );
    xor g14473 ( n4980 , n5798 , n29786 );
    or g14474 ( n10794 , n27379 , n26752 );
    or g14475 ( n514 , n9789 , n35855 );
    or g14476 ( n32692 , n28963 , n27682 );
    and g14477 ( n14865 , n10109 , n16088 );
    buf g14478 ( n2479 , n32898 );
    and g14479 ( n33015 , n21278 , n7660 );
    buf g14480 ( n27973 , n22498 );
    or g14481 ( n22863 , n15125 , n35422 );
    and g14482 ( n27979 , n26269 , n4117 );
    or g14483 ( n22832 , n9658 , n28261 );
    or g14484 ( n17420 , n30876 , n26023 );
    nor g14485 ( n4565 , n16509 , n991 );
    and g14486 ( n24740 , n9378 , n27354 );
    nor g14487 ( n25580 , n19093 , n7448 );
    nor g14488 ( n1779 , n5120 , n6842 );
    or g14489 ( n11864 , n2751 , n9328 );
    xnor g14490 ( n23587 , n35878 , n7019 );
    and g14491 ( n27730 , n12562 , n32355 );
    and g14492 ( n25508 , n16558 , n903 );
    or g14493 ( n20481 , n19551 , n4916 );
    not g14494 ( n33785 , n6288 );
    and g14495 ( n29454 , n33748 , n21492 );
    xnor g14496 ( n32016 , n1197 , n9793 );
    or g14497 ( n26538 , n19808 , n31345 );
    xnor g14498 ( n28980 , n17621 , n22014 );
    or g14499 ( n28447 , n19973 , n16345 );
    xnor g14500 ( n3591 , n28945 , n27758 );
    xnor g14501 ( n34317 , n21924 , n6779 );
    or g14502 ( n8791 , n21389 , n1763 );
    xnor g14503 ( n8413 , n11304 , n34340 );
    xnor g14504 ( n9057 , n23235 , n29933 );
    or g14505 ( n25881 , n13454 , n22501 );
    or g14506 ( n6355 , n16167 , n14988 );
    and g14507 ( n30057 , n10257 , n10679 );
    or g14508 ( n18459 , n19603 , n25831 );
    or g14509 ( n24303 , n29713 , n32822 );
    or g14510 ( n23624 , n11692 , n24696 );
    and g14511 ( n21675 , n21226 , n30387 );
    xnor g14512 ( n18626 , n5368 , n29884 );
    or g14513 ( n13208 , n12486 , n25594 );
    and g14514 ( n1057 , n18177 , n221 );
    xnor g14515 ( n10522 , n12018 , n1060 );
    xnor g14516 ( n25113 , n10454 , n13033 );
    or g14517 ( n21221 , n19148 , n35516 );
    xnor g14518 ( n6376 , n3574 , n23165 );
    xnor g14519 ( n18501 , n29512 , n33940 );
    xnor g14520 ( n23181 , n2138 , n8538 );
    or g14521 ( n2375 , n9789 , n9883 );
    xnor g14522 ( n9173 , n1037 , n10588 );
    or g14523 ( n23692 , n35736 , n22238 );
    or g14524 ( n1727 , n3087 , n35630 );
    and g14525 ( n9993 , n31681 , n36011 );
    or g14526 ( n19187 , n4552 , n11786 );
    or g14527 ( n7935 , n31799 , n10064 );
    or g14528 ( n31005 , n13751 , n34084 );
    or g14529 ( n21963 , n35351 , n7673 );
    or g14530 ( n15554 , n35927 , n22846 );
    xnor g14531 ( n22237 , n27787 , n8680 );
    or g14532 ( n5385 , n32119 , n16855 );
    not g14533 ( n26643 , n32371 );
    xnor g14534 ( n1563 , n24744 , n4288 );
    or g14535 ( n29950 , n32857 , n11058 );
    xnor g14536 ( n18289 , n32858 , n11224 );
    xnor g14537 ( n14423 , n34974 , n35370 );
    and g14538 ( n14108 , n9787 , n22605 );
    nor g14539 ( n26251 , n13553 , n34696 );
    or g14540 ( n13853 , n20873 , n3858 );
    and g14541 ( n19107 , n1457 , n3862 );
    nor g14542 ( n26942 , n17343 , n7448 );
    or g14543 ( n18714 , n11740 , n763 );
    or g14544 ( n3915 , n29268 , n15656 );
    and g14545 ( n11164 , n17229 , n34376 );
    and g14546 ( n14718 , n15816 , n14240 );
    and g14547 ( n10504 , n25140 , n30208 );
    or g14548 ( n9107 , n17218 , n17221 );
    or g14549 ( n13828 , n34724 , n9280 );
    or g14550 ( n24028 , n24501 , n19052 );
    nor g14551 ( n17303 , n24371 , n18164 );
    not g14552 ( n27091 , n7588 );
    or g14553 ( n22904 , n7637 , n33310 );
    xnor g14554 ( n24510 , n5361 , n17990 );
    or g14555 ( n2246 , n11046 , n34708 );
    and g14556 ( n34386 , n12347 , n19204 );
    nor g14557 ( n12961 , n14412 , n8997 );
    xnor g14558 ( n35537 , n27833 , n32095 );
    or g14559 ( n25046 , n16922 , n15168 );
    or g14560 ( n22768 , n22413 , n23748 );
    not g14561 ( n9280 , n2315 );
    or g14562 ( n18812 , n14520 , n25648 );
    xnor g14563 ( n25988 , n19042 , n24371 );
    or g14564 ( n24574 , n20548 , n12092 );
    not g14565 ( n32458 , n20790 );
    not g14566 ( n20443 , n7256 );
    or g14567 ( n2243 , n16332 , n12125 );
    and g14568 ( n4364 , n10606 , n35464 );
    or g14569 ( n35376 , n30737 , n35111 );
    or g14570 ( n25823 , n2352 , n6683 );
    xnor g14571 ( n18868 , n22227 , n4878 );
    and g14572 ( n2661 , n26838 , n34753 );
    xnor g14573 ( n4134 , n33550 , n13965 );
    not g14574 ( n1799 , n26257 );
    or g14575 ( n32111 , n15886 , n13326 );
    xnor g14576 ( n6040 , n12013 , n2769 );
    or g14577 ( n34931 , n17573 , n32572 );
    or g14578 ( n35464 , n30742 , n7937 );
    and g14579 ( n1741 , n29088 , n17527 );
    or g14580 ( n19974 , n6589 , n14918 );
    or g14581 ( n34058 , n7829 , n11996 );
    or g14582 ( n8303 , n16490 , n27053 );
    or g14583 ( n27044 , n34351 , n17964 );
    xnor g14584 ( n31551 , n270 , n9852 );
    and g14585 ( n4646 , n33135 , n12290 );
    not g14586 ( n12301 , n35173 );
    not g14587 ( n27725 , n30248 );
    and g14588 ( n2393 , n16182 , n11384 );
    or g14589 ( n19865 , n20051 , n20300 );
    and g14590 ( n4184 , n20081 , n2398 );
    and g14591 ( n19979 , n34184 , n16958 );
    not g14592 ( n17087 , n4311 );
    xnor g14593 ( n17983 , n18297 , n16922 );
    xnor g14594 ( n10845 , n11034 , n31799 );
    not g14595 ( n13939 , n35927 );
    not g14596 ( n529 , n19421 );
    or g14597 ( n14318 , n26712 , n34862 );
    xnor g14598 ( n25054 , n7722 , n30344 );
    or g14599 ( n19383 , n2034 , n31622 );
    and g14600 ( n21507 , n5333 , n4493 );
    or g14601 ( n32079 , n16178 , n25019 );
    xnor g14602 ( n23653 , n11654 , n27701 );
    not g14603 ( n11934 , n2682 );
    or g14604 ( n1279 , n25249 , n14699 );
    or g14605 ( n24271 , n11190 , n12409 );
    and g14606 ( n14987 , n30355 , n16378 );
    not g14607 ( n20598 , n34521 );
    or g14608 ( n26797 , n1813 , n34342 );
    xnor g14609 ( n10456 , n2892 , n19034 );
    not g14610 ( n25909 , n7054 );
    or g14611 ( n21500 , n12482 , n2955 );
    nor g14612 ( n9593 , n4878 , n35354 );
    or g14613 ( n33842 , n32280 , n24923 );
    and g14614 ( n7195 , n1857 , n3910 );
    or g14615 ( n35138 , n4880 , n2104 );
    nor g14616 ( n24565 , n27167 , n26476 );
    and g14617 ( n21937 , n8158 , n31292 );
    or g14618 ( n76 , n35927 , n24411 );
    nor g14619 ( n4010 , n22291 , n15006 );
    xnor g14620 ( n3745 , n28923 , n26527 );
    or g14621 ( n7374 , n31559 , n5704 );
    and g14622 ( n33859 , n8515 , n28620 );
    and g14623 ( n3573 , n24383 , n34060 );
    xnor g14624 ( n26861 , n31437 , n16922 );
    xnor g14625 ( n14945 , n18192 , n9789 );
    or g14626 ( n18134 , n10944 , n10913 );
    xnor g14627 ( n18483 , n10767 , n11455 );
    nor g14628 ( n13594 , n32095 , n11246 );
    and g14629 ( n13789 , n1823 , n32145 );
    or g14630 ( n810 , n12685 , n26931 );
    and g14631 ( n512 , n6799 , n6920 );
    not g14632 ( n982 , n27226 );
    or g14633 ( n23576 , n34175 , n15060 );
    and g14634 ( n18884 , n17449 , n12116 );
    or g14635 ( n748 , n34812 , n7364 );
    or g14636 ( n5994 , n2470 , n20812 );
    xnor g14637 ( n30486 , n20633 , n4522 );
    or g14638 ( n9096 , n34064 , n7353 );
    or g14639 ( n2486 , n34969 , n1435 );
    or g14640 ( n30350 , n34705 , n20181 );
    xnor g14641 ( n29165 , n31336 , n4029 );
    or g14642 ( n24197 , n32331 , n27903 );
    xnor g14643 ( n23630 , n1027 , n30602 );
    or g14644 ( n24513 , n27196 , n31261 );
    or g14645 ( n2737 , n9789 , n10320 );
    xnor g14646 ( n30833 , n19568 , n7540 );
    not g14647 ( n27872 , n25648 );
    or g14648 ( n13423 , n13376 , n14409 );
    and g14649 ( n20266 , n7958 , n10439 );
    and g14650 ( n12560 , n10787 , n14673 );
    or g14651 ( n16425 , n15464 , n26128 );
    or g14652 ( n907 , n20126 , n20308 );
    and g14653 ( n31946 , n18337 , n16883 );
    and g14654 ( n16097 , n868 , n32765 );
    xnor g14655 ( n34839 , n32492 , n34214 );
    nor g14656 ( n22195 , n3600 , n34391 );
    xnor g14657 ( n369 , n13578 , n20822 );
    and g14658 ( n29769 , n6964 , n28883 );
    and g14659 ( n8294 , n23302 , n12059 );
    xnor g14660 ( n25378 , n30630 , n26924 );
    and g14661 ( n17169 , n26583 , n22585 );
    xnor g14662 ( n3081 , n10547 , n15008 );
    not g14663 ( n12285 , n2419 );
    or g14664 ( n21020 , n30759 , n15496 );
    or g14665 ( n2558 , n11046 , n16738 );
    or g14666 ( n32949 , n29515 , n4318 );
    or g14667 ( n33775 , n247 , n23187 );
    xor g14668 ( n1566 , n4275 , n4913 );
    xnor g14669 ( n15413 , n20192 , n20187 );
    and g14670 ( n1034 , n20401 , n4693 );
    or g14671 ( n24001 , n7137 , n31627 );
    and g14672 ( n1378 , n8578 , n33824 );
    and g14673 ( n1088 , n27344 , n32763 );
    xnor g14674 ( n3788 , n28835 , n31289 );
    xnor g14675 ( n12338 , n19741 , n11046 );
    xnor g14676 ( n2154 , n580 , n12371 );
    not g14677 ( n16435 , n25765 );
    or g14678 ( n3089 , n7540 , n12354 );
    and g14679 ( n3518 , n21157 , n33814 );
    xnor g14680 ( n9417 , n4366 , n4288 );
    or g14681 ( n5491 , n15464 , n13464 );
    and g14682 ( n1629 , n18304 , n4708 );
    or g14683 ( n7879 , n2226 , n24781 );
    xnor g14684 ( n27168 , n25531 , n8840 );
    and g14685 ( n20836 , n2901 , n25925 );
    or g14686 ( n24523 , n22999 , n34075 );
    or g14687 ( n3748 , n4527 , n2981 );
    or g14688 ( n25703 , n19077 , n23377 );
    nor g14689 ( n19043 , n32095 , n24530 );
    xnor g14690 ( n23954 , n20960 , n4919 );
    or g14691 ( n14352 , n27196 , n33470 );
    or g14692 ( n2359 , n35927 , n26129 );
    xnor g14693 ( n7018 , n18063 , n3205 );
    xnor g14694 ( n8634 , n27811 , n24371 );
    or g14695 ( n29673 , n31799 , n30062 );
    or g14696 ( n29608 , n3652 , n1642 );
    or g14697 ( n22884 , n9658 , n10855 );
    or g14698 ( n15974 , n20095 , n2479 );
    or g14699 ( n29343 , n6854 , n6553 );
    and g14700 ( n19752 , n20442 , n9783 );
    and g14701 ( n33701 , n31029 , n9198 );
    or g14702 ( n11941 , n24814 , n139 );
    xnor g14703 ( n9625 , n11432 , n6725 );
    and g14704 ( n6388 , n14650 , n12755 );
    or g14705 ( n7092 , n29586 , n9551 );
    and g14706 ( n26989 , n31669 , n18324 );
    or g14707 ( n13534 , n21562 , n17233 );
    xnor g14708 ( n7001 , n11193 , n32095 );
    or g14709 ( n21898 , n19551 , n19469 );
    and g14710 ( n33911 , n11032 , n33231 );
    nor g14711 ( n34509 , n24371 , n33198 );
    and g14712 ( n16038 , n20351 , n35243 );
    or g14713 ( n16182 , n3571 , n10289 );
    xnor g14714 ( n17117 , n12696 , n8784 );
    xnor g14715 ( n6935 , n1811 , n6529 );
    and g14716 ( n19284 , n28531 , n33579 );
    and g14717 ( n2111 , n14406 , n20927 );
    and g14718 ( n3977 , n2273 , n599 );
    or g14719 ( n35677 , n7404 , n17776 );
    and g14720 ( n8300 , n855 , n30078 );
    and g14721 ( n4180 , n2142 , n25200 );
    or g14722 ( n22523 , n23864 , n27053 );
    nor g14723 ( n5967 , n4324 , n3754 );
    or g14724 ( n31480 , n16197 , n13900 );
    xnor g14725 ( n2685 , n17557 , n12136 );
    or g14726 ( n18907 , n4288 , n23701 );
    or g14727 ( n26771 , n16865 , n23323 );
    or g14728 ( n10178 , n31215 , n15678 );
    or g14729 ( n21592 , n7557 , n9257 );
    or g14730 ( n23903 , n18718 , n15538 );
    xnor g14731 ( n27290 , n29918 , n10331 );
    or g14732 ( n4200 , n3265 , n3634 );
    and g14733 ( n78 , n8130 , n18025 );
    and g14734 ( n19821 , n4943 , n28583 );
    xnor g14735 ( n25745 , n26326 , n22562 );
    xnor g14736 ( n1687 , n29274 , n14242 );
    and g14737 ( n28322 , n9427 , n29224 );
    or g14738 ( n27315 , n7455 , n4172 );
    or g14739 ( n7732 , n24509 , n1402 );
    nor g14740 ( n27003 , n27534 , n31411 );
    or g14741 ( n25868 , n5231 , n19105 );
    or g14742 ( n1470 , n8535 , n16345 );
    nor g14743 ( n11938 , n28285 , n29643 );
    or g14744 ( n33790 , n19829 , n2712 );
    not g14745 ( n34009 , n21618 );
    xnor g14746 ( n22559 , n3812 , n10275 );
    or g14747 ( n12322 , n16154 , n22501 );
    or g14748 ( n3441 , n11487 , n32329 );
    or g14749 ( n16408 , n4962 , n28361 );
    or g14750 ( n5769 , n2276 , n33310 );
    not g14751 ( n24249 , n23179 );
    or g14752 ( n24989 , n477 , n23090 );
    and g14753 ( n16809 , n34548 , n10780 );
    and g14754 ( n20689 , n27883 , n29943 );
    xnor g14755 ( n21618 , n10454 , n10411 );
    not g14756 ( n32180 , n28086 );
    or g14757 ( n13164 , n7998 , n6683 );
    and g14758 ( n9565 , n28183 , n15087 );
    and g14759 ( n11727 , n33624 , n24471 );
    or g14760 ( n17444 , n31215 , n32694 );
    or g14761 ( n14041 , n4720 , n20266 );
    xnor g14762 ( n8743 , n32168 , n15774 );
    not g14763 ( n5519 , n8953 );
    or g14764 ( n3436 , n20611 , n27973 );
    xnor g14765 ( n827 , n16966 , n18406 );
    or g14766 ( n1667 , n34045 , n5252 );
    and g14767 ( n17118 , n17185 , n22935 );
    nor g14768 ( n9985 , n1950 , n16528 );
    xnor g14769 ( n2304 , n18073 , n25776 );
    or g14770 ( n11037 , n9267 , n18255 );
    nor g14771 ( n31840 , n1950 , n22844 );
    or g14772 ( n4689 , n32857 , n4975 );
    or g14773 ( n6614 , n20818 , n20547 );
    and g14774 ( n26246 , n35361 , n11624 );
    nor g14775 ( n44 , n15095 , n18986 );
    or g14776 ( n7724 , n4102 , n18931 );
    xnor g14777 ( n18273 , n5539 , n22951 );
    or g14778 ( n2495 , n9956 , n25179 );
    and g14779 ( n33947 , n15646 , n16999 );
    and g14780 ( n22780 , n9274 , n30618 );
    not g14781 ( n12126 , n14267 );
    or g14782 ( n14539 , n9789 , n5417 );
    xnor g14783 ( n8304 , n9738 , n18938 );
    or g14784 ( n24135 , n3639 , n24801 );
    not g14785 ( n17753 , n29153 );
    xnor g14786 ( n1707 , n21874 , n8630 );
    and g14787 ( n1516 , n6563 , n10931 );
    xnor g14788 ( n1897 , n24186 , n25546 );
    or g14789 ( n13684 , n11971 , n32808 );
    xnor g14790 ( n24865 , n29595 , n24261 );
    or g14791 ( n13804 , n6567 , n33960 );
    or g14792 ( n9974 , n8461 , n15251 );
    and g14793 ( n5609 , n33839 , n19247 );
    or g14794 ( n27991 , n27899 , n13056 );
    or g14795 ( n626 , n9793 , n23594 );
    or g14796 ( n26525 , n10894 , n2359 );
    and g14797 ( n9081 , n28232 , n20627 );
    or g14798 ( n16096 , n34186 , n24505 );
    xnor g14799 ( n23400 , n20129 , n15022 );
    or g14800 ( n12537 , n17172 , n22091 );
    or g14801 ( n8830 , n32023 , n27381 );
    xnor g14802 ( n7473 , n18681 , n584 );
    and g14803 ( n28652 , n24101 , n7924 );
    and g14804 ( n20458 , n6268 , n17610 );
    or g14805 ( n33231 , n27370 , n24259 );
    or g14806 ( n9934 , n684 , n28675 );
    not g14807 ( n26070 , n26906 );
    and g14808 ( n8498 , n11436 , n16942 );
    or g14809 ( n8733 , n12920 , n4342 );
    or g14810 ( n18239 , n19205 , n33758 );
    nor g14811 ( n15887 , n25361 , n21309 );
    or g14812 ( n14544 , n16841 , n5470 );
    xnor g14813 ( n22446 , n20729 , n7512 );
    or g14814 ( n18865 , n25911 , n2479 );
    xnor g14815 ( n16933 , n26441 , n20520 );
    and g14816 ( n7172 , n23286 , n34402 );
    and g14817 ( n15429 , n31108 , n24352 );
    or g14818 ( n21906 , n8196 , n10531 );
    xnor g14819 ( n18826 , n16857 , n5160 );
    not g14820 ( n31058 , n7929 );
    xnor g14821 ( n25082 , n33996 , n4283 );
    or g14822 ( n3678 , n21986 , n3870 );
    or g14823 ( n25714 , n24365 , n7685 );
    xnor g14824 ( n31167 , n3332 , n15459 );
    or g14825 ( n6563 , n8422 , n23736 );
    xnor g14826 ( n8836 , n28399 , n16751 );
    and g14827 ( n8686 , n13227 , n12793 );
    and g14828 ( n29010 , n23051 , n8195 );
    or g14829 ( n25942 , n27850 , n33416 );
    or g14830 ( n35222 , n8969 , n12128 );
    xnor g14831 ( n7760 , n25250 , n32843 );
    or g14832 ( n1415 , n11839 , n26246 );
    nor g14833 ( n31674 , n14927 , n10127 );
    xnor g14834 ( n30246 , n24127 , n22088 );
    and g14835 ( n3592 , n4666 , n32655 );
    or g14836 ( n27660 , n771 , n20308 );
    or g14837 ( n30409 , n3222 , n13520 );
    not g14838 ( n33441 , n15182 );
    nor g14839 ( n25507 , n21535 , n32634 );
    and g14840 ( n32229 , n14122 , n29466 );
    and g14841 ( n22194 , n19941 , n21217 );
    or g14842 ( n12240 , n29713 , n15234 );
    or g14843 ( n14355 , n28835 , n33435 );
    or g14844 ( n29793 , n22620 , n6553 );
    or g14845 ( n938 , n27046 , n25773 );
    or g14846 ( n27664 , n2093 , n14841 );
    or g14847 ( n11579 , n25753 , n9096 );
    nor g14848 ( n35119 , n14660 , n548 );
    or g14849 ( n1995 , n1383 , n10634 );
    xnor g14850 ( n30184 , n7104 , n13433 );
    or g14851 ( n34405 , n32522 , n1763 );
    and g14852 ( n5187 , n16287 , n34141 );
    or g14853 ( n19962 , n17638 , n16919 );
    or g14854 ( n35849 , n13703 , n4172 );
    xnor g14855 ( n2768 , n9952 , n7125 );
    buf g14856 ( n31773 , n35981 );
    xor g14857 ( n1979 , n34566 , n15677 );
    xnor g14858 ( n3984 , n32382 , n25602 );
    xnor g14859 ( n14400 , n6185 , n31085 );
    and g14860 ( n7423 , n24472 , n6986 );
    or g14861 ( n1777 , n11284 , n4478 );
    or g14862 ( n28124 , n31303 , n34874 );
    and g14863 ( n32414 , n19893 , n13962 );
    and g14864 ( n24944 , n31275 , n15886 );
    and g14865 ( n28160 , n8453 , n2161 );
    nor g14866 ( n33461 , n30374 , n23773 );
    or g14867 ( n34288 , n5464 , n928 );
    or g14868 ( n32661 , n3250 , n544 );
    and g14869 ( n30296 , n8807 , n30141 );
    and g14870 ( n8872 , n27087 , n35898 );
    or g14871 ( n7510 , n3205 , n1113 );
    xnor g14872 ( n15332 , n27655 , n35927 );
    or g14873 ( n25585 , n18679 , n33034 );
    and g14874 ( n27195 , n28826 , n3067 );
    and g14875 ( n31928 , n11235 , n6519 );
    or g14876 ( n28216 , n35171 , n25306 );
    or g14877 ( n18190 , n12979 , n2823 );
    or g14878 ( n7279 , n7823 , n14918 );
    or g14879 ( n33022 , n22370 , n20601 );
    and g14880 ( n1350 , n6486 , n29706 );
    or g14881 ( n33294 , n29355 , n32504 );
    or g14882 ( n3110 , n28582 , n5705 );
    or g14883 ( n3567 , n21029 , n5168 );
    xnor g14884 ( n19012 , n10918 , n32046 );
    or g14885 ( n33352 , n32715 , n27160 );
    nor g14886 ( n12541 , n1842 , n22071 );
    and g14887 ( n20 , n33572 , n15954 );
    or g14888 ( n21599 , n20941 , n16762 );
    and g14889 ( n5879 , n2105 , n33327 );
    xnor g14890 ( n33959 , n25239 , n11812 );
    or g14891 ( n34377 , n32095 , n26515 );
    xnor g14892 ( n973 , n31190 , n30742 );
    or g14893 ( n1615 , n5552 , n17337 );
    or g14894 ( n16012 , n12447 , n9675 );
    or g14895 ( n35215 , n23922 , n6089 );
    nor g14896 ( n23725 , n29713 , n28634 );
    or g14897 ( n12941 , n17179 , n25332 );
    and g14898 ( n17705 , n2537 , n12527 );
    xnor g14899 ( n10372 , n22765 , n32095 );
    xnor g14900 ( n9090 , n15842 , n10995 );
    and g14901 ( n21417 , n30093 , n7210 );
    and g14902 ( n3379 , n6891 , n1443 );
    or g14903 ( n24074 , n29713 , n32143 );
    not g14904 ( n797 , n20226 );
    xnor g14905 ( n1420 , n20076 , n31984 );
    or g14906 ( n22528 , n30742 , n8686 );
    or g14907 ( n26814 , n30415 , n34537 );
    and g14908 ( n1253 , n15337 , n35345 );
    not g14909 ( n19251 , n12237 );
    xnor g14910 ( n22442 , n3406 , n20906 );
    xnor g14911 ( n13047 , n21538 , n33964 );
    xnor g14912 ( n33370 , n24790 , n4960 );
    not g14913 ( n12001 , n3015 );
    not g14914 ( n25993 , n4323 );
    or g14915 ( n28704 , n23587 , n27963 );
    not g14916 ( n18193 , n20427 );
    xnor g14917 ( n7367 , n35447 , n26404 );
    or g14918 ( n3454 , n24542 , n9555 );
    or g14919 ( n24100 , n20971 , n23090 );
    and g14920 ( n33826 , n9587 , n16442 );
    xnor g14921 ( n29910 , n18790 , n27166 );
    or g14922 ( n26741 , n16623 , n28837 );
    not g14923 ( n24000 , n16223 );
    or g14924 ( n4067 , n35927 , n29882 );
    and g14925 ( n25740 , n31489 , n29380 );
    xnor g14926 ( n1935 , n36035 , n27291 );
    not g14927 ( n15101 , n1261 );
    or g14928 ( n32028 , n11763 , n33219 );
    xnor g14929 ( n9392 , n6275 , n25951 );
    xnor g14930 ( n13514 , n4410 , n15451 );
    xnor g14931 ( n4693 , n6439 , n35326 );
    or g14932 ( n30086 , n284 , n4595 );
    or g14933 ( n19691 , n3539 , n2946 );
    or g14934 ( n25484 , n35854 , n3685 );
    or g14935 ( n4218 , n229 , n16762 );
    or g14936 ( n13839 , n994 , n23790 );
    or g14937 ( n6238 , n4960 , n13509 );
    nor g14938 ( n25150 , n34196 , n21810 );
    nor g14939 ( n14164 , n8933 , n34063 );
    or g14940 ( n18828 , n29713 , n16288 );
    and g14941 ( n35565 , n12187 , n24504 );
    or g14942 ( n1610 , n28123 , n31549 );
    or g14943 ( n19014 , n19864 , n7553 );
    or g14944 ( n32125 , n25972 , n25941 );
    or g14945 ( n162 , n17670 , n20268 );
    and g14946 ( n7439 , n30892 , n23952 );
    xnor g14947 ( n26272 , n6247 , n24165 );
    xnor g14948 ( n27834 , n17823 , n15741 );
    and g14949 ( n28212 , n24166 , n34917 );
    and g14950 ( n12257 , n10096 , n7332 );
    not g14951 ( n2609 , n17224 );
    or g14952 ( n16434 , n22291 , n4905 );
    xnor g14953 ( n13524 , n767 , n5287 );
    and g14954 ( n19636 , n17381 , n35172 );
    or g14955 ( n27466 , n10392 , n30826 );
    and g14956 ( n9520 , n35885 , n30446 );
    or g14957 ( n8578 , n4826 , n10634 );
    nor g14958 ( n17393 , n14040 , n10867 );
    nor g14959 ( n25810 , n32836 , n27096 );
    nor g14960 ( n393 , n14317 , n11021 );
    or g14961 ( n14058 , n23764 , n27574 );
    and g14962 ( n24707 , n33592 , n32396 );
    or g14963 ( n13573 , n16922 , n24331 );
    or g14964 ( n11173 , n34029 , n17974 );
    or g14965 ( n22545 , n32477 , n17162 );
    or g14966 ( n2722 , n2808 , n24943 );
    not g14967 ( n20487 , n33387 );
    not g14968 ( n28172 , n13925 );
    and g14969 ( n31024 , n10079 , n5462 );
    xnor g14970 ( n23731 , n2762 , n4135 );
    xnor g14971 ( n20668 , n34242 , n8371 );
    or g14972 ( n1985 , n24334 , n32468 );
    or g14973 ( n18077 , n9793 , n27844 );
    or g14974 ( n31553 , n5335 , n15884 );
    or g14975 ( n15709 , n6192 , n12456 );
    and g14976 ( n35986 , n29916 , n11907 );
    and g14977 ( n21336 , n19164 , n15151 );
    xnor g14978 ( n17234 , n5110 , n33542 );
    or g14979 ( n7535 , n20069 , n26894 );
    or g14980 ( n2347 , n31559 , n31112 );
    xnor g14981 ( n34475 , n19976 , n31559 );
    or g14982 ( n4107 , n6439 , n18255 );
    or g14983 ( n19067 , n8432 , n24281 );
    or g14984 ( n35416 , n14803 , n16762 );
    or g14985 ( n32564 , n17349 , n2890 );
    not g14986 ( n15799 , n14582 );
    xnor g14987 ( n27616 , n15962 , n4288 );
    and g14988 ( n10320 , n67 , n28290 );
    and g14989 ( n31523 , n3883 , n16140 );
    or g14990 ( n14333 , n20331 , n16417 );
    or g14991 ( n12646 , n1902 , n16919 );
    or g14992 ( n7066 , n19688 , n34386 );
    or g14993 ( n974 , n26581 , n128 );
    xnor g14994 ( n24119 , n33787 , n18665 );
    not g14995 ( n16516 , n3480 );
    and g14996 ( n17899 , n19325 , n33553 );
    xnor g14997 ( n13168 , n13674 , n7540 );
    and g14998 ( n22305 , n21469 , n20484 );
    or g14999 ( n24417 , n29262 , n6459 );
    or g15000 ( n10045 , n19720 , n31606 );
    or g15001 ( n13379 , n5316 , n29156 );
    xnor g15002 ( n21512 , n7004 , n19704 );
    xnor g15003 ( n33965 , n1983 , n22291 );
    and g15004 ( n17729 , n1170 , n24144 );
    or g15005 ( n15839 , n4288 , n23387 );
    or g15006 ( n31944 , n22286 , n20033 );
    nor g15007 ( n28940 , n4355 , n15345 );
    or g15008 ( n3288 , n32857 , n27919 );
    or g15009 ( n18526 , n8845 , n11712 );
    nor g15010 ( n32777 , n29166 , n28422 );
    not g15011 ( n32961 , n11996 );
    nor g15012 ( n8420 , n5335 , n9517 );
    or g15013 ( n27147 , n20073 , n12622 );
    or g15014 ( n4329 , n11616 , n4127 );
    or g15015 ( n13953 , n29529 , n21956 );
    or g15016 ( n9977 , n12714 , n14076 );
    xnor g15017 ( n34726 , n11148 , n7913 );
    and g15018 ( n23642 , n16795 , n15808 );
    and g15019 ( n331 , n3425 , n35871 );
    or g15020 ( n4887 , n29713 , n18099 );
    buf g15021 ( n13215 , n11079 );
    xnor g15022 ( n13346 , n25425 , n4188 );
    xnor g15023 ( n15698 , n31535 , n35927 );
    or g15024 ( n17410 , n9483 , n20300 );
    xnor g15025 ( n28628 , n13689 , n11455 );
    xnor g15026 ( n7199 , n21998 , n5335 );
    not g15027 ( n34012 , n22188 );
    not g15028 ( n12468 , n35972 );
    or g15029 ( n12783 , n24953 , n1511 );
    and g15030 ( n2863 , n1545 , n10118 );
    or g15031 ( n18228 , n4893 , n24653 );
    or g15032 ( n18582 , n34091 , n29172 );
    or g15033 ( n2541 , n16 , n4203 );
    or g15034 ( n6417 , n132 , n21985 );
    or g15035 ( n352 , n22175 , n16456 );
    or g15036 ( n25758 , n4807 , n30708 );
    or g15037 ( n13895 , n30865 , n16659 );
    xnor g15038 ( n5436 , n28720 , n10894 );
    and g15039 ( n11740 , n5281 , n24070 );
    xnor g15040 ( n7411 , n30523 , n5816 );
    and g15041 ( n29310 , n18369 , n33228 );
    or g15042 ( n3329 , n10497 , n554 );
    xnor g15043 ( n5910 , n32915 , n23308 );
    nor g15044 ( n6856 , n10894 , n33897 );
    nor g15045 ( n33079 , n27291 , n35386 );
    or g15046 ( n15662 , n32095 , n27151 );
    or g15047 ( n8999 , n29837 , n23462 );
    not g15048 ( n15861 , n1655 );
    and g15049 ( n26693 , n24001 , n17679 );
    xnor g15050 ( n7504 , n25172 , n31919 );
    nor g15051 ( n3221 , n14955 , n34084 );
    or g15052 ( n33602 , n24624 , n28675 );
    or g15053 ( n23501 , n35555 , n33435 );
    not g15054 ( n740 , n9209 );
    xnor g15055 ( n7630 , n12258 , n33097 );
    or g15056 ( n24096 , n313 , n16961 );
    or g15057 ( n16162 , n26197 , n24866 );
    and g15058 ( n3540 , n1508 , n4022 );
    or g15059 ( n30413 , n4499 , n12370 );
    or g15060 ( n17960 , n24216 , n29514 );
    or g15061 ( n10837 , n28142 , n21782 );
    nor g15062 ( n13974 , n1950 , n35786 );
    or g15063 ( n21289 , n15886 , n11825 );
    nor g15064 ( n8629 , n9063 , n8934 );
    and g15065 ( n27893 , n20407 , n25047 );
    xnor g15066 ( n29082 , n19790 , n35927 );
    and g15067 ( n32828 , n31882 , n3080 );
    and g15068 ( n17151 , n28002 , n24692 );
    or g15069 ( n22908 , n32857 , n32092 );
    or g15070 ( n14292 , n31205 , n13943 );
    or g15071 ( n8220 , n13275 , n5521 );
    or g15072 ( n3938 , n33874 , n3744 );
    or g15073 ( n17057 , n18379 , n18518 );
    or g15074 ( n34933 , n18581 , n31968 );
    and g15075 ( n25658 , n17683 , n20231 );
    and g15076 ( n8319 , n20131 , n170 );
    xnor g15077 ( n4469 , n35268 , n25482 );
    or g15078 ( n18701 , n24371 , n253 );
    xnor g15079 ( n10653 , n28157 , n560 );
    or g15080 ( n34854 , n7956 , n25611 );
    and g15081 ( n854 , n20345 , n24205 );
    or g15082 ( n29119 , n6646 , n27801 );
    or g15083 ( n25573 , n1950 , n16812 );
    xnor g15084 ( n26625 , n31947 , n22017 );
    and g15085 ( n12858 , n25777 , n28110 );
    and g15086 ( n31498 , n35532 , n34640 );
    or g15087 ( n33221 , n2182 , n10942 );
    and g15088 ( n7702 , n31560 , n5148 );
    or g15089 ( n27909 , n23177 , n2117 );
    and g15090 ( n32701 , n28955 , n24393 );
    and g15091 ( n8549 , n22116 , n28469 );
    or g15092 ( n19667 , n15979 , n11428 );
    xnor g15093 ( n244 , n18125 , n23204 );
    and g15094 ( n28551 , n24527 , n5642 );
    not g15095 ( n18841 , n22241 );
    or g15096 ( n12875 , n16245 , n2448 );
    xnor g15097 ( n2949 , n4021 , n32756 );
    or g15098 ( n22310 , n34 , n5868 );
    or g15099 ( n30971 , n8756 , n34451 );
    and g15100 ( n19989 , n31015 , n4961 );
    or g15101 ( n23465 , n10060 , n17190 );
    and g15102 ( n22427 , n35405 , n15865 );
    not g15103 ( n27206 , n30961 );
    and g15104 ( n14289 , n8111 , n98 );
    and g15105 ( n4580 , n8207 , n22901 );
    or g15106 ( n2664 , n2732 , n5208 );
    or g15107 ( n10578 , n22810 , n370 );
    or g15108 ( n30202 , n20098 , n20272 );
    or g15109 ( n23229 , n1950 , n1338 );
    or g15110 ( n21137 , n12458 , n8366 );
    xnor g15111 ( n11796 , n19274 , n22386 );
    or g15112 ( n14139 , n13656 , n2664 );
    xnor g15113 ( n18597 , n26010 , n15886 );
    or g15114 ( n35647 , n27779 , n24729 );
    buf g15115 ( n2823 , n25521 );
    and g15116 ( n17932 , n2947 , n12543 );
    or g15117 ( n35526 , n21147 , n20601 );
    and g15118 ( n30680 , n29111 , n26203 );
    xnor g15119 ( n362 , n28108 , n17751 );
    xnor g15120 ( n9318 , n30026 , n26108 );
    not g15121 ( n5724 , n1942 );
    or g15122 ( n6267 , n19984 , n19983 );
    xnor g15123 ( n32622 , n17338 , n21870 );
    not g15124 ( n10499 , n20840 );
    or g15125 ( n23827 , n16674 , n17861 );
    nor g15126 ( n35550 , n10153 , n908 );
    not g15127 ( n26357 , n4265 );
    and g15128 ( n15281 , n526 , n8138 );
    and g15129 ( n14458 , n29795 , n9362 );
    xnor g15130 ( n29008 , n27031 , n23604 );
    or g15131 ( n22185 , n15299 , n31707 );
    and g15132 ( n2112 , n6261 , n9201 );
    or g15133 ( n15563 , n31799 , n22531 );
    and g15134 ( n6527 , n9801 , n22828 );
    or g15135 ( n24935 , n25234 , n128 );
    or g15136 ( n22019 , n31215 , n17305 );
    and g15137 ( n6392 , n3118 , n23294 );
    nor g15138 ( n4648 , n33224 , n19619 );
    or g15139 ( n11310 , n2876 , n32329 );
    or g15140 ( n34672 , n25608 , n9194 );
    or g15141 ( n18746 , n22317 , n21338 );
    xnor g15142 ( n7981 , n6534 , n31289 );
    or g15143 ( n10144 , n5694 , n17709 );
    not g15144 ( n27436 , n5067 );
    or g15145 ( n24041 , n4288 , n19449 );
    or g15146 ( n23821 , n35414 , n30419 );
    xnor g15147 ( n9913 , n12696 , n30716 );
    xnor g15148 ( n20803 , n6643 , n9793 );
    nor g15149 ( n24173 , n31056 , n25471 );
    and g15150 ( n17812 , n7576 , n29684 );
    nor g15151 ( n33367 , n33541 , n4712 );
    and g15152 ( n23507 , n9753 , n21968 );
    and g15153 ( n22761 , n30913 , n26026 );
    or g15154 ( n3699 , n11693 , n14197 );
    not g15155 ( n28012 , n32095 );
    and g15156 ( n6701 , n3119 , n20204 );
    or g15157 ( n7715 , n27696 , n2479 );
    and g15158 ( n20912 , n16868 , n27840 );
    or g15159 ( n17987 , n36016 , n33161 );
    and g15160 ( n32080 , n29377 , n7532 );
    or g15161 ( n570 , n11058 , n9731 );
    or g15162 ( n18347 , n4962 , n32772 );
    or g15163 ( n24055 , n14861 , n16246 );
    or g15164 ( n23762 , n32576 , n24567 );
    and g15165 ( n28357 , n5308 , n25827 );
    and g15166 ( n22086 , n13052 , n19132 );
    and g15167 ( n35262 , n8397 , n15287 );
    not g15168 ( n5215 , n29713 );
    or g15169 ( n21546 , n27777 , n12069 );
    xnor g15170 ( n11632 , n34350 , n33494 );
    or g15171 ( n5433 , n3099 , n10400 );
    not g15172 ( n7842 , n28430 );
    xnor g15173 ( n7900 , n9936 , n5335 );
    xnor g15174 ( n3525 , n25975 , n28644 );
    xnor g15175 ( n17442 , n17991 , n4960 );
    or g15176 ( n9471 , n35927 , n13956 );
    nor g15177 ( n31148 , n9736 , n35969 );
    or g15178 ( n16789 , n19752 , n4772 );
    and g15179 ( n21907 , n24273 , n19027 );
    or g15180 ( n15682 , n1732 , n10548 );
    and g15181 ( n32637 , n4228 , n7562 );
    not g15182 ( n35990 , n20834 );
    not g15183 ( n16329 , n1701 );
    nor g15184 ( n9813 , n21737 , n35609 );
    xnor g15185 ( n14975 , n35687 , n14407 );
    nor g15186 ( n28062 , n32928 , n35159 );
    or g15187 ( n19764 , n34562 , n24634 );
    and g15188 ( n18862 , n21755 , n8199 );
    nor g15189 ( n9780 , n19954 , n7187 );
    and g15190 ( n22793 , n8424 , n5438 );
    buf g15191 ( n16919 , n1528 );
    xnor g15192 ( n15132 , n35707 , n12230 );
    or g15193 ( n16826 , n7957 , n32959 );
    xnor g15194 ( n17136 , n16857 , n23854 );
    and g15195 ( n13097 , n17625 , n16743 );
    xnor g15196 ( n1992 , n9228 , n4530 );
    xnor g15197 ( n28470 , n24979 , n263 );
    or g15198 ( n11659 , n31003 , n2112 );
    and g15199 ( n32963 , n3986 , n35513 );
    or g15200 ( n3451 , n19286 , n28064 );
    not g15201 ( n28196 , n29657 );
    not g15202 ( n26676 , n25032 );
    not g15203 ( n31683 , n6257 );
    or g15204 ( n13081 , n23491 , n6159 );
    and g15205 ( n20389 , n27971 , n25483 );
    or g15206 ( n21726 , n21169 , n28675 );
    or g15207 ( n10079 , n890 , n12272 );
    nor g15208 ( n7295 , n16620 , n18795 );
    not g15209 ( n26864 , n13265 );
    nor g15210 ( n9174 , n150 , n24000 );
    not g15211 ( n946 , n16620 );
    or g15212 ( n23557 , n2693 , n35036 );
    and g15213 ( n27656 , n29712 , n6729 );
    xnor g15214 ( n17431 , n8808 , n27920 );
    or g15215 ( n9713 , n32584 , n19255 );
    and g15216 ( n14437 , n14008 , n33029 );
    xnor g15217 ( n7041 , n20389 , n17568 );
    or g15218 ( n32261 , n20668 , n25404 );
    or g15219 ( n17131 , n2215 , n12901 );
    xnor g15220 ( n15739 , n5156 , n20616 );
    or g15221 ( n15772 , n27617 , n32753 );
    or g15222 ( n12825 , n30209 , n24696 );
    not g15223 ( n7562 , n18726 );
    and g15224 ( n34251 , n5943 , n23822 );
    not g15225 ( n20631 , n20976 );
    or g15226 ( n18557 , n32095 , n33170 );
    xnor g15227 ( n26725 , n32780 , n27080 );
    and g15228 ( n3215 , n20062 , n6232 );
    or g15229 ( n32483 , n6415 , n34865 );
    or g15230 ( n35941 , n11931 , n26468 );
    or g15231 ( n36032 , n1950 , n15056 );
    or g15232 ( n24881 , n15128 , n24333 );
    and g15233 ( n32093 , n30131 , n22718 );
    or g15234 ( n25349 , n17635 , n25592 );
    or g15235 ( n6839 , n31533 , n25468 );
    buf g15236 ( n16543 , n2287 );
    and g15237 ( n16314 , n26809 , n26489 );
    or g15238 ( n16581 , n25984 , n20762 );
    xnor g15239 ( n4585 , n26407 , n31215 );
    xnor g15240 ( n5955 , n33804 , n11982 );
    or g15241 ( n33679 , n8849 , n29953 );
    buf g15242 ( n28240 , n19566 );
    or g15243 ( n6305 , n18218 , n3382 );
    nor g15244 ( n34179 , n9793 , n6439 );
    nor g15245 ( n27940 , n5287 , n12487 );
    xnor g15246 ( n26868 , n26541 , n18486 );
    xnor g15247 ( n22190 , n1855 , n8039 );
    xnor g15248 ( n21197 , n13068 , n4886 );
    not g15249 ( n2235 , n22980 );
    nor g15250 ( n25898 , n28003 , n24488 );
    and g15251 ( n5234 , n332 , n3411 );
    not g15252 ( n4514 , n16326 );
    nor g15253 ( n4723 , n3205 , n150 );
    xnor g15254 ( n4122 , n25236 , n10894 );
    or g15255 ( n31872 , n20516 , n25694 );
    xnor g15256 ( n34385 , n22347 , n5806 );
    or g15257 ( n31011 , n22373 , n14414 );
    and g15258 ( n25752 , n8728 , n8668 );
    and g15259 ( n6297 , n32553 , n17704 );
    and g15260 ( n7373 , n18489 , n3238 );
    nor g15261 ( n1708 , n16620 , n16951 );
    and g15262 ( n6825 , n29115 , n2481 );
    not g15263 ( n31755 , n596 );
    not g15264 ( n34723 , n28273 );
    or g15265 ( n2336 , n5979 , n15496 );
    not g15266 ( n23708 , n14593 );
    or g15267 ( n9954 , n22491 , n16888 );
    xnor g15268 ( n32921 , n20727 , n11455 );
    nor g15269 ( n20848 , n11046 , n29911 );
    and g15270 ( n25368 , n6203 , n6905 );
    or g15271 ( n19774 , n6474 , n18841 );
    or g15272 ( n22733 , n20887 , n35935 );
    or g15273 ( n9434 , n27430 , n18488 );
    and g15274 ( n22746 , n15786 , n3857 );
    or g15275 ( n28296 , n29488 , n1176 );
    or g15276 ( n17340 , n11190 , n23020 );
    xnor g15277 ( n2214 , n5240 , n33342 );
    not g15278 ( n16090 , n18912 );
    or g15279 ( n17927 , n29232 , n24333 );
    or g15280 ( n8944 , n17983 , n6582 );
    xnor g15281 ( n16424 , n31306 , n30867 );
    or g15282 ( n17574 , n21601 , n593 );
    or g15283 ( n28845 , n738 , n25904 );
    nor g15284 ( n7243 , n18057 , n16649 );
    xnor g15285 ( n24593 , n7968 , n12208 );
    and g15286 ( n9009 , n1211 , n7501 );
    or g15287 ( n35583 , n5880 , n27728 );
    or g15288 ( n24957 , n6294 , n15534 );
    or g15289 ( n4735 , n5218 , n31587 );
    xnor g15290 ( n17950 , n29829 , n9658 );
    or g15291 ( n22759 , n29666 , n17962 );
    or g15292 ( n30760 , n16922 , n30658 );
    xnor g15293 ( n11625 , n12886 , n5335 );
    nor g15294 ( n18156 , n35927 , n15695 );
    xnor g15295 ( n17638 , n17273 , n34794 );
    and g15296 ( n33444 , n23936 , n23865 );
    or g15297 ( n16929 , n9266 , n15812 );
    and g15298 ( n29431 , n8223 , n13915 );
    or g15299 ( n22920 , n5335 , n21978 );
    not g15300 ( n12021 , n25572 );
    or g15301 ( n11189 , n11190 , n17587 );
    or g15302 ( n24780 , n12480 , n2524 );
    and g15303 ( n1135 , n8136 , n11586 );
    and g15304 ( n32477 , n11512 , n32829 );
    or g15305 ( n22486 , n143 , n28475 );
    or g15306 ( n29285 , n34972 , n35519 );
    or g15307 ( n25947 , n7200 , n33034 );
    or g15308 ( n13327 , n25988 , n9812 );
    or g15309 ( n8415 , n13956 , n33435 );
    xnor g15310 ( n10241 , n33812 , n23604 );
    or g15311 ( n21519 , n34805 , n24585 );
    xnor g15312 ( n4085 , n35640 , n23943 );
    or g15313 ( n9462 , n12630 , n9882 );
    and g15314 ( n24442 , n6923 , n24688 );
    or g15315 ( n25659 , n28646 , n9825 );
    nor g15316 ( n18994 , n10894 , n8975 );
    or g15317 ( n35101 , n35927 , n16330 );
    or g15318 ( n26484 , n4962 , n25264 );
    xnor g15319 ( n27395 , n11744 , n22291 );
    xnor g15320 ( n25265 , n15276 , n27475 );
    xnor g15321 ( n25128 , n18718 , n5837 );
    and g15322 ( n12964 , n2485 , n9566 );
    not g15323 ( n18385 , n30822 );
    xnor g15324 ( n31972 , n31307 , n4962 );
    or g15325 ( n8681 , n1950 , n10777 );
    or g15326 ( n15455 , n21092 , n32138 );
    xnor g15327 ( n14656 , n23346 , n24371 );
    and g15328 ( n21392 , n2790 , n1640 );
    not g15329 ( n12922 , n4962 );
    nor g15330 ( n20980 , n15744 , n8835 );
    or g15331 ( n23234 , n34815 , n6024 );
    or g15332 ( n14211 , n12388 , n27774 );
    or g15333 ( n31763 , n5077 , n26951 );
    xnor g15334 ( n3867 , n23963 , n33578 );
    and g15335 ( n13036 , n25600 , n22462 );
    or g15336 ( n34808 , n24998 , n9815 );
    not g15337 ( n8002 , n13318 );
    xnor g15338 ( n26078 , n16062 , n24551 );
    and g15339 ( n14855 , n23775 , n18852 );
    nor g15340 ( n26339 , n3281 , n30646 );
    or g15341 ( n17347 , n19341 , n35935 );
    or g15342 ( n10597 , n16051 , n2798 );
    or g15343 ( n16686 , n32095 , n4301 );
    and g15344 ( n2943 , n9869 , n20744 );
    xnor g15345 ( n30232 , n16935 , n26512 );
    and g15346 ( n11415 , n6378 , n14465 );
    or g15347 ( n26349 , n20343 , n6908 );
    or g15348 ( n7891 , n11498 , n5865 );
    or g15349 ( n25756 , n25269 , n33706 );
    and g15350 ( n3942 , n28297 , n33365 );
    nor g15351 ( n16901 , n30968 , n2578 );
    xor g15352 ( n32214 , n8746 , n25097 );
    xnor g15353 ( n27638 , n22541 , n17576 );
    or g15354 ( n6219 , n31272 , n8903 );
    or g15355 ( n23978 , n10768 , n29124 );
    or g15356 ( n16596 , n1950 , n26680 );
    or g15357 ( n2023 , n5616 , n10007 );
    or g15358 ( n25284 , n26068 , n35238 );
    or g15359 ( n6869 , n16202 , n2698 );
    xnor g15360 ( n3616 , n15526 , n13792 );
    buf g15361 ( n28866 , n9051 );
    and g15362 ( n28901 , n1868 , n11319 );
    nor g15363 ( n12087 , n31289 , n5304 );
    or g15364 ( n22463 , n4758 , n34763 );
    or g15365 ( n30567 , n34784 , n35425 );
    or g15366 ( n18575 , n33697 , n34484 );
    or g15367 ( n33832 , n27819 , n3577 );
    or g15368 ( n31770 , n464 , n11197 );
    or g15369 ( n15958 , n34981 , n17673 );
    or g15370 ( n16576 , n4085 , n29872 );
    or g15371 ( n35198 , n4037 , n21673 );
    or g15372 ( n13019 , n31853 , n14452 );
    or g15373 ( n1710 , n30314 , n28351 );
    and g15374 ( n15316 , n30929 , n26644 );
    or g15375 ( n28687 , n29713 , n75 );
    xnor g15376 ( n23925 , n22390 , n15249 );
    and g15377 ( n35445 , n24690 , n7824 );
    xnor g15378 ( n25162 , n10101 , n2501 );
    or g15379 ( n15549 , n26232 , n32717 );
    xnor g15380 ( n8936 , n32418 , n4488 );
    or g15381 ( n25398 , n11083 , n20200 );
    xnor g15382 ( n2413 , n13524 , n34139 );
    and g15383 ( n34323 , n1713 , n28961 );
    xnor g15384 ( n11346 , n2619 , n23604 );
    or g15385 ( n1433 , n10221 , n14582 );
    or g15386 ( n4577 , n7327 , n14572 );
    xor g15387 ( n9833 , n16532 , n28001 );
    or g15388 ( n29832 , n10894 , n28684 );
    xnor g15389 ( n8137 , n15155 , n6381 );
    and g15390 ( n23558 , n18840 , n20075 );
    and g15391 ( n13348 , n30187 , n30895 );
    or g15392 ( n21505 , n9371 , n26292 );
    and g15393 ( n5874 , n13958 , n26501 );
    and g15394 ( n14780 , n21347 , n28053 );
    and g15395 ( n15609 , n22393 , n9733 );
    or g15396 ( n32869 , n21544 , n17413 );
    and g15397 ( n25847 , n5906 , n23592 );
    or g15398 ( n27455 , n29058 , n35935 );
    or g15399 ( n8035 , n5335 , n28073 );
    xnor g15400 ( n24945 , n28834 , n34408 );
    xnor g15401 ( n34355 , n3784 , n32395 );
    or g15402 ( n32833 , n4962 , n18612 );
    xnor g15403 ( n28272 , n14279 , n6217 );
    xor g15404 ( n10910 , n31217 , n30655 );
    xnor g15405 ( n7997 , n12925 , n32584 );
    and g15406 ( n19061 , n27093 , n14828 );
    or g15407 ( n27157 , n9793 , n27985 );
    or g15408 ( n34372 , n7878 , n4445 );
    not g15409 ( n4988 , n3793 );
    or g15410 ( n26940 , n33226 , n1311 );
    and g15411 ( n16925 , n11145 , n1547 );
    and g15412 ( n23891 , n28311 , n4987 );
    and g15413 ( n6864 , n1644 , n34961 );
    xnor g15414 ( n36080 , n21758 , n7540 );
    or g15415 ( n27578 , n13617 , n9345 );
    nor g15416 ( n4882 , n1933 , n33163 );
    or g15417 ( n14923 , n30701 , n35935 );
    or g15418 ( n23797 , n33921 , n30754 );
    and g15419 ( n32893 , n28655 , n9106 );
    not g15420 ( n8983 , n28627 );
    or g15421 ( n354 , n13207 , n35630 );
    or g15422 ( n16877 , n31272 , n16750 );
    and g15423 ( n7303 , n30012 , n3712 );
    or g15424 ( n4124 , n4178 , n34472 );
    xnor g15425 ( n18439 , n25541 , n15548 );
    and g15426 ( n10829 , n5916 , n4159 );
    xnor g15427 ( n34228 , n6115 , n32968 );
    and g15428 ( n32408 , n4236 , n21123 );
    or g15429 ( n6448 , n1950 , n15829 );
    and g15430 ( n34650 , n5272 , n4060 );
    and g15431 ( n19890 , n35595 , n25192 );
    or g15432 ( n11902 , n7519 , n11601 );
    buf g15433 ( n6017 , n5592 );
    xnor g15434 ( n21184 , n22309 , n4946 );
    or g15435 ( n34851 , n29519 , n14706 );
    not g15436 ( n7268 , n28223 );
    and g15437 ( n12164 , n23054 , n722 );
    or g15438 ( n27765 , n12455 , n34235 );
    or g15439 ( n9803 , n15187 , n18488 );
    or g15440 ( n984 , n18286 , n34575 );
    or g15441 ( n14642 , n27292 , n773 );
    or g15442 ( n2989 , n15361 , n9410 );
    and g15443 ( n35089 , n29371 , n12977 );
    and g15444 ( n6907 , n15898 , n8106 );
    xnor g15445 ( n16347 , n1611 , n15599 );
    or g15446 ( n33857 , n9195 , n12575 );
    or g15447 ( n5108 , n11455 , n29976 );
    nor g15448 ( n8575 , n31486 , n876 );
    and g15449 ( n8481 , n30568 , n22787 );
    and g15450 ( n26953 , n26562 , n1690 );
    and g15451 ( n21654 , n33159 , n20322 );
    xnor g15452 ( n13858 , n29539 , n18379 );
    xnor g15453 ( n1514 , n16420 , n20849 );
    and g15454 ( n29552 , n26932 , n35661 );
    or g15455 ( n7390 , n9173 , n4172 );
    and g15456 ( n25458 , n33122 , n499 );
    or g15457 ( n18421 , n18204 , n14812 );
    nor g15458 ( n18182 , n18891 , n6548 );
    or g15459 ( n3164 , n14943 , n16543 );
    xnor g15460 ( n1149 , n18493 , n8369 );
    and g15461 ( n8851 , n14878 , n9340 );
    xnor g15462 ( n2887 , n14982 , n35565 );
    or g15463 ( n5272 , n12816 , n17162 );
    and g15464 ( n17081 , n19316 , n19183 );
    and g15465 ( n12069 , n11321 , n27155 );
    or g15466 ( n21557 , n25602 , n22303 );
    and g15467 ( n2080 , n27501 , n23022 );
    not g15468 ( n31991 , n34285 );
    not g15469 ( n19432 , n16223 );
    and g15470 ( n8614 , n627 , n3034 );
    or g15471 ( n28800 , n30774 , n11312 );
    nor g15472 ( n13486 , n4960 , n18636 );
    not g15473 ( n11987 , n5798 );
    or g15474 ( n1674 , n18871 , n10336 );
    xnor g15475 ( n14176 , n34985 , n12437 );
    and g15476 ( n593 , n24970 , n931 );
    or g15477 ( n31471 , n23770 , n5807 );
    xnor g15478 ( n15584 , n3389 , n24371 );
    nor g15479 ( n14341 , n30742 , n21322 );
    nor g15480 ( n13755 , n9425 , n29499 );
    xnor g15481 ( n9076 , n13603 , n5287 );
    xnor g15482 ( n21861 , n12696 , n31957 );
    or g15483 ( n30544 , n1747 , n10289 );
    or g15484 ( n7483 , n21311 , n4595 );
    xnor g15485 ( n28217 , n20188 , n29839 );
    or g15486 ( n26756 , n14244 , n31869 );
    or g15487 ( n35664 , n7441 , n17126 );
    or g15488 ( n5494 , n18765 , n20840 );
    and g15489 ( n20257 , n1092 , n35058 );
    or g15490 ( n11981 , n3146 , n8184 );
    or g15491 ( n33120 , n16620 , n2547 );
    or g15492 ( n32988 , n468 , n19997 );
    xnor g15493 ( n14600 , n6296 , n29713 );
    or g15494 ( n25771 , n31051 , n11589 );
    not g15495 ( n11239 , n2782 );
    xnor g15496 ( n13068 , n29868 , n12781 );
    or g15497 ( n26827 , n14820 , n30995 );
    or g15498 ( n21217 , n830 , n35371 );
    xnor g15499 ( n12263 , n2837 , n17751 );
    and g15500 ( n19076 , n2823 , n24193 );
    or g15501 ( n22372 , n12695 , n10289 );
    or g15502 ( n23510 , n27198 , n8153 );
    or g15503 ( n13874 , n17568 , n13340 );
    or g15504 ( n29777 , n15553 , n27728 );
    buf g15505 ( n8831 , n31665 );
    or g15506 ( n23733 , n29635 , n26332 );
    or g15507 ( n32824 , n9789 , n91 );
    and g15508 ( n33776 , n28660 , n11281 );
    or g15509 ( n8639 , n32225 , n32425 );
    and g15510 ( n17876 , n11289 , n5042 );
    xnor g15511 ( n35690 , n8881 , n3946 );
    or g15512 ( n14123 , n32338 , n30646 );
    xnor g15513 ( n20946 , n20564 , n32063 );
    or g15514 ( n2227 , n11172 , n9601 );
    or g15515 ( n3398 , n33333 , n29686 );
    or g15516 ( n30225 , n32095 , n20191 );
    and g15517 ( n36090 , n30882 , n12336 );
    and g15518 ( n6998 , n29236 , n6004 );
    nor g15519 ( n17286 , n34611 , n21792 );
    xnor g15520 ( n18583 , n15325 , n25974 );
    xnor g15521 ( n9665 , n11056 , n12808 );
    xnor g15522 ( n22300 , n18959 , n22112 );
    and g15523 ( n33152 , n5751 , n20753 );
    or g15524 ( n17453 , n9237 , n3832 );
    and g15525 ( n16166 , n5781 , n26596 );
    xnor g15526 ( n637 , n33715 , n2816 );
    or g15527 ( n5273 , n32107 , n2119 );
    xnor g15528 ( n19785 , n1905 , n15498 );
    or g15529 ( n29595 , n4945 , n5461 );
    buf g15530 ( n34084 , n13098 );
    or g15531 ( n497 , n27217 , n1402 );
    or g15532 ( n1013 , n22802 , n25273 );
    xnor g15533 ( n22296 , n12498 , n22291 );
    and g15534 ( n13186 , n3845 , n6190 );
    or g15535 ( n34477 , n11046 , n27484 );
    xnor g15536 ( n10491 , n17244 , n9793 );
    xnor g15537 ( n11341 , n7765 , n17769 );
    and g15538 ( n2778 , n5621 , n20674 );
    xnor g15539 ( n4390 , n17634 , n34891 );
    or g15540 ( n23622 , n30181 , n30884 );
    nor g15541 ( n34069 , n31788 , n9921 );
    xnor g15542 ( n27018 , n717 , n28751 );
    xnor g15543 ( n4304 , n27027 , n3461 );
    and g15544 ( n8323 , n3872 , n11764 );
    xnor g15545 ( n2008 , n18043 , n31799 );
    not g15546 ( n9202 , n26081 );
    and g15547 ( n26751 , n11090 , n24195 );
    and g15548 ( n75 , n28218 , n18775 );
    or g15549 ( n16535 , n36008 , n16919 );
    xnor g15550 ( n33886 , n1662 , n5116 );
    and g15551 ( n18601 , n34508 , n8987 );
    or g15552 ( n35564 , n6488 , n29411 );
    or g15553 ( n1807 , n1028 , n4478 );
    or g15554 ( n6014 , n13509 , n30708 );
    xnor g15555 ( n23422 , n25672 , n23755 );
    xnor g15556 ( n30922 , n15452 , n22086 );
    not g15557 ( n34909 , n25602 );
    or g15558 ( n12536 , n27020 , n3239 );
    and g15559 ( n20512 , n2212 , n8764 );
    or g15560 ( n19818 , n6701 , n3738 );
    and g15561 ( n21144 , n9909 , n19995 );
    and g15562 ( n29739 , n27390 , n11181 );
    or g15563 ( n1987 , n30688 , n28627 );
    and g15564 ( n14366 , n26620 , n7483 );
    xnor g15565 ( n19192 , n13638 , n17568 );
    xnor g15566 ( n4074 , n31106 , n10822 );
    or g15567 ( n24843 , n5233 , n32305 );
    and g15568 ( n4217 , n22428 , n24065 );
    xnor g15569 ( n33646 , n142 , n11046 );
    or g15570 ( n33194 , n14496 , n4965 );
    and g15571 ( n17604 , n16675 , n8773 );
    not g15572 ( n34451 , n16985 );
    or g15573 ( n14550 , n11123 , n33556 );
    or g15574 ( n29601 , n3320 , n14725 );
    or g15575 ( n14448 , n10924 , n34873 );
    or g15576 ( n26946 , n19302 , n5516 );
    or g15577 ( n1491 , n16068 , n33713 );
    xnor g15578 ( n32820 , n9949 , n7439 );
    and g15579 ( n3115 , n31309 , n18212 );
    and g15580 ( n31718 , n29700 , n4503 );
    or g15581 ( n2605 , n9658 , n24545 );
    xnor g15582 ( n11532 , n4787 , n16620 );
    and g15583 ( n33923 , n26009 , n15760 );
    or g15584 ( n24688 , n19133 , n34036 );
    xnor g15585 ( n29778 , n24286 , n25174 );
    xnor g15586 ( n16955 , n933 , n29839 );
    and g15587 ( n13795 , n1281 , n29415 );
    xnor g15588 ( n32645 , n4651 , n27793 );
    and g15589 ( n35313 , n10470 , n3656 );
    or g15590 ( n8009 , n17751 , n28108 );
    xnor g15591 ( n28838 , n14029 , n27186 );
    or g15592 ( n9707 , n5090 , n20579 );
    not g15593 ( n34620 , n1429 );
    not g15594 ( n9240 , n3168 );
    or g15595 ( n34241 , n4266 , n24505 );
    xnor g15596 ( n5979 , n34914 , n4403 );
    xnor g15597 ( n17105 , n15882 , n5161 );
    xnor g15598 ( n4245 , n1706 , n7055 );
    xnor g15599 ( n6189 , n11881 , n16922 );
    xnor g15600 ( n8373 , n33066 , n23060 );
    and g15601 ( n16840 , n26691 , n1677 );
    xnor g15602 ( n32668 , n32082 , n25593 );
    xnor g15603 ( n8777 , n2417 , n20758 );
    buf g15604 ( n3437 , n14051 );
    not g15605 ( n26263 , n29203 );
    and g15606 ( n3184 , n32398 , n30051 );
    or g15607 ( n22323 , n22715 , n12858 );
    or g15608 ( n21011 , n31394 , n4590 );
    xnor g15609 ( n33537 , n6535 , n20721 );
    and g15610 ( n23685 , n30035 , n33012 );
    xnor g15611 ( n34519 , n18847 , n9037 );
    not g15612 ( n1341 , n32095 );
    or g15613 ( n10643 , n14001 , n17915 );
    or g15614 ( n14255 , n5335 , n21102 );
    and g15615 ( n24361 , n14857 , n15674 );
    and g15616 ( n27701 , n18522 , n25325 );
    xnor g15617 ( n29507 , n9499 , n23769 );
    or g15618 ( n6171 , n6015 , n33139 );
    and g15619 ( n26243 , n27556 , n22853 );
    or g15620 ( n15192 , n31799 , n23169 );
    not g15621 ( n33302 , n25602 );
    nor g15622 ( n7297 , n22291 , n1440 );
    xnor g15623 ( n21062 , n10378 , n22967 );
    nor g15624 ( n17818 , n12202 , n21760 );
    and g15625 ( n24054 , n6808 , n11109 );
    not g15626 ( n30253 , n16620 );
    and g15627 ( n31587 , n15159 , n32951 );
    or g15628 ( n31081 , n27267 , n27973 );
    nor g15629 ( n26895 , n8432 , n5936 );
    or g15630 ( n1844 , n11046 , n4357 );
    or g15631 ( n2696 , n2138 , n24356 );
    not g15632 ( n10074 , n22980 );
    and g15633 ( n22738 , n14675 , n34773 );
    or g15634 ( n12672 , n17321 , n4254 );
    or g15635 ( n30269 , n16495 , n1605 );
    and g15636 ( n27994 , n33035 , n25590 );
    nor g15637 ( n35912 , n32857 , n25043 );
    not g15638 ( n17000 , n7801 );
    nor g15639 ( n10516 , n9789 , n1115 );
    or g15640 ( n15721 , n17487 , n9915 );
    or g15641 ( n22092 , n9950 , n18148 );
    xnor g15642 ( n17351 , n13300 , n19551 );
    xnor g15643 ( n34424 , n21799 , n24371 );
    and g15644 ( n4975 , n17734 , n1450 );
    or g15645 ( n15123 , n16135 , n25783 );
    not g15646 ( n1583 , n22501 );
    not g15647 ( n16571 , n5335 );
    not g15648 ( n25625 , n19939 );
    nor g15649 ( n29890 , n27291 , n19532 );
    and g15650 ( n7110 , n11619 , n28156 );
    or g15651 ( n17599 , n19604 , n16803 );
    and g15652 ( n1627 , n28881 , n7121 );
    or g15653 ( n26231 , n32601 , n14486 );
    or g15654 ( n30005 , n15886 , n7068 );
    or g15655 ( n21824 , n3658 , n2338 );
    xnor g15656 ( n28368 , n6759 , n6456 );
    and g15657 ( n26517 , n9402 , n18044 );
    and g15658 ( n8375 , n9608 , n25072 );
    not g15659 ( n2443 , n11190 );
    nor g15660 ( n33216 , n27603 , n24177 );
    or g15661 ( n5536 , n7399 , n20812 );
    and g15662 ( n28431 , n10059 , n21429 );
    or g15663 ( n18290 , n19397 , n21361 );
    xnor g15664 ( n19184 , n11626 , n4929 );
    not g15665 ( n3703 , n13170 );
    and g15666 ( n22280 , n1011 , n22688 );
    xnor g15667 ( n32041 , n20084 , n4960 );
    buf g15668 ( n28404 , n24513 );
    nor g15669 ( n34165 , n34988 , n7726 );
    or g15670 ( n19389 , n22429 , n908 );
    or g15671 ( n29414 , n10932 , n20722 );
    or g15672 ( n3963 , n11468 , n31606 );
    and g15673 ( n26074 , n18702 , n21341 );
    or g15674 ( n26169 , n35558 , n7726 );
    not g15675 ( n7054 , n34780 );
    and g15676 ( n6266 , n9330 , n26249 );
    and g15677 ( n19819 , n26523 , n29971 );
    or g15678 ( n19343 , n11455 , n17288 );
    or g15679 ( n14262 , n33723 , n181 );
    or g15680 ( n18447 , n23010 , n13664 );
    and g15681 ( n5093 , n33819 , n21001 );
    xnor g15682 ( n19363 , n26817 , n6489 );
    or g15683 ( n516 , n10471 , n8710 );
    or g15684 ( n5342 , n32027 , n3979 );
    or g15685 ( n17260 , n6477 , n6288 );
    not g15686 ( n23256 , n14677 );
    xnor g15687 ( n17980 , n18453 , n11351 );
    xnor g15688 ( n3929 , n23744 , n12654 );
    or g15689 ( n26066 , n28102 , n30764 );
    or g15690 ( n21341 , n2311 , n4203 );
    not g15691 ( n19556 , n6916 );
    or g15692 ( n18446 , n6465 , n17045 );
    and g15693 ( n22370 , n24223 , n24071 );
    xnor g15694 ( n18564 , n17586 , n17681 );
    not g15695 ( n15782 , n24371 );
    and g15696 ( n22483 , n27207 , n17860 );
    or g15697 ( n4602 , n3205 , n35108 );
    xnor g15698 ( n30502 , n4825 , n20277 );
    and g15699 ( n30395 , n31891 , n34426 );
    or g15700 ( n27054 , n21288 , n14746 );
    or g15701 ( n3284 , n14906 , n4706 );
    or g15702 ( n6170 , n4757 , n16213 );
    or g15703 ( n20414 , n31601 , n27501 );
    not g15704 ( n27265 , n14965 );
    or g15705 ( n31752 , n830 , n174 );
    or g15706 ( n9420 , n33752 , n4912 );
    not g15707 ( n11513 , n10221 );
    and g15708 ( n2730 , n7196 , n10949 );
    not g15709 ( n32861 , n2684 );
    and g15710 ( n7197 , n14243 , n32450 );
    or g15711 ( n809 , n27808 , n14700 );
    and g15712 ( n19718 , n1203 , n16040 );
    or g15713 ( n18335 , n14688 , n19084 );
    xnor g15714 ( n12348 , n15226 , n25602 );
    xnor g15715 ( n17261 , n21014 , n4962 );
    and g15716 ( n7636 , n14250 , n27836 );
    or g15717 ( n26213 , n21711 , n31496 );
    xor g15718 ( n35740 , n16644 , n24371 );
    and g15719 ( n5115 , n26191 , n2288 );
    nor g15720 ( n24757 , n14775 , n15980 );
    nor g15721 ( n10377 , n16620 , n32780 );
    xnor g15722 ( n31242 , n28106 , n9789 );
    xnor g15723 ( n28617 , n21980 , n18623 );
    not g15724 ( n28907 , n33499 );
    and g15725 ( n9952 , n243 , n25797 );
    or g15726 ( n6892 , n16324 , n27501 );
    or g15727 ( n13391 , n25730 , n12996 );
    xnor g15728 ( n4845 , n34283 , n31272 );
    xnor g15729 ( n12013 , n19951 , n4962 );
    and g15730 ( n26929 , n25859 , n17444 );
    and g15731 ( n23099 , n27975 , n10868 );
    and g15732 ( n20963 , n4323 , n3152 );
    xnor g15733 ( n1127 , n16302 , n5335 );
    not g15734 ( n33482 , n32619 );
    or g15735 ( n14920 , n3205 , n3379 );
    or g15736 ( n13693 , n830 , n7823 );
    and g15737 ( n780 , n10659 , n7482 );
    xnor g15738 ( n12374 , n12734 , n7540 );
    or g15739 ( n2461 , n28405 , n5208 );
    or g15740 ( n23659 , n26637 , n4239 );
    and g15741 ( n29984 , n19920 , n20248 );
    xnor g15742 ( n23519 , n10320 , n9789 );
    or g15743 ( n9519 , n15464 , n1156 );
    or g15744 ( n30191 , n32584 , n2729 );
    and g15745 ( n3803 , n14513 , n30859 );
    or g15746 ( n1559 , n7540 , n34844 );
    or g15747 ( n27654 , n29713 , n18694 );
    or g15748 ( n9458 , n14741 , n4348 );
    or g15749 ( n4791 , n21073 , n12895 );
    not g15750 ( n21631 , n9658 );
    and g15751 ( n10139 , n35444 , n3585 );
    or g15752 ( n31836 , n7772 , n8153 );
    and g15753 ( n10900 , n12145 , n8847 );
    or g15754 ( n30623 , n1938 , n8928 );
    or g15755 ( n25639 , n31289 , n12801 );
    or g15756 ( n12071 , n23687 , n15145 );
    or g15757 ( n8562 , n15469 , n12377 );
    or g15758 ( n12040 , n25174 , n34066 );
    xnor g15759 ( n14253 , n32051 , n19648 );
    or g15760 ( n9292 , n19551 , n24229 );
    or g15761 ( n12220 , n30522 , n31549 );
    or g15762 ( n7531 , n8432 , n32838 );
    nor g15763 ( n27854 , n31101 , n29448 );
    not g15764 ( n29977 , n32095 );
    or g15765 ( n24416 , n18429 , n2119 );
    and g15766 ( n20478 , n8738 , n28709 );
    or g15767 ( n603 , n24319 , n28894 );
    or g15768 ( n4158 , n4449 , n14918 );
    xnor g15769 ( n12077 , n15258 , n4930 );
    or g15770 ( n3134 , n2209 , n13028 );
    and g15771 ( n24374 , n28738 , n14772 );
    and g15772 ( n17961 , n24572 , n19352 );
    and g15773 ( n33454 , n27931 , n64 );
    nor g15774 ( n20240 , n19551 , n28834 );
    or g15775 ( n15823 , n33433 , n19464 );
    xnor g15776 ( n1808 , n11645 , n12697 );
    xnor g15777 ( n8093 , n21786 , n16582 );
    xnor g15778 ( n17804 , n24054 , n21508 );
    or g15779 ( n21545 , n5335 , n24138 );
    or g15780 ( n8040 , n25518 , n9053 );
    and g15781 ( n10087 , n9087 , n10912 );
    xnor g15782 ( n8052 , n13845 , n19664 );
    and g15783 ( n15791 , n32810 , n6813 );
    and g15784 ( n15303 , n1464 , n22528 );
    and g15785 ( n5146 , n5247 , n26487 );
    not g15786 ( n14791 , n23179 );
    not g15787 ( n12806 , n7540 );
    or g15788 ( n21291 , n34292 , n9403 );
    nor g15789 ( n34488 , n9789 , n14905 );
    or g15790 ( n1116 , n30902 , n4254 );
    or g15791 ( n20665 , n4377 , n27583 );
    and g15792 ( n34414 , n16917 , n27526 );
    or g15793 ( n4614 , n5723 , n8366 );
    xnor g15794 ( n16981 , n34439 , n283 );
    xnor g15795 ( n2281 , n13284 , n23604 );
    and g15796 ( n18881 , n12255 , n9002 );
    xnor g15797 ( n3794 , n15959 , n10894 );
    or g15798 ( n30930 , n1115 , n33275 );
    not g15799 ( n12742 , n19159 );
    xnor g15800 ( n25299 , n16563 , n18242 );
    xnor g15801 ( n18120 , n14780 , n3946 );
    nor g15802 ( n1360 , n22291 , n25644 );
    xnor g15803 ( n28767 , n25858 , n8432 );
    and g15804 ( n1181 , n31390 , n9561 );
    and g15805 ( n17259 , n32487 , n5239 );
    and g15806 ( n18106 , n1952 , n14066 );
    or g15807 ( n32034 , n3170 , n733 );
    not g15808 ( n16488 , n29879 );
    nor g15809 ( n23585 , n35927 , n941 );
    or g15810 ( n28238 , n14648 , n25831 );
    or g15811 ( n21910 , n11162 , n25648 );
    xnor g15812 ( n9172 , n3364 , n4288 );
    not g15813 ( n17761 , n22362 );
    and g15814 ( n23494 , n17473 , n5951 );
    xnor g15815 ( n17748 , n10703 , n1543 );
    or g15816 ( n5100 , n32527 , n11571 );
    xnor g15817 ( n7138 , n35163 , n25825 );
    or g15818 ( n4054 , n19186 , n10847 );
    or g15819 ( n22347 , n30633 , n20628 );
    xnor g15820 ( n28860 , n17178 , n3946 );
    or g15821 ( n23172 , n24424 , n1019 );
    or g15822 ( n19063 , n9600 , n17872 );
    or g15823 ( n12614 , n36014 , n30708 );
    or g15824 ( n10775 , n26488 , n31455 );
    or g15825 ( n34757 , n378 , n3815 );
    or g15826 ( n15681 , n23459 , n20797 );
    or g15827 ( n5147 , n33079 , n9780 );
    not g15828 ( n6276 , n12666 );
    nor g15829 ( n29047 , n4758 , n21180 );
    or g15830 ( n16931 , n19283 , n25567 );
    and g15831 ( n7571 , n27387 , n13762 );
    nor g15832 ( n6558 , n4288 , n7144 );
    or g15833 ( n23496 , n17033 , n16385 );
    or g15834 ( n28258 , n20398 , n3762 );
    and g15835 ( n21803 , n1951 , n10240 );
    not g15836 ( n1430 , n3205 );
    and g15837 ( n32641 , n27083 , n9284 );
    not g15838 ( n28566 , n9431 );
    or g15839 ( n12426 , n31559 , n27611 );
    or g15840 ( n35509 , n12521 , n14271 );
    or g15841 ( n1781 , n12212 , n7773 );
    not g15842 ( n2195 , n12667 );
    or g15843 ( n800 , n4386 , n7815 );
    nor g15844 ( n30795 , n9658 , n22975 );
    and g15845 ( n17736 , n15672 , n22925 );
    or g15846 ( n17245 , n28879 , n2823 );
    xnor g15847 ( n12740 , n31736 , n29713 );
    and g15848 ( n25927 , n28828 , n32430 );
    or g15849 ( n3464 , n7540 , n34142 );
    or g15850 ( n26644 , n26529 , n12332 );
    buf g15851 ( n17612 , n17005 );
    xnor g15852 ( n3365 , n23292 , n22455 );
    or g15853 ( n2839 , n15854 , n34501 );
    not g15854 ( n3423 , n31272 );
    nor g15855 ( n12664 , n8982 , n22657 );
    or g15856 ( n13108 , n24791 , n17354 );
    or g15857 ( n18404 , n26801 , n33279 );
    or g15858 ( n8160 , n29884 , n7139 );
    or g15859 ( n5712 , n19394 , n15517 );
    or g15860 ( n22521 , n8147 , n16905 );
    not g15861 ( n28036 , n9254 );
    xnor g15862 ( n10396 , n1370 , n25602 );
    or g15863 ( n2930 , n18224 , n28347 );
    and g15864 ( n22672 , n5449 , n23818 );
    or g15865 ( n20730 , n2887 , n23921 );
    xnor g15866 ( n28795 , n18261 , n25842 );
    or g15867 ( n14203 , n19078 , n13384 );
    and g15868 ( n34738 , n9880 , n861 );
    and g15869 ( n11897 , n5756 , n26030 );
    or g15870 ( n27988 , n11709 , n25255 );
    buf g15871 ( n6459 , n10083 );
    or g15872 ( n31280 , n8290 , n18101 );
    or g15873 ( n21876 , n24453 , n10489 );
    or g15874 ( n22033 , n5067 , n20152 );
    and g15875 ( n8008 , n5012 , n19647 );
    xnor g15876 ( n33804 , n30313 , n4962 );
    and g15877 ( n8735 , n18016 , n1844 );
    or g15878 ( n1417 , n31535 , n1557 );
    and g15879 ( n15249 , n22740 , n13237 );
    not g15880 ( n5607 , n16594 );
    and g15881 ( n13912 , n11718 , n27974 );
    or g15882 ( n21661 , n21774 , n11312 );
    xnor g15883 ( n21190 , n22301 , n4878 );
    nor g15884 ( n720 , n20881 , n3346 );
    and g15885 ( n34060 , n3469 , n15515 );
    xnor g15886 ( n21178 , n33788 , n25990 );
    xnor g15887 ( n29442 , n7382 , n4925 );
    or g15888 ( n13536 , n4878 , n19099 );
    or g15889 ( n31673 , n11872 , n13217 );
    xnor g15890 ( n15912 , n32153 , n28434 );
    and g15891 ( n1605 , n28957 , n7260 );
    and g15892 ( n30124 , n17914 , n13388 );
    xnor g15893 ( n31690 , n36036 , n24263 );
    or g15894 ( n34252 , n23065 , n21956 );
    or g15895 ( n12045 , n7282 , n1171 );
    or g15896 ( n9630 , n23558 , n25831 );
    or g15897 ( n8620 , n29839 , n27690 );
    or g15898 ( n10848 , n30630 , n26924 );
    xnor g15899 ( n9414 , n29422 , n28839 );
    and g15900 ( n20360 , n23607 , n31652 );
    or g15901 ( n8922 , n32448 , n28324 );
    and g15902 ( n32225 , n5896 , n23105 );
    or g15903 ( n32926 , n25317 , n7293 );
    and g15904 ( n3223 , n17253 , n35357 );
    nor g15905 ( n7514 , n14846 , n3808 );
    or g15906 ( n27934 , n31736 , n10336 );
    nor g15907 ( n26460 , n16620 , n17188 );
    not g15908 ( n30264 , n10147 );
    xnor g15909 ( n4908 , n3368 , n24371 );
    xnor g15910 ( n36016 , n28489 , n4960 );
    nor g15911 ( n22466 , n15228 , n16649 );
    nor g15912 ( n14904 , n9789 , n29993 );
    xnor g15913 ( n10657 , n28517 , n23819 );
    or g15914 ( n25498 , n5335 , n16000 );
    or g15915 ( n8659 , n3946 , n5612 );
    or g15916 ( n3226 , n15043 , n13165 );
    and g15917 ( n28559 , n24952 , n26742 );
    xnor g15918 ( n26304 , n1099 , n22737 );
    xnor g15919 ( n1611 , n32597 , n830 );
    and g15920 ( n24841 , n18822 , n25723 );
    or g15921 ( n11061 , n9518 , n10479 );
    and g15922 ( n30752 , n21475 , n16271 );
    xnor g15923 ( n23034 , n4842 , n11455 );
    and g15924 ( n20143 , n9127 , n12019 );
    nor g15925 ( n21236 , n24371 , n13533 );
    nor g15926 ( n19904 , n22246 , n6988 );
    or g15927 ( n32788 , n12150 , n30697 );
    not g15928 ( n7902 , n32995 );
    or g15929 ( n33437 , n27038 , n32391 );
    or g15930 ( n7012 , n8691 , n210 );
    or g15931 ( n3024 , n2155 , n32507 );
    or g15932 ( n15561 , n30434 , n9915 );
    or g15933 ( n4533 , n26556 , n2955 );
    xnor g15934 ( n17241 , n34646 , n9969 );
    and g15935 ( n24457 , n9026 , n22414 );
    xnor g15936 ( n10696 , n27718 , n20120 );
    or g15937 ( n2830 , n416 , n31687 );
    or g15938 ( n30663 , n36006 , n24756 );
    or g15939 ( n9405 , n26615 , n2712 );
    and g15940 ( n1113 , n10536 , n11405 );
    nor g15941 ( n24414 , n32857 , n24520 );
    xnor g15942 ( n26688 , n18475 , n16228 );
    not g15943 ( n18509 , n14994 );
    xnor g15944 ( n19535 , n5304 , n7830 );
    xnor g15945 ( n8260 , n5552 , n17568 );
    or g15946 ( n15430 , n28554 , n22206 );
    or g15947 ( n9802 , n24173 , n1098 );
    nor g15948 ( n24750 , n30603 , n32379 );
    not g15949 ( n1756 , n3858 );
    xnor g15950 ( n18681 , n17250 , n16135 );
    or g15951 ( n3971 , n24371 , n14842 );
    and g15952 ( n394 , n27651 , n34790 );
    or g15953 ( n10123 , n32227 , n24259 );
    or g15954 ( n29615 , n27897 , n24356 );
    not g15955 ( n33102 , n34100 );
    or g15956 ( n11032 , n11817 , n17640 );
    or g15957 ( n20496 , n2824 , n19105 );
    xnor g15958 ( n3428 , n32686 , n21233 );
    or g15959 ( n28515 , n28860 , n21301 );
    and g15960 ( n14632 , n16349 , n19160 );
    or g15961 ( n30324 , n29984 , n25773 );
    nor g15962 ( n24017 , n24932 , n29759 );
    and g15963 ( n18612 , n10413 , n9399 );
    or g15964 ( n18609 , n15959 , n33435 );
    or g15965 ( n29947 , n16818 , n18488 );
    xnor g15966 ( n1120 , n8632 , n9789 );
    or g15967 ( n5869 , n17232 , n15946 );
    or g15968 ( n21947 , n35669 , n28023 );
    or g15969 ( n35122 , n13550 , n30419 );
    or g15970 ( n25120 , n16956 , n4952 );
    or g15971 ( n3172 , n7765 , n17769 );
    and g15972 ( n5451 , n902 , n23609 );
    or g15973 ( n3331 , n30897 , n31083 );
    or g15974 ( n264 , n24311 , n10872 );
    xnor g15975 ( n15125 , n6044 , n7412 );
    or g15976 ( n22669 , n3406 , n20906 );
    or g15977 ( n29750 , n17585 , n21419 );
    or g15978 ( n25805 , n35927 , n31194 );
    not g15979 ( n35326 , n9793 );
    or g15980 ( n11983 , n32095 , n615 );
    not g15981 ( n23261 , n1111 );
    or g15982 ( n23909 , n26058 , n34287 );
    and g15983 ( n5654 , n25739 , n16706 );
    xnor g15984 ( n2982 , n9980 , n16038 );
    buf g15985 ( n6553 , n14018 );
    or g15986 ( n13166 , n3946 , n20678 );
    or g15987 ( n33316 , n8852 , n17612 );
    or g15988 ( n1788 , n32095 , n13148 );
    xnor g15989 ( n28988 , n29719 , n5103 );
    not g15990 ( n27202 , n23237 );
    or g15991 ( n7757 , n27680 , n30687 );
    xnor g15992 ( n1425 , n32127 , n20066 );
    not g15993 ( n33882 , n20061 );
    nor g15994 ( n23113 , n18943 , n13975 );
    and g15995 ( n26892 , n25085 , n32279 );
    xnor g15996 ( n1012 , n34926 , n2780 );
    xnor g15997 ( n14353 , n32241 , n34437 );
    or g15998 ( n31041 , n31141 , n5080 );
    xnor g15999 ( n8419 , n14624 , n13347 );
    or g16000 ( n11677 , n19102 , n20590 );
    xnor g16001 ( n14266 , n3488 , n368 );
    or g16002 ( n20890 , n6123 , n24412 );
    xnor g16003 ( n521 , n14435 , n21456 );
    or g16004 ( n27477 , n14735 , n14841 );
    or g16005 ( n14044 , n24371 , n6741 );
    or g16006 ( n11720 , n24183 , n6046 );
    nor g16007 ( n32076 , n33695 , n2144 );
    not g16008 ( n3847 , n7726 );
    xnor g16009 ( n29209 , n14530 , n11200 );
    not g16010 ( n27386 , n31506 );
    or g16011 ( n18355 , n4629 , n10336 );
    xnor g16012 ( n5577 , n14842 , n24371 );
    and g16013 ( n11144 , n22631 , n11900 );
    xnor g16014 ( n15000 , n34271 , n28734 );
    or g16015 ( n32653 , n20404 , n17270 );
    xnor g16016 ( n17578 , n5195 , n30742 );
    and g16017 ( n35493 , n33565 , n17738 );
    and g16018 ( n12354 , n14398 , n29219 );
    and g16019 ( n35132 , n23236 , n16584 );
    xnor g16020 ( n34469 , n12597 , n13072 );
    or g16021 ( n23615 , n27919 , n23748 );
    or g16022 ( n22021 , n26787 , n20739 );
    or g16023 ( n9608 , n29385 , n13241 );
    or g16024 ( n7764 , n1986 , n3818 );
    not g16025 ( n14264 , n31289 );
    or g16026 ( n11843 , n7030 , n4952 );
    or g16027 ( n11121 , n32739 , n17962 );
    or g16028 ( n26629 , n23945 , n22682 );
    or g16029 ( n28454 , n25 , n23319 );
    and g16030 ( n24765 , n26433 , n582 );
    and g16031 ( n27919 , n17795 , n7085 );
    or g16032 ( n19146 , n20445 , n33358 );
    and g16033 ( n3802 , n2974 , n5825 );
    nor g16034 ( n2583 , n15671 , n3437 );
    or g16035 ( n31909 , n33084 , n27728 );
    not g16036 ( n14595 , n29964 );
    xnor g16037 ( n23022 , n19225 , n28867 );
    or g16038 ( n14367 , n34221 , n5208 );
    buf g16039 ( n1414 , n19952 );
    or g16040 ( n19770 , n32715 , n8440 );
    and g16041 ( n22062 , n35026 , n35365 );
    or g16042 ( n9270 , n7392 , n29783 );
    and g16043 ( n28114 , n21597 , n16074 );
    or g16044 ( n34245 , n34602 , n35934 );
    not g16045 ( n1737 , n28482 );
    xnor g16046 ( n20751 , n7285 , n8063 );
    or g16047 ( n18663 , n18925 , n21524 );
    or g16048 ( n2395 , n31419 , n14775 );
    or g16049 ( n3767 , n32715 , n16972 );
    not g16050 ( n28816 , n25592 );
    and g16051 ( n32419 , n9300 , n21050 );
    xnor g16052 ( n17585 , n2284 , n22291 );
    or g16053 ( n34291 , n4960 , n32785 );
    and g16054 ( n2880 , n32423 , n28081 );
    nor g16055 ( n7802 , n5335 , n20132 );
    or g16056 ( n33361 , n10559 , n28404 );
    or g16057 ( n32222 , n25602 , n8103 );
    or g16058 ( n5258 , n4391 , n12595 );
    and g16059 ( n313 , n1705 , n19974 );
    not g16060 ( n27570 , n30742 );
    xnor g16061 ( n10208 , n7378 , n4512 );
    or g16062 ( n11688 , n20485 , n30419 );
    and g16063 ( n24860 , n8161 , n7652 );
    or g16064 ( n11989 , n31559 , n34150 );
    or g16065 ( n35301 , n21119 , n20813 );
    or g16066 ( n20009 , n2744 , n7289 );
    not g16067 ( n17816 , n30742 );
    and g16068 ( n6309 , n5911 , n18376 );
    nor g16069 ( n26188 , n1950 , n34212 );
    or g16070 ( n6478 , n9709 , n6543 );
    and g16071 ( n11424 , n35416 , n21969 );
    xnor g16072 ( n9718 , n1515 , n3946 );
    and g16073 ( n29707 , n31931 , n15129 );
    and g16074 ( n7943 , n1506 , n28341 );
    xnor g16075 ( n3421 , n32106 , n7315 );
    xnor g16076 ( n32945 , n11529 , n22051 );
    not g16077 ( n7817 , n18287 );
    or g16078 ( n6921 , n27245 , n26166 );
    and g16079 ( n32872 , n1025 , n8306 );
    not g16080 ( n26646 , n28287 );
    or g16081 ( n26838 , n3985 , n23281 );
    and g16082 ( n13055 , n11028 , n18379 );
    and g16083 ( n14221 , n20350 , n11974 );
    xnor g16084 ( n25203 , n2236 , n24553 );
    or g16085 ( n28118 , n1898 , n30419 );
    and g16086 ( n11827 , n6978 , n32830 );
    xnor g16087 ( n18503 , n28913 , n4432 );
    and g16088 ( n35692 , n1835 , n17496 );
    nor g16089 ( n14083 , n30160 , n14757 );
    or g16090 ( n28688 , n29839 , n4976 );
    and g16091 ( n33250 , n18311 , n17667 );
    not g16092 ( n30526 , n8638 );
    or g16093 ( n14581 , n22941 , n7553 );
    or g16094 ( n17939 , n10772 , n8587 );
    xnor g16095 ( n10062 , n26505 , n6133 );
    not g16096 ( n6050 , n22021 );
    nor g16097 ( n35983 , n13239 , n1796 );
    xnor g16098 ( n12637 , n15953 , n2538 );
    or g16099 ( n11332 , n21990 , n3352 );
    not g16100 ( n4142 , n22980 );
    and g16101 ( n32716 , n13764 , n19035 );
    and g16102 ( n21078 , n5624 , n14482 );
    xnor g16103 ( n22675 , n7442 , n5287 );
    or g16104 ( n1475 , n10841 , n1511 );
    or g16105 ( n22895 , n29713 , n25794 );
    and g16106 ( n23365 , n19393 , n19382 );
    xnor g16107 ( n17607 , n13508 , n34610 );
    or g16108 ( n28896 , n29884 , n3923 );
    or g16109 ( n6530 , n23884 , n2168 );
    or g16110 ( n13063 , n8037 , n8921 );
    or g16111 ( n31938 , n18321 , n21862 );
    or g16112 ( n19893 , n1235 , n12419 );
    nor g16113 ( n35038 , n12323 , n29941 );
    not g16114 ( n23871 , n8731 );
    and g16115 ( n26046 , n28621 , n15721 );
    or g16116 ( n32489 , n16073 , n1942 );
    and g16117 ( n26613 , n35223 , n1584 );
    xnor g16118 ( n19000 , n23754 , n31255 );
    not g16119 ( n19561 , n25387 );
    xnor g16120 ( n27636 , n15846 , n4960 );
    and g16121 ( n2757 , n3500 , n8967 );
    xnor g16122 ( n7684 , n26649 , n5440 );
    or g16123 ( n31511 , n12169 , n15496 );
    or g16124 ( n34362 , n29101 , n23113 );
    or g16125 ( n5373 , n25203 , n28668 );
    xnor g16126 ( n18262 , n8005 , n21305 );
    xnor g16127 ( n34341 , n27215 , n18080 );
    xnor g16128 ( n15949 , n1383 , n14411 );
    or g16129 ( n16558 , n12091 , n18045 );
    xnor g16130 ( n3978 , n30525 , n4722 );
    xnor g16131 ( n34978 , n25199 , n5188 );
    or g16132 ( n8460 , n5704 , n16543 );
    and g16133 ( n15982 , n24591 , n18786 );
    not g16134 ( n14736 , n6283 );
    and g16135 ( n35386 , n26387 , n20792 );
    or g16136 ( n29289 , n19545 , n34591 );
    xnor g16137 ( n18415 , n3873 , n32803 );
    or g16138 ( n32258 , n7589 , n27501 );
    and g16139 ( n14847 , n26795 , n13125 );
    and g16140 ( n17208 , n12333 , n5365 );
    xnor g16141 ( n33643 , n16219 , n23604 );
    or g16142 ( n26547 , n12207 , n11601 );
    xnor g16143 ( n18132 , n23924 , n30742 );
    or g16144 ( n24390 , n35202 , n27053 );
    and g16145 ( n5807 , n884 , n24464 );
    or g16146 ( n9149 , n21512 , n23790 );
    or g16147 ( n33385 , n3637 , n2104 );
    and g16148 ( n18871 , n28442 , n26122 );
    and g16149 ( n4129 , n21750 , n34325 );
    or g16150 ( n8385 , n18493 , n8369 );
    and g16151 ( n14073 , n30201 , n34295 );
    or g16152 ( n27148 , n18197 , n5023 );
    xnor g16153 ( n23647 , n13292 , n17170 );
    or g16154 ( n23338 , n19618 , n6012 );
    xnor g16155 ( n13438 , n3810 , n17751 );
    nor g16156 ( n19779 , n11455 , n24959 );
    not g16157 ( n15184 , n35721 );
    nor g16158 ( n28653 , n3205 , n28021 );
    and g16159 ( n16767 , n28504 , n29175 );
    and g16160 ( n22942 , n17400 , n1167 );
    nor g16161 ( n31479 , n6025 , n12107 );
    or g16162 ( n23874 , n18755 , n9672 );
    nor g16163 ( n18976 , n10370 , n34990 );
    or g16164 ( n20007 , n32016 , n138 );
    and g16165 ( n19915 , n21093 , n19774 );
    or g16166 ( n13314 , n10809 , n30204 );
    or g16167 ( n35480 , n1665 , n27728 );
    and g16168 ( n19169 , n13650 , n23765 );
    and g16169 ( n6002 , n15521 , n33479 );
    and g16170 ( n8749 , n12180 , n26343 );
    xnor g16171 ( n22739 , n9621 , n6750 );
    nor g16172 ( n3023 , n25602 , n5593 );
    and g16173 ( n13104 , n23892 , n24190 );
    or g16174 ( n26086 , n29034 , n21477 );
    xnor g16175 ( n13154 , n26424 , n30742 );
    or g16176 ( n18853 , n33232 , n27973 );
    and g16177 ( n16641 , n27477 , n30258 );
    or g16178 ( n35549 , n32304 , n25786 );
    or g16179 ( n12224 , n5335 , n19629 );
    or g16180 ( n6924 , n3205 , n29390 );
    and g16181 ( n14045 , n5978 , n18642 );
    or g16182 ( n33087 , n29512 , n33940 );
    or g16183 ( n34376 , n15637 , n11996 );
    xnor g16184 ( n13995 , n2459 , n11663 );
    and g16185 ( n1183 , n2496 , n28807 );
    not g16186 ( n16639 , n22997 );
    xnor g16187 ( n31110 , n1843 , n35466 );
    not g16188 ( n594 , n1009 );
    and g16189 ( n8192 , n31940 , n5287 );
    and g16190 ( n3165 , n32057 , n15348 );
    nor g16191 ( n14316 , n20138 , n12522 );
    and g16192 ( n14223 , n7043 , n270 );
    or g16193 ( n17904 , n10894 , n113 );
    xnor g16194 ( n15512 , n26038 , n30989 );
    or g16195 ( n13959 , n32915 , n23308 );
    xnor g16196 ( n10357 , n2045 , n33400 );
    or g16197 ( n26120 , n7413 , n33751 );
    or g16198 ( n33876 , n22700 , n35143 );
    or g16199 ( n26221 , n28217 , n27968 );
    or g16200 ( n15592 , n11359 , n24356 );
    nor g16201 ( n19583 , n31329 , n31291 );
    xnor g16202 ( n5408 , n12797 , n19551 );
    xnor g16203 ( n7499 , n4707 , n24371 );
    not g16204 ( n27705 , n9789 );
    or g16205 ( n10502 , n9658 , n31236 );
    xnor g16206 ( n34586 , n26973 , n11046 );
    xnor g16207 ( n24991 , n25954 , n8857 );
    or g16208 ( n21406 , n16922 , n32735 );
    and g16209 ( n7835 , n20533 , n1550 );
    or g16210 ( n28336 , n14904 , n32769 );
    or g16211 ( n10272 , n4723 , n22213 );
    or g16212 ( n7181 , n19914 , n4490 );
    not g16213 ( n29718 , n15233 );
    or g16214 ( n1574 , n1950 , n14674 );
    or g16215 ( n24378 , n9611 , n30621 );
    nor g16216 ( n29874 , n31056 , n25166 );
    xnor g16217 ( n14487 , n3816 , n18921 );
    or g16218 ( n6408 , n24421 , n20399 );
    or g16219 ( n11761 , n25928 , n32889 );
    and g16220 ( n33593 , n13363 , n2673 );
    not g16221 ( n5771 , n23089 );
    and g16222 ( n31453 , n29860 , n16541 );
    and g16223 ( n30399 , n6816 , n32464 );
    buf g16224 ( n32071 , n13211 );
    or g16225 ( n28491 , n29839 , n424 );
    or g16226 ( n17010 , n31559 , n27741 );
    xor g16227 ( n33068 , n12772 , n27138 );
    or g16228 ( n8331 , n16718 , n7553 );
    xnor g16229 ( n21288 , n23035 , n32750 );
    or g16230 ( n31816 , n15719 , n585 );
    nor g16231 ( n14955 , n15464 , n33919 );
    and g16232 ( n31546 , n31351 , n23124 );
    not g16233 ( n17043 , n11607 );
    and g16234 ( n20847 , n8588 , n25412 );
    xnor g16235 ( n22808 , n23418 , n17568 );
    xnor g16236 ( n30026 , n1905 , n11698 );
    and g16237 ( n18718 , n2437 , n27674 );
    or g16238 ( n33526 , n31110 , n14746 );
    not g16239 ( n16072 , n2615 );
    or g16240 ( n19811 , n14471 , n7349 );
    xnor g16241 ( n11215 , n26667 , n978 );
    or g16242 ( n26449 , n34421 , n17773 );
    xnor g16243 ( n5378 , n29080 , n27226 );
    and g16244 ( n19223 , n8076 , n25385 );
    and g16245 ( n18230 , n34881 , n22901 );
    xnor g16246 ( n29144 , n1466 , n10292 );
    or g16247 ( n21860 , n15702 , n35402 );
    and g16248 ( n13931 , n984 , n2381 );
    or g16249 ( n459 , n9607 , n20337 );
    xnor g16250 ( n11242 , n24933 , n26575 );
    or g16251 ( n10284 , n1897 , n5457 );
    or g16252 ( n33236 , n32934 , n5752 );
    or g16253 ( n24195 , n1673 , n24710 );
    and g16254 ( n22970 , n26791 , n32200 );
    or g16255 ( n4362 , n30199 , n29527 );
    or g16256 ( n21489 , n24968 , n763 );
    or g16257 ( n16764 , n18499 , n25298 );
    or g16258 ( n30524 , n16628 , n10762 );
    and g16259 ( n23300 , n16132 , n34940 );
    xnor g16260 ( n6074 , n29675 , n18547 );
    and g16261 ( n24176 , n31041 , n29186 );
    or g16262 ( n25768 , n11620 , n27821 );
    xnor g16263 ( n29665 , n12727 , n15464 );
    or g16264 ( n21885 , n11966 , n139 );
    buf g16265 ( n34600 , n30047 );
    or g16266 ( n23892 , n3921 , n8392 );
    or g16267 ( n20367 , n9060 , n5457 );
    or g16268 ( n31817 , n10894 , n25236 );
    or g16269 ( n23283 , n10052 , n20797 );
    or g16270 ( n27423 , n7835 , n11593 );
    or g16271 ( n15424 , n17568 , n7853 );
    and g16272 ( n29991 , n21831 , n24249 );
    or g16273 ( n33242 , n14098 , n2524 );
    xnor g16274 ( n23878 , n32220 , n15094 );
    or g16275 ( n11319 , n19098 , n35630 );
    or g16276 ( n17062 , n4745 , n25019 );
    xnor g16277 ( n19074 , n21618 , n671 );
    not g16278 ( n15904 , n19984 );
    or g16279 ( n638 , n2555 , n27704 );
    xnor g16280 ( n20452 , n28980 , n13118 );
    and g16281 ( n18144 , n31293 , n23520 );
    nor g16282 ( n23491 , n32584 , n32225 );
    or g16283 ( n392 , n6579 , n25306 );
    nor g16284 ( n35915 , n35927 , n1538 );
    or g16285 ( n599 , n21378 , n11996 );
    xnor g16286 ( n15340 , n28659 , n29884 );
    xnor g16287 ( n22918 , n11522 , n27878 );
    not g16288 ( n10358 , n10703 );
    buf g16289 ( n11312 , n9115 );
    xnor g16290 ( n13089 , n10317 , n19551 );
    xnor g16291 ( n10060 , n32525 , n18969 );
    or g16292 ( n32108 , n28565 , n20817 );
    or g16293 ( n17569 , n14959 , n19547 );
    or g16294 ( n15211 , n3205 , n4009 );
    nor g16295 ( n29705 , n19551 , n4598 );
    and g16296 ( n581 , n11260 , n31443 );
    or g16297 ( n13709 , n19984 , n8241 );
    or g16298 ( n12114 , n19750 , n29393 );
    or g16299 ( n27828 , n13726 , n4175 );
    and g16300 ( n12490 , n18889 , n33028 );
    or g16301 ( n29660 , n24371 , n23346 );
    xnor g16302 ( n12701 , n8767 , n10229 );
    or g16303 ( n32924 , n22988 , n2074 );
    and g16304 ( n10770 , n27055 , n30005 );
    nor g16305 ( n11464 , n32675 , n18566 );
    xnor g16306 ( n19203 , n31917 , n1368 );
    xnor g16307 ( n29173 , n34212 , n15676 );
    and g16308 ( n11985 , n35047 , n3734 );
    or g16309 ( n34803 , n3209 , n17964 );
    and g16310 ( n22736 , n2584 , n22212 );
    or g16311 ( n27035 , n22291 , n5523 );
    and g16312 ( n27611 , n4849 , n26289 );
    or g16313 ( n34886 , n2193 , n15496 );
    or g16314 ( n1483 , n14229 , n31261 );
    xnor g16315 ( n11438 , n25461 , n29252 );
    and g16316 ( n20022 , n23671 , n33478 );
    xnor g16317 ( n1106 , n32008 , n7720 );
    nor g16318 ( n23502 , n35927 , n4630 );
    buf g16319 ( n19173 , n23348 );
    or g16320 ( n2947 , n15313 , n22226 );
    or g16321 ( n15905 , n35927 , n18402 );
    xnor g16322 ( n15690 , n34313 , n4264 );
    or g16323 ( n718 , n35772 , n12950 );
    or g16324 ( n8104 , n7728 , n19671 );
    and g16325 ( n9136 , n13746 , n28817 );
    and g16326 ( n25730 , n24761 , n35066 );
    xnor g16327 ( n3957 , n20517 , n25174 );
    not g16328 ( n13436 , n23978 );
    and g16329 ( n32361 , n23839 , n33634 );
    xnor g16330 ( n11373 , n22437 , n22291 );
    xnor g16331 ( n15520 , n18339 , n26274 );
    not g16332 ( n34693 , n18572 );
    buf g16333 ( n31464 , n3842 );
    or g16334 ( n16088 , n9967 , n32608 );
    or g16335 ( n10495 , n31559 , n12480 );
    or g16336 ( n21836 , n25294 , n35402 );
    and g16337 ( n26077 , n27809 , n6403 );
    or g16338 ( n23899 , n13630 , n32329 );
    or g16339 ( n5579 , n28067 , n35043 );
    not g16340 ( n16803 , n16223 );
    xnor g16341 ( n7326 , n10858 , n18395 );
    or g16342 ( n18671 , n31056 , n16248 );
    xnor g16343 ( n4336 , n32083 , n29713 );
    or g16344 ( n21989 , n23374 , n22052 );
    or g16345 ( n359 , n22044 , n12465 );
    xnor g16346 ( n16694 , n28228 , n33039 );
    buf g16347 ( n17354 , n16728 );
    or g16348 ( n28621 , n11064 , n13307 );
    and g16349 ( n1459 , n32653 , n27366 );
    or g16350 ( n7 , n29839 , n27525 );
    or g16351 ( n30012 , n12656 , n25488 );
    xnor g16352 ( n28791 , n20470 , n33389 );
    and g16353 ( n30858 , n35685 , n6441 );
    nor g16354 ( n15195 , n14969 , n27785 );
    or g16355 ( n12081 , n1654 , n31055 );
    and g16356 ( n14481 , n2859 , n31152 );
    and g16357 ( n8932 , n15910 , n20609 );
    or g16358 ( n19719 , n21949 , n4128 );
    buf g16359 ( n11850 , n3805 );
    xnor g16360 ( n34759 , n7408 , n35457 );
    or g16361 ( n28204 , n18379 , n33284 );
    or g16362 ( n5054 , n9228 , n4530 );
    or g16363 ( n19101 , n15108 , n14637 );
    and g16364 ( n17458 , n1039 , n8532 );
    and g16365 ( n19118 , n11886 , n34768 );
    or g16366 ( n32300 , n3126 , n14554 );
    xnor g16367 ( n13600 , n32016 , n138 );
    xnor g16368 ( n20530 , n6200 , n7792 );
    not g16369 ( n15639 , n3360 );
    or g16370 ( n34572 , n2941 , n17399 );
    and g16371 ( n22994 , n29354 , n31845 );
    or g16372 ( n15583 , n28932 , n35296 );
    or g16373 ( n33801 , n7434 , n18312 );
    and g16374 ( n17902 , n24655 , n22536 );
    or g16375 ( n25380 , n7872 , n28895 );
    or g16376 ( n2069 , n11263 , n29581 );
    or g16377 ( n5203 , n32095 , n22765 );
    and g16378 ( n24381 , n3331 , n25457 );
    or g16379 ( n1305 , n20537 , n4580 );
    or g16380 ( n35236 , n1950 , n6127 );
    and g16381 ( n6991 , n28547 , n11726 );
    xnor g16382 ( n15853 , n10052 , n35800 );
    or g16383 ( n21435 , n25174 , n22080 );
    or g16384 ( n12208 , n35816 , n2124 );
    or g16385 ( n5130 , n9536 , n4184 );
    not g16386 ( n33199 , n18379 );
    and g16387 ( n1319 , n13749 , n19370 );
    or g16388 ( n4110 , n18797 , n12879 );
    xnor g16389 ( n9761 , n32544 , n5415 );
    xnor g16390 ( n12446 , n15949 , n32028 );
    xnor g16391 ( n35970 , n26561 , n30540 );
    or g16392 ( n4456 , n27683 , n26220 );
    nor g16393 ( n4028 , n31559 , n4753 );
    and g16394 ( n19982 , n23972 , n9980 );
    or g16395 ( n10109 , n21322 , n3716 );
    nor g16396 ( n8783 , n26759 , n33157 );
    xnor g16397 ( n2201 , n21759 , n19551 );
    not g16398 ( n34856 , n20925 );
    or g16399 ( n7818 , n30622 , n26292 );
    xnor g16400 ( n11150 , n3197 , n15766 );
    and g16401 ( n3141 , n22018 , n31526 );
    nor g16402 ( n29651 , n4288 , n21015 );
    xnor g16403 ( n23980 , n9321 , n21962 );
    or g16404 ( n11112 , n20597 , n15496 );
    xnor g16405 ( n18012 , n17355 , n5738 );
    and g16406 ( n16168 , n7189 , n35562 );
    not g16407 ( n10389 , n22882 );
    and g16408 ( n7436 , n18457 , n10797 );
    xnor g16409 ( n29600 , n2835 , n26347 );
    xnor g16410 ( n20256 , n13632 , n3205 );
    and g16411 ( n1970 , n15018 , n33626 );
    or g16412 ( n29609 , n4971 , n15195 );
    and g16413 ( n19953 , n167 , n11222 );
    or g16414 ( n14960 , n30954 , n3431 );
    or g16415 ( n5933 , n30974 , n22002 );
    and g16416 ( n12331 , n12027 , n31759 );
    and g16417 ( n11745 , n18771 , n15762 );
    or g16418 ( n13750 , n6430 , n15788 );
    and g16419 ( n19896 , n35403 , n8394 );
    xnor g16420 ( n19500 , n26068 , n35238 );
    xnor g16421 ( n28517 , n18258 , n3946 );
    or g16422 ( n17817 , n34547 , n30287 );
    nor g16423 ( n4838 , n24720 , n22165 );
    or g16424 ( n8676 , n10320 , n33310 );
    xnor g16425 ( n6119 , n17451 , n8432 );
    and g16426 ( n32253 , n392 , n26167 );
    or g16427 ( n29798 , n27438 , n30826 );
    and g16428 ( n29929 , n23578 , n795 );
    nor g16429 ( n27163 , n5015 , n18115 );
    and g16430 ( n20474 , n2336 , n12531 );
    and g16431 ( n27821 , n33106 , n11094 );
    or g16432 ( n24049 , n23636 , n2880 );
    or g16433 ( n11105 , n25602 , n4316 );
    not g16434 ( n10374 , n27595 );
    and g16435 ( n5112 , n31144 , n34930 );
    or g16436 ( n21445 , n4962 , n34081 );
    xnor g16437 ( n8672 , n541 , n11753 );
    or g16438 ( n22465 , n21941 , n2366 );
    or g16439 ( n33634 , n23843 , n35935 );
    or g16440 ( n19911 , n28401 , n22783 );
    xnor g16441 ( n20715 , n13667 , n20197 );
    xnor g16442 ( n739 , n19426 , n18237 );
    not g16443 ( n31395 , n6226 );
    nor g16444 ( n12901 , n28864 , n8319 );
    xnor g16445 ( n26744 , n15660 , n1078 );
    xnor g16446 ( n7594 , n9309 , n32584 );
    and g16447 ( n35708 , n22836 , n12350 );
    or g16448 ( n13507 , n35907 , n6683 );
    or g16449 ( n17124 , n15341 , n17233 );
    not g16450 ( n2535 , n3480 );
    or g16451 ( n14130 , n4079 , n24672 );
    or g16452 ( n19689 , n3055 , n19636 );
    or g16453 ( n15481 , n18631 , n21579 );
    nor g16454 ( n35934 , n13558 , n415 );
    or g16455 ( n6411 , n32722 , n7071 );
    and g16456 ( n32621 , n12905 , n2121 );
    nor g16457 ( n31249 , n34253 , n13455 );
    or g16458 ( n26518 , n11608 , n8153 );
    nor g16459 ( n5183 , n10091 , n23112 );
    xnor g16460 ( n30527 , n11534 , n7755 );
    xnor g16461 ( n19186 , n19930 , n5335 );
    and g16462 ( n24624 , n13605 , n23354 );
    and g16463 ( n22173 , n31952 , n13030 );
    or g16464 ( n10909 , n11647 , n26220 );
    or g16465 ( n13883 , n13144 , n26468 );
    or g16466 ( n27781 , n7542 , n8134 );
    or g16467 ( n12728 , n32584 , n13702 );
    or g16468 ( n12198 , n17608 , n34297 );
    or g16469 ( n10421 , n11190 , n208 );
    and g16470 ( n26526 , n30162 , n35963 );
    xnor g16471 ( n29764 , n20643 , n33476 );
    and g16472 ( n32049 , n32737 , n33506 );
    not g16473 ( n8231 , n7268 );
    or g16474 ( n1488 , n24046 , n32003 );
    or g16475 ( n21992 , n32925 , n27704 );
    and g16476 ( n19652 , n30082 , n26300 );
    or g16477 ( n4686 , n24971 , n28404 );
    and g16478 ( n22932 , n33749 , n15635 );
    xnor g16479 ( n27345 , n20448 , n2085 );
    not g16480 ( n35312 , n22980 );
    or g16481 ( n17778 , n6182 , n34997 );
    or g16482 ( n16442 , n4878 , n11808 );
    xnor g16483 ( n23867 , n9819 , n35927 );
    or g16484 ( n10830 , n17984 , n28064 );
    or g16485 ( n20691 , n8401 , n10960 );
    and g16486 ( n12457 , n5599 , n31540 );
    xnor g16487 ( n12096 , n33525 , n8305 );
    or g16488 ( n5854 , n5644 , n34865 );
    or g16489 ( n15522 , n17470 , n12035 );
    and g16490 ( n23327 , n10837 , n5177 );
    or g16491 ( n6190 , n5195 , n4751 );
    or g16492 ( n26454 , n16215 , n24856 );
    or g16493 ( n6679 , n13907 , n26468 );
    or g16494 ( n35874 , n3380 , n14361 );
    or g16495 ( n586 , n1803 , n14554 );
    and g16496 ( n30559 , n30628 , n14560 );
    nor g16497 ( n29932 , n30901 , n26189 );
    or g16498 ( n30731 , n14975 , n14076 );
    and g16499 ( n14626 , n25040 , n5203 );
    xnor g16500 ( n26731 , n29137 , n10894 );
    or g16501 ( n23893 , n25174 , n25013 );
    or g16502 ( n18311 , n35042 , n22316 );
    xnor g16503 ( n10635 , n15495 , n35927 );
    and g16504 ( n424 , n257 , n9188 );
    or g16505 ( n18735 , n10894 , n7646 );
    xnor g16506 ( n5262 , n24116 , n23692 );
    or g16507 ( n19703 , n18365 , n24672 );
    or g16508 ( n18880 , n2334 , n24517 );
    and g16509 ( n14434 , n33653 , n31161 );
    nor g16510 ( n23896 , n25711 , n30158 );
    nor g16511 ( n13466 , n4553 , n31388 );
    not g16512 ( n29224 , n9789 );
    xnor g16513 ( n9320 , n1134 , n269 );
    or g16514 ( n8854 , n22675 , n2039 );
    and g16515 ( n28693 , n6810 , n21901 );
    or g16516 ( n26994 , n25174 , n19478 );
    not g16517 ( n10783 , n7867 );
    and g16518 ( n10889 , n20999 , n9294 );
    and g16519 ( n2992 , n29781 , n31673 );
    or g16520 ( n4486 , n17261 , n4421 );
    and g16521 ( n11406 , n33062 , n20217 );
    and g16522 ( n15728 , n28625 , n26955 );
    or g16523 ( n31473 , n17336 , n10176 );
    not g16524 ( n24899 , n10273 );
    xnor g16525 ( n18763 , n15313 , n22226 );
    or g16526 ( n22389 , n9658 , n15317 );
    and g16527 ( n647 , n8082 , n34058 );
    xnor g16528 ( n16822 , n5483 , n20661 );
    or g16529 ( n25288 , n29949 , n2117 );
    xnor g16530 ( n23723 , n34622 , n5335 );
    and g16531 ( n1723 , n27197 , n33366 );
    nor g16532 ( n5653 , n15403 , n32449 );
    xnor g16533 ( n23024 , n13027 , n16620 );
    or g16534 ( n5898 , n8432 , n28479 );
    xnor g16535 ( n32421 , n22766 , n30703 );
    or g16536 ( n27798 , n23604 , n14136 );
    xnor g16537 ( n23311 , n130 , n10894 );
    or g16538 ( n33760 , n5052 , n19421 );
    or g16539 ( n18146 , n10064 , n16457 );
    buf g16540 ( n4478 , n18721 );
    or g16541 ( n8032 , n8563 , n28455 );
    and g16542 ( n4719 , n1415 , n9754 );
    and g16543 ( n5337 , n30340 , n25487 );
    or g16544 ( n33619 , n30066 , n5868 );
    or g16545 ( n17207 , n14043 , n14918 );
    or g16546 ( n15218 , n11046 , n33376 );
    nor g16547 ( n8078 , n3946 , n8486 );
    and g16548 ( n31538 , n700 , n13980 );
    xnor g16549 ( n23813 , n9002 , n12255 );
    or g16550 ( n21467 , n15464 , n35717 );
    xnor g16551 ( n18743 , n28529 , n28000 );
    or g16552 ( n1705 , n23540 , n22783 );
    or g16553 ( n1771 , n17568 , n17265 );
    nor g16554 ( n16946 , n1950 , n2037 );
    or g16555 ( n5815 , n253 , n20601 );
    or g16556 ( n15586 , n25174 , n34447 );
    and g16557 ( n35553 , n20342 , n27928 );
    xnor g16558 ( n9763 , n6344 , n19033 );
    xnor g16559 ( n19692 , n17889 , n23033 );
    or g16560 ( n30081 , n31799 , n31861 );
    xnor g16561 ( n7091 , n32224 , n4960 );
    or g16562 ( n3482 , n17151 , n9601 );
    or g16563 ( n4543 , n34927 , n17111 );
    or g16564 ( n16260 , n22054 , n14841 );
    and g16565 ( n3174 , n30579 , n32807 );
    or g16566 ( n13938 , n21520 , n12294 );
    not g16567 ( n25861 , n2928 );
    or g16568 ( n7308 , n22197 , n1783 );
    or g16569 ( n25574 , n28810 , n23790 );
    and g16570 ( n17603 , n28197 , n4205 );
    or g16571 ( n16292 , n7975 , n18482 );
    and g16572 ( n30674 , n5311 , n32761 );
    or g16573 ( n8884 , n26461 , n11497 );
    and g16574 ( n11426 , n31418 , n35192 );
    and g16575 ( n11357 , n19685 , n27597 );
    or g16576 ( n3204 , n24371 , n3389 );
    and g16577 ( n27295 , n16476 , n3879 );
    or g16578 ( n28450 , n19537 , n25392 );
    or g16579 ( n16870 , n32143 , n17162 );
    xnor g16580 ( n11797 , n17754 , n31056 );
    or g16581 ( n1891 , n10039 , n25302 );
    xnor g16582 ( n14574 , n36006 , n24756 );
    nor g16583 ( n11495 , n28742 , n12824 );
    xnor g16584 ( n4592 , n1658 , n19876 );
    or g16585 ( n11116 , n23761 , n18542 );
    or g16586 ( n6716 , n35927 , n31819 );
    and g16587 ( n3992 , n2025 , n21414 );
    or g16588 ( n9922 , n18501 , n2798 );
    xnor g16589 ( n21711 , n1488 , n3946 );
    not g16590 ( n6401 , n1078 );
    or g16591 ( n29723 , n15115 , n585 );
    xnor g16592 ( n33058 , n1412 , n19593 );
    or g16593 ( n2210 , n8706 , n2746 );
    xnor g16594 ( n35362 , n25149 , n25958 );
    and g16595 ( n21436 , n13669 , n18422 );
    or g16596 ( n21559 , n26978 , n33261 );
    and g16597 ( n20760 , n2723 , n28876 );
    xnor g16598 ( n24064 , n21877 , n26196 );
    xnor g16599 ( n33488 , n6780 , n35927 );
    not g16600 ( n9268 , n35453 );
    or g16601 ( n13422 , n4011 , n20082 );
    xor g16602 ( n11344 , n35379 , n24768 );
    xnor g16603 ( n21075 , n16857 , n13872 );
    xnor g16604 ( n16565 , n7418 , n25209 );
    or g16605 ( n5681 , n17395 , n16457 );
    or g16606 ( n21670 , n9690 , n11712 );
    or g16607 ( n7628 , n21660 , n29310 );
    or g16608 ( n35116 , n32857 , n35241 );
    or g16609 ( n30918 , n11630 , n12089 );
    or g16610 ( n31561 , n32715 , n18037 );
    xnor g16611 ( n25968 , n28472 , n22291 );
    or g16612 ( n12992 , n10845 , n21220 );
    and g16613 ( n6529 , n29931 , n24189 );
    xnor g16614 ( n33369 , n30852 , n22291 );
    or g16615 ( n2159 , n2019 , n12913 );
    nor g16616 ( n2578 , n26199 , n25962 );
    or g16617 ( n14427 , n34170 , n17845 );
    or g16618 ( n21088 , n10524 , n23836 );
    or g16619 ( n32845 , n7213 , n27963 );
    or g16620 ( n11305 , n33582 , n35644 );
    and g16621 ( n33245 , n9678 , n35919 );
    nor g16622 ( n27065 , n10894 , n4918 );
    xnor g16623 ( n25233 , n18941 , n25458 );
    xnor g16624 ( n30724 , n2909 , n22670 );
    xnor g16625 ( n18516 , n7634 , n23809 );
    or g16626 ( n28015 , n29350 , n3513 );
    and g16627 ( n15138 , n13370 , n25258 );
    buf g16628 ( n18477 , n22870 );
    not g16629 ( n11315 , n9924 );
    and g16630 ( n4627 , n5271 , n430 );
    xnor g16631 ( n31777 , n21214 , n17598 );
    or g16632 ( n563 , n4196 , n24333 );
    xnor g16633 ( n2175 , n25192 , n35595 );
    nor g16634 ( n5220 , n5727 , n30978 );
    and g16635 ( n11589 , n6154 , n29660 );
    and g16636 ( n6560 , n6695 , n14352 );
    and g16637 ( n32982 , n34115 , n17504 );
    or g16638 ( n30347 , n34441 , n31055 );
    or g16639 ( n22288 , n27441 , n17046 );
    nor g16640 ( n23130 , n10812 , n35407 );
    or g16641 ( n23506 , n31215 , n30217 );
    not g16642 ( n18088 , n15344 );
    or g16643 ( n23162 , n26622 , n15290 );
    and g16644 ( n20193 , n7395 , n1038 );
    or g16645 ( n3012 , n25367 , n17259 );
    or g16646 ( n2205 , n16620 , n4787 );
    xnor g16647 ( n32368 , n30591 , n31559 );
    and g16648 ( n11536 , n1910 , n34770 );
    xnor g16649 ( n25801 , n26665 , n28657 );
    nor g16650 ( n14115 , n4878 , n13955 );
    or g16651 ( n29906 , n5067 , n35556 );
    xnor g16652 ( n35443 , n19462 , n13113 );
    and g16653 ( n10792 , n6833 , n29399 );
    buf g16654 ( n32329 , n790 );
    or g16655 ( n30919 , n20357 , n1402 );
    or g16656 ( n11290 , n19551 , n16585 );
    or g16657 ( n11923 , n3942 , n3736 );
    or g16658 ( n6307 , n6505 , n3188 );
    xnor g16659 ( n16341 , n4268 , n3006 );
    and g16660 ( n3016 , n1035 , n30176 );
    xnor g16661 ( n4921 , n35308 , n35622 );
    or g16662 ( n18646 , n11190 , n29881 );
    and g16663 ( n15495 , n6620 , n25309 );
    or g16664 ( n23949 , n19551 , n11743 );
    or g16665 ( n23248 , n23297 , n14369 );
    nor g16666 ( n32678 , n89 , n16516 );
    or g16667 ( n18816 , n15270 , n8924 );
    or g16668 ( n33145 , n3946 , n26100 );
    or g16669 ( n3260 , n8432 , n7921 );
    not g16670 ( n30700 , n2433 );
    or g16671 ( n8339 , n7789 , n12197 );
    or g16672 ( n32974 , n32095 , n14683 );
    xnor g16673 ( n16670 , n4472 , n9802 );
    or g16674 ( n26040 , n28114 , n24489 );
    or g16675 ( n31344 , n11757 , n6919 );
    and g16676 ( n21837 , n18547 , n29675 );
    or g16677 ( n19445 , n3788 , n27944 );
    and g16678 ( n30677 , n10004 , n12842 );
    and g16679 ( n30125 , n2885 , n6028 );
    nor g16680 ( n11784 , n16620 , n26237 );
    xnor g16681 ( n16514 , n17412 , n22841 );
    or g16682 ( n32045 , n21729 , n3239 );
    nor g16683 ( n33486 , n719 , n23921 );
    and g16684 ( n31457 , n24340 , n16557 );
    xnor g16685 ( n28818 , n18750 , n17742 );
    or g16686 ( n3851 , n11438 , n31464 );
    or g16687 ( n25387 , n1686 , n6302 );
    or g16688 ( n10467 , n7937 , n20601 );
    nor g16689 ( n4564 , n34178 , n30558 );
    xnor g16690 ( n13657 , n7801 , n8501 );
    xnor g16691 ( n25495 , n13277 , n25061 );
    or g16692 ( n11220 , n4758 , n15263 );
    or g16693 ( n35904 , n13820 , n11680 );
    xnor g16694 ( n14380 , n14753 , n21685 );
    or g16695 ( n14094 , n32492 , n34214 );
    xnor g16696 ( n22645 , n14366 , n8432 );
    xnor g16697 ( n11965 , n33321 , n20380 );
    xnor g16698 ( n33631 , n20646 , n12055 );
    not g16699 ( n14998 , n20963 );
    or g16700 ( n5468 , n22381 , n9915 );
    and g16701 ( n557 , n25691 , n4371 );
    or g16702 ( n16661 , n24371 , n10485 );
    xnor g16703 ( n28199 , n8344 , n24371 );
    nor g16704 ( n14986 , n10894 , n11355 );
    and g16705 ( n2144 , n30850 , n26309 );
    not g16706 ( n23650 , n24260 );
    and g16707 ( n26195 , n33134 , n33180 );
    buf g16708 ( n19732 , n9030 );
    and g16709 ( n30575 , n28478 , n16380 );
    and g16710 ( n34717 , n20100 , n27516 );
    or g16711 ( n19592 , n12749 , n5450 );
    xnor g16712 ( n30565 , n15148 , n5795 );
    xnor g16713 ( n1999 , n35606 , n333 );
    xnor g16714 ( n31761 , n6681 , n9121 );
    xnor g16715 ( n32136 , n23014 , n35433 );
    or g16716 ( n3718 , n23487 , n32379 );
    xnor g16717 ( n35939 , n30070 , n5137 );
    xnor g16718 ( n3766 , n28920 , n1730 );
    and g16719 ( n10911 , n3665 , n9011 );
    xnor g16720 ( n10210 , n13270 , n15886 );
    or g16721 ( n25872 , n22686 , n35143 );
    or g16722 ( n31441 , n30557 , n10166 );
    or g16723 ( n8504 , n3947 , n12622 );
    or g16724 ( n5084 , n35881 , n5779 );
    or g16725 ( n32610 , n8489 , n11312 );
    or g16726 ( n4299 , n34519 , n14841 );
    and g16727 ( n26503 , n5128 , n20114 );
    xnor g16728 ( n27377 , n9980 , n22394 );
    and g16729 ( n9989 , n22728 , n23620 );
    nor g16730 ( n19131 , n24032 , n35659 );
    nor g16731 ( n35390 , n8432 , n34796 );
    or g16732 ( n11167 , n34509 , n17346 );
    or g16733 ( n13448 , n29784 , n22961 );
    and g16734 ( n23764 , n11316 , n10870 );
    xor g16735 ( n33663 , n23638 , n17852 );
    or g16736 ( n20914 , n32857 , n5478 );
    or g16737 ( n1895 , n16620 , n14816 );
    xnor g16738 ( n1221 , n16798 , n19919 );
    and g16739 ( n14723 , n29537 , n24945 );
    or g16740 ( n3646 , n32315 , n11996 );
    or g16741 ( n8996 , n11609 , n30826 );
    or g16742 ( n466 , n35286 , n25592 );
    or g16743 ( n6164 , n8616 , n4175 );
    or g16744 ( n36028 , n17663 , n28668 );
    or g16745 ( n20362 , n11744 , n122 );
    nor g16746 ( n10586 , n830 , n29499 );
    or g16747 ( n17809 , n32715 , n30144 );
    xnor g16748 ( n24630 , n32293 , n19551 );
    xnor g16749 ( n22837 , n9373 , n32095 );
    xnor g16750 ( n10786 , n35985 , n29713 );
    and g16751 ( n5111 , n14534 , n15907 );
    or g16752 ( n9582 , n8514 , n28866 );
    xnor g16753 ( n22817 , n21269 , n29839 );
    or g16754 ( n16958 , n32095 , n23579 );
    or g16755 ( n11512 , n22571 , n2384 );
    and g16756 ( n29565 , n34933 , n8681 );
    or g16757 ( n19882 , n10998 , n26864 );
    or g16758 ( n10787 , n17721 , n9995 );
    and g16759 ( n11760 , n17813 , n23003 );
    or g16760 ( n2673 , n4960 , n3223 );
    or g16761 ( n15395 , n12588 , n27973 );
    or g16762 ( n20436 , n35927 , n7998 );
    nor g16763 ( n35454 , n11455 , n30559 );
    and g16764 ( n12908 , n30903 , n28090 );
    xnor g16765 ( n9290 , n18504 , n8531 );
    or g16766 ( n4660 , n9793 , n1757 );
    and g16767 ( n24550 , n5811 , n200 );
    and g16768 ( n27171 , n2149 , n30956 );
    or g16769 ( n24800 , n9789 , n8167 );
    or g16770 ( n12814 , n5335 , n4308 );
    xnor g16771 ( n164 , n10486 , n24112 );
    nor g16772 ( n32337 , n29713 , n12640 );
    not g16773 ( n25110 , n22048 );
    or g16774 ( n28478 , n28462 , n11848 );
    nor g16775 ( n13328 , n26761 , n1603 );
    and g16776 ( n32801 , n28578 , n3760 );
    not g16777 ( n11379 , n33244 );
    and g16778 ( n32909 , n32626 , n9527 );
    or g16779 ( n33877 , n24371 , n8286 );
    or g16780 ( n8560 , n29713 , n34815 );
    not g16781 ( n20696 , n16030 );
    nor g16782 ( n32126 , n305 , n31055 );
    and g16783 ( n2927 , n14884 , n10421 );
    xnor g16784 ( n35645 , n5163 , n27226 );
    or g16785 ( n32650 , n2230 , n9832 );
    or g16786 ( n15579 , n16922 , n18297 );
    xnor g16787 ( n16046 , n15480 , n4742 );
    or g16788 ( n27846 , n550 , n5252 );
    or g16789 ( n16588 , n4878 , n396 );
    or g16790 ( n9415 , n29713 , n22514 );
    or g16791 ( n10056 , n25174 , n418 );
    or g16792 ( n21558 , n4647 , n26002 );
    or g16793 ( n3248 , n5410 , n8153 );
    or g16794 ( n6387 , n830 , n27822 );
    xnor g16795 ( n24573 , n3972 , n17133 );
    or g16796 ( n28311 , n8275 , n2802 );
    and g16797 ( n35304 , n2440 , n26330 );
    xnor g16798 ( n3541 , n33070 , n11640 );
    or g16799 ( n35734 , n33049 , n10634 );
    not g16800 ( n28746 , n32574 );
    and g16801 ( n30425 , n5016 , n432 );
    or g16802 ( n14451 , n32192 , n20 );
    or g16803 ( n16878 , n3295 , n21956 );
    or g16804 ( n9438 , n14855 , n25786 );
    or g16805 ( n17462 , n8621 , n30683 );
    or g16806 ( n12559 , n25422 , n29626 );
    and g16807 ( n34002 , n4672 , n21929 );
    xnor g16808 ( n10992 , n9980 , n26245 );
    and g16809 ( n25690 , n28597 , n3908 );
    xnor g16810 ( n14693 , n31861 , n31799 );
    or g16811 ( n4347 , n21079 , n30205 );
    not g16812 ( n35030 , n18012 );
    xor g16813 ( n5312 , n22009 , n25326 );
    not g16814 ( n3662 , n1007 );
    or g16815 ( n25996 , n208 , n27053 );
    or g16816 ( n27064 , n1932 , n15274 );
    or g16817 ( n21375 , n26004 , n20762 );
    not g16818 ( n3981 , n1494 );
    or g16819 ( n18226 , n4679 , n31773 );
    xnor g16820 ( n2314 , n29034 , n21477 );
    not g16821 ( n16667 , n20171 );
    or g16822 ( n18390 , n34985 , n24710 );
    and g16823 ( n22292 , n35752 , n24417 );
    xnor g16824 ( n8705 , n12669 , n31215 );
    xnor g16825 ( n22650 , n20465 , n21651 );
    or g16826 ( n10220 , n32050 , n34656 );
    not g16827 ( n9055 , n29954 );
    or g16828 ( n7334 , n29979 , n8580 );
    or g16829 ( n32292 , n32546 , n22322 );
    xnor g16830 ( n11454 , n20213 , n32857 );
    and g16831 ( n26515 , n22768 , n22005 );
    or g16832 ( n30261 , n31559 , n33803 );
    or g16833 ( n27836 , n3205 , n11644 );
    xnor g16834 ( n18064 , n14566 , n4960 );
    or g16835 ( n11158 , n15442 , n2798 );
    or g16836 ( n35966 , n2345 , n27181 );
    or g16837 ( n15880 , n23604 , n24243 );
    and g16838 ( n26018 , n18602 , n35331 );
    and g16839 ( n32774 , n3462 , n20693 );
    and g16840 ( n32919 , n12607 , n34143 );
    xnor g16841 ( n107 , n8540 , n27295 );
    or g16842 ( n7186 , n33288 , n578 );
    or g16843 ( n6418 , n17500 , n22858 );
    or g16844 ( n25359 , n32272 , n19421 );
    not g16845 ( n7590 , n23407 );
    and g16846 ( n25863 , n8114 , n20420 );
    and g16847 ( n1440 , n21109 , n24495 );
    or g16848 ( n32948 , n18983 , n3989 );
    or g16849 ( n23436 , n9658 , n33185 );
    xnor g16850 ( n7819 , n9611 , n30621 );
    or g16851 ( n9925 , n4878 , n36046 );
    and g16852 ( n21926 , n31338 , n12410 );
    or g16853 ( n21025 , n604 , n6950 );
    or g16854 ( n31959 , n27767 , n17068 );
    xnor g16855 ( n17222 , n32707 , n18873 );
    nor g16856 ( n6777 , n16620 , n10294 );
    or g16857 ( n22295 , n18772 , n7457 );
    and g16858 ( n15194 , n9044 , n4150 );
    not g16859 ( n35182 , n16480 );
    or g16860 ( n13125 , n25174 , n20712 );
    and g16861 ( n771 , n20831 , n31655 );
    or g16862 ( n20663 , n30742 , n24900 );
    xnor g16863 ( n1364 , n24545 , n9658 );
    or g16864 ( n10251 , n12076 , n20427 );
    not g16865 ( n24283 , n21012 );
    or g16866 ( n24705 , n7036 , n32507 );
    buf g16867 ( n35757 , n25369 );
    and g16868 ( n35317 , n17733 , n11063 );
    or g16869 ( n694 , n21167 , n4467 );
    or g16870 ( n4106 , n4878 , n20050 );
    and g16871 ( n29379 , n20791 , n7530 );
    not g16872 ( n29205 , n32095 );
    or g16873 ( n7805 , n21228 , n27740 );
    or g16874 ( n9695 , n4962 , n14481 );
    and g16875 ( n26697 , n35918 , n22895 );
    and g16876 ( n23080 , n21963 , n22216 );
    not g16877 ( n22958 , n30848 );
    not g16878 ( n34433 , n26840 );
    or g16879 ( n13365 , n4878 , n26125 );
    or g16880 ( n919 , n32529 , n4318 );
    not g16881 ( n5167 , n22009 );
    or g16882 ( n34105 , n20488 , n22858 );
    and g16883 ( n27462 , n17882 , n28838 );
    nor g16884 ( n20841 , n17568 , n4017 );
    or g16885 ( n35289 , n4960 , n4201 );
    and g16886 ( n1660 , n11491 , n21841 );
    xnor g16887 ( n5880 , n4310 , n23825 );
    or g16888 ( n12109 , n2258 , n3199 );
    xnor g16889 ( n26383 , n7470 , n20957 );
    xnor g16890 ( n14594 , n23384 , n23338 );
    and g16891 ( n8018 , n3692 , n34677 );
    and g16892 ( n27362 , n12954 , n19569 );
    and g16893 ( n29106 , n19766 , n29035 );
    and g16894 ( n33468 , n12295 , n12038 );
    xnor g16895 ( n7573 , n23118 , n10894 );
    xnor g16896 ( n20786 , n21190 , n5327 );
    xnor g16897 ( n17349 , n26915 , n830 );
    xnor g16898 ( n22211 , n33598 , n6258 );
    or g16899 ( n24409 , n5335 , n29508 );
    xnor g16900 ( n14528 , n28242 , n7540 );
    or g16901 ( n5229 , n31799 , n7003 );
    nor g16902 ( n6940 , n18137 , n15414 );
    or g16903 ( n23728 , n33027 , n24124 );
    or g16904 ( n34526 , n19972 , n9896 );
    and g16905 ( n21022 , n15902 , n1286 );
    or g16906 ( n10619 , n25476 , n4260 );
    or g16907 ( n21203 , n11730 , n2077 );
    not g16908 ( n12533 , n4477 );
    not g16909 ( n23798 , n9739 );
    or g16910 ( n15516 , n31056 , n13528 );
    not g16911 ( n12869 , n3239 );
    xnor g16912 ( n14438 , n20881 , n3346 );
    or g16913 ( n26097 , n730 , n23689 );
    or g16914 ( n30783 , n18549 , n17964 );
    or g16915 ( n1147 , n34068 , n6075 );
    nor g16916 ( n11731 , n17478 , n16007 );
    or g16917 ( n30846 , n20099 , n17354 );
    xnor g16918 ( n28098 , n6225 , n32982 );
    nor g16919 ( n20125 , n32857 , n1413 );
    not g16920 ( n13002 , n2886 );
    not g16921 ( n9058 , n20295 );
    or g16922 ( n3460 , n6504 , n7417 );
    not g16923 ( n13613 , n16069 );
    or g16924 ( n8079 , n17451 , n32821 );
    nor g16925 ( n8770 , n17568 , n18427 );
    not g16926 ( n17363 , n35523 );
    not g16927 ( n30406 , n3805 );
    not g16928 ( n3112 , n22197 );
    or g16929 ( n16109 , n4288 , n21129 );
    and g16930 ( n14885 , n1608 , n6639 );
    xnor g16931 ( n35398 , n25318 , n27291 );
    not g16932 ( n14218 , n10336 );
    or g16933 ( n12745 , n3160 , n22783 );
    xnor g16934 ( n32729 , n4030 , n33494 );
    and g16935 ( n18739 , n35409 , n15153 );
    or g16936 ( n14204 , n28795 , n32808 );
    xnor g16937 ( n9891 , n13805 , n11455 );
    not g16938 ( n33783 , n27429 );
    xnor g16939 ( n1657 , n17415 , n11046 );
    and g16940 ( n8075 , n19264 , n26996 );
    nor g16941 ( n33831 , n23337 , n25762 );
    or g16942 ( n2743 , n8454 , n4359 );
    or g16943 ( n32435 , n13420 , n3219 );
    and g16944 ( n19576 , n19157 , n12723 );
    nor g16945 ( n19776 , n31659 , n13777 );
    and g16946 ( n28564 , n30673 , n15072 );
    nor g16947 ( n26591 , n17182 , n31411 );
    or g16948 ( n2542 , n32229 , n17962 );
    and g16949 ( n25543 , n23525 , n13195 );
    and g16950 ( n13082 , n19616 , n5097 );
    and g16951 ( n2134 , n2736 , n386 );
    or g16952 ( n35945 , n19269 , n28837 );
    and g16953 ( n10311 , n21920 , n21013 );
    and g16954 ( n12727 , n32850 , n2196 );
    xnor g16955 ( n11313 , n15308 , n19551 );
    and g16956 ( n34648 , n2163 , n2205 );
    or g16957 ( n5774 , n32095 , n7888 );
    or g16958 ( n22151 , n10146 , n31055 );
    xnor g16959 ( n2397 , n9536 , n4184 );
    or g16960 ( n18704 , n32095 , n34955 );
    or g16961 ( n13399 , n33280 , n16876 );
    or g16962 ( n19501 , n7022 , n35402 );
    or g16963 ( n17824 , n4878 , n31363 );
    or g16964 ( n33516 , n14439 , n32093 );
    or g16965 ( n20761 , n7881 , n25392 );
    and g16966 ( n5593 , n11554 , n12898 );
    not g16967 ( n11309 , n24332 );
    xnor g16968 ( n36006 , n30282 , n7540 );
    xnor g16969 ( n10261 , n12507 , n18397 );
    xnor g16970 ( n33038 , n21492 , n33748 );
    and g16971 ( n25154 , n13806 , n13004 );
    or g16972 ( n32423 , n13728 , n17042 );
    buf g16973 ( n23462 , n29872 );
    xnor g16974 ( n28979 , n2217 , n31753 );
    not g16975 ( n20525 , n18404 );
    or g16976 ( n33072 , n31799 , n33569 );
    xnor g16977 ( n2103 , n16991 , n10770 );
    or g16978 ( n7076 , n11455 , n2429 );
    or g16979 ( n24644 , n9793 , n17244 );
    xnor g16980 ( n14547 , n13562 , n4288 );
    or g16981 ( n27139 , n1993 , n10730 );
    not g16982 ( n32881 , n467 );
    xnor g16983 ( n14934 , n7618 , n31700 );
    or g16984 ( n3710 , n12384 , n25051 );
    xnor g16985 ( n30251 , n29574 , n13568 );
    not g16986 ( n23378 , n7588 );
    nor g16987 ( n31004 , n4498 , n26439 );
    and g16988 ( n32725 , n35599 , n847 );
    or g16989 ( n19527 , n24950 , n23626 );
    buf g16990 ( n28438 , n3798 );
    or g16991 ( n33883 , n8552 , n20308 );
    xnor g16992 ( n20794 , n19656 , n5335 );
    xnor g16993 ( n24272 , n2539 , n18379 );
    not g16994 ( n2570 , n546 );
    or g16995 ( n35087 , n13662 , n18388 );
    and g16996 ( n32856 , n6130 , n10442 );
    and g16997 ( n4023 , n24502 , n20577 );
    not g16998 ( n15731 , n1072 );
    or g16999 ( n18315 , n9682 , n31067 );
    or g17000 ( n9276 , n28208 , n19058 );
    or g17001 ( n10120 , n3467 , n26514 );
    or g17002 ( n11602 , n7865 , n1892 );
    or g17003 ( n28152 , n24371 , n34938 );
    or g17004 ( n35670 , n5287 , n13603 );
    or g17005 ( n10778 , n23718 , n26480 );
    nor g17006 ( n29000 , n8432 , n3009 );
    xnor g17007 ( n14969 , n10545 , n15464 );
    or g17008 ( n35149 , n18273 , n6288 );
    xnor g17009 ( n21528 , n21272 , n5215 );
    or g17010 ( n251 , n1950 , n11590 );
    xnor g17011 ( n12832 , n15040 , n5335 );
    not g17012 ( n14040 , n27226 );
    and g17013 ( n5747 , n25146 , n25798 );
    or g17014 ( n30390 , n830 , n35318 );
    xnor g17015 ( n26217 , n11839 , n26246 );
    xnor g17016 ( n26587 , n1174 , n4288 );
    or g17017 ( n25634 , n34081 , n33761 );
    buf g17018 ( n19058 , n13084 );
    xnor g17019 ( n11369 , n5493 , n19730 );
    not g17020 ( n16421 , n12054 );
    xnor g17021 ( n12506 , n31450 , n26964 );
    or g17022 ( n25751 , n15869 , n11716 );
    xnor g17023 ( n20264 , n33413 , n32584 );
    not g17024 ( n34656 , n30947 );
    not g17025 ( n11104 , n16223 );
    xnor g17026 ( n18492 , n649 , n31552 );
    xnor g17027 ( n3180 , n2066 , n28868 );
    and g17028 ( n14725 , n3519 , n27134 );
    or g17029 ( n28147 , n14071 , n8295 );
    nor g17030 ( n5028 , n31559 , n13861 );
    and g17031 ( n4852 , n28213 , n24962 );
    or g17032 ( n3038 , n31289 , n22944 );
    or g17033 ( n14219 , n12408 , n8607 );
    or g17034 ( n26764 , n22291 , n15170 );
    or g17035 ( n2599 , n24111 , n34084 );
    or g17036 ( n27468 , n14156 , n16919 );
    or g17037 ( n5281 , n8650 , n13664 );
    nor g17038 ( n22612 , n31799 , n242 );
    and g17039 ( n22784 , n27828 , n18105 );
    or g17040 ( n20306 , n5092 , n26931 );
    xnor g17041 ( n15692 , n22286 , n20033 );
    or g17042 ( n23794 , n34555 , n1511 );
    xnor g17043 ( n24134 , n30142 , n25489 );
    or g17044 ( n27414 , n23800 , n20637 );
    and g17045 ( n3426 , n15280 , n28369 );
    xnor g17046 ( n31223 , n22590 , n25456 );
    and g17047 ( n8271 , n26575 , n24933 );
    xnor g17048 ( n10088 , n2516 , n17726 );
    or g17049 ( n29191 , n27226 , n32407 );
    and g17050 ( n24254 , n33756 , n11733 );
    or g17051 ( n29207 , n29573 , n18316 );
    or g17052 ( n13228 , n11114 , n15805 );
    xnor g17053 ( n33999 , n17716 , n4960 );
    or g17054 ( n3966 , n33870 , n18378 );
    nor g17055 ( n5447 , n10545 , n6548 );
    or g17056 ( n3717 , n15353 , n3056 );
    buf g17057 ( n26023 , n33262 );
    and g17058 ( n10487 , n13090 , n26681 );
    or g17059 ( n1748 , n12506 , n18264 );
    or g17060 ( n18728 , n15785 , n17724 );
    nor g17061 ( n7368 , n25602 , n13338 );
    not g17062 ( n11969 , n22980 );
    or g17063 ( n18637 , n33739 , n32505 );
    or g17064 ( n21036 , n31787 , n15109 );
    or g17065 ( n21724 , n25327 , n4172 );
    and g17066 ( n4206 , n33263 , n18909 );
    not g17067 ( n29266 , n11996 );
    xnor g17068 ( n6873 , n24387 , n12215 );
    or g17069 ( n19358 , n11190 , n17498 );
    or g17070 ( n29113 , n13189 , n17118 );
    xnor g17071 ( n31992 , n35741 , n19551 );
    or g17072 ( n15491 , n1974 , n15439 );
    xnor g17073 ( n12624 , n22280 , n19551 );
    nor g17074 ( n30252 , n8298 , n18113 );
    and g17075 ( n8247 , n31636 , n5681 );
    and g17076 ( n9853 , n13494 , n21556 );
    or g17077 ( n11840 , n14006 , n2366 );
    not g17078 ( n1201 , n23972 );
    and g17079 ( n5921 , n28949 , n21249 );
    or g17080 ( n16482 , n4662 , n17829 );
    or g17081 ( n11095 , n6576 , n33523 );
    xnor g17082 ( n12657 , n26621 , n31056 );
    nor g17083 ( n16078 , n16620 , n34246 );
    and g17084 ( n30530 , n29582 , n12216 );
    not g17085 ( n4279 , n18296 );
    or g17086 ( n11016 , n11202 , n28324 );
    and g17087 ( n26622 , n466 , n26412 );
    nor g17088 ( n15402 , n1519 , n17173 );
    and g17089 ( n22127 , n12856 , n32300 );
    or g17090 ( n26459 , n29517 , n2994 );
    or g17091 ( n4854 , n5760 , n11295 );
    nor g17092 ( n13884 , n4288 , n16538 );
    xnor g17093 ( n3768 , n875 , n9429 );
    not g17094 ( n16773 , n7540 );
    or g17095 ( n16266 , n15886 , n26047 );
    xnor g17096 ( n12650 , n15671 , n11990 );
    and g17097 ( n12857 , n28226 , n3038 );
    and g17098 ( n31848 , n26187 , n20750 );
    xnor g17099 ( n20926 , n32477 , n29839 );
    and g17100 ( n26386 , n17055 , n31504 );
    or g17101 ( n461 , n23703 , n15024 );
    xnor g17102 ( n31751 , n28182 , n4288 );
    and g17103 ( n31939 , n1733 , n30377 );
    xnor g17104 ( n25727 , n21802 , n30742 );
    or g17105 ( n24183 , n13556 , n21725 );
    not g17106 ( n3072 , n13967 );
    and g17107 ( n24240 , n32736 , n24032 );
    xnor g17108 ( n15277 , n13910 , n32095 );
    xnor g17109 ( n5539 , n29929 , n32095 );
    or g17110 ( n15576 , n22494 , n1419 );
    xnor g17111 ( n8015 , n5165 , n7734 );
    or g17112 ( n12274 , n3367 , n29585 );
    xnor g17113 ( n14607 , n4487 , n25387 );
    or g17114 ( n2785 , n31400 , n9317 );
    xnor g17115 ( n33535 , n31851 , n13518 );
    or g17116 ( n33175 , n7272 , n5868 );
    and g17117 ( n7773 , n31885 , n29217 );
    or g17118 ( n19179 , n2576 , n21349 );
    or g17119 ( n11558 , n33780 , n12026 );
    and g17120 ( n20917 , n24535 , n1186 );
    xnor g17121 ( n13188 , n25030 , n13881 );
    and g17122 ( n20920 , n23301 , n14 );
    not g17123 ( n3990 , n31125 );
    buf g17124 ( n28123 , n25629 );
    not g17125 ( n5804 , n4594 );
    or g17126 ( n20495 , n9793 , n34224 );
    or g17127 ( n24320 , n10984 , n22783 );
    and g17128 ( n32026 , n25661 , n19984 );
    or g17129 ( n24227 , n26101 , n2117 );
    and g17130 ( n29436 , n31854 , n31735 );
    and g17131 ( n15590 , n35702 , n6256 );
    nor g17132 ( n9596 , n15403 , n1663 );
    or g17133 ( n15851 , n31324 , n23128 );
    buf g17134 ( n2005 , n3239 );
    not g17135 ( n27191 , n26535 );
    xnor g17136 ( n3176 , n4357 , n11046 );
    not g17137 ( n14890 , n1041 );
    or g17138 ( n9073 , n18022 , n6394 );
    xnor g17139 ( n10351 , n34119 , n6785 );
    or g17140 ( n158 , n31799 , n8716 );
    not g17141 ( n33121 , n22980 );
    or g17142 ( n35745 , n34008 , n19939 );
    nor g17143 ( n18950 , n32857 , n16197 );
    xnor g17144 ( n16911 , n18661 , n4878 );
    nor g17145 ( n13057 , n19984 , n25661 );
    or g17146 ( n13994 , n25205 , n4610 );
    and g17147 ( n22480 , n14451 , n19792 );
    or g17148 ( n23742 , n10269 , n13217 );
    or g17149 ( n27450 , n14425 , n22276 );
    nor g17150 ( n22160 , n21717 , n27745 );
    nor g17151 ( n30963 , n32857 , n8595 );
    or g17152 ( n31886 , n31559 , n11314 );
    or g17153 ( n13111 , n9658 , n15537 );
    or g17154 ( n13946 , n26047 , n5252 );
    xnor g17155 ( n34769 , n25196 , n15090 );
    or g17156 ( n21059 , n2363 , n32961 );
    or g17157 ( n18294 , n15683 , n19123 );
    and g17158 ( n17221 , n36054 , n29291 );
    or g17159 ( n26415 , n15838 , n14076 );
    or g17160 ( n488 , n462 , n22241 );
    not g17161 ( n24570 , n30669 );
    xnor g17162 ( n4194 , n23133 , n28286 );
    nor g17163 ( n18074 , n30742 , n35666 );
    xnor g17164 ( n17863 , n12904 , n10695 );
    or g17165 ( n32709 , n30965 , n29562 );
    and g17166 ( n773 , n8589 , n1692 );
    xnor g17167 ( n262 , n7969 , n4646 );
    xnor g17168 ( n29385 , n29945 , n32095 );
    xnor g17169 ( n28942 , n17427 , n13618 );
    or g17170 ( n4005 , n12512 , n27973 );
    nor g17171 ( n33988 , n11455 , n19820 );
    xnor g17172 ( n32482 , n35517 , n10507 );
    xnor g17173 ( n24669 , n9534 , n23288 );
    or g17174 ( n4650 , n31799 , n33533 );
    not g17175 ( n35168 , n3480 );
    and g17176 ( n28702 , n33322 , n22920 );
    or g17177 ( n9365 , n27298 , n21691 );
    xnor g17178 ( n33669 , n29225 , n23604 );
    nor g17179 ( n19345 , n31289 , n1673 );
    and g17180 ( n4233 , n31717 , n9859 );
    or g17181 ( n20939 , n2421 , n15110 );
    xnor g17182 ( n28683 , n13894 , n8105 );
    not g17183 ( n12510 , n28474 );
    or g17184 ( n18764 , n25282 , n25255 );
    xnor g17185 ( n28585 , n29329 , n31093 );
    xnor g17186 ( n8767 , n26701 , n29839 );
    and g17187 ( n8210 , n30247 , n15789 );
    and g17188 ( n6579 , n10187 , n35531 );
    and g17189 ( n8352 , n9619 , n19012 );
    or g17190 ( n33636 , n2118 , n32329 );
    or g17191 ( n20569 , n9923 , n33677 );
    nor g17192 ( n6806 , n34415 , n32720 );
    and g17193 ( n9489 , n1728 , n29730 );
    nor g17194 ( n9641 , n31559 , n31966 );
    xnor g17195 ( n29509 , n28814 , n7535 );
    xnor g17196 ( n34671 , n34150 , n31559 );
    or g17197 ( n30584 , n13866 , n31134 );
    nor g17198 ( n2845 , n31314 , n28757 );
    or g17199 ( n16816 , n27265 , n9447 );
    or g17200 ( n33861 , n11059 , n35339 );
    and g17201 ( n21419 , n9823 , n6672 );
    and g17202 ( n9204 , n27141 , n25341 );
    and g17203 ( n33093 , n4144 , n788 );
    or g17204 ( n36018 , n11775 , n30419 );
    nor g17205 ( n34700 , n30345 , n34635 );
    or g17206 ( n3453 , n14947 , n5208 );
    or g17207 ( n25291 , n13879 , n28438 );
    or g17208 ( n31271 , n617 , n2667 );
    nor g17209 ( n2185 , n21409 , n19215 );
    xnor g17210 ( n2953 , n16992 , n32095 );
    xnor g17211 ( n24817 , n14879 , n22480 );
    or g17212 ( n16618 , n12686 , n5113 );
    or g17213 ( n35069 , n19407 , n16919 );
    or g17214 ( n1104 , n23077 , n20853 );
    or g17215 ( n7624 , n33052 , n28248 );
    or g17216 ( n29392 , n34665 , n10634 );
    nor g17217 ( n17044 , n9789 , n24979 );
    and g17218 ( n8045 , n24659 , n10152 );
    xnor g17219 ( n6377 , n18532 , n7369 );
    or g17220 ( n9971 , n28616 , n15805 );
    not g17221 ( n19619 , n2029 );
    or g17222 ( n19232 , n16620 , n31349 );
    or g17223 ( n24660 , n29713 , n25068 );
    or g17224 ( n8726 , n35927 , n15827 );
    not g17225 ( n11127 , n25648 );
    or g17226 ( n13416 , n17312 , n19687 );
    and g17227 ( n6285 , n7740 , n925 );
    or g17228 ( n25138 , n11455 , n6842 );
    or g17229 ( n34295 , n28349 , n28191 );
    nor g17230 ( n18205 , n31799 , n27658 );
    or g17231 ( n20089 , n10758 , n5168 );
    nor g17232 ( n111 , n23478 , n24555 );
    or g17233 ( n10719 , n5931 , n11194 );
    not g17234 ( n8892 , n20558 );
    xnor g17235 ( n9721 , n23694 , n29502 );
    or g17236 ( n1334 , n1217 , n29124 );
    not g17237 ( n5114 , n31559 );
    or g17238 ( n24384 , n2831 , n34680 );
    xnor g17239 ( n34805 , n21654 , n1950 );
    nor g17240 ( n19707 , n1331 , n7353 );
    or g17241 ( n23478 , n13377 , n31517 );
    or g17242 ( n7871 , n6506 , n3438 );
    nor g17243 ( n2431 , n4962 , n12955 );
    nor g17244 ( n15977 , n34743 , n31633 );
    and g17245 ( n27095 , n6471 , n33391 );
    and g17246 ( n29038 , n30266 , n29171 );
    xnor g17247 ( n26588 , n3854 , n27011 );
    xnor g17248 ( n2081 , n12410 , n31338 );
    or g17249 ( n13838 , n555 , n11312 );
    or g17250 ( n14902 , n7540 , n3071 );
    and g17251 ( n35249 , n33051 , n21809 );
    and g17252 ( n19575 , n13049 , n35274 );
    not g17253 ( n29365 , n3671 );
    not g17254 ( n34461 , n9793 );
    and g17255 ( n20066 , n9680 , n6238 );
    not g17256 ( n1728 , n2259 );
    or g17257 ( n20800 , n23697 , n19686 );
    xnor g17258 ( n28527 , n11134 , n1846 );
    or g17259 ( n20895 , n6059 , n20576 );
    not g17260 ( n474 , n16223 );
    xnor g17261 ( n25090 , n3739 , n2386 );
    nor g17262 ( n14749 , n16135 , n35051 );
    or g17263 ( n28950 , n6789 , n23469 );
    and g17264 ( n25825 , n9636 , n18904 );
    or g17265 ( n6986 , n3205 , n5677 );
    not g17266 ( n19664 , n3205 );
    or g17267 ( n29965 , n11280 , n25405 );
    xnor g17268 ( n12345 , n24421 , n20399 );
    xnor g17269 ( n4685 , n35876 , n27264 );
    and g17270 ( n17364 , n20545 , n24986 );
    and g17271 ( n17045 , n30643 , n11154 );
    or g17272 ( n15615 , n18532 , n7369 );
    not g17273 ( n4751 , n30732 );
    not g17274 ( n743 , n33312 );
    or g17275 ( n3413 , n20604 , n9731 );
    xnor g17276 ( n4776 , n16222 , n14976 );
    and g17277 ( n33698 , n7567 , n9333 );
    or g17278 ( n5751 , n35962 , n23101 );
    or g17279 ( n15908 , n12907 , n10140 );
    or g17280 ( n3845 , n3183 , n30732 );
    or g17281 ( n7558 , n35927 , n1660 );
    xnor g17282 ( n15683 , n15755 , n4960 );
    or g17283 ( n6301 , n28412 , n19241 );
    nor g17284 ( n1648 , n28958 , n31502 );
    and g17285 ( n10828 , n21170 , n21336 );
    nor g17286 ( n35394 , n26124 , n27583 );
    or g17287 ( n16089 , n7130 , n18811 );
    or g17288 ( n15063 , n6674 , n4470 );
    xnor g17289 ( n11637 , n12135 , n11455 );
    and g17290 ( n16417 , n22297 , n29213 );
    or g17291 ( n18467 , n10563 , n2104 );
    or g17292 ( n4417 , n12130 , n23382 );
    or g17293 ( n35194 , n4878 , n11233 );
    and g17294 ( n19001 , n30910 , n31139 );
    and g17295 ( n12949 , n30351 , n15275 );
    or g17296 ( n25891 , n31948 , n11703 );
    and g17297 ( n15398 , n24354 , n35592 );
    and g17298 ( n22719 , n10271 , n13140 );
    nor g17299 ( n34981 , n32857 , n5039 );
    buf g17300 ( n6288 , n19901 );
    and g17301 ( n9938 , n10029 , n23238 );
    or g17302 ( n2612 , n31215 , n14737 );
    nor g17303 ( n1337 , n9090 , n9921 );
    xnor g17304 ( n16914 , n11087 , n21306 );
    and g17305 ( n22244 , n34302 , n153 );
    and g17306 ( n5092 , n9393 , n2785 );
    and g17307 ( n24336 , n19613 , n12072 );
    nor g17308 ( n29290 , n11507 , n26553 );
    or g17309 ( n19382 , n17568 , n30665 );
    nor g17310 ( n1943 , n4962 , n11406 );
    and g17311 ( n146 , n15630 , n22592 );
    or g17312 ( n30437 , n33151 , n19490 );
    not g17313 ( n11155 , n29792 );
    or g17314 ( n27935 , n13270 , n26988 );
    xnor g17315 ( n24675 , n36015 , n34016 );
    xnor g17316 ( n6895 , n12196 , n22580 );
    xnor g17317 ( n29457 , n1570 , n26939 );
    nor g17318 ( n22687 , n10894 , n17458 );
    xnor g17319 ( n18768 , n25934 , n21783 );
    and g17320 ( n19170 , n21117 , n23965 );
    xnor g17321 ( n29153 , n34462 , n11013 );
    xnor g17322 ( n16848 , n33226 , n1311 );
    and g17323 ( n21494 , n9342 , n4879 );
    or g17324 ( n34831 , n6503 , n13217 );
    or g17325 ( n4455 , n28439 , n2959 );
    or g17326 ( n23778 , n21015 , n28574 );
    or g17327 ( n25000 , n22750 , n8392 );
    and g17328 ( n29318 , n7216 , n190 );
    or g17329 ( n24612 , n8026 , n10140 );
    or g17330 ( n27672 , n16232 , n21739 );
    not g17331 ( n12644 , n6793 );
    and g17332 ( n12667 , n7176 , n33574 );
    and g17333 ( n5961 , n24782 , n29653 );
    or g17334 ( n27965 , n28634 , n9915 );
    nor g17335 ( n9047 , n10596 , n31411 );
    xnor g17336 ( n21840 , n23997 , n27645 );
    or g17337 ( n13119 , n13197 , n15642 );
    not g17338 ( n29465 , n6218 );
    or g17339 ( n33081 , n34438 , n4363 );
    and g17340 ( n8537 , n19637 , n30331 );
    or g17341 ( n24638 , n28033 , n26480 );
    or g17342 ( n27967 , n24902 , n4478 );
    and g17343 ( n6556 , n21472 , n18541 );
    nor g17344 ( n14777 , n23175 , n5124 );
    xnor g17345 ( n19468 , n25835 , n8432 );
    and g17346 ( n19005 , n19452 , n29440 );
    not g17347 ( n28168 , n4962 );
    and g17348 ( n9387 , n35191 , n5131 );
    xnor g17349 ( n20470 , n15267 , n9658 );
    or g17350 ( n35252 , n2625 , n8366 );
    xnor g17351 ( n17933 , n35812 , n18049 );
    or g17352 ( n34261 , n11538 , n19058 );
    or g17353 ( n30007 , n30742 , n21261 );
    or g17354 ( n10661 , n30416 , n16345 );
    and g17355 ( n21207 , n8593 , n1573 );
    or g17356 ( n34382 , n30553 , n25189 );
    or g17357 ( n23401 , n16607 , n19594 );
    or g17358 ( n1385 , n24613 , n4069 );
    and g17359 ( n21272 , n12369 , n16683 );
    xnor g17360 ( n11697 , n3835 , n15886 );
    or g17361 ( n24494 , n1950 , n1643 );
    or g17362 ( n33611 , n29525 , n14588 );
    nor g17363 ( n13470 , n29884 , n21658 );
    xnor g17364 ( n35283 , n15597 , n32073 );
    or g17365 ( n17916 , n13308 , n16072 );
    xnor g17366 ( n8556 , n24629 , n13795 );
    or g17367 ( n26968 , n19551 , n18218 );
    and g17368 ( n36084 , n18816 , n4617 );
    nor g17369 ( n14503 , n15886 , n19630 );
    or g17370 ( n12522 , n9293 , n15028 );
    or g17371 ( n32057 , n15822 , n7547 );
    or g17372 ( n20283 , n9054 , n19910 );
    or g17373 ( n6930 , n16078 , n30620 );
    or g17374 ( n9794 , n7262 , n13015 );
    and g17375 ( n13776 , n15092 , n3567 );
    not g17376 ( n35764 , n18991 );
    nor g17377 ( n11716 , n13436 , n7565 );
    or g17378 ( n16053 , n15464 , n21588 );
    or g17379 ( n15404 , n4878 , n24302 );
    and g17380 ( n28 , n2696 , n1081 );
    or g17381 ( n35055 , n35580 , n25447 );
    xnor g17382 ( n27479 , n27734 , n24371 );
    xnor g17383 ( n12673 , n22579 , n13841 );
    or g17384 ( n6794 , n6962 , n32141 );
    xnor g17385 ( n29652 , n30407 , n31018 );
    xnor g17386 ( n10350 , n20209 , n35451 );
    xnor g17387 ( n11264 , n25803 , n6229 );
    and g17388 ( n9575 , n9743 , n1791 );
    xnor g17389 ( n1467 , n14373 , n10420 );
    or g17390 ( n86 , n20924 , n32071 );
    or g17391 ( n6754 , n1645 , n33000 );
    and g17392 ( n13394 , n17865 , n27332 );
    xnor g17393 ( n16280 , n33397 , n4878 );
    and g17394 ( n33951 , n30894 , n12631 );
    and g17395 ( n30461 , n32094 , n7080 );
    not g17396 ( n10412 , n10455 );
    or g17397 ( n1212 , n19629 , n10140 );
    and g17398 ( n7544 , n12270 , n258 );
    xnor g17399 ( n28125 , n22558 , n14447 );
    xnor g17400 ( n21639 , n26236 , n1047 );
    not g17401 ( n35525 , n6837 );
    xnor g17402 ( n9334 , n26529 , n14056 );
    not g17403 ( n8594 , n20558 );
    and g17404 ( n15209 , n28017 , n12279 );
    nor g17405 ( n19816 , n22047 , n15002 );
    and g17406 ( n27108 , n3169 , n23372 );
    and g17407 ( n10021 , n8202 , n13680 );
    xnor g17408 ( n20619 , n24842 , n28477 );
    xnor g17409 ( n27289 , n15900 , n14835 );
    and g17410 ( n17806 , n30544 , n2966 );
    xnor g17411 ( n28005 , n31620 , n20068 );
    xnor g17412 ( n35023 , n17123 , n33606 );
    or g17413 ( n10569 , n8241 , n8723 );
    or g17414 ( n20606 , n29884 , n28659 );
    and g17415 ( n14883 , n33123 , n6101 );
    xnor g17416 ( n22150 , n17526 , n4878 );
    or g17417 ( n10608 , n24371 , n34667 );
    or g17418 ( n11395 , n28713 , n6683 );
    or g17419 ( n20313 , n18958 , n2384 );
    nor g17420 ( n31562 , n18620 , n27924 );
    or g17421 ( n32542 , n11333 , n3738 );
    or g17422 ( n32552 , n8651 , n17664 );
    or g17423 ( n18128 , n24684 , n32944 );
    and g17424 ( n684 , n34984 , n3313 );
    xnor g17425 ( n12108 , n12640 , n10115 );
    and g17426 ( n11499 , n114 , n160 );
    xnor g17427 ( n11873 , n19603 , n4878 );
    or g17428 ( n21849 , n29713 , n12490 );
    or g17429 ( n22146 , n4758 , n10110 );
    xnor g17430 ( n23351 , n21245 , n388 );
    or g17431 ( n28205 , n21529 , n12927 );
    and g17432 ( n5226 , n18519 , n11696 );
    nor g17433 ( n4793 , n3205 , n15659 );
    or g17434 ( n24894 , n13476 , n22096 );
    or g17435 ( n499 , n32715 , n2650 );
    or g17436 ( n8363 , n17751 , n5549 );
    not g17437 ( n28758 , n11350 );
    and g17438 ( n18935 , n10481 , n3018 );
    xnor g17439 ( n8464 , n28367 , n7474 );
    or g17440 ( n8051 , n2318 , n33098 );
    nor g17441 ( n28276 , n17568 , n33043 );
    xnor g17442 ( n20726 , n20398 , n3762 );
    or g17443 ( n10838 , n17187 , n21977 );
    xnor g17444 ( n4494 , n20875 , n1700 );
    not g17445 ( n5204 , n35491 );
    not g17446 ( n28840 , n3205 );
    and g17447 ( n13241 , n13787 , n27210 );
    xnor g17448 ( n30438 , n16324 , n30742 );
    or g17449 ( n35090 , n35268 , n25482 );
    and g17450 ( n22614 , n7486 , n16148 );
    or g17451 ( n29930 , n4395 , n30605 );
    or g17452 ( n34116 , n24371 , n13349 );
    and g17453 ( n20775 , n2479 , n28665 );
    nor g17454 ( n27678 , n4960 , n17774 );
    or g17455 ( n29004 , n4948 , n3847 );
    or g17456 ( n5238 , n19580 , n26220 );
    or g17457 ( n5758 , n1533 , n16464 );
    and g17458 ( n29502 , n15063 , n19357 );
    xnor g17459 ( n1277 , n3751 , n11190 );
    or g17460 ( n15931 , n15886 , n14448 );
    xnor g17461 ( n17634 , n11401 , n15886 );
    or g17462 ( n5889 , n27175 , n25019 );
    or g17463 ( n30496 , n23987 , n29411 );
    or g17464 ( n23313 , n16872 , n19732 );
    xnor g17465 ( n3271 , n21067 , n29299 );
    and g17466 ( n19286 , n32514 , n27223 );
    xnor g17467 ( n129 , n25422 , n4288 );
    or g17468 ( n16815 , n4698 , n25940 );
    xnor g17469 ( n19711 , n26383 , n34222 );
    or g17470 ( n3208 , n23435 , n17974 );
    not g17471 ( n34048 , n17068 );
    and g17472 ( n3364 , n13295 , n16838 );
    xnor g17473 ( n5689 , n23057 , n10625 );
    not g17474 ( n27699 , n25436 );
    and g17475 ( n27812 , n26186 , n33131 );
    and g17476 ( n8440 , n9133 , n32767 );
    nor g17477 ( n8491 , n32857 , n14336 );
    or g17478 ( n5073 , n4845 , n30255 );
    or g17479 ( n10898 , n9789 , n839 );
    or g17480 ( n12321 , n13504 , n14818 );
    xnor g17481 ( n783 , n35727 , n32857 );
    or g17482 ( n7218 , n32295 , n3694 );
    xnor g17483 ( n4782 , n25116 , n26736 );
    or g17484 ( n23427 , n16796 , n19707 );
    and g17485 ( n5924 , n13815 , n7 );
    and g17486 ( n22477 , n31835 , n9992 );
    and g17487 ( n15820 , n8527 , n17326 );
    xnor g17488 ( n21715 , n15634 , n29962 );
    xnor g17489 ( n34786 , n33327 , n27291 );
    or g17490 ( n7911 , n22070 , n12996 );
    xnor g17491 ( n16467 , n1880 , n26656 );
    or g17492 ( n21736 , n14332 , n1796 );
    and g17493 ( n13077 , n6110 , n26042 );
    and g17494 ( n17243 , n10272 , n26093 );
    and g17495 ( n12495 , n27330 , n28195 );
    or g17496 ( n2526 , n683 , n4254 );
    and g17497 ( n25970 , n20743 , n11572 );
    and g17498 ( n18189 , n9178 , n34047 );
    or g17499 ( n2707 , n11147 , n4912 );
    xnor g17500 ( n7896 , n22675 , n2039 );
    or g17501 ( n4562 , n897 , n1942 );
    or g17502 ( n33508 , n8654 , n13132 );
    or g17503 ( n19202 , n1153 , n31514 );
    and g17504 ( n19914 , n22420 , n32616 );
    nor g17505 ( n20593 , n21281 , n16659 );
    nor g17506 ( n33719 , n19551 , n10841 );
    xnor g17507 ( n11813 , n21826 , n34614 );
    or g17508 ( n1318 , n14335 , n11816 );
    or g17509 ( n7069 , n32584 , n1343 );
    buf g17510 ( n14361 , n19754 );
    and g17511 ( n35329 , n13415 , n16157 );
    or g17512 ( n21832 , n806 , n35181 );
    xnor g17513 ( n16404 , n32183 , n12598 );
    or g17514 ( n13570 , n15886 , n21798 );
    or g17515 ( n22973 , n8824 , n26366 );
    xnor g17516 ( n14916 , n11632 , n21365 );
    not g17517 ( n19200 , n18844 );
    or g17518 ( n20263 , n5535 , n32281 );
    not g17519 ( n7287 , n4985 );
    or g17520 ( n34070 , n26316 , n17515 );
    buf g17521 ( n30646 , n29676 );
    or g17522 ( n3304 , n23900 , n33656 );
    nor g17523 ( n6576 , n5335 , n28385 );
    and g17524 ( n1312 , n15682 , n17596 );
    or g17525 ( n11627 , n4382 , n8430 );
    xnor g17526 ( n18917 , n10802 , n319 );
    and g17527 ( n31334 , n9674 , n4 );
    buf g17528 ( n2092 , n19918 );
    xnor g17529 ( n30655 , n1634 , n29839 );
    xnor g17530 ( n4280 , n20931 , n10894 );
    and g17531 ( n20104 , n27737 , n12792 );
    nor g17532 ( n31929 , n31799 , n34455 );
    xnor g17533 ( n16718 , n12360 , n8954 );
    xnor g17534 ( n28733 , n25118 , n25984 );
    or g17535 ( n4263 , n4333 , n33908 );
    or g17536 ( n30410 , n899 , n21956 );
    and g17537 ( n30095 , n27932 , n13814 );
    or g17538 ( n5508 , n18263 , n11703 );
    xnor g17539 ( n5334 , n19077 , n13051 );
    xnor g17540 ( n32525 , n20687 , n22575 );
    not g17541 ( n35961 , n28078 );
    or g17542 ( n32209 , n5413 , n3683 );
    xnor g17543 ( n3615 , n30460 , n30357 );
    nor g17544 ( n26825 , n25602 , n27095 );
    or g17545 ( n7059 , n9758 , n6181 );
    not g17546 ( n21358 , n31799 );
    or g17547 ( n2891 , n13867 , n21579 );
    xnor g17548 ( n26843 , n22784 , n3205 );
    or g17549 ( n93 , n18707 , n4058 );
    or g17550 ( n29129 , n2678 , n14382 );
    xnor g17551 ( n10194 , n26156 , n19143 );
    or g17552 ( n19938 , n17568 , n26632 );
    nor g17553 ( n23942 , n24353 , n29393 );
    and g17554 ( n21014 , n19854 , n20451 );
    or g17555 ( n7977 , n16951 , n30646 );
    xnor g17556 ( n35261 , n29878 , n23599 );
    or g17557 ( n10037 , n14421 , n30405 );
    nor g17558 ( n20111 , n31272 , n17182 );
    or g17559 ( n31274 , n28383 , n2111 );
    or g17560 ( n16022 , n15886 , n5609 );
    or g17561 ( n14404 , n23556 , n15344 );
    xnor g17562 ( n21063 , n31802 , n29383 );
    or g17563 ( n28010 , n12586 , n23209 );
    xnor g17564 ( n16968 , n29418 , n21754 );
    or g17565 ( n27248 , n10132 , n23546 );
    xnor g17566 ( n17421 , n33370 , n31140 );
    xnor g17567 ( n30331 , n32255 , n7543 );
    xnor g17568 ( n34514 , n18612 , n4962 );
    and g17569 ( n103 , n35745 , n28916 );
    or g17570 ( n8649 , n14551 , n21634 );
    nor g17571 ( n7728 , n31272 , n34578 );
    xnor g17572 ( n33119 , n9048 , n12457 );
    and g17573 ( n25405 , n8507 , n3049 );
    or g17574 ( n7614 , n5066 , n4490 );
    xnor g17575 ( n15442 , n4585 , n373 );
    xnor g17576 ( n25119 , n33169 , n24795 );
    and g17577 ( n27160 , n1953 , n20978 );
    and g17578 ( n8174 , n27150 , n5973 );
    or g17579 ( n12789 , n17436 , n26737 );
    xnor g17580 ( n4773 , n19833 , n16809 );
    and g17581 ( n22111 , n26831 , n38 );
    or g17582 ( n32755 , n10469 , n13817 );
    and g17583 ( n18794 , n20396 , n11294 );
    or g17584 ( n29943 , n5742 , n29315 );
    xnor g17585 ( n21119 , n18220 , n19257 );
    nor g17586 ( n20723 , n31215 , n3596 );
    or g17587 ( n24388 , n3814 , n14800 );
    or g17588 ( n4431 , n33666 , n5779 );
    or g17589 ( n30827 , n3737 , n34977 );
    and g17590 ( n13975 , n12665 , n19735 );
    or g17591 ( n31857 , n25167 , n20844 );
    and g17592 ( n26407 , n25981 , n19935 );
    or g17593 ( n2498 , n12142 , n7647 );
    nor g17594 ( n33519 , n35523 , n18100 );
    xnor g17595 ( n7505 , n21890 , n6785 );
    or g17596 ( n2491 , n34365 , n33362 );
    or g17597 ( n27093 , n28039 , n32909 );
    or g17598 ( n2836 , n3210 , n29366 );
    or g17599 ( n27110 , n19401 , n24489 );
    and g17600 ( n35633 , n34936 , n31553 );
    or g17601 ( n29951 , n16620 , n28972 );
    or g17602 ( n27219 , n5335 , n11326 );
    xnor g17603 ( n12704 , n12276 , n16486 );
    or g17604 ( n2073 , n18408 , n19732 );
    or g17605 ( n31666 , n24080 , n31134 );
    or g17606 ( n30294 , n34587 , n5752 );
    or g17607 ( n1858 , n30065 , n17070 );
    or g17608 ( n30326 , n18523 , n4790 );
    and g17609 ( n20592 , n32848 , n28239 );
    xnor g17610 ( n14685 , n8586 , n35927 );
    and g17611 ( n13177 , n12220 , n19903 );
    not g17612 ( n9200 , n18596 );
    not g17613 ( n27910 , n30957 );
    and g17614 ( n12595 , n9737 , n13532 );
    or g17615 ( n2816 , n27024 , n16304 );
    or g17616 ( n15352 , n28480 , n30732 );
    buf g17617 ( n23790 , n33013 );
    not g17618 ( n32046 , n4960 );
    and g17619 ( n8627 , n15385 , n34734 );
    xnor g17620 ( n19290 , n14336 , n5289 );
    or g17621 ( n28226 , n9683 , n22869 );
    or g17622 ( n17636 , n4353 , n24479 );
    and g17623 ( n500 , n19313 , n33997 );
    or g17624 ( n20725 , n33522 , n16345 );
    or g17625 ( n11937 , n29836 , n216 );
    not g17626 ( n24981 , n31300 );
    xnor g17627 ( n13445 , n27657 , n15464 );
    and g17628 ( n667 , n269 , n1134 );
    not g17629 ( n34196 , n15158 );
    and g17630 ( n1352 , n31279 , n15437 );
    or g17631 ( n21395 , n27164 , n17354 );
    xnor g17632 ( n27138 , n5015 , n15464 );
    and g17633 ( n9878 , n23053 , n35548 );
    nor g17634 ( n35250 , n5106 , n33157 );
    xnor g17635 ( n1821 , n2141 , n10356 );
    and g17636 ( n7046 , n9826 , n16422 );
    nor g17637 ( n13937 , n19070 , n13610 );
    or g17638 ( n2139 , n11727 , n9194 );
    xnor g17639 ( n31040 , n15924 , n5335 );
    not g17640 ( n34406 , n15578 );
    and g17641 ( n29735 , n32342 , n9639 );
    xnor g17642 ( n35052 , n35432 , n31559 );
    xnor g17643 ( n17889 , n2300 , n23604 );
    xnor g17644 ( n3689 , n13885 , n24691 );
    or g17645 ( n11108 , n7847 , n10432 );
    or g17646 ( n186 , n3889 , n29125 );
    or g17647 ( n17590 , n29713 , n16884 );
    or g17648 ( n21915 , n8846 , n15344 );
    and g17649 ( n16644 , n8504 , n20569 );
    or g17650 ( n10727 , n17995 , n33513 );
    and g17651 ( n29066 , n18256 , n11093 );
    or g17652 ( n18759 , n16465 , n4478 );
    not g17653 ( n27325 , n4960 );
    xnor g17654 ( n8584 , n21662 , n29335 );
    and g17655 ( n9161 , n15823 , n9196 );
    or g17656 ( n9461 , n16367 , n18264 );
    nor g17657 ( n17629 , n7281 , n33826 );
    or g17658 ( n12577 , n30523 , n5816 );
    buf g17659 ( n544 , n9822 );
    or g17660 ( n3289 , n16547 , n16543 );
    and g17661 ( n905 , n32308 , n26975 );
    xnor g17662 ( n34613 , n31131 , n9860 );
    not g17663 ( n34781 , n10894 );
    or g17664 ( n5950 , n22514 , n15290 );
    nor g17665 ( n17572 , n31387 , n18095 );
    and g17666 ( n24759 , n12243 , n32346 );
    nor g17667 ( n29064 , n4288 , n31131 );
    or g17668 ( n26131 , n10010 , n30646 );
    or g17669 ( n8561 , n22227 , n27447 );
    xnor g17670 ( n26733 , n2201 , n2813 );
    or g17671 ( n22893 , n15468 , n31627 );
    or g17672 ( n4136 , n10595 , n4055 );
    nor g17673 ( n547 , n8682 , n14625 );
    and g17674 ( n17322 , n29204 , n19312 );
    and g17675 ( n7587 , n31909 , n9484 );
    and g17676 ( n30373 , n25669 , n6001 );
    or g17677 ( n34321 , n3237 , n9555 );
    or g17678 ( n32365 , n28806 , n19556 );
    nor g17679 ( n11123 , n31799 , n15768 );
    or g17680 ( n25182 , n32095 , n24360 );
    and g17681 ( n30293 , n15152 , n13816 );
    or g17682 ( n21665 , n15045 , n10570 );
    xnor g17683 ( n13489 , n5613 , n27291 );
    and g17684 ( n33706 , n30831 , n1879 );
    not g17685 ( n11954 , n10894 );
    not g17686 ( n18267 , n17568 );
    and g17687 ( n2386 , n9785 , n29682 );
    or g17688 ( n17678 , n3226 , n11831 );
    or g17689 ( n14722 , n4960 , n21410 );
    or g17690 ( n21996 , n35334 , n2845 );
    nor g17691 ( n31501 , n1950 , n5441 );
    or g17692 ( n23434 , n31509 , n1866 );
    or g17693 ( n16529 , n34350 , n15144 );
    xnor g17694 ( n11775 , n25850 , n22691 );
    not g17695 ( n20475 , n17427 );
    or g17696 ( n1177 , n32931 , n4399 );
    and g17697 ( n6698 , n20297 , n25001 );
    and g17698 ( n2300 , n30063 , n14204 );
    and g17699 ( n30084 , n33241 , n25966 );
    xnor g17700 ( n35415 , n685 , n27609 );
    and g17701 ( n15541 , n8097 , n32648 );
    and g17702 ( n22843 , n20385 , n25156 );
    or g17703 ( n21764 , n9609 , n34939 );
    not g17704 ( n4550 , n29799 );
    not g17705 ( n29327 , n1326 );
    and g17706 ( n13562 , n35142 , n3920 );
    or g17707 ( n19564 , n33611 , n13245 );
    buf g17708 ( n8392 , n22924 );
    or g17709 ( n33948 , n1678 , n35297 );
    or g17710 ( n30165 , n14710 , n24505 );
    xnor g17711 ( n8662 , n3295 , n4288 );
    and g17712 ( n29921 , n16603 , n22980 );
    or g17713 ( n3358 , n15825 , n24139 );
    or g17714 ( n1709 , n26743 , n26292 );
    or g17715 ( n35733 , n8462 , n17612 );
    buf g17716 ( n33310 , n28816 );
    not g17717 ( n19946 , n8637 );
    and g17718 ( n15788 , n10711 , n34422 );
    and g17719 ( n6690 , n2023 , n4531 );
    and g17720 ( n12991 , n16921 , n17497 );
    or g17721 ( n31785 , n23590 , n10644 );
    nor g17722 ( n8031 , n17568 , n23115 );
    or g17723 ( n32424 , n9658 , n21012 );
    or g17724 ( n21367 , n31559 , n1500 );
    xnor g17725 ( n12192 , n30036 , n27407 );
    or g17726 ( n9239 , n19304 , n35186 );
    xnor g17727 ( n9321 , n8348 , n23604 );
    xnor g17728 ( n8616 , n1959 , n15675 );
    xnor g17729 ( n4406 , n27399 , n32930 );
    or g17730 ( n26432 , n11046 , n19781 );
    and g17731 ( n23008 , n22716 , n35399 );
    or g17732 ( n1032 , n4960 , n32322 );
    or g17733 ( n33640 , n12334 , n27574 );
    or g17734 ( n10929 , n9137 , n6511 );
    and g17735 ( n25171 , n11761 , n35125 );
    or g17736 ( n26470 , n16924 , n24025 );
    xnor g17737 ( n33446 , n895 , n29185 );
    xnor g17738 ( n24270 , n16319 , n24091 );
    and g17739 ( n24132 , n22957 , n35139 );
    or g17740 ( n19937 , n10894 , n410 );
    or g17741 ( n30288 , n23363 , n9030 );
    xnor g17742 ( n13716 , n9105 , n11046 );
    or g17743 ( n21811 , n18282 , n15109 );
    and g17744 ( n25164 , n7088 , n28506 );
    or g17745 ( n15131 , n27500 , n9213 );
    or g17746 ( n28144 , n3946 , n9827 );
    and g17747 ( n14912 , n10619 , n10284 );
    or g17748 ( n29568 , n8428 , n17068 );
    xnor g17749 ( n11467 , n34072 , n11659 );
    or g17750 ( n15239 , n7003 , n25355 );
    xnor g17751 ( n18246 , n18610 , n4288 );
    xnor g17752 ( n20878 , n11852 , n4288 );
    or g17753 ( n16371 , n5697 , n33833 );
    or g17754 ( n21909 , n27533 , n34700 );
    nor g17755 ( n11496 , n25174 , n35846 );
    or g17756 ( n31791 , n3217 , n12622 );
    and g17757 ( n10662 , n10641 , n22769 );
    nor g17758 ( n3484 , n4758 , n27831 );
    nor g17759 ( n13286 , n35169 , n32387 );
    or g17760 ( n33426 , n3222 , n27046 );
    and g17761 ( n34334 , n24359 , n16789 );
    or g17762 ( n16478 , n8432 , n14366 );
    or g17763 ( n10774 , n29216 , n20966 );
    or g17764 ( n61 , n15987 , n28240 );
    xnor g17765 ( n34052 , n10737 , n32095 );
    or g17766 ( n22395 , n26303 , n32505 );
    not g17767 ( n32588 , n23604 );
    and g17768 ( n16479 , n2642 , n19921 );
    xnor g17769 ( n32633 , n22745 , n21608 );
    or g17770 ( n1991 , n5335 , n9918 );
    or g17771 ( n26586 , n8792 , n10872 );
    and g17772 ( n19446 , n5400 , n26281 );
    xnor g17773 ( n26069 , n1993 , n10730 );
    and g17774 ( n8503 , n23385 , n11953 );
    or g17775 ( n515 , n18247 , n33848 );
    nor g17776 ( n35703 , n22291 , n26910 );
    or g17777 ( n8202 , n26995 , n27695 );
    not g17778 ( n16431 , n21350 );
    and g17779 ( n19485 , n15920 , n11628 );
    not g17780 ( n28993 , n22200 );
    xnor g17781 ( n21104 , n144 , n18333 );
    xor g17782 ( n34255 , n32266 , n4288 );
    or g17783 ( n31526 , n4074 , n16115 );
    not g17784 ( n27404 , n18121 );
    xnor g17785 ( n13014 , n10454 , n26521 );
    and g17786 ( n25301 , n1714 , n12365 );
    xnor g17787 ( n33415 , n34545 , n530 );
    or g17788 ( n10565 , n27190 , n18264 );
    or g17789 ( n26181 , n33911 , n2955 );
    or g17790 ( n18687 , n13071 , n29007 );
    and g17791 ( n13337 , n8099 , n30169 );
    xnor g17792 ( n4105 , n23107 , n34616 );
    xnor g17793 ( n3403 , n14037 , n2727 );
    or g17794 ( n12884 , n32543 , n25594 );
    buf g17795 ( n8153 , n5752 );
    or g17796 ( n32993 , n6011 , n34431 );
    or g17797 ( n1336 , n7610 , n25810 );
    xnor g17798 ( n34499 , n21769 , n12304 );
    or g17799 ( n18702 , n17285 , n26659 );
    xnor g17800 ( n6438 , n10434 , n8886 );
    xnor g17801 ( n32109 , n29410 , n2683 );
    xnor g17802 ( n21090 , n8793 , n32414 );
    or g17803 ( n15510 , n4898 , n20797 );
    nor g17804 ( n22763 , n4960 , n17899 );
    or g17805 ( n26775 , n14217 , n9308 );
    or g17806 ( n24640 , n13196 , n35977 );
    or g17807 ( n17645 , n32502 , n22646 );
    or g17808 ( n21259 , n19551 , n28490 );
    not g17809 ( n4661 , n30732 );
    xnor g17810 ( n22842 , n28007 , n25419 );
    or g17811 ( n8127 , n20952 , n5868 );
    and g17812 ( n8324 , n20003 , n34642 );
    not g17813 ( n5866 , n20851 );
    and g17814 ( n20651 , n32079 , n7067 );
    and g17815 ( n2894 , n30083 , n29173 );
    xnor g17816 ( n11505 , n16583 , n24371 );
    nor g17817 ( n10403 , n22511 , n16007 );
    xnor g17818 ( n2402 , n10454 , n16087 );
    or g17819 ( n24153 , n4667 , n12326 );
    not g17820 ( n27327 , n31056 );
    or g17821 ( n8545 , n6055 , n742 );
    xnor g17822 ( n7502 , n17886 , n26048 );
    not g17823 ( n19602 , n27851 );
    or g17824 ( n8810 , n3255 , n26890 );
    or g17825 ( n10846 , n10621 , n35764 );
    and g17826 ( n18769 , n24293 , n11009 );
    or g17827 ( n13061 , n24444 , n24262 );
    or g17828 ( n10790 , n9578 , n8300 );
    and g17829 ( n27657 , n4312 , n1748 );
    xnor g17830 ( n17786 , n29887 , n3205 );
    xnor g17831 ( n19397 , n8044 , n1950 );
    and g17832 ( n27785 , n33283 , n25464 );
    not g17833 ( n8937 , n2092 );
    and g17834 ( n7061 , n23366 , n8998 );
    and g17835 ( n20159 , n9043 , n23243 );
    or g17836 ( n13115 , n31594 , n31896 );
    nor g17837 ( n4075 , n16620 , n5009 );
    or g17838 ( n6905 , n18778 , n26365 );
    and g17839 ( n27472 , n14615 , n17011 );
    xnor g17840 ( n15843 , n18448 , n16217 );
    xnor g17841 ( n12408 , n5773 , n32095 );
    xnor g17842 ( n17823 , n24422 , n20877 );
    and g17843 ( n16647 , n9436 , n31197 );
    xnor g17844 ( n21378 , n31223 , n2015 );
    or g17845 ( n6379 , n23579 , n27447 );
    xnor g17846 ( n27230 , n23954 , n25547 );
    xnor g17847 ( n9829 , n28661 , n8092 );
    and g17848 ( n21604 , n7899 , n20409 );
    not g17849 ( n25354 , n18925 );
    or g17850 ( n34871 , n24105 , n614 );
    xnor g17851 ( n23855 , n16788 , n11952 );
    and g17852 ( n13490 , n6750 , n9621 );
    nor g17853 ( n27342 , n31272 , n7705 );
    or g17854 ( n9186 , n9547 , n26023 );
    or g17855 ( n34211 , n6047 , n30287 );
    xnor g17856 ( n30022 , n25088 , n31744 );
    or g17857 ( n13248 , n5026 , n13449 );
    or g17858 ( n5638 , n19478 , n19421 );
    nor g17859 ( n1280 , n29839 , n31332 );
    xnor g17860 ( n22838 , n27849 , n9789 );
    or g17861 ( n30543 , n30116 , n1763 );
    or g17862 ( n3449 , n25025 , n27704 );
    and g17863 ( n32058 , n16861 , n13242 );
    or g17864 ( n24671 , n31012 , n33310 );
    or g17865 ( n22462 , n18139 , n3188 );
    or g17866 ( n35145 , n21700 , n19218 );
    or g17867 ( n25707 , n27804 , n9675 );
    or g17868 ( n295 , n32520 , n12332 );
    and g17869 ( n15047 , n18607 , n22333 );
    or g17870 ( n32398 , n10174 , n11252 );
    or g17871 ( n9941 , n33905 , n26642 );
    xnor g17872 ( n33945 , n25249 , n25602 );
    and g17873 ( n2039 , n26218 , n32888 );
    xnor g17874 ( n6315 , n19204 , n12347 );
    or g17875 ( n31579 , n27288 , n11977 );
    and g17876 ( n17774 , n11720 , n30694 );
    or g17877 ( n31341 , n15403 , n20488 );
    xnor g17878 ( n25030 , n25740 , n1479 );
    or g17879 ( n18733 , n7760 , n22682 );
    or g17880 ( n22009 , n33463 , n16390 );
    or g17881 ( n34338 , n10894 , n20931 );
    or g17882 ( n5427 , n6134 , n13307 );
    or g17883 ( n11286 , n23840 , n15486 );
    or g17884 ( n34692 , n7540 , n15559 );
    and g17885 ( n25742 , n17392 , n8390 );
    or g17886 ( n25532 , n19013 , n13664 );
    xnor g17887 ( n22020 , n34491 , n31289 );
    and g17888 ( n27590 , n18595 , n24482 );
    or g17889 ( n16645 , n13812 , n19575 );
    not g17890 ( n22583 , n22120 );
    not g17891 ( n33248 , n2433 );
    and g17892 ( n35523 , n1641 , n22980 );
    xnor g17893 ( n16872 , n22526 , n16569 );
    or g17894 ( n14583 , n29839 , n20188 );
    and g17895 ( n13702 , n34233 , n17909 );
    not g17896 ( n35048 , n10602 );
    xnor g17897 ( n32174 , n19191 , n511 );
    and g17898 ( n17682 , n29556 , n19004 );
    nor g17899 ( n23469 , n16280 , n27257 );
    xnor g17900 ( n1936 , n29892 , n22318 );
    buf g17901 ( n10762 , n35422 );
    xnor g17902 ( n7868 , n17836 , n24323 );
    and g17903 ( n20206 , n31519 , n20672 );
    or g17904 ( n25028 , n29648 , n6340 );
    nor g17905 ( n18703 , n15334 , n31699 );
    nor g17906 ( n11292 , n25174 , n2221 );
    nor g17907 ( n7693 , n15886 , n32774 );
    not g17908 ( n25910 , n29462 );
    or g17909 ( n30966 , n2455 , n7153 );
    or g17910 ( n2390 , n31703 , n7113 );
    nor g17911 ( n4193 , n8325 , n20905 );
    or g17912 ( n31904 , n4080 , n28159 );
    and g17913 ( n12015 , n19014 , n11088 );
    or g17914 ( n29690 , n22291 , n13348 );
    xnor g17915 ( n26671 , n26238 , n31215 );
    or g17916 ( n18324 , n18915 , n1320 );
    xnor g17917 ( n25377 , n29320 , n16640 );
    or g17918 ( n2378 , n5987 , n9668 );
    or g17919 ( n7462 , n25998 , n30700 );
    or g17920 ( n18971 , n5738 , n3729 );
    not g17921 ( n6791 , n32857 );
    or g17922 ( n215 , n8513 , n4254 );
    or g17923 ( n4356 , n16922 , n35802 );
    xnor g17924 ( n33967 , n8274 , n30742 );
    xnor g17925 ( n18453 , n15733 , n31799 );
    or g17926 ( n2582 , n9658 , n25543 );
    xnor g17927 ( n33567 , n23971 , n35547 );
    or g17928 ( n18058 , n1855 , n8039 );
    and g17929 ( n3543 , n9286 , n21578 );
    or g17930 ( n10135 , n10206 , n25837 );
    or g17931 ( n25014 , n15464 , n9190 );
    or g17932 ( n3729 , n29496 , n31435 );
    or g17933 ( n1324 , n12639 , n30010 );
    or g17934 ( n27103 , n21121 , n11312 );
    and g17935 ( n17885 , n20335 , n28426 );
    or g17936 ( n16900 , n16024 , n1796 );
    or g17937 ( n35487 , n4835 , n27574 );
    and g17938 ( n4454 , n33998 , n28508 );
    nor g17939 ( n27500 , n3729 , n31411 );
    xnor g17940 ( n30881 , n30085 , n15435 );
    xnor g17941 ( n23923 , n25118 , n34172 );
    and g17942 ( n36039 , n5759 , n9292 );
    not g17943 ( n16656 , n4960 );
    or g17944 ( n28948 , n35927 , n3316 );
    and g17945 ( n33655 , n21919 , n34358 );
    not g17946 ( n32167 , n14292 );
    nor g17947 ( n32185 , n33650 , n35965 );
    or g17948 ( n31697 , n27291 , n22272 );
    and g17949 ( n878 , n14521 , n8436 );
    and g17950 ( n22846 , n23705 , n21617 );
    not g17951 ( n25314 , n11502 );
    or g17952 ( n15513 , n3493 , n17988 );
    or g17953 ( n34904 , n3956 , n18255 );
    xnor g17954 ( n18977 , n30184 , n8730 );
    and g17955 ( n9534 , n30757 , n340 );
    or g17956 ( n31918 , n11722 , n28406 );
    not g17957 ( n33822 , n21087 );
    or g17958 ( n24809 , n14603 , n29411 );
    and g17959 ( n28113 , n34304 , n5983 );
    not g17960 ( n5008 , n30292 );
    or g17961 ( n3644 , n10579 , n286 );
    or g17962 ( n30257 , n20402 , n26737 );
    or g17963 ( n23835 , n28750 , n5618 );
    xnor g17964 ( n29243 , n10449 , n10110 );
    xnor g17965 ( n25432 , n29456 , n33430 );
    and g17966 ( n876 , n18856 , n6387 );
    and g17967 ( n31012 , n25254 , n32566 );
    and g17968 ( n23825 , n23999 , n21632 );
    and g17969 ( n14696 , n25522 , n17947 );
    xnor g17970 ( n15286 , n28647 , n23604 );
    or g17971 ( n12051 , n20855 , n3680 );
    and g17972 ( n32703 , n13440 , n28732 );
    or g17973 ( n23263 , n16489 , n13451 );
    and g17974 ( n1840 , n24995 , n21517 );
    or g17975 ( n34478 , n31799 , n13010 );
    or g17976 ( n9215 , n32584 , n19217 );
    or g17977 ( n2062 , n30742 , n16733 );
    or g17978 ( n4569 , n20700 , n23090 );
    xnor g17979 ( n35246 , n25414 , n17751 );
    and g17980 ( n15784 , n1569 , n2154 );
    and g17981 ( n1505 , n5994 , n6446 );
    or g17982 ( n24089 , n19985 , n15109 );
    and g17983 ( n30987 , n15223 , n6886 );
    or g17984 ( n11107 , n830 , n26915 );
    and g17985 ( n35696 , n24158 , n4211 );
    nor g17986 ( n12751 , n32568 , n3847 );
    nor g17987 ( n7071 , n6499 , n8953 );
    and g17988 ( n21159 , n21779 , n12689 );
    or g17989 ( n10501 , n30215 , n8153 );
    not g17990 ( n30969 , n28500 );
    and g17991 ( n22082 , n6853 , n35218 );
    or g17992 ( n6300 , n28302 , n21977 );
    xor g17993 ( n30614 , n1409 , n19229 );
    xnor g17994 ( n34566 , n4500 , n21631 );
    or g17995 ( n21066 , n18677 , n29445 );
    xnor g17996 ( n17938 , n20492 , n11455 );
    and g17997 ( n8636 , n26086 , n13330 );
    nor g17998 ( n26813 , n35793 , n26826 );
    or g17999 ( n27609 , n22298 , n23572 );
    nor g18000 ( n12175 , n29097 , n3550 );
    and g18001 ( n33558 , n34330 , n17079 );
    or g18002 ( n31778 , n20043 , n1165 );
    and g18003 ( n31049 , n34299 , n11131 );
    or g18004 ( n10779 , n4878 , n30737 );
    and g18005 ( n118 , n14856 , n24139 );
    or g18006 ( n14491 , n17568 , n13315 );
    or g18007 ( n10270 , n30312 , n12465 );
    or g18008 ( n10811 , n28856 , n4175 );
    not g18009 ( n4260 , n26192 );
    or g18010 ( n12403 , n5335 , n11470 );
    or g18011 ( n6243 , n35625 , n14505 );
    or g18012 ( n4270 , n29868 , n21644 );
    nor g18013 ( n6883 , n9658 , n19077 );
    or g18014 ( n1146 , n10427 , n32608 );
    or g18015 ( n30824 , n15412 , n13768 );
    or g18016 ( n5390 , n28169 , n14620 );
    or g18017 ( n22407 , n4750 , n4203 );
    or g18018 ( n28132 , n31647 , n20866 );
    not g18019 ( n9896 , n1528 );
    or g18020 ( n11516 , n24411 , n27447 );
    xnor g18021 ( n14435 , n14578 , n15403 );
    nor g18022 ( n5543 , n35927 , n26539 );
    and g18023 ( n33844 , n8296 , n14493 );
    or g18024 ( n21290 , n5335 , n1428 );
    xnor g18025 ( n26532 , n12024 , n31289 );
    xnor g18026 ( n26247 , n23926 , n7443 );
    xnor g18027 ( n8935 , n22429 , n17115 );
    xnor g18028 ( n7322 , n4724 , n32408 );
    or g18029 ( n26870 , n4878 , n3121 );
    xnor g18030 ( n30053 , n7739 , n28716 );
    and g18031 ( n13210 , n35233 , n1788 );
    nor g18032 ( n29014 , n29876 , n415 );
    and g18033 ( n15128 , n3164 , n34136 );
    buf g18034 ( n714 , n19120 );
    xor g18035 ( n23838 , n2006 , n32527 );
    or g18036 ( n5813 , n15413 , n11518 );
    xnor g18037 ( n23203 , n30061 , n35826 );
    or g18038 ( n9282 , n31949 , n3694 );
    or g18039 ( n33394 , n19551 , n33142 );
    xnor g18040 ( n21083 , n19420 , n4288 );
    or g18041 ( n11138 , n6696 , n26002 );
    and g18042 ( n10433 , n35583 , n19006 );
    or g18043 ( n8786 , n32857 , n6829 );
    or g18044 ( n13216 , n33914 , n11495 );
    and g18045 ( n8255 , n4618 , n32794 );
    and g18046 ( n24027 , n33087 , n4518 );
    and g18047 ( n21106 , n5714 , n20555 );
    or g18048 ( n9171 , n27891 , n32071 );
    and g18049 ( n2458 , n5053 , n26397 );
    xnor g18050 ( n16984 , n27422 , n34396 );
    and g18051 ( n9360 , n31859 , n35610 );
    or g18052 ( n34574 , n29410 , n2683 );
    and g18053 ( n32632 , n17365 , n26917 );
    or g18054 ( n7738 , n32918 , n12596 );
    or g18055 ( n27926 , n21107 , n19722 );
    or g18056 ( n29114 , n30192 , n20177 );
    not g18057 ( n7267 , n33186 );
    xnor g18058 ( n7157 , n30587 , n20458 );
    and g18059 ( n15559 , n22122 , n5673 );
    xnor g18060 ( n7441 , n5166 , n25174 );
    xnor g18061 ( n23662 , n4369 , n24332 );
    and g18062 ( n5275 , n22779 , n14527 );
    xnor g18063 ( n14358 , n15294 , n17450 );
    or g18064 ( n13026 , n6823 , n34656 );
    or g18065 ( n24269 , n1565 , n17354 );
    xnor g18066 ( n28020 , n4494 , n15546 );
    and g18067 ( n29624 , n1444 , n26663 );
    or g18068 ( n7570 , n31799 , n15841 );
    xnor g18069 ( n35268 , n26313 , n19551 );
    not g18070 ( n33398 , n29839 );
    or g18071 ( n1394 , n5335 , n31775 );
    xnor g18072 ( n31061 , n35383 , n33952 );
    or g18073 ( n16597 , n4631 , n11258 );
    or g18074 ( n27270 , n9895 , n32991 );
    buf g18075 ( n35748 , n19058 );
    and g18076 ( n10430 , n13063 , n30726 );
    or g18077 ( n29528 , n18527 , n5868 );
    or g18078 ( n30330 , n4878 , n3349 );
    xnor g18079 ( n17370 , n32995 , n33312 );
    nor g18080 ( n27694 , n2956 , n30753 );
    or g18081 ( n2497 , n17858 , n6288 );
    or g18082 ( n24515 , n4370 , n31134 );
    and g18083 ( n16207 , n29758 , n36037 );
    xnor g18084 ( n2824 , n8494 , n16445 );
    or g18085 ( n17825 , n29588 , n35476 );
    not g18086 ( n28787 , n19939 );
    buf g18087 ( n12596 , n32837 );
    xnor g18088 ( n34333 , n15960 , n15993 );
    nor g18089 ( n15297 , n32095 , n29952 );
    and g18090 ( n11442 , n718 , n20163 );
    not g18091 ( n23279 , n9686 );
    or g18092 ( n30355 , n12014 , n30476 );
    and g18093 ( n31622 , n33406 , n14606 );
    xnor g18094 ( n21049 , n19850 , n22720 );
    xnor g18095 ( n5940 , n31356 , n5287 );
    or g18096 ( n21678 , n20437 , n5457 );
    or g18097 ( n25989 , n2735 , n17233 );
    and g18098 ( n20403 , n32779 , n28447 );
    and g18099 ( n26037 , n10677 , n18172 );
    or g18100 ( n30035 , n13594 , n824 );
    or g18101 ( n8072 , n5959 , n15109 );
    xnor g18102 ( n5248 , n33291 , n31484 );
    and g18103 ( n3962 , n23808 , n10766 );
    and g18104 ( n10986 , n10649 , n4795 );
    not g18105 ( n9767 , n31411 );
    and g18106 ( n27250 , n9041 , n19912 );
    and g18107 ( n25476 , n22656 , n12045 );
    or g18108 ( n98 , n15886 , n33044 );
    or g18109 ( n11669 , n19363 , n22961 );
    xnor g18110 ( n5086 , n16692 , n32584 );
    or g18111 ( n3880 , n35301 , n35764 );
    xor g18112 ( n8345 , n8533 , n29823 );
    or g18113 ( n29313 , n10894 , n32469 );
    or g18114 ( n30946 , n1805 , n2119 );
    and g18115 ( n3477 , n4573 , n26492 );
    xnor g18116 ( n27718 , n15055 , n11455 );
    and g18117 ( n21954 , n4329 , n18262 );
    not g18118 ( n12747 , n2317 );
    xnor g18119 ( n25746 , n34224 , n9793 );
    xnor g18120 ( n20956 , n660 , n29630 );
    xnor g18121 ( n13848 , n12677 , n32095 );
    and g18122 ( n12557 , n2324 , n644 );
    and g18123 ( n30683 , n10482 , n1262 );
    or g18124 ( n22919 , n20453 , n27625 );
    and g18125 ( n19955 , n2938 , n10130 );
    or g18126 ( n16241 , n18507 , n31055 );
    nor g18127 ( n19188 , n29713 , n23744 );
    xnor g18128 ( n32561 , n3362 , n35927 );
    or g18129 ( n4902 , n27158 , n26365 );
    or g18130 ( n31859 , n5773 , n1942 );
    or g18131 ( n22095 , n12669 , n30431 );
    and g18132 ( n32275 , n2297 , n10496 );
    and g18133 ( n6658 , n17231 , n23129 );
    or g18134 ( n16441 , n362 , n15363 );
    and g18135 ( n25418 , n3172 , n18420 );
    or g18136 ( n26795 , n5582 , n31656 );
    not g18137 ( n8725 , n5411 );
    buf g18138 ( n21579 , n15638 );
    xnor g18139 ( n13622 , n8650 , n29571 );
    or g18140 ( n3700 , n3070 , n20690 );
    xnor g18141 ( n161 , n21488 , n3205 );
    and g18142 ( n25753 , n19031 , n24128 );
    or g18143 ( n12094 , n15886 , n35028 );
    or g18144 ( n9976 , n13672 , n32329 );
    and g18145 ( n27257 , n18663 , n36083 );
    or g18146 ( n28040 , n25026 , n24710 );
    xnor g18147 ( n27548 , n34324 , n24069 );
    xnor g18148 ( n23415 , n26688 , n13983 );
    or g18149 ( n31385 , n25081 , n35228 );
    xnor g18150 ( n11953 , n15904 , n21907 );
    and g18151 ( n20368 , n10836 , n5787 );
    or g18152 ( n22674 , n5702 , n32808 );
    or g18153 ( n12295 , n18279 , n27687 );
    not g18154 ( n21524 , n289 );
    or g18155 ( n14392 , n2399 , n17046 );
    xnor g18156 ( n20700 , n9206 , n16593 );
    xnor g18157 ( n16143 , n35627 , n13224 );
    or g18158 ( n20908 , n1256 , n30204 );
    or g18159 ( n13519 , n5777 , n3922 );
    xnor g18160 ( n34220 , n7355 , n17408 );
    xnor g18161 ( n823 , n3569 , n6179 );
    nor g18162 ( n6894 , n8255 , n24666 );
    or g18163 ( n33322 , n27326 , n31359 );
    nor g18164 ( n35427 , n18344 , n7448 );
    or g18165 ( n31495 , n34662 , n19069 );
    or g18166 ( n13927 , n20764 , n19952 );
    nor g18167 ( n23284 , n35917 , n34014 );
    and g18168 ( n18555 , n25018 , n12806 );
    and g18169 ( n11781 , n19765 , n12604 );
    not g18170 ( n1862 , n7026 );
    xnor g18171 ( n15964 , n15904 , n33467 );
    nor g18172 ( n24622 , n6282 , n17067 );
    and g18173 ( n24697 , n34886 , n24152 );
    and g18174 ( n20462 , n30651 , n14948 );
    not g18175 ( n29533 , n30607 );
    xnor g18176 ( n4651 , n25645 , n31799 );
    and g18177 ( n7262 , n18568 , n6805 );
    not g18178 ( n13187 , n12238 );
    or g18179 ( n22930 , n17189 , n34537 );
    or g18180 ( n16020 , n32401 , n24427 );
    or g18181 ( n14096 , n19367 , n4691 );
    or g18182 ( n16335 , n6434 , n19435 );
    and g18183 ( n28560 , n12256 , n32085 );
    or g18184 ( n28127 , n34676 , n20308 );
    or g18185 ( n26694 , n27803 , n34472 );
    not g18186 ( n7672 , n15886 );
    or g18187 ( n16190 , n3205 , n31124 );
    xnor g18188 ( n32672 , n34496 , n25360 );
    and g18189 ( n18087 , n12786 , n7606 );
    or g18190 ( n20533 , n25227 , n10289 );
    and g18191 ( n31175 , n18890 , n32318 );
    and g18192 ( n26157 , n20078 , n35479 );
    not g18193 ( n24193 , n4201 );
    or g18194 ( n34956 , n32095 , n10737 );
    or g18195 ( n29744 , n6743 , n26630 );
    xnor g18196 ( n14591 , n34149 , n18582 );
    or g18197 ( n2135 , n3149 , n1763 );
    not g18198 ( n19265 , n6257 );
    xnor g18199 ( n10160 , n23120 , n15577 );
    and g18200 ( n1541 , n4349 , n24615 );
    or g18201 ( n25027 , n940 , n13307 );
    xnor g18202 ( n36053 , n28637 , n7511 );
    xnor g18203 ( n11623 , n16752 , n9789 );
    or g18204 ( n13265 , n5835 , n8789 );
    or g18205 ( n7743 , n26623 , n11601 );
    xnor g18206 ( n2906 , n19578 , n30563 );
    and g18207 ( n32466 , n12761 , n28284 );
    or g18208 ( n22601 , n9786 , n20300 );
    xnor g18209 ( n19147 , n1352 , n16175 );
    or g18210 ( n19116 , n9789 , n632 );
    or g18211 ( n874 , n9658 , n12331 );
    and g18212 ( n33850 , n25562 , n16203 );
    or g18213 ( n19083 , n22291 , n16925 );
    xnor g18214 ( n21277 , n5464 , n928 );
    or g18215 ( n34911 , n8270 , n20817 );
    or g18216 ( n22207 , n12756 , n12910 );
    or g18217 ( n25802 , n9244 , n14397 );
    or g18218 ( n9620 , n7498 , n578 );
    nor g18219 ( n7304 , n15886 , n14648 );
    or g18220 ( n35567 , n13903 , n17612 );
    or g18221 ( n17084 , n33438 , n27963 );
    or g18222 ( n23445 , n22932 , n17354 );
    or g18223 ( n29286 , n27283 , n28240 );
    or g18224 ( n14692 , n30742 , n566 );
    xnor g18225 ( n23194 , n26376 , n15185 );
    and g18226 ( n2470 , n10756 , n18041 );
    or g18227 ( n34101 , n10324 , n4595 );
    and g18228 ( n7523 , n30263 , n26130 );
    nor g18229 ( n25550 , n3069 , n11757 );
    and g18230 ( n4042 , n24028 , n19278 );
    or g18231 ( n4781 , n31446 , n22783 );
    or g18232 ( n11235 , n30556 , n9555 );
    xnor g18233 ( n17696 , n28365 , n32095 );
    xnor g18234 ( n31211 , n32571 , n11167 );
    buf g18235 ( n17046 , n22793 );
    nor g18236 ( n10391 , n4960 , n19429 );
    or g18237 ( n12097 , n7615 , n11460 );
    and g18238 ( n10363 , n3724 , n1468 );
    not g18239 ( n28669 , n7588 );
    and g18240 ( n4444 , n15410 , n17547 );
    not g18241 ( n34425 , n16502 );
    nor g18242 ( n22611 , n4651 , n27793 );
    xnor g18243 ( n31771 , n5071 , n11471 );
    or g18244 ( n24224 , n9511 , n16688 );
    xnor g18245 ( n11413 , n2506 , n10894 );
    or g18246 ( n31404 , n8190 , n3239 );
    or g18247 ( n32854 , n20910 , n14847 );
    or g18248 ( n33267 , n32885 , n8446 );
    or g18249 ( n22420 , n3017 , n12326 );
    or g18250 ( n33817 , n31364 , n19690 );
    or g18251 ( n1457 , n12000 , n9009 );
    xnor g18252 ( n32577 , n3949 , n4288 );
    or g18253 ( n34466 , n7785 , n27671 );
    or g18254 ( n19849 , n3205 , n31586 );
    not g18255 ( n811 , n30155 );
    and g18256 ( n29294 , n17251 , n32424 );
    or g18257 ( n8426 , n28348 , n2823 );
    or g18258 ( n16801 , n31138 , n10760 );
    nor g18259 ( n8926 , n4288 , n12269 );
    and g18260 ( n33961 , n7114 , n5318 );
    and g18261 ( n5066 , n33026 , n25443 );
    xnor g18262 ( n2022 , n17458 , n10894 );
    xnor g18263 ( n26641 , n11953 , n23385 );
    or g18264 ( n27301 , n21421 , n19241 );
    nor g18265 ( n7602 , n4288 , n26968 );
    xnor g18266 ( n4429 , n13944 , n2260 );
    or g18267 ( n29667 , n146 , n34484 );
    or g18268 ( n19831 , n8456 , n12067 );
    or g18269 ( n35184 , n14424 , n22241 );
    and g18270 ( n29138 , n3082 , n27235 );
    and g18271 ( n25236 , n10859 , n25707 );
    xnor g18272 ( n13843 , n28016 , n22472 );
    xnor g18273 ( n12616 , n15853 , n25439 );
    nor g18274 ( n13834 , n23604 , n20983 );
    nor g18275 ( n9970 , n7727 , n25507 );
    or g18276 ( n33366 , n1572 , n21977 );
    nor g18277 ( n24922 , n29713 , n30027 );
    or g18278 ( n16706 , n33109 , n20318 );
    and g18279 ( n30492 , n250 , n5141 );
    and g18280 ( n32730 , n9705 , n18747 );
    xnor g18281 ( n27067 , n23334 , n17568 );
    or g18282 ( n6142 , n5436 , n27624 );
    or g18283 ( n34896 , n4694 , n6553 );
    or g18284 ( n8370 , n11190 , n32667 );
    nor g18285 ( n11820 , n31215 , n1118 );
    xnor g18286 ( n29475 , n35712 , n17568 );
    xnor g18287 ( n32285 , n13260 , n11876 );
    or g18288 ( n30283 , n35706 , n20840 );
    nor g18289 ( n23538 , n28819 , n30608 );
    or g18290 ( n35501 , n32530 , n27704 );
    or g18291 ( n19747 , n29197 , n2613 );
    or g18292 ( n21534 , n17008 , n6900 );
    or g18293 ( n35599 , n34632 , n17964 );
    or g18294 ( n17620 , n22838 , n2932 );
    or g18295 ( n31665 , n30553 , n32243 );
    xnor g18296 ( n19407 , n33150 , n35165 );
    not g18297 ( n22084 , n19520 );
    or g18298 ( n21140 , n24332 , n12164 );
    and g18299 ( n28804 , n31667 , n6271 );
    or g18300 ( n10704 , n29887 , n18255 );
    or g18301 ( n15670 , n18551 , n7423 );
    or g18302 ( n34861 , n12093 , n11703 );
    xnor g18303 ( n27884 , n1676 , n17306 );
    and g18304 ( n19249 , n21933 , n31192 );
    nor g18305 ( n9109 , n32857 , n18181 );
    or g18306 ( n18817 , n32041 , n21061 );
    not g18307 ( n26877 , n7540 );
    and g18308 ( n20879 , n21558 , n9209 );
    or g18309 ( n8835 , n28566 , n6288 );
    or g18310 ( n26478 , n7314 , n9546 );
    or g18311 ( n9733 , n15755 , n17337 );
    and g18312 ( n33918 , n3549 , n9622 );
    and g18313 ( n6318 , n22562 , n26326 );
    xnor g18314 ( n32479 , n15914 , n26877 );
    or g18315 ( n30301 , n24371 , n16840 );
    or g18316 ( n31733 , n9376 , n28089 );
    or g18317 ( n32013 , n24665 , n3274 );
    or g18318 ( n8360 , n14552 , n14841 );
    and g18319 ( n4610 , n34185 , n30626 );
    and g18320 ( n24458 , n6631 , n34495 );
    not g18321 ( n26543 , n16691 );
    and g18322 ( n8349 , n31730 , n4358 );
    and g18323 ( n33762 , n28969 , n21720 );
    or g18324 ( n34809 , n18950 , n30449 );
    or g18325 ( n4155 , n2663 , n11258 );
    or g18326 ( n7085 , n4180 , n7293 );
    not g18327 ( n33896 , n11996 );
    or g18328 ( n9444 , n1192 , n12879 );
    and g18329 ( n11640 , n3666 , n15525 );
    or g18330 ( n22034 , n21758 , n7417 );
    and g18331 ( n35649 , n8757 , n17021 );
    xnor g18332 ( n2274 , n24211 , n12201 );
    or g18333 ( n19312 , n2435 , n27963 );
    xnor g18334 ( n5391 , n14536 , n32191 );
    or g18335 ( n27205 , n30933 , n34493 );
    nor g18336 ( n11916 , n4962 , n24132 );
    and g18337 ( n16888 , n22963 , n29857 );
    and g18338 ( n7481 , n1182 , n9283 );
    and g18339 ( n13350 , n1388 , n19072 );
    xnor g18340 ( n31897 , n16915 , n25174 );
    nor g18341 ( n10961 , n15226 , n16348 );
    and g18342 ( n7982 , n29961 , n7234 );
    and g18343 ( n14171 , n28132 , n29999 );
    or g18344 ( n24876 , n13192 , n29872 );
    xnor g18345 ( n5075 , n26755 , n34219 );
    or g18346 ( n3935 , n8374 , n26306 );
    nor g18347 ( n617 , n31799 , n18300 );
    xnor g18348 ( n13479 , n7242 , n1950 );
    and g18349 ( n17481 , n3339 , n16509 );
    and g18350 ( n1567 , n33361 , n5805 );
    xnor g18351 ( n10832 , n35605 , n10894 );
    and g18352 ( n33376 , n11140 , n25614 );
    or g18353 ( n19705 , n5772 , n3631 );
    and g18354 ( n27185 , n1163 , n1501 );
    or g18355 ( n33954 , n30233 , n10634 );
    or g18356 ( n4290 , n28581 , n27973 );
    or g18357 ( n15029 , n12025 , n3761 );
    xnor g18358 ( n29696 , n21112 , n3222 );
    or g18359 ( n28256 , n29486 , n12622 );
    and g18360 ( n5720 , n27162 , n5762 );
    xnor g18361 ( n13637 , n18508 , n19652 );
    xnor g18362 ( n25076 , n25382 , n30667 );
    and g18363 ( n19091 , n4815 , n15453 );
    or g18364 ( n18386 , n28091 , n9555 );
    or g18365 ( n17069 , n14552 , n12606 );
    or g18366 ( n445 , n33646 , n11577 );
    and g18367 ( n26705 , n31471 , n21612 );
    and g18368 ( n14726 , n33293 , n31330 );
    or g18369 ( n32681 , n13731 , n27511 );
    and g18370 ( n33388 , n4886 , n13068 );
    and g18371 ( n20155 , n24762 , n10956 );
    xnor g18372 ( n1719 , n5111 , n10894 );
    and g18373 ( n13877 , n10741 , n14014 );
    nor g18374 ( n11266 , n23604 , n101 );
    or g18375 ( n3828 , n32469 , n34484 );
    or g18376 ( n24838 , n20425 , n31755 );
    or g18377 ( n27957 , n30600 , n21644 );
    not g18378 ( n14145 , n18445 );
    xnor g18379 ( n43 , n29243 , n31073 );
    buf g18380 ( n20576 , n28404 );
    or g18381 ( n32405 , n32857 , n25589 );
    nor g18382 ( n31922 , n11241 , n19125 );
    or g18383 ( n17484 , n4142 , n12146 );
    or g18384 ( n480 , n20918 , n29735 );
    and g18385 ( n14077 , n23797 , n16483 );
    not g18386 ( n34532 , n9957 );
    or g18387 ( n11861 , n1109 , n25648 );
    or g18388 ( n24429 , n31947 , n18542 );
    or g18389 ( n14007 , n4915 , n34557 );
    or g18390 ( n13607 , n26585 , n6374 );
    xnor g18391 ( n19434 , n5921 , n4758 );
    xnor g18392 ( n35381 , n6368 , n3651 );
    or g18393 ( n1238 , n27456 , n8723 );
    and g18394 ( n26090 , n4110 , n2298 );
    or g18395 ( n15573 , n22396 , n20932 );
    xnor g18396 ( n7722 , n29748 , n13254 );
    buf g18397 ( n30431 , n21418 );
    or g18398 ( n13531 , n26921 , n7417 );
    or g18399 ( n15470 , n22149 , n3188 );
    not g18400 ( n16501 , n34415 );
    or g18401 ( n19007 , n19621 , n33889 );
    and g18402 ( n11849 , n21766 , n2557 );
    and g18403 ( n22268 , n30288 , n25872 );
    nor g18404 ( n32189 , n8231 , n25153 );
    or g18405 ( n10338 , n4960 , n5884 );
    and g18406 ( n2633 , n22204 , n36066 );
    nor g18407 ( n31517 , n8958 , n24827 );
    and g18408 ( n8238 , n30394 , n16721 );
    or g18409 ( n24604 , n7084 , n6374 );
    and g18410 ( n16608 , n2638 , n20984 );
    xnor g18411 ( n11928 , n32103 , n31776 );
    and g18412 ( n32278 , n904 , n18464 );
    not g18413 ( n12535 , n19559 );
    xnor g18414 ( n30836 , n18438 , n10975 );
    or g18415 ( n25480 , n4316 , n949 );
    or g18416 ( n12700 , n23997 , n27645 );
    or g18417 ( n4385 , n24229 , n1454 );
    or g18418 ( n30378 , n8238 , n32329 );
    not g18419 ( n281 , n1950 );
    and g18420 ( n6296 , n15550 , n21692 );
    xnor g18421 ( n28971 , n16168 , n22291 );
    xnor g18422 ( n1986 , n3278 , n30742 );
    xnor g18423 ( n30934 , n811 , n24332 );
    or g18424 ( n21399 , n34258 , n20797 );
    nor g18425 ( n22118 , n10989 , n7306 );
    or g18426 ( n16070 , n4277 , n21977 );
    or g18427 ( n3617 , n1546 , n32959 );
    and g18428 ( n914 , n27200 , n12403 );
    or g18429 ( n11362 , n25299 , n26002 );
    or g18430 ( n19436 , n10894 , n12171 );
    xnor g18431 ( n3149 , n2447 , n33969 );
    not g18432 ( n28846 , n4878 );
    or g18433 ( n11012 , n1802 , n21155 );
    or g18434 ( n10104 , n8432 , n17451 );
    or g18435 ( n9216 , n418 , n2955 );
    or g18436 ( n18903 , n30742 , n12621 );
    or g18437 ( n6404 , n21788 , n5972 );
    nor g18438 ( n35033 , n3205 , n35923 );
    or g18439 ( n23097 , n27712 , n15439 );
    not g18440 ( n96 , n24371 );
    or g18441 ( n2715 , n28617 , n30732 );
    not g18442 ( n31765 , n9192 );
    or g18443 ( n33110 , n23026 , n1511 );
    xnor g18444 ( n9804 , n22527 , n9840 );
    and g18445 ( n25842 , n28381 , n17948 );
    and g18446 ( n7546 , n22878 , n11686 );
    nor g18447 ( n7789 , n30742 , n19259 );
    xnor g18448 ( n30816 , n36034 , n19814 );
    xnor g18449 ( n9064 , n13407 , n25304 );
    and g18450 ( n22829 , n31889 , n16931 );
    or g18451 ( n20535 , n23787 , n4648 );
    and g18452 ( n8710 , n17254 , n21183 );
    not g18453 ( n27952 , n15260 );
    and g18454 ( n19609 , n15078 , n28501 );
    or g18455 ( n31880 , n3966 , n16516 );
    xnor g18456 ( n29218 , n32401 , n24427 );
    or g18457 ( n2983 , n13284 , n9601 );
    and g18458 ( n11156 , n25901 , n7980 );
    xnor g18459 ( n17378 , n4935 , n28873 );
    or g18460 ( n22360 , n2539 , n15538 );
    or g18461 ( n10705 , n25165 , n7726 );
    xnor g18462 ( n1134 , n10454 , n20173 );
    xnor g18463 ( n9919 , n23213 , n9658 );
    or g18464 ( n10029 , n33065 , n30023 );
    nor g18465 ( n13238 , n17568 , n24646 );
    or g18466 ( n5497 , n1376 , n26292 );
    not g18467 ( n27601 , n31825 );
    nor g18468 ( n15050 , n29713 , n2608 );
    or g18469 ( n29511 , n18503 , n27704 );
    nor g18470 ( n12396 , n7814 , n30656 );
    not g18471 ( n2878 , n19851 );
    and g18472 ( n8288 , n12479 , n18806 );
    or g18473 ( n30857 , n25177 , n8203 );
    or g18474 ( n1623 , n35229 , n28191 );
    or g18475 ( n27931 , n9379 , n34484 );
    or g18476 ( n11278 , n25035 , n21956 );
    or g18477 ( n18833 , n32332 , n20747 );
    xnor g18478 ( n6588 , n26293 , n15381 );
    or g18479 ( n12750 , n31426 , n12596 );
    and g18480 ( n33901 , n25017 , n24812 );
    and g18481 ( n130 , n10032 , n30916 );
    not g18482 ( n11483 , n9969 );
    or g18483 ( n29221 , n18700 , n15256 );
    or g18484 ( n34307 , n3795 , n16919 );
    not g18485 ( n5149 , n19551 );
    or g18486 ( n26387 , n3113 , n6075 );
    and g18487 ( n9995 , n32756 , n4021 );
    xnor g18488 ( n21355 , n21227 , n27226 );
    and g18489 ( n6692 , n26714 , n32355 );
    or g18490 ( n35081 , n11233 , n9675 );
    not g18491 ( n22047 , n27060 );
    xnor g18492 ( n31878 , n6371 , n31477 );
    or g18493 ( n1303 , n18404 , n15295 );
    or g18494 ( n9754 , n830 , n29570 );
    or g18495 ( n16601 , n29075 , n34600 );
    or g18496 ( n35721 , n2928 , n10960 );
    or g18497 ( n2156 , n21230 , n32182 );
    xnor g18498 ( n9038 , n3191 , n27226 );
    or g18499 ( n18328 , n8432 , n35514 );
    and g18500 ( n8624 , n6202 , n19804 );
    buf g18501 ( n11996 , n27006 );
    or g18502 ( n22122 , n8948 , n25255 );
    and g18503 ( n33513 , n24425 , n7855 );
    and g18504 ( n14340 , n32651 , n14647 );
    or g18505 ( n27975 , n34242 , n8371 );
    or g18506 ( n29789 , n20406 , n11593 );
    nor g18507 ( n6325 , n11190 , n25799 );
    or g18508 ( n31540 , n4960 , n36038 );
    or g18509 ( n28352 , n13634 , n11518 );
    or g18510 ( n11279 , n28425 , n1909 );
    and g18511 ( n15230 , n20544 , n22872 );
    and g18512 ( n29847 , n7628 , n4465 );
    and g18513 ( n28174 , n11069 , n30920 );
    nor g18514 ( n15984 , n19551 , n8642 );
    xnor g18515 ( n21539 , n20746 , n7931 );
    and g18516 ( n2270 , n8760 , n24906 );
    or g18517 ( n8047 , n31272 , n20328 );
    xnor g18518 ( n31580 , n29 , n8256 );
    xnor g18519 ( n33040 , n24613 , n4962 );
    not g18520 ( n17591 , n2648 );
    not g18521 ( n16263 , n24226 );
    or g18522 ( n32470 , n19551 , n8489 );
    xnor g18523 ( n10370 , n21106 , n31215 );
    or g18524 ( n1775 , n4911 , n23717 );
    or g18525 ( n4699 , n1076 , n4912 );
    or g18526 ( n10796 , n28971 , n21010 );
    and g18527 ( n15298 , n18229 , n32868 );
    xnor g18528 ( n11331 , n5029 , n6821 );
    or g18529 ( n20182 , n4335 , n33034 );
    or g18530 ( n19754 , n26968 , n8255 );
    xnor g18531 ( n33943 , n12753 , n830 );
    xnor g18532 ( n19057 , n31884 , n2057 );
    and g18533 ( n18954 , n3401 , n7010 );
    or g18534 ( n31008 , n23403 , n34084 );
    xnor g18535 ( n19932 , n32876 , n10637 );
    and g18536 ( n7906 , n8143 , n21761 );
    and g18537 ( n1900 , n7128 , n35081 );
    and g18538 ( n22774 , n4483 , n11937 );
    xnor g18539 ( n23202 , n7265 , n21651 );
    and g18540 ( n29917 , n3717 , n8560 );
    or g18541 ( n10078 , n25792 , n23093 );
    or g18542 ( n15560 , n24956 , n16854 );
    and g18543 ( n35985 , n10000 , n10014 );
    or g18544 ( n22032 , n18754 , n10161 );
    or g18545 ( n26527 , n21513 , n8064 );
    or g18546 ( n18320 , n9222 , n20780 );
    xnor g18547 ( n19985 , n10091 , n23112 );
    or g18548 ( n18093 , n15254 , n12428 );
    or g18549 ( n11710 , n23604 , n2361 );
    or g18550 ( n5211 , n28441 , n10762 );
    xnor g18551 ( n3171 , n24410 , n1725 );
    or g18552 ( n8806 , n20504 , n25831 );
    or g18553 ( n19303 , n3121 , n14285 );
    xnor g18554 ( n29683 , n22559 , n21665 );
    or g18555 ( n12561 , n8484 , n19952 );
    and g18556 ( n6336 , n26142 , n28543 );
    not g18557 ( n15178 , n3744 );
    xnor g18558 ( n13225 , n19535 , n27711 );
    or g18559 ( n35277 , n27698 , n20776 );
    not g18560 ( n19730 , n16922 );
    buf g18561 ( n29592 , n14627 );
    and g18562 ( n28613 , n16227 , n22185 );
    xnor g18563 ( n6367 , n6527 , n12652 );
    buf g18564 ( n31411 , n32983 );
    nor g18565 ( n798 , n32095 , n11147 );
    not g18566 ( n8493 , n7588 );
    xnor g18567 ( n30189 , n35067 , n32091 );
    or g18568 ( n21506 , n32584 , n9309 );
    xnor g18569 ( n18150 , n6192 , n12456 );
    or g18570 ( n8145 , n12883 , n33416 );
    and g18571 ( n8684 , n35146 , n6834 );
    and g18572 ( n4893 , n29768 , n5638 );
    or g18573 ( n11236 , n9940 , n30419 );
    xnor g18574 ( n20503 , n29008 , n26892 );
    or g18575 ( n17925 , n33195 , n23852 );
    and g18576 ( n29036 , n18713 , n49 );
    or g18577 ( n17326 , n31220 , n35748 );
    or g18578 ( n32070 , n24332 , n7699 );
    and g18579 ( n6680 , n28264 , n12892 );
    and g18580 ( n18487 , n22525 , n2846 );
    xnor g18581 ( n31216 , n31863 , n22291 );
    and g18582 ( n17616 , n4861 , n26375 );
    nor g18583 ( n7090 , n25584 , n11074 );
    and g18584 ( n16632 , n20970 , n27315 );
    nor g18585 ( n2405 , n35728 , n4271 );
    and g18586 ( n20498 , n29227 , n35094 );
    and g18587 ( n31131 , n30487 , n34944 );
    or g18588 ( n2485 , n10585 , n16734 );
    or g18589 ( n17512 , n29839 , n3143 );
    not g18590 ( n2613 , n714 );
    xnor g18591 ( n15399 , n14882 , n19551 );
    or g18592 ( n26204 , n15119 , n31514 );
    or g18593 ( n7839 , n31000 , n34086 );
    or g18594 ( n9650 , n17957 , n763 );
    or g18595 ( n19905 , n9658 , n16616 );
    or g18596 ( n6056 , n17940 , n24554 );
    nor g18597 ( n2999 , n29279 , n24030 );
    or g18598 ( n15680 , n32061 , n25786 );
    or g18599 ( n35588 , n9768 , n26105 );
    or g18600 ( n31366 , n24332 , n23621 );
    xnor g18601 ( n20919 , n17404 , n17150 );
    xnor g18602 ( n7822 , n17788 , n9793 );
    xnor g18603 ( n31772 , n29488 , n31215 );
    or g18604 ( n29192 , n16424 , n8203 );
    or g18605 ( n11356 , n22106 , n25940 );
    or g18606 ( n24067 , n4983 , n4532 );
    nor g18607 ( n24085 , n35927 , n20030 );
    or g18608 ( n625 , n20455 , n24672 );
    and g18609 ( n35259 , n26318 , n35628 );
    or g18610 ( n35544 , n18419 , n25648 );
    not g18611 ( n10153 , n14136 );
    and g18612 ( n4135 , n30464 , n32084 );
    xnor g18613 ( n267 , n12352 , n4804 );
    and g18614 ( n19524 , n12893 , n24620 );
    and g18615 ( n32485 , n4248 , n15598 );
    xnor g18616 ( n27874 , n11314 , n31559 );
    xnor g18617 ( n25609 , n9673 , n1950 );
    or g18618 ( n9908 , n23704 , n14746 );
    or g18619 ( n2452 , n4288 , n28051 );
    xnor g18620 ( n29123 , n14801 , n30013 );
    and g18621 ( n9443 , n18036 , n5898 );
    or g18622 ( n18461 , n4962 , n11901 );
    xnor g18623 ( n14879 , n13567 , n15886 );
    and g18624 ( n27741 , n2088 , n32108 );
    xnor g18625 ( n12355 , n13509 , n4960 );
    and g18626 ( n7589 , n12716 , n9616 );
    and g18627 ( n1795 , n25935 , n16546 );
    and g18628 ( n32811 , n18479 , n5551 );
    and g18629 ( n25987 , n35155 , n28040 );
    and g18630 ( n33458 , n8957 , n23291 );
    xnor g18631 ( n9132 , n623 , n9658 );
    and g18632 ( n32795 , n20295 , n19948 );
    and g18633 ( n8658 , n30935 , n16560 );
    or g18634 ( n16739 , n24438 , n14671 );
    or g18635 ( n9343 , n17751 , n7941 );
    or g18636 ( n18879 , n34867 , n18845 );
    xnor g18637 ( n28399 , n15272 , n3222 );
    or g18638 ( n21383 , n16243 , n21237 );
    or g18639 ( n1543 , n8550 , n32087 );
    and g18640 ( n29020 , n19517 , n18129 );
    and g18641 ( n4009 , n19660 , n14843 );
    and g18642 ( n13603 , n17714 , n23738 );
    or g18643 ( n6745 , n34450 , n10577 );
    or g18644 ( n21103 , n2344 , n26468 );
    xnor g18645 ( n21107 , n12632 , n31028 );
    xnor g18646 ( n27487 , n28902 , n29322 );
    or g18647 ( n24980 , n33858 , n17434 );
    nor g18648 ( n11489 , n9658 , n23914 );
    nor g18649 ( n24179 , n23081 , n21514 );
    or g18650 ( n14593 , n13316 , n28120 );
    and g18651 ( n18722 , n3664 , n35156 );
    or g18652 ( n2368 , n15886 , n13270 );
    or g18653 ( n153 , n4534 , n32039 );
    xnor g18654 ( n6615 , n17907 , n1950 );
    or g18655 ( n20891 , n12830 , n35935 );
    xnor g18656 ( n15285 , n24044 , n33551 );
    xnor g18657 ( n23946 , n27615 , n25174 );
    and g18658 ( n5690 , n25601 , n33866 );
    and g18659 ( n22571 , n28681 , n28976 );
    xnor g18660 ( n5740 , n34096 , n9658 );
    and g18661 ( n33227 , n17085 , n7132 );
    or g18662 ( n104 , n29318 , n11977 );
    or g18663 ( n26685 , n13325 , n29195 );
    or g18664 ( n333 , n2312 , n22530 );
    nor g18665 ( n19618 , n15886 , n22766 );
    or g18666 ( n31462 , n34173 , n15145 );
    xnor g18667 ( n22821 , n12385 , n25638 );
    or g18668 ( n13323 , n32629 , n21691 );
    not g18669 ( n12132 , n2099 );
    xnor g18670 ( n31361 , n695 , n4130 );
    xnor g18671 ( n34517 , n6660 , n31799 );
    xnor g18672 ( n19041 , n19914 , n27291 );
    nor g18673 ( n6933 , n4962 , n22672 );
    not g18674 ( n23288 , n31289 );
    or g18675 ( n21238 , n14142 , n11295 );
    and g18676 ( n30485 , n24236 , n226 );
    not g18677 ( n31753 , n22291 );
    xnor g18678 ( n5446 , n519 , n35097 );
    and g18679 ( n14682 , n16009 , n35751 );
    or g18680 ( n13873 , n14459 , n32071 );
    xnor g18681 ( n30821 , n32844 , n34648 );
    not g18682 ( n16141 , n23604 );
    xnor g18683 ( n25131 , n22975 , n9658 );
    or g18684 ( n8859 , n9831 , n33435 );
    and g18685 ( n25705 , n31369 , n3953 );
    or g18686 ( n26820 , n10894 , n14589 );
    xnor g18687 ( n9870 , n980 , n4878 );
    and g18688 ( n29866 , n1164 , n26495 );
    or g18689 ( n4374 , n35424 , n19490 );
    and g18690 ( n7187 , n21777 , n25014 );
    or g18691 ( n9632 , n33407 , n8392 );
    not g18692 ( n29492 , n11926 );
    xnor g18693 ( n1304 , n23387 , n4288 );
    or g18694 ( n31373 , n12744 , n12112 );
    xnor g18695 ( n27346 , n10809 , n32043 );
    or g18696 ( n18346 , n19794 , n13307 );
    xnor g18697 ( n786 , n9578 , n8300 );
    xnor g18698 ( n33341 , n27880 , n31056 );
    xnor g18699 ( n19950 , n15822 , n7547 );
    or g18700 ( n28185 , n33729 , n22613 );
    xnor g18701 ( n22114 , n13037 , n4288 );
    xnor g18702 ( n10884 , n27456 , n31272 );
    or g18703 ( n2158 , n21052 , n11601 );
    or g18704 ( n15223 , n25633 , n11218 );
    buf g18705 ( n35402 , n11785 );
    and g18706 ( n18173 , n4584 , n9416 );
    and g18707 ( n19787 , n27012 , n1746 );
    xnor g18708 ( n33276 , n4308 , n5335 );
    xnor g18709 ( n16669 , n36068 , n27812 );
    or g18710 ( n21976 , n11958 , n2660 );
    or g18711 ( n27906 , n19984 , n13368 );
    xnor g18712 ( n2356 , n32326 , n19872 );
    or g18713 ( n5825 , n29183 , n5752 );
    xnor g18714 ( n16026 , n27237 , n1645 );
    xnor g18715 ( n25275 , n33319 , n34738 );
    not g18716 ( n24262 , n32054 );
    xnor g18717 ( n4701 , n13521 , n7352 );
    xnor g18718 ( n35345 , n35584 , n28852 );
    or g18719 ( n7384 , n24675 , n20840 );
    or g18720 ( n24917 , n31105 , n16464 );
    and g18721 ( n5423 , n4850 , n15071 );
    or g18722 ( n1760 , n30756 , n20811 );
    and g18723 ( n25976 , n21066 , n18249 );
    or g18724 ( n16317 , n5067 , n22843 );
    xnor g18725 ( n18232 , n25774 , n34247 );
    not g18726 ( n18533 , n12428 );
    and g18727 ( n7677 , n10330 , n33801 );
    xnor g18728 ( n11525 , n9829 , n28885 );
    xnor g18729 ( n7269 , n3819 , n9905 );
    or g18730 ( n9061 , n18202 , n13011 );
    xnor g18731 ( n26651 , n644 , n2324 );
    xnor g18732 ( n6196 , n21015 , n16361 );
    or g18733 ( n17687 , n25870 , n17385 );
    or g18734 ( n2322 , n32584 , n12053 );
    and g18735 ( n28181 , n22741 , n21552 );
    and g18736 ( n36033 , n6198 , n20730 );
    and g18737 ( n10076 , n34345 , n31680 );
    or g18738 ( n8546 , n32584 , n21373 );
    and g18739 ( n17957 , n33074 , n21589 );
    or g18740 ( n13694 , n14631 , n35657 );
    xnor g18741 ( n14329 , n6979 , n4878 );
    and g18742 ( n11170 , n33005 , n23758 );
    or g18743 ( n22706 , n2468 , n17829 );
    or g18744 ( n25503 , n30362 , n13057 );
    or g18745 ( n35601 , n22291 , n3448 );
    or g18746 ( n27204 , n9075 , n25567 );
    xnor g18747 ( n15903 , n30682 , n4919 );
    or g18748 ( n591 , n32699 , n15109 );
    or g18749 ( n20508 , n12338 , n27527 );
    xnor g18750 ( n35671 , n14953 , n21659 );
    xnor g18751 ( n15966 , n13728 , n17042 );
    xnor g18752 ( n12372 , n33043 , n17898 );
    or g18753 ( n14930 , n11565 , n25123 );
    or g18754 ( n33290 , n9247 , n22312 );
    or g18755 ( n487 , n21866 , n16762 );
    and g18756 ( n30091 , n34966 , n13809 );
    or g18757 ( n20233 , n29851 , n13250 );
    xnor g18758 ( n10621 , n30022 , n7686 );
    not g18759 ( n437 , n12622 );
    nor g18760 ( n28635 , n9658 , n5379 );
    or g18761 ( n35835 , n25696 , n31549 );
    or g18762 ( n34675 , n11834 , n2490 );
    or g18763 ( n9533 , n17537 , n16464 );
    and g18764 ( n12775 , n32273 , n4331 );
    or g18765 ( n10592 , n25531 , n8840 );
    nor g18766 ( n6289 , n23604 , n27231 );
    xnor g18767 ( n10966 , n4009 , n3205 );
    or g18768 ( n7605 , n22195 , n35572 );
    or g18769 ( n20083 , n8432 , n21638 );
    or g18770 ( n10515 , n16780 , n34727 );
    and g18771 ( n12067 , n2378 , n29471 );
    or g18772 ( n451 , n22574 , n25831 );
    and g18773 ( n15804 , n14869 , n26243 );
    xnor g18774 ( n17858 , n15698 , n17932 );
    xnor g18775 ( n2865 , n30090 , n23977 );
    xnor g18776 ( n28231 , n14324 , n241 );
    or g18777 ( n24452 , n23151 , n3611 );
    xnor g18778 ( n4748 , n5446 , n11660 );
    or g18779 ( n3401 , n8579 , n4016 );
    not g18780 ( n18017 , n16064 );
    or g18781 ( n1040 , n17095 , n15497 );
    or g18782 ( n9766 , n12545 , n20308 );
    or g18783 ( n5916 , n8257 , n2119 );
    or g18784 ( n32551 , n30486 , n12596 );
    or g18785 ( n26064 , n14987 , n20358 );
    or g18786 ( n11380 , n4423 , n20308 );
    or g18787 ( n24657 , n22291 , n1983 );
    and g18788 ( n25032 , n23191 , n21674 );
    xnor g18789 ( n6757 , n34837 , n10061 );
    or g18790 ( n7438 , n3946 , n1649 );
    or g18791 ( n4084 , n34663 , n32505 );
    or g18792 ( n33442 , n13937 , n18471 );
    and g18793 ( n34280 , n15564 , n33973 );
    not g18794 ( n33541 , n7540 );
    and g18795 ( n5826 , n27832 , n16993 );
    xnor g18796 ( n15476 , n20242 , n32268 );
    or g18797 ( n26885 , n24922 , n15870 );
    and g18798 ( n28909 , n24318 , n7351 );
    or g18799 ( n28153 , n1185 , n21042 );
    nor g18800 ( n10040 , n16620 , n5095 );
    xnor g18801 ( n29501 , n35017 , n11190 );
    and g18802 ( n29661 , n35779 , n3728 );
    xnor g18803 ( n10559 , n26368 , n28959 );
    xnor g18804 ( n29500 , n5553 , n28890 );
    not g18805 ( n31820 , n36042 );
    and g18806 ( n19971 , n26463 , n1976 );
    xnor g18807 ( n22889 , n23427 , n25086 );
    or g18808 ( n23780 , n30515 , n30204 );
    xnor g18809 ( n18886 , n24363 , n4288 );
    or g18810 ( n35287 , n3362 , n6024 );
    xnor g18811 ( n6200 , n32466 , n25174 );
    or g18812 ( n22332 , n23502 , n33205 );
    and g18813 ( n34746 , n32988 , n14212 );
    or g18814 ( n13060 , n24279 , n11712 );
    not g18815 ( n381 , n25130 );
    xnor g18816 ( n8612 , n20328 , n31272 );
    nor g18817 ( n24406 , n3205 , n7894 );
    or g18818 ( n12177 , n1950 , n21703 );
    or g18819 ( n11103 , n8708 , n406 );
    not g18820 ( n14754 , n20721 );
    nor g18821 ( n30995 , n34312 , n9856 );
    or g18822 ( n21047 , n11251 , n7212 );
    or g18823 ( n15013 , n18205 , n10572 );
    or g18824 ( n15550 , n32674 , n21002 );
    xnor g18825 ( n17331 , n19211 , n8107 );
    xnor g18826 ( n3913 , n5765 , n23288 );
    or g18827 ( n3390 , n23218 , n2241 );
    xnor g18828 ( n27208 , n4391 , n12595 );
    xnor g18829 ( n1848 , n8776 , n25602 );
    and g18830 ( n13810 , n20243 , n23239 );
    or g18831 ( n15556 , n30117 , n16659 );
    and g18832 ( n19999 , n5285 , n35442 );
    xnor g18833 ( n24151 , n33965 , n14129 );
    or g18834 ( n727 , n7429 , n6819 );
    or g18835 ( n8952 , n34568 , n6212 );
    and g18836 ( n2630 , n8248 , n33946 );
    not g18837 ( n26779 , n16922 );
    xnor g18838 ( n13686 , n12407 , n28222 );
    xnor g18839 ( n33641 , n23337 , n21922 );
    or g18840 ( n20967 , n27291 , n21510 );
    xnor g18841 ( n2320 , n31421 , n26459 );
    xnor g18842 ( n34974 , n13955 , n23355 );
    or g18843 ( n27547 , n10506 , n4478 );
    xnor g18844 ( n34327 , n16215 , n24856 );
    and g18845 ( n6645 , n25675 , n19364 );
    not g18846 ( n16060 , n25451 );
    not g18847 ( n1592 , n25602 );
    and g18848 ( n396 , n13223 , n14139 );
    and g18849 ( n4057 , n6824 , n2183 );
    nor g18850 ( n16510 , n9580 , n16855 );
    and g18851 ( n5894 , n33270 , n26011 );
    xnor g18852 ( n2776 , n32445 , n7945 );
    or g18853 ( n3519 , n16119 , n28295 );
    and g18854 ( n29716 , n20380 , n33321 );
    xnor g18855 ( n20438 , n11313 , n8423 );
    and g18856 ( n16943 , n28258 , n19165 );
    nor g18857 ( n31290 , n23261 , n5284 );
    xnor g18858 ( n20445 , n24906 , n8760 );
    xnor g18859 ( n31973 , n8212 , n23729 );
    xnor g18860 ( n13783 , n33185 , n9658 );
    or g18861 ( n26278 , n1173 , n35920 );
    or g18862 ( n26534 , n23311 , n34249 );
    xnor g18863 ( n17132 , n29911 , n573 );
    nor g18864 ( n26440 , n1950 , n1446 );
    and g18865 ( n16505 , n27714 , n19825 );
    xnor g18866 ( n25400 , n3652 , n10894 );
    or g18867 ( n29292 , n31746 , n27437 );
    or g18868 ( n11869 , n6482 , n35271 );
    or g18869 ( n28496 , n35408 , n35141 );
    and g18870 ( n15003 , n4294 , n34131 );
    or g18871 ( n4859 , n30452 , n8924 );
    or g18872 ( n6944 , n24371 , n22321 );
    and g18873 ( n10450 , n22326 , n15492 );
    or g18874 ( n7426 , n9665 , n8090 );
    or g18875 ( n18952 , n7568 , n29393 );
    and g18876 ( n12808 , n31942 , n33145 );
    xnor g18877 ( n21421 , n27238 , n33796 );
    and g18878 ( n24744 , n17689 , n12924 );
    or g18879 ( n2967 , n1736 , n22501 );
    or g18880 ( n29196 , n9593 , n27642 );
    nor g18881 ( n33009 , n3222 , n36042 );
    or g18882 ( n4413 , n19284 , n16594 );
    nor g18883 ( n33505 , n22548 , n13141 );
    or g18884 ( n35169 , n8432 , n1919 );
    and g18885 ( n15700 , n13832 , n34957 );
    or g18886 ( n21458 , n3064 , n30287 );
    xnor g18887 ( n3702 , n11141 , n2078 );
    or g18888 ( n9436 , n6363 , n34360 );
    and g18889 ( n17988 , n5445 , n25697 );
    xnor g18890 ( n8343 , n28211 , n11190 );
    or g18891 ( n7922 , n25918 , n21080 );
    or g18892 ( n10904 , n10653 , n16296 );
    or g18893 ( n23041 , n25602 , n7302 );
    and g18894 ( n29381 , n6005 , n17452 );
    or g18895 ( n30669 , n32955 , n32114 );
    or g18896 ( n13813 , n7140 , n26818 );
    and g18897 ( n21998 , n26144 , n32033 );
    nor g18898 ( n32141 , n8068 , n24955 );
    or g18899 ( n34106 , n9723 , n19561 );
    or g18900 ( n24799 , n19467 , n26697 );
    or g18901 ( n23858 , n6592 , n32313 );
    nor g18902 ( n24518 , n12323 , n16568 );
    xnor g18903 ( n3467 , n5045 , n31289 );
    or g18904 ( n32426 , n26754 , n22682 );
    or g18905 ( n9709 , n26897 , n22950 );
    or g18906 ( n3030 , n1950 , n13629 );
    and g18907 ( n6133 , n33502 , n3894 );
    or g18908 ( n26456 , n2831 , n11780 );
    nor g18909 ( n35780 , n17568 , n7470 );
    or g18910 ( n34721 , n10350 , n19403 );
    nor g18911 ( n3432 , n8743 , n28493 );
    xnor g18912 ( n22618 , n35921 , n11472 );
    not g18913 ( n29560 , n26263 );
    or g18914 ( n25790 , n1093 , n16457 );
    or g18915 ( n4019 , n24607 , n29629 );
    nor g18916 ( n28606 , n26867 , n6017 );
    buf g18917 ( n28668 , n3842 );
    xnor g18918 ( n26162 , n19988 , n29917 );
    xnor g18919 ( n4973 , n4468 , n27226 );
    xnor g18920 ( n35962 , n11415 , n4288 );
    nor g18921 ( n3998 , n24721 , n18115 );
    xnor g18922 ( n361 , n33 , n21807 );
    or g18923 ( n6253 , n25607 , n32071 );
    or g18924 ( n5812 , n32486 , n26468 );
    or g18925 ( n22752 , n8337 , n2104 );
    and g18926 ( n34968 , n22551 , n14088 );
    or g18927 ( n28271 , n505 , n4490 );
    xnor g18928 ( n26765 , n31760 , n6473 );
    or g18929 ( n2267 , n10427 , n22241 );
    xnor g18930 ( n32065 , n28752 , n28939 );
    and g18931 ( n20521 , n32022 , n31503 );
    and g18932 ( n9214 , n22606 , n31528 );
    nor g18933 ( n3786 , n10207 , n30365 );
    not g18934 ( n24666 , n22980 );
    and g18935 ( n24790 , n13087 , n27670 );
    or g18936 ( n11025 , n25174 , n30399 );
    and g18937 ( n4918 , n5266 , n9582 );
    and g18938 ( n4551 , n3828 , n24122 );
    or g18939 ( n22695 , n28199 , n13453 );
    and g18940 ( n32669 , n20757 , n6997 );
    or g18941 ( n14131 , n16031 , n13307 );
    or g18942 ( n31491 , n3609 , n676 );
    or g18943 ( n10476 , n26985 , n1251 );
    xnor g18944 ( n9206 , n762 , n15623 );
    or g18945 ( n14212 , n9789 , n15358 );
    xnor g18946 ( n12191 , n2489 , n32584 );
    and g18947 ( n1812 , n30344 , n7722 );
    or g18948 ( n5870 , n29867 , n4230 );
    buf g18949 ( n12950 , n5713 );
    or g18950 ( n4234 , n27864 , n16033 );
    xnor g18951 ( n31486 , n29800 , n31215 );
    or g18952 ( n8675 , n19243 , n35973 );
    or g18953 ( n32762 , n18201 , n19421 );
    or g18954 ( n4936 , n3205 , n3637 );
    xnor g18955 ( n31105 , n12681 , n4477 );
    or g18956 ( n35102 , n4044 , n25255 );
    or g18957 ( n25522 , n19248 , n17974 );
    or g18958 ( n26081 , n22492 , n28904 );
    or g18959 ( n2206 , n28176 , n12428 );
    and g18960 ( n28397 , n29838 , n32426 );
    and g18961 ( n29132 , n3333 , n29901 );
    or g18962 ( n36082 , n7540 , n18130 );
    xnor g18963 ( n19923 , n22968 , n17751 );
    and g18964 ( n16724 , n33718 , n18434 );
    not g18965 ( n32386 , n20393 );
    xnor g18966 ( n35607 , n26995 , n4288 );
    xnor g18967 ( n21409 , n14439 , n32093 );
    or g18968 ( n23932 , n20490 , n34472 );
    nor g18969 ( n4282 , n31215 , n30297 );
    xnor g18970 ( n29 , n24777 , n35756 );
    nor g18971 ( n6518 , n33025 , n20172 );
    xnor g18972 ( n6646 , n34726 , n35957 );
    or g18973 ( n16040 , n20651 , n17337 );
    or g18974 ( n15425 , n15048 , n27405 );
    or g18975 ( n765 , n13775 , n12879 );
    or g18976 ( n19157 , n15286 , n32797 );
    and g18977 ( n25282 , n35774 , n33383 );
    not g18978 ( n35909 , n4288 );
    xnor g18979 ( n28423 , n27680 , n30687 );
    or g18980 ( n13040 , n27806 , n28440 );
    xnor g18981 ( n18532 , n22292 , n11190 );
    not g18982 ( n21054 , n22980 );
    xnor g18983 ( n2311 , n3259 , n2792 );
    and g18984 ( n35967 , n12114 , n26509 );
    or g18985 ( n11434 , n16330 , n9675 );
    xnor g18986 ( n9530 , n12251 , n16019 );
    or g18987 ( n4512 , n35484 , n31498 );
    and g18988 ( n15004 , n15806 , n5002 );
    or g18989 ( n2286 , n17545 , n28668 );
    or g18990 ( n29131 , n10078 , n19402 );
    xnor g18991 ( n4951 , n5066 , n31289 );
    or g18992 ( n22333 , n33536 , n3979 );
    or g18993 ( n385 , n11190 , n5079 );
    and g18994 ( n17244 , n7174 , n10671 );
    or g18995 ( n33922 , n15397 , n20300 );
    or g18996 ( n30998 , n11735 , n22160 );
    or g18997 ( n8388 , n6226 , n25629 );
    nor g18998 ( n5512 , n32715 , n2647 );
    xnor g18999 ( n18057 , n26093 , n10272 );
    and g19000 ( n9953 , n10715 , n2942 );
    xnor g19001 ( n21949 , n18694 , n29713 );
    and g19002 ( n14506 , n24960 , n16236 );
    or g19003 ( n25535 , n35108 , n27447 );
    and g19004 ( n17976 , n3915 , n27377 );
    or g19005 ( n12246 , n9618 , n6553 );
    or g19006 ( n17418 , n35637 , n10762 );
    or g19007 ( n11580 , n27565 , n11789 );
    or g19008 ( n17880 , n17568 , n17435 );
    or g19009 ( n30941 , n16219 , n14918 );
    and g19010 ( n15895 , n12592 , n30191 );
    and g19011 ( n11621 , n1405 , n16748 );
    or g19012 ( n29863 , n29271 , n22736 );
    not g19013 ( n9006 , n25761 );
    and g19014 ( n26004 , n9 , n28101 );
    or g19015 ( n2414 , n16922 , n23894 );
    or g19016 ( n20186 , n18466 , n28248 );
    not g19017 ( n1145 , n9789 );
    xnor g19018 ( n5366 , n28199 , n13453 );
    xnor g19019 ( n10996 , n28546 , n19992 );
    xnor g19020 ( n27411 , n337 , n23032 );
    or g19021 ( n22729 , n32533 , n10289 );
    xnor g19022 ( n5363 , n20983 , n32588 );
    or g19023 ( n2617 , n32095 , n26556 );
    xnor g19024 ( n7245 , n28830 , n7540 );
    xnor g19025 ( n27263 , n34665 , n16017 );
    or g19026 ( n22053 , n830 , n6051 );
    nor g19027 ( n19409 , n7509 , n16649 );
    or g19028 ( n13793 , n11046 , n6828 );
    or g19029 ( n3755 , n24702 , n35306 );
    or g19030 ( n21548 , n30742 , n4740 );
    nor g19031 ( n5865 , n16799 , n28072 );
    xnor g19032 ( n25821 , n1718 , n4288 );
    or g19033 ( n224 , n14220 , n19095 );
    and g19034 ( n5976 , n25221 , n24854 );
    or g19035 ( n21348 , n24528 , n25447 );
    and g19036 ( n8105 , n30758 , n5083 );
    or g19037 ( n2810 , n18266 , n2712 );
    or g19038 ( n8097 , n23830 , n4917 );
    and g19039 ( n19028 , n34506 , n447 );
    and g19040 ( n18761 , n26790 , n10338 );
    xnor g19041 ( n12570 , n21465 , n8432 );
    or g19042 ( n34339 , n13676 , n27728 );
    xnor g19043 ( n13854 , n7379 , n5887 );
    and g19044 ( n26447 , n35646 , n7938 );
    nor g19045 ( n23390 , n27388 , n21149 );
    and g19046 ( n15766 , n26405 , n27017 );
    or g19047 ( n25621 , n17568 , n13186 );
    and g19048 ( n12860 , n15001 , n12144 );
    xnor g19049 ( n28982 , n2361 , n1884 );
    xnor g19050 ( n36022 , n29396 , n22295 );
    or g19051 ( n9777 , n35534 , n22641 );
    and g19052 ( n24559 , n23617 , n30259 );
    or g19053 ( n29641 , n12044 , n31563 );
    or g19054 ( n25736 , n8692 , n26002 );
    and g19055 ( n29967 , n28918 , n23803 );
    not g19056 ( n29871 , n29839 );
    and g19057 ( n28429 , n10232 , n12572 );
    or g19058 ( n14492 , n5899 , n20692 );
    xnor g19059 ( n8742 , n33485 , n11455 );
    nor g19060 ( n993 , n31559 , n8488 );
    and g19061 ( n28855 , n20323 , n15725 );
    or g19062 ( n4671 , n3036 , n4716 );
    not g19063 ( n4077 , n32451 );
    or g19064 ( n19315 , n970 , n23209 );
    not g19065 ( n11708 , n2414 );
    and g19066 ( n35846 , n23356 , n34498 );
    or g19067 ( n7910 , n13628 , n17531 );
    or g19068 ( n6750 , n4282 , n29687 );
    or g19069 ( n3060 , n15886 , n23369 );
    and g19070 ( n20504 , n17137 , n35068 );
    and g19071 ( n21964 , n15666 , n4593 );
    xnor g19072 ( n782 , n6572 , n22291 );
    xnor g19073 ( n15930 , n26074 , n9793 );
    xnor g19074 ( n15684 , n30855 , n32943 );
    not g19075 ( n11174 , n9385 );
    or g19076 ( n32440 , n10508 , n16139 );
    or g19077 ( n16999 , n2776 , n16345 );
    and g19078 ( n6480 , n20160 , n69 );
    or g19079 ( n28824 , n5568 , n7673 );
    xnor g19080 ( n32527 , n12601 , n4878 );
    and g19081 ( n14671 , n18630 , n3650 );
    xnor g19082 ( n10471 , n6388 , n31056 );
    and g19083 ( n25912 , n32910 , n25790 );
    and g19084 ( n22514 , n34624 , n14455 );
    or g19085 ( n33594 , n30881 , n2340 );
    or g19086 ( n18786 , n16585 , n34923 );
    or g19087 ( n25692 , n14127 , n31055 );
    nor g19088 ( n10478 , n34111 , n22270 );
    xnor g19089 ( n12084 , n350 , n103 );
    xnor g19090 ( n2750 , n14108 , n4288 );
    and g19091 ( n26973 , n8079 , n21376 );
    or g19092 ( n13985 , n20920 , n14812 );
    or g19093 ( n16962 , n24852 , n5343 );
    xnor g19094 ( n9243 , n6999 , n25817 );
    xnor g19095 ( n13461 , n6482 , n35271 );
    or g19096 ( n17689 , n28229 , n24672 );
    xnor g19097 ( n13276 , n35740 , n2734 );
    or g19098 ( n18396 , n4179 , n26931 );
    xnor g19099 ( n32264 , n25118 , n4492 );
    or g19100 ( n3855 , n16852 , n28837 );
    nor g19101 ( n15043 , n2800 , n5635 );
    and g19102 ( n31114 , n7849 , n12952 );
    or g19103 ( n18036 , n15432 , n26121 );
    and g19104 ( n699 , n19075 , n81 );
    and g19105 ( n2606 , n3527 , n9980 );
    and g19106 ( n12016 , n18860 , n27345 );
    and g19107 ( n30089 , n31512 , n24794 );
    or g19108 ( n11090 , n9649 , n24672 );
    and g19109 ( n348 , n18335 , n26617 );
    not g19110 ( n1982 , n25873 );
    or g19111 ( n30788 , n9623 , n27053 );
    xnor g19112 ( n8713 , n2136 , n32584 );
    and g19113 ( n20094 , n16550 , n29245 );
    or g19114 ( n32611 , n20980 , n1688 );
    or g19115 ( n904 , n12819 , n9629 );
    or g19116 ( n10105 , n17751 , n12949 );
    or g19117 ( n3625 , n24476 , n16797 );
    or g19118 ( n1284 , n33300 , n6374 );
    not g19119 ( n18148 , n2247 );
    or g19120 ( n9826 , n4560 , n140 );
    or g19121 ( n18215 , n7540 , n11055 );
    and g19122 ( n17308 , n9532 , n23083 );
    or g19123 ( n12184 , n9179 , n11578 );
    xnor g19124 ( n6034 , n31475 , n22111 );
    xnor g19125 ( n9235 , n26232 , n32717 );
    or g19126 ( n933 , n29259 , n24180 );
    xnor g19127 ( n35257 , n7857 , n11455 );
    and g19128 ( n14882 , n193 , n14010 );
    or g19129 ( n21093 , n4433 , n12622 );
    or g19130 ( n8962 , n27291 , n5961 );
    xnor g19131 ( n30429 , n35884 , n6163 );
    xnor g19132 ( n13024 , n6287 , n480 );
    not g19133 ( n17628 , n4725 );
    and g19134 ( n3005 , n31529 , n6177 );
    xnor g19135 ( n28706 , n30099 , n12912 );
    xnor g19136 ( n1441 , n21255 , n33271 );
    or g19137 ( n32595 , n31799 , n20244 );
    and g19138 ( n8954 , n35350 , n35790 );
    xnor g19139 ( n16258 , n11091 , n35927 );
    or g19140 ( n33260 , n15464 , n32476 );
    and g19141 ( n20490 , n34133 , n34526 );
    or g19142 ( n1047 , n13890 , n30190 );
    or g19143 ( n34169 , n22291 , n30149 );
    and g19144 ( n33647 , n34843 , n18646 );
    or g19145 ( n11230 , n22272 , n21002 );
    or g19146 ( n33893 , n14214 , n17612 );
    and g19147 ( n7511 , n224 , n14228 );
    not g19148 ( n106 , n12428 );
    and g19149 ( n34192 , n23104 , n10704 );
    xnor g19150 ( n213 , n24435 , n1884 );
    not g19151 ( n31699 , n22471 );
    not g19152 ( n25401 , n31692 );
    and g19153 ( n2842 , n11412 , n8860 );
    and g19154 ( n22274 , n25396 , n27852 );
    and g19155 ( n12674 , n17145 , n25242 );
    and g19156 ( n35744 , n27659 , n14934 );
    xnor g19157 ( n14117 , n29549 , n12402 );
    and g19158 ( n19333 , n23598 , n22588 );
    or g19159 ( n33583 , n33332 , n28455 );
    and g19160 ( n20676 , n6195 , n28144 );
    or g19161 ( n34387 , n19295 , n1849 );
    not g19162 ( n1458 , n24371 );
    nor g19163 ( n13623 , n17568 , n12514 );
    buf g19164 ( n31134 , n6075 );
    buf g19165 ( n21042 , n2005 );
    not g19166 ( n9439 , n7817 );
    or g19167 ( n12478 , n20444 , n27704 );
    buf g19168 ( n2384 , n9297 );
    or g19169 ( n23782 , n22229 , n31758 );
    or g19170 ( n33534 , n35324 , n4254 );
    nor g19171 ( n8789 , n30026 , n26108 );
    and g19172 ( n25729 , n10811 , n25822 );
    not g19173 ( n20467 , n2029 );
    and g19174 ( n31964 , n29424 , n2373 );
    and g19175 ( n19144 , n34564 , n21135 );
    buf g19176 ( n36000 , n33200 );
    or g19177 ( n26135 , n32584 , n17642 );
    or g19178 ( n4832 , n24477 , n29562 );
    and g19179 ( n12529 , n2828 , n29960 );
    not g19180 ( n34551 , n2417 );
    not g19181 ( n24397 , n36075 );
    not g19182 ( n11187 , n2172 );
    and g19183 ( n17657 , n27964 , n36012 );
    or g19184 ( n1164 , n27479 , n19728 );
    and g19185 ( n31032 , n7156 , n1348 );
    xnor g19186 ( n8969 , n1332 , n27630 );
    and g19187 ( n10335 , n25039 , n6623 );
    not g19188 ( n1411 , n1528 );
    and g19189 ( n32138 , n27421 , n31513 );
    or g19190 ( n35710 , n8491 , n18691 );
    nor g19191 ( n6101 , n14670 , n2801 );
    or g19192 ( n6902 , n17971 , n15439 );
    or g19193 ( n4786 , n8661 , n5607 );
    and g19194 ( n6498 , n26401 , n23951 );
    xnor g19195 ( n31439 , n35042 , n9658 );
    or g19196 ( n26679 , n26321 , n11703 );
    and g19197 ( n745 , n34247 , n25774 );
    or g19198 ( n32307 , n3222 , n7621 );
    or g19199 ( n9492 , n21197 , n15109 );
    or g19200 ( n29228 , n7629 , n8122 );
    nor g19201 ( n14461 , n4962 , n791 );
    and g19202 ( n30405 , n19775 , n34490 );
    or g19203 ( n29170 , n24626 , n19421 );
    xnor g19204 ( n14225 , n15829 , n1950 );
    or g19205 ( n3154 , n33981 , n32505 );
    and g19206 ( n8286 , n22848 , n4173 );
    or g19207 ( n26603 , n35249 , n14918 );
    nor g19208 ( n31650 , n5287 , n28315 );
    xnor g19209 ( n30064 , n418 , n25174 );
    or g19210 ( n33755 , n23604 , n1616 );
    nor g19211 ( n23660 , n10894 , n15540 );
    or g19212 ( n13700 , n17419 , n29872 );
    or g19213 ( n16864 , n19118 , n33034 );
    nor g19214 ( n34892 , n1178 , n9440 );
    xnor g19215 ( n32129 , n9964 , n1018 );
    or g19216 ( n17813 , n21889 , n3842 );
    and g19217 ( n14589 , n9027 , n9276 );
    not g19218 ( n8702 , n30459 );
    or g19219 ( n269 , n28076 , n14719 );
    or g19220 ( n24081 , n26262 , n25940 );
    or g19221 ( n13616 , n817 , n13891 );
    xnor g19222 ( n2113 , n35371 , n830 );
    xnor g19223 ( n14897 , n4587 , n4960 );
    not g19224 ( n1534 , n26352 );
    or g19225 ( n30211 , n32844 , n34648 );
    not g19226 ( n3424 , n34477 );
    xnor g19227 ( n18758 , n21193 , n19551 );
    or g19228 ( n3597 , n13992 , n4515 );
    or g19229 ( n32776 , n32095 , n28365 );
    or g19230 ( n17277 , n35282 , n25567 );
    nor g19231 ( n10681 , n29713 , n4835 );
    or g19232 ( n8240 , n15253 , n27030 );
    or g19233 ( n32805 , n13615 , n33310 );
    nor g19234 ( n16567 , n28394 , n21792 );
    or g19235 ( n14529 , n2091 , n29393 );
    xnor g19236 ( n27891 , n35118 , n14215 );
    not g19237 ( n9955 , n8637 );
    not g19238 ( n14954 , n32168 );
    nor g19239 ( n33061 , n13957 , n16649 );
    and g19240 ( n14739 , n16268 , n19960 );
    or g19241 ( n33525 , n21094 , n18810 );
    nor g19242 ( n6604 , n16620 , n34976 );
    or g19243 ( n24122 , n26784 , n17612 );
    xnor g19244 ( n22906 , n23485 , n5335 );
    or g19245 ( n21740 , n15403 , n5022 );
    xnor g19246 ( n10460 , n30398 , n22323 );
    or g19247 ( n34460 , n28320 , n29379 );
    or g19248 ( n27223 , n14000 , n26365 );
    and g19249 ( n13578 , n34010 , n11913 );
    or g19250 ( n31222 , n31272 , n8695 );
    or g19251 ( n257 , n24759 , n29592 );
    and g19252 ( n5209 , n4894 , n11353 );
    xnor g19253 ( n19677 , n1045 , n18851 );
    not g19254 ( n35337 , n6021 );
    or g19255 ( n23230 , n2106 , n19105 );
    and g19256 ( n27820 , n32789 , n20499 );
    xnor g19257 ( n28171 , n8889 , n25022 );
    or g19258 ( n1562 , n29478 , n4595 );
    xnor g19259 ( n14500 , n24132 , n4962 );
    or g19260 ( n620 , n35386 , n3694 );
    or g19261 ( n19020 , n19273 , n26919 );
    or g19262 ( n1481 , n11637 , n6632 );
    or g19263 ( n18497 , n4162 , n12622 );
    and g19264 ( n27563 , n14297 , n679 );
    or g19265 ( n30513 , n21583 , n6106 );
    xnor g19266 ( n34080 , n24344 , n25180 );
    and g19267 ( n10528 , n19672 , n20359 );
    or g19268 ( n7487 , n36090 , n23626 );
    xnor g19269 ( n12282 , n21875 , n7309 );
    or g19270 ( n28773 , n8049 , n31749 );
    and g19271 ( n30158 , n14362 , n4848 );
    or g19272 ( n6672 , n9793 , n35907 );
    xnor g19273 ( n30160 , n31807 , n2253 );
    or g19274 ( n30709 , n22966 , n34688 );
    not g19275 ( n15044 , n35443 );
    or g19276 ( n31635 , n7304 , n29023 );
    and g19277 ( n30448 , n1461 , n19161 );
    and g19278 ( n6153 , n9425 , n11561 );
    not g19279 ( n12826 , n11046 );
    or g19280 ( n14572 , n34512 , n16762 );
    or g19281 ( n34306 , n1467 , n1756 );
    xnor g19282 ( n32877 , n22038 , n3688 );
    not g19283 ( n19945 , n30204 );
    or g19284 ( n19966 , n1950 , n8317 );
    xnor g19285 ( n16119 , n10596 , n4962 );
    nor g19286 ( n20953 , n27910 , n34723 );
    nor g19287 ( n27698 , n5335 , n25104 );
    and g19288 ( n12480 , n31666 , n17019 );
    not g19289 ( n32837 , n13216 );
    or g19290 ( n10507 , n29413 , n19223 );
    xnor g19291 ( n21980 , n24229 , n19551 );
    or g19292 ( n23110 , n8432 , n27978 );
    not g19293 ( n7653 , n12393 );
    or g19294 ( n14243 , n14817 , n10432 );
    and g19295 ( n31966 , n17418 , n4261 );
    or g19296 ( n13653 , n30337 , n11977 );
    xnor g19297 ( n19059 , n14485 , n32584 );
    or g19298 ( n7476 , n3521 , n14554 );
    or g19299 ( n108 , n30977 , n10765 );
    or g19300 ( n34920 , n35607 , n10484 );
    xnor g19301 ( n6653 , n1616 , n8582 );
    or g19302 ( n34884 , n4222 , n17629 );
    xnor g19303 ( n1993 , n30399 , n25174 );
    xnor g19304 ( n29969 , n32385 , n4758 );
    nor g19305 ( n20170 , n11190 , n33053 );
    or g19306 ( n22928 , n12476 , n24355 );
    xnor g19307 ( n34301 , n35870 , n32038 );
    xnor g19308 ( n24275 , n19051 , n13743 );
    or g19309 ( n8135 , n34034 , n5752 );
    and g19310 ( n370 , n4051 , n34748 );
    and g19311 ( n10997 , n24884 , n23841 );
    xnor g19312 ( n16024 , n30102 , n3840 );
    or g19313 ( n28998 , n1950 , n13407 );
    or g19314 ( n14114 , n31056 , n5684 );
    or g19315 ( n18859 , n7967 , n16464 );
    or g19316 ( n15898 , n22742 , n31134 );
    or g19317 ( n15259 , n20973 , n6340 );
    xnor g19318 ( n18029 , n35493 , n25686 );
    xnor g19319 ( n31449 , n26985 , n1251 );
    xnor g19320 ( n15957 , n30809 , n5335 );
    xnor g19321 ( n15696 , n24765 , n25174 );
    xnor g19322 ( n19140 , n14907 , n11891 );
    and g19323 ( n23627 , n4278 , n13439 );
    not g19324 ( n28503 , n1989 );
    xnor g19325 ( n9122 , n14682 , n7698 );
    xnor g19326 ( n25607 , n18462 , n2580 );
    and g19327 ( n7495 , n12233 , n30443 );
    or g19328 ( n34401 , n1877 , n16919 );
    nor g19329 ( n20279 , n7540 , n12685 );
    or g19330 ( n7370 , n1940 , n9112 );
    xnor g19331 ( n3676 , n10405 , n34745 );
    or g19332 ( n4261 , n18534 , n30646 );
    xnor g19333 ( n3959 , n28784 , n23259 );
    not g19334 ( n10038 , n13906 );
    xnor g19335 ( n12548 , n31060 , n3864 );
    or g19336 ( n24060 , n19932 , n28404 );
    or g19337 ( n12241 , n17568 , n31619 );
    or g19338 ( n5757 , n5154 , n25648 );
    and g19339 ( n30161 , n21994 , n15995 );
    not g19340 ( n11161 , n16223 );
    or g19341 ( n16375 , n3222 , n35827 );
    or g19342 ( n23730 , n12166 , n11774 );
    nor g19343 ( n19686 , n35817 , n3683 );
    or g19344 ( n28505 , n32137 , n24548 );
    and g19345 ( n9918 , n3690 , n33452 );
    or g19346 ( n14552 , n33588 , n18798 );
    xnor g19347 ( n20324 , n10595 , n4055 );
    or g19348 ( n30103 , n17568 , n20453 );
    or g19349 ( n31713 , n26842 , n27728 );
    not g19350 ( n35570 , n2535 );
    or g19351 ( n7640 , n29420 , n3979 );
    not g19352 ( n10191 , n29203 );
    or g19353 ( n21128 , n30373 , n34484 );
    and g19354 ( n1736 , n29723 , n34947 );
    xnor g19355 ( n10640 , n29531 , n29713 );
    or g19356 ( n26841 , n9332 , n22682 );
    and g19357 ( n10367 , n28723 , n18285 );
    and g19358 ( n31550 , n4866 , n24074 );
    xnor g19359 ( n14496 , n16230 , n30742 );
    and g19360 ( n7646 , n26014 , n21407 );
    and g19361 ( n31133 , n26223 , n26901 );
    buf g19362 ( n15290 , n1183 );
    xnor g19363 ( n13617 , n7050 , n31799 );
    or g19364 ( n12116 , n29884 , n31715 );
    or g19365 ( n16063 , n13695 , n35043 );
    or g19366 ( n35191 , n34074 , n28324 );
    or g19367 ( n25851 , n27291 , n27715 );
    and g19368 ( n176 , n3722 , n22403 );
    or g19369 ( n20123 , n3222 , n33138 );
    xnor g19370 ( n7292 , n27326 , n31359 );
    or g19371 ( n1023 , n11525 , n29585 );
    and g19372 ( n21588 , n17192 , n27799 );
    and g19373 ( n24427 , n31668 , n35705 );
    xnor g19374 ( n20564 , n32841 , n27226 );
    not g19375 ( n20811 , n16292 );
    nor g19376 ( n26052 , n16879 , n30883 );
    xnor g19377 ( n3282 , n30805 , n10363 );
    or g19378 ( n20979 , n20178 , n21953 );
    or g19379 ( n15916 , n17081 , n20797 );
    not g19380 ( n32274 , n16938 );
    xnor g19381 ( n31571 , n26969 , n24586 );
    or g19382 ( n26570 , n27884 , n578 );
    or g19383 ( n9765 , n3876 , n25306 );
    nor g19384 ( n13420 , n16922 , n21893 );
    or g19385 ( n6357 , n18427 , n15538 );
    not g19386 ( n16651 , n32857 );
    and g19387 ( n10622 , n21365 , n11632 );
    and g19388 ( n25835 , n29553 , n34500 );
    or g19389 ( n7406 , n3732 , n16464 );
    and g19390 ( n18958 , n21515 , n9841 );
    and g19391 ( n15274 , n1073 , n27 );
    or g19392 ( n23003 , n14179 , n28323 );
    xnor g19393 ( n6211 , n3311 , n35005 );
    and g19394 ( n5345 , n25578 , n3476 );
    or g19395 ( n14053 , n27193 , n27963 );
    or g19396 ( n5430 , n17040 , n30654 );
    or g19397 ( n6523 , n35397 , n34273 );
    or g19398 ( n27398 , n20503 , n32959 );
    and g19399 ( n10663 , n15615 , n6943 );
    not g19400 ( n16115 , n7730 );
    or g19401 ( n22971 , n32541 , n4175 );
    or g19402 ( n3280 , n9008 , n3759 );
    not g19403 ( n4847 , n8157 );
    nor g19404 ( n21555 , n21212 , n25247 );
    or g19405 ( n2988 , n30527 , n28248 );
    xnor g19406 ( n13029 , n90 , n10718 );
    and g19407 ( n17805 , n6826 , n8530 );
    or g19408 ( n22712 , n1140 , n5588 );
    and g19409 ( n29848 , n21947 , n29596 );
    xnor g19410 ( n26817 , n22313 , n10573 );
    and g19411 ( n29949 , n8301 , n10069 );
    and g19412 ( n21441 , n18792 , n15123 );
    or g19413 ( n21614 , n29620 , n3842 );
    xnor g19414 ( n14678 , n4771 , n830 );
    or g19415 ( n17930 , n31289 , n10324 );
    or g19416 ( n1937 , n32095 , n28356 );
    or g19417 ( n28625 , n29485 , n24160 );
    xnor g19418 ( n10945 , n13732 , n3205 );
    not g19419 ( n9102 , n17982 );
    not g19420 ( n9137 , n444 );
    and g19421 ( n17353 , n10566 , n14577 );
    or g19422 ( n10014 , n10352 , n18488 );
    or g19423 ( n15061 , n16922 , n5076 );
    xnor g19424 ( n17171 , n21026 , n4962 );
    xnor g19425 ( n34544 , n31746 , n10894 );
    or g19426 ( n25936 , n3735 , n21691 );
    xnor g19427 ( n30714 , n34976 , n15073 );
    or g19428 ( n19320 , n380 , n21977 );
    or g19429 ( n34772 , n22483 , n24653 );
    and g19430 ( n7063 , n26576 , n24469 );
    or g19431 ( n23686 , n11055 , n10336 );
    and g19432 ( n21328 , n22058 , n17340 );
    or g19433 ( n22161 , n7366 , n20521 );
    xnor g19434 ( n31737 , n11271 , n3319 );
    or g19435 ( n17579 , n20328 , n19058 );
    or g19436 ( n34182 , n31107 , n5252 );
    xnor g19437 ( n13695 , n698 , n16985 );
    or g19438 ( n3080 , n31272 , n11223 );
    xnor g19439 ( n32995 , n15658 , n24394 );
    or g19440 ( n15233 , n210 , n32562 );
    not g19441 ( n20553 , n4822 );
    xnor g19442 ( n24225 , n14831 , n8471 );
    or g19443 ( n11440 , n11714 , n3634 );
    or g19444 ( n6070 , n30742 , n1046 );
    not g19445 ( n14425 , n26072 );
    or g19446 ( n27543 , n16881 , n3348 );
    nor g19447 ( n4116 , n4878 , n22301 );
    and g19448 ( n16532 , n25807 , n16511 );
    or g19449 ( n23457 , n35247 , n29643 );
    xnor g19450 ( n2719 , n20952 , n9789 );
    xnor g19451 ( n28145 , n34331 , n35927 );
    not g19452 ( n35859 , n26027 );
    buf g19453 ( n17962 , n21785 );
    not g19454 ( n26769 , n33401 );
    or g19455 ( n24359 , n17319 , n32505 );
    and g19456 ( n27866 , n12265 , n19080 );
    and g19457 ( n15841 , n25349 , n30274 );
    xnor g19458 ( n15844 , n6703 , n31559 );
    xnor g19459 ( n11529 , n24816 , n15464 );
    nor g19460 ( n25619 , n18282 , n9528 );
    xnor g19461 ( n5706 , n15463 , n18379 );
    and g19462 ( n4470 , n13412 , n33425 );
    and g19463 ( n7310 , n32551 , n25155 );
    or g19464 ( n25248 , n19589 , n5252 );
    or g19465 ( n22271 , n35319 , n11477 );
    or g19466 ( n22487 , n19010 , n12596 );
    and g19467 ( n10721 , n17778 , n16047 );
    or g19468 ( n9894 , n7994 , n26357 );
    or g19469 ( n33616 , n33902 , n11977 );
    nor g19470 ( n9699 , n4878 , n5064 );
    xnor g19471 ( n9509 , n5555 , n3746 );
    nor g19472 ( n34089 , n30061 , n35826 );
    or g19473 ( n1886 , n20492 , n7647 );
    or g19474 ( n20429 , n22400 , n8405 );
    or g19475 ( n32848 , n32493 , n34971 );
    nor g19476 ( n23537 , n18413 , n18654 );
    xnor g19477 ( n15415 , n17096 , n14119 );
    and g19478 ( n19603 , n17488 , n33679 );
    and g19479 ( n26290 , n10790 , n34169 );
    or g19480 ( n5665 , n28227 , n32572 );
    or g19481 ( n22651 , n5335 , n9936 );
    and g19482 ( n17402 , n27435 , n4317 );
    nor g19483 ( n26563 , n23604 , n23846 );
    nor g19484 ( n32438 , n30742 , n25888 );
    nor g19485 ( n9855 , n24210 , n19044 );
    or g19486 ( n12937 , n24235 , n20576 );
    xnor g19487 ( n26498 , n7158 , n25959 );
    and g19488 ( n28678 , n21734 , n10468 );
    or g19489 ( n8218 , n25452 , n11851 );
    and g19490 ( n23761 , n13321 , n19826 );
    or g19491 ( n2382 , n3900 , n14759 );
    xnor g19492 ( n12000 , n17677 , n32715 );
    and g19493 ( n16037 , n22510 , n29973 );
    nor g19494 ( n1265 , n90 , n10718 );
    or g19495 ( n6208 , n7250 , n6683 );
    xnor g19496 ( n4667 , n8717 , n31621 );
    xnor g19497 ( n19195 , n35354 , n4878 );
    or g19498 ( n35333 , n17570 , n35422 );
    or g19499 ( n4946 , n24921 , n33018 );
    xnor g19500 ( n14846 , n3664 , n36005 );
    or g19501 ( n35871 , n17382 , n28675 );
    not g19502 ( n20469 , n31799 );
    and g19503 ( n10563 , n22987 , n20052 );
    or g19504 ( n16912 , n28420 , n21176 );
    nor g19505 ( n2751 , n3946 , n21630 );
    or g19506 ( n8206 , n23604 , n29713 );
    and g19507 ( n22975 , n869 , n30497 );
    or g19508 ( n31028 , n11348 , n14429 );
    not g19509 ( n4800 , n30755 );
    or g19510 ( n4215 , n28166 , n14841 );
    or g19511 ( n32946 , n32964 , n24356 );
    or g19512 ( n13574 , n33197 , n7293 );
    or g19513 ( n5400 , n30938 , n21056 );
    or g19514 ( n35751 , n21371 , n17337 );
    not g19515 ( n33155 , n3480 );
    or g19516 ( n17167 , n8058 , n35332 );
    or g19517 ( n5300 , n34758 , n34452 );
    not g19518 ( n30607 , n33262 );
    xnor g19519 ( n11425 , n20666 , n27592 );
    or g19520 ( n31066 , n17740 , n4231 );
    and g19521 ( n14687 , n5430 , n3902 );
    xnor g19522 ( n12307 , n8049 , n31749 );
    xnor g19523 ( n29892 , n24934 , n4962 );
    and g19524 ( n4590 , n3012 , n12397 );
    and g19525 ( n33114 , n34946 , n7146 );
    not g19526 ( n334 , n14063 );
    or g19527 ( n18741 , n35573 , n7151 );
    not g19528 ( n6157 , n8101 );
    not g19529 ( n34912 , n6257 );
    or g19530 ( n28194 , n12446 , n27963 );
    and g19531 ( n4945 , n13685 , n22980 );
    or g19532 ( n22673 , n31799 , n3802 );
    xnor g19533 ( n3087 , n2367 , n1840 );
    or g19534 ( n1923 , n16595 , n22322 );
    and g19535 ( n2222 , n32166 , n32524 );
    xnor g19536 ( n6911 , n28593 , n4962 );
    or g19537 ( n10695 , n20170 , n13130 );
    xnor g19538 ( n34953 , n397 , n24610 );
    not g19539 ( n29464 , n32734 );
    nor g19540 ( n27607 , n3205 , n8005 );
    and g19541 ( n12966 , n17093 , n31156 );
    xnor g19542 ( n23877 , n5378 , n22717 );
    nor g19543 ( n26316 , n25839 , n30871 );
    and g19544 ( n15163 , n18315 , n8391 );
    or g19545 ( n30349 , n29713 , n33676 );
    not g19546 ( n23667 , n6505 );
    and g19547 ( n32520 , n2362 , n12868 );
    or g19548 ( n19620 , n34829 , n34923 );
    or g19549 ( n34653 , n9893 , n28909 );
    not g19550 ( n17892 , n24054 );
    xnor g19551 ( n24109 , n14288 , n24317 );
    or g19552 ( n32683 , n3946 , n18015 );
    nor g19553 ( n29923 , n26245 , n29203 );
    or g19554 ( n19788 , n25157 , n27963 );
    or g19555 ( n33579 , n8400 , n35402 );
    not g19556 ( n27890 , n4210 );
    or g19557 ( n1426 , n9658 , n10168 );
    nor g19558 ( n8934 , n643 , n24208 );
    nor g19559 ( n28148 , n35479 , n33034 );
    and g19560 ( n25606 , n32941 , n24429 );
    nor g19561 ( n63 , n17767 , n7375 );
    nor g19562 ( n29007 , n23081 , n34542 );
    or g19563 ( n20767 , n28317 , n28438 );
    or g19564 ( n19231 , n34533 , n12428 );
    or g19565 ( n26228 , n19346 , n16660 );
    buf g19566 ( n25567 , n93 );
    or g19567 ( n5698 , n27206 , n15351 );
    not g19568 ( n22097 , n33435 );
    xnor g19569 ( n25016 , n10134 , n21212 );
    or g19570 ( n13706 , n1998 , n5779 );
    and g19571 ( n33765 , n25532 , n7643 );
    nor g19572 ( n1014 , n14856 , n27728 );
    and g19573 ( n17698 , n35725 , n25145 );
    not g19574 ( n12163 , n18555 );
    or g19575 ( n6700 , n26175 , n24025 );
    xnor g19576 ( n1173 , n8552 , n16922 );
    or g19577 ( n18251 , n15884 , n23748 );
    and g19578 ( n25441 , n15379 , n20430 );
    xnor g19579 ( n9347 , n23132 , n29015 );
    or g19580 ( n34940 , n29713 , n9565 );
    and g19581 ( n30985 , n12530 , n31846 );
    and g19582 ( n12317 , n28644 , n25975 );
    or g19583 ( n3118 , n27638 , n10872 );
    xnor g19584 ( n21357 , n14138 , n31215 );
    or g19585 ( n16778 , n4056 , n16602 );
    or g19586 ( n8574 , n13657 , n25940 );
    xnor g19587 ( n35777 , n28175 , n7845 );
    and g19588 ( n24985 , n7870 , n25632 );
    or g19589 ( n5442 , n22846 , n1511 );
    or g19590 ( n30926 , n27787 , n8680 );
    xnor g19591 ( n26677 , n1222 , n17568 );
    xnor g19592 ( n27716 , n26083 , n14946 );
    and g19593 ( n24760 , n28967 , n7006 );
    or g19594 ( n23372 , n32857 , n4827 );
    xnor g19595 ( n4745 , n2965 , n11101 );
    or g19596 ( n35729 , n25558 , n26365 );
    or g19597 ( n19672 , n18072 , n19403 );
    not g19598 ( n1419 , n16223 );
    or g19599 ( n18882 , n9641 , n21144 );
    or g19600 ( n17092 , n13522 , n5561 );
    xnor g19601 ( n32642 , n10454 , n9111 );
    or g19602 ( n2604 , n6814 , n30826 );
    xnor g19603 ( n2102 , n36019 , n16110 );
    or g19604 ( n27581 , n8432 , n35249 );
    or g19605 ( n2935 , n12554 , n9731 );
    nor g19606 ( n20178 , n3443 , n18115 );
    or g19607 ( n2327 , n11931 , n3979 );
    or g19608 ( n4933 , n29495 , n29258 );
    or g19609 ( n16918 , n12267 , n21653 );
    or g19610 ( n4767 , n28545 , n8392 );
    xnor g19611 ( n932 , n6072 , n33210 );
    or g19612 ( n10590 , n4288 , n26208 );
    and g19613 ( n3882 , n14668 , n6630 );
    xnor g19614 ( n19168 , n28196 , n18678 );
    xnor g19615 ( n28899 , n25282 , n1950 );
    not g19616 ( n35895 , n29713 );
    or g19617 ( n27210 , n24371 , n4510 );
    or g19618 ( n22450 , n449 , n9410 );
    xnor g19619 ( n10211 , n3792 , n5375 );
    nor g19620 ( n4097 , n31272 , n11955 );
    and g19621 ( n19155 , n29337 , n15968 );
    and g19622 ( n35869 , n165 , n22355 );
    xnor g19623 ( n22168 , n6970 , n31711 );
    or g19624 ( n17459 , n20517 , n13900 );
    not g19625 ( n25638 , n35927 );
    nor g19626 ( n17544 , n7274 , n14221 );
    xnor g19627 ( n23875 , n2335 , n3222 );
    xnor g19628 ( n20514 , n29589 , n32584 );
    and g19629 ( n25247 , n32608 , n9590 );
    or g19630 ( n20792 , n2024 , n7647 );
    or g19631 ( n10470 , n9172 , n28601 );
    and g19632 ( n22386 , n12804 , n22506 );
    or g19633 ( n18002 , n14503 , n28449 );
    or g19634 ( n2588 , n5435 , n28262 );
    or g19635 ( n28469 , n32095 , n29929 );
    or g19636 ( n6733 , n23186 , n12824 );
    xnor g19637 ( n3889 , n329 , n11455 );
    xnor g19638 ( n1570 , n14680 , n11046 );
    or g19639 ( n12002 , n21447 , n34600 );
    or g19640 ( n23832 , n1525 , n15144 );
    and g19641 ( n4716 , n27414 , n31769 );
    or g19642 ( n13692 , n15787 , n19105 );
    or g19643 ( n25797 , n22864 , n35630 );
    nor g19644 ( n4566 , n34543 , n8404 );
    nor g19645 ( n27871 , n23604 , n14907 );
    and g19646 ( n18498 , n14758 , n8787 );
    and g19647 ( n17901 , n12737 , n19699 );
    xnor g19648 ( n5123 , n15759 , n8322 );
    or g19649 ( n6875 , n3752 , n26813 );
    nor g19650 ( n29439 , n35833 , n14545 );
    xnor g19651 ( n15116 , n35669 , n28023 );
    and g19652 ( n19690 , n17205 , n25388 );
    xnor g19653 ( n18234 , n4670 , n29839 );
    or g19654 ( n19164 , n8542 , n21042 );
    or g19655 ( n28359 , n6269 , n20579 );
    xnor g19656 ( n16672 , n30967 , n25174 );
    xnor g19657 ( n10876 , n27850 , n6321 );
    or g19658 ( n7467 , n15914 , n3437 );
    nor g19659 ( n18599 , n4962 , n2455 );
    or g19660 ( n34697 , n25160 , n22685 );
    or g19661 ( n12689 , n22442 , n32808 );
    xnor g19662 ( n25708 , n12850 , n24382 );
    or g19663 ( n64 , n30785 , n17612 );
    and g19664 ( n26729 , n7185 , n2881 );
    xnor g19665 ( n10776 , n9245 , n16587 );
    or g19666 ( n30668 , n22291 , n28472 );
    and g19667 ( n15501 , n6223 , n35266 );
    xnor g19668 ( n16394 , n6822 , n15377 );
    or g19669 ( n12290 , n29884 , n5368 );
    or g19670 ( n21302 , n24371 , n6316 );
    or g19671 ( n8700 , n17159 , n25594 );
    xnor g19672 ( n20398 , n17395 , n24371 );
    or g19673 ( n4810 , n22747 , n16457 );
    or g19674 ( n15107 , n26606 , n5534 );
    xnor g19675 ( n26887 , n31897 , n18207 );
    xnor g19676 ( n2140 , n20910 , n14847 );
    or g19677 ( n14614 , n4878 , n3686 );
    and g19678 ( n18899 , n11273 , n24398 );
    or g19679 ( n20432 , n13160 , n8245 );
    nor g19680 ( n35056 , n28624 , n1864 );
    xnor g19681 ( n32973 , n17525 , n32095 );
    nor g19682 ( n26323 , n24371 , n5324 );
    and g19683 ( n12774 , n20600 , n13288 );
    nor g19684 ( n34722 , n4999 , n29934 );
    or g19685 ( n34366 , n29816 , n16331 );
    or g19686 ( n16239 , n3663 , n27396 );
    xnor g19687 ( n34845 , n33456 , n26109 );
    or g19688 ( n27928 , n34265 , n7212 );
    nor g19689 ( n6833 , n26504 , n2823 );
    or g19690 ( n23451 , n19930 , n26737 );
    or g19691 ( n36052 , n29500 , n10548 );
    or g19692 ( n22921 , n25495 , n22961 );
    xnor g19693 ( n5318 , n16857 , n33765 );
    or g19694 ( n15418 , n32 , n31606 );
    nor g19695 ( n26876 , n31799 , n33968 );
    or g19696 ( n6147 , n2822 , n33615 );
    xnor g19697 ( n4035 , n33705 , n405 );
    or g19698 ( n1085 , n16922 , n30736 );
    or g19699 ( n9390 , n23622 , n25492 );
    and g19700 ( n4740 , n20884 , n27889 );
    or g19701 ( n4576 , n29767 , n25036 );
    not g19702 ( n10526 , n8865 );
    or g19703 ( n15852 , n19171 , n15250 );
    and g19704 ( n23959 , n1298 , n25758 );
    xnor g19705 ( n34837 , n16250 , n8432 );
    or g19706 ( n1568 , n13142 , n28969 );
    or g19707 ( n33371 , n12574 , n9033 );
    and g19708 ( n8241 , n17463 , n14862 );
    and g19709 ( n19537 , n32687 , n26403 );
    and g19710 ( n11737 , n5100 , n34335 );
    and g19711 ( n25589 , n12186 , n29619 );
    or g19712 ( n26717 , n19551 , n32328 );
    xnor g19713 ( n35347 , n12238 , n32480 );
    nor g19714 ( n22943 , n5335 , n18778 );
    or g19715 ( n4229 , n31099 , n9601 );
    and g19716 ( n16083 , n14756 , n17089 );
    or g19717 ( n34489 , n20765 , n17069 );
    or g19718 ( n6346 , n24331 , n7417 );
    xnor g19719 ( n3645 , n17995 , n33513 );
    xnor g19720 ( n10789 , n6917 , n28859 );
    or g19721 ( n20826 , n1652 , n19421 );
    xnor g19722 ( n23244 , n30112 , n12432 );
    and g19723 ( n22750 , n18609 , n4571 );
    nor g19724 ( n13628 , n3284 , n18115 );
    and g19725 ( n11211 , n870 , n35803 );
    and g19726 ( n23741 , n15451 , n4410 );
    or g19727 ( n4573 , n20087 , n22003 );
    buf g19728 ( n17162 , n17313 );
    and g19729 ( n518 , n501 , n35674 );
    or g19730 ( n33179 , n7178 , n3239 );
    xnor g19731 ( n1399 , n33789 , n24466 );
    and g19732 ( n34191 , n22501 , n12644 );
    or g19733 ( n11898 , n1950 , n21045 );
    or g19734 ( n2591 , n9085 , n21582 );
    or g19735 ( n21327 , n1316 , n3115 );
    xnor g19736 ( n32042 , n12740 , n3414 );
    xnor g19737 ( n7296 , n33853 , n16922 );
    or g19738 ( n27213 , n15460 , n15310 );
    or g19739 ( n27324 , n26895 , n12827 );
    not g19740 ( n10736 , n24364 );
    not g19741 ( n24463 , n32898 );
    or g19742 ( n22103 , n17866 , n30419 );
    or g19743 ( n33823 , n18633 , n32697 );
    or g19744 ( n13919 , n3551 , n33923 );
    and g19745 ( n8107 , n4735 , n18828 );
    nor g19746 ( n751 , n11455 , n32485 );
    or g19747 ( n25506 , n3157 , n30204 );
    xnor g19748 ( n994 , n20525 , n29934 );
    or g19749 ( n6084 , n4748 , n31514 );
    nor g19750 ( n22359 , n22447 , n34183 );
    or g19751 ( n9157 , n4255 , n19952 );
    or g19752 ( n8599 , n23052 , n34912 );
    or g19753 ( n21408 , n17622 , n17337 );
    and g19754 ( n25548 , n15242 , n31063 );
    and g19755 ( n4546 , n10755 , n1882 );
    or g19756 ( n1347 , n24302 , n31606 );
    xnor g19757 ( n29934 , n17470 , n16620 );
    and g19758 ( n20805 , n28761 , n23856 );
    xnor g19759 ( n15057 , n3210 , n29839 );
    or g19760 ( n6103 , n32417 , n21862 );
    or g19761 ( n32902 , n16538 , n12332 );
    and g19762 ( n27225 , n25528 , n34129 );
    xnor g19763 ( n12594 , n22689 , n32584 );
    or g19764 ( n24962 , n17043 , n7434 );
    nor g19765 ( n14371 , n35019 , n12913 );
    not g19766 ( n27074 , n22705 );
    xnor g19767 ( n25908 , n18915 , n18379 );
    nor g19768 ( n13887 , n12848 , n21935 );
    or g19769 ( n11701 , n31693 , n3523 );
    and g19770 ( n6338 , n8592 , n31170 );
    and g19771 ( n19925 , n11293 , n24601 );
    and g19772 ( n11204 , n11876 , n13260 );
    or g19773 ( n13267 , n6365 , n6938 );
    or g19774 ( n22654 , n13660 , n10914 );
    or g19775 ( n10850 , n22291 , n26101 );
    not g19776 ( n14757 , n22200 );
    buf g19777 ( n10634 , n13015 );
    and g19778 ( n26730 , n17595 , n299 );
    or g19779 ( n17465 , n9810 , n18811 );
    xnor g19780 ( n30479 , n27815 , n27226 );
    or g19781 ( n6942 , n35831 , n5972 );
    and g19782 ( n9990 , n24882 , n20378 );
    xnor g19783 ( n15595 , n25968 , n15371 );
    not g19784 ( n12035 , n915 );
    not g19785 ( n33469 , n2310 );
    or g19786 ( n21110 , n11292 , n10905 );
    or g19787 ( n29986 , n13872 , n128 );
    or g19788 ( n23505 , n30531 , n25866 );
    and g19789 ( n25887 , n7659 , n8786 );
    not g19790 ( n24753 , n7588 );
    not g19791 ( n5675 , n16389 );
    and g19792 ( n24161 , n28745 , n17828 );
    or g19793 ( n34032 , n1313 , n14554 );
    xnor g19794 ( n30241 , n8505 , n30721 );
    or g19795 ( n16383 , n30677 , n12538 );
    and g19796 ( n31843 , n8850 , n24907 );
    or g19797 ( n25566 , n12840 , n16543 );
    nor g19798 ( n12923 , n3078 , n9241 );
    not g19799 ( n268 , n1482 );
    xnor g19800 ( n16552 , n11872 , n11455 );
    or g19801 ( n35380 , n13512 , n20840 );
    or g19802 ( n14892 , n24908 , n3805 );
    xnor g19803 ( n13189 , n29984 , n11046 );
    xnor g19804 ( n27984 , n34953 , n27324 );
    or g19805 ( n35761 , n23812 , n6288 );
    nor g19806 ( n21462 , n19858 , n4774 );
    or g19807 ( n19585 , n28020 , n20427 );
    nor g19808 ( n35276 , n30578 , n17235 );
    xnor g19809 ( n9649 , n23343 , n8653 );
    and g19810 ( n6229 , n25450 , n13942 );
    and g19811 ( n18066 , n23232 , n17676 );
    not g19812 ( n4283 , n30742 );
    or g19813 ( n6792 , n11046 , n2076 );
    xnor g19814 ( n3312 , n2726 , n16620 );
    or g19815 ( n35179 , n2395 , n11295 );
    or g19816 ( n35452 , n19549 , n32959 );
    or g19817 ( n9311 , n6351 , n25941 );
    or g19818 ( n7508 , n15886 , n22256 );
    xnor g19819 ( n22363 , n31267 , n25164 );
    or g19820 ( n7465 , n25602 , n8776 );
    or g19821 ( n32602 , n2636 , n32329 );
    and g19822 ( n16579 , n11387 , n2643 );
    and g19823 ( n9626 , n17234 , n12644 );
    or g19824 ( n25937 , n9326 , n3383 );
    and g19825 ( n24315 , n2480 , n13551 );
    nor g19826 ( n7366 , n32715 , n5648 );
    not g19827 ( n33272 , n8977 );
    or g19828 ( n16203 , n29839 , n33256 );
    and g19829 ( n20961 , n18741 , n29893 );
    xnor g19830 ( n22503 , n35649 , n35927 );
    xnor g19831 ( n19578 , n15235 , n25602 );
    or g19832 ( n31158 , n11999 , n26192 );
    or g19833 ( n30765 , n18208 , n13217 );
    not g19834 ( n16338 , n23434 );
    or g19835 ( n15012 , n15738 , n30617 );
    nor g19836 ( n20291 , n32642 , n16849 );
    and g19837 ( n13648 , n24395 , n16053 );
    and g19838 ( n23276 , n31432 , n9461 );
    xnor g19839 ( n13427 , n7594 , n10557 );
    and g19840 ( n2232 , n21727 , n12079 );
    and g19841 ( n34737 , n5950 , n27517 );
    or g19842 ( n13297 , n17188 , n32425 );
    or g19843 ( n17323 , n4213 , n35143 );
    or g19844 ( n27165 , n20755 , n9097 );
    or g19845 ( n35302 , n7286 , n8090 );
    and g19846 ( n11892 , n6724 , n16629 );
    and g19847 ( n11501 , n8510 , n32724 );
    or g19848 ( n35774 , n32825 , n30204 );
    or g19849 ( n3605 , n32120 , n31710 );
    and g19850 ( n22993 , n13236 , n27293 );
    and g19851 ( n3489 , n8011 , n7193 );
    or g19852 ( n7148 , n22291 , n12803 );
    xnor g19853 ( n20677 , n25383 , n18364 );
    xnor g19854 ( n29808 , n27327 , n29552 );
    or g19855 ( n10596 , n4865 , n2739 );
    or g19856 ( n14781 , n35985 , n16457 );
    nor g19857 ( n24357 , n29752 , n16497 );
    or g19858 ( n11876 , n20944 , n34777 );
    or g19859 ( n24062 , n12850 , n26336 );
    or g19860 ( n29566 , n4960 , n20084 );
    or g19861 ( n23344 , n2395 , n32959 );
    and g19862 ( n8784 , n7533 , n4808 );
    xnor g19863 ( n14704 , n14220 , n19095 );
    or g19864 ( n28381 , n17299 , n19666 );
    and g19865 ( n16388 , n16066 , n25496 );
    xor g19866 ( n35760 , n14533 , n19551 );
    xnor g19867 ( n24633 , n6830 , n26781 );
    or g19868 ( n19109 , n5555 , n3746 );
    xnor g19869 ( n9493 , n34708 , n11046 );
    and g19870 ( n27518 , n9531 , n20145 );
    or g19871 ( n7633 , n25838 , n29411 );
    or g19872 ( n29189 , n10894 , n20912 );
    and g19873 ( n24822 , n27063 , n22046 );
    or g19874 ( n5471 , n32715 , n14148 );
    and g19875 ( n27212 , n21250 , n16452 );
    or g19876 ( n18892 , n30791 , n27719 );
    xnor g19877 ( n5920 , n34842 , n11455 );
    or g19878 ( n2976 , n34544 , n9529 );
    or g19879 ( n23166 , n19695 , n34702 );
    or g19880 ( n8861 , n3052 , n18274 );
    and g19881 ( n27031 , n1851 , n8226 );
    buf g19882 ( n27801 , n25761 );
    or g19883 ( n32233 , n18846 , n27704 );
    and g19884 ( n10380 , n15472 , n135 );
    xnor g19885 ( n23250 , n19457 , n31559 );
    xnor g19886 ( n8425 , n27611 , n31559 );
    or g19887 ( n21772 , n9997 , n19490 );
    not g19888 ( n20647 , n22544 );
    and g19889 ( n30206 , n24966 , n19582 );
    or g19890 ( n15988 , n4682 , n21956 );
    xnor g19891 ( n16155 , n22889 , n30341 );
    or g19892 ( n34619 , n11046 , n142 );
    or g19893 ( n23056 , n3753 , n1856 );
    and g19894 ( n27950 , n1814 , n5140 );
    xnor g19895 ( n12160 , n17659 , n35718 );
    or g19896 ( n9557 , n16135 , n19470 );
    or g19897 ( n14951 , n27226 , n15820 );
    xnor g19898 ( n20166 , n31422 , n18046 );
    xnor g19899 ( n4690 , n14043 , n25602 );
    xnor g19900 ( n27538 , n26759 , n18379 );
    xnor g19901 ( n36041 , n20913 , n29839 );
    and g19902 ( n5119 , n26402 , n6173 );
    xnor g19903 ( n15166 , n26183 , n4288 );
    or g19904 ( n5340 , n17177 , n2327 );
    or g19905 ( n6891 , n7742 , n32697 );
    and g19906 ( n978 , n31078 , n35819 );
    xnor g19907 ( n15945 , n24867 , n9793 );
    xnor g19908 ( n25688 , n24717 , n6947 );
    xnor g19909 ( n6193 , n32684 , n32427 );
    xnor g19910 ( n18742 , n35262 , n10894 );
    not g19911 ( n11646 , n34318 );
    or g19912 ( n21710 , n292 , n25241 );
    xnor g19913 ( n17474 , n12532 , n4962 );
    or g19914 ( n33135 , n18626 , n29118 );
    or g19915 ( n15862 , n13496 , n4952 );
    or g19916 ( n28930 , n10789 , n5972 );
    xnor g19917 ( n26266 , n33324 , n26209 );
    and g19918 ( n16152 , n28339 , n24084 );
    or g19919 ( n28522 , n20588 , n12495 );
    and g19920 ( n28539 , n31058 , n18555 );
    xnor g19921 ( n4061 , n17007 , n33622 );
    or g19922 ( n24323 , n20568 , n613 );
    and g19923 ( n22105 , n18138 , n29729 );
    and g19924 ( n16972 , n8017 , n34536 );
    xnor g19925 ( n7893 , n21881 , n34811 );
    xnor g19926 ( n18748 , n14655 , n3222 );
    or g19927 ( n33077 , n11881 , n27501 );
    or g19928 ( n34399 , n4457 , n10762 );
    and g19929 ( n10112 , n35734 , n17477 );
    or g19930 ( n24358 , n16922 , n19374 );
    buf g19931 ( n14841 , n34458 );
    xnor g19932 ( n17546 , n2717 , n14411 );
    xnor g19933 ( n18100 , n14537 , n16620 );
    xnor g19934 ( n17031 , n35328 , n9658 );
    and g19935 ( n26208 , n7241 , n84 );
    or g19936 ( n27898 , n11435 , n1402 );
    and g19937 ( n14808 , n2272 , n20449 );
    xnor g19938 ( n20223 , n150 , n7851 );
    or g19939 ( n29403 , n33374 , n18280 );
    or g19940 ( n17039 , n825 , n12758 );
    not g19941 ( n18137 , n22705 );
    xnor g19942 ( n32146 , n3793 , n8050 );
    or g19943 ( n22840 , n31339 , n27408 );
    and g19944 ( n30488 , n12274 , n810 );
    not g19945 ( n11126 , n2339 );
    or g19946 ( n35651 , n16708 , n3415 );
    and g19947 ( n7479 , n21656 , n16198 );
    and g19948 ( n16569 , n32432 , n11948 );
    or g19949 ( n5896 , n35377 , n3344 );
    and g19950 ( n12569 , n9369 , n10298 );
    and g19951 ( n16820 , n26640 , n28825 );
    or g19952 ( n29768 , n13346 , n22783 );
    or g19953 ( n32713 , n21888 , n32507 );
    or g19954 ( n19758 , n20293 , n33338 );
    xnor g19955 ( n12756 , n24104 , n27291 );
    xnor g19956 ( n8150 , n33376 , n11046 );
    and g19957 ( n35557 , n7181 , n13137 );
    or g19958 ( n29982 , n25174 , n15875 );
    xnor g19959 ( n34740 , n23706 , n3426 );
    or g19960 ( n34148 , n2453 , n28248 );
    nor g19961 ( n1321 , n29713 , n8614 );
    or g19962 ( n23931 , n8027 , n862 );
    or g19963 ( n21855 , n25602 , n32452 );
    or g19964 ( n21920 , n29765 , n15145 );
    and g19965 ( n20228 , n1243 , n10186 );
    or g19966 ( n24616 , n12320 , n30431 );
    or g19967 ( n27829 , n32645 , n28248 );
    or g19968 ( n13707 , n9994 , n27343 );
    or g19969 ( n32301 , n14039 , n31554 );
    or g19970 ( n6110 , n15699 , n10662 );
    or g19971 ( n2571 , n19449 , n22858 );
    or g19972 ( n22156 , n19275 , n5833 );
    or g19973 ( n28321 , n25148 , n16797 );
    not g19974 ( n20450 , n7795 );
    and g19975 ( n5096 , n15269 , n25848 );
    or g19976 ( n10215 , n8103 , n22206 );
    xnor g19977 ( n22166 , n35724 , n23604 );
    and g19978 ( n31999 , n26558 , n25359 );
    nor g19979 ( n16952 , n4878 , n22236 );
    xnor g19980 ( n22065 , n32287 , n31613 );
    or g19981 ( n3034 , n23699 , n29953 );
    or g19982 ( n5439 , n30661 , n20427 );
    or g19983 ( n3555 , n21129 , n1176 );
    not g19984 ( n14182 , n33442 );
    or g19985 ( n33992 , n27089 , n5868 );
    or g19986 ( n17948 , n15886 , n22127 );
    and g19987 ( n25414 , n2499 , n25996 );
    or g19988 ( n23784 , n1671 , n20002 );
    xnor g19989 ( n4242 , n27319 , n5507 );
    and g19990 ( n34481 , n27112 , n5572 );
    or g19991 ( n2747 , n18531 , n29302 );
    xnor g19992 ( n16990 , n19488 , n6669 );
    or g19993 ( n234 , n18278 , n5064 );
    or g19994 ( n28044 , n12451 , n4436 );
    or g19995 ( n11504 , n12590 , n8587 );
    or g19996 ( n24997 , n7670 , n25831 );
    xnor g19997 ( n14065 , n26967 , n30156 );
    not g19998 ( n10177 , n32857 );
    or g19999 ( n29894 , n32879 , n19989 );
    or g20000 ( n13543 , n30566 , n26195 );
    xnor g20001 ( n2589 , n3929 , n23391 );
    or g20002 ( n3585 , n7540 , n32778 );
    xnor g20003 ( n11253 , n15657 , n10894 );
    or g20004 ( n24058 , n27594 , n33618 );
    xnor g20005 ( n22539 , n22626 , n3222 );
    and g20006 ( n4359 , n10937 , n16187 );
    and g20007 ( n18946 , n36073 , n17269 );
    xnor g20008 ( n21428 , n4345 , n26342 );
    or g20009 ( n4836 , n18109 , n2122 );
    buf g20010 ( n3634 , n16863 );
    buf g20011 ( n30292 , n3610 );
    or g20012 ( n5822 , n34346 , n24672 );
    nor g20013 ( n25417 , n31799 , n35383 );
    or g20014 ( n7731 , n15526 , n13792 );
    xnor g20015 ( n5297 , n12920 , n4342 );
    and g20016 ( n6996 , n14314 , n11751 );
    xnor g20017 ( n31693 , n21231 , n5679 );
    and g20018 ( n23605 , n2000 , n22635 );
    or g20019 ( n30078 , n9793 , n35914 );
    or g20020 ( n10964 , n11455 , n24445 );
    and g20021 ( n17018 , n8 , n24308 );
    or g20022 ( n23286 , n6714 , n9832 );
    and g20023 ( n3761 , n18049 , n35812 );
    xnor g20024 ( n26268 , n1305 , n14979 );
    or g20025 ( n9475 , n24040 , n14706 );
    and g20026 ( n23735 , n17039 , n33234 );
    xnor g20027 ( n2952 , n35865 , n3205 );
    or g20028 ( n15407 , n7540 , n22070 );
    or g20029 ( n34633 , n28851 , n18829 );
    or g20030 ( n13474 , n12330 , n9361 );
    xnor g20031 ( n8110 , n8260 , n26595 );
    or g20032 ( n17734 , n32685 , n17829 );
    or g20033 ( n5750 , n26074 , n437 );
    or g20034 ( n27920 , n11879 , n29987 );
    nor g20035 ( n13504 , n19551 , n1712 );
    or g20036 ( n30118 , n512 , n17829 );
    not g20037 ( n1905 , n4758 );
    and g20038 ( n2733 , n23031 , n16369 );
    or g20039 ( n31803 , n23908 , n6961 );
    xnor g20040 ( n31534 , n28971 , n21010 );
    and g20041 ( n18235 , n25650 , n2675 );
    xnor g20042 ( n16885 , n9266 , n15812 );
    and g20043 ( n4515 , n17341 , n31925 );
    and g20044 ( n26569 , n30627 , n22042 );
    nor g20045 ( n26606 , n5287 , n35465 );
    xnor g20046 ( n9031 , n203 , n24529 );
    or g20047 ( n12333 , n7291 , n14841 );
    not g20048 ( n29607 , n29628 );
    or g20049 ( n33966 , n14494 , n837 );
    or g20050 ( n26645 , n22994 , n26105 );
    or g20051 ( n2381 , n11046 , n19851 );
    nor g20052 ( n19214 , n18379 , n3701 );
    not g20053 ( n32243 , n8171 );
    and g20054 ( n13075 , n21198 , n27153 );
    and g20055 ( n4771 , n20742 , n10830 );
    or g20056 ( n32870 , n13889 , n23187 );
    not g20057 ( n28712 , n31126 );
    or g20058 ( n4225 , n12039 , n30296 );
    and g20059 ( n22353 , n18140 , n7794 );
    or g20060 ( n22481 , n27252 , n11295 );
    and g20061 ( n14984 , n35987 , n14433 );
    or g20062 ( n24399 , n6143 , n19403 );
    or g20063 ( n8193 , n22560 , n25019 );
    xnor g20064 ( n12915 , n17983 , n6582 );
    or g20065 ( n34788 , n25174 , n27534 );
    or g20066 ( n6608 , n19777 , n20546 );
    xnor g20067 ( n13239 , n17602 , n33468 );
    or g20068 ( n9756 , n21615 , n7221 );
    nor g20069 ( n25262 , n20647 , n8000 );
    or g20070 ( n16080 , n18099 , n12996 );
    and g20071 ( n31147 , n11908 , n622 );
    and g20072 ( n19151 , n4632 , n4993 );
    or g20073 ( n8053 , n26253 , n3437 );
    and g20074 ( n35057 , n10234 , n14367 );
    or g20075 ( n35153 , n27874 , n25657 );
    xnor g20076 ( n3315 , n29029 , n21676 );
    not g20077 ( n20822 , n31799 );
    or g20078 ( n22414 , n5242 , n30431 );
    or g20079 ( n15961 , n12247 , n35763 );
    and g20080 ( n26947 , n8341 , n26726 );
    xnor g20081 ( n25102 , n5350 , n640 );
    and g20082 ( n32853 , n5404 , n23017 );
    and g20083 ( n28034 , n34372 , n5334 );
    not g20084 ( n20959 , n15886 );
    xnor g20085 ( n28374 , n1712 , n19551 );
    and g20086 ( n33101 , n3612 , n30283 );
    xnor g20087 ( n20660 , n27297 , n272 );
    or g20088 ( n16998 , n34277 , n6487 );
    or g20089 ( n27882 , n22451 , n3595 );
    or g20090 ( n16727 , n22722 , n12557 );
    and g20091 ( n23981 , n32323 , n22778 );
    or g20092 ( n30959 , n18411 , n9317 );
    or g20093 ( n2919 , n2214 , n16326 );
    and g20094 ( n34370 , n25138 , n23476 );
    or g20095 ( n25800 , n4962 , n34159 );
    or g20096 ( n9548 , n30062 , n9930 );
    and g20097 ( n3708 , n10476 , n22805 );
    xnor g20098 ( n19011 , n11157 , n15886 );
    xnor g20099 ( n33958 , n3360 , n22907 );
    xnor g20100 ( n35831 , n17588 , n9575 );
    and g20101 ( n14021 , n2186 , n19498 );
    xnor g20102 ( n21293 , n7023 , n1021 );
    or g20103 ( n33308 , n19042 , n33310 );
    and g20104 ( n10408 , n33092 , n25986 );
    not g20105 ( n7697 , n19159 );
    or g20106 ( n24882 , n31824 , n29842 );
    or g20107 ( n5575 , n17128 , n9194 );
    or g20108 ( n8758 , n31715 , n3352 );
    xnor g20109 ( n34662 , n28678 , n32857 );
    and g20110 ( n20637 , n20207 , n31342 );
    nor g20111 ( n29853 , n2973 , n2653 );
    or g20112 ( n34200 , n8140 , n17409 );
    and g20113 ( n31194 , n27664 , n5000 );
    nor g20114 ( n27612 , n17355 , n33956 );
    or g20115 ( n25428 , n16230 , n30299 );
    or g20116 ( n24891 , n4962 , n25317 );
    xnor g20117 ( n9621 , n31926 , n7115 );
    or g20118 ( n25770 , n29713 , n34767 );
    xnor g20119 ( n11317 , n18981 , n21130 );
    or g20120 ( n25072 , n32095 , n29945 );
    and g20121 ( n6369 , n3263 , n30742 );
    xnor g20122 ( n21877 , n9693 , n20469 );
    or g20123 ( n30043 , n11702 , n23748 );
    nor g20124 ( n10497 , n10894 , n30117 );
    xnor g20125 ( n35034 , n14458 , n30140 );
    not g20126 ( n27649 , n8870 );
    or g20127 ( n9835 , n2081 , n8090 );
    or g20128 ( n13120 , n24790 , n18255 );
    or g20129 ( n2109 , n13278 , n29953 );
    or g20130 ( n19053 , n21596 , n36007 );
    or g20131 ( n19240 , n4981 , n13900 );
    or g20132 ( n1368 , n17325 , n8684 );
    nor g20133 ( n7874 , n35927 , n20095 );
    or g20134 ( n28741 , n32136 , n10960 );
    xnor g20135 ( n29968 , n5039 , n27294 );
    or g20136 ( n14816 , n35115 , n22458 );
    xnor g20137 ( n11414 , n25729 , n29713 );
    and g20138 ( n23532 , n6850 , n874 );
    xnor g20139 ( n8780 , n34568 , n6212 );
    or g20140 ( n21438 , n10145 , n18255 );
    or g20141 ( n28408 , n18381 , n20318 );
    xnor g20142 ( n15601 , n34030 , n830 );
    xnor g20143 ( n23793 , n32600 , n9702 );
    or g20144 ( n30484 , n4288 , n22610 );
    and g20145 ( n9373 , n9505 , n23860 );
    or g20146 ( n35114 , n8595 , n31773 );
    or g20147 ( n10626 , n34541 , n18477 );
    or g20148 ( n28771 , n14067 , n11771 );
    or g20149 ( n12709 , n16591 , n29565 );
    nor g20150 ( n15715 , n30742 , n28661 );
    or g20151 ( n19613 , n34400 , n8057 );
    or g20152 ( n16593 , n20513 , n6318 );
    not g20153 ( n21619 , n19458 );
    nor g20154 ( n14504 , n24873 , n35417 );
    and g20155 ( n4842 , n15935 , n6353 );
    xnor g20156 ( n31187 , n15332 , n32701 );
    xnor g20157 ( n25008 , n21663 , n8432 );
    xnor g20158 ( n4720 , n30290 , n10894 );
    not g20159 ( n6424 , n22200 );
    or g20160 ( n15837 , n9793 , n23708 );
    or g20161 ( n4641 , n304 , n9679 );
    nor g20162 ( n18119 , n9793 , n34918 );
    and g20163 ( n3774 , n7182 , n1895 );
    or g20164 ( n19704 , n8016 , n3156 );
    or g20165 ( n9828 , n19639 , n7864 );
    or g20166 ( n11231 , n26440 , n15585 );
    xnor g20167 ( n23121 , n15406 , n9482 );
    or g20168 ( n12304 , n31057 , n22719 );
    or g20169 ( n33894 , n9477 , n9428 );
    xnor g20170 ( n11502 , n21733 , n10982 );
    or g20171 ( n24405 , n3946 , n10620 );
    and g20172 ( n14688 , n32986 , n33797 );
    or g20173 ( n6985 , n7041 , n15303 );
    or g20174 ( n26227 , n24371 , n32614 );
    or g20175 ( n35595 , n15947 , n6607 );
    or g20176 ( n5759 , n21980 , n18623 );
    or g20177 ( n10667 , n4288 , n24820 );
    and g20178 ( n21108 , n12031 , n33802 );
    xnor g20179 ( n890 , n34618 , n24371 );
    xnor g20180 ( n17072 , n23177 , n31289 );
    or g20181 ( n10614 , n17565 , n1404 );
    nor g20182 ( n27474 , n35927 , n15590 );
    xnor g20183 ( n4353 , n33488 , n9301 );
    xnor g20184 ( n16485 , n17136 , n32303 );
    nor g20185 ( n28035 , n31799 , n18231 );
    nor g20186 ( n11821 , n30742 , n17095 );
    or g20187 ( n27413 , n5287 , n28206 );
    and g20188 ( n17429 , n3871 , n33130 );
    and g20189 ( n15714 , n16235 , n21898 );
    nor g20190 ( n8268 , n24610 , n34501 );
    xnor g20191 ( n34979 , n11368 , n22496 );
    and g20192 ( n10317 , n25743 , n34584 );
    not g20193 ( n11474 , n4878 );
    or g20194 ( n7280 , n13407 , n28866 );
    or g20195 ( n29751 , n8432 , n12458 );
    or g20196 ( n11109 , n10768 , n1176 );
    nor g20197 ( n2689 , n31822 , n32199 );
    xnor g20198 ( n11618 , n4753 , n31559 );
    not g20199 ( n6927 , n17363 );
    or g20200 ( n179 , n17525 , n20318 );
    xnor g20201 ( n17691 , n31546 , n19551 );
    nor g20202 ( n35188 , n30742 , n2470 );
    or g20203 ( n25297 , n16769 , n4203 );
    or g20204 ( n14028 , n8432 , n12545 );
    xor g20205 ( n27375 , n8547 , n33040 );
    or g20206 ( n13500 , n36084 , n1557 );
    and g20207 ( n31784 , n34368 , n33351 );
    or g20208 ( n33312 , n3023 , n30238 );
    or g20209 ( n36062 , n11888 , n32071 );
    xnor g20210 ( n25926 , n28174 , n9658 );
    or g20211 ( n27945 , n29444 , n3694 );
    xnor g20212 ( n4654 , n29490 , n25154 );
    or g20213 ( n21917 , n32857 , n34162 );
    not g20214 ( n17886 , n27226 );
    xnor g20215 ( n23666 , n31932 , n33364 );
    and g20216 ( n17357 , n16549 , n26036 );
    or g20217 ( n34442 , n26916 , n18477 );
    nor g20218 ( n8814 , n32857 , n30036 );
    nor g20219 ( n30949 , n24011 , n3710 );
    or g20220 ( n1526 , n3946 , n1515 );
    xnor g20221 ( n3070 , n18022 , n6394 );
    xor g20222 ( n34274 , n2926 , n18908 );
    or g20223 ( n28858 , n25141 , n21540 );
    xnor g20224 ( n26212 , n35368 , n16620 );
    or g20225 ( n31196 , n21352 , n6340 );
    or g20226 ( n7156 , n9218 , n29624 );
    xnor g20227 ( n10941 , n8834 , n32857 );
    buf g20228 ( n26112 , n3437 );
    or g20229 ( n5375 , n10058 , n5119 );
    or g20230 ( n28003 , n24177 , n9058 );
    or g20231 ( n30411 , n22734 , n31554 );
    or g20232 ( n19313 , n31797 , n29880 );
    and g20233 ( n12853 , n10744 , n16655 );
    or g20234 ( n28006 , n16922 , n34258 );
    and g20235 ( n27645 , n9845 , n21498 );
    or g20236 ( n19960 , n23684 , n25648 );
    nor g20237 ( n19362 , n8432 , n16937 );
    xnor g20238 ( n28908 , n16044 , n1755 );
    xnor g20239 ( n22702 , n24608 , n31287 );
    or g20240 ( n19525 , n5029 , n6821 );
    nor g20241 ( n6131 , n11190 , n12667 );
    xnor g20242 ( n27805 , n5577 , n16461 );
    and g20243 ( n14805 , n27775 , n10907 );
    or g20244 ( n35993 , n34979 , n17068 );
    or g20245 ( n33013 , n9078 , n27720 );
    or g20246 ( n5847 , n25882 , n4363 );
    xnor g20247 ( n25147 , n32219 , n14086 );
    or g20248 ( n14711 , n17016 , n9317 );
    nor g20249 ( n33639 , n7540 , n35598 );
    not g20250 ( n31926 , n15464 );
    or g20251 ( n21163 , n31424 , n29716 );
    or g20252 ( n20635 , n8437 , n15256 );
    and g20253 ( n28799 , n25287 , n10100 );
    or g20254 ( n12786 , n18999 , n30287 );
    xnor g20255 ( n3503 , n16874 , n29839 );
    nor g20256 ( n6847 , n22155 , n33157 );
    or g20257 ( n12079 , n25122 , n10960 );
    xnor g20258 ( n1427 , n3223 , n4960 );
    or g20259 ( n30844 , n31999 , n24653 );
    and g20260 ( n35727 , n16455 , n20891 );
    or g20261 ( n17359 , n27317 , n10961 );
    and g20262 ( n32911 , n24060 , n815 );
    or g20263 ( n21407 , n11743 , n29052 );
    or g20264 ( n24267 , n24068 , n3257 );
    nor g20265 ( n24068 , n4174 , n9921 );
    or g20266 ( n4207 , n473 , n32388 );
    or g20267 ( n8530 , n28098 , n11996 );
    or g20268 ( n4676 , n8432 , n28187 );
    or g20269 ( n9198 , n22050 , n19421 );
    nor g20270 ( n21303 , n19702 , n7448 );
    and g20271 ( n30328 , n35461 , n26547 );
    not g20272 ( n7198 , n25301 );
    or g20273 ( n33211 , n11911 , n677 );
    xnor g20274 ( n17641 , n23202 , n29530 );
    or g20275 ( n967 , n17746 , n29626 );
    and g20276 ( n20127 , n858 , n33613 );
    not g20277 ( n172 , n33085 );
    not g20278 ( n20172 , n28273 );
    xnor g20279 ( n21138 , n18562 , n16079 );
    xnor g20280 ( n20867 , n11530 , n29650 );
    xnor g20281 ( n9154 , n7999 , n15969 );
    or g20282 ( n22820 , n18341 , n8197 );
    not g20283 ( n29867 , n13822 );
    and g20284 ( n14575 , n2565 , n27374 );
    or g20285 ( n14834 , n97 , n35630 );
    or g20286 ( n23720 , n29278 , n19421 );
    xnor g20287 ( n7343 , n2954 , n17554 );
    and g20288 ( n34527 , n16267 , n977 );
    or g20289 ( n25449 , n12556 , n34552 );
    or g20290 ( n3254 , n7410 , n26930 );
    or g20291 ( n5514 , n6003 , n1414 );
    not g20292 ( n28603 , n15368 );
    xnor g20293 ( n4346 , n30515 , n30742 );
    not g20294 ( n27300 , n17568 );
    and g20295 ( n5090 , n17626 , n8072 );
    and g20296 ( n29693 , n10503 , n2401 );
    or g20297 ( n8738 , n14118 , n21151 );
    or g20298 ( n24547 , n10825 , n34199 );
    nor g20299 ( n15100 , n7477 , n4338 );
    xnor g20300 ( n29859 , n30670 , n5335 );
    or g20301 ( n28193 , n24109 , n31627 );
    and g20302 ( n7344 , n15851 , n17149 );
    or g20303 ( n17090 , n23063 , n13786 );
    or g20304 ( n6758 , n26359 , n27963 );
    or g20305 ( n29112 , n34447 , n32329 );
    xnor g20306 ( n1633 , n16505 , n25602 );
    xnor g20307 ( n14634 , n23064 , n4962 );
    and g20308 ( n21757 , n27998 , n19520 );
    or g20309 ( n26750 , n33073 , n17046 );
    and g20310 ( n1663 , n10750 , n27749 );
    or g20311 ( n14615 , n1590 , n28324 );
    not g20312 ( n18332 , n31289 );
    or g20313 ( n25371 , n15535 , n19614 );
    and g20314 ( n35579 , n18391 , n11003 );
    or g20315 ( n6770 , n16891 , n28255 );
    nor g20316 ( n6431 , n19551 , n10287 );
    and g20317 ( n27056 , n283 , n34439 );
    or g20318 ( n33827 , n33884 , n54 );
    or g20319 ( n7026 , n2172 , n19198 );
    xnor g20320 ( n24221 , n30311 , n22959 );
    and g20321 ( n35992 , n34616 , n23107 );
    xnor g20322 ( n24444 , n23800 , n20637 );
    or g20323 ( n1434 , n8432 , n32546 );
    and g20324 ( n3210 , n31872 , n30450 );
    or g20325 ( n29217 , n35927 , n4180 );
    not g20326 ( n17659 , n5738 );
    not g20327 ( n1554 , n3347 );
    and g20328 ( n384 , n2151 , n1210 );
    nor g20329 ( n1315 , n15940 , n2261 );
    and g20330 ( n13462 , n4909 , n35611 );
    or g20331 ( n21325 , n24573 , n14841 );
    or g20332 ( n30394 , n28564 , n20308 );
    xnor g20333 ( n7739 , n24450 , n19551 );
    xnor g20334 ( n19963 , n35641 , n2293 );
    and g20335 ( n30736 , n22743 , n8496 );
    or g20336 ( n18951 , n23115 , n34484 );
    xnor g20337 ( n9451 , n21927 , n35093 );
    and g20338 ( n22923 , n20695 , n22113 );
    or g20339 ( n6570 , n23604 , n25760 );
    or g20340 ( n30869 , n17086 , n32866 );
    not g20341 ( n16897 , n1950 );
    or g20342 ( n5192 , n1852 , n26737 );
    or g20343 ( n27419 , n21175 , n10960 );
    not g20344 ( n31153 , n1574 );
    or g20345 ( n29544 , n34314 , n6082 );
    or g20346 ( n5878 , n5541 , n26468 );
    and g20347 ( n18364 , n192 , n26080 );
    xnor g20348 ( n32082 , n8323 , n1145 );
    xor g20349 ( n24654 , n26535 , n2532 );
    or g20350 ( n34789 , n4009 , n30292 );
    and g20351 ( n33346 , n17669 , n10926 );
    and g20352 ( n2890 , n27278 , n33953 );
    xnor g20353 ( n33067 , n1068 , n22374 );
    and g20354 ( n16248 , n14022 , n7843 );
    and g20355 ( n9850 , n488 , n34916 );
    or g20356 ( n13977 , n17568 , n25918 );
    or g20357 ( n31592 , n9827 , n22858 );
    or g20358 ( n29669 , n32095 , n8244 );
    or g20359 ( n1464 , n26165 , n524 );
    or g20360 ( n26682 , n9389 , n35458 );
    nor g20361 ( n1802 , n16620 , n34462 );
    or g20362 ( n28511 , n22687 , n29341 );
    and g20363 ( n18615 , n893 , n23168 );
    or g20364 ( n20000 , n19927 , n32274 );
    or g20365 ( n29177 , n21731 , n27764 );
    or g20366 ( n31717 , n35004 , n21002 );
    xnor g20367 ( n17537 , n26053 , n17153 );
    or g20368 ( n17615 , n28571 , n17125 );
    not g20369 ( n27923 , n3515 );
    or g20370 ( n11099 , n26364 , n28953 );
    nor g20371 ( n30581 , n10894 , n35262 );
    nor g20372 ( n18245 , n4960 , n7273 );
    or g20373 ( n8946 , n17129 , n34135 );
    xnor g20374 ( n24703 , n7110 , n30742 );
    or g20375 ( n14228 , n32857 , n18102 );
    xnor g20376 ( n16865 , n25081 , n35228 );
    nor g20377 ( n19531 , n19551 , n20159 );
    or g20378 ( n6007 , n6976 , n27501 );
    and g20379 ( n18944 , n18685 , n21948 );
    or g20380 ( n31122 , n4740 , n18255 );
    and g20381 ( n25725 , n24072 , n11153 );
    and g20382 ( n20790 , n12839 , n23285 );
    or g20383 ( n29401 , n34978 , n19952 );
    or g20384 ( n893 , n27461 , n19433 );
    not g20385 ( n33025 , n20535 );
    xnor g20386 ( n28082 , n11975 , n16608 );
    xnor g20387 ( n32036 , n9120 , n2728 );
    not g20388 ( n14535 , n26459 );
    xnor g20389 ( n34751 , n27658 , n21358 );
    or g20390 ( n6776 , n7540 , n24048 );
    xnor g20391 ( n33657 , n34623 , n31215 );
    and g20392 ( n27995 , n15592 , n4005 );
    buf g20393 ( n19834 , n9554 );
    or g20394 ( n12397 , n17751 , n4423 );
    xnor g20395 ( n1767 , n21521 , n31799 );
    xnor g20396 ( n33743 , n9136 , n32857 );
    nor g20397 ( n13129 , n31065 , n29203 );
    not g20398 ( n20644 , n27471 );
    or g20399 ( n22497 , n19086 , n26190 );
    or g20400 ( n35094 , n23604 , n33911 );
    and g20401 ( n26237 , n26082 , n1084 );
    and g20402 ( n7242 , n31483 , n16195 );
    or g20403 ( n10458 , n27226 , n35557 );
    and g20404 ( n27337 , n29858 , n17920 );
    or g20405 ( n8433 , n1083 , n34472 );
    or g20406 ( n29252 , n6113 , n25372 );
    and g20407 ( n13956 , n12449 , n32615 );
    and g20408 ( n29557 , n16346 , n9375 );
    not g20409 ( n7478 , n27156 );
    not g20410 ( n17855 , n32620 );
    not g20411 ( n721 , n4962 );
    or g20412 ( n11915 , n21928 , n25036 );
    or g20413 ( n5762 , n8432 , n19333 );
    and g20414 ( n34816 , n25284 , n15389 );
    and g20415 ( n27254 , n14992 , n31315 );
    or g20416 ( n9027 , n33537 , n2119 );
    or g20417 ( n5063 , n23198 , n8153 );
    not g20418 ( n30711 , n16052 );
    or g20419 ( n11050 , n22782 , n15805 );
    or g20420 ( n18937 , n35511 , n3604 );
    or g20421 ( n12156 , n26524 , n16435 );
    and g20422 ( n3575 , n32188 , n7510 );
    or g20423 ( n3898 , n5067 , n21846 );
    or g20424 ( n9059 , n23265 , n7726 );
    xnor g20425 ( n15941 , n3951 , n3205 );
    nor g20426 ( n10668 , n14140 , n21105 );
    or g20427 ( n31655 , n24312 , n24124 );
    and g20428 ( n21518 , n29763 , n22653 );
    and g20429 ( n4423 , n10994 , n22430 );
    or g20430 ( n6520 , n658 , n2104 );
    and g20431 ( n5855 , n30990 , n1548 );
    and g20432 ( n19721 , n659 , n21435 );
    or g20433 ( n32623 , n24371 , n425 );
    and g20434 ( n13364 , n8744 , n24316 );
    or g20435 ( n17723 , n4288 , n26995 );
    xnor g20436 ( n20464 , n16415 , n4288 );
    and g20437 ( n17746 , n14469 , n24738 );
    nor g20438 ( n35208 , n31559 , n2325 );
    and g20439 ( n26689 , n11420 , n27640 );
    nor g20440 ( n30280 , n1680 , n35834 );
    and g20441 ( n9209 , n11583 , n1933 );
    or g20442 ( n24461 , n7540 , n6735 );
    or g20443 ( n10679 , n32095 , n692 );
    and g20444 ( n36058 , n12655 , n25032 );
    or g20445 ( n28319 , n32584 , n29276 );
    xnor g20446 ( n19029 , n26783 , n20284 );
    nor g20447 ( n4796 , n15886 , n23067 );
    or g20448 ( n31023 , n32095 , n2191 );
    xnor g20449 ( n2072 , n24206 , n35873 );
    nor g20450 ( n22542 , n34637 , n16649 );
    or g20451 ( n3333 , n31422 , n18046 );
    and g20452 ( n8907 , n18112 , n22330 );
    buf g20453 ( n23323 , n16863 );
    and g20454 ( n17422 , n27987 , n10086 );
    or g20455 ( n7860 , n19726 , n17078 );
    nor g20456 ( n11638 , n26266 , n24287 );
    or g20457 ( n5517 , n20279 , n24663 );
    nor g20458 ( n28410 , n1066 , n17944 );
    or g20459 ( n15396 , n23057 , n10625 );
    xnor g20460 ( n16422 , n13162 , n117 );
    and g20461 ( n33716 , n16482 , n18821 );
    or g20462 ( n35524 , n18334 , n9601 );
    xnor g20463 ( n7527 , n32964 , n35310 );
    or g20464 ( n7678 , n8346 , n10693 );
    xnor g20465 ( n22801 , n2986 , n4878 );
    not g20466 ( n4809 , n27496 );
    xnor g20467 ( n19178 , n11959 , n3205 );
    nor g20468 ( n6941 , n26641 , n16649 );
    and g20469 ( n19095 , n7923 , n7317 );
    xnor g20470 ( n7688 , n30790 , n9021 );
    buf g20471 ( n28837 , n15344 );
    or g20472 ( n31326 , n8903 , n18477 );
    or g20473 ( n1243 , n7458 , n17931 );
    xnor g20474 ( n17737 , n32648 , n8097 );
    or g20475 ( n10009 , n18055 , n19609 );
    and g20476 ( n12907 , n29840 , n25235 );
    or g20477 ( n24126 , n10158 , n7417 );
    not g20478 ( n15222 , n16894 );
    or g20479 ( n27852 , n7495 , n20579 );
    xnor g20480 ( n13998 , n25118 , n20093 );
    or g20481 ( n21233 , n7503 , n19151 );
    nor g20482 ( n22037 , n32715 , n8008 );
    or g20483 ( n13430 , n23534 , n6666 );
    and g20484 ( n10031 , n35153 , n31886 );
    xnor g20485 ( n29504 , n22162 , n24027 );
    xnor g20486 ( n19607 , n29141 , n7943 );
    xnor g20487 ( n28519 , n28107 , n1955 );
    and g20488 ( n18242 , n2302 , n17015 );
    and g20489 ( n9820 , n5305 , n34951 );
    or g20490 ( n20278 , n35780 , n12829 );
    not g20491 ( n31566 , n35938 );
    or g20492 ( n31892 , n13447 , n28668 );
    and g20493 ( n29160 , n27750 , n6843 );
    and g20494 ( n20562 , n23172 , n11398 );
    or g20495 ( n33355 , n31215 , n29488 );
    not g20496 ( n8305 , n16620 );
    and g20497 ( n16934 , n28248 , n2861 );
    or g20498 ( n14645 , n26903 , n19403 );
    and g20499 ( n14866 , n7936 , n27406 );
    or g20500 ( n25840 , n15590 , n4254 );
    or g20501 ( n13980 , n9442 , n5457 );
    or g20502 ( n24316 , n932 , n26468 );
    or g20503 ( n12785 , n30036 , n3738 );
    or g20504 ( n7593 , n1950 , n28640 );
    xnor g20505 ( n19717 , n24898 , n6338 );
    or g20506 ( n25450 , n27514 , n319 );
    or g20507 ( n16412 , n15464 , n15456 );
    or g20508 ( n33975 , n1524 , n7417 );
    and g20509 ( n15381 , n19103 , n13693 );
    and g20510 ( n948 , n1354 , n20691 );
    or g20511 ( n1743 , n3205 , n15341 );
    or g20512 ( n27467 , n17352 , n4619 );
    and g20513 ( n33973 , n22546 , n11946 );
    and g20514 ( n21598 , n5849 , n1432 );
    or g20515 ( n10150 , n8838 , n24672 );
    or g20516 ( n17253 , n28986 , n31337 );
    xnor g20517 ( n18754 , n5894 , n24371 );
    or g20518 ( n14160 , n14391 , n10085 );
    or g20519 ( n18807 , n14721 , n25338 );
    xnor g20520 ( n11033 , n22817 , n18974 );
    or g20521 ( n28889 , n17311 , n2410 );
    xnor g20522 ( n30801 , n10339 , n13939 );
    or g20523 ( n18285 , n20324 , n3188 );
    and g20524 ( n23919 , n22395 , n24006 );
    nor g20525 ( n14287 , n22209 , n18115 );
    xnor g20526 ( n22512 , n20289 , n10487 );
    or g20527 ( n6261 , n6319 , n4485 );
    and g20528 ( n6139 , n17310 , n17432 );
    nor g20529 ( n14452 , n22040 , n9208 );
    or g20530 ( n11053 , n25934 , n21783 );
    or g20531 ( n30539 , n14558 , n34070 );
    not g20532 ( n13411 , n9344 );
    and g20533 ( n27004 , n34884 , n35970 );
    nor g20534 ( n27779 , n29713 , n21272 );
    or g20535 ( n35370 , n28498 , n9626 );
    and g20536 ( n1673 , n13152 , n6109 );
    xnor g20537 ( n26792 , n31072 , n3205 );
    or g20538 ( n21401 , n15520 , n19490 );
    and g20539 ( n29563 , n32513 , n22072 );
    xnor g20540 ( n3985 , n23065 , n31799 );
    or g20541 ( n18825 , n11522 , n35107 );
    not g20542 ( n16356 , n25113 );
    or g20543 ( n29321 , n16512 , n2479 );
    nor g20544 ( n14303 , n7540 , n4889 );
    or g20545 ( n21776 , n35322 , n22783 );
    xnor g20546 ( n34497 , n22701 , n17568 );
    or g20547 ( n28792 , n35927 , n23010 );
    or g20548 ( n18766 , n6466 , n20690 );
    and g20549 ( n25423 , n18662 , n4245 );
    or g20550 ( n17470 , n32749 , n1961 );
    or g20551 ( n28825 , n32584 , n22244 );
    nor g20552 ( n24164 , n4960 , n29136 );
    not g20553 ( n18514 , n16777 );
    or g20554 ( n1597 , n24371 , n28997 );
    xnor g20555 ( n8534 , n34168 , n23604 );
    and g20556 ( n27897 , n4922 , n1685 );
    or g20557 ( n20097 , n24460 , n2454 );
    not g20558 ( n27745 , n18296 );
    and g20559 ( n23711 , n29250 , n17410 );
    xnor g20560 ( n35691 , n723 , n22427 );
    or g20561 ( n26652 , n17044 , n29547 );
    or g20562 ( n2437 , n690 , n32572 );
    or g20563 ( n2302 , n19838 , n28331 );
    or g20564 ( n26096 , n31289 , n18780 );
    buf g20565 ( n33435 , n3252 );
    nor g20566 ( n29578 , n23604 , n22030 );
    or g20567 ( n9521 , n20383 , n9571 );
    or g20568 ( n5620 , n13834 , n3510 );
    xnor g20569 ( n29141 , n30468 , n4758 );
    or g20570 ( n390 , n18356 , n19241 );
    buf g20571 ( n32572 , n6255 );
    not g20572 ( n33031 , n17065 );
    or g20573 ( n26050 , n19468 , n25976 );
    or g20574 ( n4770 , n29082 , n16041 );
    or g20575 ( n20843 , n9530 , n31067 );
    xnor g20576 ( n12023 , n35948 , n17568 );
    or g20577 ( n10921 , n19984 , n6624 );
    or g20578 ( n31299 , n23336 , n2168 );
    or g20579 ( n15106 , n3076 , n18811 );
    or g20580 ( n6727 , n27980 , n3736 );
    and g20581 ( n17060 , n26430 , n19505 );
    and g20582 ( n35290 , n6839 , n22696 );
    xnor g20583 ( n1448 , n32725 , n19984 );
    or g20584 ( n3926 , n9789 , n19485 );
    nor g20585 ( n13928 , n33999 , n33685 );
    and g20586 ( n30621 , n34539 , n1031 );
    not g20587 ( n6715 , n7183 );
    or g20588 ( n27522 , n32584 , n6820 );
    or g20589 ( n9285 , n12874 , n1474 );
    xnor g20590 ( n32107 , n31082 , n21704 );
    or g20591 ( n22628 , n30702 , n21042 );
    and g20592 ( n20021 , n21448 , n17403 );
    xnor g20593 ( n28430 , n19949 , n17881 );
    or g20594 ( n8967 , n16135 , n10408 );
    or g20595 ( n15867 , n1712 , n18193 );
    or g20596 ( n19437 , n19751 , n4203 );
    xnor g20597 ( n24776 , n1139 , n4234 );
    nor g20598 ( n34216 , n14097 , n27747 );
    or g20599 ( n13013 , n29579 , n1433 );
    xnor g20600 ( n19124 , n20705 , n25725 );
    or g20601 ( n25546 , n11661 , n25475 );
    xnor g20602 ( n14660 , n1639 , n4288 );
    or g20603 ( n9000 , n9883 , n26737 );
    xnor g20604 ( n21982 , n22598 , n14356 );
    xnor g20605 ( n3533 , n33276 , n17698 );
    and g20606 ( n25013 , n5913 , n35530 );
    or g20607 ( n33283 , n30142 , n25489 );
    nor g20608 ( n2950 , n13318 , n16468 );
    xnor g20609 ( n19088 , n21079 , n30205 );
    and g20610 ( n14943 , n21095 , n28919 );
    or g20611 ( n22963 , n2035 , n16097 );
    xnor g20612 ( n15115 , n1986 , n3818 );
    and g20613 ( n4050 , n27660 , n9514 );
    xnor g20614 ( n9332 , n29475 , n20559 );
    or g20615 ( n34593 , n22703 , n28584 );
    or g20616 ( n13488 , n25111 , n7673 );
    xnor g20617 ( n24798 , n2189 , n1130 );
    or g20618 ( n26727 , n6873 , n19490 );
    or g20619 ( n13424 , n4825 , n20277 );
    or g20620 ( n8652 , n3369 , n28438 );
    nor g20621 ( n24030 , n11664 , n24565 );
    or g20622 ( n32410 , n19540 , n11241 );
    or g20623 ( n30939 , n29001 , n19135 );
    and g20624 ( n18562 , n15478 , n29463 );
    or g20625 ( n16949 , n2953 , n1026 );
    buf g20626 ( n10336 , n603 );
    and g20627 ( n26244 , n11185 , n10674 );
    or g20628 ( n19857 , n21647 , n27728 );
    or g20629 ( n30875 , n5259 , n21712 );
    xnor g20630 ( n3563 , n18514 , n15299 );
    xnor g20631 ( n4694 , n34371 , n18819 );
    xnor g20632 ( n29075 , n1261 , n26918 );
    or g20633 ( n5973 , n3222 , n2335 );
    xnor g20634 ( n17783 , n35318 , n830 );
    or g20635 ( n5943 , n3535 , n10707 );
    and g20636 ( n21547 , n31826 , n3027 );
    or g20637 ( n20468 , n20783 , n2374 );
    or g20638 ( n24459 , n19635 , n31173 );
    or g20639 ( n33075 , n11046 , n14680 );
    not g20640 ( n35107 , n10266 );
    or g20641 ( n13596 , n24295 , n23090 );
    not g20642 ( n31204 , n27050 );
    and g20643 ( n11877 , n16790 , n5191 );
    not g20644 ( n23348 , n29872 );
    or g20645 ( n21756 , n9763 , n6340 );
    and g20646 ( n897 , n1973 , n23845 );
    or g20647 ( n9192 , n34046 , n28703 );
    or g20648 ( n14738 , n31272 , n31375 );
    and g20649 ( n30563 , n31678 , n25316 );
    or g20650 ( n33083 , n4855 , n28248 );
    and g20651 ( n11790 , n34087 , n33392 );
    or g20652 ( n35367 , n32785 , n12950 );
    and g20653 ( n3483 , n27424 , n10308 );
    xnor g20654 ( n3530 , n5436 , n27624 );
    xnor g20655 ( n11612 , n12289 , n34467 );
    or g20656 ( n16428 , n16135 , n21464 );
    nor g20657 ( n34363 , n30470 , n3850 );
    buf g20658 ( n18296 , n4241 );
    not g20659 ( n33750 , n16659 );
    or g20660 ( n12256 , n3602 , n1414 );
    and g20661 ( n23212 , n10815 , n26200 );
    and g20662 ( n29647 , n34887 , n23445 );
    or g20663 ( n23216 , n25684 , n14918 );
    or g20664 ( n34616 , n32733 , n22679 );
    xnor g20665 ( n19886 , n35307 , n11455 );
    and g20666 ( n32199 , n16320 , n14490 );
    or g20667 ( n28418 , n18683 , n35339 );
    xnor g20668 ( n7754 , n24728 , n11113 );
    nor g20669 ( n25160 , n4519 , n28870 );
    or g20670 ( n25040 , n10372 , n13525 );
    or g20671 ( n9313 , n32857 , n20213 );
    or g20672 ( n17840 , n15055 , n9915 );
    not g20673 ( n5315 , n33791 );
    nor g20674 ( n6333 , n11502 , n5387 );
    xnor g20675 ( n25850 , n5020 , n5287 );
    or g20676 ( n18191 , n32515 , n20762 );
    or g20677 ( n25224 , n8628 , n13883 );
    not g20678 ( n29571 , n29713 );
    not g20679 ( n24839 , n35927 );
    or g20680 ( n13605 , n14661 , n14841 );
    nor g20681 ( n109 , n10894 , n28941 );
    xnor g20682 ( n34085 , n34447 , n25174 );
    or g20683 ( n30656 , n4950 , n28324 );
    not g20684 ( n23851 , n31177 );
    or g20685 ( n16211 , n35923 , n2010 );
    or g20686 ( n15260 , n11017 , n28502 );
    xnor g20687 ( n18697 , n16332 , n12125 );
    or g20688 ( n19156 , n34585 , n29592 );
    xnor g20689 ( n6475 , n25908 , n2256 );
    and g20690 ( n29195 , n18985 , n7027 );
    or g20691 ( n5970 , n8623 , n25036 );
    nor g20692 ( n2179 , n24981 , n35625 );
    or g20693 ( n12033 , n8413 , n16762 );
    xnor g20694 ( n6122 , n22569 , n24371 );
    or g20695 ( n2309 , n19011 , n26419 );
    not g20696 ( n3274 , n15290 );
    not g20697 ( n3142 , n24271 );
    xnor g20698 ( n121 , n21829 , n6390 );
    and g20699 ( n19949 , n23783 , n12246 );
    or g20700 ( n33381 , n34905 , n29739 );
    or g20701 ( n22726 , n31164 , n11996 );
    xnor g20702 ( n15228 , n12769 , n35647 );
    and g20703 ( n6035 , n16756 , n20801 );
    nor g20704 ( n14743 , n9789 , n13708 );
    and g20705 ( n17731 , n20187 , n20192 );
    or g20706 ( n10257 , n27078 , n2748 );
    xnor g20707 ( n19098 , n12277 , n16343 );
    and g20708 ( n25099 , n22258 , n32536 );
    xnor g20709 ( n28043 , n30492 , n31215 );
    and g20710 ( n27401 , n13258 , n15726 );
    or g20711 ( n6858 , n29713 , n1576 );
    xnor g20712 ( n15596 , n3073 , n16791 );
    and g20713 ( n29478 , n15763 , n10505 );
    xnor g20714 ( n32332 , n17002 , n23604 );
    not g20715 ( n9591 , n828 );
    xnor g20716 ( n16804 , n4061 , n7678 );
    and g20717 ( n29367 , n9762 , n27965 );
    and g20718 ( n329 , n35810 , n30068 );
    and g20719 ( n12353 , n5532 , n23400 );
    or g20720 ( n6988 , n14045 , n21037 );
    xnor g20721 ( n33347 , n12686 , n5113 );
    or g20722 ( n17296 , n10454 , n22851 );
    nor g20723 ( n11247 , n22500 , n32379 );
    or g20724 ( n5212 , n13837 , n4318 );
    or g20725 ( n5988 , n29709 , n25594 );
    xnor g20726 ( n12236 , n28462 , n11848 );
    xnor g20727 ( n20098 , n24819 , n22291 );
    or g20728 ( n22183 , n31958 , n24408 );
    xnor g20729 ( n2516 , n35855 , n9789 );
    and g20730 ( n18316 , n30937 , n11306 );
    xnor g20731 ( n16044 , n11120 , n10894 );
    and g20732 ( n715 , n26946 , n26198 );
    nor g20733 ( n32316 , n30742 , n34992 );
    or g20734 ( n8864 , n20585 , n13518 );
    or g20735 ( n17610 , n32095 , n27212 );
    not g20736 ( n32090 , n19551 );
    or g20737 ( n13555 , n17755 , n27053 );
    or g20738 ( n33700 , n12483 , n35473 );
    xnor g20739 ( n19635 , n20516 , n16922 );
    or g20740 ( n30323 , n4288 , n8311 );
    and g20741 ( n16989 , n12882 , n19427 );
    and g20742 ( n13548 , n23794 , n21564 );
    or g20743 ( n5863 , n2532 , n27191 );
    or g20744 ( n15811 , n26678 , n18253 );
    or g20745 ( n1857 , n29975 , n24489 );
    or g20746 ( n34227 , n6422 , n34746 );
    not g20747 ( n33810 , n28807 );
    or g20748 ( n15315 , n28385 , n28240 );
    or g20749 ( n9864 , n20925 , n31134 );
    not g20750 ( n31184 , n18296 );
    and g20751 ( n22159 , n25874 , n11994 );
    xnor g20752 ( n34051 , n26524 , n25765 );
    or g20753 ( n5984 , n34566 , n15677 );
    or g20754 ( n33744 , n26580 , n33265 );
    and g20755 ( n19291 , n74 , n22444 );
    xnor g20756 ( n9032 , n22047 , n17568 );
    and g20757 ( n31589 , n32410 , n32734 );
    xnor g20758 ( n24715 , n21995 , n7851 );
    or g20759 ( n26405 , n4247 , n6470 );
    and g20760 ( n4763 , n892 , n13899 );
    and g20761 ( n2207 , n12741 , n16651 );
    or g20762 ( n11180 , n25602 , n10544 );
    and g20763 ( n27008 , n33937 , n33828 );
    nor g20764 ( n22346 , n25602 , n11859 );
    or g20765 ( n1594 , n20518 , n28240 );
    or g20766 ( n20431 , n15464 , n24941 );
    or g20767 ( n32512 , n22962 , n27996 );
    not g20768 ( n11739 , n29470 );
    nor g20769 ( n29885 , n35385 , n19834 );
    xnor g20770 ( n29864 , n13520 , n3222 );
    or g20771 ( n18515 , n16922 , n11881 );
    xnor g20772 ( n9002 , n22334 , n33863 );
    or g20773 ( n22506 , n30742 , n5195 );
    xnor g20774 ( n7028 , n20443 , n19551 );
    xnor g20775 ( n10508 , n28212 , n32095 );
    xnor g20776 ( n13101 , n6539 , n10212 );
    not g20777 ( n27851 , n8388 );
    xnor g20778 ( n11446 , n20636 , n830 );
    and g20779 ( n13035 , n19627 , n1226 );
    buf g20780 ( n12913 , n7448 );
    xnor g20781 ( n23522 , n7150 , n8731 );
    or g20782 ( n29026 , n20311 , n7147 );
    not g20783 ( n28493 , n17396 );
    or g20784 ( n24708 , n16620 , n15671 );
    nor g20785 ( n6994 , n1429 , n21043 );
    xnor g20786 ( n17658 , n2483 , n20021 );
    or g20787 ( n15027 , n11046 , n10075 );
    xnor g20788 ( n27647 , n4890 , n34017 );
    and g20789 ( n6565 , n23977 , n30090 );
    xnor g20790 ( n32401 , n33099 , n30742 );
    xnor g20791 ( n25697 , n367 , n13021 );
    and g20792 ( n14445 , n31970 , n379 );
    or g20793 ( n32922 , n12838 , n11295 );
    xnor g20794 ( n24246 , n12707 , n30762 );
    xnor g20795 ( n14047 , n3579 , n29277 );
    or g20796 ( n4453 , n31992 , n3 );
    nor g20797 ( n33543 , n13545 , n25171 );
    not g20798 ( n31389 , n20045 );
    not g20799 ( n9394 , n8865 );
    and g20800 ( n35623 , n34392 , n15483 );
    xnor g20801 ( n17718 , n30207 , n4531 );
    or g20802 ( n9151 , n1618 , n23323 );
    or g20803 ( n22253 , n1054 , n28314 );
    or g20804 ( n191 , n0 , n29441 );
    or g20805 ( n29503 , n23362 , n3842 );
    nor g20806 ( n20588 , n32857 , n3485 );
    xnor g20807 ( n16761 , n18708 , n7891 );
    or g20808 ( n9455 , n19097 , n10140 );
    xnor g20809 ( n28960 , n25519 , n17878 );
    not g20810 ( n19121 , n32794 );
    or g20811 ( n11272 , n14816 , n26737 );
    buf g20812 ( n12996 , n30292 );
    or g20813 ( n3811 , n2573 , n139 );
    and g20814 ( n34687 , n25751 , n24314 );
    and g20815 ( n13915 , n34241 , n10828 );
    nor g20816 ( n3852 , n1891 , n18115 );
    or g20817 ( n32377 , n3229 , n30216 );
    or g20818 ( n15134 , n23604 , n30084 );
    or g20819 ( n10931 , n24371 , n23333 );
    xnor g20820 ( n30800 , n31407 , n30198 );
    xnor g20821 ( n20214 , n35607 , n10484 );
    xnor g20822 ( n23992 , n35722 , n17568 );
    and g20823 ( n7265 , n5666 , n9759 );
    or g20824 ( n32317 , n1228 , n7647 );
    and g20825 ( n28453 , n30469 , n5011 );
    xnor g20826 ( n12423 , n2973 , n2653 );
    or g20827 ( n7923 , n32561 , n12873 );
    or g20828 ( n6879 , n18919 , n31067 );
    or g20829 ( n26914 , n15105 , n27116 );
    and g20830 ( n18318 , n34146 , n27286 );
    not g20831 ( n24124 , n3805 );
    nor g20832 ( n8972 , n15951 , n7327 );
    and g20833 ( n20457 , n12428 , n32386 );
    and g20834 ( n26103 , n21221 , n30323 );
    not g20835 ( n15295 , n26907 );
    nor g20836 ( n3779 , n5738 , n30993 );
    or g20837 ( n33212 , n4947 , n4206 );
    xnor g20838 ( n23551 , n36038 , n4960 );
    and g20839 ( n20244 , n6420 , n30510 );
    not g20840 ( n10115 , n29713 );
    and g20841 ( n19733 , n11044 , n35070 );
    or g20842 ( n28373 , n19991 , n34484 );
    or g20843 ( n5050 , n15716 , n24479 );
    or g20844 ( n3667 , n4288 , n9183 );
    xnor g20845 ( n23970 , n3931 , n32095 );
    or g20846 ( n14513 , n15900 , n18845 );
    nor g20847 ( n19359 , n19551 , n13667 );
    xnor g20848 ( n28228 , n21606 , n3222 );
    xnor g20849 ( n8938 , n9637 , n7540 );
    and g20850 ( n35432 , n18384 , n27236 );
    xnor g20851 ( n26156 , n7003 , n31799 );
    and g20852 ( n23410 , n7463 , n654 );
    or g20853 ( n34471 , n27559 , n12096 );
    xnor g20854 ( n29876 , n19990 , n9730 );
    xnor g20855 ( n3814 , n18015 , n3946 );
    or g20856 ( n15453 , n5335 , n32529 );
    xnor g20857 ( n28058 , n29912 , n18265 );
    or g20858 ( n12936 , n20438 , n28668 );
    or g20859 ( n3912 , n8576 , n25592 );
    not g20860 ( n26811 , n6596 );
    xnor g20861 ( n18648 , n688 , n7087 );
    xnor g20862 ( n154 , n30530 , n23604 );
    and g20863 ( n26404 , n22669 , n33258 );
    or g20864 ( n31468 , n4878 , n32603 );
    or g20865 ( n123 , n8597 , n27963 );
    and g20866 ( n15085 , n8751 , n22556 );
    nor g20867 ( n35806 , n23604 , n20465 );
    xnor g20868 ( n20225 , n1827 , n8174 );
    or g20869 ( n13982 , n22527 , n9840 );
    or g20870 ( n531 , n3205 , n23919 );
    and g20871 ( n35802 , n35025 , n29947 );
    nor g20872 ( n35288 , n652 , n27447 );
    not g20873 ( n30940 , n2092 );
    nor g20874 ( n21381 , n27291 , n1252 );
    or g20875 ( n8138 , n4960 , n14827 );
    xnor g20876 ( n25266 , n14965 , n33381 );
    or g20877 ( n12870 , n4878 , n1093 );
    or g20878 ( n15382 , n14592 , n15538 );
    and g20879 ( n22081 , n24878 , n58 );
    xnor g20880 ( n4583 , n12696 , n5089 );
    xnor g20881 ( n12330 , n26624 , n5403 );
    or g20882 ( n15627 , n16715 , n27447 );
    xnor g20883 ( n34049 , n7199 , n10537 );
    or g20884 ( n35251 , n8632 , n24345 );
    or g20885 ( n9662 , n8984 , n5208 );
    xnor g20886 ( n22117 , n9010 , n4288 );
    or g20887 ( n6882 , n34618 , n31606 );
    or g20888 ( n8521 , n24332 , n14585 );
    and g20889 ( n23183 , n8922 , n29099 );
    buf g20890 ( n34865 , n32329 );
    not g20891 ( n30619 , n13421 );
    and g20892 ( n2251 , n19595 , n19795 );
    and g20893 ( n25249 , n16104 , n20026 );
    and g20894 ( n26529 , n30074 , n211 );
    and g20895 ( n1393 , n7549 , n13918 );
    not g20896 ( n29104 , n10191 );
    or g20897 ( n34353 , n4398 , n24465 );
    or g20898 ( n13602 , n35465 , n19421 );
    xnor g20899 ( n2089 , n29391 , n32584 );
    and g20900 ( n14138 , n28370 , n23911 );
    not g20901 ( n3936 , n15290 );
    or g20902 ( n32640 , n9658 , n9910 );
    or g20903 ( n13330 , n15464 , n23749 );
    xnor g20904 ( n3114 , n10491 , n5005 );
    not g20905 ( n11751 , n24026 );
    or g20906 ( n14799 , n4962 , n25912 );
    or g20907 ( n32791 , n31289 , n32559 );
    or g20908 ( n440 , n21995 , n8392 );
    and g20909 ( n9867 , n17386 , n4181 );
    not g20910 ( n34036 , n12428 );
    and g20911 ( n34762 , n4577 , n3240 );
    not g20912 ( n25715 , n12132 );
    or g20913 ( n34570 , n15558 , n22746 );
    xnor g20914 ( n29079 , n18574 , n12228 );
    or g20915 ( n14462 , n25243 , n8090 );
    not g20916 ( n19507 , n21461 );
    or g20917 ( n28821 , n21916 , n24653 );
    or g20918 ( n1780 , n31070 , n12879 );
    xnor g20919 ( n5162 , n9961 , n11046 );
    not g20920 ( n15215 , n2092 );
    and g20921 ( n19750 , n29251 , n5871 );
    xnor g20922 ( n7161 , n20514 , n7261 );
    or g20923 ( n21972 , n35557 , n27501 );
    or g20924 ( n30726 , n22291 , n35967 );
    or g20925 ( n15423 , n9985 , n9631 );
    or g20926 ( n28718 , n17568 , n22799 );
    and g20927 ( n6427 , n3706 , n2934 );
    nor g20928 ( n1374 , n16155 , n7175 );
    or g20929 ( n23267 , n22291 , n7745 );
    xnor g20930 ( n29583 , n3100 , n15464 );
    and g20931 ( n9409 , n2741 , n29905 );
    or g20932 ( n21750 , n1349 , n10550 );
    or g20933 ( n21556 , n11031 , n20690 );
    xnor g20934 ( n27279 , n32156 , n20133 );
    or g20935 ( n962 , n5560 , n15194 );
    xnor g20936 ( n28195 , n3485 , n11782 );
    or g20937 ( n30371 , n29677 , n12128 );
    and g20938 ( n8478 , n34598 , n21865 );
    nor g20939 ( n9046 , n33899 , n22305 );
    or g20940 ( n19981 , n649 , n31552 );
    not g20941 ( n15255 , n23604 );
    and g20942 ( n26539 , n25446 , n20224 );
    or g20943 ( n975 , n8186 , n9675 );
    or g20944 ( n33506 , n3222 , n22626 );
    and g20945 ( n24900 , n25505 , n26750 );
    and g20946 ( n2726 , n14505 , n9974 );
    and g20947 ( n4818 , n6000 , n18211 );
    or g20948 ( n30193 , n16084 , n13526 );
    nor g20949 ( n13043 , n4878 , n980 );
    and g20950 ( n34990 , n34651 , n24830 );
    or g20951 ( n18342 , n29839 , n31948 );
    and g20952 ( n9730 , n15709 , n3898 );
    and g20953 ( n26313 , n24036 , n16878 );
    xnor g20954 ( n4926 , n1312 , n35927 );
    or g20955 ( n934 , n5543 , n35504 );
    xnor g20956 ( n1540 , n32611 , n11599 );
    xnor g20957 ( n11523 , n6533 , n32539 );
    nor g20958 ( n20783 , n26275 , n33956 );
    or g20959 ( n2850 , n16244 , n8723 );
    or g20960 ( n25339 , n13674 , n9440 );
    or g20961 ( n9180 , n31799 , n18043 );
    or g20962 ( n432 , n13148 , n3694 );
    or g20963 ( n20940 , n15360 , n27356 );
    and g20964 ( n9800 , n3608 , n33893 );
    or g20965 ( n19929 , n25267 , n30431 );
    or g20966 ( n13860 , n20945 , n6017 );
    and g20967 ( n14901 , n28959 , n26368 );
    or g20968 ( n45 , n31416 , n18615 );
    not g20969 ( n17668 , n23280 );
    xnor g20970 ( n4177 , n4746 , n11844 );
    xnor g20971 ( n30270 , n34867 , n10894 );
    and g20972 ( n425 , n708 , n31644 );
    or g20973 ( n1966 , n23604 , n33326 );
    xnor g20974 ( n34187 , n941 , n3004 );
    or g20975 ( n16476 , n22739 , n27728 );
    xnor g20976 ( n26358 , n33189 , n10894 );
    nor g20977 ( n13499 , n16971 , n7339 );
    xnor g20978 ( n13662 , n30985 , n32095 );
    or g20979 ( n30860 , n502 , n26458 );
    or g20980 ( n18890 , n2346 , n32537 );
    or g20981 ( n24071 , n2525 , n14554 );
    xnor g20982 ( n8753 , n2686 , n14226 );
    xnor g20983 ( n26068 , n10285 , n29713 );
    or g20984 ( n34246 , n7444 , n3891 );
    or g20985 ( n29663 , n6755 , n31902 );
    not g20986 ( n29061 , n26538 );
    or g20987 ( n18590 , n31322 , n15329 );
    and g20988 ( n24861 , n16791 , n3073 );
    or g20989 ( n12041 , n3946 , n29117 );
    and g20990 ( n31715 , n29307 , n32306 );
    xnor g20991 ( n33536 , n1850 , n11128 );
    and g20992 ( n13520 , n32713 , n24253 );
    and g20993 ( n3968 , n12634 , n22857 );
    buf g20994 ( n28574 , n12436 );
    and g20995 ( n15263 , n17048 , n22468 );
    not g20996 ( n5538 , n25592 );
    xnor g20997 ( n649 , n7385 , n25602 );
    or g20998 ( n23571 , n24267 , n29106 );
    and g20999 ( n1755 , n843 , n25719 );
    or g21000 ( n29443 , n2066 , n28868 );
    xnor g21001 ( n31294 , n8372 , n23066 );
    and g21002 ( n30610 , n18112 , n385 );
    xnor g21003 ( n20833 , n20477 , n19338 );
    and g21004 ( n5076 , n7524 , n26394 );
    or g21005 ( n24830 , n830 , n4771 );
    and g21006 ( n35667 , n23234 , n6788 );
    or g21007 ( n26494 , n32056 , n11295 );
    or g21008 ( n14213 , n8432 , n25878 );
    not g21009 ( n34546 , n33830 );
    or g21010 ( n21646 , n16450 , n28404 );
    and g21011 ( n1447 , n13180 , n9707 );
    xnor g21012 ( n32906 , n70 , n35900 );
    or g21013 ( n20744 , n8074 , n26112 );
    or g21014 ( n33970 , n4288 , n35772 );
    and g21015 ( n7485 , n22460 , n20879 );
    xnor g21016 ( n1356 , n22222 , n3946 );
    or g21017 ( n22741 , n21160 , n4081 );
    or g21018 ( n5454 , n3890 , n35043 );
    or g21019 ( n21181 , n18834 , n19776 );
    or g21020 ( n23381 , n13485 , n29843 );
    not g21021 ( n25389 , n2827 );
    or g21022 ( n19296 , n2899 , n35230 );
    and g21023 ( n16244 , n26307 , n8754 );
    and g21024 ( n35852 , n14227 , n16312 );
    and g21025 ( n8539 , n23931 , n29849 );
    not g21026 ( n23179 , n7435 );
    xnor g21027 ( n12213 , n1498 , n13464 );
    buf g21028 ( n23626 , n22561 );
    or g21029 ( n30781 , n28451 , n35111 );
    nor g21030 ( n22201 , n31289 , n30488 );
    and g21031 ( n8833 , n30874 , n19938 );
    nor g21032 ( n27445 , n16620 , n4629 );
    xnor g21033 ( n468 , n15358 , n9789 );
    xnor g21034 ( n34151 , n27109 , n1371 );
    nor g21035 ( n806 , n33103 , n32379 );
    xnor g21036 ( n1754 , n5932 , n7665 );
    or g21037 ( n33343 , n7540 , n18195 );
    or g21038 ( n35166 , n5112 , n5252 );
    xnor g21039 ( n27104 , n15286 , n32797 );
    and g21040 ( n27696 , n28805 , n11915 );
    and g21041 ( n23112 , n24087 , n6766 );
    nor g21042 ( n18737 , n20494 , n13935 );
    and g21043 ( n5170 , n11212 , n30801 );
    not g21044 ( n665 , n1409 );
    or g21045 ( n5031 , n3222 , n899 );
    and g21046 ( n26632 , n25623 , n30592 );
    or g21047 ( n2840 , n31289 , n12944 );
    nor g21048 ( n32826 , n31590 , n11831 );
    and g21049 ( n22192 , n4101 , n3464 );
    or g21050 ( n33839 , n6402 , n20308 );
    or g21051 ( n13964 , n19026 , n8549 );
    xnor g21052 ( n28320 , n4858 , n31289 );
    or g21053 ( n19759 , n27291 , n34414 );
    not g21054 ( n22794 , n9232 );
    and g21055 ( n18968 , n10554 , n32207 );
    xnor g21056 ( n25520 , n14009 , n19551 );
    or g21057 ( n15493 , n22809 , n16697 );
    xnor g21058 ( n27341 , n31507 , n27291 );
    and g21059 ( n24194 , n21838 , n32460 );
    nor g21060 ( n7025 , n3951 , n3754 );
    or g21061 ( n1636 , n30429 , n4363 );
    and g21062 ( n16598 , n26057 , n16092 );
    and g21063 ( n18423 , n4674 , n17262 );
    and g21064 ( n16652 , n34699 , n14926 );
    xnor g21065 ( n14603 , n14658 , n17951 );
    and g21066 ( n5523 , n15901 , n20549 );
    or g21067 ( n7536 , n6119 , n31596 );
    or g21068 ( n14422 , n16620 , n16370 );
    or g21069 ( n27137 , n8584 , n544 );
    xnor g21070 ( n16578 , n16857 , n427 );
    or g21071 ( n20248 , n27127 , n23323 );
    or g21072 ( n17914 , n17536 , n25019 );
    not g21073 ( n23347 , n13 );
    xnor g21074 ( n26389 , n5723 , n24371 );
    and g21075 ( n17075 , n20150 , n21698 );
    or g21076 ( n15920 , n16885 , n30732 );
    nor g21077 ( n29268 , n32584 , n26608 );
    and g21078 ( n24005 , n34766 , n33133 );
    and g21079 ( n7529 , n8322 , n15759 );
    xnor g21080 ( n35311 , n22188 , n558 );
    xnor g21081 ( n25808 , n24607 , n29629 );
    and g21082 ( n15361 , n24747 , n27867 );
    or g21083 ( n21695 , n8974 , n28866 );
    not g21084 ( n14143 , n30381 );
    not g21085 ( n34560 , n6490 );
    and g21086 ( n27077 , n9089 , n15627 );
    and g21087 ( n7086 , n35248 , n14972 );
    or g21088 ( n21005 , n8151 , n18264 );
    and g21089 ( n30993 , n1080 , n6330 );
    or g21090 ( n33553 , n7701 , n3979 );
    not g21091 ( n33287 , n22200 );
    and g21092 ( n388 , n22181 , n14799 );
    or g21093 ( n27662 , n29346 , n31923 );
    or g21094 ( n32369 , n19127 , n35971 );
    xnor g21095 ( n13798 , n31284 , n4288 );
    or g21096 ( n32415 , n15388 , n5457 );
    and g21097 ( n6259 , n31905 , n32032 );
    and g21098 ( n22713 , n13401 , n11086 );
    or g21099 ( n3131 , n11858 , n1856 );
    nor g21100 ( n9363 , n9789 , n22777 );
    or g21101 ( n6492 , n32445 , n7945 );
    xnor g21102 ( n761 , n32890 , n35253 );
    or g21103 ( n35083 , n8829 , n8796 );
    xnor g21104 ( n11329 , n15982 , n10894 );
    or g21105 ( n6058 , n15464 , n20541 );
    or g21106 ( n34515 , n3376 , n18970 );
    or g21107 ( n26150 , n1120 , n12515 );
    nor g21108 ( n33986 , n35401 , n15849 );
    xor g21109 ( n33103 , n20501 , n34756 );
    nor g21110 ( n5544 , n19018 , n12996 );
    not g21111 ( n23453 , n13319 );
    or g21112 ( n4272 , n5078 , n28192 );
    or g21113 ( n33209 , n1913 , n18874 );
    xnor g21114 ( n23514 , n11042 , n4878 );
    or g21115 ( n21971 , n6399 , n780 );
    or g21116 ( n28484 , n18782 , n12089 );
    xnor g21117 ( n5745 , n17786 , n2621 );
    and g21118 ( n7577 , n34890 , n12918 );
    or g21119 ( n29902 , n21765 , n34626 );
    or g21120 ( n33903 , n19599 , n22682 );
    or g21121 ( n3410 , n15047 , n33435 );
    xnor g21122 ( n35256 , n19104 , n24332 );
    and g21123 ( n20188 , n5133 , n8939 );
    or g21124 ( n10089 , n35232 , n16518 );
    or g21125 ( n34160 , n24534 , n22501 );
    and g21126 ( n21213 , n26734 , n2571 );
    or g21127 ( n10051 , n10522 , n27973 );
    and g21128 ( n3050 , n31713 , n5237 );
    or g21129 ( n10582 , n2963 , n7427 );
    and g21130 ( n9345 , n495 , n18308 );
    and g21131 ( n13204 , n16090 , n22980 );
    buf g21132 ( n3352 , n17793 );
    not g21133 ( n4053 , n20644 );
    and g21134 ( n27615 , n31978 , n27916 );
    or g21135 ( n23480 , n26211 , n15256 );
    and g21136 ( n29830 , n16460 , n33857 );
    not g21137 ( n553 , n11904 );
    or g21138 ( n2828 , n17230 , n4570 );
    or g21139 ( n22772 , n8705 , n14249 );
    and g21140 ( n9005 , n33793 , n22980 );
    xnor g21141 ( n7078 , n11728 , n1351 );
    and g21142 ( n18745 , n30919 , n28777 );
    or g21143 ( n3272 , n5877 , n8723 );
    not g21144 ( n19845 , n11633 );
    or g21145 ( n16372 , n29683 , n28455 );
    or g21146 ( n22627 , n9658 , n12565 );
    xnor g21147 ( n7480 , n26532 , n22192 );
    or g21148 ( n6722 , n17322 , n28648 );
    xnor g21149 ( n22043 , n11822 , n16123 );
    or g21150 ( n17280 , n34443 , n32260 );
    or g21151 ( n14758 , n32727 , n16464 );
    and g21152 ( n11269 , n8861 , n9439 );
    and g21153 ( n5864 , n8689 , n17700 );
    or g21154 ( n31260 , n27095 , n26659 );
    xnor g21155 ( n7829 , n15505 , n12464 );
    or g21156 ( n20476 , n3222 , n14340 );
    or g21157 ( n28782 , n781 , n14706 );
    or g21158 ( n20373 , n4962 , n30045 );
    and g21159 ( n31487 , n23316 , n17631 );
    or g21160 ( n6515 , n21463 , n19336 );
    or g21161 ( n36037 , n5093 , n11833 );
    not g21162 ( n22255 , n16831 );
    not g21163 ( n16603 , n35479 );
    nor g21164 ( n24942 , n29713 , n9605 );
    and g21165 ( n25608 , n14961 , n8444 );
    or g21166 ( n11733 , n25174 , n19772 );
    and g21167 ( n11548 , n5431 , n25994 );
    nor g21168 ( n20002 , n13691 , n30077 );
    and g21169 ( n13769 , n32100 , n2519 );
    not g21170 ( n14540 , n13744 );
    xnor g21171 ( n28227 , n26702 , n28522 );
    or g21172 ( n14664 , n24857 , n28104 );
    or g21173 ( n29198 , n22170 , n30650 );
    and g21174 ( n17360 , n10312 , n23575 );
    xnor g21175 ( n18114 , n29647 , n15299 );
    or g21176 ( n297 , n13826 , n35027 );
    and g21177 ( n11205 , n13627 , n31224 );
    and g21178 ( n16924 , n24597 , n10193 );
    or g21179 ( n28670 , n11528 , n11850 );
    or g21180 ( n1588 , n31442 , n14586 );
    and g21181 ( n25558 , n20153 , n13356 );
    or g21182 ( n9050 , n14099 , n20812 );
    xnor g21183 ( n28485 , n32907 , n239 );
    xnor g21184 ( n19460 , n33012 , n30035 );
    or g21185 ( n10949 , n10894 , n3897 );
    not g21186 ( n33006 , n2861 );
    xnor g21187 ( n12342 , n35431 , n28900 );
    xnor g21188 ( n1553 , n3045 , n31848 );
    and g21189 ( n34811 , n4227 , n6993 );
    or g21190 ( n25656 , n34847 , n19955 );
    or g21191 ( n34457 , n11446 , n8398 );
    or g21192 ( n28290 , n29603 , n33034 );
    xnor g21193 ( n28877 , n23511 , n4217 );
    or g21194 ( n8689 , n1161 , n24505 );
    or g21195 ( n12604 , n29713 , n4938 );
    buf g21196 ( n22858 , n26365 );
    and g21197 ( n28252 , n27784 , n14016 );
    and g21198 ( n25127 , n12651 , n32307 );
    and g21199 ( n7547 , n6953 , n29301 );
    or g21200 ( n9982 , n17633 , n35111 );
    xnor g21201 ( n917 , n9838 , n4758 );
    or g21202 ( n23845 , n4711 , n34923 );
    or g21203 ( n19491 , n34050 , n23565 );
    or g21204 ( n35726 , n25602 , n7014 );
    xnor g21205 ( n36015 , n14683 , n32095 );
    not g21206 ( n32855 , n12612 );
    or g21207 ( n28961 , n10894 , n9647 );
    or g21208 ( n8653 , n19327 , n17859 );
    xnor g21209 ( n28494 , n10553 , n5287 );
    not g21210 ( n23028 , n2805 );
    or g21211 ( n26674 , n4858 , n24259 );
    and g21212 ( n2446 , n20321 , n17644 );
    or g21213 ( n30500 , n3946 , n6183 );
    nor g21214 ( n25712 , n7424 , n759 );
    nor g21215 ( n11323 , n31289 , n15740 );
    xnor g21216 ( n13414 , n23542 , n1050 );
    or g21217 ( n26798 , n4962 , n15900 );
    or g21218 ( n29598 , n19255 , n18542 );
    and g21219 ( n20402 , n29986 , n21730 );
    or g21220 ( n11811 , n4962 , n10269 );
    and g21221 ( n8369 , n27543 , n22023 );
    buf g21222 ( n20817 , n18488 );
    or g21223 ( n30453 , n3901 , n7361 );
    or g21224 ( n950 , n35640 , n23943 );
    and g21225 ( n12554 , n13022 , n14522 );
    and g21226 ( n29993 , n18505 , n25502 );
    or g21227 ( n18547 , n18380 , n6194 );
    and g21228 ( n169 , n17843 , n2908 );
    or g21229 ( n25278 , n12417 , n4478 );
    or g21230 ( n32062 , n19711 , n19490 );
    xnor g21231 ( n23509 , n11002 , n946 );
    xnor g21232 ( n27238 , n15361 , n27226 );
    nor g21233 ( n10556 , n17091 , n26578 );
    or g21234 ( n17077 , n15512 , n15805 );
    or g21235 ( n17488 , n28972 , n25255 );
    or g21236 ( n30248 , n8420 , n27490 );
    and g21237 ( n25166 , n10539 , n35860 );
    xnor g21238 ( n16023 , n2628 , n16673 );
    or g21239 ( n26824 , n20353 , n2600 );
    xnor g21240 ( n35377 , n2545 , n23533 );
    and g21241 ( n30953 , n7579 , n10806 );
    and g21242 ( n20577 , n26955 , n20354 );
    xnor g21243 ( n27090 , n27154 , n30553 );
    or g21244 ( n21812 , n16159 , n441 );
    not g21245 ( n15350 , n1528 );
    or g21246 ( n27545 , n12677 , n17337 );
    and g21247 ( n4976 , n16277 , n15470 );
    and g21248 ( n18780 , n9976 , n4155 );
    or g21249 ( n32606 , n21826 , n34614 );
    nor g21250 ( n23529 , n13479 , n32874 );
    or g21251 ( n693 , n19497 , n20690 );
    or g21252 ( n16477 , n25602 , n5275 );
    not g21253 ( n35310 , n16620 );
    or g21254 ( n25403 , n1244 , n6018 );
    nor g21255 ( n32280 , n24034 , n12100 );
    or g21256 ( n5121 , n35912 , n16499 );
    nor g21257 ( n34760 , n31799 , n9693 );
    xnor g21258 ( n11550 , n31926 , n32682 );
    xnor g21259 ( n6449 , n5794 , n19984 );
    or g21260 ( n21600 , n15284 , n12465 );
    or g21261 ( n22284 , n3389 , n24259 );
    xnor g21262 ( n2970 , n11914 , n32715 );
    not g21263 ( n5455 , n16620 );
    nor g21264 ( n26411 , n11182 , n23564 );
    or g21265 ( n11764 , n33665 , n26468 );
    and g21266 ( n31949 , n23341 , n22770 );
    xnor g21267 ( n3116 , n20627 , n28232 );
    and g21268 ( n15991 , n11494 , n9142 );
    not g21269 ( n26577 , n24371 );
    or g21270 ( n32868 , n4151 , n5972 );
    or g21271 ( n5014 , n22341 , n8735 );
    or g21272 ( n34957 , n32857 , n32825 );
    and g21273 ( n3388 , n8483 , n21503 );
    xnor g21274 ( n9627 , n20072 , n8432 );
    or g21275 ( n9212 , n15065 , n20840 );
    or g21276 ( n20707 , n9658 , n23574 );
    xnor g21277 ( n22341 , n32 , n11455 );
    buf g21278 ( n9194 , n3325 );
    and g21279 ( n17450 , n32630 , n20261 );
    and g21280 ( n22959 , n9395 , n5480 );
    xnor g21281 ( n35022 , n32950 , n32095 );
    nor g21282 ( n31002 , n31559 , n17671 );
    not g21283 ( n26022 , n18296 );
    xnor g21284 ( n22558 , n25035 , n3205 );
    and g21285 ( n1229 , n10395 , n27697 );
    and g21286 ( n15358 , n12066 , n14216 );
    xnor g21287 ( n30522 , n21048 , n35922 );
    not g21288 ( n19367 , n31209 );
    or g21289 ( n25062 , n35349 , n33462 );
    or g21290 ( n10169 , n24875 , n15496 );
    not g21291 ( n32967 , n17359 );
    nor g21292 ( n33466 , n29151 , n16717 );
    or g21293 ( n33055 , n15263 , n24333 );
    or g21294 ( n19745 , n31080 , n28191 );
    and g21295 ( n28591 , n8393 , n14255 );
    and g21296 ( n35716 , n15888 , n19548 );
    not g21297 ( n16763 , n26526 );
    nor g21298 ( n1913 , n31799 , n9692 );
    not g21299 ( n28507 , n16223 );
    and g21300 ( n14586 , n30196 , n28534 );
    or g21301 ( n1914 , n536 , n9555 );
    or g21302 ( n35968 , n31559 , n22891 );
    xnor g21303 ( n34008 , n28049 , n12717 );
    buf g21304 ( n33416 , n5713 );
    or g21305 ( n22995 , n17568 , n3463 );
    xnor g21306 ( n13050 , n30566 , n26195 );
    and g21307 ( n29516 , n19227 , n10768 );
    nor g21308 ( n22379 , n2548 , n6548 );
    and g21309 ( n33752 , n13131 , n7848 );
    xnor g21310 ( n29536 , n21096 , n5279 );
    not g21311 ( n33581 , n30586 );
    not g21312 ( n18495 , n4962 );
    or g21313 ( n6016 , n830 , n15213 );
    and g21314 ( n13037 , n15186 , n31097 );
    xnor g21315 ( n28307 , n1403 , n830 );
    or g21316 ( n12153 , n22723 , n13480 );
    or g21317 ( n5778 , n27795 , n30134 );
    or g21318 ( n10975 , n26899 , n34864 );
    or g21319 ( n12425 , n16146 , n2432 );
    and g21320 ( n13925 , n3201 , n8249 );
    not g21321 ( n16014 , n25830 );
    xnor g21322 ( n18999 , n30473 , n5355 );
    or g21323 ( n31971 , n33185 , n20601 );
    and g21324 ( n28608 , n12085 , n26452 );
    or g21325 ( n9231 , n9943 , n19732 );
    or g21326 ( n33141 , n5930 , n31532 );
    or g21327 ( n15252 , n12653 , n27872 );
    and g21328 ( n30851 , n13273 , n17809 );
    or g21329 ( n4623 , n25195 , n34862 );
    or g21330 ( n315 , n11437 , n34084 );
    or g21331 ( n25158 , n10488 , n9672 );
    or g21332 ( n34453 , n26692 , n11518 );
    not g21333 ( n33076 , n8386 );
    not g21334 ( n28778 , n20558 );
    and g21335 ( n34518 , n12425 , n4782 );
    buf g21336 ( n26931 , n26365 );
    xnor g21337 ( n4223 , n16711 , n11046 );
    or g21338 ( n6467 , n13285 , n21757 );
    or g21339 ( n7190 , n2141 , n10356 );
    xnor g21340 ( n15054 , n31486 , n876 );
    nor g21341 ( n29985 , n29713 , n28695 );
    xnor g21342 ( n11419 , n31416 , n18615 );
    or g21343 ( n5271 , n15288 , n33257 );
    xnor g21344 ( n21897 , n9446 , n15790 );
    and g21345 ( n22668 , n25844 , n29766 );
    or g21346 ( n20028 , n34719 , n1414 );
    xnor g21347 ( n12822 , n4972 , n9617 );
    or g21348 ( n14419 , n4122 , n7692 );
    or g21349 ( n10388 , n10894 , n35587 );
    xnor g21350 ( n21834 , n24546 , n18711 );
    or g21351 ( n19426 , n32896 , n13465 );
    xnor g21352 ( n4418 , n4414 , n10603 );
    or g21353 ( n31160 , n12003 , n9030 );
    or g21354 ( n31726 , n24380 , n11605 );
    not g21355 ( n24998 , n29649 );
    buf g21356 ( n35111 , n34048 );
    or g21357 ( n2234 , n33101 , n28586 );
    and g21358 ( n734 , n7825 , n6158 );
    or g21359 ( n1224 , n23848 , n27574 );
    not g21360 ( n3577 , n30459 );
    and g21361 ( n2293 , n26789 , n22331 );
    or g21362 ( n20449 , n15886 , n29821 );
    or g21363 ( n14157 , n25084 , n15394 );
    or g21364 ( n14210 , n25764 , n10432 );
    and g21365 ( n32130 , n8381 , n15095 );
    or g21366 ( n22408 , n32678 , n3104 );
    and g21367 ( n30652 , n32795 , n34487 );
    or g21368 ( n12365 , n8432 , n7812 );
    xnor g21369 ( n19127 , n25292 , n25602 );
    or g21370 ( n18852 , n3660 , n27963 );
    or g21371 ( n32387 , n30560 , n35591 );
    and g21372 ( n31087 , n14932 , n4812 );
    xnor g21373 ( n36068 , n2047 , n9793 );
    or g21374 ( n11073 , n35927 , n32465 );
    not g21375 ( n3799 , n24263 );
    or g21376 ( n12963 , n4125 , n7553 );
    or g21377 ( n18464 , n7540 , n6569 );
    or g21378 ( n2969 , n24544 , n27963 );
    xnor g21379 ( n32965 , n32092 , n32857 );
    or g21380 ( n1828 , n1152 , n27963 );
    and g21381 ( n837 , n30743 , n9131 );
    xnor g21382 ( n28676 , n22918 , n19399 );
    or g21383 ( n7783 , n18710 , n27053 );
    or g21384 ( n14733 , n28765 , n34084 );
    nor g21385 ( n32473 , n30629 , n33956 );
    xnor g21386 ( n31156 , n34203 , n21305 );
    not g21387 ( n34208 , n11190 );
    and g21388 ( n8480 , n22004 , n14755 );
    and g21389 ( n23736 , n19388 , n3726 );
    xnor g21390 ( n29574 , n25998 , n29771 );
    or g21391 ( n7596 , n20059 , n9317 );
    or g21392 ( n11149 , n32157 , n17125 );
    xnor g21393 ( n21120 , n3838 , n31799 );
    xnor g21394 ( n13715 , n17382 , n2064 );
    or g21395 ( n19224 , n4026 , n10417 );
    or g21396 ( n5188 , n7297 , n12317 );
    not g21397 ( n20996 , n17674 );
    or g21398 ( n14900 , n27160 , n34472 );
    and g21399 ( n4495 , n6860 , n15934 );
    and g21400 ( n9944 , n35273 , n29542 );
    xnor g21401 ( n32248 , n17622 , n32715 );
    or g21402 ( n8030 , n19550 , n11593 );
    or g21403 ( n19208 , n8170 , n32634 );
    xnor g21404 ( n29398 , n13197 , n15642 );
    or g21405 ( n491 , n22524 , n30674 );
    xnor g21406 ( n34494 , n27385 , n25456 );
    and g21407 ( n33109 , n3086 , n29627 );
    not g21408 ( n1187 , n3598 );
    or g21409 ( n15466 , n36038 , n14706 );
    xnor g21410 ( n8042 , n29395 , n15886 );
    xnor g21411 ( n20971 , n9893 , n28909 );
    or g21412 ( n13856 , n23035 , n32750 );
    or g21413 ( n22088 , n29044 , n18305 );
    or g21414 ( n34946 , n16634 , n1402 );
    xnor g21415 ( n19467 , n28545 , n23604 );
    xnor g21416 ( n16286 , n8470 , n19953 );
    not g21417 ( n20029 , n34094 );
    not g21418 ( n24586 , n16620 );
    xnor g21419 ( n34035 , n20378 , n24882 );
    and g21420 ( n19509 , n28785 , n3620 );
    xnor g21421 ( n1938 , n983 , n8432 );
    or g21422 ( n26572 , n33119 , n3680 );
    xnor g21423 ( n30626 , n13770 , n17376 );
    or g21424 ( n540 , n10894 , n27863 );
    not g21425 ( n19198 , n29431 );
    or g21426 ( n2297 , n35789 , n1511 );
    nor g21427 ( n12324 , n933 , n31411 );
    and g21428 ( n16542 , n11386 , n18355 );
    xnor g21429 ( n24879 , n24353 , n3148 );
    nor g21430 ( n29623 , n5287 , n29273 );
    and g21431 ( n9162 , n28362 , n35760 );
    xnor g21432 ( n10101 , n6828 , n11046 );
    and g21433 ( n27796 , n3932 , n29608 );
    nor g21434 ( n19410 , n30702 , n4104 );
    xnor g21435 ( n11336 , n3299 , n24433 );
    or g21436 ( n2779 , n21118 , n16762 );
    and g21437 ( n5355 , n24835 , n15424 );
    xnor g21438 ( n22157 , n4827 , n32857 );
    or g21439 ( n84 , n4001 , n11518 );
    nor g21440 ( n1380 , n11190 , n5477 );
    xnor g21441 ( n1028 , n13263 , n29267 );
    and g21442 ( n833 , n8102 , n3166 );
    or g21443 ( n30351 , n6377 , n28404 );
    xnor g21444 ( n30819 , n2402 , n22915 );
    or g21445 ( n35350 , n18868 , n16294 );
    xnor g21446 ( n13558 , n23636 , n2880 );
    and g21447 ( n15262 , n29621 , n4795 );
    and g21448 ( n24086 , n1291 , n28691 );
    xnor g21449 ( n14128 , n33645 , n24172 );
    xnor g21450 ( n32695 , n26072 , n26683 );
    nor g21451 ( n27894 , n20327 , n10556 );
    or g21452 ( n29763 , n12740 , n3414 );
    or g21453 ( n4392 , n31799 , n3327 );
    or g21454 ( n34582 , n16620 , n19347 );
    and g21455 ( n7872 , n32148 , n3112 );
    or g21456 ( n25492 , n16922 , n13652 );
    and g21457 ( n10475 , n29196 , n33259 );
    or g21458 ( n4313 , n25265 , n29953 );
    not g21459 ( n12254 , n16223 );
    not g21460 ( n16339 , n2562 );
    and g21461 ( n29172 , n12208 , n7968 );
    or g21462 ( n25528 , n3794 , n32963 );
    nor g21463 ( n20573 , n19510 , n1470 );
    and g21464 ( n5195 , n30958 , n26415 );
    xnor g21465 ( n16705 , n20755 , n9097 );
    or g21466 ( n6460 , n35797 , n32872 );
    or g21467 ( n23752 , n15474 , n18477 );
    or g21468 ( n3057 , n7842 , n27725 );
    or g21469 ( n30937 , n36026 , n5139 );
    xnor g21470 ( n18136 , n13168 , n26184 );
    and g21471 ( n4911 , n12995 , n25297 );
    xnor g21472 ( n23006 , n1837 , n27300 );
    or g21473 ( n34348 , n17568 , n14405 );
    xnor g21474 ( n16284 , n28372 , n23730 );
    and g21475 ( n25652 , n16593 , n9206 );
    and g21476 ( n21112 , n2742 , n12887 );
    and g21477 ( n28434 , n23381 , n32819 );
    and g21478 ( n16910 , n23061 , n12746 );
    or g21479 ( n10649 , n33455 , n25898 );
    and g21480 ( n29188 , n13692 , n3390 );
    nor g21481 ( n5384 , n19984 , n16703 );
    or g21482 ( n1506 , n10218 , n11071 );
    xnor g21483 ( n27084 , n35833 , n14545 );
    and g21484 ( n18588 , n34720 , n9329 );
    xnor g21485 ( n28347 , n652 , n16620 );
    xnor g21486 ( n35668 , n36013 , n2351 );
    and g21487 ( n12677 , n3925 , n32444 );
    or g21488 ( n21310 , n22479 , n25255 );
    nor g21489 ( n1932 , n15886 , n11359 );
    and g21490 ( n28822 , n13835 , n28725 );
    or g21491 ( n16295 , n3927 , n3518 );
    and g21492 ( n9576 , n21455 , n32163 );
    buf g21493 ( n12791 , n30519 );
    or g21494 ( n29933 , n23109 , n23677 );
    or g21495 ( n8949 , n35105 , n29036 );
    xnor g21496 ( n14468 , n16857 , n15991 );
    or g21497 ( n20614 , n22291 , n20960 );
    or g21498 ( n2874 , n9168 , n17601 );
    xnor g21499 ( n24241 , n16793 , n2888 );
    or g21500 ( n30666 , n35927 , n32442 );
    xnor g21501 ( n31830 , n23886 , n13966 );
    or g21502 ( n24242 , n3317 , n17852 );
    or g21503 ( n20369 , n28117 , n22783 );
    and g21504 ( n29080 , n23488 , n11340 );
    or g21505 ( n21141 , n10657 , n24672 );
    or g21506 ( n9011 , n16922 , n17575 );
    and g21507 ( n12649 , n12469 , n28731 );
    or g21508 ( n14695 , n17379 , n26365 );
    or g21509 ( n23732 , n31799 , n28712 );
    or g21510 ( n6901 , n30742 , n25982 );
    or g21511 ( n10305 , n30553 , n14106 );
    or g21512 ( n13766 , n32975 , n15344 );
    or g21513 ( n7433 , n2341 , n7788 );
    or g21514 ( n31738 , n25512 , n8283 );
    and g21515 ( n14978 , n6612 , n27455 );
    and g21516 ( n32092 , n22205 , n22365 );
    xnor g21517 ( n15359 , n12000 , n9009 );
    xnor g21518 ( n35606 , n18263 , n22751 );
    or g21519 ( n33818 , n26744 , n1763 );
    or g21520 ( n20243 , n19852 , n5186 );
    or g21521 ( n23088 , n24403 , n2823 );
    or g21522 ( n1163 , n11330 , n33036 );
    xnor g21523 ( n20202 , n12636 , n34556 );
    and g21524 ( n681 , n3869 , n13754 );
    or g21525 ( n13003 , n29097 , n14746 );
    and g21526 ( n21962 , n18330 , n12508 );
    xnor g21527 ( n5985 , n13971 , n34161 );
    or g21528 ( n4388 , n4960 , n17991 );
    or g21529 ( n30316 , n35209 , n14075 );
    not g21530 ( n439 , n11455 );
    and g21531 ( n18981 , n28233 , n14559 );
    or g21532 ( n8856 , n22066 , n15144 );
    not g21533 ( n18596 , n10195 );
    or g21534 ( n21172 , n9793 , n21981 );
    not g21535 ( n22681 , n25708 );
    nor g21536 ( n18705 , n10945 , n4065 );
    or g21537 ( n24366 , n15733 , n6683 );
    xnor g21538 ( n21323 , n33882 , n20341 );
    or g21539 ( n24078 , n32715 , n30953 );
    or g21540 ( n27357 , n15464 , n7170 );
    xnor g21541 ( n14259 , n4981 , n24741 );
    and g21542 ( n29715 , n30572 , n15710 );
    or g21543 ( n2391 , n4288 , n7564 );
    nor g21544 ( n17467 , n9793 , n3579 );
    or g21545 ( n32720 , n6927 , n24672 );
    buf g21546 ( n26737 , n11712 );
    or g21547 ( n16746 , n12117 , n34084 );
    not g21548 ( n22866 , n8431 );
    or g21549 ( n29263 , n672 , n6374 );
    and g21550 ( n3463 , n17530 , n13698 );
    or g21551 ( n20801 , n9789 , n20952 );
    not g21552 ( n33489 , n34739 );
    xnor g21553 ( n11738 , n26226 , n17978 );
    or g21554 ( n31574 , n10979 , n4637 );
    xnor g21555 ( n4286 , n19140 , n29634 );
    not g21556 ( n23714 , n16533 );
    or g21557 ( n34486 , n10450 , n19084 );
    xnor g21558 ( n8178 , n6440 , n27113 );
    xnor g21559 ( n21844 , n19959 , n12198 );
    or g21560 ( n30305 , n16970 , n2330 );
    and g21561 ( n16069 , n21972 , n16400 );
    or g21562 ( n233 , n20249 , n16133 );
    or g21563 ( n16590 , n29457 , n18264 );
    xnor g21564 ( n17471 , n31878 , n4040 );
    or g21565 ( n14378 , n13005 , n578 );
    xnor g21566 ( n35360 , n29864 , n23489 );
    xnor g21567 ( n25928 , n16403 , n15464 );
    or g21568 ( n4966 , n2992 , n9675 );
    or g21569 ( n31113 , n34246 , n35748 );
    not g21570 ( n17166 , n13438 );
    and g21571 ( n14507 , n9691 , n2627 );
    or g21572 ( n29394 , n11461 , n12021 );
    xnor g21573 ( n1496 , n17902 , n31559 );
    or g21574 ( n32998 , n1420 , n27728 );
    or g21575 ( n20396 , n3236 , n22206 );
    not g21576 ( n24431 , n16223 );
    not g21577 ( n628 , n28866 );
    or g21578 ( n16315 , n21188 , n8389 );
    xnor g21579 ( n21826 , n33164 , n32095 );
    and g21580 ( n3391 , n24912 , n12074 );
    and g21581 ( n23879 , n12297 , n31661 );
    xnor g21582 ( n24737 , n16616 , n9658 );
    xnor g21583 ( n16945 , n19271 , n31559 );
    or g21584 ( n13579 , n2718 , n25924 );
    or g21585 ( n33410 , n18516 , n2168 );
    or g21586 ( n11734 , n26493 , n28837 );
    xnor g21587 ( n72 , n6586 , n31559 );
    or g21588 ( n21879 , n19551 , n24450 );
    or g21589 ( n11342 , n16095 , n544 );
    and g21590 ( n1200 , n8036 , n20042 );
    or g21591 ( n22653 , n29713 , n31736 );
    xnor g21592 ( n6533 , n26208 , n4288 );
    or g21593 ( n11857 , n23155 , n25940 );
    and g21594 ( n16451 , n16830 , n35418 );
    and g21595 ( n33364 , n491 , n28590 );
    xnor g21596 ( n19988 , n22774 , n23604 );
    not g21597 ( n13058 , n714 );
    and g21598 ( n29352 , n28991 , n27073 );
    or g21599 ( n24773 , n35927 , n4757 );
    and g21600 ( n20039 , n6538 , n32722 );
    or g21601 ( n16352 , n25118 , n6153 );
    or g21602 ( n1211 , n20264 , n14984 );
    or g21603 ( n13233 , n4962 , n7363 );
    or g21604 ( n13218 , n11787 , n25392 );
    or g21605 ( n30990 , n17785 , n23626 );
    and g21606 ( n14039 , n16313 , n2426 );
    or g21607 ( n28492 , n32584 , n7346 );
    xnor g21608 ( n13929 , n8748 , n15886 );
    xnor g21609 ( n22289 , n7235 , n34973 );
    or g21610 ( n1206 , n9793 , n17052 );
    and g21611 ( n8358 , n4156 , n10599 );
    xnor g21612 ( n29856 , n4679 , n4878 );
    xnor g21613 ( n23176 , n9614 , n19166 );
    or g21614 ( n17448 , n36042 , n30370 );
    xnor g21615 ( n17215 , n24415 , n5200 );
    and g21616 ( n29208 , n12880 , n35496 );
    and g21617 ( n35051 , n20282 , n33798 );
    or g21618 ( n16500 , n18529 , n3962 );
    or g21619 ( n4060 , n19237 , n20840 );
    or g21620 ( n2734 , n31185 , n22485 );
    or g21621 ( n31237 , n4223 , n20909 );
    xnor g21622 ( n30545 , n13366 , n17877 );
    not g21623 ( n10065 , n28273 );
    xnor g21624 ( n15691 , n3957 , n10745 );
    xnor g21625 ( n6613 , n31436 , n11990 );
    or g21626 ( n4166 , n4284 , n31554 );
    or g21627 ( n16032 , n17265 , n949 );
    or g21628 ( n32591 , n18697 , n11850 );
    and g21629 ( n5530 , n25525 , n13248 );
    and g21630 ( n8905 , n23726 , n107 );
    xnor g21631 ( n4125 , n8093 , n574 );
    xnor g21632 ( n17609 , n34255 , n19798 );
    or g21633 ( n25654 , n8511 , n24679 );
    and g21634 ( n18248 , n13644 , n21385 );
    xnor g21635 ( n7984 , n7495 , n12402 );
    xnor g21636 ( n34824 , n1327 , n3222 );
    or g21637 ( n29580 , n4288 , n1627 );
    not g21638 ( n31065 , n31928 );
    or g21639 ( n4412 , n8609 , n19336 );
    or g21640 ( n16308 , n11070 , n19403 );
    or g21641 ( n15015 , n29617 , n26737 );
    and g21642 ( n34172 , n3991 , n9700 );
    or g21643 ( n27321 , n5262 , n5821 );
    xnor g21644 ( n235 , n28766 , n17018 );
    buf g21645 ( n16457 , n33469 );
    and g21646 ( n10107 , n26848 , n33651 );
    xnor g21647 ( n2665 , n18037 , n32715 );
    xnor g21648 ( n30735 , n2576 , n21349 );
    not g21649 ( n30893 , n20029 );
    or g21650 ( n2724 , n9038 , n3950 );
    or g21651 ( n10671 , n28143 , n11593 );
    or g21652 ( n13658 , n5690 , n25447 );
    and g21653 ( n3132 , n12941 , n7677 );
    or g21654 ( n8471 , n26778 , n33725 );
    nor g21655 ( n21800 , n18537 , n30444 );
    or g21656 ( n16256 , n5335 , n6503 );
    not g21657 ( n3158 , n5738 );
    and g21658 ( n10670 , n2720 , n19693 );
    xnor g21659 ( n15284 , n10318 , n32806 );
    or g21660 ( n21380 , n5335 , n20025 );
    or g21661 ( n25022 , n28635 , n18591 );
    or g21662 ( n22925 , n8748 , n14918 );
    and g21663 ( n3989 , n2390 , n21482 );
    or g21664 ( n33375 , n3353 , n2117 );
    xnor g21665 ( n30215 , n24063 , n6531 );
    or g21666 ( n19681 , n5613 , n13900 );
    not g21667 ( n5339 , n33272 );
    and g21668 ( n20909 , n30414 , n6455 );
    xnor g21669 ( n18049 , n26335 , n23755 );
    or g21670 ( n23082 , n32584 , n2136 );
    xnor g21671 ( n34023 , n16249 , n28852 );
    xnor g21672 ( n23151 , n24589 , n5287 );
    or g21673 ( n6734 , n18734 , n8648 );
    or g21674 ( n27566 , n5998 , n34110 );
    or g21675 ( n10384 , n33146 , n18542 );
    or g21676 ( n6265 , n5961 , n14706 );
    and g21677 ( n24745 , n17113 , n28492 );
    and g21678 ( n23914 , n13228 , n3878 );
    and g21679 ( n24104 , n25692 , n2028 );
    and g21680 ( n12046 , n3408 , n28487 );
    nor g21681 ( n23836 , n11969 , n1595 );
    xnor g21682 ( n35447 , n27046 , n3222 );
    xnor g21683 ( n10048 , n16205 , n2668 );
    and g21684 ( n14472 , n12697 , n11645 );
    or g21685 ( n328 , n29226 , n28836 );
    and g21686 ( n6790 , n33688 , n26114 );
    or g21687 ( n4228 , n17844 , n27973 );
    or g21688 ( n22431 , n25174 , n34731 );
    xnor g21689 ( n4079 , n12019 , n9127 );
    or g21690 ( n27492 , n18379 , n24514 );
    or g21691 ( n5153 , n7461 , n30617 );
    and g21692 ( n9401 , n7165 , n21483 );
    or g21693 ( n18731 , n5065 , n8149 );
    or g21694 ( n17908 , n668 , n25447 );
    or g21695 ( n13412 , n28844 , n17876 );
    and g21696 ( n5242 , n20799 , n25028 );
    or g21697 ( n6354 , n19074 , n544 );
    and g21698 ( n34103 , n24099 , n11550 );
    not g21699 ( n21134 , n1825 );
    xnor g21700 ( n24677 , n31598 , n20094 );
    and g21701 ( n8122 , n31539 , n32656 );
    and g21702 ( n24793 , n18565 , n15903 );
    or g21703 ( n21222 , n17568 , n15005 );
    or g21704 ( n19685 , n16911 , n29465 );
    or g21705 ( n3632 , n14720 , n139 );
    or g21706 ( n9806 , n4640 , n12128 );
    and g21707 ( n24317 , n18517 , n2671 );
    nor g21708 ( n2946 , n17594 , n29092 );
    nor g21709 ( n21742 , n34432 , n4508 );
    not g21710 ( n13193 , n7588 );
    or g21711 ( n6889 , n9658 , n15267 );
    or g21712 ( n6952 , n11456 , n10432 );
    and g21713 ( n7259 , n16662 , n2882 );
    and g21714 ( n27734 , n1301 , n25685 );
    and g21715 ( n33317 , n1667 , n33548 );
    nor g21716 ( n911 , n31799 , n13578 );
    and g21717 ( n25596 , n25112 , n7761 );
    not g21718 ( n8242 , n22980 );
    or g21719 ( n13136 , n996 , n23122 );
    or g21720 ( n15533 , n32472 , n139 );
    or g21721 ( n25252 , n2975 , n23368 );
    and g21722 ( n32778 , n30015 , n16844 );
    or g21723 ( n12158 , n11509 , n25831 );
    or g21724 ( n11021 , n27537 , n19005 );
    and g21725 ( n26108 , n15176 , n29191 );
    or g21726 ( n18617 , n32715 , n20402 );
    and g21727 ( n27688 , n33386 , n32899 );
    xnor g21728 ( n16799 , n30724 , n17131 );
    or g21729 ( n195 , n17568 , n6675 );
    xnor g21730 ( n17061 , n22373 , n14414 );
    xnor g21731 ( n6732 , n23770 , n5807 );
    and g21732 ( n13162 , n20355 , n992 );
    or g21733 ( n10806 , n29391 , n24333 );
    xnor g21734 ( n27235 , n14239 , n12826 );
    and g21735 ( n12135 , n12280 , n26668 );
    and g21736 ( n4308 , n33938 , n19698 );
    or g21737 ( n32000 , n18669 , n1198 );
    or g21738 ( n26352 , n31692 , n29411 );
    or g21739 ( n19623 , n33269 , n13664 );
    or g21740 ( n18673 , n25119 , n25592 );
    nor g21741 ( n23374 , n25174 , n33093 );
    or g21742 ( n30014 , n28917 , n4788 );
    or g21743 ( n22392 , n15079 , n10140 );
    nor g21744 ( n7899 , n16610 , n6333 );
    xnor g21745 ( n3792 , n31651 , n29296 );
    xnor g21746 ( n3594 , n21337 , n28124 );
    or g21747 ( n6496 , n8803 , n585 );
    xnor g21748 ( n2532 , n33109 , n10894 );
    and g21749 ( n16054 , n1539 , n116 );
    or g21750 ( n29770 , n24243 , n14706 );
    and g21751 ( n20911 , n34504 , n30106 );
    or g21752 ( n32007 , n3205 , n668 );
    or g21753 ( n14564 , n5852 , n21177 );
    or g21754 ( n21842 , n35441 , n20049 );
    not g21755 ( n11261 , n30204 );
    or g21756 ( n21683 , n10201 , n20840 );
    xnor g21757 ( n35482 , n6495 , n12124 );
    xnor g21758 ( n25097 , n27288 , n23604 );
    not g21759 ( n17898 , n17568 );
    xnor g21760 ( n19324 , n26126 , n35927 );
    nor g21761 ( n31455 , n11485 , n18964 );
    xnor g21762 ( n22167 , n7005 , n21819 );
    buf g21763 ( n19105 , n19939 );
    or g21764 ( n11421 , n11294 , n23870 );
    or g21765 ( n14478 , n5919 , n3805 );
    and g21766 ( n4621 , n16701 , n1937 );
    and g21767 ( n18266 , n12783 , n11769 );
    not g21768 ( n32059 , n30292 );
    or g21769 ( n4678 , n18182 , n33486 );
    or g21770 ( n5974 , n26410 , n2823 );
    xnor g21771 ( n201 , n20392 , n20917 );
    and g21772 ( n18305 , n30453 , n34355 );
    or g21773 ( n12147 , n103 , n3738 );
    or g21774 ( n29471 , n19551 , n35791 );
    or g21775 ( n18653 , n26270 , n9555 );
    nor g21776 ( n14244 , n15886 , n23196 );
    and g21777 ( n24548 , n20814 , n19117 );
    or g21778 ( n24984 , n8804 , n22322 );
    and g21779 ( n25984 , n18480 , n7783 );
    not g21780 ( n5662 , n19982 );
    or g21781 ( n2862 , n5287 , n10553 );
    or g21782 ( n1696 , n17568 , n3136 );
    or g21783 ( n20988 , n9793 , n1197 );
    or g21784 ( n14406 , n23723 , n14778 );
    and g21785 ( n26719 , n4238 , n16416 );
    and g21786 ( n28456 , n22374 , n1068 );
    and g21787 ( n14988 , n32598 , n3427 );
    xnor g21788 ( n13726 , n21391 , n11459 );
    and g21789 ( n12540 , n19176 , n14715 );
    or g21790 ( n1580 , n19714 , n10348 );
    xnor g21791 ( n34666 , n32348 , n4878 );
    or g21792 ( n25591 , n35649 , n20318 );
    xnor g21793 ( n8651 , n13186 , n17568 );
    or g21794 ( n29861 , n9752 , n28404 );
    not g21795 ( n33723 , n12650 );
    and g21796 ( n10967 , n25585 , n18788 );
    xnor g21797 ( n22962 , n27690 , n29839 );
    and g21798 ( n18052 , n2888 , n16793 );
    or g21799 ( n6574 , n35927 , n35259 );
    or g21800 ( n17279 , n1624 , n10122 );
    or g21801 ( n32773 , n23654 , n1042 );
    xnor g21802 ( n23265 , n35614 , n28357 );
    or g21803 ( n33412 , n30742 , n16763 );
    or g21804 ( n8262 , n28579 , n21837 );
    or g21805 ( n13237 , n4962 , n12532 );
    and g21806 ( n9403 , n32256 , n1 );
    xnor g21807 ( n880 , n21638 , n8432 );
    or g21808 ( n6292 , n27015 , n4821 );
    xnor g21809 ( n19026 , n18667 , n4288 );
    or g21810 ( n4278 , n17433 , n29323 );
    xnor g21811 ( n30226 , n13929 , n12453 );
    nor g21812 ( n14906 , n20239 , n33956 );
    xnor g21813 ( n7466 , n35830 , n26503 );
    or g21814 ( n22012 , n19551 , n13300 );
    or g21815 ( n35890 , n19376 , n9915 );
    xnor g21816 ( n24044 , n18235 , n35927 );
    or g21817 ( n32084 , n11190 , n8437 );
    or g21818 ( n27012 , n25239 , n11812 );
    or g21819 ( n17977 , n28350 , n5779 );
    xnor g21820 ( n23640 , n31513 , n27421 );
    xnor g21821 ( n28596 , n13769 , n15886 );
    xnor g21822 ( n3324 , n19162 , n9872 );
    not g21823 ( n33384 , n28781 );
    or g21824 ( n34651 , n14678 , n17226 );
    or g21825 ( n23117 , n5118 , n35935 );
    and g21826 ( n12944 , n4942 , n6520 );
    and g21827 ( n34702 , n33881 , n14054 );
    or g21828 ( n20510 , n9724 , n23921 );
    not g21829 ( n18913 , n22980 );
    not g21830 ( n21113 , n12681 );
    or g21831 ( n20282 , n7133 , n2174 );
    nor g21832 ( n464 , n27226 , n15361 );
    or g21833 ( n15865 , n11046 , n17356 );
    and g21834 ( n3106 , n31159 , n2123 );
    or g21835 ( n883 , n235 , n28668 );
    and g21836 ( n28594 , n20557 , n16758 );
    and g21837 ( n22052 , n10643 , n32357 );
    or g21838 ( n23657 , n28444 , n15581 );
    xnor g21839 ( n25144 , n3637 , n3205 );
    or g21840 ( n25101 , n19461 , n14716 );
    buf g21841 ( n10432 , n27404 );
    xnor g21842 ( n3073 , n24315 , n15872 );
    or g21843 ( n26918 , n15607 , n24793 );
    and g21844 ( n4258 , n17636 , n15551 );
    or g21845 ( n31537 , n31619 , n15290 );
    xnor g21846 ( n30542 , n1268 , n16519 );
    and g21847 ( n23259 , n30647 , n26240 );
    or g21848 ( n25352 , n4878 , n34994 );
    and g21849 ( n4700 , n11701 , n8457 );
    and g21850 ( n10616 , n30088 , n13373 );
    nor g21851 ( n305 , n15403 , n24967 );
    or g21852 ( n20608 , n30545 , n12596 );
    or g21853 ( n25864 , n13158 , n20797 );
    xnor g21854 ( n1376 , n25047 , n20407 );
    and g21855 ( n3396 , n1769 , n12328 );
    not g21856 ( n14931 , n32857 );
    xnor g21857 ( n28609 , n16971 , n7339 );
    or g21858 ( n8367 , n6586 , n33310 );
    xnor g21859 ( n26502 , n8100 , n4288 );
    xnor g21860 ( n21769 , n13127 , n33630 );
    xnor g21861 ( n29701 , n10145 , n11455 );
    not g21862 ( n8855 , n9789 );
    or g21863 ( n24284 , n16922 , n13456 );
    nor g21864 ( n31094 , n561 , n7096 );
    xnor g21865 ( n34134 , n24900 , n30742 );
    or g21866 ( n20570 , n4288 , n6684 );
    and g21867 ( n24837 , n25656 , n32521 );
    nor g21868 ( n5437 , n24371 , n26561 );
    and g21869 ( n33335 , n34841 , n34338 );
    or g21870 ( n12008 , n25602 , n4405 );
    or g21871 ( n27406 , n5335 , n5580 );
    and g21872 ( n26512 , n6728 , n21623 );
    or g21873 ( n10304 , n7621 , n6683 );
    xnor g21874 ( n21852 , n7262 , n11455 );
    xnor g21875 ( n30391 , n21098 , n9540 );
    or g21876 ( n26976 , n24545 , n10336 );
    or g21877 ( n8693 , n20870 , n28507 );
    and g21878 ( n31531 , n32292 , n23683 );
    or g21879 ( n21001 , n17788 , n35111 );
    or g21880 ( n19817 , n13375 , n31053 );
    nor g21881 ( n23601 , n28966 , n14137 );
    or g21882 ( n14238 , n27291 , n28551 );
    or g21883 ( n29726 , n31289 , n4830 );
    nor g21884 ( n31321 , n17484 , n32005 );
    not g21885 ( n8781 , n35927 );
    not g21886 ( n20152 , n2676 );
    or g21887 ( n35488 , n3205 , n16177 );
    xnor g21888 ( n3677 , n16522 , n16729 );
    and g21889 ( n15829 , n33495 , n31045 );
    or g21890 ( n2162 , n29839 , n1634 );
    and g21891 ( n21463 , n19003 , n15764 );
    or g21892 ( n14768 , n22291 , n7546 );
    and g21893 ( n12844 , n4798 , n7821 );
    xnor g21894 ( n12517 , n1009 , n6490 );
    or g21895 ( n33678 , n30805 , n10363 );
    xnor g21896 ( n10218 , n26966 , n27226 );
    or g21897 ( n30551 , n32158 , n17862 );
    or g21898 ( n14348 , n21666 , n29866 );
    or g21899 ( n12856 , n18192 , n34971 );
    xnor g21900 ( n30102 , n7170 , n15464 );
    or g21901 ( n22403 , n448 , n29626 );
    or g21902 ( n6564 , n10894 , n31746 );
    and g21903 ( n20621 , n35234 , n20532 );
    or g21904 ( n31730 , n10214 , n3483 );
    not g21905 ( n14056 , n32095 );
    or g21906 ( n35070 , n7540 , n11188 );
    and g21907 ( n4603 , n2199 , n26409 );
    not g21908 ( n3490 , n7352 );
    or g21909 ( n32193 , n9793 , n18891 );
    and g21910 ( n16806 , n18176 , n14769 );
    or g21911 ( n23367 , n26180 , n18811 );
    xnor g21912 ( n5085 , n7907 , n1950 );
    or g21913 ( n14724 , n25326 , n5167 );
    or g21914 ( n31712 , n35586 , n1100 );
    xnor g21915 ( n29206 , n19679 , n32105 );
    or g21916 ( n10117 , n7963 , n9921 );
    and g21917 ( n19555 , n8653 , n23343 );
    or g21918 ( n3682 , n24371 , n647 );
    xnor g21919 ( n31801 , n22518 , n32721 );
    or g21920 ( n29247 , n25277 , n10289 );
    xnor g21921 ( n20708 , n8435 , n7540 );
    or g21922 ( n1908 , n35927 , n32290 );
    and g21923 ( n14099 , n9305 , n14669 );
    xnor g21924 ( n12527 , n35204 , n31273 );
    and g21925 ( n10485 , n19610 , n25634 );
    and g21926 ( n24546 , n24199 , n23631 );
    xnor g21927 ( n19009 , n2225 , n21266 );
    or g21928 ( n3843 , n8814 , n24628 );
    or g21929 ( n105 , n16922 , n5402 );
    or g21930 ( n10574 , n7930 , n3338 );
    or g21931 ( n24239 , n13344 , n33000 );
    or g21932 ( n20142 , n16620 , n5883 );
    xnor g21933 ( n19236 , n4233 , n23604 );
    or g21934 ( n13257 , n12767 , n27462 );
    or g21935 ( n33560 , n14029 , n31773 );
    or g21936 ( n26635 , n26833 , n25831 );
    nor g21937 ( n35007 , n16922 , n14571 );
    xnor g21938 ( n1261 , n18374 , n20079 );
    or g21939 ( n25412 , n15201 , n22732 );
    xnor g21940 ( n24343 , n4923 , n16757 );
    xnor g21941 ( n163 , n4026 , n27291 );
    xnor g21942 ( n12003 , n24603 , n10277 );
    and g21943 ( n23315 , n29412 , n11581 );
    xnor g21944 ( n5033 , n30713 , n28336 );
    nor g21945 ( n17895 , n14116 , n20915 );
    not g21946 ( n2860 , n31799 );
    or g21947 ( n23619 , n16207 , n30646 );
    and g21948 ( n2295 , n33290 , n1006 );
    and g21949 ( n9037 , n445 , n34619 );
    or g21950 ( n12497 , n11085 , n13217 );
    nor g21951 ( n15947 , n35927 , n23483 );
    nor g21952 ( n35115 , n25767 , n30950 );
    or g21953 ( n18627 , n31467 , n13305 );
    nor g21954 ( n8346 , n4878 , n28500 );
    or g21955 ( n31323 , n19551 , n13925 );
    or g21956 ( n31135 , n14187 , n17964 );
    or g21957 ( n22064 , n23662 , n26555 );
    nor g21958 ( n30620 , n21413 , n19190 );
    or g21959 ( n10274 , n24349 , n12332 );
    nor g21960 ( n27246 , n10586 , n25594 );
    or g21961 ( n16977 , n32857 , n8834 );
    and g21962 ( n24968 , n23774 , n24244 );
    and g21963 ( n928 , n11393 , n32903 );
    or g21964 ( n18155 , n2274 , n26220 );
    or g21965 ( n12368 , n17332 , n26866 );
    or g21966 ( n1208 , n17820 , n35630 );
    xnor g21967 ( n9383 , n21213 , n20197 );
    and g21968 ( n13028 , n7859 , n28727 );
    xnor g21969 ( n26571 , n5625 , n18393 );
    xnor g21970 ( n19536 , n9126 , n1274 );
    xnor g21971 ( n25584 , n15209 , n35927 );
    xnor g21972 ( n28412 , n4879 , n9342 );
    not g21973 ( n10490 , n7588 );
    or g21974 ( n5237 , n10553 , n2814 );
    and g21975 ( n24294 , n17645 , n25851 );
    or g21976 ( n24019 , n3324 , n12622 );
    or g21977 ( n23215 , n8168 , n34727 );
    or g21978 ( n2595 , n31289 , n12358 );
    or g21979 ( n18793 , n6680 , n3858 );
    not g21980 ( n28031 , n34095 );
    xnor g21981 ( n14968 , n4884 , n25953 );
    xnor g21982 ( n7325 , n17839 , n830 );
    or g21983 ( n9374 , n29194 , n13900 );
    and g21984 ( n31596 , n5652 , n1141 );
    xnor g21985 ( n7408 , n17436 , n32857 );
    or g21986 ( n10258 , n3205 , n35865 );
    or g21987 ( n4034 , n2369 , n9030 );
    and g21988 ( n1934 , n2645 , n34099 );
    xnor g21989 ( n12874 , n13671 , n30864 );
    not g21990 ( n8025 , n19510 );
    buf g21991 ( n19490 , n9210 );
    or g21992 ( n2537 , n2505 , n29454 );
    not g21993 ( n17782 , n16223 );
    or g21994 ( n231 , n24371 , n13731 );
    and g21995 ( n12433 , n11972 , n9934 );
    or g21996 ( n15936 , n8469 , n288 );
    xnor g21997 ( n15699 , n1436 , n11046 );
    nor g21998 ( n24569 , n10894 , n25476 );
    or g21999 ( n6904 , n9838 , n24710 );
    nor g22000 ( n2410 , n31690 , n25197 );
    and g22001 ( n11921 , n26141 , n9296 );
    xnor g22002 ( n17293 , n13479 , n32874 );
    and g22003 ( n34635 , n33607 , n12475 );
    nor g22004 ( n5876 , n9793 , n31417 );
    or g22005 ( n21692 , n5372 , n27801 );
    nor g22006 ( n2811 , n17568 , n15975 );
    or g22007 ( n21309 , n5782 , n12030 );
    and g22008 ( n25234 , n1279 , n22617 );
    xnor g22009 ( n1787 , n31124 , n3205 );
    xnor g22010 ( n6148 , n8056 , n3946 );
    or g22011 ( n23671 , n25400 , n17447 );
    xnor g22012 ( n6231 , n36046 , n4878 );
    or g22013 ( n21563 , n23464 , n5972 );
    or g22014 ( n28504 , n15698 , n17932 );
    nor g22015 ( n3668 , n30396 , n4508 );
    or g22016 ( n15671 , n31200 , n25334 );
    xnor g22017 ( n18827 , n8829 , n8796 );
    or g22018 ( n4798 , n34066 , n19336 );
    and g22019 ( n2735 , n32591 , n24780 );
    or g22020 ( n8321 , n29342 , n29643 );
    or g22021 ( n9169 , n4373 , n25940 );
    or g22022 ( n35379 , n14115 , n35478 );
    or g22023 ( n10442 , n31149 , n7293 );
    nor g22024 ( n15607 , n22291 , n30682 );
    xnor g22025 ( n9900 , n32816 , n4962 );
    not g22026 ( n1957 , n26918 );
    xnor g22027 ( n20146 , n8621 , n30683 );
    buf g22028 ( n4772 , n3560 );
    or g22029 ( n30201 , n14873 , n22946 );
    nor g22030 ( n25003 , n2902 , n32379 );
    or g22031 ( n8421 , n26725 , n36057 );
    and g22032 ( n188 , n28077 , n1032 );
    and g22033 ( n22989 , n26898 , n2246 );
    or g22034 ( n2194 , n31893 , n25398 );
    or g22035 ( n30426 , n5437 , n27004 );
    or g22036 ( n17276 , n29304 , n34433 );
    and g22037 ( n4830 , n20479 , n7818 );
    or g22038 ( n10756 , n35786 , n24356 );
    and g22039 ( n32322 , n2810 , n26952 );
    buf g22040 ( n20308 , n22870 );
    and g22041 ( n682 , n26361 , n21489 );
    or g22042 ( n20062 , n27215 , n18080 );
    and g22043 ( n4673 , n5176 , n14781 );
    and g22044 ( n32382 , n30524 , n35785 );
    nor g22045 ( n23681 , n3205 , n29748 );
    not g22046 ( n35963 , n17568 );
    and g22047 ( n25346 , n15237 , n21314 );
    and g22048 ( n7965 , n27495 , n31530 );
    nor g22049 ( n9597 , n32857 , n28292 );
    xnor g22050 ( n21544 , n10027 , n15464 );
    or g22051 ( n7450 , n19551 , n33015 );
    or g22052 ( n8631 , n1267 , n8755 );
    or g22053 ( n7786 , n16776 , n5771 );
    or g22054 ( n15091 , n7634 , n23809 );
    or g22055 ( n25309 , n11419 , n6340 );
    or g22056 ( n26198 , n25174 , n35847 );
    xnor g22057 ( n15624 , n6055 , n742 );
    or g22058 ( n24475 , n5162 , n31401 );
    nor g22059 ( n17864 , n3222 , n23183 );
    or g22060 ( n15417 , n20389 , n12950 );
    or g22061 ( n14514 , n182 , n29066 );
    or g22062 ( n27738 , n10852 , n24011 );
    not g22063 ( n31581 , n4960 );
    or g22064 ( n1547 , n12278 , n5607 );
    xnor g22065 ( n11724 , n35534 , n22641 );
    or g22066 ( n26124 , n12843 , n10535 );
    xnor g22067 ( n25338 , n28947 , n35310 );
    xnor g22068 ( n13799 , n33167 , n1950 );
    xnor g22069 ( n21196 , n882 , n30689 );
    xnor g22070 ( n10163 , n14837 , n4962 );
    xnor g22071 ( n13469 , n25687 , n5626 );
    or g22072 ( n22631 , n4045 , n2955 );
    and g22073 ( n18171 , n4872 , n18060 );
    or g22074 ( n26186 , n17121 , n26627 );
    not g22075 ( n10122 , n30193 );
    nor g22076 ( n2218 , n34992 , n18115 );
    and g22077 ( n27102 , n5104 , n32712 );
    or g22078 ( n20938 , n2192 , n24130 );
    nor g22079 ( n2739 , n27606 , n22124 );
    buf g22080 ( n22316 , n17313 );
    or g22081 ( n2920 , n24327 , n18059 );
    nor g22082 ( n5909 , n29607 , n22036 );
    not g22083 ( n17305 , n3498 );
    xnor g22084 ( n18160 , n4180 , n35927 );
    and g22085 ( n6725 , n22607 , n33566 );
    or g22086 ( n27083 , n24363 , n10336 );
    xnor g22087 ( n15960 , n2325 , n5114 );
    or g22088 ( n7421 , n21565 , n26953 );
    and g22089 ( n11509 , n19626 , n21229 );
    nor g22090 ( n17325 , n25602 , n5949 );
    xnor g22091 ( n30576 , n2656 , n34088 );
    or g22092 ( n33721 , n24777 , n31773 );
    or g22093 ( n3400 , n4913 , n3430 );
    xnor g22094 ( n15526 , n28551 , n27291 );
    xnor g22095 ( n30493 , n16512 , n15704 );
    buf g22096 ( n10417 , n15350 );
    and g22097 ( n9983 , n18730 , n15449 );
    nor g22098 ( n9563 , n34771 , n34711 );
    or g22099 ( n6953 , n10923 , n23446 );
    or g22100 ( n6273 , n11190 , n10873 );
    or g22101 ( n34992 , n35189 , n3341 );
    or g22102 ( n10189 , n22570 , n21673 );
    xnor g22103 ( n14941 , n13036 , n32715 );
    nor g22104 ( n31998 , n10017 , n5699 );
    or g22105 ( n17316 , n11820 , n23611 );
    or g22106 ( n19665 , n13941 , n14570 );
    and g22107 ( n33585 , n34942 , n33182 );
    or g22108 ( n11642 , n18861 , n19631 );
    xnor g22109 ( n23922 , n16738 , n11046 );
    and g22110 ( n2361 , n9973 , n28468 );
    or g22111 ( n15816 , n12354 , n13215 );
    and g22112 ( n33544 , n45 , n20422 );
    or g22113 ( n8526 , n31556 , n27476 );
    or g22114 ( n26075 , n12364 , n34826 );
    or g22115 ( n6766 , n32095 , n20832 );
    xnor g22116 ( n35346 , n30710 , n34001 );
    or g22117 ( n21265 , n6829 , n8392 );
    or g22118 ( n35103 , n13244 , n34472 );
    or g22119 ( n20160 , n18158 , n2384 );
    or g22120 ( n5415 , n14276 , n29656 );
    or g22121 ( n9906 , n9387 , n30646 );
    xnor g22122 ( n30105 , n8988 , n29839 );
    or g22123 ( n4294 , n12549 , n19939 );
    or g22124 ( n5603 , n12443 , n2927 );
    or g22125 ( n3564 , n23914 , n22858 );
    and g22126 ( n18700 , n31518 , n33337 );
    and g22127 ( n33751 , n2177 , n15300 );
    or g22128 ( n29115 , n4073 , n3502 );
    and g22129 ( n22035 , n12980 , n4854 );
    nor g22130 ( n959 , n30020 , n34022 );
    xnor g22131 ( n19126 , n13858 , n3964 );
    not g22132 ( n29216 , n32463 );
    or g22133 ( n8957 , n23025 , n34600 );
    and g22134 ( n15499 , n22486 , n3926 );
    or g22135 ( n19427 , n3368 , n3694 );
    or g22136 ( n24821 , n31559 , n7847 );
    xnor g22137 ( n18513 , n23183 , n3222 );
    xnor g22138 ( n26692 , n21132 , n859 );
    or g22139 ( n9700 , n30819 , n3634 );
    xnor g22140 ( n29149 , n22358 , n30454 );
    or g22141 ( n27069 , n3860 , n27893 );
    xnor g22142 ( n3126 , n14945 , n301 );
    and g22143 ( n8750 , n25408 , n30157 );
    and g22144 ( n2580 , n29541 , n14172 );
    or g22145 ( n15523 , n21083 , n32178 );
    xnor g22146 ( n10146 , n23758 , n33005 );
    or g22147 ( n31097 , n19669 , n19490 );
    or g22148 ( n4501 , n24949 , n19519 );
    or g22149 ( n2428 , n29255 , n14841 );
    or g22150 ( n1876 , n31289 , n5045 );
    or g22151 ( n26972 , n24296 , n33741 );
    xnor g22152 ( n7973 , n22070 , n7540 );
    or g22153 ( n24504 , n19551 , n8624 );
    xnor g22154 ( n16420 , n17736 , n29713 );
    or g22155 ( n5364 , n35436 , n27152 );
    xnor g22156 ( n13139 , n6503 , n5335 );
    not g22157 ( n5730 , n4407 );
    and g22158 ( n34898 , n33033 , n29728 );
    or g22159 ( n27229 , n18675 , n13480 );
    or g22160 ( n33955 , n9251 , n8375 );
    or g22161 ( n20655 , n10134 , n26931 );
    and g22162 ( n11841 , n1064 , n19966 );
    not g22163 ( n4653 , n33571 );
    or g22164 ( n15792 , n29116 , n4081 );
    xnor g22165 ( n5954 , n18551 , n7423 );
    and g22166 ( n35580 , n9806 , n6149 );
    or g22167 ( n2031 , n32400 , n5709 );
    xnor g22168 ( n14231 , n31675 , n25602 );
    or g22169 ( n5349 , n12105 , n4446 );
    and g22170 ( n26752 , n4219 , n11376 );
    or g22171 ( n5645 , n16021 , n9096 );
    nor g22172 ( n28747 , n35927 , n30677 );
    xnor g22173 ( n6851 , n16857 , n20239 );
    and g22174 ( n6151 , n5302 , n23772 );
    or g22175 ( n5193 , n3841 , n25263 );
    xnor g22176 ( n19956 , n25893 , n2984 );
    xnor g22177 ( n20597 , n6196 , n31188 );
    or g22178 ( n24804 , n22324 , n17640 );
    and g22179 ( n18406 , n1255 , n251 );
    and g22180 ( n20132 , n28815 , n11311 );
    xnor g22181 ( n20269 , n18920 , n26225 );
    and g22182 ( n29102 , n15338 , n11721 );
    or g22183 ( n2723 , n7906 , n29366 );
    and g22184 ( n27037 , n8408 , n17207 );
    not g22185 ( n25185 , n29203 );
    or g22186 ( n8923 , n7873 , n12664 );
    or g22187 ( n23513 , n4301 , n13900 );
    nor g22188 ( n14985 , n17687 , n3437 );
    xnor g22189 ( n31414 , n6474 , n9658 );
    or g22190 ( n1798 , n26573 , n21579 );
    not g22191 ( n20013 , n31574 );
    not g22192 ( n14024 , n19551 );
    xnor g22193 ( n26353 , n10449 , n17169 );
    or g22194 ( n28109 , n13567 , n30292 );
    xnor g22195 ( n5736 , n4250 , n28613 );
    and g22196 ( n30591 , n33992 , n25879 );
    and g22197 ( n15537 , n1912 , n14368 );
    or g22198 ( n27597 , n4878 , n18661 );
    or g22199 ( n15847 , n23552 , n26002 );
    or g22200 ( n8917 , n35262 , n25306 );
    and g22201 ( n10331 , n4347 , n28037 );
    and g22202 ( n11851 , n7225 , n438 );
    or g22203 ( n16790 , n20708 , n13810 );
    not g22204 ( n9984 , n5664 );
    or g22205 ( n33193 , n16530 , n31464 );
    not g22206 ( n25086 , n9658 );
    or g22207 ( n11311 , n9534 , n30646 );
    or g22208 ( n33599 , n17071 , n34423 );
    or g22209 ( n17160 , n16448 , n24505 );
    or g22210 ( n30074 , n31898 , n27756 );
    xnor g22211 ( n29164 , n28767 , n15490 );
    or g22212 ( n11184 , n30861 , n2829 );
    or g22213 ( n14207 , n14497 , n7448 );
    and g22214 ( n27089 , n4528 , n1765 );
    nor g22215 ( n22535 , n25233 , n4508 );
    and g22216 ( n29117 , n7415 , n33851 );
    xnor g22217 ( n5839 , n16048 , n8432 );
    or g22218 ( n31664 , n30852 , n30204 );
    not g22219 ( n23377 , n30732 );
    and g22220 ( n30468 , n2989 , n27301 );
    not g22221 ( n2299 , n3239 );
    xnor g22222 ( n1519 , n17524 , n15886 );
    or g22223 ( n14349 , n24496 , n34862 );
    not g22224 ( n26067 , n7605 );
    or g22225 ( n28570 , n18796 , n20958 );
    or g22226 ( n10473 , n3946 , n32217 );
    xnor g22227 ( n28358 , n14448 , n15886 );
    or g22228 ( n27999 , n25536 , n7844 );
    and g22229 ( n33960 , n13934 , n20218 );
    or g22230 ( n32471 , n22391 , n5972 );
    or g22231 ( n3119 , n24246 , n19105 );
    and g22232 ( n33413 , n29041 , n35761 );
    and g22233 ( n18510 , n31714 , n15149 );
    or g22234 ( n25853 , n4878 , n23900 );
    and g22235 ( n18689 , n29861 , n32439 );
    and g22236 ( n19413 , n20496 , n9650 );
    and g22237 ( n31140 , n6501 , n32595 );
    not g22238 ( n24053 , n9658 );
    xnor g22239 ( n9510 , n21232 , n5335 );
    xnor g22240 ( n11822 , n11246 , n29205 );
    or g22241 ( n15629 , n19697 , n6950 );
    and g22242 ( n21707 , n29568 , n15927 );
    or g22243 ( n6235 , n25602 , n18633 );
    xnor g22244 ( n18410 , n14071 , n10275 );
    nor g22245 ( n21239 , n34813 , n26095 );
    nor g22246 ( n808 , n14639 , n4108 );
    nor g22247 ( n22874 , n25503 , n9225 );
    not g22248 ( n8966 , n24265 );
    xnor g22249 ( n25460 , n4976 , n29839 );
    and g22250 ( n9238 , n26997 , n11356 );
    and g22251 ( n20776 , n7412 , n6044 );
    and g22252 ( n17037 , n34919 , n12728 );
    or g22253 ( n2358 , n15705 , n34735 );
    and g22254 ( n15086 , n9954 , n22825 );
    or g22255 ( n27883 , n2910 , n27641 );
    nor g22256 ( n26696 , n3020 , n21714 );
    or g22257 ( n5545 , n15403 , n863 );
    or g22258 ( n34948 , n15875 , n24259 );
    xnor g22259 ( n18674 , n28779 , n31704 );
    or g22260 ( n10686 , n23306 , n22241 );
    nor g22261 ( n5591 , n18233 , n27214 );
    and g22262 ( n10052 , n18048 , n21571 );
    xnor g22263 ( n24106 , n255 , n25086 );
    or g22264 ( n28674 , n10894 , n23602 );
    or g22265 ( n32506 , n2240 , n11755 );
    and g22266 ( n7915 , n21939 , n30122 );
    xnor g22267 ( n34511 , n7346 , n32584 );
    or g22268 ( n33168 , n2895 , n429 );
    nor g22269 ( n29341 , n2022 , n36030 );
    xnor g22270 ( n1037 , n12955 , n36005 );
    or g22271 ( n32124 , n28123 , n597 );
    and g22272 ( n35907 , n14581 , n12322 );
    or g22273 ( n5537 , n1650 , n23130 );
    xnor g22274 ( n11249 , n342 , n8237 );
    not g22275 ( n3570 , n16075 );
    nor g22276 ( n10971 , n31056 , n20067 );
    xnor g22277 ( n19049 , n19589 , n4878 );
    or g22278 ( n26196 , n9080 , n10128 );
    or g22279 ( n2094 , n19124 , n25940 );
    not g22280 ( n25637 , n29884 );
    xnor g22281 ( n31584 , n8696 , n8657 );
    or g22282 ( n30325 , n9793 , n30328 );
    and g22283 ( n5127 , n11062 , n34306 );
    and g22284 ( n15900 , n5398 , n27028 );
    not g22285 ( n16175 , n4962 );
    nor g22286 ( n30505 , n4878 , n33173 );
    or g22287 ( n16871 , n22189 , n12833 );
    or g22288 ( n6768 , n32567 , n23187 );
    not g22289 ( n32897 , n25602 );
    or g22290 ( n10580 , n11543 , n35943 );
    or g22291 ( n20845 , n25048 , n27704 );
    or g22292 ( n8667 , n35802 , n16457 );
    or g22293 ( n4252 , n4758 , n29262 );
    xnor g22294 ( n18432 , n8123 , n6640 );
    xnor g22295 ( n25668 , n20972 , n1218 );
    and g22296 ( n33403 , n29551 , n29024 );
    xnor g22297 ( n28421 , n25926 , n16548 );
    or g22298 ( n30072 , n1768 , n23748 );
    or g22299 ( n192 , n22952 , n12389 );
    not g22300 ( n2518 , n6930 );
    xnor g22301 ( n29956 , n6790 , n32095 );
    or g22302 ( n34739 , n12711 , n33491 );
    and g22303 ( n21928 , n8272 , n30733 );
    and g22304 ( n25699 , n22345 , n3566 );
    xnor g22305 ( n26368 , n935 , n8879 );
    xnor g22306 ( n14676 , n25021 , n18026 );
    nor g22307 ( n26660 , n35645 , n11794 );
    not g22308 ( n19070 , n8432 );
    and g22309 ( n21126 , n4234 , n1139 );
    and g22310 ( n18209 , n29948 , n19597 );
    not g22311 ( n510 , n30181 );
    or g22312 ( n4202 , n29348 , n35043 );
    or g22313 ( n10443 , n8372 , n35748 );
    xnor g22314 ( n18252 , n21965 , n19984 );
    or g22315 ( n20618 , n31276 , n6397 );
    and g22316 ( n32116 , n25785 , n4572 );
    or g22317 ( n12168 , n29839 , n4670 );
    not g22318 ( n8720 , n15953 );
    xnor g22319 ( n31060 , n15603 , n10894 );
    not g22320 ( n24022 , n12326 );
    xnor g22321 ( n25977 , n20985 , n4779 );
    not g22322 ( n1498 , n15464 );
    xnor g22323 ( n4497 , n7645 , n1950 );
    and g22324 ( n34098 , n27059 , n11267 );
    not g22325 ( n8535 , n31472 );
    or g22326 ( n20951 , n9789 , n18192 );
    nor g22327 ( n29833 , n4758 , n17169 );
    or g22328 ( n1910 , n26531 , n29300 );
    nor g22329 ( n10138 , n24410 , n18934 );
    and g22330 ( n29913 , n6095 , n26708 );
    and g22331 ( n35438 , n17539 , n17801 );
    xnor g22332 ( n23361 , n11901 , n4962 );
    xnor g22333 ( n14720 , n18483 , n29810 );
    xnor g22334 ( n18139 , n9667 , n8362 );
    or g22335 ( n864 , n32095 , n21774 );
    or g22336 ( n18081 , n16882 , n36000 );
    or g22337 ( n12373 , n7420 , n1474 );
    not g22338 ( n7013 , n34897 );
    and g22339 ( n24491 , n7008 , n4212 );
    not g22340 ( n17190 , n32054 );
    or g22341 ( n29712 , n8479 , n17360 );
    or g22342 ( n28881 , n1745 , n9194 );
    or g22343 ( n23808 , n32179 , n14901 );
    and g22344 ( n32923 , n307 , n18779 );
    or g22345 ( n27655 , n34043 , n2980 );
    and g22346 ( n29599 , n35195 , n16864 );
    or g22347 ( n30019 , n24332 , n32419 );
    and g22348 ( n20636 , n18325 , n32754 );
    not g22349 ( n12064 , n21894 );
    or g22350 ( n11203 , n25043 , n28648 );
    and g22351 ( n32370 , n22028 , n2406 );
    or g22352 ( n4780 , n5306 , n28248 );
    and g22353 ( n15874 , n7039 , n18400 );
    or g22354 ( n31565 , n1697 , n3277 );
    xnor g22355 ( n7461 , n30493 , n32134 );
    xnor g22356 ( n10005 , n12832 , n18877 );
    buf g22357 ( n10400 , n4725 );
    and g22358 ( n566 , n32852 , n624 );
    or g22359 ( n23222 , n3852 , n3095 );
    or g22360 ( n20347 , n10514 , n21862 );
    xnor g22361 ( n24735 , n10716 , n11805 );
    nor g22362 ( n25240 , n2172 , n1236 );
    xnor g22363 ( n4484 , n31398 , n4626 );
    and g22364 ( n5402 , n28153 , n1212 );
    or g22365 ( n33549 , n2509 , n16594 );
    not g22366 ( n1320 , n3842 );
    nor g22367 ( n30277 , n4960 , n6275 );
    xnor g22368 ( n27149 , n22159 , n439 );
    or g22369 ( n14792 , n9993 , n17692 );
    or g22370 ( n28738 , n4926 , n384 );
    or g22371 ( n22104 , n10894 , n15376 );
    and g22372 ( n17155 , n33521 , n18222 );
    or g22373 ( n6281 , n3205 , n11927 );
    or g22374 ( n6086 , n3809 , n26473 );
    or g22375 ( n14012 , n20582 , n25255 );
    xnor g22376 ( n25385 , n33668 , n31700 );
    and g22377 ( n8685 , n20835 , n2987 );
    nor g22378 ( n5741 , n21190 , n5327 );
    or g22379 ( n24199 , n285 , n25592 );
    or g22380 ( n30981 , n20820 , n12128 );
    and g22381 ( n33149 , n34638 , n14114 );
    or g22382 ( n14810 , n32095 , n33844 );
    or g22383 ( n35903 , n23796 , n23930 );
    not g22384 ( n16017 , n9789 );
    or g22385 ( n21426 , n19219 , n14083 );
    and g22386 ( n36021 , n33418 , n21076 );
    and g22387 ( n8101 , n20136 , n28168 );
    xnor g22388 ( n16845 , n16065 , n4878 );
    or g22389 ( n15244 , n18379 , n29539 );
    and g22390 ( n13511 , n1610 , n13413 );
    or g22391 ( n3932 , n35964 , n4175 );
    buf g22392 ( n4912 , n9232 );
    and g22393 ( n22256 , n24927 , n13807 );
    xor g22394 ( n26099 , n28167 , n34666 );
    or g22395 ( n11674 , n5761 , n11781 );
    and g22396 ( n18270 , n30632 , n6801 );
    or g22397 ( n22935 , n8432 , n16250 );
    or g22398 ( n11947 , n33138 , n34537 );
    or g22399 ( n15980 , n7928 , n18059 );
    and g22400 ( n6272 , n2916 , n3179 );
    or g22401 ( n26832 , n34290 , n435 );
    and g22402 ( n21625 , n20770 , n21195 );
    and g22403 ( n14014 , n29131 , n11297 );
    xnor g22404 ( n24424 , n30130 , n11190 );
    and g22405 ( n25895 , n16589 , n30905 );
    or g22406 ( n30839 , n7754 , n14361 );
    or g22407 ( n26935 , n36010 , n14938 );
    nor g22408 ( n3713 , n16652 , n24625 );
    xnor g22409 ( n13252 , n33716 , n23604 );
    or g22410 ( n35161 , n1950 , n8044 );
    nor g22411 ( n7680 , n30099 , n12912 );
    and g22412 ( n33118 , n962 , n16493 );
    and g22413 ( n18321 , n21797 , n11588 );
    xnor g22414 ( n10706 , n35882 , n32351 );
    or g22415 ( n15264 , n6168 , n24672 );
    or g22416 ( n3705 , n4878 , n7173 );
    or g22417 ( n35662 , n2079 , n32507 );
    nor g22418 ( n28797 , n26083 , n14946 );
    or g22419 ( n11714 , n25767 , n28123 );
    or g22420 ( n8299 , n17611 , n12273 );
    xnor g22421 ( n13875 , n28004 , n31559 );
    and g22422 ( n9782 , n10280 , n21773 );
    or g22423 ( n2228 , n20712 , n20601 );
    xnor g22424 ( n8332 , n35167 , n16413 );
    and g22425 ( n20922 , n2233 , n21694 );
    and g22426 ( n2284 , n34144 , n5030 );
    and g22427 ( n32290 , n4218 , n28850 );
    xnor g22428 ( n23025 , n17262 , n4674 );
    and g22429 ( n28759 , n17925 , n10733 );
    and g22430 ( n29897 , n33212 , n15326 );
    xnor g22431 ( n34927 , n8334 , n33558 );
    or g22432 ( n33614 , n18141 , n19403 );
    or g22433 ( n11903 , n15886 , n18366 );
    or g22434 ( n30339 , n20899 , n14076 );
    not g22435 ( n13541 , n6132 );
    not g22436 ( n22498 , n30033 );
    or g22437 ( n2835 , n20085 , n2767 );
    or g22438 ( n19199 , n27690 , n14918 );
    xnor g22439 ( n12636 , n17322 , n19551 );
    and g22440 ( n35473 , n23917 , n5875 );
    and g22441 ( n35585 , n25386 , n17589 );
    and g22442 ( n31746 , n15897 , n6300 );
    or g22443 ( n4669 , n14607 , n24672 );
    or g22444 ( n855 , n24764 , n16388 );
    and g22445 ( n17133 , n21215 , n19220 );
    xnor g22446 ( n590 , n17691 , n27782 );
    or g22447 ( n10552 , n9549 , n20579 );
    xnor g22448 ( n28422 , n24218 , n16620 );
    and g22449 ( n16518 , n13966 , n23886 );
    or g22450 ( n25502 , n10211 , n2903 );
    and g22451 ( n29880 , n29100 , n4824 );
    or g22452 ( n7866 , n30952 , n35046 );
    not g22453 ( n20863 , n29808 );
    or g22454 ( n17501 , n9511 , n1375 );
    xnor g22455 ( n30385 , n32331 , n22291 );
    and g22456 ( n12319 , n30930 , n7595 );
    or g22457 ( n21414 , n18636 , n10417 );
    xnor g22458 ( n9564 , n9325 , n15403 );
    or g22459 ( n30580 , n6533 , n32539 );
    or g22460 ( n23889 , n27018 , n24479 );
    or g22461 ( n15794 , n20154 , n32071 );
    or g22462 ( n13800 , n23759 , n4490 );
    and g22463 ( n17535 , n29544 , n21834 );
    or g22464 ( n26490 , n22505 , n17829 );
    nor g22465 ( n3374 , n11432 , n6725 );
    or g22466 ( n13846 , n4878 , n25717 );
    or g22467 ( n4003 , n31272 , n31022 );
    or g22468 ( n258 , n32584 , n3002 );
    or g22469 ( n5764 , n15886 , n176 );
    nor g22470 ( n6800 , n10154 , n12500 );
    or g22471 ( n5207 , n9789 , n22994 );
    and g22472 ( n24976 , n13013 , n5836 );
    not g22473 ( n2607 , n3988 );
    xnor g22474 ( n12229 , n31086 , n20529 );
    and g22475 ( n23843 , n34093 , n29402 );
    or g22476 ( n25719 , n19551 , n21916 );
    or g22477 ( n3674 , n10697 , n26480 );
    or g22478 ( n9888 , n33648 , n25355 );
    not g22479 ( n20519 , n28982 );
    nor g22480 ( n5601 , n16225 , n9099 );
    or g22481 ( n28442 , n20448 , n18512 );
    or g22482 ( n33531 , n11445 , n20817 );
    nor g22483 ( n13493 , n17707 , n28184 );
    or g22484 ( n2900 , n1959 , n15675 );
    nor g22485 ( n27344 , n35288 , n219 );
    xnor g22486 ( n24664 , n11727 , n23604 );
    or g22487 ( n26722 , n8772 , n21154 );
    xnor g22488 ( n30516 , n4389 , n5996 );
    or g22489 ( n12682 , n18977 , n36000 );
    and g22490 ( n13132 , n18460 , n16477 );
    or g22491 ( n33984 , n1502 , n24592 );
    or g22492 ( n2147 , n24371 , n3803 );
    or g22493 ( n26233 , n3193 , n31128 );
    or g22494 ( n645 , n6937 , n20797 );
    or g22495 ( n589 , n18006 , n6502 );
    xnor g22496 ( n11018 , n16377 , n24371 );
    xnor g22497 ( n8660 , n3245 , n1104 );
    xnor g22498 ( n4435 , n28320 , n29379 );
    nor g22499 ( n32847 , n18917 , n20558 );
    or g22500 ( n17252 , n11508 , n6035 );
    or g22501 ( n17097 , n5287 , n10306 );
    and g22502 ( n23225 , n10828 , n11187 );
    xnor g22503 ( n14661 , n3984 , n15713 );
    and g22504 ( n3614 , n7619 , n24823 );
    or g22505 ( n20927 , n5335 , n34622 );
    or g22506 ( n34388 , n25602 , n8337 );
    or g22507 ( n27889 , n26680 , n30708 );
    buf g22508 ( n7726 , n34076 );
    xnor g22509 ( n10869 , n31183 , n13869 );
    not g22510 ( n20520 , n15886 );
    or g22511 ( n21794 , n28641 , n12162 );
    or g22512 ( n16637 , n28102 , n32412 );
    or g22513 ( n19563 , n30438 , n28652 );
    or g22514 ( n13339 , n33384 , n32359 );
    and g22515 ( n19653 , n28461 , n2593 );
    not g22516 ( n5222 , n16326 );
    or g22517 ( n23895 , n9327 , n33961 );
    xnor g22518 ( n31137 , n15923 , n18416 );
    or g22519 ( n33806 , n31772 , n13767 );
    xnor g22520 ( n14616 , n2647 , n32715 );
    xnor g22521 ( n16027 , n9454 , n23890 );
    not g22522 ( n22602 , n13416 );
    xnor g22523 ( n24483 , n23029 , n22332 );
    and g22524 ( n10602 , n7974 , n6754 );
    or g22525 ( n29576 , n12111 , n21977 );
    not g22526 ( n31300 , n12126 );
    not g22527 ( n31662 , n14983 );
    or g22528 ( n35130 , n27291 , n23740 );
    xnor g22529 ( n4578 , n28388 , n7215 );
    or g22530 ( n30895 , n17244 , n30646 );
    and g22531 ( n4095 , n19817 , n16282 );
    or g22532 ( n9822 , n3981 , n7877 );
    xnor g22533 ( n13078 , n9980 , n7388 );
    or g22534 ( n414 , n16016 , n27501 );
    buf g22535 ( n22322 , n22561 );
    or g22536 ( n6486 , n30460 , n30357 );
    and g22537 ( n8650 , n29028 , n17583 );
    xnor g22538 ( n25595 , n32349 , n12259 );
    or g22539 ( n8678 , n11505 , n22456 );
    or g22540 ( n31374 , n25836 , n14918 );
    or g22541 ( n24797 , n22285 , n6929 );
    and g22542 ( n2931 , n14462 , n18922 );
    or g22543 ( n29780 , n163 , n35211 );
    or g22544 ( n2177 , n30067 , n7955 );
    and g22545 ( n4840 , n1659 , n6974 );
    and g22546 ( n22621 , n4152 , n26328 );
    or g22547 ( n14701 , n3409 , n19241 );
    or g22548 ( n31504 , n20931 , n35143 );
    and g22549 ( n23535 , n1921 , n32261 );
    and g22550 ( n1098 , n29930 , n22287 );
    xnor g22551 ( n4008 , n31013 , n24704 );
    or g22552 ( n26489 , n25814 , n24259 );
    and g22553 ( n22070 , n13441 , n23619 );
    or g22554 ( n6188 , n17722 , n29626 );
    or g22555 ( n11768 , n5335 , n4641 );
    xnor g22556 ( n35495 , n26242 , n117 );
    not g22557 ( n21130 , n25602 );
    or g22558 ( n24887 , n1627 , n16457 );
    and g22559 ( n5611 , n9903 , n11416 );
    or g22560 ( n18306 , n3429 , n13059 );
    and g22561 ( n35931 , n31135 , n34851 );
    and g22562 ( n17250 , n20986 , n3211 );
    or g22563 ( n3706 , n23350 , n11312 );
    or g22564 ( n1751 , n5475 , n6613 );
    nor g22565 ( n5732 , n10329 , n14757 );
    and g22566 ( n23512 , n34445 , n10850 );
    or g22567 ( n13559 , n29084 , n5890 );
    xnor g22568 ( n10441 , n5612 , n3946 );
    and g22569 ( n11816 , n24163 , n15734 );
    or g22570 ( n9294 , n4288 , n3295 );
    or g22571 ( n869 , n24819 , n13015 );
    xnor g22572 ( n5306 , n31992 , n3 );
    and g22573 ( n7742 , n15239 , n31576 );
    or g22574 ( n10907 , n7540 , n27077 );
    or g22575 ( n6010 , n293 , n25728 );
    xnor g22576 ( n30080 , n21707 , n1950 );
    and g22577 ( n15603 , n11450 , n10111 );
    xnor g22578 ( n21273 , n9066 , n31799 );
    or g22579 ( n29351 , n14929 , n25567 );
    xnor g22580 ( n11125 , n24859 , n20964 );
    not g22581 ( n21342 , n25174 );
    and g22582 ( n5956 , n2260 , n13944 );
    and g22583 ( n21783 , n16449 , n17424 );
    nor g22584 ( n1522 , n21795 , n27091 );
    or g22585 ( n32813 , n23242 , n9153 );
    buf g22586 ( n9317 , n26112 );
    not g22587 ( n34310 , n18359 );
    nor g22588 ( n5221 , n9708 , n33956 );
    and g22589 ( n20887 , n16233 , n9381 );
    or g22590 ( n19529 , n14837 , n30292 );
    and g22591 ( n30515 , n19334 , n6679 );
    or g22592 ( n12995 , n29103 , n16594 );
    xnor g22593 ( n16373 , n3875 , n4727 );
    or g22594 ( n17694 , n1441 , n17111 );
    not g22595 ( n22732 , n22471 );
    nor g22596 ( n20954 , n23386 , n30904 );
    xnor g22597 ( n5888 , n1649 , n3946 );
    or g22598 ( n23904 , n24439 , n32634 );
    and g22599 ( n24890 , n8953 , n3599 );
    or g22600 ( n1249 , n33967 , n3489 );
    or g22601 ( n34468 , n25602 , n23507 );
    and g22602 ( n15172 , n7377 , n23893 );
    and g22603 ( n13817 , n31237 , n17796 );
    not g22604 ( n13960 , n10457 );
    xnor g22605 ( n16018 , n29701 , n25596 );
    or g22606 ( n11371 , n2714 , n3437 );
    xnor g22607 ( n6759 , n7944 , n4878 );
    or g22608 ( n28183 , n32818 , n31627 );
    or g22609 ( n6951 , n13055 , n19206 );
    or g22610 ( n12316 , n33878 , n32425 );
    or g22611 ( n10234 , n13689 , n29393 );
    or g22612 ( n31882 , n12352 , n4804 );
    nor g22613 ( n17025 , n11656 , n17757 );
    xnor g22614 ( n10329 , n27565 , n11789 );
    or g22615 ( n8853 , n34012 , n3863 );
    xnor g22616 ( n11296 , n9779 , n31272 );
    xnor g22617 ( n9454 , n22244 , n32584 );
    nor g22618 ( n4907 , n33324 , n10382 );
    and g22619 ( n8888 , n646 , n105 );
    and g22620 ( n15502 , n26123 , n13970 );
    or g22621 ( n5873 , n25005 , n29953 );
    or g22622 ( n25464 , n31215 , n6286 );
    and g22623 ( n30006 , n19818 , n23075 );
    or g22624 ( n24420 , n19274 , n22386 );
    or g22625 ( n8453 , n23863 , n2063 );
    or g22626 ( n16994 , n18848 , n19946 );
    xnor g22627 ( n30923 , n3737 , n34977 );
    or g22628 ( n6654 , n21087 , n5976 );
    xnor g22629 ( n1898 , n532 , n29926 );
    xnor g22630 ( n29458 , n26861 , n32801 );
    xnor g22631 ( n30136 , n32560 , n34112 );
    xnor g22632 ( n19371 , n26762 , n14808 );
    and g22633 ( n17335 , n25060 , n20424 );
    or g22634 ( n3018 , n29946 , n19241 );
    or g22635 ( n25905 , n4960 , n4587 );
    or g22636 ( n15420 , n11705 , n32226 );
    xnor g22637 ( n5614 , n23867 , n24170 );
    or g22638 ( n6165 , n7630 , n35043 );
    not g22639 ( n8000 , n2029 );
    or g22640 ( n25155 , n25690 , n2104 );
    or g22641 ( n19698 , n29123 , n34084 );
    nor g22642 ( n7994 , n21282 , n32386 );
    xnor g22643 ( n13748 , n8437 , n11190 );
    not g22644 ( n20798 , n30999 );
    not g22645 ( n31372 , n4367 );
    or g22646 ( n15127 , n14168 , n12511 );
    xnor g22647 ( n36077 , n253 , n24371 );
    nor g22648 ( n35217 , n8038 , n23257 );
    xnor g22649 ( n2435 , n19712 , n3704 );
    or g22650 ( n22581 , n2587 , n31310 );
    xnor g22651 ( n18000 , n32284 , n8432 );
    or g22652 ( n15508 , n4141 , n16744 );
    nor g22653 ( n34688 , n24954 , n16976 );
    or g22654 ( n18369 , n34497 , n26770 );
    or g22655 ( n33418 , n6982 , n24185 );
    xnor g22656 ( n28915 , n21775 , n20642 );
    or g22657 ( n12271 , n16641 , n2104 );
    or g22658 ( n7889 , n16620 , n1305 );
    and g22659 ( n410 , n1759 , n29785 );
    not g22660 ( n9617 , n23604 );
    xnor g22661 ( n3830 , n5360 , n32716 );
    not g22662 ( n7785 , n28853 );
    or g22663 ( n19364 , n827 , n4478 );
    or g22664 ( n34500 , n4176 , n17354 );
    or g22665 ( n24561 , n32438 , n9990 );
    nor g22666 ( n23517 , n31799 , n30256 );
    and g22667 ( n17494 , n22263 , n9382 );
    nor g22668 ( n28257 , n25852 , n18993 );
    xnor g22669 ( n6067 , n16578 , n21746 );
    and g22670 ( n35212 , n4160 , n14470 );
    and g22671 ( n31068 , n30518 , n28619 );
    xnor g22672 ( n29677 , n29851 , n13250 );
    xnor g22673 ( n2710 , n22006 , n6023 );
    or g22674 ( n3102 , n4288 , n32431 );
    or g22675 ( n6619 , n17623 , n28404 );
    xnor g22676 ( n9992 , n16114 , n13262 );
    nor g22677 ( n14154 , n10894 , n6371 );
    and g22678 ( n16343 , n22566 , n3820 );
    not g22679 ( n30444 , n18296 );
    xnor g22680 ( n16194 , n21396 , n11046 );
    xnor g22681 ( n20844 , n16279 , n16620 );
    and g22682 ( n35476 , n11243 , n17624 );
    and g22683 ( n21307 , n6723 , n12712 );
    or g22684 ( n12627 , n19217 , n19058 );
    or g22685 ( n20769 , n30401 , n20308 );
    or g22686 ( n20892 , n1000 , n33229 );
    or g22687 ( n34184 , n35325 , n11060 );
    or g22688 ( n20385 , n12524 , n2005 );
    xnor g22689 ( n2898 , n35939 , n724 );
    buf g22690 ( n20690 , n29533 );
    or g22691 ( n25442 , n12860 , n28631 );
    or g22692 ( n23100 , n16314 , n16543 );
    and g22693 ( n11014 , n27092 , n32311 );
    or g22694 ( n8264 , n11424 , n34971 );
    and g22695 ( n13731 , n30300 , n29142 );
    or g22696 ( n6603 , n2970 , n20629 );
    or g22697 ( n16091 , n17568 , n2091 );
    and g22698 ( n7273 , n31494 , n5882 );
    or g22699 ( n22984 , n18412 , n6760 );
    xnor g22700 ( n6823 , n10791 , n25106 );
    nor g22701 ( n35511 , n23953 , n16329 );
    or g22702 ( n16947 , n10968 , n34084 );
    not g22703 ( n21944 , n1950 );
    nor g22704 ( n15336 , n10894 , n13718 );
    and g22705 ( n19606 , n12965 , n2184 );
    or g22706 ( n10240 , n18379 , n18915 );
    or g22707 ( n7088 , n23461 , n33950 );
    or g22708 ( n34006 , n35375 , n14746 );
    and g22709 ( n30589 , n16056 , n22980 );
    or g22710 ( n20035 , n34897 , n23933 );
    or g22711 ( n15318 , n28594 , n17233 );
    not g22712 ( n17661 , n13198 );
    or g22713 ( n26618 , n32742 , n19105 );
    nor g22714 ( n16379 , n31289 , n18527 );
    or g22715 ( n5310 , n6765 , n29384 );
    xnor g22716 ( n32638 , n25746 , n16409 );
    and g22717 ( n28060 , n17922 , n32795 );
    or g22718 ( n1778 , n11455 , n21392 );
    or g22719 ( n10148 , n6296 , n128 );
    and g22720 ( n31359 , n15652 , n22792 );
    or g22721 ( n1226 , n32095 , n30175 );
    or g22722 ( n30418 , n34281 , n35543 );
    nor g22723 ( n19714 , n32095 , n35171 );
    xnor g22724 ( n24728 , n15197 , n4962 );
    and g22725 ( n29928 , n25582 , n9776 );
    or g22726 ( n23702 , n31172 , n18811 );
    xnor g22727 ( n19864 , n3654 , n3906 );
    and g22728 ( n35196 , n21181 , n11335 );
    nor g22729 ( n22934 , n6193 , n2105 );
    or g22730 ( n25650 , n31239 , n25831 );
    xnor g22731 ( n6652 , n9790 , n7540 );
    xnor g22732 ( n23087 , n10408 , n16135 );
    xnor g22733 ( n35765 , n28340 , n26517 );
    xnor g22734 ( n22174 , n6906 , n9658 );
    nor g22735 ( n37 , n19948 , n29954 );
    and g22736 ( n1046 , n576 , n630 );
    not g22737 ( n13390 , n18296 );
    nor g22738 ( n18995 , n19324 , n7639 );
    and g22739 ( n16249 , n21886 , n3272 );
    nor g22740 ( n25586 , n1600 , n13395 );
    or g22741 ( n3473 , n5886 , n13307 );
    nor g22742 ( n24636 , n8386 , n916 );
    not g22743 ( n2241 , n19939 );
    or g22744 ( n22266 , n20514 , n7261 );
    xnor g22745 ( n3618 , n11830 , n28287 );
    xnor g22746 ( n19577 , n16421 , n9789 );
    or g22747 ( n12722 , n7242 , n128 );
    or g22748 ( n5326 , n10673 , n28854 );
    or g22749 ( n33504 , n21796 , n11295 );
    or g22750 ( n28530 , n24999 , n16326 );
    or g22751 ( n15427 , n15299 , n12916 );
    or g22752 ( n20339 , n34009 , n11912 );
    and g22753 ( n31433 , n28097 , n8673 );
    and g22754 ( n23281 , n18863 , n10970 );
    or g22755 ( n6531 , n16379 , n3351 );
    not g22756 ( n33200 , n26365 );
    xnor g22757 ( n7838 , n11324 , n31368 );
    and g22758 ( n23157 , n16625 , n35364 );
    xnor g22759 ( n5253 , n12841 , n6349 );
    and g22760 ( n21496 , n26420 , n31026 );
    or g22761 ( n21955 , n28907 , n585 );
    and g22762 ( n34311 , n32366 , n26091 );
    and g22763 ( n34806 , n30202 , n11343 );
    or g22764 ( n818 , n20344 , n22946 );
    and g22765 ( n25836 , n5426 , n13406 );
    or g22766 ( n31528 , n25174 , n27089 );
    xnor g22767 ( n34271 , n25139 , n31289 );
    xnor g22768 ( n29271 , n3565 , n19984 );
    and g22769 ( n17750 , n35731 , n29828 );
    or g22770 ( n10513 , n6781 , n19490 );
    or g22771 ( n30699 , n22708 , n9507 );
    or g22772 ( n8593 , n2364 , n29896 );
    nor g22773 ( n25749 , n32095 , n9193 );
    xnor g22774 ( n6746 , n11363 , n34673 );
    or g22775 ( n27293 , n35927 , n27796 );
    or g22776 ( n31296 , n4357 , n9832 );
    not g22777 ( n21439 , n7730 );
    and g22778 ( n23177 , n27977 , n10713 );
    or g22779 ( n9114 , n1649 , n24333 );
    xnor g22780 ( n13671 , n23420 , n8701 );
    or g22781 ( n3246 , n32095 , n27897 );
    and g22782 ( n11794 , n7731 , n14238 );
    xnor g22783 ( n30352 , n12696 , n29273 );
    xnor g22784 ( n8001 , n22150 , n7105 );
    nor g22785 ( n29101 , n30742 , n8845 );
    xnor g22786 ( n31378 , n19467 , n26697 );
    or g22787 ( n31935 , n9550 , n26365 );
    and g22788 ( n24585 , n30350 , n3288 );
    xnor g22789 ( n17033 , n7350 , n9789 );
    xnor g22790 ( n3146 , n35802 , n16922 );
    and g22791 ( n6675 , n24848 , n20288 );
    not g22792 ( n13670 , n7699 );
    not g22793 ( n5549 , n471 );
    or g22794 ( n14752 , n13104 , n20797 );
    or g22795 ( n23468 , n20785 , n9675 );
    and g22796 ( n2024 , n32380 , n16089 );
    nor g22797 ( n16642 , n12393 , n32922 );
    or g22798 ( n4831 , n29060 , n2563 );
    or g22799 ( n17013 , n33515 , n16543 );
    or g22800 ( n26528 , n19551 , n21759 );
    nor g22801 ( n10812 , n15464 , n33317 );
    nor g22802 ( n8028 , n16922 , n31437 );
    or g22803 ( n10043 , n33304 , n11258 );
    nor g22804 ( n23305 , n32715 , n5670 );
    and g22805 ( n31624 , n2854 , n21895 );
    not g22806 ( n2353 , n26525 );
    or g22807 ( n1684 , n16922 , n8380 );
    xor g22808 ( n8250 , n3904 , n10532 );
    and g22809 ( n30289 , n7454 , n25118 );
    xnor g22810 ( n3916 , n13476 , n22096 );
    and g22811 ( n34578 , n6661 , n26185 );
    not g22812 ( n1096 , n33977 );
    and g22813 ( n21995 , n15434 , n10121 );
    or g22814 ( n19840 , n18823 , n9975 );
    and g22815 ( n7812 , n6673 , n31814 );
    and g22816 ( n35712 , n31244 , n35723 );
    not g22817 ( n25952 , n21042 );
    or g22818 ( n14198 , n4538 , n9030 );
    or g22819 ( n14136 , n25877 , n31773 );
    and g22820 ( n8655 , n34399 , n9906 );
    or g22821 ( n7403 , n22291 , n5093 );
    xnor g22822 ( n15818 , n7835 , n10424 );
    and g22823 ( n31336 , n30017 , n32208 );
    nor g22824 ( n30370 , n9539 , n13307 );
    or g22825 ( n6083 , n4288 , n11852 );
    or g22826 ( n1342 , n9005 , n8163 );
    or g22827 ( n7160 , n2818 , n28843 );
    and g22828 ( n32834 , n8033 , n25481 );
    or g22829 ( n30087 , n20109 , n13305 );
    and g22830 ( n15317 , n23669 , n15259 );
    or g22831 ( n20679 , n23482 , n29953 );
    and g22832 ( n23196 , n34678 , n29340 );
    or g22833 ( n6464 , n23919 , n22322 );
    and g22834 ( n33829 , n18294 , n13868 );
    and g22835 ( n30456 , n26775 , n26971 );
    nor g22836 ( n27691 , n35627 , n5138 );
    or g22837 ( n16828 , n13018 , n23365 );
    or g22838 ( n18751 , n5335 , n2863 );
    or g22839 ( n35413 , n33874 , n20765 );
    or g22840 ( n14501 , n10435 , n503 );
    or g22841 ( n35700 , n10864 , n29643 );
    or g22842 ( n19472 , n25465 , n22322 );
    xnor g22843 ( n18982 , n32433 , n28260 );
    or g22844 ( n14226 , n4351 , n28973 );
    nor g22845 ( n22534 , n35927 , n4841 );
    nor g22846 ( n31034 , n19551 , n13801 );
    or g22847 ( n4489 , n30634 , n23139 );
    or g22848 ( n32323 , n11349 , n25201 );
    or g22849 ( n12905 , n36064 , n11473 );
    xnor g22850 ( n31899 , n25465 , n30742 );
    or g22851 ( n5449 , n6427 , n26032 );
    nor g22852 ( n2933 , n24192 , n31962 );
    nor g22853 ( n21918 , n14291 , n20905 );
    and g22854 ( n575 , n10959 , n7620 );
    not g22855 ( n34305 , n7404 );
    not g22856 ( n20316 , n20716 );
    nor g22857 ( n9303 , n15279 , n10289 );
    or g22858 ( n7530 , n7540 , n9790 );
    and g22859 ( n3121 , n18656 , n28604 );
    or g22860 ( n8308 , n15298 , n22316 );
    xnor g22861 ( n29295 , n19236 , n8600 );
    xnor g22862 ( n12398 , n18132 , n35660 );
    and g22863 ( n8523 , n23767 , n16085 );
    and g22864 ( n13306 , n31726 , n32251 );
    not g22865 ( n31774 , n10902 );
    xnor g22866 ( n35152 , n32834 , n9789 );
    not g22867 ( n18686 , n7726 );
    nor g22868 ( n31181 , n8624 , n6548 );
    not g22869 ( n18849 , n6252 );
    and g22870 ( n6339 , n589 , n32613 );
    or g22871 ( n10474 , n2635 , n8663 );
    buf g22872 ( n2029 , n23651 );
    xnor g22873 ( n2188 , n5737 , n7471 );
    and g22874 ( n7905 , n17089 , n16651 );
    or g22875 ( n18035 , n17568 , n29381 );
    xnor g22876 ( n8740 , n15353 , n3056 );
    and g22877 ( n15240 , n20759 , n18011 );
    or g22878 ( n22435 , n18379 , n16631 );
    or g22879 ( n23009 , n6588 , n35141 );
    or g22880 ( n27747 , n12547 , n31067 );
    buf g22881 ( n7647 , n3681 );
    xnor g22882 ( n21479 , n24419 , n24371 );
    or g22883 ( n19815 , n2136 , n24653 );
    xnor g22884 ( n22391 , n26854 , n7066 );
    xnor g22885 ( n12714 , n29362 , n29330 );
    or g22886 ( n24815 , n5630 , n6950 );
    or g22887 ( n1473 , n19630 , n34484 );
    or g22888 ( n27639 , n4603 , n17974 );
    or g22889 ( n22216 , n6807 , n8723 );
    and g22890 ( n6116 , n14369 , n18687 );
    or g22891 ( n35433 , n22564 , n4937 );
    and g22892 ( n2647 , n26471 , n12584 );
    or g22893 ( n25551 , n29701 , n25596 );
    or g22894 ( n35975 , n19051 , n13743 );
    and g22895 ( n5044 , n2213 , n35353 );
    or g22896 ( n25300 , n24347 , n454 );
    not g22897 ( n30702 , n9431 );
    and g22898 ( n35280 , n35179 , n23553 );
    and g22899 ( n2639 , n32242 , n3528 );
    or g22900 ( n8441 , n6842 , n29592 );
    xnor g22901 ( n13336 , n16959 , n10894 );
    xnor g22902 ( n8214 , n2554 , n11231 );
    and g22903 ( n1251 , n18966 , n27802 );
    xnor g22904 ( n6634 , n21261 , n30742 );
    or g22905 ( n1659 , n27122 , n27625 );
    or g22906 ( n14331 , n27528 , n8963 );
    or g22907 ( n9712 , n14301 , n4203 );
    or g22908 ( n9887 , n27833 , n11712 );
    or g22909 ( n15436 , n17529 , n33113 );
    xnor g22910 ( n8414 , n19752 , n34161 );
    or g22911 ( n29254 , n36078 , n4439 );
    and g22912 ( n26852 , n31907 , n34468 );
    xnor g22913 ( n13205 , n9939 , n19337 );
    not g22914 ( n14908 , n8206 );
    and g22915 ( n21102 , n414 , n19056 );
    and g22916 ( n6503 , n17894 , n13597 );
    or g22917 ( n4843 , n32518 , n27447 );
    or g22918 ( n2807 , n4960 , n15649 );
    and g22919 ( n6114 , n22756 , n5335 );
    and g22920 ( n29831 , n29449 , n9455 );
    xnor g22921 ( n13922 , n14660 , n548 );
    xnor g22922 ( n16469 , n1935 , n9553 );
    or g22923 ( n12145 , n6009 , n20562 );
    and g22924 ( n9696 , n20583 , n4936 );
    xnor g22925 ( n22952 , n24035 , n11455 );
    and g22926 ( n25052 , n21825 , n1394 );
    xnor g22927 ( n10469 , n22013 , n11455 );
    or g22928 ( n30353 , n32516 , n31250 );
    or g22929 ( n22225 , n28878 , n22961 );
    nor g22930 ( n31536 , n25207 , n35616 );
    nor g22931 ( n27748 , n11455 , n30739 );
    or g22932 ( n6445 , n5417 , n30708 );
    or g22933 ( n4471 , n13779 , n29872 );
    or g22934 ( n3498 , n6153 , n27246 );
    or g22935 ( n6489 , n976 , n14342 );
    or g22936 ( n29548 , n14364 , n32680 );
    or g22937 ( n5948 , n18901 , n19945 );
    nor g22938 ( n26391 , n16620 , n35280 );
    and g22939 ( n5773 , n21599 , n31790 );
    nor g22940 ( n17814 , n23638 , n26826 );
    nor g22941 ( n25268 , n19762 , n2633 );
    or g22942 ( n5857 , n972 , n14076 );
    xnor g22943 ( n19497 , n2941 , n17399 );
    or g22944 ( n5668 , n16526 , n23069 );
    or g22945 ( n6623 , n24371 , n9385 );
    xnor g22946 ( n16788 , n14728 , n4962 );
    or g22947 ( n29828 , n26567 , n26023 );
    nor g22948 ( n5515 , n29316 , n8493 );
    or g22949 ( n21672 , n1297 , n27053 );
    not g22950 ( n26116 , n5377 );
    or g22951 ( n33064 , n18345 , n21977 );
    and g22952 ( n19429 , n31096 , n14893 );
    or g22953 ( n27042 , n14124 , n31549 );
    xnor g22954 ( n1581 , n35197 , n32095 );
    or g22955 ( n12400 , n26205 , n23713 );
    not g22956 ( n8376 , n32857 );
    or g22957 ( n4309 , n31439 , n33931 );
    or g22958 ( n4574 , n21054 , n14610 );
    or g22959 ( n26700 , n23838 , n5779 );
    and g22960 ( n1197 , n12439 , n6 );
    or g22961 ( n307 , n11821 , n16058 );
    or g22962 ( n23485 , n34344 , n21931 );
    or g22963 ( n19877 , n11046 , n2546 );
    and g22964 ( n27858 , n23140 , n14207 );
    and g22965 ( n14958 , n25120 , n32496 );
    xnor g22966 ( n14631 , n26622 , n3222 );
    and g22967 ( n17123 , n25946 , n9624 );
    not g22968 ( n29990 , n15886 );
    and g22969 ( n7209 , n32489 , n22164 );
    or g22970 ( n22073 , n10761 , n18477 );
    and g22971 ( n13760 , n29997 , n8858 );
    and g22972 ( n11188 , n1594 , n126 );
    and g22973 ( n25998 , n14210 , n32345 );
    and g22974 ( n7072 , n30198 , n31407 );
    or g22975 ( n6150 , n10155 , n20292 );
    not g22976 ( n11510 , n3488 );
    xor g22977 ( n28317 , n15873 , n31322 );
    xnor g22978 ( n34322 , n34790 , n27651 );
    or g22979 ( n7222 , n24159 , n3805 );
    or g22980 ( n27179 , n1648 , n19700 );
    xnor g22981 ( n6134 , n34134 , n19521 );
    and g22982 ( n22313 , n3983 , n571 );
    not g22983 ( n1230 , n7542 );
    or g22984 ( n1193 , n16692 , n16457 );
    nor g22985 ( n14300 , n16620 , n17382 );
    xnor g22986 ( n25181 , n1007 , n2339 );
    or g22987 ( n27256 , n15056 , n1557 );
    xnor g22988 ( n3731 , n3802 , n31799 );
    or g22989 ( n30336 , n8800 , n13886 );
    or g22990 ( n9196 , n9017 , n34084 );
    or g22991 ( n20772 , n17178 , n4318 );
    and g22992 ( n33604 , n11342 , n23513 );
    or g22993 ( n3825 , n9789 , n17499 );
    or g22994 ( n18740 , n19162 , n9872 );
    and g22995 ( n7709 , n27360 , n5633 );
    not g22996 ( n3782 , n6478 );
    xnor g22997 ( n25804 , n20527 , n2295 );
    or g22998 ( n28313 , n15429 , n17962 );
    or g22999 ( n11283 , n18359 , n34559 );
    or g23000 ( n13981 , n22979 , n8702 );
    and g23001 ( n2996 , n36063 , n13166 );
    or g23002 ( n21574 , n32095 , n13910 );
    nor g23003 ( n395 , n4962 , n26687 );
    or g23004 ( n30887 , n32816 , n26659 );
    nor g23005 ( n13114 , n9789 , n13776 );
    xnor g23006 ( n20229 , n13485 , n29843 );
    not g23007 ( n16802 , n26972 );
    or g23008 ( n17671 , n33831 , n29264 );
    or g23009 ( n27451 , n32235 , n3954 );
    and g23010 ( n7144 , n27373 , n27666 );
    or g23011 ( n2519 , n8167 , n35935 );
    or g23012 ( n28768 , n4541 , n15805 );
    or g23013 ( n25044 , n31215 , n14138 );
    xnor g23014 ( n26844 , n3320 , n14725 );
    xnor g23015 ( n1784 , n5065 , n8149 );
    and g23016 ( n15248 , n6166 , n33480 );
    and g23017 ( n19532 , n17077 , n26959 );
    or g23018 ( n26952 , n30749 , n30826 );
    and g23019 ( n5245 , n10426 , n33120 );
    not g23020 ( n12787 , n30742 );
    or g23021 ( n29399 , n5591 , n29672 );
    nor g23022 ( n8707 , n20464 , n19 );
    and g23023 ( n12648 , n10813 , n912 );
    and g23024 ( n10459 , n898 , n19144 );
    xnor g23025 ( n10114 , n21986 , n3870 );
    or g23026 ( n1486 , n13177 , n2299 );
    or g23027 ( n1123 , n10894 , n8088 );
    or g23028 ( n15868 , n35587 , n4595 );
    and g23029 ( n27804 , n15636 , n336 );
    not g23030 ( n21218 , n3884 );
    or g23031 ( n34332 , n20960 , n15256 );
    not g23032 ( n9431 , n12473 );
    and g23033 ( n26177 , n13143 , n22726 );
    and g23034 ( n3353 , n31988 , n5467 );
    or g23035 ( n36025 , n4582 , n27963 );
    or g23036 ( n21434 , n21303 , n1472 );
    and g23037 ( n16392 , n32173 , n34478 );
    nor g23038 ( n27491 , n1758 , n27667 );
    or g23039 ( n5068 , n2511 , n19336 );
    xnor g23040 ( n3265 , n13773 , n22604 );
    not g23041 ( n6663 , n3349 );
    or g23042 ( n1429 , n16090 , n3713 );
    and g23043 ( n469 , n25748 , n16351 );
    and g23044 ( n3870 , n20149 , n6901 );
    or g23045 ( n24184 , n26579 , n3575 );
    xnor g23046 ( n17967 , n14589 , n10894 );
    and g23047 ( n13059 , n9073 , n25985 );
    and g23048 ( n3414 , n26145 , n887 );
    or g23049 ( n28081 , n16135 , n22209 );
    xnor g23050 ( n969 , n25118 , n25742 );
    or g23051 ( n20736 , n1754 , n28837 );
    xnor g23052 ( n8803 , n20878 , n21547 );
    or g23053 ( n35510 , n8239 , n3188 );
    or g23054 ( n24762 , n24519 , n12596 );
    and g23055 ( n14106 , n3359 , n13706 );
    and g23056 ( n803 , n15396 , n14479 );
    and g23057 ( n50 , n6484 , n2478 );
    or g23058 ( n17103 , n22291 , n33746 );
    or g23059 ( n23124 , n24820 , n1320 );
    and g23060 ( n32272 , n4713 , n11057 );
    xnor g23061 ( n4174 , n12160 , n34353 );
    or g23062 ( n3844 , n16517 , n26023 );
    xnor g23063 ( n25331 , n29671 , n10582 );
    and g23064 ( n28553 , n15347 , n31682 );
    xnor g23065 ( n1805 , n5236 , n6972 );
    or g23066 ( n27534 , n10896 , n16567 );
    or g23067 ( n19369 , n28337 , n27827 );
    nor g23068 ( n21984 , n35927 , n17643 );
    not g23069 ( n13341 , n10355 );
    or g23070 ( n25069 , n9793 , n35737 );
    or g23071 ( n32767 , n11738 , n2798 );
    and g23072 ( n17879 , n24373 , n27183 );
    xnor g23073 ( n29269 , n18411 , n19984 );
    xnor g23074 ( n4089 , n3794 , n32963 );
    nor g23075 ( n4974 , n9789 , n25541 );
    xnor g23076 ( n14254 , n9351 , n19755 );
    and g23077 ( n19970 , n6217 , n14279 );
    or g23078 ( n9083 , n21847 , n10762 );
    or g23079 ( n25485 , n18418 , n29411 );
    or g23080 ( n34185 , n23517 , n15198 );
    or g23081 ( n21755 , n16644 , n25392 );
    and g23082 ( n33796 , n14514 , n31697 );
    xnor g23083 ( n18664 , n1940 , n9112 );
    and g23084 ( n2959 , n32028 , n15949 );
    xnor g23085 ( n33739 , n21120 , n3296 );
    not g23086 ( n19171 , n31662 );
    or g23087 ( n29093 , n16365 , n21673 );
    xnor g23088 ( n23190 , n4245 , n18662 );
    xnor g23089 ( n28532 , n309 , n33115 );
    or g23090 ( n14771 , n29390 , n21002 );
    not g23091 ( n32565 , n7238 );
    not g23092 ( n14563 , n3205 );
    and g23093 ( n17194 , n25826 , n30496 );
    or g23094 ( n1504 , n29833 , n12851 );
    or g23095 ( n34303 , n723 , n22427 );
    or g23096 ( n23620 , n19551 , n7256 );
    and g23097 ( n17677 , n15817 , n19185 );
    or g23098 ( n30495 , n27546 , n10289 );
    xnor g23099 ( n19300 , n2510 , n32688 );
    or g23100 ( n27784 , n25231 , n13085 );
    or g23101 ( n1604 , n13763 , n25052 );
    or g23102 ( n10890 , n31056 , n5428 );
    or g23103 ( n28612 , n23352 , n19173 );
    or g23104 ( n16772 , n22745 , n21608 );
    or g23105 ( n25439 , n15686 , n15717 );
    not g23106 ( n7913 , n1950 );
    xnor g23107 ( n33232 , n11514 , n33942 );
    xnor g23108 ( n3711 , n32102 , n27308 );
    or g23109 ( n15196 , n25930 , n19155 );
    or g23110 ( n23898 , n8432 , n23918 );
    nor g23111 ( n10903 , n4878 , n36078 );
    and g23112 ( n25832 , n25959 , n7158 );
    or g23113 ( n15133 , n6979 , n35935 );
    and g23114 ( n11567 , n21511 , n24366 );
    or g23115 ( n13334 , n16922 , n19050 );
    xnor g23116 ( n8049 , n16585 , n19551 );
    or g23117 ( n28891 , n28074 , n1856 );
    or g23118 ( n13191 , n32403 , n4952 );
    or g23119 ( n14180 , n27428 , n29407 );
    and g23120 ( n24729 , n26805 , n21528 );
    and g23121 ( n22475 , n3597 , n23181 );
    or g23122 ( n35839 , n9476 , n35630 );
    and g23123 ( n7289 , n30567 , n13331 );
    or g23124 ( n1670 , n3751 , n949 );
    nor g23125 ( n6845 , n30802 , n32379 );
    and g23126 ( n24339 , n20241 , n5873 );
    or g23127 ( n23285 , n21619 , n19089 );
    or g23128 ( n5012 , n15064 , n13664 );
    and g23129 ( n11120 , n11275 , n8942 );
    and g23130 ( n24355 , n4501 , n25082 );
    or g23131 ( n6382 , n28519 , n4203 );
    or g23132 ( n21446 , n12375 , n585 );
    nor g23133 ( n29279 , n5335 , n22756 );
    xnor g23134 ( n34836 , n24857 , n28104 );
    or g23135 ( n24244 , n11942 , n27963 );
    or g23136 ( n14470 , n17324 , n12996 );
    or g23137 ( n34617 , n5169 , n20817 );
    and g23138 ( n34397 , n33625 , n5074 );
    nor g23139 ( n7354 , n15956 , n6276 );
    xnor g23140 ( n8176 , n4011 , n20082 );
    or g23141 ( n2754 , n9140 , n32425 );
    or g23142 ( n25643 , n21113 , n12533 );
    and g23143 ( n13797 , n33966 , n30104 );
    or g23144 ( n24903 , n17889 , n23033 );
    or g23145 ( n872 , n6074 , n5972 );
    and g23146 ( n22272 , n26542 , n5524 );
    xnor g23147 ( n26376 , n14654 , n4288 );
    or g23148 ( n15193 , n1739 , n20601 );
    nor g23149 ( n11282 , n4960 , n17716 );
    or g23150 ( n26901 , n24015 , n24299 );
    xnor g23151 ( n25518 , n25448 , n4288 );
    or g23152 ( n5805 , n935 , n15538 );
    or g23153 ( n29440 , n5067 , n4800 );
    not g23154 ( n9308 , n35710 );
    nor g23155 ( n9539 , n3770 , n21294 );
    and g23156 ( n13299 , n10263 , n35316 );
    or g23157 ( n2668 , n27614 , n15188 );
    or g23158 ( n29180 , n21591 , n26480 );
    xnor g23159 ( n24280 , n6172 , n8432 );
    or g23160 ( n13172 , n31289 , n35580 );
    nor g23161 ( n140 , n5475 , n32928 );
    nor g23162 ( n2075 , n11046 , n29361 );
    or g23163 ( n10447 , n31229 , n4254 );
    xnor g23164 ( n32055 , n636 , n17751 );
    or g23165 ( n34755 , n4960 , n9020 );
    xnor g23166 ( n10492 , n8655 , n35927 );
    or g23167 ( n11009 , n20222 , n8153 );
    and g23168 ( n15975 , n35020 , n7735 );
    and g23169 ( n22320 , n18287 , n2353 );
    or g23170 ( n22880 , n13349 , n14699 );
    xnor g23171 ( n19663 , n11413 , n24549 );
    or g23172 ( n26804 , n25204 , n11996 );
    or g23173 ( n190 , n4243 , n13203 );
    or g23174 ( n12584 , n30185 , n31554 );
    or g23175 ( n23831 , n31559 , n30591 );
    not g23176 ( n15529 , n28561 );
    or g23177 ( n27366 , n4878 , n3416 );
    or g23178 ( n5784 , n25150 , n13912 );
    and g23179 ( n18033 , n30472 , n31789 );
    or g23180 ( n16779 , n15464 , n16102 );
    or g23181 ( n20578 , n18897 , n28438 );
    and g23182 ( n19441 , n6893 , n3698 );
    or g23183 ( n22028 , n22100 , n29562 );
    buf g23184 ( n5972 , n4478 );
    or g23185 ( n3439 , n469 , n22858 );
    or g23186 ( n28146 , n33538 , n7288 );
    and g23187 ( n3517 , n6838 , n33877 );
    not g23188 ( n26261 , n1761 );
    or g23189 ( n3688 , n13385 , n33466 );
    and g23190 ( n33676 , n27147 , n2291 );
    nor g23191 ( n20871 , n17568 , n25997 );
    or g23192 ( n26451 , n6215 , n32329 );
    xor g23193 ( n5737 , n33582 , n35927 );
    or g23194 ( n26138 , n31289 , n4858 );
    xnor g23195 ( n1391 , n5318 , n7114 );
    and g23196 ( n11756 , n21257 , n35976 );
    and g23197 ( n30960 , n8729 , n17528 );
    or g23198 ( n20976 , n8268 , n3424 );
    xnor g23199 ( n24933 , n7318 , n17376 );
    and g23200 ( n28159 , n35932 , n14147 );
    xnor g23201 ( n33207 , n12331 , n9658 );
    and g23202 ( n32336 , n3140 , n6301 );
    or g23203 ( n8572 , n29418 , n26653 );
    or g23204 ( n7750 , n12570 , n19560 );
    nor g23205 ( n17651 , n27135 , n26103 );
    or g23206 ( n16233 , n22353 , n25447 );
    xnor g23207 ( n204 , n35576 , n11936 );
    and g23208 ( n2701 , n11355 , n10894 );
    or g23209 ( n20045 , n25555 , n34657 );
    and g23210 ( n17505 , n19212 , n20632 );
    or g23211 ( n15983 , n28599 , n4363 );
    and g23212 ( n13677 , n29877 , n13382 );
    and g23213 ( n3818 , n13865 , n11898 );
    and g23214 ( n35200 , n30402 , n1523 );
    or g23215 ( n22617 , n16833 , n19241 );
    or g23216 ( n10665 , n9647 , n17233 );
    or g23217 ( n32831 , n6664 , n7192 );
    nor g23218 ( n21513 , n32857 , n16512 );
    or g23219 ( n22731 , n23359 , n19241 );
    or g23220 ( n24398 , n29884 , n27176 );
    and g23221 ( n16490 , n28528 , n16358 );
    or g23222 ( n16281 , n26541 , n18486 );
    not g23223 ( n33863 , n24371 );
    nor g23224 ( n13395 , n35682 , n21811 );
    or g23225 ( n27128 , n396 , n27501 );
    xnor g23226 ( n12226 , n15182 , n27633 );
    not g23227 ( n25304 , n1950 );
    xnor g23228 ( n3209 , n12173 , n32812 );
    or g23229 ( n34126 , n15886 , n19447 );
    or g23230 ( n22460 , n30367 , n27801 );
    or g23231 ( n232 , n1575 , n17111 );
    or g23232 ( n7475 , n9238 , n9915 );
    xnor g23233 ( n26842 , n28494 , n26429 );
    or g23234 ( n11815 , n24407 , n11850 );
    nor g23235 ( n16059 , n15696 , n6995 );
    nor g23236 ( n24204 , n34021 , n20675 );
    xor g23237 ( n27613 , n20009 , n31594 );
    and g23238 ( n19612 , n34833 , n19083 );
    and g23239 ( n35547 , n6242 , n16224 );
    or g23240 ( n8279 , n5954 , n11850 );
    or g23241 ( n33620 , n33334 , n23299 );
    or g23242 ( n9904 , n32597 , n14903 );
    or g23243 ( n11482 , n852 , n9930 );
    or g23244 ( n7736 , n25181 , n23921 );
    or g23245 ( n13906 , n12648 , n31536 );
    and g23246 ( n29136 , n30886 , n11865 );
    or g23247 ( n4705 , n4288 , n28182 );
    xnor g23248 ( n34793 , n8247 , n32095 );
    or g23249 ( n27389 , n25033 , n25592 );
    xnor g23250 ( n1248 , n36075 , n7649 );
    nor g23251 ( n27464 , n6161 , n16503 );
    or g23252 ( n29200 , n12433 , n9194 );
    and g23253 ( n4804 , n15618 , n35612 );
    xnor g23254 ( n13580 , n26001 , n4960 );
    not g23255 ( n9858 , n4960 );
    and g23256 ( n14356 , n27182 , n31023 );
    not g23257 ( n30397 , n4960 );
    or g23258 ( n21730 , n5753 , n23462 );
    xnor g23259 ( n29089 , n10834 , n18393 );
    or g23260 ( n1348 , n24371 , n21603 );
    not g23261 ( n10275 , n31799 );
    xnor g23262 ( n2954 , n32989 , n29713 );
    not g23263 ( n13823 , n31808 );
    or g23264 ( n30474 , n4801 , n11593 );
    xnor g23265 ( n9483 , n5353 , n6336 );
    or g23266 ( n20965 , n31289 , n30133 );
    or g23267 ( n11503 , n12514 , n23655 );
    or g23268 ( n21364 , n9047 , n634 );
    or g23269 ( n14580 , n10645 , n35304 );
    xnor g23270 ( n31956 , n2714 , n5287 );
    or g23271 ( n32807 , n19607 , n23462 );
    or g23272 ( n32213 , n11455 , n329 );
    xnor g23273 ( n6488 , n16810 , n25824 );
    and g23274 ( n32625 , n23700 , n8115 );
    or g23275 ( n35530 , n22254 , n20817 );
    and g23276 ( n21606 , n22225 , n27255 );
    and g23277 ( n33161 , n29443 , n31030 );
    and g23278 ( n29178 , n14498 , n13365 );
    or g23279 ( n16138 , n20660 , n19241 );
    or g23280 ( n32012 , n10114 , n24696 );
    or g23281 ( n23341 , n23793 , n16797 );
    or g23282 ( n5848 , n24646 , n763 );
    and g23283 ( n17643 , n273 , n33303 );
    or g23284 ( n11213 , n4288 , n19248 );
    xnor g23285 ( n25457 , n22632 , n16293 );
    or g23286 ( n22430 , n17498 , n3736 );
    and g23287 ( n24185 , n15217 , n6967 );
    xnor g23288 ( n17635 , n26677 , n9108 );
    and g23289 ( n34235 , n7092 , n11979 );
    or g23290 ( n6865 , n6299 , n20253 );
    or g23291 ( n34202 , n10894 , n21463 );
    or g23292 ( n33095 , n33369 , n4249 );
    nor g23293 ( n7515 , n27571 , n32697 );
    xnor g23294 ( n15881 , n23181 , n3597 );
    not g23295 ( n14887 , n16252 );
    and g23296 ( n17178 , n8825 , n23932 );
    or g23297 ( n12765 , n25602 , n16505 );
    or g23298 ( n21743 , n25913 , n4175 );
    or g23299 ( n11145 , n9265 , n26659 );
    or g23300 ( n23473 , n25174 , n27122 );
    and g23301 ( n6820 , n25989 , n13103 );
    or g23302 ( n6573 , n13129 , n33561 );
    xnor g23303 ( n8290 , n28827 , n5335 );
    and g23304 ( n17769 , n13641 , n4888 );
    and g23305 ( n11360 , n33807 , n16022 );
    or g23306 ( n27987 , n23740 , n17233 );
    xnor g23307 ( n19646 , n783 , n20285 );
    not g23308 ( n18749 , n23554 );
    or g23309 ( n28644 , n34179 , n1034 );
    and g23310 ( n32567 , n26635 , n13921 );
    and g23311 ( n23387 , n5536 , n7040 );
    or g23312 ( n31560 , n5999 , n7673 );
    and g23313 ( n20216 , n28755 , n13398 );
    xnor g23314 ( n13818 , n20652 , n7169 );
    or g23315 ( n31615 , n2385 , n4246 );
    and g23316 ( n2394 , n4559 , n5265 );
    and g23317 ( n23060 , n9807 , n24056 );
    xnor g23318 ( n22633 , n7272 , n29713 );
    nor g23319 ( n31384 , n27226 , n5163 );
    or g23320 ( n6204 , n13673 , n23503 );
    and g23321 ( n2960 , n15508 , n10388 );
    not g23322 ( n16635 , n833 );
    or g23323 ( n22083 , n5726 , n13000 );
    nor g23324 ( n2277 , n7540 , n15914 );
    and g23325 ( n530 , n11417 , n4197 );
    xnor g23326 ( n4527 , n25608 , n24371 );
    or g23327 ( n11650 , n5581 , n25418 );
    not g23328 ( n33360 , n25909 );
    or g23329 ( n8267 , n21152 , n1558 );
    xnor g23330 ( n6605 , n33015 , n19551 );
    or g23331 ( n34576 , n30422 , n12465 );
    or g23332 ( n21334 , n1126 , n8159 );
    or g23333 ( n23639 , n4442 , n3856 );
    or g23334 ( n13398 , n34941 , n578 );
    or g23335 ( n27463 , n16373 , n34342 );
    or g23336 ( n12939 , n8432 , n5460 );
    xnor g23337 ( n1829 , n34705 , n20181 );
    xnor g23338 ( n16366 , n34349 , n14264 );
    and g23339 ( n31356 , n35213 , n25278 );
    xnor g23340 ( n26115 , n28979 , n3474 );
    xnor g23341 ( n3231 , n28145 , n34413 );
    or g23342 ( n25679 , n13294 , n21173 );
    or g23343 ( n12020 , n31783 , n10315 );
    or g23344 ( n7740 , n29890 , n5570 );
    nor g23345 ( n18529 , n7540 , n15375 );
    or g23346 ( n28823 , n7299 , n19241 );
    not g23347 ( n31370 , n25174 );
    and g23348 ( n21040 , n19472 , n4332 );
    or g23349 ( n11124 , n19936 , n33177 );
    and g23350 ( n29882 , n33329 , n9086 );
    and g23351 ( n30223 , n6636 , n21335 );
    or g23352 ( n33794 , n7540 , n9637 );
    xnor g23353 ( n12455 , n6589 , n1950 );
    xnor g23354 ( n9547 , n28966 , n14137 );
    or g23355 ( n33481 , n34524 , n9951 );
    or g23356 ( n35785 , n18063 , n30646 );
    or g23357 ( n9656 , n14842 , n22858 );
    not g23358 ( n25133 , n24694 );
    not g23359 ( n8430 , n26781 );
    xnor g23360 ( n9583 , n27844 , n9793 );
    xnor g23361 ( n24662 , n30322 , n1207 );
    nor g23362 ( n26197 , n17568 , n29253 );
    xnor g23363 ( n6031 , n5704 , n31559 );
    or g23364 ( n26381 , n4878 , n18576 );
    xnor g23365 ( n21209 , n35681 , n13161 );
    or g23366 ( n14282 , n19875 , n4772 );
    and g23367 ( n32348 , n34975 , n7335 );
    not g23368 ( n1815 , n4878 );
    and g23369 ( n3277 , n5121 , n7799 );
    or g23370 ( n28218 , n1687 , n585 );
    and g23371 ( n4722 , n12990 , n8335 );
    or g23372 ( n27608 , n29865 , n26919 );
    nor g23373 ( n19632 , n8182 , n17354 );
    and g23374 ( n11666 , n21487 , n31222 );
    not g23375 ( n32969 , n30204 );
    or g23376 ( n399 , n11046 , n27283 );
    not g23377 ( n12654 , n29713 );
    not g23378 ( n26455 , n15729 );
    not g23379 ( n1884 , n23604 );
    xnor g23380 ( n14252 , n4993 , n4632 );
    and g23381 ( n19159 , n2419 , n14908 );
    xnor g23382 ( n4216 , n33148 , n10894 );
    and g23383 ( n13564 , n9412 , n11322 );
    or g23384 ( n21642 , n5122 , n25773 );
    or g23385 ( n3412 , n26247 , n31627 );
    and g23386 ( n2962 , n29359 , n31295 );
    not g23387 ( n21212 , n31289 );
    not g23388 ( n8597 , n22980 );
    xnor g23389 ( n20329 , n31239 , n10894 );
    nor g23390 ( n9085 , n24054 , n29203 );
    and g23391 ( n13270 , n29616 , n21161 );
    not g23392 ( n11527 , n8610 );
    and g23393 ( n32597 , n8519 , n30031 );
    xnor g23394 ( n8224 , n25708 , n13784 );
    nor g23395 ( n8263 , n4288 , n21928 );
    nor g23396 ( n21582 , n34679 , n23280 );
    and g23397 ( n22158 , n2976 , n6564 );
    xnor g23398 ( n2417 , n7058 , n32857 );
    nor g23399 ( n33586 , n7540 , n5301 );
    or g23400 ( n10209 , n35933 , n9930 );
    buf g23401 ( n9915 , n8366 );
    and g23402 ( n6115 , n27999 , n32471 );
    or g23403 ( n624 , n15132 , n8203 );
    and g23404 ( n6077 , n34466 , n14175 );
    and g23405 ( n290 , n26092 , n7452 );
    and g23406 ( n5507 , n33371 , n15134 );
    and g23407 ( n17267 , n600 , n619 );
    nor g23408 ( n32321 , n35479 , n17945 );
    not g23409 ( n3595 , n35051 );
    xnor g23410 ( n1099 , n10021 , n19551 );
    and g23411 ( n5166 , n30347 , n27648 );
    or g23412 ( n21516 , n33965 , n14129 );
    nor g23413 ( n4281 , n3946 , n7310 );
    not g23414 ( n29237 , n23604 );
    or g23415 ( n35453 , n16254 , n16749 );
    not g23416 ( n35572 , n34256 );
    and g23417 ( n20213 , n18295 , n6175 );
    xnor g23418 ( n23268 , n1656 , n11190 );
    nor g23419 ( n34531 , n19984 , n11478 );
    and g23420 ( n22129 , n10237 , n35031 );
    or g23421 ( n16544 , n4015 , n28404 );
    or g23422 ( n32334 , n29839 , n32477 );
    or g23423 ( n23214 , n11654 , n27701 );
    or g23424 ( n9208 , n10627 , n13936 );
    not g23425 ( n23219 , n31799 );
    or g23426 ( n23350 , n31575 , n7500 );
    and g23427 ( n6714 , n6102 , n35945 );
    not g23428 ( n17109 , n19200 );
    or g23429 ( n2857 , n8432 , n9500 );
    or g23430 ( n3067 , n16173 , n14554 );
    or g23431 ( n1111 , n21281 , n33121 );
    nor g23432 ( n5224 , n29713 , n23233 );
    or g23433 ( n24448 , n30107 , n908 );
    or g23434 ( n23553 , n8084 , n21859 );
    or g23435 ( n34588 , n909 , n23287 );
    or g23436 ( n579 , n35356 , n30708 );
    or g23437 ( n1527 , n7540 , n29478 );
    or g23438 ( n21871 , n32857 , n33728 );
    not g23439 ( n23037 , n23422 );
    or g23440 ( n22384 , n8890 , n24259 );
    or g23441 ( n8995 , n15886 , n13769 );
    or g23442 ( n26492 , n8831 , n12843 );
    xnor g23443 ( n18781 , n29881 , n11190 );
    not g23444 ( n20074 , n33596 );
    not g23445 ( n29659 , n32089 );
    not g23446 ( n25067 , n1511 );
    xnor g23447 ( n25231 , n35746 , n19551 );
    or g23448 ( n25733 , n12319 , n10336 );
    or g23449 ( n24584 , n8015 , n24696 );
    and g23450 ( n28666 , n14703 , n31329 );
    and g23451 ( n12823 , n27768 , n5525 );
    or g23452 ( n11649 , n4258 , n14706 );
    or g23453 ( n18753 , n32672 , n19490 );
    xnor g23454 ( n9277 , n30471 , n1264 );
    or g23455 ( n21086 , n10976 , n34745 );
    or g23456 ( n26986 , n15464 , n12727 );
    or g23457 ( n28042 , n24546 , n19336 );
    or g23458 ( n33033 , n25747 , n34989 );
    xnor g23459 ( n8068 , n17986 , n19551 );
    or g23460 ( n31519 , n10425 , n9194 );
    xnor g23461 ( n25972 , n9184 , n16399 );
    and g23462 ( n28096 , n34428 , n25736 );
    or g23463 ( n30856 , n15861 , n34822 );
    xnor g23464 ( n29274 , n11846 , n15886 );
    and g23465 ( n24040 , n10969 , n32690 );
    and g23466 ( n3704 , n33484 , n34956 );
    xnor g23467 ( n19246 , n5363 , n4049 );
    or g23468 ( n4964 , n19984 , n29628 );
    or g23469 ( n23426 , n24305 , n5515 );
    or g23470 ( n7210 , n18379 , n5937 );
    not g23471 ( n8677 , n30742 );
    xnor g23472 ( n29586 , n32272 , n32857 );
    or g23473 ( n14297 , n8688 , n16166 );
    and g23474 ( n11605 , n18880 , n15327 );
    or g23475 ( n10844 , n18935 , n19173 );
    and g23476 ( n21227 , n30841 , n6265 );
    xnor g23477 ( n28903 , n31775 , n5335 );
    xnor g23478 ( n17482 , n14623 , n3205 );
    or g23479 ( n35185 , n5669 , n9103 );
    or g23480 ( n25360 , n1124 , n20620 );
    xnor g23481 ( n28954 , n24596 , n7657 );
    xnor g23482 ( n21160 , n31210 , n31048 );
    or g23483 ( n28785 , n11796 , n12879 );
    not g23484 ( n29065 , n27780 );
    and g23485 ( n9623 , n23272 , n10046 );
    not g23486 ( n10734 , n17751 );
    and g23487 ( n178 , n5853 , n15837 );
    xor g23488 ( n8692 , n12537 , n25727 );
    xnor g23489 ( n33286 , n6396 , n25965 );
    and g23490 ( n2625 , n27830 , n8021 );
    and g23491 ( n23218 , n2695 , n14053 );
    not g23492 ( n24634 , n20558 );
    or g23493 ( n7600 , n9789 , n448 );
    buf g23494 ( n19948 , n8179 );
    or g23495 ( n31347 , n26582 , n4478 );
    or g23496 ( n30548 , n17650 , n31627 );
    or g23497 ( n1929 , n29713 , n6296 );
    xnor g23498 ( n7752 , n25911 , n28512 );
    and g23499 ( n5456 , n18731 , n34669 );
    not g23500 ( n1841 , n18471 );
    and g23501 ( n12042 , n2239 , n33692 );
    or g23502 ( n16677 , n10268 , n35841 );
    and g23503 ( n4338 , n32768 , n18328 );
    xnor g23504 ( n33274 , n10454 , n15213 );
    or g23505 ( n3534 , n10894 , n20785 );
    or g23506 ( n23302 , n31137 , n28404 );
    and g23507 ( n1156 , n26152 , n20089 );
    xnor g23508 ( n21668 , n28956 , n31117 );
    or g23509 ( n1838 , n30115 , n3239 );
    xnor g23510 ( n23967 , n16880 , n23532 );
    xnor g23511 ( n4169 , n12624 , n31198 );
    xnor g23512 ( n16825 , n11604 , n28799 );
    xnor g23513 ( n26623 , n30573 , n8293 );
    or g23514 ( n18363 , n29940 , n32782 );
    nor g23515 ( n1671 , n16620 , n11798 );
    or g23516 ( n2086 , n5067 , n8154 );
    or g23517 ( n23964 , n29136 , n10634 );
    nor g23518 ( n27051 , n32857 , n10288 );
    nor g23519 ( n3860 , n29839 , n4954 );
    or g23520 ( n31431 , n23481 , n30988 );
    or g23521 ( n28086 , n784 , n19812 );
    not g23522 ( n27620 , n31056 );
    xnor g23523 ( n15719 , n25665 , n277 );
    or g23524 ( n23104 , n5745 , n1414 );
    buf g23525 ( n16659 , n3276 );
    and g23526 ( n33815 , n12061 , n10883 );
    and g23527 ( n21450 , n32599 , n18421 );
    or g23528 ( n31351 , n19459 , n28668 );
    xnor g23529 ( n35436 , n3837 , n24371 );
    or g23530 ( n5082 , n10011 , n7448 );
    or g23531 ( n23683 , n7016 , n11518 );
    or g23532 ( n16355 , n30546 , n16423 );
    xnor g23533 ( n30164 , n28465 , n15886 );
    xnor g23534 ( n28446 , n35345 , n15337 );
    xnor g23535 ( n23675 , n6710 , n30448 );
    and g23536 ( n8283 , n25551 , n3047 );
    not g23537 ( n22856 , n28987 );
    or g23538 ( n26720 , n7940 , n11666 );
    and g23539 ( n3465 , n27350 , n18340 );
    or g23540 ( n14060 , n19578 , n30563 );
    or g23541 ( n35981 , n4100 , n26988 );
    not g23542 ( n30807 , n1578 );
    xnor g23543 ( n291 , n1925 , n28134 );
    buf g23544 ( n29562 , n13905 );
    xnor g23545 ( n26540 , n155 , n4870 );
    or g23546 ( n29694 , n16534 , n13305 );
    xnor g23547 ( n1573 , n33632 , n1341 );
    or g23548 ( n19183 , n9249 , n28248 );
    or g23549 ( n26934 , n25041 , n10432 );
    not g23550 ( n13886 , n28969 );
    or g23551 ( n19181 , n22774 , n19547 );
    or g23552 ( n1782 , n25541 , n19084 );
    and g23553 ( n15084 , n28201 , n2181 );
    buf g23554 ( n22200 , n32983 );
    or g23555 ( n5001 , n17373 , n6950 );
    or g23556 ( n25504 , n11537 , n23187 );
    xnor g23557 ( n14294 , n27352 , n27570 );
    or g23558 ( n23772 , n30742 , n28099 );
    or g23559 ( n30706 , n3895 , n34537 );
    not g23560 ( n2287 , n6220 );
    or g23561 ( n35582 , n20302 , n26002 );
    nor g23562 ( n30968 , n4372 , n26023 );
    and g23563 ( n11113 , n9898 , n26870 );
    and g23564 ( n32793 , n35922 , n21048 );
    and g23565 ( n5561 , n6621 , n19611 );
    xnor g23566 ( n6176 , n33943 , n19189 );
    and g23567 ( n6054 , n15121 , n11408 );
    and g23568 ( n27444 , n2978 , n8996 );
    xnor g23569 ( n15986 , n30475 , n8310 );
    xnor g23570 ( n10236 , n10881 , n35820 );
    nor g23571 ( n12311 , n25174 , n24765 );
    and g23572 ( n18978 , n27908 , n1227 );
    xnor g23573 ( n25537 , n23958 , n35203 );
    or g23574 ( n8054 , n25672 , n11833 );
    not g23575 ( n19560 , n32692 );
    and g23576 ( n13340 , n2296 , n18872 );
    not g23577 ( n1911 , n22980 );
    xnor g23578 ( n35899 , n546 , n29727 );
    xnor g23579 ( n18824 , n24941 , n15464 );
    or g23580 ( n21752 , n4497 , n33331 );
    xnor g23581 ( n8870 , n3921 , n15094 );
    and g23582 ( n12958 , n31723 , n35563 );
    not g23583 ( n18566 , n181 );
    nor g23584 ( n29573 , n17568 , n14991 );
    xnor g23585 ( n27949 , n24086 , n4288 );
    or g23586 ( n33608 , n4113 , n9675 );
    nor g23587 ( n29157 , n30817 , n32379 );
    or g23588 ( n30831 , n13505 , n5260 );
    not g23589 ( n35237 , n28404 );
    or g23590 ( n11695 , n2515 , n25940 );
    or g23591 ( n22981 , n35927 , n15503 );
    and g23592 ( n33011 , n19725 , n1930 );
    or g23593 ( n30104 , n4960 , n25730 );
    and g23594 ( n34092 , n13694 , n22140 );
    xnor g23595 ( n13979 , n34555 , n29713 );
    xnor g23596 ( n3887 , n2521 , n31289 );
    or g23597 ( n23844 , n34156 , n17111 );
    or g23598 ( n2146 , n26035 , n544 );
    and g23599 ( n33556 , n16162 , n1889 );
    and g23600 ( n16898 , n29339 , n23094 );
    and g23601 ( n4857 , n17342 , n9186 );
    or g23602 ( n23860 , n1180 , n29953 );
    xnor g23603 ( n31722 , n18652 , n16135 );
    and g23604 ( n20758 , n22083 , n32892 );
    nor g23605 ( n1126 , n31799 , n32625 );
    nor g23606 ( n34840 , n27226 , n20920 );
    and g23607 ( n8039 , n9262 , n16726 );
    or g23608 ( n20686 , n10894 , n34867 );
    and g23609 ( n4030 , n12785 , n31618 );
    not g23610 ( n8869 , n28539 );
    nor g23611 ( n13073 , n27753 , n6950 );
    and g23612 ( n7318 , n16679 , n21199 );
    or g23613 ( n13988 , n1617 , n2198 );
    or g23614 ( n5030 , n11617 , n27447 );
    and g23615 ( n16048 , n6734 , n4511 );
    or g23616 ( n11175 , n28572 , n16919 );
    not g23617 ( n33372 , n32458 );
    nor g23618 ( n27490 , n11448 , n8075 );
    xnor g23619 ( n5999 , n28195 , n27330 );
    or g23620 ( n2642 , n11188 , n1511 );
    not g23621 ( n26698 , n30742 );
    or g23622 ( n30533 , n22291 , n5044 );
    nor g23623 ( n6294 , n3946 , n18675 );
    or g23624 ( n6641 , n24763 , n18803 );
    or g23625 ( n13682 , n1272 , n12602 );
    or g23626 ( n5862 , n31258 , n20948 );
    or g23627 ( n15701 , n34761 , n443 );
    or g23628 ( n4341 , n9793 , n6463 );
    not g23629 ( n17557 , n19984 );
    or g23630 ( n4171 , n19656 , n20797 );
    xnor g23631 ( n29140 , n6403 , n27809 );
    nor g23632 ( n20189 , n8119 , n9928 );
    xnor g23633 ( n33559 , n24447 , n30825 );
    xnor g23634 ( n9145 , n9273 , n11046 );
    nor g23635 ( n8820 , n4878 , n13082 );
    or g23636 ( n587 , n2717 , n28323 );
    or g23637 ( n18616 , n7380 , n14918 );
    or g23638 ( n14590 , n5287 , n8980 );
    or g23639 ( n20799 , n3191 , n11712 );
    not g23640 ( n3452 , n3205 );
    and g23641 ( n10171 , n15440 , n8843 );
    xnor g23642 ( n3287 , n3327 , n31799 );
    or g23643 ( n12625 , n6851 , n14636 );
    or g23644 ( n2463 , n8348 , n3694 );
    or g23645 ( n16405 , n32029 , n18811 );
    xnor g23646 ( n1359 , n1191 , n12703 );
    not g23647 ( n35437 , n12042 );
    or g23648 ( n31111 , n830 , n26312 );
    xnor g23649 ( n13366 , n10563 , n1950 );
    or g23650 ( n20113 , n29080 , n24025 );
    or g23651 ( n24588 , n18674 , n11518 );
    or g23652 ( n21706 , n32206 , n19807 );
    and g23653 ( n15753 , n15513 , n19536 );
    not g23654 ( n15645 , n2029 );
    and g23655 ( n34154 , n28555 , n3330 );
    or g23656 ( n23102 , n30635 , n4303 );
    or g23657 ( n34336 , n11854 , n11518 );
    xnor g23658 ( n11466 , n22290 , n26685 );
    xnor g23659 ( n32925 , n1453 , n10383 );
    xor g23660 ( n15605 , n31000 , n34086 );
    and g23661 ( n4179 , n15798 , n14262 );
    or g23662 ( n10637 , n35214 , n12618 );
    and g23663 ( n610 , n31119 , n5219 );
    xnor g23664 ( n16708 , n35028 , n15886 );
    or g23665 ( n35594 , n31215 , n26407 );
    nor g23666 ( n20201 , n2477 , n5138 );
    or g23667 ( n18044 , n3205 , n31072 );
    or g23668 ( n25559 , n14865 , n10336 );
    and g23669 ( n12351 , n31316 , n7070 );
    nor g23670 ( n6161 , n34462 , n15256 );
    xnor g23671 ( n1150 , n6054 , n1941 );
    nor g23672 ( n13209 , n25602 , n10809 );
    and g23673 ( n11744 , n34932 , n7749 );
    or g23674 ( n27001 , n4960 , n25740 );
    or g23675 ( n24694 , n19742 , n14164 );
    and g23676 ( n2813 , n4019 , n18577 );
    or g23677 ( n33342 , n10283 , n31611 );
    and g23678 ( n10164 , n22804 , n6483 );
    and g23679 ( n14025 , n23392 , n24532 );
    or g23680 ( n14515 , n11523 , n20300 );
    xnor g23681 ( n16836 , n28610 , n19551 );
    or g23682 ( n21943 , n14613 , n2119 );
    xnor g23683 ( n22366 , n9032 , n24013 );
    or g23684 ( n21377 , n15463 , n24333 );
    or g23685 ( n3973 , n20506 , n13664 );
    or g23686 ( n26583 , n9836 , n16762 );
    nor g23687 ( n24021 , n11190 , n19286 );
    or g23688 ( n27873 , n33422 , n31514 );
    or g23689 ( n29590 , n27983 , n11258 );
    or g23690 ( n29462 , n35550 , n32270 );
    xnor g23691 ( n28831 , n15574 , n28355 );
    or g23692 ( n22778 , n11455 , n16794 );
    xnor g23693 ( n8400 , n2263 , n29873 );
    or g23694 ( n7575 , n1057 , n14706 );
    not g23695 ( n13301 , n26112 );
    xnor g23696 ( n24186 , n25476 , n4430 );
    or g23697 ( n27772 , n5473 , n4172 );
    or g23698 ( n9727 , n29248 , n30292 );
    or g23699 ( n14291 , n25003 , n7025 );
    nor g23700 ( n17172 , n1950 , n6115 );
    or g23701 ( n14017 , n34196 , n15339 );
    and g23702 ( n1903 , n35906 , n16144 );
    xnor g23703 ( n3376 , n17499 , n9789 );
    and g23704 ( n14681 , n19149 , n13044 );
    or g23705 ( n22532 , n14440 , n31150 );
    or g23706 ( n30194 , n10561 , n17243 );
    and g23707 ( n19991 , n2659 , n1818 );
    nor g23708 ( n30771 , n30141 , n11234 );
    and g23709 ( n14536 , n34906 , n9035 );
    or g23710 ( n23002 , n24218 , n33435 );
    and g23711 ( n12299 , n11075 , n20634 );
    or g23712 ( n14569 , n25174 , n32466 );
    xnor g23713 ( n3299 , n35259 , n35927 );
    or g23714 ( n10137 , n16922 , n33006 );
    and g23715 ( n35072 , n15613 , n21125 );
    or g23716 ( n12957 , n4787 , n16457 );
    and g23717 ( n8606 , n19389 , n6659 );
    or g23718 ( n21422 , n24603 , n10277 );
    xnor g23719 ( n8579 , n22676 , n1950 );
    and g23720 ( n25817 , n30359 , n33534 );
    or g23721 ( n9283 , n31559 , n35432 );
    xnor g23722 ( n11971 , n12820 , n4939 );
    xnor g23723 ( n25581 , n942 , n31116 );
    or g23724 ( n26904 , n6468 , n9915 );
    not g23725 ( n17368 , n134 );
    or g23726 ( n22162 , n4967 , n34832 );
    and g23727 ( n4649 , n20118 , n6060 );
    or g23728 ( n20750 , n9789 , n16595 );
    nor g23729 ( n7537 , n8443 , n4161 );
    or g23730 ( n2184 , n22159 , n26365 );
    or g23731 ( n11541 , n23993 , n11205 );
    xnor g23732 ( n35613 , n4583 , n8442 );
    and g23733 ( n7784 , n17142 , n31037 );
    and g23734 ( n30853 , n4946 , n22309 );
    or g23735 ( n16318 , n33812 , n1511 );
    or g23736 ( n32121 , n12151 , n2730 );
    not g23737 ( n20930 , n9802 );
    and g23738 ( n10683 , n9728 , n34409 );
    or g23739 ( n30653 , n1829 , n28191 );
    or g23740 ( n11887 , n22542 , n21145 );
    xnor g23741 ( n19229 , n18130 , n7540 );
    or g23742 ( n8477 , n20326 , n31094 );
    xnor g23743 ( n11051 , n27713 , n10908 );
    or g23744 ( n17935 , n29549 , n7892 );
    or g23745 ( n33421 , n1950 , n31999 );
    or g23746 ( n9464 , n22117 , n13306 );
    or g23747 ( n2238 , n22264 , n25567 );
    and g23748 ( n16751 , n27014 , n1778 );
    xnor g23749 ( n5353 , n21611 , n32857 );
    not g23750 ( n13071 , n34269 );
    not g23751 ( n23894 , n27672 );
    and g23752 ( n6568 , n2392 , n29655 );
    xnor g23753 ( n20293 , n10311 , n9793 );
    nor g23754 ( n25126 , n32715 , n4284 );
    not g23755 ( n23355 , n4878 );
    or g23756 ( n20421 , n28869 , n20840 );
    not g23757 ( n14721 , n20316 );
    or g23758 ( n25681 , n520 , n7553 );
    not g23759 ( n26594 , n22980 );
    xnor g23760 ( n6290 , n7029 , n13452 );
    and g23761 ( n8668 , n7905 , n841 );
    xnor g23762 ( n29364 , n27696 , n31544 );
    or g23763 ( n13110 , n877 , n4363 );
    xnor g23764 ( n18983 , n13344 , n5067 );
    or g23765 ( n24092 , n25595 , n6374 );
    or g23766 ( n16509 , n20058 , n2444 );
    not g23767 ( n34045 , n17305 );
    and g23768 ( n16232 , n29072 , n3554 );
    and g23769 ( n23420 , n7440 , n18390 );
    xnor g23770 ( n35704 , n35128 , n4962 );
    not g23771 ( n8429 , n22980 );
    or g23772 ( n9070 , n5067 , n13344 );
    or g23773 ( n30267 , n980 , n19084 );
    or g23774 ( n11303 , n16857 , n5019 );
    or g23775 ( n13614 , n27629 , n28837 );
    or g23776 ( n15633 , n25189 , n17962 );
    or g23777 ( n15471 , n15114 , n585 );
    and g23778 ( n25489 , n6608 , n6087 );
    and g23779 ( n25088 , n2257 , n18185 );
    and g23780 ( n3835 , n23012 , n14404 );
    or g23781 ( n21284 , n23182 , n29334 );
    xnor g23782 ( n23079 , n25374 , n15911 );
    xnor g23783 ( n24105 , n9946 , n28950 );
    and g23784 ( n19790 , n30996 , n4229 );
    not g23785 ( n3486 , n11596 );
    xnor g23786 ( n20885 , n35284 , n8520 );
    and g23787 ( n12499 , n25768 , n5774 );
    xnor g23788 ( n12769 , n31387 , n20141 );
    or g23789 ( n27363 , n10022 , n3026 );
    nor g23790 ( n28425 , n9789 , n22479 );
    or g23791 ( n34685 , n34398 , n2524 );
    or g23792 ( n34479 , n26537 , n11170 );
    or g23793 ( n26285 , n4960 , n5118 );
    xnor g23794 ( n31827 , n12387 , n12470 );
    nor g23795 ( n22883 , n15886 , n15906 );
    and g23796 ( n33908 , n22840 , n14622 );
    or g23797 ( n25833 , n27065 , n27693 );
    or g23798 ( n10692 , n16829 , n17068 );
    and g23799 ( n27831 , n32104 , n2110 );
    or g23800 ( n14260 , n9658 , n34810 );
    buf g23801 ( n15344 , n32096 );
    or g23802 ( n3944 , n30828 , n12428 );
    or g23803 ( n3836 , n35520 , n26002 );
    xnor g23804 ( n1389 , n24272 , n2251 );
    or g23805 ( n27348 , n23424 , n4363 );
    and g23806 ( n8465 , n25407 , n33672 );
    not g23807 ( n7437 , n31355 );
    or g23808 ( n662 , n29497 , n10140 );
    or g23809 ( n29107 , n17467 , n25469 );
    or g23810 ( n22278 , n566 , n8392 );
    or g23811 ( n15849 , n25389 , n8924 );
    xnor g23812 ( n12885 , n29821 , n15886 );
    and g23813 ( n436 , n10796 , n25556 );
    or g23814 ( n32097 , n10624 , n23921 );
    or g23815 ( n35597 , n10751 , n27580 );
    xnor g23816 ( n26633 , n14418 , n16620 );
    or g23817 ( n21117 , n28598 , n6950 );
    nor g23818 ( n35619 , n10454 , n13755 );
    or g23819 ( n31037 , n1950 , n29081 );
    xnor g23820 ( n12946 , n3543 , n24695 );
    xnor g23821 ( n2367 , n10528 , n9793 );
    nor g23822 ( n27336 , n10894 , n29549 );
    xnor g23823 ( n26724 , n20129 , n7507 );
    xnor g23824 ( n18466 , n27245 , n3636 );
    and g23825 ( n13285 , n17344 , n4962 );
    or g23826 ( n35532 , n26188 , n2894 );
    or g23827 ( n19318 , n14698 , n2518 );
    xnor g23828 ( n21360 , n29427 , n5397 );
    nor g23829 ( n32664 , n32095 , n987 );
    and g23830 ( n18334 , n11687 , n16354 );
    or g23831 ( n2482 , n14728 , n30646 );
    xnor g23832 ( n22745 , n18862 , n32095 );
    or g23833 ( n28327 , n27521 , n27735 );
    and g23834 ( n20906 , n29113 , n5831 );
    xnor g23835 ( n31172 , n27540 , n1484 );
    or g23836 ( n22470 , n7540 , n20338 );
    or g23837 ( n35551 , n29201 , n13402 );
    xnor g23838 ( n21888 , n28047 , n25530 );
    xnor g23839 ( n18313 , n22755 , n16622 );
    not g23840 ( n7251 , n13943 );
    xnor g23841 ( n10494 , n14277 , n33053 );
    xnor g23842 ( n110 , n1119 , n32584 );
    and g23843 ( n27693 , n24466 , n33789 );
    not g23844 ( n31583 , n8341 );
    or g23845 ( n29817 , n31289 , n2610 );
    and g23846 ( n19133 , n3120 , n32987 );
    xnor g23847 ( n33321 , n32239 , n27124 );
    xnor g23848 ( n28562 , n5867 , n35200 );
    and g23849 ( n30024 , n23580 , n14989 );
    nor g23850 ( n2963 , n32095 , n24842 );
    xnor g23851 ( n8452 , n13529 , n16620 );
    or g23852 ( n32462 , n9658 , n23608 );
    or g23853 ( n18998 , n10391 , n33983 );
    nor g23854 ( n10039 , n2835 , n29203 );
    or g23855 ( n28085 , n26234 , n12250 );
    and g23856 ( n28571 , n15015 , n13697 );
    xnor g23857 ( n25416 , n21928 , n4288 );
    xnor g23858 ( n1412 , n3897 , n10894 );
    nor g23859 ( n12029 , n16620 , n11002 );
    xnor g23860 ( n10697 , n10884 , n545 );
    nor g23861 ( n10754 , n9789 , n29983 );
    and g23862 ( n1845 , n35805 , n6871 );
    and g23863 ( n32 , n30324 , n19640 );
    and g23864 ( n8024 , n30079 , n32021 );
    nor g23865 ( n21823 , n29713 , n8487 );
    nor g23866 ( n8832 , n13226 , n12332 );
    and g23867 ( n781 , n12810 , n29244 );
    or g23868 ( n13401 , n3686 , n24356 );
    and g23869 ( n19628 , n8917 , n5270 );
    or g23870 ( n2805 , n16083 , n1397 );
    xnor g23871 ( n26475 , n7612 , n25658 );
    or g23872 ( n21476 , n17356 , n2117 );
    xnor g23873 ( n31164 , n22554 , n21163 );
    xnor g23874 ( n22006 , n8074 , n27705 );
    not g23875 ( n8100 , n23701 );
    and g23876 ( n30049 , n26905 , n34659 );
    or g23877 ( n6057 , n1916 , n12791 );
    xnor g23878 ( n1695 , n18106 , n19551 );
    or g23879 ( n1967 , n24361 , n29626 );
    or g23880 ( n23814 , n6591 , n15538 );
    nor g23881 ( n20613 , n10310 , n12913 );
    or g23882 ( n2699 , n27226 , n23312 );
    and g23883 ( n6779 , n1988 , n2449 );
    or g23884 ( n21633 , n31414 , n19612 );
    and g23885 ( n7618 , n9377 , n26727 );
    or g23886 ( n7114 , n18051 , n13499 );
    or g23887 ( n31259 , n11382 , n26292 );
    not g23888 ( n15688 , n19984 );
    xnor g23889 ( n29851 , n31203 , n31559 );
    and g23890 ( n4554 , n14930 , n30760 );
    and g23891 ( n7966 , n14573 , n35887 );
    and g23892 ( n7934 , n22915 , n2402 );
    not g23893 ( n13198 , n5339 );
    and g23894 ( n26615 , n5442 , n12587 );
    nor g23895 ( n19040 , n35927 , n12385 );
    xnor g23896 ( n5506 , n12984 , n1351 );
    or g23897 ( n9844 , n24371 , n8344 );
    xnor g23898 ( n10675 , n35856 , n2494 );
    and g23899 ( n25226 , n22319 , n18984 );
    and g23900 ( n30772 , n10033 , n35679 );
    xnor g23901 ( n2376 , n9992 , n31835 );
    xnor g23902 ( n29452 , n3686 , n34369 );
    or g23903 ( n23084 , n10829 , n27053 );
    xnor g23904 ( n8533 , n29752 , n33606 );
    or g23905 ( n31698 , n30742 , n25664 );
    xnor g23906 ( n16178 , n20536 , n32215 );
    or g23907 ( n11494 , n22222 , n19464 );
    xnor g23908 ( n696 , n11004 , n10463 );
    or g23909 ( n32496 , n1113 , n23187 );
    or g23910 ( n7625 , n30553 , n1229 );
    or g23911 ( n33637 , n6790 , n5868 );
    or g23912 ( n11957 , n32827 , n25592 );
    or g23913 ( n24174 , n24589 , n34472 );
    xnor g23914 ( n1590 , n14656 , n4014 );
    and g23915 ( n13230 , n12615 , n10720 );
    and g23916 ( n32038 , n3335 , n28400 );
    and g23917 ( n33766 , n9242 , n20046 );
    or g23918 ( n1954 , n12466 , n23626 );
    or g23919 ( n22710 , n30742 , n4377 );
    or g23920 ( n22135 , n1497 , n12660 );
    not g23921 ( n10066 , n25776 );
    xnor g23922 ( n24681 , n19883 , n35317 );
    or g23923 ( n27814 , n32058 , n26112 );
    or g23924 ( n14010 , n1406 , n527 );
    and g23925 ( n27471 , n19416 , n30755 );
    xnor g23926 ( n12582 , n27985 , n9793 );
    not g23927 ( n27760 , n16620 );
    or g23928 ( n25286 , n5160 , n2104 );
    and g23929 ( n13008 , n23573 , n29875 );
    xnor g23930 ( n35929 , n10324 , n31289 );
    nor g23931 ( n19526 , n31215 , n21106 );
    and g23932 ( n14251 , n33885 , n4288 );
    or g23933 ( n22985 , n12217 , n5168 );
    xnor g23934 ( n13277 , n12320 , n8432 );
    xnor g23935 ( n8528 , n16387 , n32857 );
    or g23936 ( n22176 , n26087 , n13808 );
    or g23937 ( n30894 , n6884 , n30851 );
    xnor g23938 ( n35867 , n486 , n23438 );
    nor g23939 ( n28963 , n29839 , n18165 );
    or g23940 ( n13606 , n13609 , n31549 );
    or g23941 ( n9948 , n4288 , n6753 );
    xnor g23942 ( n34969 , n3780 , n25602 );
    nor g23943 ( n13400 , n28941 , n1176 );
    not g23944 ( n29097 , n22980 );
    nor g23945 ( n13247 , n13790 , n28246 );
    and g23946 ( n13924 , n7211 , n20179 );
    and g23947 ( n12436 , n35677 , n7619 );
    xnor g23948 ( n6707 , n10218 , n11071 );
    and g23949 ( n33049 , n13182 , n22250 );
    and g23950 ( n22261 , n11688 , n20655 );
    xnor g23951 ( n141 , n11492 , n18005 );
    and g23952 ( n29083 , n7681 , n1669 );
    nor g23953 ( n31920 , n27436 , n13318 );
    not g23954 ( n17692 , n16376 );
    xnor g23955 ( n7299 , n182 , n29066 );
    or g23956 ( n886 , n15886 , n3835 );
    xnor g23957 ( n20694 , n7441 , n17126 );
    not g23958 ( n18502 , n9568 );
    or g23959 ( n31769 , n4288 , n7577 );
    or g23960 ( n32756 , n6883 , n28034 );
    or g23961 ( n14522 , n28651 , n28837 );
    and g23962 ( n4642 , n11941 , n11746 );
    not g23963 ( n20408 , n23923 );
    or g23964 ( n8439 , n31305 , n20013 );
    or g23965 ( n19393 , n4923 , n16757 );
    xnor g23966 ( n10102 , n3138 , n24371 );
    and g23967 ( n9838 , n35206 , n21375 );
    buf g23968 ( n7417 , n24581 );
    or g23969 ( n29954 , n24926 , n25580 );
    and g23970 ( n30386 , n14237 , n35252 );
    or g23971 ( n17787 , n12866 , n30725 );
    nor g23972 ( n4971 , n15464 , n10545 );
    and g23973 ( n4545 , n14580 , n14510 );
    or g23974 ( n20370 , n4962 , n18978 );
    xnor g23975 ( n236 , n26773 , n25602 );
    or g23976 ( n15763 , n27722 , n20797 );
    or g23977 ( n34868 , n29622 , n10634 );
    nor g23978 ( n32179 , n9658 , n935 );
    not g23979 ( n18931 , n34625 );
    and g23980 ( n3143 , n32575 , n31856 );
    xnor g23981 ( n30312 , n16398 , n6056 );
    xnor g23982 ( n99 , n36041 , n6139 );
    or g23983 ( n19356 , n15856 , n32828 );
    or g23984 ( n21609 , n19884 , n6178 );
    xnor g23985 ( n10214 , n34590 , n32095 );
    xnor g23986 ( n19414 , n22568 , n34809 );
    xnor g23987 ( n30818 , n33932 , n18676 );
    or g23988 ( n32381 , n21428 , n36000 );
    nor g23989 ( n23547 , n19551 , n28608 );
    or g23990 ( n22306 , n8432 , n12320 );
    or g23991 ( n30629 , n7243 , n14504 );
    xnor g23992 ( n23406 , n6180 , n12774 );
    or g23993 ( n26289 , n9391 , n26023 );
    buf g23994 ( n9951 , n2609 );
    buf g23995 ( n21977 , n7787 );
    or g23996 ( n35790 , n4878 , n22227 );
    xnor g23997 ( n34701 , n35180 , n23349 );
    or g23998 ( n21734 , n22228 , n21210 );
    or g23999 ( n21549 , n10160 , n6288 );
    or g24000 ( n9778 , n2931 , n26931 );
    not g24001 ( n27262 , n11996 );
    xnor g24002 ( n15594 , n34268 , n12302 );
    or g24003 ( n16165 , n9793 , n23883 );
    nor g24004 ( n31747 , n32857 , n25536 );
    and g24005 ( n7775 , n26111 , n29755 );
    not g24006 ( n26902 , n33429 );
    not g24007 ( n34549 , n33805 );
    xnor g24008 ( n16316 , n2618 , n8959 );
    xnor g24009 ( n29722 , n29497 , n32075 );
    or g24010 ( n23973 , n35328 , n3685 );
    or g24011 ( n1241 , n22303 , n9731 );
    or g24012 ( n33406 , n31084 , n31147 );
    xnor g24013 ( n17284 , n14440 , n31150 );
    or g24014 ( n3053 , n3918 , n6950 );
    nor g24015 ( n11023 , n22508 , n578 );
    or g24016 ( n32763 , n28347 , n4235 );
    or g24017 ( n35711 , n13577 , n10872 );
    and g24018 ( n3763 , n35264 , n15218 );
    and g24019 ( n29614 , n27187 , n22639 );
    or g24020 ( n11054 , n6409 , n15496 );
    or g24021 ( n24236 , n20592 , n20601 );
    or g24022 ( n27826 , n3574 , n23165 );
    or g24023 ( n5414 , n31272 , n7380 );
    and g24024 ( n28985 , n15013 , n9392 );
    xnor g24025 ( n29733 , n11055 , n7540 );
    nor g24026 ( n8152 , n13469 , n6017 );
    not g24027 ( n4950 , n11287 );
    or g24028 ( n4148 , n2794 , n19464 );
    not g24029 ( n19086 , n22980 );
    and g24030 ( n12125 , n23160 , n24467 );
    xnor g24031 ( n19879 , n30494 , n809 );
    buf g24032 ( n15145 , n17111 );
    or g24033 ( n26533 , n7901 , n3858 );
    and g24034 ( n19449 , n10842 , n12567 );
    or g24035 ( n2638 , n21096 , n5279 );
    or g24036 ( n20683 , n11178 , n35064 );
    and g24037 ( n30605 , n35185 , n15964 );
    not g24038 ( n1904 , n28044 );
    not g24039 ( n25694 , n6288 );
    or g24040 ( n22644 , n3946 , n6579 );
    or g24041 ( n13178 , n19551 , n12133 );
    or g24042 ( n26355 , n32239 , n16259 );
    nor g24043 ( n27795 , n30742 , n24697 );
    not g24044 ( n33761 , n9361 );
    and g24045 ( n683 , n12435 , n18191 );
    and g24046 ( n16781 , n10963 , n28279 );
    xnor g24047 ( n24020 , n34918 , n7543 );
    and g24048 ( n29425 , n33137 , n8329 );
    buf g24049 ( n28064 , n17184 );
    and g24050 ( n20589 , n1442 , n12969 );
    not g24051 ( n32491 , n8920 );
    or g24052 ( n27115 , n4878 , n19589 );
    or g24053 ( n29674 , n5687 , n1158 );
    not g24054 ( n14275 , n17725 );
    nor g24055 ( n13345 , n35927 , n22632 );
    xnor g24056 ( n22598 , n30025 , n4288 );
    or g24057 ( n15640 , n2356 , n19125 );
    xnor g24058 ( n1551 , n7621 , n3222 );
    or g24059 ( n4883 , n16654 , n9520 );
    or g24060 ( n32150 , n24969 , n30260 );
    xnor g24061 ( n18709 , n18668 , n4288 );
    and g24062 ( n23759 , n14163 , n7020 );
    xnor g24063 ( n28388 , n20683 , n19551 );
    nor g24064 ( n22715 , n29713 , n17278 );
    or g24065 ( n34047 , n19551 , n11442 );
    xnor g24066 ( n27269 , n18383 , n11954 );
    or g24067 ( n801 , n15890 , n15256 );
    xnor g24068 ( n34138 , n9359 , n4428 );
    and g24069 ( n22968 , n2173 , n29091 );
    or g24070 ( n16043 , n5335 , n18498 );
    or g24071 ( n33692 , n6877 , n23921 );
    or g24072 ( n27255 , n32580 , n17125 );
    or g24073 ( n17051 , n35303 , n34537 );
    or g24074 ( n19935 , n25121 , n31514 );
    or g24075 ( n21664 , n33925 , n26482 );
    xnor g24076 ( n24859 , n17475 , n5149 );
    xnor g24077 ( n825 , n26581 , n9793 );
    or g24078 ( n3450 , n29839 , n1518 );
    and g24079 ( n4188 , n88 , n35893 );
    xnor g24080 ( n27326 , n21978 , n5335 );
    or g24081 ( n25628 , n2394 , n11977 );
    nor g24082 ( n7503 , n16922 , n20418 );
    or g24083 ( n27651 , n28558 , n18881 );
    nor g24084 ( n34644 , n29561 , n26856 );
    and g24085 ( n2351 , n26560 , n12168 );
    and g24086 ( n33712 , n35433 , n23014 );
    nor g24087 ( n21230 , n4878 , n4679 );
    and g24088 ( n1520 , n18019 , n21548 );
    or g24089 ( n21125 , n5287 , n2714 );
    and g24090 ( n20712 , n4562 , n26771 );
    or g24091 ( n22536 , n24264 , n5779 );
    or g24092 ( n19655 , n4678 , n14486 );
    or g24093 ( n356 , n12226 , n23090 );
    xnor g24094 ( n2236 , n5313 , n4758 );
    xnor g24095 ( n17157 , n35694 , n16922 );
    and g24096 ( n33902 , n3442 , n24143 );
    nor g24097 ( n19543 , n13670 , n15486 );
    or g24098 ( n31518 , n7252 , n31055 );
    or g24099 ( n28604 , n30380 , n344 );
    or g24100 ( n3659 , n33978 , n5956 );
    xnor g24101 ( n11609 , n33374 , n18280 );
    or g24102 ( n23876 , n17007 , n10264 );
    xnor g24103 ( n21662 , n26719 , n8805 );
    xnor g24104 ( n10108 , n10174 , n11252 );
    and g24105 ( n20030 , n16643 , n631 );
    or g24106 ( n33021 , n28272 , n27973 );
    xnor g24107 ( n17521 , n19908 , n35313 );
    and g24108 ( n19521 , n23433 , n3001 );
    or g24109 ( n5256 , n11751 , n32576 );
    or g24110 ( n21206 , n28527 , n4081 );
    and g24111 ( n21339 , n18008 , n2982 );
    and g24112 ( n5663 , n12709 , n31698 );
    xnor g24113 ( n25426 , n3769 , n19984 );
    xnor g24114 ( n34276 , n26716 , n3420 );
    not g24115 ( n12725 , n14627 );
    and g24116 ( n30577 , n31286 , n13240 );
    or g24117 ( n1184 , n5648 , n13664 );
    and g24118 ( n10269 , n23695 , n23885 );
    or g24119 ( n13627 , n29575 , n1810 );
    or g24120 ( n10539 , n1753 , n30478 );
    xnor g24121 ( n35747 , n23759 , n31272 );
    or g24122 ( n14186 , n27503 , n28330 );
    xnor g24123 ( n18456 , n9565 , n29713 );
    or g24124 ( n9787 , n24360 , n20797 );
    xnor g24125 ( n31415 , n29557 , n22291 );
    nor g24126 ( n34764 , n19837 , n9915 );
    or g24127 ( n22342 , n20536 , n32215 );
    and g24128 ( n8311 , n25967 , n27918 );
    not g24129 ( n11922 , n31457 );
    and g24130 ( n1228 , n149 , n8602 );
    or g24131 ( n10740 , n2148 , n16457 );
    and g24132 ( n5441 , n3944 , n16055 );
    nor g24133 ( n1322 , n14221 , n17029 );
    nor g24134 ( n28974 , n32671 , n21044 );
    nor g24135 ( n7591 , n1950 , n35553 );
    and g24136 ( n20846 , n23866 , n19529 );
    or g24137 ( n22321 , n24750 , n5967 );
    xnor g24138 ( n4147 , n24281 , n8432 );
    or g24139 ( n15314 , n25644 , n4772 );
    and g24140 ( n12294 , n21936 , n20900 );
    and g24141 ( n24795 , n29815 , n34145 );
    and g24142 ( n34423 , n35634 , n6570 );
    nor g24143 ( n21567 , n17435 , n18115 );
    xnor g24144 ( n22286 , n7762 , n9658 );
    or g24145 ( n32428 , n8432 , n6094 );
    or g24146 ( n20323 , n35204 , n11977 );
    not g24147 ( n20585 , n31851 );
    and g24148 ( n28997 , n17929 , n30793 );
    xnor g24149 ( n21345 , n34355 , n30453 );
    xnor g24150 ( n32934 , n26587 , n189 );
    nor g24151 ( n23077 , n29839 , n24602 );
    or g24152 ( n3442 , n21604 , n908 );
    xnor g24153 ( n29662 , n6015 , n33139 );
    xnor g24154 ( n9271 , n33458 , n34461 );
    or g24155 ( n19539 , n15832 , n35265 );
    or g24156 ( n32237 , n10326 , n25594 );
    xnor g24157 ( n14439 , n27534 , n25174 );
    or g24158 ( n13746 , n1538 , n13305 );
    or g24159 ( n6095 , n14712 , n4454 );
    or g24160 ( n17920 , n17812 , n122 );
    or g24161 ( n34548 , n33360 , n11776 );
    and g24162 ( n17587 , n3973 , n15238 );
    nor g24163 ( n3562 , n35927 , n14929 );
    xnor g24164 ( n31742 , n7296 , n966 );
    and g24165 ( n3327 , n17627 , n35862 );
    or g24166 ( n32628 , n23535 , n30204 );
    not g24167 ( n28705 , n25761 );
    or g24168 ( n13733 , n33716 , n24635 );
    xnor g24169 ( n10366 , n29280 , n27226 );
    xnor g24170 ( n26270 , n31772 , n13767 );
    xnor g24171 ( n14851 , n32234 , n12448 );
    nor g24172 ( n25274 , n19551 , n24777 );
    nor g24173 ( n19045 , n30742 , n25149 );
    or g24174 ( n22816 , n28047 , n25530 );
    or g24175 ( n29405 , n338 , n32618 );
    and g24176 ( n28136 , n10871 , n27346 );
    or g24177 ( n13581 , n10367 , n19464 );
    buf g24178 ( n10454 , n19573 );
    xnor g24179 ( n10352 , n15273 , n36003 );
    or g24180 ( n22666 , n32102 , n27308 );
    nor g24181 ( n10375 , n17568 , n31743 );
    or g24182 ( n28209 , n25968 , n15371 );
    or g24183 ( n32302 , n27885 , n5168 );
    or g24184 ( n9877 , n11433 , n24485 );
    xnor g24185 ( n13676 , n16968 , n14432 );
    buf g24186 ( n34484 , n8666 );
    and g24187 ( n28331 , n31031 , n33675 );
    not g24188 ( n34728 , n15299 );
    xnor g24189 ( n14057 , n19065 , n15826 );
    xnor g24190 ( n25651 , n12266 , n35650 );
    or g24191 ( n28501 , n10540 , n24973 );
    or g24192 ( n17963 , n6400 , n22027 );
    or g24193 ( n34198 , n15626 , n4508 );
    or g24194 ( n8492 , n19360 , n20576 );
    nor g24195 ( n19412 , n34276 , n9921 );
    xnor g24196 ( n26299 , n27090 , n12143 );
    and g24197 ( n35936 , n32397 , n7689 );
    xnor g24198 ( n18762 , n4504 , n13855 );
    and g24199 ( n35504 , n1177 , n26377 );
    xnor g24200 ( n23126 , n11791 , n8154 );
    xnor g24201 ( n35640 , n27994 , n7540 );
    or g24202 ( n11686 , n5749 , n1763 );
    or g24203 ( n3185 , n22879 , n35170 );
    and g24204 ( n34542 , n705 , n1721 );
    or g24205 ( n12749 , n15989 , n20824 );
    or g24206 ( n15225 , n20787 , n28513 );
    or g24207 ( n34031 , n33631 , n10289 );
    xnor g24208 ( n24786 , n3193 , n31128 );
    or g24209 ( n4612 , n4435 , n12128 );
    not g24210 ( n17372 , n22501 );
    xnor g24211 ( n7795 , n2511 , n28536 );
    xnor g24212 ( n24533 , n14532 , n3800 );
    buf g24213 ( n578 , n11773 );
    and g24214 ( n5644 , n28127 , n2349 );
    or g24215 ( n34799 , n24872 , n29897 );
    not g24216 ( n16298 , n5320 );
    nor g24217 ( n7094 , n9789 , n10300 );
    xor g24218 ( n13194 , n27857 , n10748 );
    xnor g24219 ( n20043 , n10199 , n18379 );
    xnor g24220 ( n15065 , n34320 , n4525 );
    and g24221 ( n35425 , n24547 , n856 );
    not g24222 ( n7453 , n18481 );
    nor g24223 ( n6682 , n14595 , n4495 );
    nor g24224 ( n22099 , n15403 , n18593 );
    or g24225 ( n4666 , n12023 , n5663 );
    and g24226 ( n13629 , n14519 , n8220 );
    or g24227 ( n18785 , n32095 , n8778 );
    xnor g24228 ( n23590 , n17713 , n19551 );
    not g24229 ( n3600 , n15886 );
    xnor g24230 ( n28765 , n23721 , n26686 );
    and g24231 ( n9147 , n26228 , n13570 );
    xnor g24232 ( n23428 , n17114 , n22589 );
    or g24233 ( n18813 , n4960 , n3629 );
    or g24234 ( n14384 , n6773 , n30242 );
    or g24235 ( n2603 , n3596 , n4490 );
    and g24236 ( n17601 , n5193 , n12962 );
    or g24237 ( n25049 , n25575 , n7647 );
    or g24238 ( n9156 , n32638 , n17964 );
    or g24239 ( n539 , n18632 , n29592 );
    or g24240 ( n6025 , n27291 , n15464 );
    and g24241 ( n19271 , n10778 , n8303 );
    xnor g24242 ( n33898 , n15449 , n18730 );
    xnor g24243 ( n27249 , n3696 , n35927 );
    xnor g24244 ( n8445 , n19291 , n4878 );
    or g24245 ( n15760 , n5335 , n22370 );
    nor g24246 ( n422 , n27226 , n24713 );
    or g24247 ( n24482 , n3946 , n1015 );
    xnor g24248 ( n13207 , n14165 , n885 );
    and g24249 ( n21019 , n19141 , n27843 );
    xnor g24250 ( n31720 , n24919 , n4288 );
    or g24251 ( n6378 , n15606 , n17964 );
    not g24252 ( n26340 , n1342 );
    xnor g24253 ( n15452 , n27434 , n25174 );
    or g24254 ( n19683 , n26621 , n24710 );
    not g24255 ( n22048 , n34800 );
    or g24256 ( n21784 , n4758 , n10602 );
    or g24257 ( n9127 , n19252 , n14640 );
    nor g24258 ( n22273 , n29713 , n28889 );
    or g24259 ( n21997 , n28877 , n578 );
    and g24260 ( n6415 , n7609 , n4292 );
    or g24261 ( n2499 , n10244 , n32572 );
    or g24262 ( n25446 , n35369 , n23089 );
    xnor g24263 ( n34694 , n1627 , n4288 );
    xnor g24264 ( n9366 , n320 , n22291 );
    xnor g24265 ( n4373 , n5435 , n28262 );
    or g24266 ( n21612 , n15403 , n20211 );
    or g24267 ( n3919 , n12461 , n4334 );
    or g24268 ( n25053 , n25514 , n24333 );
    xnor g24269 ( n9453 , n11997 , n4076 );
    nor g24270 ( n27864 , n32715 , n4857 );
    or g24271 ( n25965 , n9363 , n1001 );
    and g24272 ( n17553 , n184 , n14312 );
    xnor g24273 ( n11956 , n13454 , n1950 );
    or g24274 ( n16274 , n11046 , n2625 );
    xnor g24275 ( n31649 , n32264 , n21291 );
    or g24276 ( n1035 , n10881 , n35820 );
    and g24277 ( n36029 , n23730 , n28372 );
    or g24278 ( n28056 , n8244 , n8392 );
    not g24279 ( n20079 , n9658 );
    and g24280 ( n21234 , n28726 , n16839 );
    xnor g24281 ( n10486 , n12803 , n22291 );
    or g24282 ( n7006 , n17524 , n23187 );
    and g24283 ( n17526 , n25506 , n29057 );
    or g24284 ( n7283 , n7813 , n24025 );
    and g24285 ( n1001 , n35509 , n22406 );
    or g24286 ( n27553 , n28361 , n33034 );
    or g24287 ( n21276 , n8775 , n24653 );
    xnor g24288 ( n19139 , n12172 , n5335 );
    and g24289 ( n6332 , n24594 , n21276 );
    and g24290 ( n14286 , n13115 , n35342 );
    or g24291 ( n23153 , n23849 , n14328 );
    or g24292 ( n14135 , n18318 , n35107 );
    and g24293 ( n11067 , n29915 , n7143 );
    or g24294 ( n3075 , n25604 , n26244 );
    xnor g24295 ( n20245 , n28892 , n30752 );
    or g24296 ( n16592 , n259 , n19952 );
    not g24297 ( n28870 , n11021 );
    or g24298 ( n4931 , n35521 , n22946 );
    or g24299 ( n26788 , n10012 , n20817 );
    xor g24300 ( n18344 , n21219 , n2705 );
    not g24301 ( n21231 , n27226 );
    or g24302 ( n31865 , n9658 , n2998 );
    not g24303 ( n21266 , n4878 );
    nor g24304 ( n28121 , n27156 , n35337 );
    or g24305 ( n27241 , n12191 , n34922 );
    not g24306 ( n20227 , n18224 );
    and g24307 ( n11172 , n16913 , n28391 );
    or g24308 ( n5682 , n27710 , n28064 );
    and g24309 ( n4297 , n23409 , n14044 );
    or g24310 ( n29251 , n30649 , n10872 );
    and g24311 ( n19444 , n25618 , n4747 );
    and g24312 ( n21869 , n33238 , n30358 );
    or g24313 ( n9545 , n27530 , n16797 );
    nor g24314 ( n12660 , n17660 , n2629 );
    nor g24315 ( n28557 , n24371 , n4955 );
    or g24316 ( n31376 , n15340 , n21803 );
    not g24317 ( n3481 , n24371 );
    or g24318 ( n11453 , n27291 , n33327 );
    not g24319 ( n16855 , n3858 );
    or g24320 ( n35353 , n10062 , n34727 );
    and g24321 ( n24024 , n13435 , n30585 );
    or g24322 ( n6739 , n4755 , n19241 );
    not g24323 ( n4430 , n10894 );
    and g24324 ( n13689 , n264 , n31218 );
    or g24325 ( n27059 , n13960 , n25392 );
    xnor g24326 ( n8841 , n27644 , n15499 );
    or g24327 ( n9671 , n23415 , n3842 );
    or g24328 ( n19114 , n12122 , n10656 );
    nor g24329 ( n4056 , n27471 , n23103 );
    xnor g24330 ( n11271 , n10454 , n24024 );
    xnor g24331 ( n24603 , n5412 , n9793 );
    nor g24332 ( n28092 , n22291 , n4668 );
    not g24333 ( n33249 , n24127 );
    not g24334 ( n27886 , n7951 );
    xnor g24335 ( n24159 , n28217 , n27968 );
    or g24336 ( n34078 , n19984 , n1195 );
    or g24337 ( n22375 , n34473 , n7966 );
    or g24338 ( n2166 , n16922 , n1948 );
    and g24339 ( n10075 , n18494 , n13711 );
    nor g24340 ( n14886 , n10404 , n3730 );
    xnor g24341 ( n23789 , n12558 , n12540 );
    xnor g24342 ( n13274 , n34192 , n25602 );
    not g24343 ( n9856 , n14617 );
    or g24344 ( n953 , n7590 , n26214 );
    xnor g24345 ( n20258 , n2982 , n18008 );
    and g24346 ( n22776 , n33294 , n34264 );
    or g24347 ( n31658 , n35927 , n18235 );
    or g24348 ( n24709 , n29839 , n18061 );
    xnor g24349 ( n27721 , n11637 , n6632 );
    or g24350 ( n15023 , n12713 , n5309 );
    or g24351 ( n9166 , n26566 , n3979 );
    nor g24352 ( n9225 , n26942 , n19386 );
    xnor g24353 ( n33190 , n22399 , n95 );
    or g24354 ( n18926 , n19419 , n18163 );
    and g24355 ( n7639 , n8512 , n19242 );
    or g24356 ( n21300 , n5921 , n14918 );
    or g24357 ( n28280 , n1287 , n10872 );
    or g24358 ( n30093 , n21460 , n13337 );
    xnor g24359 ( n8124 , n23169 , n31799 );
    and g24360 ( n22505 , n6464 , n3139 );
    or g24361 ( n13625 , n19859 , n5900 );
    and g24362 ( n26974 , n12600 , n25770 );
    buf g24363 ( n16857 , n9981 );
    xnor g24364 ( n13609 , n27628 , n467 );
    or g24365 ( n23298 , n26938 , n19241 );
    or g24366 ( n31117 , n12087 , n11704 );
    or g24367 ( n30455 , n11697 , n4818 );
    not g24368 ( n17384 , n30742 );
    nor g24369 ( n33156 , n9658 , n24546 );
    or g24370 ( n30770 , n30619 , n25019 );
    not g24371 ( n21853 , n3842 );
    not g24372 ( n6867 , n30998 );
    and g24373 ( n29300 , n30194 , n13864 );
    xnor g24374 ( n8813 , n32643 , n22557 );
    and g24375 ( n5495 , n29773 , n29978 );
    and g24376 ( n34801 , n17282 , n30528 );
    or g24377 ( n8787 , n20176 , n34923 );
    and g24378 ( n18851 , n29414 , n2870 );
    or g24379 ( n23477 , n7507 , n29366 );
    not g24380 ( n8171 , n16725 );
    xnor g24381 ( n13612 , n5981 , n25174 );
    or g24382 ( n30408 , n23597 , n23566 );
    or g24383 ( n15039 , n29910 , n25592 );
    nor g24384 ( n32087 , n31050 , n3800 );
    or g24385 ( n21051 , n16922 , n8552 );
    xnor g24386 ( n23913 , n26579 , n3575 );
    nor g24387 ( n6043 , n31289 , n9534 );
    or g24388 ( n5605 , n19923 , n492 );
    or g24389 ( n32927 , n23583 , n15921 );
    or g24390 ( n10991 , n32293 , n27695 );
    or g24391 ( n9745 , n2008 , n11665 );
    and g24392 ( n31989 , n5326 , n17012 );
    and g24393 ( n21981 , n15031 , n6803 );
    xnor g24394 ( n9808 , n31126 , n31799 );
    or g24395 ( n14149 , n28486 , n25761 );
    and g24396 ( n35150 , n23873 , n2541 );
    and g24397 ( n18099 , n22410 , n26276 );
    xnor g24398 ( n28176 , n34021 , n20675 );
    and g24399 ( n6572 , n9050 , n32221 );
    nor g24400 ( n12010 , n26827 , n22874 );
    and g24401 ( n35521 , n27097 , n24507 );
    and g24402 ( n9140 , n11328 , n8561 );
    xnor g24403 ( n23665 , n23922 , n6089 );
    and g24404 ( n5379 , n33500 , n1967 );
    or g24405 ( n33313 , n10917 , n12791 );
    and g24406 ( n28255 , n19967 , n14095 );
    not g24407 ( n4999 , n18404 );
    xnor g24408 ( n4433 , n31414 , n19612 );
    nor g24409 ( n3572 , n5287 , n767 );
    xnor g24410 ( n4140 , n2921 , n30095 );
    or g24411 ( n30843 , n31844 , n4952 );
    not g24412 ( n18358 , n22241 );
    xnor g24413 ( n6092 , n10766 , n23808 );
    and g24414 ( n34001 , n15126 , n22093 );
    xnor g24415 ( n7797 , n4916 , n19551 );
    xnor g24416 ( n4015 , n33408 , n404 );
    and g24417 ( n35383 , n25559 , n4696 );
    or g24418 ( n18200 , n35199 , n5151 );
    xnor g24419 ( n3675 , n30107 , n21459 );
    xnor g24420 ( n22974 , n32479 , n31654 );
    xnor g24421 ( n4063 , n28130 , n14000 );
    or g24422 ( n32667 , n34069 , n30812 );
    xnor g24423 ( n23085 , n26237 , n23549 );
    or g24424 ( n2 , n26956 , n27960 );
    xnor g24425 ( n11257 , n2998 , n9658 );
    and g24426 ( n28827 , n5293 , n3181 );
    and g24427 ( n983 , n32709 , n27499 );
    and g24428 ( n29602 , n25360 , n34496 );
    not g24429 ( n19830 , n3041 );
    and g24430 ( n11484 , n26 , n4063 );
    and g24431 ( n14845 , n5863 , n29022 );
    or g24432 ( n15269 , n28005 , n20427 );
    xnor g24433 ( n14977 , n22261 , n33910 );
    or g24434 ( n26298 , n10888 , n23921 );
    xnor g24435 ( n10951 , n14605 , n17751 );
    xor g24436 ( n16892 , n25434 , n19924 );
    and g24437 ( n7993 , n3787 , n21402 );
    or g24438 ( n34942 , n3657 , n12118 );
    xnor g24439 ( n6422 , n19447 , n15886 );
    and g24440 ( n17998 , n6007 , n16008 );
    and g24441 ( n2061 , n4298 , n13721 );
    or g24442 ( n11217 , n24057 , n6553 );
    xnor g24443 ( n23710 , n7001 , n29633 );
    xor g24444 ( n9014 , n12908 , n10261 );
    and g24445 ( n32293 , n8925 , n21047 );
    xnor g24446 ( n735 , n9980 , n5670 );
    and g24447 ( n6316 , n33616 , n4374 );
    or g24448 ( n28426 , n32715 , n6733 );
    and g24449 ( n6828 , n26311 , n30823 );
    or g24450 ( n17100 , n26069 , n34600 );
    and g24451 ( n34815 , n15458 , n359 );
    or g24452 ( n5744 , n35017 , n23209 );
    nor g24453 ( n27388 , n27562 , n17314 );
    or g24454 ( n5177 , n4288 , n19118 );
    and g24455 ( n9355 , n13032 , n21408 );
    xnor g24456 ( n28708 , n26464 , n20439 );
    or g24457 ( n2675 , n30123 , n6553 );
    nor g24458 ( n12043 , n4878 , n29692 );
    xnor g24459 ( n53 , n19324 , n7639 );
    and g24460 ( n8552 , n5331 , n23682 );
    or g24461 ( n1550 , n12205 , n9601 );
    and g24462 ( n2521 , n9083 , n15562 );
    or g24463 ( n12988 , n4288 , n5052 );
    or g24464 ( n31367 , n3916 , n3072 );
    xnor g24465 ( n32416 , n2370 , n25466 );
    and g24466 ( n345 , n1854 , n5134 );
    nor g24467 ( n33065 , n35927 , n25441 );
    nor g24468 ( n8601 , n18468 , n4508 );
    and g24469 ( n35514 , n2836 , n25399 );
    or g24470 ( n23184 , n5378 , n22717 );
    or g24471 ( n21226 , n16238 , n19079 );
    buf g24472 ( n21644 , n26418 );
    or g24473 ( n12631 , n5287 , n18769 );
    or g24474 ( n4462 , n25074 , n15895 );
    and g24475 ( n17258 , n3233 , n8116 );
    or g24476 ( n7813 , n14174 , n6478 );
    and g24477 ( n3241 , n11080 , n10853 );
    nor g24478 ( n18767 , n14487 , n6017 );
    or g24479 ( n35566 , n35605 , n7417 );
    and g24480 ( n26371 , n7879 , n16428 );
    or g24481 ( n18116 , n15051 , n29872 );
    or g24482 ( n24472 , n32040 , n28189 );
    or g24483 ( n32327 , n1888 , n28804 );
    xnor g24484 ( n16174 , n35300 , n3117 );
    and g24485 ( n24924 , n27508 , n27620 );
    nor g24486 ( n7516 , n28707 , n19446 );
    or g24487 ( n35996 , n2367 , n1840 );
    and g24488 ( n8974 , n16545 , n26636 );
    or g24489 ( n19301 , n17568 , n2230 );
    xnor g24490 ( n19884 , n47 , n12974 );
    xnor g24491 ( n32742 , n13014 , n22438 );
    or g24492 ( n4123 , n4960 , n15295 );
    or g24493 ( n3198 , n14448 , n19968 );
    and g24494 ( n9875 , n7471 , n5737 );
    or g24495 ( n12513 , n28231 , n30826 );
    not g24496 ( n15809 , n2092 );
    and g24497 ( n13451 , n23600 , n349 );
    and g24498 ( n7369 , n7780 , n25091 );
    xnor g24499 ( n29816 , n8685 , n16922 );
    xnor g24500 ( n13660 , n36084 , n29713 );
    and g24501 ( n34142 , n19538 , n6264 );
    xnor g24502 ( n27050 , n913 , n28510 );
    xnor g24503 ( n33635 , n10654 , n8795 );
    xnor g24504 ( n9795 , n21570 , n24118 );
    not g24505 ( n14567 , n21706 );
    and g24506 ( n31796 , n10929 , n26607 );
    and g24507 ( n367 , n17523 , n18350 );
    xnor g24508 ( n27431 , n34578 , n31272 );
    or g24509 ( n12675 , n30742 , n19819 );
    and g24510 ( n22437 , n16401 , n4302 );
    xnor g24511 ( n32392 , n22229 , n31758 );
    xnor g24512 ( n24295 , n30404 , n12828 );
    xnor g24513 ( n8643 , n7741 , n29990 );
    or g24514 ( n7196 , n1412 , n19593 );
    and g24515 ( n35505 , n14892 , n26654 );
    not g24516 ( n27121 , n29839 );
    nor g24517 ( n6324 , n19984 , n3769 );
    or g24518 ( n9484 , n15991 , n2814 );
    and g24519 ( n14619 , n17210 , n17752 );
    xnor g24520 ( n35176 , n1695 , n19836 );
    or g24521 ( n33330 , n9125 , n19732 );
    or g24522 ( n19337 , n33719 , n21970 );
    xnor g24523 ( n28214 , n32350 , n30742 );
    or g24524 ( n27194 , n15456 , n11712 );
    or g24525 ( n5292 , n20452 , n16762 );
    or g24526 ( n2427 , n142 , n12996 );
    or g24527 ( n27061 , n16794 , n763 );
    and g24528 ( n34258 , n24325 , n12539 );
    and g24529 ( n4807 , n18346 , n35569 );
    or g24530 ( n32596 , n30742 , n26424 );
    and g24531 ( n17128 , n34454 , n22752 );
    or g24532 ( n20023 , n9789 , n16752 );
    not g24533 ( n35314 , n4288 );
    nor g24534 ( n14116 , n28343 , n6017 );
    or g24535 ( n6005 , n25664 , n2955 );
    or g24536 ( n10720 , n15464 , n23916 );
    or g24537 ( n31064 , n8627 , n30646 );
    or g24538 ( n8739 , n1356 , n22129 );
    xnor g24539 ( n27318 , n35580 , n31289 );
    or g24540 ( n32510 , n17101 , n15100 );
    or g24541 ( n2337 , n11373 , n35157 );
    or g24542 ( n2324 , n31384 , n26660 );
    and g24543 ( n33338 , n25178 , n7341 );
    or g24544 ( n18023 , n10410 , n2712 );
    or g24545 ( n5790 , n27498 , n1317 );
    or g24546 ( n32459 , n10676 , n30708 );
    xnor g24547 ( n543 , n29862 , n18371 );
    not g24548 ( n10235 , n16620 );
    xnor g24549 ( n16881 , n19413 , n27226 );
    or g24550 ( n22263 , n11002 , n11977 );
    not g24551 ( n34369 , n4878 );
    and g24552 ( n3162 , n34140 , n9059 );
    nor g24553 ( n31440 , n15886 , n7741 );
    or g24554 ( n22573 , n35059 , n11850 );
    xnor g24555 ( n26678 , n16240 , n29839 );
    xnor g24556 ( n32957 , n19948 , n19013 );
    and g24557 ( n24934 , n19891 , n3617 );
    and g24558 ( n14405 , n20703 , n28577 );
    nor g24559 ( n4790 , n33621 , n20379 );
    or g24560 ( n22011 , n33108 , n3188 );
    xnor g24561 ( n25552 , n23164 , n4138 );
    or g24562 ( n28528 , n33082 , n34600 );
    or g24563 ( n12531 , n25441 , n28574 );
    not g24564 ( n35834 , n22200 );
    or g24565 ( n375 , n23604 , n16219 );
    and g24566 ( n14029 , n4699 , n19853 );
    or g24567 ( n10871 , n28653 , n31930 );
    or g24568 ( n24918 , n18313 , n4478 );
    or g24569 ( n25807 , n16514 , n5129 );
    or g24570 ( n2790 , n31090 , n24869 );
    or g24571 ( n4182 , n20025 , n16457 );
    or g24572 ( n21312 , n13097 , n21002 );
    not g24573 ( n32612 , n20713 );
    nor g24574 ( n2490 , n2236 , n24553 );
    or g24575 ( n30874 , n32585 , n11673 );
    and g24576 ( n12845 , n27369 , n7717 );
    or g24577 ( n14638 , n11046 , n12155 );
    or g24578 ( n9585 , n32857 , n16387 );
    buf g24579 ( n2117 , n12275 );
    or g24580 ( n29377 , n4041 , n1474 );
    or g24581 ( n12843 , n16468 , n4289 );
    or g24582 ( n15998 , n11455 , n20734 );
    or g24583 ( n33660 , n8432 , n16212 );
    and g24584 ( n32841 , n10650 , n7506 );
    and g24585 ( n5597 , n13616 , n20274 );
    or g24586 ( n8089 , n1119 , n22858 );
    xnor g24587 ( n1869 , n30342 , n4269 );
    or g24588 ( n10926 , n4814 , n5972 );
    or g24589 ( n22343 , n11046 , n20468 );
    not g24590 ( n29761 , n21105 );
    xnor g24591 ( n23164 , n33269 , n20138 );
    or g24592 ( n15543 , n13633 , n25499 );
    and g24593 ( n1997 , n31688 , n5799 );
    nor g24594 ( n17715 , n32715 , n6254 );
    xnor g24595 ( n34743 , n2468 , n4878 );
    xnor g24596 ( n26707 , n13592 , n23442 );
    or g24597 ( n13847 , n5422 , n13230 );
    and g24598 ( n18343 , n7721 , n23050 );
    and g24599 ( n15490 , n10906 , n28688 );
    or g24600 ( n3181 , n17361 , n28837 );
    or g24601 ( n27599 , n20593 , n31290 );
    or g24602 ( n7747 , n8958 , n26480 );
    xnor g24603 ( n29575 , n5122 , n19551 );
    and g24604 ( n7005 , n32409 , n2920 );
    nor g24605 ( n14836 , n7540 , n18760 );
    or g24606 ( n4903 , n5564 , n6711 );
    or g24607 ( n9876 , n22291 , n7666 );
    xnor g24608 ( n21219 , n34312 , n11142 );
    or g24609 ( n22172 , n13884 , n5010 );
    xnor g24610 ( n27959 , n30664 , n25548 );
    or g24611 ( n16410 , n33847 , n18488 );
    xnor g24612 ( n30537 , n12408 , n8607 );
    or g24613 ( n3107 , n22689 , n25306 );
    or g24614 ( n33479 , n31559 , n26390 );
    or g24615 ( n19050 , n23335 , n13904 );
    xnor g24616 ( n7662 , n26748 , n9789 );
    not g24617 ( n31921 , n19812 );
    xnor g24618 ( n22594 , n14481 , n4962 );
    nor g24619 ( n8801 , n31215 , n16113 );
    and g24620 ( n21121 , n29694 , n7236 );
    or g24621 ( n6532 , n31355 , n19490 );
    xnor g24622 ( n27376 , n1448 , n2825 );
    or g24623 ( n35490 , n23131 , n1535 );
    and g24624 ( n556 , n22695 , n9844 );
    or g24625 ( n13086 , n4962 , n3141 );
    or g24626 ( n22964 , n13071 , n24179 );
    not g24627 ( n21180 , n5060 );
    and g24628 ( n20033 , n30163 , n3945 );
    or g24629 ( n20420 , n31799 , n6660 );
    not g24630 ( n33654 , n14160 );
    and g24631 ( n3579 , n31059 , n13428 );
    xnor g24632 ( n25565 , n7416 , n35937 );
    xnor g24633 ( n34661 , n33695 , n2144 );
    or g24634 ( n16732 , n10860 , n51 );
    not g24635 ( n20338 , n27699 );
    xnor g24636 ( n5700 , n35747 , n7436 );
    nor g24637 ( n31291 , n30210 , n16961 );
    and g24638 ( n29372 , n34647 , n11220 );
    or g24639 ( n35902 , n10894 , n11144 );
    and g24640 ( n4743 , n11853 , n21263 );
    or g24641 ( n7840 , n27224 , n20441 );
    not g24642 ( n2170 , n29791 );
    or g24643 ( n29534 , n31425 , n28135 );
    and g24644 ( n12841 , n25071 , n5970 );
    xnor g24645 ( n25020 , n26916 , n31559 );
    nor g24646 ( n28935 , n3205 , n23848 );
    and g24647 ( n13638 , n20560 , n25428 );
    or g24648 ( n16643 , n785 , n908 );
    or g24649 ( n22369 , n25920 , n3419 );
    or g24650 ( n6186 , n3180 , n11518 );
    or g24651 ( n34302 , n6183 , n17974 );
    or g24652 ( n5808 , n22978 , n29953 );
    and g24653 ( n19288 , n13688 , n15563 );
    xnor g24654 ( n2922 , n1364 , n14681 );
    and g24655 ( n3199 , n11214 , n30409 );
    or g24656 ( n13918 , n23210 , n21977 );
    xnor g24657 ( n20378 , n25888 , n889 );
    xnor g24658 ( n20353 , n21068 , n10335 );
    or g24659 ( n13945 , n32792 , n25276 );
    or g24660 ( n8589 , n23867 , n24170 );
    or g24661 ( n17508 , n36044 , n308 );
    or g24662 ( n30274 , n1222 , n5538 );
    and g24663 ( n21510 , n35515 , n20994 );
    buf g24664 ( n15144 , n19120 );
    not g24665 ( n36017 , n13159 );
    nor g24666 ( n14391 , n25174 , n27434 );
    or g24667 ( n3690 , n20919 , n585 );
    and g24668 ( n25644 , n2475 , n10282 );
    xnor g24669 ( n4476 , n23577 , n33152 );
    or g24670 ( n6752 , n34668 , n29459 );
    nor g24671 ( n30569 , n27358 , n6686 );
    xnor g24672 ( n26785 , n31017 , n10171 );
    or g24673 ( n23777 , n110 , n20676 );
    not g24674 ( n12357 , n11455 );
    and g24675 ( n2829 , n1504 , n18600 );
    and g24676 ( n8389 , n11028 , n3423 );
    and g24677 ( n4037 , n18190 , n23023 );
    or g24678 ( n32444 , n26561 , n34537 );
    xnor g24679 ( n6731 , n8974 , n10894 );
    xnor g24680 ( n12284 , n29904 , n25246 );
    xnor g24681 ( n30142 , n6286 , n31215 );
    xnor g24682 ( n32497 , n27796 , n35927 );
    xnor g24683 ( n2155 , n6274 , n16862 );
    or g24684 ( n12119 , n1958 , n28455 );
    or g24685 ( n28815 , n28630 , n35422 );
    xnor g24686 ( n26165 , n8686 , n30742 );
    or g24687 ( n12670 , n32636 , n12035 );
    and g24688 ( n1379 , n19187 , n1691 );
    xnor g24689 ( n19835 , n24931 , n23733 );
    nor g24690 ( n23863 , n35927 , n5654 );
    or g24691 ( n11779 , n17588 , n9575 );
    and g24692 ( n16692 , n30657 , n16362 );
    and g24693 ( n26680 , n8485 , n24722 );
    and g24694 ( n11361 , n10727 , n14920 );
    buf g24695 ( n7293 , n4595 );
    xnor g24696 ( n3846 , n30114 , n4962 );
    xnor g24697 ( n34704 , n28429 , n29713 );
    or g24698 ( n2418 , n8432 , n21663 );
    or g24699 ( n5201 , n33681 , n7177 );
    xnor g24700 ( n19954 , n35386 , n27291 );
    and g24701 ( n24292 , n31654 , n32479 );
    or g24702 ( n14483 , n30686 , n17469 );
    or g24703 ( n21109 , n11466 , n28438 );
    or g24704 ( n7761 , n11046 , n4335 );
    or g24705 ( n21346 , n875 , n9429 );
    or g24706 ( n25191 , n35877 , n28324 );
    or g24707 ( n32803 , n14303 , n2134 );
    not g24708 ( n7771 , n26439 );
    nor g24709 ( n32955 , n9789 , n35782 );
    or g24710 ( n5811 , n25589 , n19173 );
    or g24711 ( n12508 , n29713 , n14978 );
    not g24712 ( n22451 , n16135 );
    or g24713 ( n7534 , n30955 , n18161 );
    not g24714 ( n4324 , n25264 );
    not g24715 ( n9773 , n10598 );
    or g24716 ( n15365 , n34596 , n34862 );
    nor g24717 ( n15102 , n28566 , n13656 );
    xnor g24718 ( n23915 , n18001 , n14319 );
    nor g24719 ( n23859 , n16620 , n32804 );
    nor g24720 ( n28390 , n1950 , n4178 );
    xnor g24721 ( n24385 , n35667 , n23604 );
    xnor g24722 ( n2040 , n7300 , n5780 );
    or g24723 ( n34476 , n23791 , n6951 );
    not g24724 ( n1326 , n2805 );
    and g24725 ( n2057 , n15103 , n366 );
    nor g24726 ( n7897 , n20356 , n33759 );
    and g24727 ( n15040 , n22060 , n14307 );
    or g24728 ( n20466 , n8517 , n17818 );
    xnor g24729 ( n22139 , n9493 , n19544 );
    or g24730 ( n7386 , n24959 , n30947 );
    and g24731 ( n33174 , n18833 , n2634 );
    or g24732 ( n35658 , n15332 , n32701 );
    or g24733 ( n24774 , n8566 , n32581 );
    and g24734 ( n24769 , n28672 , n7129 );
    or g24735 ( n23580 , n34374 , n18272 );
    and g24736 ( n6470 , n8318 , n9560 );
    not g24737 ( n14964 , n30969 );
    or g24738 ( n9643 , n33144 , n8452 );
    and g24739 ( n27099 , n35456 , n7283 );
    or g24740 ( n30157 , n11046 , n11487 );
    and g24741 ( n27844 , n19181 , n32244 );
    or g24742 ( n24142 , n27216 , n1763 );
    or g24743 ( n14432 , n35454 , n15070 );
    and g24744 ( n924 , n35903 , n32111 );
    and g24745 ( n34209 , n34305 , n32654 );
    or g24746 ( n6295 , n30304 , n5826 );
    or g24747 ( n24724 , n30440 , n5752 );
    and g24748 ( n21893 , n5822 , n12672 );
    or g24749 ( n9570 , n4288 , n1087 );
    or g24750 ( n33574 , n43 , n7448 );
    xnor g24751 ( n29637 , n13776 , n30126 );
    xnor g24752 ( n30692 , n19570 , n19553 );
    or g24753 ( n14465 , n27401 , n9675 );
    xnor g24754 ( n3737 , n13789 , n4288 );
    not g24755 ( n8666 , n17005 );
    or g24756 ( n33824 , n13729 , n5900 );
    or g24757 ( n6846 , n10030 , n26371 );
    xnor g24758 ( n24629 , n9657 , n32857 );
    or g24759 ( n7275 , n29839 , n16874 );
    or g24760 ( n10886 , n3689 , n14076 );
    nor g24761 ( n15167 , n5287 , n31957 );
    and g24762 ( n4916 , n11500 , n30543 );
    or g24763 ( n24952 , n26783 , n20284 );
    xnor g24764 ( n22308 , n27037 , n9789 );
    or g24765 ( n33547 , n16194 , n7127 );
    not g24766 ( n1267 , n1254 );
    xnor g24767 ( n47 , n948 , n1941 );
    and g24768 ( n14242 , n2120 , n20023 );
    and g24769 ( n18837 , n27486 , n16719 );
    or g24770 ( n17476 , n31272 , n31928 );
    or g24771 ( n11939 , n24196 , n21439 );
    nor g24772 ( n31824 , n1950 , n22429 );
    and g24773 ( n15924 , n4612 , n26674 );
    or g24774 ( n30021 , n1695 , n19836 );
    xnor g24775 ( n19102 , n6912 , n24371 );
    xnor g24776 ( n12597 , n29993 , n15877 );
    or g24777 ( n3980 , n34166 , n8153 );
    or g24778 ( n26421 , n19900 , n5779 );
    not g24779 ( n21780 , n19939 );
    or g24780 ( n1681 , n32877 , n17612 );
    xor g24781 ( n28105 , n5390 , n26041 );
    xnor g24782 ( n7252 , n17803 , n31868 );
    or g24783 ( n28244 , n9457 , n28455 );
    or g24784 ( n9988 , n24371 , n17054 );
    or g24785 ( n29720 , n15886 , n29639 );
    or g24786 ( n16323 , n18760 , n1642 );
    nor g24787 ( n6026 , n19246 , n4899 );
    or g24788 ( n10588 , n23290 , n33766 );
    and g24789 ( n19042 , n31779 , n27553 );
    or g24790 ( n33595 , n10358 , n27159 );
    nor g24791 ( n24180 , n20699 , n799 );
    and g24792 ( n18161 , n14702 , n11710 );
    or g24793 ( n35742 , n29878 , n23599 );
    and g24794 ( n6172 , n14475 , n18360 );
    or g24795 ( n5710 , n31289 , n27353 );
    and g24796 ( n6632 , n29521 , n21946 );
    xnor g24797 ( n18323 , n21457 , n9789 );
    xnor g24798 ( n12835 , n30 , n11169 );
    and g24799 ( n12388 , n20621 , n12261 );
    not g24800 ( n31902 , n28438 );
    or g24801 ( n33345 , n28431 , n9731 );
    or g24802 ( n35035 , n21420 , n21644 );
    nor g24803 ( n7864 , n32745 , n7448 );
    nor g24804 ( n15602 , n28043 , n20486 );
    or g24805 ( n14205 , n9068 , n2446 );
    or g24806 ( n23083 , n8432 , n21502 );
    nor g24807 ( n16146 , n23604 , n24435 );
    and g24808 ( n36087 , n13842 , n33703 );
    xnor g24809 ( n5600 , n24521 , n32979 );
    and g24810 ( n807 , n774 , n16432 );
    not g24811 ( n3928 , n31799 );
    or g24812 ( n4877 , n812 , n17974 );
    and g24813 ( n3104 , n6675 , n17568 );
    not g24814 ( n15372 , n4472 );
    not g24815 ( n31273 , n25602 );
    nor g24816 ( n3790 , n11455 , n12205 );
    or g24817 ( n4394 , n28693 , n13664 );
    or g24818 ( n14066 , n6438 , n6553 );
    xnor g24819 ( n32029 , n2133 , n11613 );
    or g24820 ( n23031 , n13456 , n28987 );
    xnor g24821 ( n6080 , n284 , n35895 );
    or g24822 ( n31661 , n31799 , n3838 );
    and g24823 ( n24892 , n35874 , n1005 );
    not g24824 ( n6279 , n4960 );
    or g24825 ( n36004 , n9949 , n7439 );
    xnor g24826 ( n5802 , n33333 , n29686 );
    and g24827 ( n14098 , n24515 , n31208 );
    and g24828 ( n34622 , n3719 , n18236 );
    or g24829 ( n10658 , n30102 , n3840 );
    or g24830 ( n3105 , n4960 , n10158 );
    xnor g24831 ( n28923 , n14209 , n16897 );
    nor g24832 ( n4775 , n14128 , n35834 );
    xnor g24833 ( n6059 , n34054 , n12088 );
    or g24834 ( n30491 , n27226 , n22814 );
    or g24835 ( n20012 , n28962 , n7647 );
    nor g24836 ( n8878 , n18150 , n7700 );
    and g24837 ( n20784 , n17092 , n22586 );
    nor g24838 ( n32887 , n4960 , n7318 );
    not g24839 ( n21781 , n15403 );
    xnor g24840 ( n32009 , n15316 , n1260 );
    and g24841 ( n26242 , n31648 , n24939 );
    and g24842 ( n5723 , n8145 , n8574 );
    xnor g24843 ( n19280 , n31953 , n18379 );
    or g24844 ( n9865 , n30715 , n21644 );
    or g24845 ( n35898 , n17568 , n1736 );
    xnor g24846 ( n5169 , n13078 , n731 );
    or g24847 ( n6824 , n14982 , n35565 );
    or g24848 ( n11788 , n23604 , n8348 );
    xnor g24849 ( n11942 , n11618 , n3106 );
    or g24850 ( n27097 , n34725 , n5618 );
    and g24851 ( n12903 , n4099 , n7154 );
    nor g24852 ( n27875 , n4960 , n26211 );
    not g24853 ( n14386 , n31799 );
    or g24854 ( n4861 , n7608 , n12281 );
    nor g24855 ( n14208 , n23749 , n15835 );
    and g24856 ( n29323 , n7106 , n21174 );
    or g24857 ( n7017 , n11806 , n18811 );
    xnor g24858 ( n35778 , n32442 , n35927 );
    or g24859 ( n16117 , n8409 , n20817 );
    xnor g24860 ( n21352 , n5667 , n11864 );
    not g24861 ( n31295 , n24371 );
    xnor g24862 ( n26226 , n6820 , n32584 );
    and g24863 ( n33148 , n2833 , n30731 );
    or g24864 ( n32794 , n4288 , n28009 );
    buf g24865 ( n21673 , n33206 );
    not g24866 ( n3177 , n29902 );
    or g24867 ( n32494 , n32083 , n2814 );
    xnor g24868 ( n17466 , n31603 , n568 );
    not g24869 ( n23071 , n4962 );
    or g24870 ( n35889 , n35104 , n4695 );
    xnor g24871 ( n26257 , n22451 , n21699 );
    nor g24872 ( n4941 , n17662 , n30400 );
    or g24873 ( n24813 , n11873 , n32799 );
    and g24874 ( n12432 , n6135 , n34116 );
    xnor g24875 ( n30562 , n21430 , n25343 );
    and g24876 ( n23332 , n6747 , n32009 );
    or g24877 ( n29482 , n30798 , n22501 );
    or g24878 ( n23539 , n18379 , n31362 );
    or g24879 ( n31228 , n31897 , n18207 );
    or g24880 ( n28673 , n11949 , n18264 );
    or g24881 ( n4620 , n11455 , n19668 );
    not g24882 ( n34785 , n4517 );
    or g24883 ( n8158 , n25821 , n4621 );
    and g24884 ( n25209 , n7604 , n17057 );
    xnor g24885 ( n33332 , n26030 , n5756 );
    or g24886 ( n28009 , n33885 , n8752 );
    and g24887 ( n5476 , n6312 , n9356 );
    or g24888 ( n21932 , n21026 , n1557 );
    and g24889 ( n23483 , n2692 , n19869 );
    or g24890 ( n26209 , n6561 , n28013 );
    not g24891 ( n29134 , n29713 );
    nor g24892 ( n17740 , n3946 , n19013 );
    xnor g24893 ( n10759 , n17146 , n15120 );
    not g24894 ( n5890 , n24691 );
    or g24895 ( n18104 , n16707 , n12879 );
    and g24896 ( n1837 , n11682 , n33816 );
    and g24897 ( n35211 , n1579 , n21368 );
    or g24898 ( n1053 , n15291 , n3858 );
    and g24899 ( n17324 , n20156 , n23423 );
    or g24900 ( n7333 , n17072 , n803 );
    nor g24901 ( n8396 , n3222 , n13332 );
    or g24902 ( n22209 , n11250 , n9217 );
    and g24903 ( n17294 , n8986 , n16317 );
    or g24904 ( n32166 , n7898 , n6950 );
    or g24905 ( n13025 , n34866 , n33590 );
    or g24906 ( n30197 , n27291 , n849 );
    or g24907 ( n23493 , n2331 , n23509 );
    nor g24908 ( n13385 , n32857 , n25788 );
    or g24909 ( n10842 , n26709 , n1474 );
    xnor g24910 ( n3212 , n78 , n19551 );
    buf g24911 ( n19336 , n15290 );
    nor g24912 ( n26537 , n4960 , n16771 );
    not g24913 ( n19983 , n18934 );
    or g24914 ( n3182 , n15464 , n34792 );
    not g24915 ( n27145 , n32095 );
    nor g24916 ( n17764 , n30742 , n12743 );
    xnor g24917 ( n31516 , n4475 , n28711 );
    xnor g24918 ( n23591 , n15856 , n32828 );
    not g24919 ( n382 , n9789 );
    nor g24920 ( n16103 , n32857 , n9136 );
    not g24921 ( n28807 , n2882 );
    and g24922 ( n34061 , n13811 , n35293 );
    or g24923 ( n23441 , n5488 , n33416 );
    xnor g24924 ( n4352 , n13702 , n32584 );
    xnor g24925 ( n13409 , n34585 , n9789 );
    and g24926 ( n18591 , n12219 , n2169 );
    or g24927 ( n29474 , n3205 , n29887 );
    and g24928 ( n23848 , n23480 , n9248 );
    buf g24929 ( n5868 , n19566 );
    or g24930 ( n13450 , n19622 , n15805 );
    or g24931 ( n7298 , n11455 , n7262 );
    and g24932 ( n6818 , n19068 , n6036 );
    and g24933 ( n2977 , n21150 , n27313 );
    or g24934 ( n14996 , n24385 , n21518 );
    and g24935 ( n28740 , n6162 , n2147 );
    buf g24936 ( n2119 , n23545 );
    and g24937 ( n23352 , n20014 , n19965 );
    or g24938 ( n6505 , n4461 , n860 );
    or g24939 ( n16940 , n8793 , n32414 );
    not g24940 ( n33737 , n29727 );
    nor g24941 ( n22170 , n21918 , n17248 );
    or g24942 ( n7576 , n14574 , n3842 );
    buf g24943 ( n22241 , n6037 );
    not g24944 ( n14285 , n8725 );
    xnor g24945 ( n9639 , n14269 , n33398 );
    and g24946 ( n20531 , n14776 , n29119 );
    nor g24947 ( n22132 , n32095 , n10997 );
    xnor g24948 ( n4947 , n24040 , n32584 );
    and g24949 ( n19235 , n33281 , n21401 );
    and g24950 ( n15304 , n2844 , n15801 );
    not g24951 ( n34937 , n4960 );
    or g24952 ( n23951 , n3222 , n9065 );
    and g24953 ( n17499 , n24029 , n18455 );
    buf g24954 ( n28969 , n4023 );
    nor g24955 ( n16811 , n26696 , n12428 );
    xnor g24956 ( n7202 , n19397 , n21361 );
    xnor g24957 ( n12684 , n16834 , n24371 );
    and g24958 ( n9267 , n25253 , n19943 );
    and g24959 ( n27944 , n5595 , n6362 );
    not g24960 ( n25762 , n3480 );
    or g24961 ( n6775 , n33731 , n16847 );
    and g24962 ( n19228 , n27270 , n22627 );
    not g24963 ( n31541 , n16223 );
    or g24964 ( n14867 , n22035 , n2384 );
    xnor g24965 ( n32952 , n30597 , n29846 );
    or g24966 ( n3031 , n35360 , n26480 );
    not g24967 ( n6156 , n31272 );
    and g24968 ( n2042 , n2016 , n36071 );
    or g24969 ( n5383 , n23194 , n26002 );
    or g24970 ( n19352 , n22154 , n18065 );
    xnor g24971 ( n9942 , n20929 , n19335 );
    and g24972 ( n1472 , n24033 , n19418 );
    or g24973 ( n4511 , n33949 , n25761 );
    or g24974 ( n92 , n14739 , n32329 );
    nor g24975 ( n2408 , n32584 , n15064 );
    xnor g24976 ( n25994 , n7894 , n27391 );
    or g24977 ( n31567 , n19071 , n18065 );
    nor g24978 ( n34885 , n25767 , n9358 );
    xnor g24979 ( n8454 , n5804 , n32191 );
    or g24980 ( n21256 , n30235 , n34361 );
    nor g24981 ( n34765 , n26844 , n28993 );
    or g24982 ( n25117 , n15320 , n32039 );
    or g24983 ( n181 , n26229 , n1474 );
    or g24984 ( n12567 , n615 , n26112 );
    xnor g24985 ( n3890 , n11285 , n29352 );
    xnor g24986 ( n1000 , n23173 , n35927 );
    or g24987 ( n25395 , n29038 , n19336 );
    xnor g24988 ( n26938 , n30879 , n596 );
    or g24989 ( n16556 , n6786 , n1783 );
    nor g24990 ( n26136 , n17568 , n688 );
    xnor g24991 ( n17703 , n34763 , n4758 );
    or g24992 ( n1239 , n26407 , n32329 );
    or g24993 ( n29704 , n29713 , n5695 );
    nor g24994 ( n9376 , n15886 , n2394 );
    or g24995 ( n31256 , n21032 , n22961 );
    not g24996 ( n29084 , n13885 );
    and g24997 ( n4979 , n23562 , n34267 );
    not g24998 ( n11967 , n17568 );
    and g24999 ( n20559 , n32534 , n17924 );
    or g25000 ( n23295 , n4878 , n34762 );
    or g25001 ( n14548 , n8936 , n19952 );
    and g25002 ( n35230 , n12157 , n13157 );
    or g25003 ( n12183 , n10219 , n9772 );
    not g25004 ( n12474 , n10975 );
    or g25005 ( n15437 , n10529 , n33034 );
    xnor g25006 ( n31393 , n24697 , n25958 );
    and g25007 ( n34804 , n3377 , n17214 );
    or g25008 ( n19588 , n4962 , n29715 );
    nor g25009 ( n16835 , n15183 , n7163 );
    and g25010 ( n11568 , n31409 , n32936 );
    or g25011 ( n29280 , n4789 , n20271 );
    and g25012 ( n492 , n11562 , n33724 );
    or g25013 ( n18131 , n1950 , n17961 );
    xnor g25014 ( n1770 , n15697 , n17816 );
    or g25015 ( n19558 , n22412 , n28288 );
    xnor g25016 ( n5156 , n30334 , n35927 );
    xnor g25017 ( n10302 , n9334 , n16506 );
    and g25018 ( n25468 , n34645 , n14511 );
    or g25019 ( n8964 , n23956 , n27580 );
    or g25020 ( n17597 , n27376 , n21579 );
    xnor g25021 ( n5227 , n21082 , n7914 );
    or g25022 ( n28576 , n1867 , n3437 );
    and g25023 ( n7619 , n13560 , n24699 );
    or g25024 ( n9131 , n31799 , n9066 );
    or g25025 ( n29301 , n18379 , n14098 );
    or g25026 ( n23525 , n28614 , n29562 );
    or g25027 ( n20994 , n32573 , n23462 );
    or g25028 ( n12598 , n18914 , n10478 );
    or g25029 ( n33609 , n15624 , n34084 );
    xnor g25030 ( n7820 , n2943 , n533 );
    and g25031 ( n10212 , n30227 , n28122 );
    or g25032 ( n21777 , n31525 , n15732 );
    or g25033 ( n14309 , n34962 , n8153 );
    or g25034 ( n1664 , n29713 , n25729 );
    xnor g25035 ( n6884 , n18769 , n5287 );
    or g25036 ( n19032 , n28315 , n13217 );
    and g25037 ( n17771 , n6795 , n30972 );
    and g25038 ( n33680 , n2551 , n3216 );
    nor g25039 ( n33833 , n3957 , n10745 );
    and g25040 ( n10081 , n8284 , n35278 );
    nor g25041 ( n24007 , n25602 , n2717 );
    or g25042 ( n5829 , n6495 , n12124 );
    or g25043 ( n29972 , n26207 , n35445 );
    and g25044 ( n8348 , n26416 , n9710 );
    or g25045 ( n23988 , n13987 , n31067 );
    or g25046 ( n35316 , n10462 , n4172 );
    or g25047 ( n12210 , n34810 , n33416 );
    or g25048 ( n34980 , n24241 , n31055 );
    xnor g25049 ( n660 , n3050 , n830 );
    nor g25050 ( n35676 , n8345 , n32379 );
    xnor g25051 ( n28039 , n22571 , n16922 );
    and g25052 ( n29262 , n3588 , n12773 );
    xnor g25053 ( n26350 , n2812 , n26633 );
    or g25054 ( n9129 , n17761 , n178 );
    xnor g25055 ( n3536 , n20582 , n7540 );
    xnor g25056 ( n18317 , n12599 , n7601 );
    or g25057 ( n8132 , n2055 , n30763 );
    xnor g25058 ( n23059 , n25772 , n32621 );
    or g25059 ( n18720 , n11798 , n4426 );
    nor g25060 ( n17230 , n31799 , n19394 );
    or g25061 ( n4498 , n30615 , n24138 );
    or g25062 ( n5819 , n22321 , n24108 );
    nor g25063 ( n1964 , n7515 , n11732 );
    xnor g25064 ( n30314 , n28451 , n30742 );
    nor g25065 ( n17203 , n34371 , n18819 );
    or g25066 ( n9659 , n28780 , n24141 );
    not g25067 ( n11924 , n21258 );
    not g25068 ( n12273 , n14902 );
    or g25069 ( n10312 , n302 , n24088 );
    xnor g25070 ( n17004 , n6269 , n12144 );
    xnor g25071 ( n17506 , n10996 , n31522 );
    and g25072 ( n23131 , n16242 , n32658 );
    xnor g25073 ( n33151 , n13710 , n21937 );
    not g25074 ( n34528 , n19811 );
    xnor g25075 ( n3744 , n19018 , n29855 );
    not g25076 ( n519 , n4758 );
    xnor g25077 ( n14440 , n35212 , n15886 );
    xnor g25078 ( n24872 , n14575 , n32715 );
    xnor g25079 ( n16419 , n16638 , n7247 );
    or g25080 ( n28156 , n36053 , n32608 );
    not g25081 ( n1129 , n9187 );
    or g25082 ( n32099 , n28107 , n1955 );
    and g25083 ( n8827 , n11700 , n11117 );
    not g25084 ( n16819 , n21594 );
    not g25085 ( n9873 , n18941 );
    xnor g25086 ( n16821 , n7777 , n29048 );
    and g25087 ( n24673 , n11981 , n4356 );
    and g25088 ( n30994 , n1622 , n11203 );
    xnor g25089 ( n18585 , n9001 , n31066 );
    xnor g25090 ( n18992 , n28299 , n17234 );
    nor g25091 ( n6319 , n31289 , n11172 );
    or g25092 ( n25826 , n12984 , n21862 );
    not g25093 ( n24595 , n35067 );
    or g25094 ( n4064 , n17096 , n14119 );
    or g25095 ( n5849 , n7068 , n19336 );
    xnor g25096 ( n11565 , n30658 , n16922 );
    xnor g25097 ( n22210 , n18299 , n9015 );
    or g25098 ( n19417 , n6027 , n11308 );
    or g25099 ( n28542 , n4960 , n11567 );
    and g25100 ( n996 , n30839 , n26837 );
    and g25101 ( n13889 , n12158 , n2856 );
    or g25102 ( n6729 , n9568 , n30224 );
    and g25103 ( n6906 , n27506 , n24230 );
    xnor g25104 ( n35637 , n5409 , n2017 );
    nor g25105 ( n21152 , n16620 , n35697 );
    or g25106 ( n27105 , n15477 , n10400 );
    or g25107 ( n35554 , n17442 , n10861 );
    xnor g25108 ( n5541 , n6299 , n20253 );
    or g25109 ( n23304 , n20032 , n8366 );
    nor g25110 ( n22619 , n3776 , n31411 );
    or g25111 ( n28645 , n7893 , n36000 );
    or g25112 ( n29429 , n3222 , n14021 );
    and g25113 ( n31368 , n23777 , n30642 );
    or g25114 ( n34394 , n22291 , n27850 );
    and g25115 ( n4337 , n17762 , n31798 );
    or g25116 ( n9077 , n34835 , n6690 );
    or g25117 ( n25949 , n4962 , n8387 );
    and g25118 ( n16843 , n5047 , n33662 );
    and g25119 ( n27536 , n2415 , n8449 );
    and g25120 ( n32636 , n7732 , n16340 );
    and g25121 ( n16197 , n17439 , n12478 );
    and g25122 ( n33420 , n6049 , n11983 );
    not g25123 ( n5058 , n10216 );
    or g25124 ( n10530 , n30818 , n17964 );
    and g25125 ( n6929 , n7840 , n8160 );
    and g25126 ( n7050 , n15417 , n13171 );
    buf g25127 ( n25118 , n5469 );
    or g25128 ( n20150 , n13231 , n30287 );
    not g25129 ( n29909 , n3404 );
    or g25130 ( n34800 , n9291 , n21018 );
    or g25131 ( n35624 , n27291 , n31507 );
    or g25132 ( n12892 , n25217 , n8153 );
    and g25133 ( n27275 , n15892 , n34689 );
    nor g25134 ( n20993 , n32857 , n2363 );
    buf g25135 ( n14076 , n12725 );
    and g25136 ( n27630 , n9777 , n7077 );
    or g25137 ( n21365 , n19763 , n15378 );
    nor g25138 ( n10924 , n26222 , n9921 );
    or g25139 ( n21657 , n30616 , n33762 );
    xnor g25140 ( n16851 , n13138 , n25927 );
    or g25141 ( n9917 , n34631 , n28248 );
    nor g25142 ( n22988 , n4209 , n26634 );
    and g25143 ( n19013 , n17003 , n11149 );
    or g25144 ( n25146 , n20110 , n24005 );
    nor g25145 ( n12711 , n830 , n17141 );
    or g25146 ( n32511 , n9175 , n26648 );
    or g25147 ( n31813 , n24371 , n3368 );
    and g25148 ( n36079 , n28580 , n12253 );
    or g25149 ( n14585 , n8209 , n6459 );
    or g25150 ( n18528 , n9658 , n25684 );
    xnor g25151 ( n27680 , n8380 , n16922 );
    and g25152 ( n22693 , n3283 , n10025 );
    or g25153 ( n23938 , n26651 , n3239 );
    and g25154 ( n10570 , n9422 , n31516 );
    or g25155 ( n31914 , n33458 , n6459 );
    xnor g25156 ( n19572 , n30565 , n34318 );
    or g25157 ( n16599 , n15464 , n11929 );
    or g25158 ( n23816 , n6116 , n33034 );
    or g25159 ( n22728 , n29430 , n23254 );
    or g25160 ( n13087 , n17658 , n4081 );
    and g25161 ( n11240 , n3834 , n14766 );
    or g25162 ( n4934 , n16615 , n8352 );
    or g25163 ( n10854 , n32732 , n31389 );
    and g25164 ( n27860 , n8310 , n30475 );
    not g25165 ( n24408 , n2156 );
    or g25166 ( n33718 , n30100 , n7808 );
    xnor g25167 ( n4879 , n19800 , n12922 );
    xnor g25168 ( n16827 , n839 , n9789 );
    xnor g25169 ( n29886 , n19217 , n32584 );
    or g25170 ( n7395 , n3598 , n19501 );
    or g25171 ( n1971 , n33284 , n18542 );
    and g25172 ( n5816 , n27139 , n11025 );
    and g25173 ( n16473 , n14100 , n25900 );
    or g25174 ( n34603 , n17907 , n10634 );
    xnor g25175 ( n33974 , n26941 , n18761 );
    xnor g25176 ( n22616 , n31349 , n16620 );
    not g25177 ( n15009 , n13881 );
    xnor g25178 ( n22234 , n1000 , n33229 );
    or g25179 ( n13443 , n25151 , n35141 );
    or g25180 ( n1717 , n17568 , n4997 );
    or g25181 ( n9227 , n14968 , n5208 );
    not g25182 ( n183 , n23440 );
    nor g25183 ( n11475 , n10768 , n32893 );
    or g25184 ( n15806 , n11363 , n34673 );
    or g25185 ( n11092 , n19256 , n27488 );
    xnor g25186 ( n12820 , n7937 , n30742 );
    or g25187 ( n34513 , n4878 , n21604 );
    and g25188 ( n9273 , n31847 , n8053 );
    or g25189 ( n19160 , n1950 , n13454 );
    xnor g25190 ( n15450 , n34066 , n25174 );
    or g25191 ( n30696 , n34529 , n29106 );
    xnor g25192 ( n36091 , n2970 , n20629 );
    and g25193 ( n10265 , n9229 , n8377 );
    and g25194 ( n25997 , n20347 , n13134 );
    not g25195 ( n18919 , n35917 );
    xnor g25196 ( n32775 , n23902 , n7711 );
    or g25197 ( n18124 , n35118 , n14215 );
    xnor g25198 ( n33291 , n9413 , n10894 );
    or g25199 ( n24047 , n6726 , n5610 );
    or g25200 ( n16236 , n10894 , n15657 );
    xnor g25201 ( n29912 , n812 , n32715 );
    or g25202 ( n9026 , n19661 , n22961 );
    or g25203 ( n16867 , n9791 , n3583 );
    not g25204 ( n31756 , n1950 );
    or g25205 ( n14190 , n25126 , n12964 );
    xnor g25206 ( n155 , n30027 , n31429 );
    xnor g25207 ( n23238 , n28292 , n1438 );
    xnor g25208 ( n34641 , n31149 , n1950 );
    and g25209 ( n5440 , n11674 , n3495 );
    or g25210 ( n5107 , n2400 , n35766 );
    xnor g25211 ( n14142 , n34037 , n10205 );
    and g25212 ( n17095 , n28629 , n2084 );
    or g25213 ( n29700 , n19002 , n8043 );
    and g25214 ( n10356 , n17318 , n34157 );
    nor g25215 ( n3891 , n15097 , n1534 );
    or g25216 ( n11895 , n13553 , n20212 );
    or g25217 ( n2755 , n8429 , n35757 );
    or g25218 ( n34237 , n31289 , n9556 );
    and g25219 ( n33373 , n28118 , n6418 );
    or g25220 ( n16493 , n24332 , n30155 );
    or g25221 ( n3032 , n23967 , n21579 );
    xnor g25222 ( n21613 , n21344 , n21974 );
    or g25223 ( n27052 , n30742 , n3099 );
    nor g25224 ( n1100 , n29089 , n20330 );
    xnor g25225 ( n30003 , n20829 , n10894 );
    or g25226 ( n7854 , n12616 , n9951 );
    or g25227 ( n35006 , n23589 , n30287 );
    xnor g25228 ( n34111 , n29611 , n11455 );
    or g25229 ( n6934 , n30742 , n32856 );
    and g25230 ( n32469 , n2278 , n18392 );
    and g25231 ( n30069 , n8649 , n17156 );
    or g25232 ( n20900 , n22291 , n32133 );
    or g25233 ( n450 , n19551 , n6627 );
    and g25234 ( n16041 , n14041 , n8327 );
    buf g25235 ( n5457 , n14017 );
    nor g25236 ( n10435 , n29713 , n8650 );
    or g25237 ( n18276 , n19551 , n4045 );
    or g25238 ( n27026 , n4954 , n23626 );
    not g25239 ( n27770 , n2029 );
    and g25240 ( n29650 , n7942 , n25880 );
    xnor g25241 ( n9391 , n19554 , n21569 );
    or g25242 ( n28379 , n33198 , n25036 );
    xnor g25243 ( n8889 , n20869 , n16773 );
    xnor g25244 ( n5789 , n12611 , n6395 );
    nor g25245 ( n4378 , n33524 , n27178 );
    xnor g25246 ( n19150 , n7984 , n6794 );
    and g25247 ( n36085 , n30681 , n14151 );
    nor g25248 ( n33914 , n2882 , n23186 );
    and g25249 ( n34383 , n30087 , n33064 );
    or g25250 ( n992 , n18992 , n26002 );
    xnor g25251 ( n7586 , n27479 , n19728 );
    or g25252 ( n32022 , n2408 , n23811 );
    and g25253 ( n34897 , n22602 , n9350 );
    and g25254 ( n19433 , n28015 , n22854 );
    xnor g25255 ( n17772 , n338 , n32618 );
    not g25256 ( n17600 , n29145 );
    nor g25257 ( n21151 , n1719 , n20096 );
    and g25258 ( n8630 , n25869 , n23110 );
    or g25259 ( n7146 , n33996 , n25567 );
    or g25260 ( n28041 , n30161 , n23626 );
    xnor g25261 ( n32600 , n11927 , n3205 );
    not g25262 ( n6321 , n22291 );
    or g25263 ( n20721 , n12859 , n35608 );
    xnor g25264 ( n22526 , n29796 , n31799 );
    or g25265 ( n11222 , n11455 , n32538 );
    or g25266 ( n15929 , n28960 , n3188 );
    or g25267 ( n6878 , n30290 , n11593 );
    or g25268 ( n25622 , n25429 , n4363 );
    or g25269 ( n4112 , n13969 , n15109 );
    and g25270 ( n28770 , n27320 , n27419 );
    nor g25271 ( n12872 , n5067 , n19452 );
    xnor g25272 ( n28921 , n15584 , n18398 );
    not g25273 ( n6720 , n3205 );
    not g25274 ( n15117 , n11996 );
    nor g25275 ( n9574 , n99 , n19834 );
    xnor g25276 ( n13941 , n30485 , n3946 );
    or g25277 ( n16364 , n955 , n2090 );
    and g25278 ( n10651 , n8562 , n35502 );
    or g25279 ( n10891 , n34934 , n8090 );
    not g25280 ( n27903 , n35422 );
    or g25281 ( n34300 , n35224 , n11703 );
    or g25282 ( n35234 , n32813 , n17992 );
    xnor g25283 ( n16735 , n5441 , n25304 );
    and g25284 ( n7315 , n26215 , n9925 );
    nor g25285 ( n4187 , n2342 , n31541 );
    xnor g25286 ( n25811 , n18238 , n11046 );
    and g25287 ( n9702 , n32327 , n26285 );
    nor g25288 ( n23481 , n30742 , n25911 );
    or g25289 ( n32873 , n12409 , n471 );
    or g25290 ( n6108 , n4288 , n13789 );
    or g25291 ( n31465 , n17696 , n1516 );
    or g25292 ( n28607 , n4962 , n25793 );
    or g25293 ( n7794 , n27470 , n14706 );
    and g25294 ( n28275 , n24522 , n16960 );
    xnor g25295 ( n22815 , n5478 , n32857 );
    or g25296 ( n29215 , n5155 , n27728 );
    or g25297 ( n20770 , n33783 , n24570 );
    or g25298 ( n9965 , n20751 , n29872 );
    not g25299 ( n20070 , n3196 );
    xnor g25300 ( n18159 , n17670 , n20268 );
    xnor g25301 ( n11492 , n11442 , n19551 );
    not g25302 ( n3892 , n2606 );
    or g25303 ( n35683 , n15906 , n20812 );
    and g25304 ( n32250 , n11160 , n26824 );
    or g25305 ( n12615 , n17890 , n11089 );
    and g25306 ( n308 , n17870 , n26201 );
    or g25307 ( n15008 , n22883 , n14774 );
    or g25308 ( n6959 , n32124 , n33042 );
    nor g25309 ( n28854 , n33169 , n24795 );
    or g25310 ( n29901 , n9793 , n30034 );
    xnor g25311 ( n33997 , n2363 , n25194 );
    and g25312 ( n11470 , n20908 , n15830 );
    not g25313 ( n760 , n5315 );
    or g25314 ( n25436 , n31289 , n15136 );
    xnor g25315 ( n34319 , n12696 , n18918 );
    not g25316 ( n18787 , n3770 );
    nor g25317 ( n17237 , n21942 , n24505 );
    and g25318 ( n4774 , n4452 , n15990 );
    not g25319 ( n32128 , n22200 );
    or g25320 ( n26318 , n23038 , n4081 );
    not g25321 ( n4024 , n2029 );
    nor g25322 ( n36027 , n776 , n2313 );
    and g25323 ( n15781 , n24449 , n8915 );
    and g25324 ( n6206 , n20608 , n18467 );
    or g25325 ( n27013 , n24368 , n2137 );
    or g25326 ( n25640 , n11852 , n2814 );
    or g25327 ( n10033 , n4827 , n1557 );
    not g25328 ( n350 , n15464 );
    and g25329 ( n1476 , n11998 , n31676 );
    and g25330 ( n28546 , n16627 , n34459 );
    or g25331 ( n30153 , n31086 , n20529 );
    or g25332 ( n12697 , n13238 , n7529 );
    xnor g25333 ( n5240 , n19171 , n9860 );
    xnor g25334 ( n16769 , n11730 , n2077 );
    or g25335 ( n17440 , n21808 , n17233 );
    and g25336 ( n11982 , n30824 , n5715 );
    or g25337 ( n11397 , n19368 , n22858 );
    and g25338 ( n36078 , n22415 , n32115 );
    xnor g25339 ( n90 , n20067 , n31056 );
    and g25340 ( n27144 , n31257 , n23786 );
    xor g25341 ( n25587 , n5683 , n8523 );
    or g25342 ( n9515 , n30742 , n5991 );
    not g25343 ( n15096 , n11379 );
    nor g25344 ( n28769 , n31799 , n17577 );
    or g25345 ( n9711 , n27434 , n17962 );
    and g25346 ( n18675 , n7462 , n17268 );
    nor g25347 ( n9628 , n25147 , n9555 );
    xor g25348 ( n4183 , n10576 , n6911 );
    not g25349 ( n776 , n2533 );
    xnor g25350 ( n31089 , n30660 , n7540 );
    xnor g25351 ( n17853 , n9296 , n26141 );
    not g25352 ( n15519 , n6308 );
    and g25353 ( n20547 , n13431 , n33260 );
    or g25354 ( n815 , n8187 , n3352 );
    xor g25355 ( n28210 , n29522 , n12152 );
    xnor g25356 ( n14201 , n26508 , n29713 );
    and g25357 ( n3479 , n27920 , n8808 );
    not g25358 ( n23805 , n3239 );
    and g25359 ( n9874 , n25224 , n28207 );
    or g25360 ( n2050 , n4878 , n5026 );
    or g25361 ( n22845 , n3003 , n29545 );
    or g25362 ( n21878 , n35931 , n2955 );
    not g25363 ( n12144 , n16620 );
    or g25364 ( n35126 , n6774 , n33098 );
    xnor g25365 ( n5743 , n19147 , n25572 );
    not g25366 ( n30540 , n24371 );
    or g25367 ( n30151 , n5653 , n5925 );
    or g25368 ( n23672 , n23602 , n32697 );
    and g25369 ( n6592 , n19559 , n15706 );
    or g25370 ( n12982 , n11190 , n28550 );
    or g25371 ( n27334 , n5520 , n28933 );
    or g25372 ( n1915 , n25378 , n25594 );
    or g25373 ( n6443 , n15886 , n29395 );
    or g25374 ( n21136 , n12385 , n19058 );
    or g25375 ( n27802 , n35927 , n10010 );
    and g25376 ( n4265 , n10330 , n34464 );
    xnor g25377 ( n7884 , n20311 , n7147 );
    nor g25378 ( n11732 , n8278 , n13757 );
    or g25379 ( n11232 , n12462 , n5965 );
    and g25380 ( n35318 , n758 , n11116 );
    not g25381 ( n13221 , n12141 );
    or g25382 ( n34279 , n15358 , n22316 );
    and g25383 ( n32676 , n6783 , n5962 );
    xnor g25384 ( n16818 , n29979 , n8580 );
    or g25385 ( n8095 , n28898 , n9268 );
    and g25386 ( n1296 , n15628 , n28402 );
    nor g25387 ( n17196 , n30268 , n30353 );
    xnor g25388 ( n31809 , n32970 , n8450 );
    xnor g25389 ( n17129 , n28684 , n10894 );
    or g25390 ( n6853 , n20936 , n31464 );
    xnor g25391 ( n34173 , n8425 , n27253 );
    and g25392 ( n19579 , n17106 , n17117 );
    and g25393 ( n20669 , n26164 , n24012 );
    or g25394 ( n3319 , n23901 , n17024 );
    or g25395 ( n19967 , n16723 , n21641 );
    or g25396 ( n27832 , n9846 , n15304 );
    or g25397 ( n3393 , n7838 , n30419 );
    or g25398 ( n9784 , n23604 , n4273 );
    nor g25399 ( n10673 , n9793 , n7637 );
    or g25400 ( n21347 , n4840 , n2384 );
    xnor g25401 ( n27127 , n1938 , n8928 );
    or g25402 ( n3933 , n13259 , n15805 );
    or g25403 ( n19134 , n28748 , n1762 );
    or g25404 ( n3411 , n4878 , n25172 );
    or g25405 ( n9473 , n35694 , n34971 );
    or g25406 ( n31888 , n4149 , n1997 );
    or g25407 ( n26014 , n9341 , n15145 );
    or g25408 ( n29745 , n35384 , n35757 );
    and g25409 ( n25340 , n22563 , n8962 );
    or g25410 ( n2296 , n3456 , n19403 );
    or g25411 ( n32211 , n23369 , n19464 );
    or g25412 ( n29284 , n19371 , n28438 );
    xnor g25413 ( n21816 , n20793 , n6748 );
    or g25414 ( n706 , n31799 , n23185 );
    and g25415 ( n31203 , n23889 , n17110 );
    and g25416 ( n21243 , n2355 , n5244 );
    or g25417 ( n24023 , n26846 , n16820 );
    or g25418 ( n23395 , n30112 , n12432 );
    or g25419 ( n1266 , n25174 , n15928 );
    and g25420 ( n9022 , n6676 , n30271 );
    xnor g25421 ( n6982 , n20216 , n3946 );
    and g25422 ( n17884 , n6056 , n16398 );
    or g25423 ( n23935 , n8247 , n10432 );
    nor g25424 ( n5164 , n33085 , n15202 );
    or g25425 ( n11998 , n19354 , n14246 );
    or g25426 ( n26971 , n1950 , n26703 );
    xnor g25427 ( n34358 , n25223 , n25686 );
    and g25428 ( n22954 , n3134 , n31637 );
    xnor g25429 ( n1598 , n17128 , n9789 );
    or g25430 ( n1257 , n24964 , n32808 );
    or g25431 ( n24794 , n24371 , n24415 );
    or g25432 ( n24031 , n8083 , n4639 );
    not g25433 ( n8211 , n15007 );
    xnor g25434 ( n13521 , n6663 , n11474 );
    or g25435 ( n31834 , n35097 , n20308 );
    or g25436 ( n32501 , n1950 , n1282 );
    xnor g25437 ( n24212 , n30066 , n14024 );
    and g25438 ( n5711 , n7927 , n2595 );
    or g25439 ( n6177 , n26256 , n2814 );
    or g25440 ( n29319 , n32095 , n8247 );
    or g25441 ( n26185 , n32449 , n7647 );
    or g25442 ( n26385 , n16922 , n8685 );
    or g25443 ( n16756 , n2719 , n3807 );
    xnor g25444 ( n29151 , n25788 , n32857 );
    nor g25445 ( n3267 , n17492 , n2912 );
    or g25446 ( n6631 , n5609 , n34865 );
    or g25447 ( n26061 , n19718 , n5868 );
    xnor g25448 ( n24015 , n10579 , n286 );
    and g25449 ( n24943 , n7421 , n18563 );
    xnor g25450 ( n10766 , n15375 , n947 );
    not g25451 ( n29804 , n23712 );
    and g25452 ( n8184 , n28858 , n21380 );
    or g25453 ( n1233 , n19434 , n5587 );
    or g25454 ( n5646 , n21454 , n965 );
    or g25455 ( n30574 , n31799 , n10407 );
    or g25456 ( n28861 , n11141 , n2078 );
    or g25457 ( n27974 , n4760 , n31249 );
    xnor g25458 ( n2985 , n5581 , n25418 );
    and g25459 ( n11381 , n8128 , n32729 );
    and g25460 ( n22413 , n28905 , n32926 );
    nor g25461 ( n4865 , n16242 , n33956 );
    or g25462 ( n9781 , n27939 , n22961 );
    or g25463 ( n23039 , n20329 , n19263 );
    or g25464 ( n14961 , n15257 , n30287 );
    and g25465 ( n30175 , n28116 , n7009 );
    not g25466 ( n17231 , n12575 );
    or g25467 ( n29702 , n32972 , n1411 );
    or g25468 ( n7031 , n36080 , n1132 );
    or g25469 ( n8920 , n31318 , n23976 );
    or g25470 ( n12283 , n14849 , n2955 );
    nor g25471 ( n17766 , n23604 , n13837 );
    or g25472 ( n15214 , n23387 , n26659 );
    and g25473 ( n18829 , n9756 , n33963 );
    nor g25474 ( n36044 , n1950 , n19133 );
    and g25475 ( n35449 , n22580 , n12196 );
    xnor g25476 ( n10050 , n20834 , n13978 );
    not g25477 ( n25351 , n9568 );
    or g25478 ( n22860 , n11667 , n9951 );
    and g25479 ( n29311 , n18715 , n29506 );
    or g25480 ( n16271 , n19551 , n17771 );
    buf g25481 ( n11977 , n341 );
    or g25482 ( n14888 , n2313 , n11440 );
    not g25483 ( n17618 , n2477 );
    xnor g25484 ( n13545 , n23008 , n27291 );
    or g25485 ( n4986 , n16419 , n13307 );
    and g25486 ( n3056 , n30262 , n15346 );
    and g25487 ( n1195 , n6619 , n31609 );
    not g25488 ( n28987 , n3480 );
    or g25489 ( n6519 , n1663 , n17782 );
    or g25490 ( n26997 , n19291 , n33416 );
    or g25491 ( n28167 , n10248 , n30672 );
    xnor g25492 ( n23004 , n23055 , n33292 );
    xnor g25493 ( n4243 , n26377 , n1177 );
    or g25494 ( n32534 , n4346 , n32632 );
    xnor g25495 ( n7611 , n10841 , n35756 );
    or g25496 ( n7082 , n30536 , n25592 );
    or g25497 ( n13865 , n4220 , n30481 );
    and g25498 ( n4892 , n11255 , n31658 );
    xnor g25499 ( n27717 , n22672 , n4962 );
    xnor g25500 ( n35136 , n13381 , n29110 );
    not g25501 ( n24177 , n22980 );
    and g25502 ( n33428 , n19944 , n30738 );
    and g25503 ( n15191 , n29528 , n3124 );
    or g25504 ( n8204 , n26313 , n19336 );
    or g25505 ( n10203 , n35778 , n25663 );
    xnor g25506 ( n24157 , n33395 , n26132 );
    or g25507 ( n30684 , n14980 , n3016 );
    or g25508 ( n26173 , n11837 , n14027 );
    xnor g25509 ( n22524 , n36014 , n8432 );
    or g25510 ( n24680 , n22558 , n14447 );
    or g25511 ( n829 , n19551 , n17633 );
    nor g25512 ( n24305 , n1890 , n18115 );
    or g25513 ( n12940 , n31557 , n11539 );
    not g25514 ( n35538 , n34300 );
    not g25515 ( n927 , n30742 );
    or g25516 ( n13156 , n27868 , n1715 );
    not g25517 ( n4895 , n11833 );
    or g25518 ( n24474 , n32284 , n23209 );
    and g25519 ( n23065 , n7517 , n34019 );
    not g25520 ( n4036 , n32071 );
    xnor g25521 ( n20073 , n35365 , n35026 );
    and g25522 ( n7755 , n306 , n29669 );
    or g25523 ( n2411 , n24844 , n18884 );
    or g25524 ( n7995 , n20041 , n33118 );
    or g25525 ( n2938 , n12152 , n26382 );
    or g25526 ( n27244 , n15464 , n27470 );
    or g25527 ( n29889 , n3428 , n19732 );
    or g25528 ( n34658 , n2837 , n32329 );
    or g25529 ( n18624 , n18867 , n6341 );
    or g25530 ( n5969 , n21372 , n3738 );
    and g25531 ( n8909 , n15113 , n16730 );
    or g25532 ( n33306 , n10021 , n10336 );
    or g25533 ( n28017 , n27361 , n17872 );
    xnor g25534 ( n33774 , n605 , n31631 );
    xnor g25535 ( n34313 , n1757 , n9793 );
    or g25536 ( n12009 , n31289 , n14444 );
    or g25537 ( n29747 , n9804 , n19732 );
    or g25538 ( n19680 , n25174 , n22972 );
    or g25539 ( n14939 , n4400 , n11601 );
    or g25540 ( n20645 , n16922 , n12678 );
    or g25541 ( n16196 , n10628 , n25999 );
    and g25542 ( n4445 , n8112 , n6230 );
    xnor g25543 ( n6027 , n2657 , n9658 );
    nor g25544 ( n24567 , n24621 , n1763 );
    or g25545 ( n2116 , n23926 , n7443 );
    not g25546 ( n19314 , n26283 );
    or g25547 ( n27557 , n14324 , n241 );
    and g25548 ( n1634 , n30946 , n26043 );
    or g25549 ( n17211 , n9279 , n10289 );
    xnor g25550 ( n33715 , n11740 , n15255 );
    or g25551 ( n23975 , n26224 , n3188 );
    xnor g25552 ( n20107 , n7688 , n25323 );
    and g25553 ( n34621 , n19082 , n31858 );
    or g25554 ( n1561 , n32431 , n19173 );
    or g25555 ( n2049 , n4969 , n16464 );
    nor g25556 ( n17582 , n26268 , n13141 );
    nor g25557 ( n27541 , n31002 , n20428 );
    or g25558 ( n13730 , n17751 , n32535 );
    or g25559 ( n32886 , n32375 , n34727 );
    and g25560 ( n21999 , n34293 , n24660 );
    or g25561 ( n26229 , n32675 , n4142 );
    xnor g25562 ( n28624 , n18567 , n15299 );
    or g25563 ( n22240 , n31559 , n22246 );
    or g25564 ( n35656 , n31082 , n21704 );
    and g25565 ( n19998 , n28600 , n16101 );
    not g25566 ( n13976 , n7540 );
    or g25567 ( n5573 , n20174 , n26023 );
    and g25568 ( n16717 , n11973 , n33862 );
    nor g25569 ( n27915 , n32584 , n28219 );
    not g25570 ( n8844 , n1950 );
    xnor g25571 ( n34109 , n23740 , n27291 );
    and g25572 ( n34043 , n1198 , n28822 );
    or g25573 ( n35661 , n12136 , n17354 );
    or g25574 ( n13538 , n31056 , n12894 );
    and g25575 ( n2684 , n22537 , n17935 );
    xnor g25576 ( n12558 , n5580 , n5335 );
    or g25577 ( n36001 , n8274 , n18477 );
    or g25578 ( n25483 , n30542 , n27580 );
    xnor g25579 ( n12483 , n32088 , n15886 );
    and g25580 ( n632 , n21607 , n15465 );
    or g25581 ( n26147 , n6189 , n11849 );
    or g25582 ( n33318 , n23959 , n18255 );
    not g25583 ( n16607 , n737 );
    and g25584 ( n17802 , n20684 , n32004 );
    or g25585 ( n8195 , n32900 , n27580 );
    or g25586 ( n21198 , n22866 , n26891 );
    or g25587 ( n20168 , n4955 , n14285 );
    xnor g25588 ( n8168 , n35489 , n18961 );
    xnor g25589 ( n23461 , n11925 , n32095 );
    or g25590 ( n5480 , n31799 , n18266 );
    xnor g25591 ( n4226 , n35767 , n12046 );
    xnor g25592 ( n9354 , n32190 , n26174 );
    not g25593 ( n19766 , n11234 );
    buf g25594 ( n25761 , n6977 );
    or g25595 ( n1442 , n30279 , n7669 );
    or g25596 ( n16545 , n1452 , n16659 );
    or g25597 ( n25716 , n34701 , n25592 );
    or g25598 ( n17329 , n22405 , n27728 );
    not g25599 ( n35100 , n28746 );
    nor g25600 ( n19931 , n1463 , n23148 );
    xnor g25601 ( n30128 , n34231 , n10533 );
    and g25602 ( n13158 , n3952 , n26012 );
    xnor g25603 ( n18782 , n21722 , n34804 );
    xnor g25604 ( n17747 , n9238 , n4962 );
    xnor g25605 ( n9525 , n9692 , n7348 );
    xnor g25606 ( n26232 , n25373 , n4960 );
    and g25607 ( n23621 , n678 , n18319 );
    xnor g25608 ( n20174 , n8290 , n18101 );
    xnor g25609 ( n35193 , n16936 , n7578 );
    and g25610 ( n33405 , n27410 , n27349 );
    or g25611 ( n16252 , n12225 , n4556 );
    or g25612 ( n33134 , n16759 , n30779 );
    xnor g25613 ( n14343 , n19518 , n3096 );
    not g25614 ( n32731 , n25338 );
    xnor g25615 ( n16025 , n10997 , n32095 );
    or g25616 ( n25781 , n15403 , n16180 );
    or g25617 ( n33228 , n17568 , n22701 );
    xnor g25618 ( n20392 , n330 , n3946 );
    and g25619 ( n23593 , n711 , n29211 );
    xnor g25620 ( n9676 , n2226 , n24781 );
    or g25621 ( n31934 , n25665 , n277 );
    or g25622 ( n3462 , n8323 , n30204 );
    nor g25623 ( n12585 , n12406 , n10038 );
    not g25624 ( n29349 , n29104 );
    nor g25625 ( n19419 , n1950 , n14209 );
    or g25626 ( n31309 , n29558 , n30898 );
    or g25627 ( n6326 , n2456 , n20902 );
    and g25628 ( n20654 , n5531 , n10947 );
    nor g25629 ( n30113 , n1950 , n30994 );
    nor g25630 ( n5303 , n25174 , n2352 );
    xnor g25631 ( n32714 , n21636 , n12481 );
    or g25632 ( n26215 , n6231 , n3774 );
    not g25633 ( n6513 , n15660 );
    or g25634 ( n31430 , n14280 , n10872 );
    and g25635 ( n6258 , n19400 , n31524 );
    nor g25636 ( n26768 , n9740 , n9921 );
    or g25637 ( n19094 , n19984 , n7987 );
    and g25638 ( n22597 , n22973 , n433 );
    nor g25639 ( n2997 , n19439 , n12913 );
    or g25640 ( n14307 , n34491 , n13217 );
    or g25641 ( n35697 , n29870 , n702 );
    or g25642 ( n33653 , n29476 , n11458 );
    and g25643 ( n1586 , n7676 , n19424 );
    not g25644 ( n2380 , n4544 );
    or g25645 ( n24181 , n22567 , n21977 );
    xnor g25646 ( n3055 , n30161 , n10894 );
    and g25647 ( n24229 , n17366 , n14515 );
    or g25648 ( n1493 , n16620 , n21088 );
    xnor g25649 ( n18520 , n10494 , n16727 );
    or g25650 ( n3869 , n32277 , n17872 );
    or g25651 ( n2669 , n23315 , n24356 );
    xnor g25652 ( n23766 , n22906 , n34236 );
    or g25653 ( n29554 , n16922 , n15890 );
    or g25654 ( n9619 , n23586 , n22611 );
    or g25655 ( n26167 , n22193 , n4478 );
    or g25656 ( n31593 , n9596 , n5874 );
    or g25657 ( n32990 , n4962 , n3532 );
    not g25658 ( n24261 , n16620 );
    xnor g25659 ( n34847 , n11713 , n3222 );
    xnor g25660 ( n27736 , n5241 , n29039 );
    nor g25661 ( n9916 , n18932 , n30463 );
    or g25662 ( n30266 , n15062 , n35043 );
    or g25663 ( n19533 , n35927 , n15495 );
    or g25664 ( n26829 , n3835 , n9731 );
    xnor g25665 ( n19073 , n16528 , n33328 );
    or g25666 ( n30750 , n32509 , n28493 );
    or g25667 ( n27287 , n3205 , n24339 );
    not g25668 ( n11773 , n15290 );
    or g25669 ( n21199 , n31202 , n21977 );
    and g25670 ( n11252 , n15670 , n26925 );
    or g25671 ( n4039 , n27757 , n22241 );
    nor g25672 ( n24351 , n2467 , n31184 );
    or g25673 ( n19582 , n24371 , n19071 );
    and g25674 ( n150 , n25818 , n32475 );
    or g25675 ( n11408 , n17307 , n2817 );
    and g25676 ( n22939 , n25000 , n9917 );
    or g25677 ( n31074 , n18864 , n19952 );
    or g25678 ( n26249 , n5335 , n12886 );
    and g25679 ( n28014 , n21568 , n2604 );
    and g25680 ( n11234 , n15175 , n28914 );
    or g25681 ( n2212 , n18252 , n31939 );
    xnor g25682 ( n20209 , n9543 , n19551 );
    or g25683 ( n19801 , n3372 , n27801 );
    or g25684 ( n27264 , n21484 , n30483 );
    nor g25685 ( n8245 , n10743 , n24753 );
    or g25686 ( n35462 , n32857 , n15085 );
    not g25687 ( n23755 , n16620 );
    or g25688 ( n6593 , n4288 , n25422 );
    and g25689 ( n18593 , n29114 , n6221 );
    or g25690 ( n35165 , n16561 , n25841 );
    or g25691 ( n28377 , n33995 , n14554 );
    and g25692 ( n2939 , n5453 , n3142 );
    xnor g25693 ( n32349 , n35494 , n32857 );
    or g25694 ( n13640 , n18383 , n14699 );
    and g25695 ( n5301 , n30889 , n11573 );
    or g25696 ( n29426 , n27291 , n17957 );
    or g25697 ( n34007 , n20556 , n22788 );
    or g25698 ( n1794 , n4878 , n31624 );
    xnor g25699 ( n14324 , n16479 , n31289 );
    not g25700 ( n9928 , n22501 );
    xnor g25701 ( n35431 , n10943 , n5335 );
    buf g25702 ( n25648 , n6560 );
    not g25703 ( n11757 , n22767 );
    or g25704 ( n7979 , n13565 , n22206 );
    or g25705 ( n20208 , n24371 , n24222 );
    nor g25706 ( n4499 , n29839 , n214 );
    not g25707 ( n8538 , n4960 );
    and g25708 ( n34381 , n29168 , n35768 );
    not g25709 ( n11035 , n4240 );
    or g25710 ( n21363 , n16694 , n16456 );
    xnor g25711 ( n21636 , n16261 , n24332 );
    and g25712 ( n9523 , n9302 , n28161 );
    and g25713 ( n767 , n16171 , n17291 );
    and g25714 ( n35598 , n29401 , n10019 );
    xnor g25715 ( n27190 , n17332 , n26866 );
    or g25716 ( n34954 , n25057 , n10960 );
    xnor g25717 ( n24978 , n13139 , n14950 );
    not g25718 ( n3663 , n18448 );
    nor g25719 ( n5925 , n30777 , n79 );
    or g25720 ( n21766 , n23309 , n17438 );
    and g25721 ( n29444 , n31266 , n563 );
    and g25722 ( n25545 , n6594 , n33343 );
    xnor g25723 ( n31806 , n5839 , n8766 );
    xnor g25724 ( n26574 , n19645 , n20957 );
    or g25725 ( n16439 , n30285 , n35784 );
    or g25726 ( n26523 , n10777 , n25447 );
    nor g25727 ( n9346 , n32584 , n21869 );
    or g25728 ( n33270 , n22621 , n13215 );
    xnor g25729 ( n30749 , n34553 , n4557 );
    or g25730 ( n6419 , n9076 , n14798 );
    or g25731 ( n27006 , n12742 , n15202 );
    and g25732 ( n8313 , n34071 , n18243 );
    or g25733 ( n33851 , n30254 , n26002 );
    or g25734 ( n12525 , n12594 , n21787 );
    xnor g25735 ( n39 , n35970 , n34884 );
    and g25736 ( n30825 , n19525 , n1266 );
    xnor g25737 ( n35286 , n18796 , n20958 );
    or g25738 ( n18479 , n11814 , n9030 );
    and g25739 ( n31632 , n34574 , n28664 );
    xnor g25740 ( n26005 , n11010 , n1950 );
    or g25741 ( n15746 , n4878 , n28882 );
    xnor g25742 ( n11435 , n5074 , n33625 );
    nor g25743 ( n18367 , n5287 , n12494 );
    and g25744 ( n31955 , n8051 , n33273 );
    and g25745 ( n17859 , n30582 , n23431 );
    or g25746 ( n20889 , n10894 , n6215 );
    or g25747 ( n15121 , n22065 , n21042 );
    or g25748 ( n33953 , n5287 , n5020 );
    or g25749 ( n12977 , n33485 , n6459 );
    or g25750 ( n34579 , n32095 , n5115 );
    nor g25751 ( n2171 , n3205 , n28 );
    or g25752 ( n20984 , n3205 , n17300 );
    xnor g25753 ( n21829 , n14959 , n27391 );
    xnor g25754 ( n25613 , n9145 , n5720 );
    and g25755 ( n20852 , n36089 , n5108 );
    xnor g25756 ( n17548 , n29163 , n24371 );
    or g25757 ( n22790 , n35321 , n21550 );
    xnor g25758 ( n10988 , n11487 , n11046 );
    not g25759 ( n10982 , n16620 );
    and g25760 ( n32135 , n22064 , n32759 );
    and g25761 ( n19248 , n20898 , n14349 );
    and g25762 ( n20546 , n17999 , n20505 );
    or g25763 ( n8451 , n32855 , n17604 );
    or g25764 ( n9969 , n35568 , n12752 );
    or g25765 ( n4340 , n16620 , n13529 );
    xnor g25766 ( n7255 , n1220 , n28591 );
    or g25767 ( n10947 , n31559 , n19976 );
    nor g25768 ( n17873 , n9260 , n33956 );
    or g25769 ( n2288 , n32129 , n14076 );
    not g25770 ( n21839 , n7357 );
    or g25771 ( n9178 , n11492 , n18005 );
    and g25772 ( n22448 , n25246 , n29904 );
    xnor g25773 ( n1888 , n5118 , n4960 );
    nor g25774 ( n7397 , n4962 , n19800 );
    or g25775 ( n31170 , n29713 , n33875 );
    xnor g25776 ( n34337 , n33166 , n9811 );
    xnor g25777 ( n4900 , n18868 , n16294 );
    and g25778 ( n21318 , n17279 , n33755 );
    or g25779 ( n17735 , n198 , n26292 );
    or g25780 ( n1038 , n11790 , n20812 );
    xnor g25781 ( n16617 , n30934 , n15194 );
    or g25782 ( n12211 , n35927 , n18601 );
    or g25783 ( n8291 , n16667 , n24093 );
    or g25784 ( n35626 , n15502 , n21780 );
    and g25785 ( n14759 , n461 , n11811 );
    and g25786 ( n22899 , n3843 , n35788 );
    nor g25787 ( n25855 , n19418 , n17668 );
    or g25788 ( n11777 , n4878 , n17842 );
    not g25789 ( n862 , n14501 );
    xnor g25790 ( n21847 , n21523 , n25695 );
    xnor g25791 ( n19392 , n32336 , n1458 );
    or g25792 ( n29678 , n5194 , n17060 );
    or g25793 ( n20731 , n34121 , n35038 );
    or g25794 ( n30814 , n22466 , n17572 );
    xnor g25795 ( n32970 , n12813 , n23604 );
    and g25796 ( n21759 , n29086 , n13061 );
    not g25797 ( n6760 , n21287 );
    or g25798 ( n24149 , n13280 , n2127 );
    nor g25799 ( n4596 , n30742 , n23307 );
    and g25800 ( n20440 , n16210 , n15965 );
    xnor g25801 ( n943 , n13848 , n12553 );
    or g25802 ( n18715 , n7762 , n8392 );
    and g25803 ( n13302 , n32550 , n9233 );
    xnor g25804 ( n7912 , n33976 , n15782 );
    and g25805 ( n8434 , n35526 , n3855 );
    xnor g25806 ( n26207 , n23312 , n27226 );
    and g25807 ( n1978 , n3334 , n25063 );
    not g25808 ( n433 , n14747 );
    nor g25809 ( n6550 , n15261 , n32128 );
    or g25810 ( n35117 , n34796 , n27625 );
    xnor g25811 ( n26559 , n29428 , n34675 );
    and g25812 ( n5048 , n36052 , n20761 );
    xnor g25813 ( n34221 , n28628 , n18269 );
    or g25814 ( n29811 , n9516 , n27418 );
    xnor g25815 ( n5344 , n408 , n10176 );
    or g25816 ( n15324 , n33442 , n2556 );
    xnor g25817 ( n29593 , n9718 , n18855 );
    and g25818 ( n20515 , n22862 , n10729 );
    xnor g25819 ( n21775 , n14739 , n4758 );
    or g25820 ( n7699 , n23762 , n7647 );
    or g25821 ( n1621 , n30573 , n8293 );
    and g25822 ( n9950 , n10610 , n3306 );
    xnor g25823 ( n10748 , n33044 , n15886 );
    nor g25824 ( n17745 , n10587 , n21135 );
    or g25825 ( n22680 , n7907 , n30204 );
    xnor g25826 ( n17784 , n32935 , n23604 );
    and g25827 ( n34268 , n31260 , n9712 );
    or g25828 ( n6810 , n21099 , n544 );
    xnor g25829 ( n34597 , n23583 , n15921 );
    nor g25830 ( n371 , n24332 , n19977 );
    and g25831 ( n19861 , n23174 , n9415 );
    or g25832 ( n25178 , n77 , n20805 );
    or g25833 ( n20078 , n879 , n19952 );
    xnor g25834 ( n29520 , n30175 , n32095 );
    nor g25835 ( n4821 , n33456 , n26109 );
    and g25836 ( n11577 , n12875 , n7097 );
    or g25837 ( n29869 , n31751 , n4718 );
    or g25838 ( n24291 , n228 , n7293 );
    nor g25839 ( n34097 , n26878 , n13390 );
    or g25840 ( n24770 , n10983 , n1278 );
    and g25841 ( n19034 , n17653 , n20431 );
    and g25842 ( n13106 , n27329 , n34859 );
    xnor g25843 ( n23394 , n2953 , n1026 );
    xnor g25844 ( n9184 , n12363 , n9793 );
    or g25845 ( n13143 , n34894 , n33896 );
    and g25846 ( n4488 , n26497 , n28495 );
    nor g25847 ( n1381 , n31289 , n580 );
    buf g25848 ( n9030 , n15233 );
    or g25849 ( n15041 , n32715 , n7347 );
    or g25850 ( n3804 , n16620 , n14418 );
    xnor g25851 ( n18559 , n25020 , n12798 );
    xnor g25852 ( n13331 , n12816 , n31227 );
    not g25853 ( n30751 , n19939 );
    or g25854 ( n7400 , n11190 , n3174 );
    or g25855 ( n3945 , n22291 , n29557 );
    not g25856 ( n3513 , n35466 );
    xnor g25857 ( n4766 , n11144 , n10894 );
    or g25858 ( n23140 , n22955 , n7271 );
    or g25859 ( n12975 , n25174 , n15240 );
    or g25860 ( n11288 , n28695 , n12950 );
    or g25861 ( n25691 , n21255 , n33271 );
    or g25862 ( n22897 , n18343 , n11977 );
    xnor g25863 ( n17522 , n22020 , n481 );
    or g25864 ( n13273 , n31183 , n13869 );
    and g25865 ( n17141 , n22039 , n27045 );
    or g25866 ( n18420 , n31056 , n33060 );
    or g25867 ( n20575 , n20815 , n3858 );
    xnor g25868 ( n17655 , n10629 , n194 );
    and g25869 ( n22494 , n17777 , n24886 );
    xnor g25870 ( n35797 , n22637 , n9789 );
    or g25871 ( n31009 , n31267 , n25164 );
    xnor g25872 ( n2019 , n8819 , n31718 );
    xnor g25873 ( n15294 , n15800 , n8432 );
    and g25874 ( n26508 , n26279 , n12613 );
    or g25875 ( n5935 , n5187 , n31563 );
    xnor g25876 ( n21827 , n35397 , n34273 );
    and g25877 ( n3556 , n455 , n20928 );
    or g25878 ( n8731 , n12120 , n15831 );
    and g25879 ( n23890 , n17238 , n12579 );
    or g25880 ( n13723 , n20613 , n22408 );
    or g25881 ( n493 , n33094 , n9951 );
    or g25882 ( n9841 , n33567 , n34656 );
    or g25883 ( n30487 , n3116 , n19125 );
    or g25884 ( n13739 , n10894 , n18383 );
    or g25885 ( n22219 , n21688 , n15496 );
    and g25886 ( n17577 , n30174 , n11007 );
    and g25887 ( n24792 , n34181 , n19948 );
    and g25888 ( n34249 , n2210 , n13178 );
    xnor g25889 ( n33981 , n7917 , n15899 );
    or g25890 ( n24175 , n21806 , n10345 );
    xnor g25891 ( n35833 , n27831 , n4758 );
    and g25892 ( n15267 , n13095 , n16410 );
    xnor g25893 ( n17613 , n2596 , n12710 );
    and g25894 ( n19934 , n25395 , n10646 );
    or g25895 ( n29446 , n798 , n23776 );
    xnor g25896 ( n8875 , n21355 , n22970 );
    and g25897 ( n7792 , n12700 , n23448 );
    or g25898 ( n31995 , n2985 , n17872 );
    or g25899 ( n28293 , n5022 , n14918 );
    or g25900 ( n10414 , n21088 , n4772 );
    or g25901 ( n12738 , n12955 , n19173 );
    and g25902 ( n29054 , n15202 , n22189 );
    nor g25903 ( n29974 , n4962 , n28247 );
    xnor g25904 ( n13864 , n23880 , n263 );
    and g25905 ( n1606 , n18179 , n13311 );
    nor g25906 ( n29130 , n32180 , n31946 );
    and g25907 ( n34152 , n27634 , n16204 );
    not g25908 ( n24651 , n4288 );
    and g25909 ( n12391 , n13038 , n28602 );
    or g25910 ( n15159 , n12276 , n16486 );
    or g25911 ( n21035 , n18689 , n4254 );
    or g25912 ( n9040 , n29776 , n31253 );
    and g25913 ( n34356 , n22220 , n27810 );
    nor g25914 ( n4792 , n22497 , n8266 );
    and g25915 ( n31354 , n1604 , n13573 );
    and g25916 ( n10625 , n28263 , n33994 );
    or g25917 ( n25242 , n31289 , n5719 );
    nor g25918 ( n21324 , n25602 , n35204 );
    nor g25919 ( n34776 , n30742 , n34894 );
    or g25920 ( n8602 , n9310 , n18811 );
    or g25921 ( n10237 , n15011 , n6831 );
    and g25922 ( n5684 , n31894 , n34104 );
    and g25923 ( n31069 , n17617 , n8030 );
    xnor g25924 ( n18431 , n1094 , n20540 );
    not g25925 ( n8365 , n3884 );
    or g25926 ( n22441 , n33853 , n7293 );
    xnor g25927 ( n28335 , n17802 , n31799 );
    or g25928 ( n13816 , n15143 , n6459 );
    and g25929 ( n16606 , n9337 , n30019 );
    or g25930 ( n12757 , n23430 , n30893 );
    or g25931 ( n22718 , n3222 , n22336 );
    or g25932 ( n4049 , n22273 , n9579 );
    not g25933 ( n597 , n23786 );
    xnor g25934 ( n21615 , n6556 , n15886 );
    xnor g25935 ( n4813 , n23307 , n22281 );
    and g25936 ( n9629 , n30723 , n29293 );
    or g25937 ( n13784 , n28557 , n12649 );
    and g25938 ( n5635 , n11601 , n303 );
    xnor g25939 ( n10256 , n14099 , n9793 );
    or g25940 ( n10152 , n15054 , n25648 );
    or g25941 ( n23042 , n35260 , n2005 );
    xnor g25942 ( n4797 , n32248 , n24745 );
    nor g25943 ( n35232 , n29839 , n21169 );
    xnor g25944 ( n20400 , n4833 , n24176 );
    and g25945 ( n35937 , n9107 , n30678 );
    or g25946 ( n552 , n10792 , n19076 );
    or g25947 ( n1721 , n25174 , n17448 );
    and g25948 ( n19368 , n1283 , n27814 );
    or g25949 ( n6256 , n8975 , n15538 );
    or g25950 ( n6637 , n7499 , n11985 );
    xnor g25951 ( n14270 , n7396 , n5941 );
    xnor g25952 ( n19549 , n31841 , n9079 );
    or g25953 ( n13370 , n22958 , n20024 );
    or g25954 ( n15764 , n29599 , n21956 );
    and g25955 ( n10287 , n22349 , n1894 );
    not g25956 ( n2056 , n31559 );
    and g25957 ( n33198 , n23876 , n1766 );
    or g25958 ( n10453 , n3907 , n2168 );
    and g25959 ( n31283 , n27088 , n4689 );
    or g25960 ( n28689 , n18658 , n2340 );
    not g25961 ( n2409 , n14456 );
    or g25962 ( n33365 , n16000 , n35935 );
    or g25963 ( n34340 , n6670 , n14315 );
    xnor g25964 ( n8583 , n16954 , n32913 );
    and g25965 ( n18426 , n18809 , n4605 );
    nor g25966 ( n23290 , n4878 , n23658 );
    or g25967 ( n23530 , n5163 , n2117 );
    xnor g25968 ( n32748 , n21373 , n32584 );
    and g25969 ( n22799 , n11669 , n34872 );
    or g25970 ( n30170 , n32715 , n18689 );
    or g25971 ( n20128 , n29713 , n5187 );
    xnor g25972 ( n26619 , n34595 , n22519 );
    nor g25973 ( n1924 , n17119 , n4508 );
    not g25974 ( n26565 , n31799 );
    or g25975 ( n11347 , n17869 , n20762 );
    or g25976 ( n20288 , n30742 , n3263 );
    and g25977 ( n18887 , n20622 , n27157 );
    and g25978 ( n23809 , n33907 , n1597 );
    or g25979 ( n1286 , n28446 , n8282 );
    buf g25980 ( n34971 , n1942 );
    xnor g25981 ( n15819 , n10214 , n3483 );
    or g25982 ( n3238 , n16922 , n33049 );
    or g25983 ( n16648 , n17058 , n34898 );
    or g25984 ( n31805 , n14813 , n5598 );
    and g25985 ( n14983 , n31671 , n26064 );
    xnor g25986 ( n18765 , n25 , n23319 );
    and g25987 ( n12867 , n31971 , n15364 );
    not g25988 ( n14612 , n30742 );
    or g25989 ( n15326 , n32584 , n24040 );
    and g25990 ( n34413 , n4295 , n540 );
    and g25991 ( n34922 , n34387 , n32175 );
    xnor g25992 ( n25232 , n34612 , n9022 );
    not g25993 ( n29220 , n22907 );
    or g25994 ( n22764 , n22244 , n14918 );
    or g25995 ( n11884 , n3530 , n4952 );
    or g25996 ( n24736 , n32857 , n24940 );
    nor g25997 ( n34639 , n21738 , n25127 );
    nor g25998 ( n24818 , n23604 , n11740 );
    not g25999 ( n21651 , n23604 );
    or g26000 ( n32001 , n510 , n18409 );
    nor g26001 ( n20428 , n28514 , n31186 );
    or g26002 ( n937 , n20147 , n30549 );
    xnor g26003 ( n5746 , n4975 , n32857 );
    and g26004 ( n341 , n6380 , n5332 );
    or g26005 ( n9408 , n17568 , n19860 );
    and g26006 ( n4779 , n18945 , n32914 );
    xnor g26007 ( n27685 , n34994 , n11974 );
    xnor g26008 ( n32863 , n13123 , n25174 );
    or g26009 ( n34817 , n16341 , n33098 );
    or g26010 ( n26252 , n32590 , n28064 );
    and g26011 ( n27853 , n32014 , n29189 );
    xnor g26012 ( n8083 , n28962 , n31056 );
    and g26013 ( n2387 , n15367 , n13102 );
    or g26014 ( n32242 , n26271 , n31055 );
    xnor g26015 ( n31874 , n31114 , n32095 );
    and g26016 ( n12618 , n5295 , n34023 );
    not g26017 ( n16979 , n29327 );
    or g26018 ( n7512 , n15984 , n7926 );
    nor g26019 ( n24296 , n17751 , n11225 );
    nor g26020 ( n8059 , n25602 , n8985 );
    xnor g26021 ( n16623 , n33096 , n16463 );
    or g26022 ( n31870 , n22291 , n31782 );
    and g26023 ( n10300 , n5314 , n20864 );
    not g26024 ( n35441 , n34510 );
    nor g26025 ( n7136 , n32857 , n2128 );
    xnor g26026 ( n15261 , n34385 , n3207 );
    and g26027 ( n7692 , n35799 , n18276 );
    or g26028 ( n29572 , n20977 , n2955 );
    not g26029 ( n35027 , n31277 );
    or g26030 ( n2659 , n30695 , n19084 );
    not g26031 ( n3091 , n35927 );
    and g26032 ( n966 , n12676 , n3934 );
    or g26033 ( n34120 , n23906 , n12996 );
    xnor g26034 ( n26601 , n2886 , n16299 );
    xnor g26035 ( n8608 , n5162 , n31401 );
    xnor g26036 ( n8647 , n14797 , n20091 );
    or g26037 ( n30272 , n641 , n21042 );
    or g26038 ( n20056 , n9589 , n16456 );
    or g26039 ( n26853 , n18235 , n4772 );
    nor g26040 ( n5554 , n17568 , n7479 );
    or g26041 ( n26920 , n32341 , n16875 );
    xnor g26042 ( n16563 , n32020 , n5335 );
    not g26043 ( n27902 , n32699 );
    and g26044 ( n34086 , n3253 , n22146 );
    or g26045 ( n6277 , n33056 , n25773 );
    nor g26046 ( n27727 , n18699 , n115 );
    not g26047 ( n8701 , n9793 );
    and g26048 ( n1421 , n9157 , n18451 );
    buf g26049 ( n7448 , n6017 );
    nor g26050 ( n4386 , n12078 , n31411 );
    and g26051 ( n26109 , n10144 , n6611 );
    nor g26052 ( n13947 , n32095 , n3028 );
    not g26053 ( n15835 , n28273 );
    xnor g26054 ( n22978 , n3536 , n30200 );
    or g26055 ( n3881 , n33641 , n1051 );
    not g26056 ( n21810 , n1629 );
    or g26057 ( n7989 , n18504 , n3405 );
    or g26058 ( n22469 , n4405 , n16543 );
    xnor g26059 ( n30116 , n35962 , n23101 );
    and g26060 ( n31282 , n25714 , n26753 );
    or g26061 ( n10773 , n3939 , n25761 );
    xnor g26062 ( n23336 , n9895 , n32991 );
    or g26063 ( n11003 , n22123 , n4772 );
    and g26064 ( n24538 , n6745 , n26735 );
    not g26065 ( n16697 , n31474 );
    xnor g26066 ( n6667 , n2863 , n5335 );
    or g26067 ( n27509 , n3109 , n3466 );
    and g26068 ( n5223 , n6117 , n12846 );
    or g26069 ( n21825 , n28903 , n4546 );
    or g26070 ( n28112 , n10418 , n29626 );
    or g26071 ( n21843 , n4758 , n32385 );
    or g26072 ( n29051 , n569 , n31773 );
    xnor g26073 ( n11514 , n22690 , n927 );
    and g26074 ( n28728 , n14157 , n2391 );
    xnor g26075 ( n25376 , n19071 , n24371 );
    xnor g26076 ( n25324 , n12782 , n11455 );
    or g26077 ( n28038 , n26868 , n25592 );
    or g26078 ( n5755 , n10997 , n26365 );
    not g26079 ( n10147 , n23186 );
    or g26080 ( n34136 , n14107 , n18811 );
    xnor g26081 ( n20766 , n30557 , n10166 );
    or g26082 ( n80 , n31792 , n30431 );
    or g26083 ( n32010 , n19064 , n8324 );
    xnor g26084 ( n20942 , n5024 , n3514 );
    or g26085 ( n31974 , n2447 , n33969 );
    or g26086 ( n26401 , n15639 , n29220 );
    xnor g26087 ( n24880 , n14829 , n9568 );
    or g26088 ( n15245 , n5335 , n19930 );
    nor g26089 ( n29587 , n17665 , n28867 );
    and g26090 ( n20441 , n8810 , n26816 );
    and g26091 ( n27502 , n10457 , n12371 );
    xnor g26092 ( n30718 , n4920 , n21320 );
    and g26093 ( n28873 , n13070 , n25362 );
    xnor g26094 ( n20947 , n11855 , n12654 );
    and g26095 ( n1616 , n5526 , n25676 );
    or g26096 ( n4383 , n20191 , n34923 );
    or g26097 ( n16868 , n28610 , n12950 );
    and g26098 ( n14232 , n16439 , n11566 );
    and g26099 ( n33471 , n31007 , n20410 );
    xnor g26100 ( n11465 , n1944 , n12823 );
    and g26101 ( n1625 , n12373 , n15093 );
    and g26102 ( n14215 , n7603 , n13483 );
    xnor g26103 ( n7971 , n24948 , n35693 );
    nor g26104 ( n33610 , n16620 , n32061 );
    buf g26105 ( n3756 , n32071 );
    or g26106 ( n33971 , n1965 , n34727 );
    xnor g26107 ( n3036 , n6629 , n19551 );
    not g26108 ( n7834 , n11307 );
    or g26109 ( n26141 , n30113 , n22899 );
    not g26110 ( n17861 , n33435 );
    xnor g26111 ( n34050 , n8088 , n10894 );
    not g26112 ( n14351 , n22180 );
    nor g26113 ( n5930 , n16620 , n25679 );
    or g26114 ( n4799 , n15957 , n10882 );
    and g26115 ( n19097 , n21885 , n17520 );
    or g26116 ( n29606 , n34313 , n4264 );
    or g26117 ( n22957 , n33173 , n8392 );
    or g26118 ( n5087 , n32052 , n34427 );
    or g26119 ( n8826 , n20158 , n23157 );
    and g26120 ( n24613 , n294 , n19303 );
    and g26121 ( n5477 , n23938 , n4376 );
    or g26122 ( n29697 , n19184 , n31464 );
    xnor g26123 ( n1747 , n33538 , n7288 );
    or g26124 ( n16792 , n17082 , n27053 );
    or g26125 ( n20810 , n19551 , n28208 );
    or g26126 ( n22835 , n11455 , n23080 );
    xnor g26127 ( n21881 , n9827 , n3946 );
    not g26128 ( n912 , n23604 );
    xnor g26129 ( n30100 , n22268 , n1950 );
    and g26130 ( n26473 , n29063 , n6080 );
    nor g26131 ( n11614 , n4758 , n30468 );
    and g26132 ( n25663 , n10700 , n20580 );
    xnor g26133 ( n13822 , n7387 , n1465 );
    and g26134 ( n12816 , n4068 , n872 );
    or g26135 ( n14191 , n29713 , n23212 );
    xnor g26136 ( n2964 , n25245 , n24788 );
    and g26137 ( n11825 , n25919 , n2032 );
    or g26138 ( n28268 , n13462 , n4254 );
    or g26139 ( n11011 , n33765 , n30751 );
    xnor g26140 ( n29989 , n14634 , n746 );
    xnor g26141 ( n35707 , n27820 , n1950 );
    or g26142 ( n4181 , n16620 , n20815 );
    xnor g26143 ( n30597 , n30256 , n14386 );
    not g26144 ( n33888 , n10895 );
    xnor g26145 ( n33869 , n6116 , n27080 );
    or g26146 ( n2614 , n5301 , n18255 );
    xnor g26147 ( n12007 , n13734 , n6259 );
    xnor g26148 ( n16628 , n7018 , n20897 );
    xnor g26149 ( n21350 , n9980 , n27160 );
    nor g26150 ( n21725 , n35121 , n6017 );
    xnor g26151 ( n20501 , n2909 , n11924 );
    xnor g26152 ( n8696 , n9831 , n17568 );
    not g26153 ( n14698 , n5606 );
    nor g26154 ( n33086 , n4574 , n1701 );
    and g26155 ( n1525 , n31511 , n23458 );
    or g26156 ( n14177 , n9175 , n14313 );
    buf g26157 ( n10960 , n2666 );
    nor g26158 ( n4647 , n27226 , n16930 );
    or g26159 ( n7211 , n33183 , n34621 );
    or g26160 ( n13765 , n11046 , n32446 );
    or g26161 ( n9144 , n23971 , n35547 );
    xnor g26162 ( n6311 , n1302 , n14322 );
    or g26163 ( n21577 , n3854 , n27011 );
    or g26164 ( n21854 , n830 , n20760 );
    or g26165 ( n18021 , n5044 , n34537 );
    and g26166 ( n18196 , n13838 , n3772 );
    and g26167 ( n16893 , n6523 , n864 );
    and g26168 ( n20340 , n26786 , n18957 );
    and g26169 ( n9010 , n4533 , n9497 );
    or g26170 ( n33727 , n30936 , n26480 );
    or g26171 ( n30797 , n17026 , n17405 );
    xnor g26172 ( n30622 , n29792 , n12477 );
    nor g26173 ( n5548 , n3205 , n6297 );
    or g26174 ( n12552 , n10764 , n20427 );
    xnor g26175 ( n12930 , n35929 , n24102 );
    or g26176 ( n7779 , n18703 , n2591 );
    not g26177 ( n16129 , n6185 );
    not g26178 ( n19215 , n7588 );
    and g26179 ( n8071 , n27765 , n12404 );
    not g26180 ( n4368 , n13204 );
    nor g26181 ( n22868 , n24432 , n7544 );
    not g26182 ( n35965 , n11024 );
    or g26183 ( n29992 , n17295 , n27108 );
    nor g26184 ( n14915 , n4962 , n32636 );
    and g26185 ( n22089 , n33110 , n6224 );
    and g26186 ( n24172 , n21628 , n2418 );
    or g26187 ( n8785 , n35773 , n4364 );
    or g26188 ( n27320 , n31538 , n31773 );
    or g26189 ( n19266 , n5423 , n3352 );
    or g26190 ( n12297 , n21120 , n3296 );
    not g26191 ( n17170 , n1950 );
    and g26192 ( n3687 , n21614 , n29055 );
    nor g26193 ( n21154 , n26548 , n26022 );
    or g26194 ( n3328 , n19925 , n2712 );
    and g26195 ( n29133 , n18696 , n13813 );
    xnor g26196 ( n10932 , n35951 , n31799 );
    and g26197 ( n3096 , n32140 , n13765 );
    nor g26198 ( n9849 , n16620 , n25215 );
    nor g26199 ( n3095 , n23004 , n7648 );
    nor g26200 ( n13325 , n23604 , n29367 );
    xnor g26201 ( n28302 , n13109 , n17402 );
    or g26202 ( n10566 , n17981 , n12596 );
    not g26203 ( n2745 , n20840 );
    not g26204 ( n20008 , n26801 );
    or g26205 ( n10919 , n16169 , n29592 );
    and g26206 ( n2215 , n28906 , n26448 );
    or g26207 ( n19778 , n25138 , n14310 );
    and g26208 ( n15659 , n23832 , n19146 );
    or g26209 ( n24137 , n31204 , n26341 );
    or g26210 ( n5398 , n34994 , n27437 );
    nor g26211 ( n27908 , n35574 , n31161 );
    xnor g26212 ( n11692 , n22474 , n8416 );
    or g26213 ( n27073 , n15886 , n28465 );
    or g26214 ( n19247 , n26500 , n31514 );
    or g26215 ( n17116 , n19023 , n22351 );
    or g26216 ( n12245 , n22758 , n9303 );
    xnor g26217 ( n12979 , n23361 , n29535 );
    or g26218 ( n32397 , n13064 , n17872 );
    and g26219 ( n12412 , n1602 , n15905 );
    xnor g26220 ( n18107 , n28383 , n2111 );
    xnor g26221 ( n30085 , n8719 , n20469 );
    or g26222 ( n12723 , n23604 , n28647 );
    xnor g26223 ( n35459 , n31586 , n3205 );
    or g26224 ( n26054 , n20251 , n2689 );
    xnor g26225 ( n1546 , n20404 , n17270 );
    xnor g26226 ( n14374 , n550 , n29839 );
    and g26227 ( n25633 , n23874 , n17047 );
    not g26228 ( n28843 , n26365 );
    or g26229 ( n11955 , n21813 , n31838 );
    and g26230 ( n19456 , n31488 , n20230 );
    nor g26231 ( n513 , n24670 , n12328 );
    and g26232 ( n29214 , n12305 , n17590 );
    and g26233 ( n22010 , n32406 , n11553 );
    and g26234 ( n16573 , n23935 , n14834 );
    not g26235 ( n2190 , n4758 );
    or g26236 ( n19355 , n3917 , n26659 );
    xnor g26237 ( n27438 , n26522 , n16252 );
    and g26238 ( n435 , n13353 , n18135 );
    nor g26239 ( n7002 , n28482 , n4214 );
    or g26240 ( n25285 , n16737 , n2531 );
    nor g26241 ( n4043 , n33434 , n16037 );
    or g26242 ( n9633 , n6463 , n21002 );
    or g26243 ( n35076 , n1302 , n14322 );
    nor g26244 ( n19540 , n13416 , n24751 );
    and g26245 ( n6512 , n21246 , n32802 );
    or g26246 ( n5725 , n15619 , n4784 );
    xnor g26247 ( n25 , n32253 , n32584 );
    and g26248 ( n19106 , n25709 , n4158 );
    xnor g26249 ( n32604 , n19456 , n31215 );
    xnor g26250 ( n14293 , n16537 , n32354 );
    or g26251 ( n9236 , n9503 , n2179 );
    or g26252 ( n20534 , n9658 , n14840 );
    not g26253 ( n10083 , n32572 );
    xnor g26254 ( n36036 , n34326 , n7672 );
    xnor g26255 ( n32314 , n19392 , n31987 );
    and g26256 ( n31116 , n10987 , n8763 );
    and g26257 ( n24587 , n507 , n25573 );
    not g26258 ( n1351 , n9789 );
    or g26259 ( n20742 , n27459 , n16919 );
    xnor g26260 ( n9516 , n32580 , n11455 );
    and g26261 ( n5279 , n18281 , n21572 );
    or g26262 ( n28531 , n22713 , n20812 );
    nor g26263 ( n21953 , n19405 , n13926 );
    xnor g26264 ( n30188 , n30902 , n31727 );
    buf g26265 ( n31606 , n9731 );
    not g26266 ( n5289 , n32857 );
    xnor g26267 ( n22038 , n29397 , n6651 );
    or g26268 ( n24563 , n30217 , n5501 );
    xnor g26269 ( n13866 , n31317 , n33647 );
    nor g26270 ( n30182 , n4962 , n33864 );
    and g26271 ( n21379 , n5869 , n1303 );
    or g26272 ( n31383 , n11046 , n20987 );
    and g26273 ( n10550 , n1246 , n595 );
    or g26274 ( n8046 , n30105 , n10911 );
    or g26275 ( n32809 , n14241 , n9921 );
    or g26276 ( n13006 , n2964 , n7726 );
    xnor g26277 ( n34741 , n30728 , n2229 );
    xnor g26278 ( n12588 , n20947 , n27064 );
    and g26279 ( n24785 , n23153 , n28792 );
    or g26280 ( n34201 , n27003 , n2185 );
    nor g26281 ( n4834 , n7540 , n2393 );
    or g26282 ( n27700 , n26819 , n8349 );
    nor g26283 ( n19129 , n9789 , n8074 );
    or g26284 ( n9234 , n1950 , n23711 );
    and g26285 ( n30762 , n31011 , n19567 );
    or g26286 ( n1011 , n26481 , n9975 );
    and g26287 ( n18040 , n12193 , n30526 );
    and g26288 ( n32674 , n34279 , n35582 );
    or g26289 ( n24308 , n31289 , n6314 );
    or g26290 ( n12421 , n31412 , n25392 );
    or g26291 ( n14657 , n15886 , n32088 );
    xnor g26292 ( n3225 , n31582 , n17568 );
    nor g26293 ( n18776 , n16620 , n27179 );
    or g26294 ( n32592 , n10396 , n4444 );
    or g26295 ( n3727 , n21252 , n18509 );
    or g26296 ( n7053 , n14665 , n33251 );
    and g26297 ( n23760 , n4062 , n1704 );
    or g26298 ( n30119 , n28261 , n35143 );
    or g26299 ( n10813 , n29212 , n1416 );
    xnor g26300 ( n16001 , n26046 , n5335 );
    and g26301 ( n4492 , n35166 , n22443 );
    nor g26302 ( n27030 , n6615 , n30223 );
    and g26303 ( n33173 , n23002 , n3695 );
    and g26304 ( n25267 , n24639 , n638 );
    and g26305 ( n15540 , n12260 , n20992 );
    xnor g26306 ( n20434 , n27457 , n5245 );
    or g26307 ( n29402 , n25455 , n1763 );
    not g26308 ( n17330 , n33042 );
    and g26309 ( n3813 , n34993 , n4425 );
    or g26310 ( n8130 , n35 , n16797 );
    or g26311 ( n6453 , n11455 , n4711 );
    xnor g26312 ( n33408 , n18427 , n27878 );
    or g26313 ( n2594 , n18001 , n14319 );
    or g26314 ( n16523 , n34085 , n6966 );
    or g26315 ( n2691 , n28212 , n10412 );
    or g26316 ( n22607 , n35837 , n3636 );
    nor g26317 ( n17594 , n14976 , n33795 );
    and g26318 ( n9588 , n3632 , n16604 );
    or g26319 ( n7451 , n23744 , n3738 );
    not g26320 ( n21817 , n29731 );
    or g26321 ( n4451 , n7229 , n21780 );
    not g26322 ( n28649 , n17454 );
    xnor g26323 ( n30008 , n4497 , n33331 );
    and g26324 ( n4475 , n12081 , n31543 );
    and g26325 ( n27397 , n14598 , n34525 );
    or g26326 ( n452 , n17345 , n7293 );
    and g26327 ( n18278 , n25442 , n2484 );
    or g26328 ( n19196 , n1950 , n33167 );
    or g26329 ( n26111 , n15305 , n29366 );
    nor g26330 ( n17510 , n32584 , n23854 );
    or g26331 ( n27167 , n20312 , n24652 );
    or g26332 ( n17710 , n30660 , n8392 );
    or g26333 ( n4493 , n34502 , n8594 );
    or g26334 ( n9134 , n32775 , n32959 );
    or g26335 ( n29788 , n26591 , n7537 );
    xnor g26336 ( n19824 , n24950 , n1950 );
    and g26337 ( n12363 , n24828 , n2983 );
    or g26338 ( n34345 , n34680 , n7494 );
    or g26339 ( n30265 , n15886 , n3218 );
    or g26340 ( n23573 , n34879 , n31024 );
    and g26341 ( n20528 , n12564 , n17193 );
    nor g26342 ( n24501 , n4288 , n32250 );
    xor g26343 ( n3237 , n25300 , n27395 );
    or g26344 ( n16887 , n22166 , n35866 );
    xnor g26345 ( n34959 , n13 , n25107 );
    not g26346 ( n32821 , n25761 );
    and g26347 ( n14874 , n12501 , n8052 );
    or g26348 ( n2559 , n973 , n16724 );
    or g26349 ( n17380 , n35927 , n34331 );
    and g26350 ( n9861 , n19705 , n7820 );
    or g26351 ( n6583 , n267 , n16919 );
    or g26352 ( n25060 , n6681 , n9121 );
    or g26353 ( n13914 , n25519 , n17878 );
    or g26354 ( n7632 , n22826 , n5909 );
    or g26355 ( n14714 , n11151 , n6968 );
    or g26356 ( n32244 , n26162 , n7726 );
    not g26357 ( n26647 , n9658 );
    or g26358 ( n898 , n2396 , n1049 );
    xnor g26359 ( n11437 , n9251 , n8375 );
    xnor g26360 ( n15273 , n32110 , n15886 );
    and g26361 ( n35855 , n12051 , n29404 );
    and g26362 ( n16381 , n2623 , n17686 );
    or g26363 ( n31248 , n2815 , n6447 );
    nor g26364 ( n11715 , n37 , n27541 );
    xnor g26365 ( n26550 , n18381 , n30742 );
    xnor g26366 ( n28383 , n3058 , n16922 );
    or g26367 ( n24202 , n18546 , n20817 );
    or g26368 ( n15893 , n11925 , n25255 );
    or g26369 ( n25986 , n21271 , n10417 );
    or g26370 ( n20381 , n17991 , n9915 );
    or g26371 ( n22336 , n17873 , n22855 );
    or g26372 ( n33008 , n23154 , n2798 );
    xnor g26373 ( n29382 , n10393 , n6749 );
    and g26374 ( n35093 , n1138 , n2852 );
    or g26375 ( n29612 , n22632 , n20579 );
    and g26376 ( n10285 , n16071 , n17533 );
    not g26377 ( n21747 , n11960 );
    nor g26378 ( n34899 , n29713 , n7104 );
    or g26379 ( n33521 , n6931 , n2842 );
    or g26380 ( n35810 , n5557 , n4175 );
    xnor g26381 ( n14801 , n17139 , n31289 );
    and g26382 ( n18411 , n28075 , n31335 );
    nor g26383 ( n35973 , n7485 , n8907 );
    or g26384 ( n20088 , n10894 , n33148 );
    and g26385 ( n24589 , n35086 , n22985 );
    not g26386 ( n17412 , n30761 );
    and g26387 ( n1645 , n9671 , n3457 );
    or g26388 ( n13212 , n28997 , n34865 );
    or g26389 ( n17921 , n8614 , n25831 );
    not g26390 ( n29585 , n26365 );
    and g26391 ( n17532 , n16300 , n23973 );
    not g26392 ( n21922 , n25174 );
    xnor g26393 ( n13661 , n32965 , n20257 );
    xnor g26394 ( n25005 , n13713 , n29425 );
    or g26395 ( n29230 , n7662 , n4606 );
    xnor g26396 ( n32744 , n30498 , n26453 );
    and g26397 ( n27111 , n34194 , n4878 );
    and g26398 ( n20687 , n35588 , n26804 );
    or g26399 ( n23965 , n12218 , n14918 );
    xnor g26400 ( n28802 , n21271 , n24332 );
    or g26401 ( n13220 , n14113 , n1384 );
    not g26402 ( n23456 , n24371 );
    xnor g26403 ( n8351 , n28266 , n14612 );
    nor g26404 ( n23019 , n22291 , n866 );
    and g26405 ( n29802 , n33496 , n26062 );
    xnor g26406 ( n20724 , n4785 , n34781 );
    and g26407 ( n6381 , n8570 , n1722 );
    not g26408 ( n22455 , n22291 );
    or g26409 ( n33160 , n3897 , n3736 );
    and g26410 ( n25124 , n8521 , n11283 );
    or g26411 ( n15935 , n8553 , n28668 );
    nor g26412 ( n6738 , n3242 , n12622 );
    xnor g26413 ( n12249 , n6610 , n17508 );
    and g26414 ( n25459 , n31974 , n28152 );
    or g26415 ( n4117 , n22233 , n20840 );
    or g26416 ( n2199 , n19019 , n20308 );
    not g26417 ( n32328 , n19144 );
    xnor g26418 ( n20698 , n5791 , n23456 );
    xnor g26419 ( n32164 , n3788 , n27944 );
    and g26420 ( n34529 , n5059 , n28476 );
    or g26421 ( n24167 , n22045 , n31067 );
    or g26422 ( n35503 , n10939 , n22682 );
    and g26423 ( n3807 , n33305 , n24503 );
    and g26424 ( n4127 , n18969 , n32525 );
    or g26425 ( n23629 , n29295 , n23462 );
    or g26426 ( n7338 , n35712 , n30204 );
    or g26427 ( n11900 , n4476 , n1763 );
    not g26428 ( n13459 , n12477 );
    not g26429 ( n11791 , n5067 );
    or g26430 ( n23533 , n35208 , n27679 );
    or g26431 ( n17369 , n31395 , n13012 );
    or g26432 ( n30250 , n6128 , n1196 );
    nor g26433 ( n10315 , n3397 , n15278 );
    and g26434 ( n4619 , n21760 , n29431 );
    and g26435 ( n13525 , n16466 , n26102 );
    or g26436 ( n35444 , n22223 , n23820 );
    or g26437 ( n10242 , n5770 , n3437 );
    xnor g26438 ( n26956 , n22939 , n32857 );
    or g26439 ( n26200 , n176 , n9601 );
    and g26440 ( n27527 , n26050 , n16928 );
    xnor g26441 ( n11276 , n24279 , n1430 );
    or g26442 ( n6815 , n34780 , n24696 );
    xnor g26443 ( n11047 , n18234 , n3556 );
    or g26444 ( n16680 , n24842 , n15144 );
    xnor g26445 ( n21391 , n3629 , n4960 );
    xnor g26446 ( n14067 , n28181 , n32857 );
    nor g26447 ( n17311 , n34326 , n29203 );
    xnor g26448 ( n25111 , n31258 , n20948 );
    xnor g26449 ( n6331 , n7876 , n4878 );
    xnor g26450 ( n25326 , n26760 , n29839 );
    xnor g26451 ( n6241 , n18209 , n21097 );
    or g26452 ( n3487 , n5738 , n19998 );
    or g26453 ( n26598 , n9658 , n22381 );
    nor g26454 ( n35715 , n9789 , n228 );
    or g26455 ( n7532 , n10339 , n3437 );
    or g26456 ( n27750 , n31437 , n23626 );
    nor g26457 ( n22426 , n28926 , n18287 );
    xor g26458 ( n29620 , n254 , n8452 );
    buf g26459 ( n25831 , n35225 );
    or g26460 ( n4819 , n34429 , n29953 );
    xnor g26461 ( n23467 , n20474 , n10177 );
    and g26462 ( n33056 , n8264 , n25012 );
    xnor g26463 ( n4982 , n3975 , n3019 );
    or g26464 ( n16703 , n25095 , n3432 );
    and g26465 ( n1920 , n17581 , n4103 );
    and g26466 ( n31586 , n25230 , n8506 );
    or g26467 ( n35621 , n26998 , n21579 );
    or g26468 ( n26344 , n32030 , n24861 );
    or g26469 ( n6097 , n14634 , n746 );
    nor g26470 ( n34771 , n18937 , n12563 );
    or g26471 ( n3576 , n28717 , n22206 );
    not g26472 ( n7869 , n25434 );
    and g26473 ( n25482 , n8040 , n11122 );
    or g26474 ( n33401 , n34780 , n11601 );
    or g26475 ( n5322 , n9481 , n14283 );
    or g26476 ( n20667 , n24664 , n17152 );
    xnor g26477 ( n33436 , n34290 , n435 );
    or g26478 ( n17080 , n18379 , n10860 );
    not g26479 ( n18655 , n22980 );
    or g26480 ( n24155 , n29839 , n3895 );
    and g26481 ( n5782 , n35718 , n3158 );
    xnor g26482 ( n22055 , n13672 , n7540 );
    or g26483 ( n6433 , n10544 , n5252 );
    and g26484 ( n5052 , n33726 , n33410 );
    or g26485 ( n8326 , n11046 , n14742 );
    not g26486 ( n8756 , n698 );
    xnor g26487 ( n6451 , n7294 , n15770 );
    or g26488 ( n25490 , n12581 , n1715 );
    or g26489 ( n16907 , n4960 , n32361 );
    and g26490 ( n6468 , n9562 , n14599 );
    xnor g26491 ( n608 , n8479 , n17360 );
    nor g26492 ( n10920 , n11046 , n5152 );
    xnor g26493 ( n25337 , n20332 , n26794 );
    or g26494 ( n2793 , n31799 , n15733 );
    and g26495 ( n26988 , n16639 , n23858 );
    or g26496 ( n29013 , n31559 , n657 );
    and g26497 ( n5623 , n2707 , n21678 );
    or g26498 ( n17463 , n24462 , n32507 );
    nor g26499 ( n6931 , n31799 , n5490 );
    or g26500 ( n20163 , n15415 , n17046 );
    xnor g26501 ( n1613 , n36074 , n23788 );
    xnor g26502 ( n5155 , n8551 , n21084 );
    or g26503 ( n30970 , n32350 , n23187 );
    or g26504 ( n7816 , n4878 , n4880 );
    xnor g26505 ( n22560 , n16167 , n14988 );
    or g26506 ( n24214 , n19551 , n8613 );
    nor g26507 ( n13467 , n9789 , n12078 );
    or g26508 ( n2149 , n1487 , n10381 );
    and g26509 ( n6607 , n17168 , n8183 );
    or g26510 ( n22873 , n6994 , n30808 );
    buf g26511 ( n11258 , n7446 );
    nor g26512 ( n11824 , n15886 , n28367 );
    or g26513 ( n20321 , n23511 , n4217 );
    xnor g26514 ( n27416 , n36065 , n26120 );
    and g26515 ( n11537 , n9630 , n12050 );
    xnor g26516 ( n8456 , n16696 , n10894 );
    nor g26517 ( n22613 , n35431 , n28900 );
    nor g26518 ( n31685 , n32857 , n29318 );
    or g26519 ( n8023 , n7540 , n22123 );
    or g26520 ( n24252 , n15584 , n18398 );
    nor g26521 ( n15614 , n8365 , n7919 );
    not g26522 ( n4440 , n7872 );
    and g26523 ( n17183 , n10200 , n20649 );
    xnor g26524 ( n7634 , n27151 , n32095 );
    and g26525 ( n2721 , n28488 , n6722 );
    or g26526 ( n3427 , n1950 , n24897 );
    or g26527 ( n15082 , n9349 , n443 );
    and g26528 ( n25728 , n5310 , n9584 );
    or g26529 ( n1761 , n2172 , n30141 );
    or g26530 ( n5032 , n10567 , n9951 );
    xnor g26531 ( n12202 , n22110 , n15369 );
    xnor g26532 ( n32684 , n23339 , n32090 );
    and g26533 ( n27021 , n33883 , n27873 );
    or g26534 ( n33147 , n15155 , n6381 );
    or g26535 ( n23123 , n10894 , n15603 );
    and g26536 ( n7654 , n26780 , n23947 );
    and g26537 ( n33728 , n31145 , n35567 );
    not g26538 ( n2658 , n4241 );
    or g26539 ( n19597 , n24999 , n33750 );
    and g26540 ( n31401 , n2958 , n31701 );
    xnor g26541 ( n12117 , n8456 , n12067 );
    xnor g26542 ( n26991 , n19259 , n26726 );
    and g26543 ( n148 , n26147 , n18515 );
    nor g26544 ( n19756 , n24583 , n25922 );
    and g26545 ( n26710 , n23623 , n5596 );
    and g26546 ( n2610 , n7635 , n3032 );
    and g26547 ( n32750 , n5126 , n19234 );
    xnor g26548 ( n18901 , n3147 , n21284 );
    and g26549 ( n12159 , n8795 , n10654 );
    and g26550 ( n166 , n21468 , n12161 );
    or g26551 ( n7717 , n23569 , n9951 );
    and g26552 ( n10314 , n22248 , n25781 );
    xnor g26553 ( n11530 , n21588 , n15464 );
    or g26554 ( n18565 , n18119 , n28857 );
    not g26555 ( n33069 , n18164 );
    and g26556 ( n20537 , n7306 , n30911 );
    or g26557 ( n11628 , n19796 , n24635 );
    or g26558 ( n12065 , n20867 , n31067 );
    and g26559 ( n9958 , n2309 , n8314 );
    and g26560 ( n25523 , n3880 , n35648 );
    or g26561 ( n28380 , n9892 , n35043 );
    and g26562 ( n6749 , n16637 , n27458 );
    and g26563 ( n33491 , n7665 , n5932 );
    or g26564 ( n33449 , n29713 , n26508 );
    and g26565 ( n26916 , n28891 , n11286 );
    nor g26566 ( n30890 , n19634 , n111 );
    and g26567 ( n10630 , n5369 , n2162 );
    and g26568 ( n6973 , n6165 , n26807 );
    xnor g26569 ( n11656 , n11887 , n31429 );
    or g26570 ( n5367 , n7999 , n15969 );
    not g26571 ( n23534 , n7981 );
    xnor g26572 ( n28844 , n2794 , n9793 );
    xnor g26573 ( n5939 , n21893 , n20877 );
    or g26574 ( n14163 , n17965 , n8924 );
    xnor g26575 ( n6508 , n13048 , n35822 );
    not g26576 ( n18397 , n9658 );
    and g26577 ( n24554 , n27264 , n35876 );
    or g26578 ( n35158 , n6425 , n20840 );
    or g26579 ( n10086 , n15342 , n31514 );
    and g26580 ( n34391 , n15109 , n36045 );
    xnor g26581 ( n8654 , n5417 , n9789 );
    not g26582 ( n3850 , n31571 );
    not g26583 ( n20129 , n27291 );
    or g26584 ( n11289 , n29008 , n26892 );
    or g26585 ( n5399 , n34693 , n6307 );
    xnor g26586 ( n3749 , n25995 , n423 );
    and g26587 ( n6807 , n11385 , n34261 );
    or g26588 ( n13999 , n5056 , n22682 );
    nor g26589 ( n15475 , n3041 , n26634 );
    xnor g26590 ( n24596 , n12315 , n15886 );
    nor g26591 ( n33463 , n16922 , n21330 );
    and g26592 ( n14003 , n16846 , n14790 );
    or g26593 ( n506 , n112 , n10526 );
    or g26594 ( n34099 , n4878 , n9684 );
    or g26595 ( n3722 , n22242 , n30732 );
    xnor g26596 ( n10747 , n13389 , n9696 );
    or g26597 ( n7626 , n10042 , n23379 );
    xnor g26598 ( n29765 , n17121 , n26627 );
    and g26599 ( n28900 , n33678 , n31527 );
    or g26600 ( n14095 , n4878 , n16222 );
    nor g26601 ( n21565 , n1950 , n8080 );
    or g26602 ( n17683 , n33341 , n16396 );
    and g26603 ( n35253 , n23039 , n2441 );
    not g26604 ( n17765 , n24739 );
    xnor g26605 ( n11904 , n27250 , n14835 );
    xnor g26606 ( n27751 , n32748 , n26106 );
    or g26607 ( n2449 , n15299 , n32335 );
    and g26608 ( n16250 , n25791 , n19326 );
    or g26609 ( n24014 , n8716 , n14689 );
    xnor g26610 ( n23062 , n23233 , n35895 );
    or g26611 ( n13463 , n20723 , n27114 );
    and g26612 ( n8398 , n27071 , n30281 );
    and g26613 ( n16058 , n6395 , n12611 );
    or g26614 ( n21526 , n15032 , n2823 );
    or g26615 ( n3042 , n2076 , n11104 );
    or g26616 ( n7180 , n78 , n3694 );
    or g26617 ( n35020 , n31793 , n11312 );
    or g26618 ( n10322 , n8993 , n9916 );
    xnor g26619 ( n819 , n13633 , n25499 );
    not g26620 ( n4108 , n20558 );
    not g26621 ( n9123 , n34072 );
    or g26622 ( n7332 , n18066 , n24710 );
    not g26623 ( n22482 , n19641 );
    or g26624 ( n26193 , n13475 , n1133 );
    or g26625 ( n33100 , n4962 , n21014 );
    xnor g26626 ( n26551 , n28312 , n25710 );
    nor g26627 ( n31399 , n15886 , n9401 );
    or g26628 ( n13317 , n13821 , n26958 );
    and g26629 ( n14269 , n24808 , n21925 );
    and g26630 ( n31245 , n9111 , n10454 );
    nor g26631 ( n17174 , n25602 , n9205 );
    nor g26632 ( n29493 , n15301 , n25610 );
    or g26633 ( n6066 , n23725 , n8618 );
    not g26634 ( n4104 , n1396 );
    and g26635 ( n14659 , n20133 , n32156 );
    xnor g26636 ( n28480 , n5657 , n2651 );
    or g26637 ( n34417 , n21000 , n22977 );
    not g26638 ( n2389 , n12374 );
    or g26639 ( n28466 , n22859 , n17125 );
    and g26640 ( n9418 , n21423 , n5385 );
    and g26641 ( n23918 , n23497 , n18727 );
    or g26642 ( n5255 , n24371 , n19284 );
    or g26643 ( n34573 , n23375 , n25019 );
    or g26644 ( n13917 , n26588 , n11850 );
    and g26645 ( n15697 , n24605 , n21036 );
    or g26646 ( n2257 , n26628 , n9672 );
    xnor g26647 ( n35743 , n18300 , n7348 );
    xnor g26648 ( n24619 , n6080 , n29063 );
    xnor g26649 ( n17513 , n11551 , n3553 );
    or g26650 ( n16720 , n3992 , n2117 );
    nor g26651 ( n10793 , n16025 , n33605 );
    or g26652 ( n22297 , n30042 , n20605 );
    buf g26653 ( n18121 , n905 );
    and g26654 ( n24756 , n5540 , n31865 );
    or g26655 ( n30915 , n16116 , n21627 );
    xnor g26656 ( n19275 , n17094 , n19377 );
    xnor g26657 ( n17262 , n23846 , n29237 );
    not g26658 ( n23986 , n35507 );
    or g26659 ( n1489 , n19000 , n21691 );
    or g26660 ( n34654 , n9789 , n32101 );
    and g26661 ( n19478 , n17821 , n28588 );
    and g26662 ( n34889 , n8442 , n4583 );
    or g26663 ( n18747 , n25174 , n20406 );
    nor g26664 ( n18110 , n4288 , n23920 );
    or g26665 ( n226 , n2140 , n32808 );
    and g26666 ( n1484 , n30803 , n17614 );
    or g26667 ( n20704 , n35340 , n6879 );
    and g26668 ( n14441 , n30038 , n6234 );
    or g26669 ( n18312 , n18310 , n14167 );
    and g26670 ( n16953 , n1223 , n26421 );
    or g26671 ( n6547 , n19934 , n34537 );
    xnor g26672 ( n31505 , n5085 , n15700 );
    or g26673 ( n494 , n29513 , n13495 );
    or g26674 ( n28497 , n7124 , n19131 );
    and g26675 ( n5634 , n31653 , n12312 );
    xnor g26676 ( n1052 , n32431 , n35314 );
    or g26677 ( n34996 , n4380 , n14841 );
    xnor g26678 ( n10833 , n13457 , n29839 );
    not g26679 ( n8273 , n16620 );
    not g26680 ( n30884 , n22980 );
    or g26681 ( n25235 , n33373 , n10417 );
    xnor g26682 ( n35325 , n23579 , n32095 );
    or g26683 ( n23885 , n32549 , n23209 );
    not g26684 ( n26418 , n4852 );
    and g26685 ( n17699 , n19344 , n17032 );
    or g26686 ( n18428 , n29362 , n29330 );
    and g26687 ( n19553 , n21605 , n7203 );
    and g26688 ( n2044 , n31663 , n16076 );
    nor g26689 ( n28013 , n27823 , n27351 );
    or g26690 ( n33570 , n19844 , n5709 );
    or g26691 ( n8128 , n6454 , n1293 );
    xnor g26692 ( n20550 , n6761 , n24741 );
    buf g26693 ( n32505 , n15871 );
    or g26694 ( n26425 , n19605 , n2523 );
    and g26695 ( n18224 , n30982 , n22980 );
    xnor g26696 ( n2197 , n3985 , n23281 );
    or g26697 ( n25960 , n15729 , n2706 );
    or g26698 ( n9728 , n33528 , n1920 );
    or g26699 ( n28158 , n15673 , n16797 );
    or g26700 ( n26999 , n13461 , n27973 );
    and g26701 ( n33983 , n21334 , n35024 );
    or g26702 ( n14152 , n19917 , n26883 );
    and g26703 ( n15518 , n32552 , n25621 );
    and g26704 ( n21311 , n21399 , n7743 );
    xnor g26705 ( n34631 , n34374 , n18272 );
    and g26706 ( n14620 , n33869 , n25809 );
    xnor g26707 ( n35590 , n11807 , n8319 );
    or g26708 ( n2650 , n34430 , n14787 );
    or g26709 ( n18773 , n30742 , n18927 );
    buf g26710 ( n15439 , n28893 );
    not g26711 ( n34487 , n26977 );
    not g26712 ( n16186 , n11174 );
    or g26713 ( n30815 , n17542 , n33448 );
    not g26714 ( n17958 , n11190 );
    xnor g26715 ( n25549 , n1254 , n33786 );
    and g26716 ( n26048 , n5292 , n10483 );
    nor g26717 ( n32746 , n1160 , n18739 );
    or g26718 ( n11045 , n5174 , n20478 );
    or g26719 ( n22603 , n29929 , n4490 );
    or g26720 ( n11631 , n25163 , n11850 );
    or g26721 ( n8166 , n20238 , n21684 );
    and g26722 ( n7301 , n5812 , n13218 );
    or g26723 ( n35406 , n29398 , n34862 );
    xnor g26724 ( n12090 , n31371 , n13824 );
    and g26725 ( n30467 , n3053 , n27494 );
    or g26726 ( n34384 , n20400 , n20576 );
    or g26727 ( n29063 , n26294 , n20301 );
    nor g26728 ( n14818 , n28374 , n19430 );
    not g26729 ( n7320 , n30501 );
    xnor g26730 ( n25636 , n3146 , n8184 );
    not g26731 ( n17887 , n25174 );
    and g26732 ( n11182 , n18989 , n16620 );
    or g26733 ( n3108 , n29713 , n26906 );
    nor g26734 ( n35334 , n7891 , n22200 );
    xnor g26735 ( n11004 , n25982 , n30742 );
    or g26736 ( n21846 , n29491 , n35109 );
    and g26737 ( n23270 , n13645 , n26904 );
    not g26738 ( n30917 , n31289 );
    or g26739 ( n30259 , n25174 , n20336 );
    xnor g26740 ( n13282 , n5706 , n11570 );
    xnor g26741 ( n33492 , n24107 , n7709 );
    and g26742 ( n31936 , n33267 , n30265 );
    or g26743 ( n32765 , n32095 , n7399 );
    nor g26744 ( n31724 , n29839 , n29160 );
    or g26745 ( n2268 , n22173 , n34814 );
    xnor g26746 ( n27258 , n17498 , n11190 );
    and g26747 ( n23614 , n24259 , n9558 );
    or g26748 ( n27329 , n1632 , n24582 );
    not g26749 ( n17089 , n6566 );
    nor g26750 ( n1697 , n1950 , n8121 );
    not g26751 ( n15855 , n12146 );
    xnor g26752 ( n35517 , n7140 , n29134 );
    xnor g26753 ( n24852 , n632 , n9789 );
    nor g26754 ( n18055 , n15917 , n28065 );
    not g26755 ( n24026 , n7940 );
    or g26756 ( n25632 , n11406 , n2479 );
    xnor g26757 ( n36074 , n9760 , n18603 );
    or g26758 ( n4605 , n29957 , n15109 );
    or g26759 ( n10899 , n4288 , n9010 );
    and g26760 ( n22402 , n570 , n34137 );
    or g26761 ( n1820 , n821 , n19241 );
    xnor g26762 ( n33985 , n27773 , n927 );
    or g26763 ( n17639 , n20766 , n31627 );
    xnor g26764 ( n12721 , n21897 , n23806 );
    xnor g26765 ( n22208 , n12756 , n12910 );
    or g26766 ( n33184 , n3875 , n4727 );
    xnor g26767 ( n13508 , n5115 , n32095 );
    xnor g26768 ( n33084 , n14468 , n24957 );
    xnor g26769 ( n30878 , n23467 , n12609 );
    or g26770 ( n6555 , n8985 , n34484 );
    or g26771 ( n20992 , n28055 , n33358 );
    nor g26772 ( n1686 , n4962 , n6761 );
    or g26773 ( n17182 , n5221 , n19351 );
    or g26774 ( n17929 , n27250 , n17233 );
    or g26775 ( n7375 , n33888 , n1763 );
    not g26776 ( n27294 , n32857 );
    or g26777 ( n8048 , n16920 , n32505 );
    or g26778 ( n9660 , n25382 , n30667 );
    xnor g26779 ( n22229 , n17699 , n5335 );
    and g26780 ( n8963 , n7686 , n30022 );
    or g26781 ( n2569 , n35346 , n17872 );
    or g26782 ( n19569 , n320 , n13900 );
    or g26783 ( n32105 , n23691 , n10953 );
    and g26784 ( n30382 , n31252 , n8698 );
    or g26785 ( n30602 , n34232 , n31912 );
    and g26786 ( n8600 , n17213 , n1929 );
    and g26787 ( n23869 , n1368 , n31917 );
    or g26788 ( n14372 , n6200 , n7792 );
    xnor g26789 ( n25933 , n8358 , n3205 );
    xnor g26790 ( n11281 , n6644 , n5171 );
    or g26791 ( n35435 , n7442 , n17974 );
    and g26792 ( n9764 , n20278 , n6184 );
    or g26793 ( n193 , n6753 , n2712 );
    or g26794 ( n26714 , n34821 , n14651 );
    buf g26795 ( n27437 , n27890 );
    xnor g26796 ( n27577 , n25346 , n2472 );
    and g26797 ( n12131 , n2445 , n5813 );
    or g26798 ( n6202 , n18667 , n33785 );
    or g26799 ( n13698 , n19819 , n35935 );
    xnor g26800 ( n16973 , n4977 , n10840 );
    xnor g26801 ( n10698 , n8933 , n34063 );
    or g26802 ( n14857 , n12131 , n17829 );
    or g26803 ( n32708 , n32715 , n11914 );
    xnor g26804 ( n15883 , n3888 , n9135 );
    and g26805 ( n25026 , n20895 , n35689 );
    or g26806 ( n33690 , n32857 , n421 );
    xnor g26807 ( n16002 , n30948 , n10267 );
    not g26808 ( n30616 , n11269 );
    xnor g26809 ( n33825 , n12461 , n4334 );
    or g26810 ( n26094 , n34741 , n3842 );
    or g26811 ( n28488 , n20202 , n19105 );
    or g26812 ( n5333 , n7667 , n32379 );
    xnor g26813 ( n35079 , n8382 , n15547 );
    or g26814 ( n3084 , n3822 , n24259 );
    xnor g26815 ( n13429 , n19002 , n8043 );
    nor g26816 ( n25527 , n31289 , n27211 );
    or g26817 ( n21913 , n6028 , n2885 );
    or g26818 ( n2671 , n4962 , n3005 );
    or g26819 ( n26462 , n15539 , n26212 );
    or g26820 ( n2855 , n9834 , n5124 );
    or g26821 ( n32249 , n2271 , n14706 );
    or g26822 ( n6842 , n27484 , n24772 );
    xnor g26823 ( n8621 , n32058 , n18379 );
    and g26824 ( n29539 , n6583 , n35091 );
    nor g26825 ( n17352 , n7026 , n16389 );
    or g26826 ( n13289 , n17104 , n8109 );
    or g26827 ( n34895 , n30742 , n30798 );
    or g26828 ( n12610 , n35927 , n19790 );
    not g26829 ( n8092 , n30742 );
    or g26830 ( n32061 , n27400 , n23284 );
    or g26831 ( n28353 , n30084 , n5868 );
    and g26832 ( n1801 , n8568 , n8633 );
    xnor g26833 ( n24763 , n7142 , n33557 );
    not g26834 ( n9558 , n31692 );
    and g26835 ( n6972 , n18604 , n6798 );
    xnor g26836 ( n3927 , n27950 , n32857 );
    or g26837 ( n32195 , n15813 , n26737 );
    or g26838 ( n24391 , n16220 , n25761 );
    or g26839 ( n9013 , n35667 , n10336 );
    or g26840 ( n31405 , n9384 , n28324 );
    not g26841 ( n35410 , n23909 );
    or g26842 ( n29819 , n4192 , n16326 );
    or g26843 ( n13272 , n3327 , n34814 );
    xnor g26844 ( n34473 , n31362 , n18379 );
    or g26845 ( n25221 , n14383 , n14390 );
    nor g26846 ( n407 , n760 , n31557 );
    buf g26847 ( n5252 , n27404 );
    or g26848 ( n12770 , n8250 , n12596 );
    nor g26849 ( n7796 , n32715 , n22394 );
    and g26850 ( n34030 , n22352 , n33289 );
    or g26851 ( n7506 , n28551 , n28788 );
    or g26852 ( n20286 , n9744 , n20851 );
    xnor g26853 ( n10173 , n20821 , n7122 );
    not g26854 ( n23407 , n2409 );
    or g26855 ( n15458 , n1393 , n11312 );
    xnor g26856 ( n6287 , n3009 , n6909 );
    or g26857 ( n23607 , n14879 , n22480 );
    or g26858 ( n13882 , n27985 , n1511 );
    xnor g26859 ( n8257 , n23161 , n30906 );
    xnor g26860 ( n23531 , n13069 , n35864 );
    or g26861 ( n22960 , n15476 , n31514 );
    or g26862 ( n19797 , n11040 , n6008 );
    nor g26863 ( n1373 , n24599 , n8493 );
    and g26864 ( n27880 , n35861 , n12776 );
    and g26865 ( n17339 , n29374 , n26999 );
    xnor g26866 ( n8212 , n30401 , n11046 );
    or g26867 ( n21216 , n34005 , n11996 );
    xnor g26868 ( n33928 , n15150 , n16922 );
    or g26869 ( n34901 , n15085 , n30708 );
    xnor g26870 ( n25819 , n30594 , n28710 );
    xnor g26871 ( n1410 , n23114 , n1588 );
    or g26872 ( n29749 , n682 , n21862 );
    nor g26873 ( n7349 , n13848 , n12553 );
    or g26874 ( n34396 , n55 , n33498 );
    or g26875 ( n22917 , n10527 , n14866 );
    or g26876 ( n13968 , n32857 , n12262 );
    and g26877 ( n32539 , n16949 , n2425 );
    or g26878 ( n8316 , n35590 , n115 );
    buf g26879 ( n9980 , n33840 );
    nor g26880 ( n2422 , n6325 , n23323 );
    xnor g26881 ( n583 , n31392 , n12922 );
    xnor g26882 ( n7661 , n32290 , n35927 );
    and g26883 ( n26915 , n9971 , n11371 );
    and g26884 ( n33124 , n12378 , n8508 );
    or g26885 ( n29067 , n4288 , n14687 );
    and g26886 ( n24608 , n24045 , n31914 );
    xnor g26887 ( n5241 , n29318 , n7712 );
    or g26888 ( n18608 , n10941 , n27512 );
    and g26889 ( n23707 , n516 , n9176 );
    and g26890 ( n31793 , n20923 , n29576 );
    not g26891 ( n20140 , n3437 );
    or g26892 ( n11063 , n9793 , n3548 );
    or g26893 ( n8598 , n1563 , n33420 );
    not g26894 ( n24400 , n18596 );
    or g26895 ( n2500 , n11259 , n27853 );
    and g26896 ( n6254 , n13208 , n1193 );
    xnor g26897 ( n2161 , n16805 , n27407 );
    xnor g26898 ( n34819 , n3475 , n4822 );
    and g26899 ( n32493 , n11519 , n10304 );
    or g26900 ( n10399 , n22922 , n4561 );
    or g26901 ( n3656 , n4288 , n3364 );
    or g26902 ( n25784 , n28219 , n11703 );
    or g26903 ( n11080 , n18756 , n35258 );
    and g26904 ( n4965 , n7522 , n16596 );
    or g26905 ( n16055 , n26609 , n18533 );
    not g26906 ( n6984 , n35804 );
    not g26907 ( n25889 , n24371 );
    or g26908 ( n16813 , n28943 , n25648 );
    or g26909 ( n20442 , n24435 , n25831 );
    xnor g26910 ( n990 , n32338 , n1950 );
    xnor g26911 ( n851 , n9599 , n27724 );
    not g26912 ( n26726 , n30742 );
    xnor g26913 ( n23583 , n1745 , n32095 );
    xnor g26914 ( n22488 , n23875 , n16609 );
    and g26915 ( n21012 , n21461 , n21527 );
    or g26916 ( n7335 , n19190 , n2682 );
    or g26917 ( n25962 , n8388 , n26023 );
    or g26918 ( n19230 , n27611 , n7417 );
    not g26919 ( n7022 , n21594 );
    or g26920 ( n32966 , n29422 , n28839 );
    xnor g26921 ( n22474 , n34527 , n19551 );
    or g26922 ( n2995 , n6421 , n15552 );
    xnor g26923 ( n21060 , n5985 , n1482 );
    xnor g26924 ( n13794 , n33844 , n32095 );
    or g26925 ( n30685 , n28367 , n3352 );
    and g26926 ( n15168 , n23376 , n2068 );
    not g26927 ( n755 , n27289 );
    xnor g26928 ( n7559 , n33049 , n16922 );
    or g26929 ( n27307 , n9894 , n21714 );
    xnor g26930 ( n3873 , n4830 , n13452 );
    or g26931 ( n35918 , n31608 , n25193 );
    and g26932 ( n31107 , n30847 , n18146 );
    or g26933 ( n32296 , n13229 , n24356 );
    or g26934 ( n6198 , n12683 , n27501 );
    or g26935 ( n32490 , n2626 , n15737 );
    or g26936 ( n3425 , n13715 , n22487 );
    and g26937 ( n22589 , n12109 , n20433 );
    or g26938 ( n26363 , n17568 , n1451 );
    xnor g26939 ( n33438 , n16575 , n25830 );
    or g26940 ( n32962 , n17421 , n19952 );
    or g26941 ( n28893 , n34534 , n3132 );
    or g26942 ( n1025 , n4690 , n9604 );
    or g26943 ( n12530 , n1155 , n11218 );
    and g26944 ( n27833 , n27483 , n33080 );
    not g26945 ( n30333 , n13198 );
    or g26946 ( n2265 , n7573 , n17483 );
    or g26947 ( n14426 , n30562 , n16456 );
    xnor g26948 ( n32686 , n18165 , n29871 );
    xnor g26949 ( n14279 , n9800 , n9165 );
    xnor g26950 ( n1632 , n23761 , n5287 );
    or g26951 ( n29825 , n5662 , n2849 );
    not g26952 ( n23625 , n35938 );
    xnor g26953 ( n3113 , n8982 , n22657 );
    or g26954 ( n15593 , n4766 , n20001 );
    or g26955 ( n18629 , n25174 , n1181 );
    and g26956 ( n28342 , n28841 , n25929 );
    or g26957 ( n13067 , n31799 , n29796 );
    or g26958 ( n1536 , n6698 , n18477 );
    and g26959 ( n5376 , n32162 , n12314 );
    not g26960 ( n15872 , n17568 );
    or g26961 ( n22385 , n5553 , n28890 );
    nor g26962 ( n5078 , n31559 , n18263 );
    xnor g26963 ( n13611 , n154 , n16192 );
    and g26964 ( n20001 , n20788 , n20481 );
    xnor g26965 ( n846 , n2276 , n29839 );
    or g26966 ( n28129 , n29188 , n21862 );
    and g26967 ( n12036 , n30148 , n30261 );
    or g26968 ( n15280 , n6595 , n1048 );
    xnor g26969 ( n29068 , n6332 , n9789 );
    nor g26970 ( n15542 , n18062 , n29349 );
    not g26971 ( n1494 , n7435 );
    not g26972 ( n947 , n7540 );
    or g26973 ( n19055 , n4226 , n22783 );
    nor g26974 ( n13160 , n14037 , n31411 );
    or g26975 ( n10827 , n14358 , n3188 );
    and g26976 ( n15034 , n7920 , n29147 );
    xnor g26977 ( n10387 , n13820 , n11680 );
    not g26978 ( n34505 , n3166 );
    or g26979 ( n3150 , n18695 , n30519 );
    and g26980 ( n34796 , n6303 , n1284 );
    nor g26981 ( n1600 , n2547 , n21644 );
    xnor g26982 ( n27277 , n8103 , n34254 );
    xnor g26983 ( n17373 , n35797 , n32872 );
    or g26984 ( n15331 , n26949 , n29703 );
    or g26985 ( n18168 , n16952 , n9298 );
    or g26986 ( n12861 , n25549 , n21042 );
    or g26987 ( n18172 , n22803 , n3634 );
    nor g26988 ( n14787 , n10452 , n32186 );
    not g26989 ( n34821 , n29037 );
    or g26990 ( n8730 , n10549 , n9861 );
    or g26991 ( n3027 , n32095 , n31762 );
    and g26992 ( n16519 , n21519 , n31980 );
    xnor g26993 ( n9618 , n15957 , n10882 );
    or g26994 ( n4704 , n32569 , n19084 );
    and g26995 ( n5488 , n4931 , n15387 );
    or g26996 ( n1262 , n31272 , n878 );
    nor g26997 ( n5705 , n22822 , n21701 );
    or g26998 ( n31942 , n9095 , n19281 );
    and g26999 ( n31412 , n31490 , n29254 );
    xnor g27000 ( n9994 , n17478 , n6349 );
    xnor g27001 ( n22069 , n33993 , n9658 );
    or g27002 ( n2577 , n30614 , n19939 );
    or g27003 ( n20077 , n16135 , n653 );
    not g27004 ( n6736 , n21017 );
    or g27005 ( n18902 , n30308 , n30419 );
    and g27006 ( n19447 , n17272 , n30412 );
    xnor g27007 ( n14105 , n8870 , n24739 );
    or g27008 ( n8496 , n12580 , n23323 );
    or g27009 ( n2908 , n2013 , n3634 );
    or g27010 ( n20599 , n23961 , n3756 );
    and g27011 ( n24008 , n26120 , n36065 );
    or g27012 ( n16753 , n29713 , n28429 );
    or g27013 ( n5267 , n32234 , n12448 );
    or g27014 ( n20456 , n18981 , n8392 );
    and g27015 ( n8807 , n32149 , n30696 );
    or g27016 ( n17477 , n5562 , n5900 );
    not g27017 ( n792 , n22579 );
    or g27018 ( n24874 , n3877 , n19733 );
    or g27019 ( n6928 , n32154 , n9555 );
    or g27020 ( n14250 , n3311 , n35005 );
    or g27021 ( n6283 , n35813 , n1379 );
    or g27022 ( n22197 , n19984 , n17751 );
    and g27023 ( n5022 , n9459 , n1024 );
    xnor g27024 ( n21814 , n29469 , n850 );
    xnor g27025 ( n7178 , n34915 , n18157 );
    and g27026 ( n4120 , n17908 , n26322 );
    not g27027 ( n4823 , n1721 );
    and g27028 ( n18101 , n14690 , n34237 );
    or g27029 ( n26152 , n29206 , n139 );
    xnor g27030 ( n57 , n20206 , n1950 );
    and g27031 ( n28634 , n17550 , n25029 );
    or g27032 ( n26948 , n1512 , n3805 );
    and g27033 ( n22130 , n32854 , n19254 );
    or g27034 ( n31029 , n10071 , n6950 );
    or g27035 ( n6577 , n17613 , n29033 );
    and g27036 ( n10647 , n18454 , n10985 );
    or g27037 ( n33253 , n17568 , n18201 );
    or g27038 ( n18400 , n12358 , n763 );
    and g27039 ( n9758 , n26516 , n9935 );
    xnor g27040 ( n29518 , n23647 , n12933 );
    nor g27041 ( n28403 , n3205 , n12127 );
    xnor g27042 ( n28345 , n19827 , n32095 );
    nor g27043 ( n26134 , n3715 , n18115 );
    xnor g27044 ( n30588 , n24360 , n32095 );
    xnor g27045 ( n5555 , n3143 , n29839 );
    or g27046 ( n10000 , n32110 , n24489 );
    or g27047 ( n31226 , n31133 , n34537 );
    xnor g27048 ( n30 , n21330 , n11678 );
    not g27049 ( n32732 , n35495 );
    nor g27050 ( n18090 , n33888 , n34406 );
    nor g27051 ( n10585 , n32584 , n30185 );
    xnor g27052 ( n1453 , n7583 , n11046 );
    or g27053 ( n15078 , n14610 , n28719 );
    xnor g27054 ( n34706 , n4551 , n35927 );
    and g27055 ( n19335 , n29750 , n4404 );
    or g27056 ( n35752 , n26765 , n26480 );
    or g27057 ( n32846 , n29821 , n30708 );
    xnor g27058 ( n26604 , n33811 , n9960 );
    not g27059 ( n1518 , n24383 );
    and g27060 ( n7484 , n15418 , n20105 );
    xor g27061 ( n28343 , n35784 , n30285 );
    or g27062 ( n27100 , n30949 , n25855 );
    xnor g27063 ( n18222 , n18871 , n25951 );
    or g27064 ( n15679 , n27658 , n21644 );
    and g27065 ( n28449 , n26395 , n9902 );
    or g27066 ( n1701 , n20571 , n35619 );
    and g27067 ( n27070 , n10735 , n5357 );
    xnor g27068 ( n14373 , n152 , n25602 );
    or g27069 ( n35714 , n2928 , n1386 );
    and g27070 ( n18923 , n18142 , n13602 );
    or g27071 ( n32723 , n4300 , n21210 );
    or g27072 ( n35513 , n19551 , n32641 );
    or g27073 ( n4696 , n5307 , n25583 );
    or g27074 ( n14669 , n30836 , n27973 );
    not g27075 ( n2889 , n19322 );
    and g27076 ( n205 , n34875 , n6219 );
    and g27077 ( n16114 , n26230 , n1157 );
    xnor g27078 ( n17022 , n512 , n5335 );
    or g27079 ( n11314 , n12049 , n32006 );
    or g27080 ( n32947 , n23013 , n18477 );
    xnor g27081 ( n25330 , n28692 , n16904 );
    not g27082 ( n6008 , n14564 );
    and g27083 ( n35995 , n23344 , n35305 );
    and g27084 ( n20460 , n10692 , n32994 );
    or g27085 ( n25186 , n750 , n30680 );
    and g27086 ( n25241 , n30815 , n24821 );
    xnor g27087 ( n20154 , n21610 , n31936 );
    or g27088 ( n29936 , n19551 , n6629 );
    or g27089 ( n24649 , n30128 , n35422 );
    and g27090 ( n26690 , n21665 , n22559 );
    nor g27091 ( n24438 , n1950 , n569 );
    or g27092 ( n6903 , n1129 , n27759 );
    buf g27093 ( n139 , n31549 );
    not g27094 ( n21397 , n17751 );
    not g27095 ( n25390 , n22471 );
    buf g27096 ( n24025 , n4036 );
    and g27097 ( n15774 , n31016 , n8973 );
    or g27098 ( n25675 , n27444 , n19265 );
    nor g27099 ( n22896 , n11046 , n9273 );
    xnor g27100 ( n1153 , n6373 , n3647 );
    and g27101 ( n31792 , n34861 , n16957 );
    and g27102 ( n22144 , n25529 , n3030 );
    xnor g27103 ( n23017 , n4598 , n34408 );
    xnor g27104 ( n25677 , n29467 , n28078 );
    or g27105 ( n18592 , n7014 , n27625 );
    xnor g27106 ( n5658 , n15448 , n9239 );
    xnor g27107 ( n7832 , n19152 , n32676 );
    or g27108 ( n33289 , n28206 , n20762 );
    or g27109 ( n19916 , n3838 , n4772 );
    or g27110 ( n18175 , n12519 , n30732 );
    and g27111 ( n1174 , n31445 , n27545 );
    or g27112 ( n12687 , n32095 , n32275 );
    and g27113 ( n6064 , n2797 , n12056 );
    or g27114 ( n30082 , n9388 , n34806 );
    not g27115 ( n34040 , n11607 );
    or g27116 ( n26 , n35483 , n6285 );
    not g27117 ( n30088 , n27656 );
    xnor g27118 ( n1889 , n15768 , n29249 );
    or g27119 ( n18619 , n16944 , n5395 );
    and g27120 ( n648 , n13737 , n26907 );
    or g27121 ( n15864 , n28888 , n25036 );
    or g27122 ( n1669 , n21978 , n33034 );
    nor g27123 ( n35131 , n4960 , n2138 );
    or g27124 ( n13650 , n28794 , n17855 );
    not g27125 ( n26818 , n19939 );
    xnor g27126 ( n34429 , n28899 , n5209 );
    or g27127 ( n12427 , n20205 , n1642 );
    and g27128 ( n21464 , n3302 , n5828 );
    not g27129 ( n18097 , n25602 );
    xnor g27130 ( n30304 , n23883 , n9793 );
    or g27131 ( n30340 , n5204 , n6509 );
    or g27132 ( n8615 , n3554 , n22356 );
    and g27133 ( n34455 , n3381 , n30363 );
    not g27134 ( n15544 , n12384 );
    not g27135 ( n34609 , n17891 );
    xnor g27136 ( n16265 , n27741 , n31559 );
    not g27137 ( n24454 , n7677 );
    xnor g27138 ( n13476 , n22649 , n32857 );
    or g27139 ( n35527 , n25329 , n20194 );
    xnor g27140 ( n16759 , n36081 , n3205 );
    and g27141 ( n18643 , n10574 , n7545 );
    xnor g27142 ( n18414 , n35062 , n25836 );
    and g27143 ( n33189 , n10170 , n16807 );
    or g27144 ( n32562 , n8192 , n17781 );
    xnor g27145 ( n22311 , n8564 , n3222 );
    or g27146 ( n5053 , n28784 , n23259 );
    or g27147 ( n31894 , n16046 , n34600 );
    or g27148 ( n24163 , n1943 , n8478 );
    or g27149 ( n32134 , n7874 , n15541 );
    and g27150 ( n25903 , n36031 , n24106 );
    or g27151 ( n32474 , n27834 , n30519 );
    or g27152 ( n2692 , n12573 , n12428 );
    or g27153 ( n558 , n24147 , n10475 );
    or g27154 ( n16713 , n10222 , n28248 );
    or g27155 ( n22936 , n26100 , n3437 );
    not g27156 ( n31684 , n24788 );
    not g27157 ( n15706 , n29713 );
    or g27158 ( n9176 , n31056 , n6388 );
    or g27159 ( n17065 , n26229 , n2168 );
    or g27160 ( n14173 , n18118 , n28438 );
    xnor g27161 ( n32023 , n15878 , n4960 );
    and g27162 ( n658 , n26957 , n4864 );
    xnor g27163 ( n15293 , n25997 , n9021 );
    not g27164 ( n27560 , n25073 );
    or g27165 ( n17504 , n19551 , n22280 );
    or g27166 ( n6914 , n27739 , n13215 );
    xnor g27167 ( n12848 , n33864 , n4962 );
    nor g27168 ( n2074 , n17241 , n7448 );
    xnor g27169 ( n14288 , n24222 , n24371 );
    nor g27170 ( n10464 , n32189 , n13735 );
    or g27171 ( n3817 , n19551 , n26313 );
    xnor g27172 ( n23812 , n26021 , n26443 );
    or g27173 ( n25213 , n11455 , n5597 );
    xnor g27174 ( n30094 , n18252 , n31939 );
    xnor g27175 ( n30239 , n6060 , n20118 );
    nor g27176 ( n3135 , n4878 , n6427 );
    xnor g27177 ( n5760 , n30147 , n27990 );
    not g27178 ( n10769 , n31799 );
    or g27179 ( n18577 , n4288 , n20403 );
    or g27180 ( n24825 , n16922 , n26729 );
    or g27181 ( n495 , n2907 , n22834 );
    and g27182 ( n14578 , n4643 , n34772 );
    not g27183 ( n1236 , n5989 );
    or g27184 ( n28053 , n3094 , n4478 );
    or g27185 ( n16333 , n26887 , n1414 );
    nor g27186 ( n10151 , n7159 , n14512 );
    xnor g27187 ( n22137 , n16342 , n6721 );
    or g27188 ( n21939 , n32202 , n2535 );
    and g27189 ( n8722 , n15120 , n17146 );
    or g27190 ( n8390 , n9320 , n28455 );
    xnor g27191 ( n21447 , n8612 , n35388 );
    and g27192 ( n1105 , n27609 , n685 );
    xnor g27193 ( n21815 , n24280 , n5924 );
    not g27194 ( n29174 , n28866 );
    or g27195 ( n4644 , n10799 , n6374 );
    nor g27196 ( n19502 , n25845 , n24841 );
    xnor g27197 ( n2152 , n27442 , n8904 );
    or g27198 ( n29281 , n32633 , n22682 );
    xnor g27199 ( n8118 , n24106 , n36031 );
    nor g27200 ( n32733 , n31799 , n5090 );
    or g27201 ( n29542 , n14575 , n24259 );
    or g27202 ( n24805 , n19551 , n17258 );
    or g27203 ( n67 , n5070 , n1414 );
    or g27204 ( n30321 , n20225 , n12596 );
    xnor g27205 ( n4001 , n27078 , n2748 );
    xnor g27206 ( n13192 , n34111 , n22270 );
    or g27207 ( n19056 , n11425 , n4279 );
    or g27208 ( n31176 , n32715 , n30417 );
    or g27209 ( n1144 , n20821 , n23187 );
    xnor g27210 ( n14999 , n4893 , n31559 );
    xnor g27211 ( n8899 , n362 , n15363 );
    nor g27212 ( n12370 , n19841 , n19061 );
    or g27213 ( n787 , n19311 , n12585 );
    and g27214 ( n6384 , n5636 , n17426 );
    and g27215 ( n35920 , n28080 , n1285 );
    or g27216 ( n11622 , n14446 , n12622 );
    nor g27217 ( n29496 , n22457 , n33956 );
    and g27218 ( n29468 , n2712 , n12903 );
    xnor g27219 ( n29786 , n21129 , n4288 );
    or g27220 ( n25631 , n31691 , n6550 );
    or g27221 ( n5225 , n28818 , n12622 );
    xnor g27222 ( n11445 , n13336 , n29913 );
    not g27223 ( n32528 , n9864 );
    and g27224 ( n13211 , n17493 , n30001 );
    or g27225 ( n26497 , n9962 , n12724 );
    xnor g27226 ( n24496 , n6063 , n20515 );
    and g27227 ( n16075 , n9348 , n32252 );
    and g27228 ( n10420 , n17411 , n28069 );
    or g27229 ( n11717 , n14038 , n20512 );
    or g27230 ( n30863 , n27230 , n28455 );
    nor g27231 ( n29264 , n14871 , n4508 );
    or g27232 ( n30822 , n6324 , n9207 );
    not g27233 ( n26129 , n20577 );
    or g27234 ( n25966 , n25729 , n17337 );
    and g27235 ( n30027 , n11072 , n6910 );
    or g27236 ( n20857 , n5299 , n13480 );
    and g27237 ( n20821 , n17921 , n29793 );
    not g27238 ( n10510 , n25030 );
    xnor g27239 ( n2515 , n23746 , n1831 );
    and g27240 ( n35080 , n20771 , n7555 );
    and g27241 ( n32950 , n4413 , n28484 );
    xnor g27242 ( n8123 , n18487 , n24789 );
    and g27243 ( n16137 , n15331 , n17088 );
    nor g27244 ( n17844 , n9798 , n34423 );
    or g27245 ( n14668 , n14547 , n34528 );
    and g27246 ( n9338 , n25439 , n15853 );
    or g27247 ( n5232 , n26127 , n31331 );
    or g27248 ( n11978 , n32857 , n1204 );
    xnor g27249 ( n32885 , n3218 , n15886 );
    and g27250 ( n26003 , n30532 , n5200 );
    or g27251 ( n14267 , n27627 , n2235 );
    xnor g27252 ( n25157 , n749 , n24785 );
    xnor g27253 ( n14124 , n17548 , n31796 );
    xnor g27254 ( n28278 , n11306 , n30937 );
    or g27255 ( n793 , n3222 , n18574 );
    not g27256 ( n10423 , n15096 );
    and g27257 ( n21758 , n26435 , n21270 );
    or g27258 ( n24916 , n16160 , n23689 );
    xnor g27259 ( n10881 , n24626 , n7540 );
    or g27260 ( n4822 , n6933 , n28363 );
    xnor g27261 ( n3603 , n12696 , n33224 );
    or g27262 ( n5853 , n8720 , n2538 );
    or g27263 ( n19987 , n7746 , n20817 );
    or g27264 ( n11679 , n12048 , n10340 );
    or g27265 ( n16506 , n32764 , n2416 );
    or g27266 ( n6088 , n19889 , n32644 );
    or g27267 ( n15467 , n5670 , n32425 );
    and g27268 ( n34183 , n8782 , n29538 );
    or g27269 ( n30454 , n5384 , n26051 );
    not g27270 ( n29249 , n31799 );
    or g27271 ( n23783 , n30809 , n25831 );
    and g27272 ( n30769 , n31079 , n829 );
    not g27273 ( n30617 , n8637 );
    or g27274 ( n12356 , n4568 , n35630 );
    or g27275 ( n20380 , n20993 , n500 );
    or g27276 ( n23635 , n20426 , n13215 );
    or g27277 ( n22345 , n10472 , n33098 );
    xnor g27278 ( n14156 , n29903 , n14697 );
    or g27279 ( n7676 , n15644 , n1792 );
    or g27280 ( n25290 , n4857 , n7417 );
    or g27281 ( n7329 , n5803 , n1474 );
    or g27282 ( n25979 , n10099 , n7417 );
    or g27283 ( n33572 , n3984 , n15713 );
    or g27284 ( n14862 , n23040 , n35748 );
    xnor g27285 ( n11572 , n10300 , n382 );
    and g27286 ( n2076 , n10023 , n11121 );
    or g27287 ( n18210 , n14528 , n4305 );
    not g27288 ( n7429 , n144 );
    or g27289 ( n30295 , n31046 , n5611 );
    xnor g27290 ( n9481 , n22202 , n19551 );
    or g27291 ( n3261 , n22612 , n225 );
    or g27292 ( n27681 , n33968 , n23089 );
    or g27293 ( n14830 , n19551 , n78 );
    xnor g27294 ( n2467 , n5559 , n19867 );
    or g27295 ( n35987 , n17647 , n17543 );
    xnor g27296 ( n18062 , n27823 , n33744 );
    nor g27297 ( n2864 , n15886 , n32417 );
    buf g27298 ( n9930 , n13523 );
    and g27299 ( n25611 , n35536 , n31118 );
    or g27300 ( n23358 , n5091 , n16919 );
    and g27301 ( n34970 , n5842 , n602 );
    or g27302 ( n21883 , n12661 , n23327 );
    and g27303 ( n1833 , n21932 , n16745 );
    and g27304 ( n9693 , n28525 , n33021 );
    or g27305 ( n35946 , n10894 , n9192 );
    or g27306 ( n14178 , n22974 , n15805 );
    or g27307 ( n11137 , n20038 , n25773 );
    xnor g27308 ( n1960 , n24700 , n12162 );
    nor g27309 ( n31575 , n2764 , n27126 );
    not g27310 ( n25799 , n1504 );
    not g27311 ( n6220 , n28783 );
    nor g27312 ( n23111 , n29037 , n7251 );
    and g27313 ( n15308 , n32905 , n32760 );
    buf g27314 ( n28273 , n29437 );
    xnor g27315 ( n17953 , n9683 , n22869 );
    nor g27316 ( n9498 , n12341 , n28669 );
    xnor g27317 ( n12707 , n17587 , n11190 );
    or g27318 ( n17779 , n2264 , n28668 );
    and g27319 ( n16974 , n3881 , n22431 );
    xnor g27320 ( n6898 , n8706 , n2746 );
    and g27321 ( n31220 , n12147 , n14876 );
    or g27322 ( n1952 , n212 , n25831 );
    or g27323 ( n26276 , n31069 , n30646 );
    and g27324 ( n1130 , n8830 , n33687 );
    or g27325 ( n1092 , n1811 , n6529 );
    or g27326 ( n33378 , n16992 , n17829 );
    or g27327 ( n31224 , n19551 , n5122 );
    nor g27328 ( n26900 , n25602 , n3977 );
    or g27329 ( n24812 , n24371 , n35789 );
    or g27330 ( n12309 , n27341 , n1549 );
    and g27331 ( n10010 , n26020 , n6878 );
    not g27332 ( n8993 , n30306 );
    not g27333 ( n3069 , n24441 );
    xnor g27334 ( n22421 , n12698 , n29783 );
    xnor g27335 ( n5231 , n10955 , n2157 );
    xnor g27336 ( n32840 , n17750 , n15886 );
    not g27337 ( n15486 , n3805 );
    and g27338 ( n31143 , n6065 , n17255 );
    and g27339 ( n35042 , n222 , n21563 );
    or g27340 ( n5680 , n28549 , n13305 );
    not g27341 ( n26347 , n3205 );
    and g27342 ( n7808 , n9868 , n7959 );
    or g27343 ( n12148 , n1738 , n12913 );
    or g27344 ( n14370 , n24298 , n3395 );
    or g27345 ( n1578 , n33061 , n12244 );
    or g27346 ( n20014 , n24698 , n14699 );
    and g27347 ( n3629 , n14431 , n14378 );
    xnor g27348 ( n5070 , n24727 , n27813 );
    xnor g27349 ( n1749 , n2575 , n15403 );
    not g27350 ( n1609 , n22980 );
    or g27351 ( n280 , n28796 , n14746 );
    xnor g27352 ( n13505 , n30659 , n32715 );
    xnor g27353 ( n1357 , n27249 , n22572 );
    or g27354 ( n22910 , n4733 , n17872 );
    xnor g27355 ( n14694 , n14788 , n4960 );
    and g27356 ( n30066 , n5904 , n19473 );
    and g27357 ( n27352 , n7953 , n6030 );
    or g27358 ( n8527 , n4401 , n34600 );
    not g27359 ( n14639 , n36033 );
    or g27360 ( n31342 , n32095 , n31114 );
    xnor g27361 ( n1584 , n25644 , n12778 );
    and g27362 ( n5695 , n5988 , n10740 );
    and g27363 ( n14946 , n21794 , n7409 );
    or g27364 ( n34435 , n958 , n16762 );
    xnor g27365 ( n16626 , n15502 , n21266 );
    or g27366 ( n21006 , n34212 , n9317 );
    or g27367 ( n32480 , n31605 , n31638 );
    or g27368 ( n28664 , n7540 , n31792 );
    nor g27369 ( n29743 , n14593 , n4024 );
    not g27370 ( n25511 , n11830 );
    nor g27371 ( n20200 , n17163 , n29830 );
    xnor g27372 ( n23926 , n24411 , n35927 );
    or g27373 ( n15161 , n15886 , n15565 );
    and g27374 ( n23382 , n5051 , n24796 );
    xnor g27375 ( n35958 , n4616 , n27859 );
    not g27376 ( n3808 , n35490 );
    not g27377 ( n35029 , n20070 );
    or g27378 ( n22901 , n13659 , n9479 );
    and g27379 ( n2253 , n28245 , n4326 );
    nor g27380 ( n31046 , n3946 , n13677 );
    and g27381 ( n16980 , n8788 , n3782 );
    or g27382 ( n2260 , n17763 , n11381 );
    and g27383 ( n19876 , n11717 , n13538 );
    or g27384 ( n20756 , n13783 , n8851 );
    xnor g27385 ( n3819 , n27525 , n27121 );
    xnor g27386 ( n20235 , n30438 , n28652 );
    not g27387 ( n24011 , n22980 );
    or g27388 ( n13757 , n19483 , n15344 );
    and g27389 ( n4606 , n24184 , n23041 );
    and g27390 ( n2636 , n35014 , n26204 );
    or g27391 ( n1921 , n21354 , n25392 );
    and g27392 ( n7250 , n2924 , n3839 );
    xnor g27393 ( n28405 , n22311 , n7679 );
    or g27394 ( n25892 , n28182 , n11833 );
    or g27395 ( n30598 , n2358 , n27053 );
    or g27396 ( n3831 , n24225 , n25761 );
    or g27397 ( n13549 , n28001 , n16532 );
    xnor g27398 ( n10731 , n11349 , n25201 );
    nor g27399 ( n5034 , n24371 , n18180 );
    not g27400 ( n8490 , n3842 );
    xnor g27401 ( n32530 , n22223 , n23820 );
    and g27402 ( n29408 , n34401 , n3451 );
    or g27403 ( n13173 , n13533 , n29077 );
    or g27404 ( n4071 , n25539 , n31883 );
    xnor g27405 ( n14402 , n12348 , n24801 );
    or g27406 ( n18169 , n881 , n27778 );
    or g27407 ( n15232 , n32747 , n15145 );
    and g27408 ( n32465 , n24571 , n693 );
    and g27409 ( n24265 , n36017 , n22980 );
    or g27410 ( n7225 , n4191 , n13094 );
    or g27411 ( n32455 , n9288 , n949 );
    or g27412 ( n7377 , n15747 , n13478 );
    or g27413 ( n6826 , n25228 , n27262 );
    or g27414 ( n22511 , n16470 , n11475 );
    or g27415 ( n5595 , n31306 , n30867 );
    or g27416 ( n8815 , n15482 , n9338 );
    xnor g27417 ( n58 , n4178 , n6651 );
    xnor g27418 ( n10799 , n187 , n4763 );
    xnor g27419 ( n8819 , n22321 , n24371 );
    or g27420 ( n34316 , n29839 , n16240 );
    xnor g27421 ( n28639 , n19852 , n5186 );
    or g27422 ( n12776 , n4995 , n18649 );
    or g27423 ( n21480 , n3205 , n2636 );
    or g27424 ( n23448 , n3222 , n7484 );
    not g27425 ( n3951 , n16177 );
    xnor g27426 ( n12277 , n14284 , n31289 );
    not g27427 ( n7446 , n32329 );
    or g27428 ( n12496 , n4419 , n28837 );
    or g27429 ( n15913 , n15157 , n17233 );
    or g27430 ( n35448 , n29884 , n14567 );
    or g27431 ( n8077 , n34982 , n9118 );
    xnor g27432 ( n18053 , n18370 , n5145 );
    nor g27433 ( n28251 , n17992 , n22097 );
    xnor g27434 ( n21048 , n866 , n16307 );
    or g27435 ( n23917 , n13409 , n15894 );
    or g27436 ( n20412 , n24776 , n15145 );
    and g27437 ( n17226 , n24452 , n9004 );
    xnor g27438 ( n30525 , n19283 , n4962 );
    xnor g27439 ( n34053 , n31812 , n3946 );
    and g27440 ( n26424 , n23036 , n401 );
    or g27441 ( n26395 , n35348 , n10632 );
    xnor g27442 ( n29935 , n23923 , n34739 );
    not g27443 ( n11463 , n29839 );
    and g27444 ( n6414 , n18605 , n3269 );
    and g27445 ( n32143 , n25969 , n27881 );
    or g27446 ( n14030 , n22075 , n4172 );
    and g27447 ( n13714 , n29938 , n29369 );
    or g27448 ( n274 , n26847 , n16297 );
    or g27449 ( n32002 , n10040 , n12123 );
    or g27450 ( n29532 , n16028 , n31464 );
    or g27451 ( n6897 , n3562 , n30382 );
    and g27452 ( n33996 , n9458 , n25100 );
    or g27453 ( n1599 , n13201 , n30832 );
    or g27454 ( n15622 , n8439 , n16979 );
    nor g27455 ( n12123 , n16819 , n1230 );
    or g27456 ( n29550 , n21965 , n3736 );
    nor g27457 ( n3227 , n4288 , n16415 );
    xnor g27458 ( n1676 , n21463 , n10894 );
    or g27459 ( n14819 , n11324 , n31368 );
    or g27460 ( n18086 , n30214 , n28404 );
    or g27461 ( n30242 , n21413 , n34600 );
    or g27462 ( n4201 , n2242 , n31922 );
    and g27463 ( n33689 , n9258 , n7246 );
    xnor g27464 ( n30435 , n20363 , n13076 );
    or g27465 ( n4211 , n830 , n34030 );
    and g27466 ( n6061 , n19299 , n20165 );
    xnor g27467 ( n24231 , n10163 , n35692 );
    xnor g27468 ( n18430 , n5936 , n22294 );
    xnor g27469 ( n5608 , n18082 , n22271 );
    nor g27470 ( n9956 , n16620 , n32964 );
    xnor g27471 ( n29358 , n18538 , n16272 );
    or g27472 ( n34869 , n27539 , n9921 );
    or g27473 ( n34841 , n4280 , n21585 );
    or g27474 ( n18771 , n26177 , n19084 );
    or g27475 ( n5331 , n9331 , n3805 );
    or g27476 ( n10118 , n25563 , n31514 );
    or g27477 ( n26133 , n1613 , n8282 );
    and g27478 ( n18039 , n19986 , n14304 );
    or g27479 ( n28951 , n6741 , n8723 );
    and g27480 ( n25263 , n19399 , n22918 );
    or g27481 ( n23227 , n5872 , n5223 );
    and g27482 ( n10276 , n34362 , n27577 );
    and g27483 ( n10752 , n6650 , n11427 );
    or g27484 ( n35095 , n66 , n31514 );
    or g27485 ( n16515 , n8224 , n14361 );
    xnor g27486 ( n11096 , n23514 , n16357 );
    or g27487 ( n24097 , n3607 , n16525 );
    or g27488 ( n25667 , n31311 , n35168 );
    and g27489 ( n30707 , n34649 , n18642 );
    or g27490 ( n14134 , n25602 , n22505 );
    xnor g27491 ( n20413 , n6765 , n29384 );
    not g27492 ( n21892 , n18073 );
    or g27493 ( n8897 , n12601 , n1557 );
    xor g27494 ( n35508 , n8610 , n3287 );
    or g27495 ( n2687 , n35152 , n27243 );
    xnor g27496 ( n6557 , n14042 , n24004 );
    and g27497 ( n885 , n10474 , n29704 );
    or g27498 ( n3642 , n24725 , n4460 );
    or g27499 ( n35045 , n7073 , n25594 );
    and g27500 ( n12149 , n6071 , n10327 );
    or g27501 ( n10722 , n471 , n7308 );
    and g27502 ( n21808 , n3823 , n12504 );
    and g27503 ( n9579 , n36002 , n34608 );
    or g27504 ( n21027 , n7075 , n1373 );
    or g27505 ( n3273 , n24042 , n32276 );
    and g27506 ( n8344 , n4046 , n10051 );
    xnor g27507 ( n2624 , n15527 , n8923 );
    or g27508 ( n15530 , n21702 , n27580 );
    and g27509 ( n14399 , n34863 , n31941 );
    and g27510 ( n8890 , n13232 , n2348 );
    xnor g27511 ( n25222 , n20159 , n9155 );
    or g27512 ( n10534 , n8124 , n13933 );
    xnor g27513 ( n4977 , n9349 , n32897 );
    or g27514 ( n20105 , n2269 , n26220 );
    or g27515 ( n32751 , n357 , n21042 );
    and g27516 ( n26457 , n23401 , n35959 );
    xnor g27517 ( n15574 , n30772 , n1950 );
    xnor g27518 ( n2961 , n34492 , n15937 );
    or g27519 ( n12942 , n7590 , n2562 );
    xnor g27520 ( n15545 , n28929 , n11752 );
    or g27521 ( n27790 , n1334 , n5618 );
    xnor g27522 ( n5409 , n18534 , n21342 );
    or g27523 ( n31711 , n22382 , n29003 );
    xnor g27524 ( n20416 , n9878 , n16922 );
    or g27525 ( n7790 , n23079 , n15109 );
    or g27526 ( n35612 , n15403 , n14437 );
    xnor g27527 ( n6719 , n15066 , n35927 );
    nor g27528 ( n4555 , n32243 , n8002 );
    or g27529 ( n12416 , n18100 , n4293 );
    or g27530 ( n14416 , n34742 , n4318 );
    xnor g27531 ( n4414 , n6817 , n29839 );
    or g27532 ( n8782 , n27540 , n1484 );
    xnor g27533 ( n30460 , n10099 , n3205 );
    or g27534 ( n653 , n19412 , n16149 );
    or g27535 ( n14257 , n33309 , n8203 );
    nor g27536 ( n31214 , n30742 , n32515 );
    xnor g27537 ( n14325 , n32041 , n21061 );
    xnor g27538 ( n7263 , n28802 , n33924 );
    nor g27539 ( n9747 , n28384 , n11179 );
    or g27540 ( n1074 , n486 , n23438 );
    and g27541 ( n3136 , n15916 , n6948 );
    or g27542 ( n17739 , n32095 , n8623 );
    not g27543 ( n10206 , n35257 );
    or g27544 ( n35735 , n32267 , n3188 );
    not g27545 ( n13651 , n2597 );
    or g27546 ( n28826 , n23418 , n25355 );
    xnor g27547 ( n16159 , n12015 , n10894 );
    xnor g27548 ( n27228 , n1787 , n9504 );
    nor g27549 ( n21074 , n27451 , n14889 );
    or g27550 ( n11277 , n14379 , n25036 );
    and g27551 ( n1436 , n22921 , n24616 );
    xnor g27552 ( n23161 , n10454 , n29059 );
    or g27553 ( n9412 , n24198 , n5505 );
    or g27554 ( n20230 , n9019 , n27801 );
    or g27555 ( n6041 , n34671 , n3465 );
    not g27556 ( n8325 , n28457 );
    xnor g27557 ( n6317 , n9095 , n19281 );
    and g27558 ( n1560 , n13257 , n13296 );
    or g27559 ( n3899 , n1950 , n32338 );
    or g27560 ( n9573 , n30369 , n19939 );
    and g27561 ( n256 , n35201 , n14894 );
    xnor g27562 ( n2369 , n3913 , n16402 );
    not g27563 ( n6968 , n20348 );
    xnor g27564 ( n34962 , n27896 , n35663 );
    not g27565 ( n34367 , n32857 );
    or g27566 ( n6544 , n34041 , n1715 );
    or g27567 ( n8189 , n5523 , n23748 );
    or g27568 ( n31618 , n25170 , n29411 );
    and g27569 ( n2991 , n34721 , n33638 );
    or g27570 ( n16507 , n14667 , n3239 );
    and g27571 ( n10601 , n7372 , n6702 );
    and g27572 ( n24698 , n18836 , n17712 );
    xnor g27573 ( n33949 , n8142 , n17446 );
    or g27574 ( n21122 , n31272 , n19604 );
    or g27575 ( n27520 , n15403 , n8215 );
    xnor g27576 ( n23570 , n18018 , n281 );
    nor g27577 ( n27482 , n16699 , n16649 );
    or g27578 ( n19298 , n32603 , n29626 );
    or g27579 ( n25741 , n29945 , n33248 );
    and g27580 ( n7261 , n8739 , n1065 );
    buf g27581 ( n15256 , n21862 );
    nor g27582 ( n21813 , n12414 , n9921 );
    and g27583 ( n10593 , n23659 , n20436 );
    or g27584 ( n14505 , n14267 , n12428 );
    xnor g27585 ( n10521 , n14021 , n19992 );
    and g27586 ( n5887 , n24023 , n19770 );
    not g27587 ( n9092 , n6507 );
    and g27588 ( n23165 , n13993 , n14321 );
    or g27589 ( n23950 , n17805 , n19084 );
    xnor g27590 ( n2066 , n11488 , n31799 );
    xnor g27591 ( n21470 , n26724 , n29609 );
    and g27592 ( n3263 , n25667 , n13860 );
    xnor g27593 ( n31867 , n32685 , n35927 );
    xnor g27594 ( n18941 , n22953 , n5287 );
    and g27595 ( n31236 , n34321 , n20362 );
    or g27596 ( n3586 , n201 , n2005 );
    not g27597 ( n31448 , n32857 );
    or g27598 ( n25353 , n7029 , n3352 );
    and g27599 ( n4898 , n11655 , n20186 );
    or g27600 ( n17491 , n22251 , n5779 );
    or g27601 ( n13593 , n15299 , n28463 );
    xnor g27602 ( n28221 , n19073 , n15958 );
    and g27603 ( n28361 , n20767 , n17789 );
    or g27604 ( n17017 , n30942 , n3239 );
    or g27605 ( n33239 , n12915 , n14746 );
    or g27606 ( n31543 , n25149 , n763 );
    and g27607 ( n31345 , n1104 , n3245 );
    and g27608 ( n32457 , n11092 , n13871 );
    or g27609 ( n2014 , n27554 , n19732 );
    and g27610 ( n31739 , n26982 , n7508 );
    not g27611 ( n23122 , n11633 );
    xnor g27612 ( n34072 , n3455 , n26779 );
    and g27613 ( n28222 , n5300 , n31010 );
    or g27614 ( n22415 , n25215 , n16594 );
    not g27615 ( n26510 , n26532 );
    and g27616 ( n3281 , n23714 , n22423 );
    or g27617 ( n21085 , n28393 , n28064 );
    or g27618 ( n25017 , n34364 , n9879 );
    xnor g27619 ( n747 , n2394 , n18103 );
    and g27620 ( n10161 , n34593 , n9681 );
    xnor g27621 ( n4287 , n6437 , n5335 );
    or g27622 ( n25693 , n16800 , n28248 );
    or g27623 ( n34828 , n29884 , n21200 );
    or g27624 ( n20693 , n32668 , n22682 );
    and g27625 ( n20620 , n921 , n9397 );
    or g27626 ( n9254 , n22658 , n15572 );
    or g27627 ( n5019 , n7674 , n26339 );
    and g27628 ( n8293 , n25670 , n34123 );
    or g27629 ( n16303 , n27542 , n7162 );
    or g27630 ( n27888 , n23314 , n24559 );
    or g27631 ( n5381 , n35368 , n1102 );
    or g27632 ( n2445 , n15985 , n22322 );
    not g27633 ( n12734 , n34142 );
    nor g27634 ( n28087 , n27291 , n15022 );
    or g27635 ( n22438 , n29623 , n33320 );
    nor g27636 ( n7413 , n3205 , n1135 );
    and g27637 ( n5717 , n8842 , n19262 );
    xnor g27638 ( n16634 , n25082 , n4501 );
    or g27639 ( n8874 , n31469 , n16464 );
    or g27640 ( n30068 , n9105 , n1642 );
    or g27641 ( n21656 , n34155 , n28668 );
    xnor g27642 ( n28049 , n25118 , n1118 );
    or g27643 ( n17556 , n12017 , n17046 );
    xnor g27644 ( n22948 , n21852 , n13077 );
    or g27645 ( n32376 , n17568 , n29519 );
    or g27646 ( n31308 , n25835 , n1557 );
    not g27647 ( n33921 , n8902 );
    or g27648 ( n27867 , n3033 , n26002 );
    or g27649 ( n3476 , n11000 , n26881 );
    xnor g27650 ( n19085 , n11147 , n32095 );
    or g27651 ( n17936 , n34113 , n3239 );
    xnor g27652 ( n6011 , n34972 , n35519 );
    xnor g27653 ( n1786 , n11315 , n7125 );
    or g27654 ( n11491 , n11159 , n19173 );
    xor g27655 ( n1830 , n3168 , n6731 );
    xnor g27656 ( n15301 , n19319 , n31559 );
    xnor g27657 ( n28026 , n17246 , n29839 );
    or g27658 ( n3588 , n18469 , n34600 );
    or g27659 ( n31871 , n32253 , n17162 );
    and g27660 ( n16105 , n4613 , n35158 );
    not g27661 ( n27740 , n23089 );
    or g27662 ( n8011 , n27713 , n10908 );
    nor g27663 ( n28703 , n20443 , n15645 );
    or g27664 ( n5270 , n33348 , n4478 );
    and g27665 ( n10933 , n5073 , n15891 );
    nor g27666 ( n2711 , n8432 , n12581 );
    or g27667 ( n17680 , n9568 , n27188 );
    xnor g27668 ( n30747 , n17830 , n6485 );
    nor g27669 ( n10896 , n23986 , n33956 );
    and g27670 ( n20191 , n28193 , n5057 );
    nor g27671 ( n9168 , n31799 , n18144 );
    xnor g27672 ( n10724 , n14648 , n29098 );
    or g27673 ( n15160 , n5312 , n36000 );
    or g27674 ( n21626 , n14353 , n24299 );
    xnor g27675 ( n24807 , n20550 , n18728 );
    or g27676 ( n27387 , n5522 , n12288 );
    or g27677 ( n33786 , n19526 , n18976 );
    or g27678 ( n33344 , n2207 , n23260 );
    or g27679 ( n5325 , n8899 , n31055 );
    xnor g27680 ( n29467 , n3423 , n22677 );
    or g27681 ( n11 , n23444 , n5752 );
    or g27682 ( n11036 , n22291 , n11509 );
    not g27683 ( n15329 , n15873 );
    or g27684 ( n22508 , n10560 , n24778 );
    or g27685 ( n10598 , n254 , n23921 );
    xnor g27686 ( n24432 , n6254 , n32715 );
    and g27687 ( n2749 , n24813 , n31708 );
    nor g27688 ( n20405 , n17568 , n14865 );
    or g27689 ( n34112 , n12429 , n29818 );
    and g27690 ( n18027 , n11429 , n24181 );
    or g27691 ( n9382 , n23493 , n19490 );
    not g27692 ( n30999 , n26720 );
    or g27693 ( n34659 , n9407 , n15344 );
    xnor g27694 ( n7887 , n33011 , n32857 );
    nor g27695 ( n29212 , n15722 , n16649 );
    xnor g27696 ( n9611 , n30062 , n31799 );
    xnor g27697 ( n6060 , n10008 , n11474 );
    or g27698 ( n10015 , n25430 , n1402 );
    xnor g27699 ( n32992 , n5421 , n35927 );
    and g27700 ( n28737 , n13801 , n19551 );
    or g27701 ( n27749 , n25471 , n17962 );
    or g27702 ( n19017 , n1903 , n34865 );
    xnor g27703 ( n9757 , n27378 , n20280 );
    not g27704 ( n12329 , n16026 );
    or g27705 ( n29691 , n28683 , n10762 );
    or g27706 ( n35274 , n30742 , n12938 );
    or g27707 ( n25884 , n187 , n4763 );
    or g27708 ( n12366 , n15886 , n20873 );
    xnor g27709 ( n18905 , n34228 , n8968 );
    and g27710 ( n31163 , n3301 , n10726 );
    or g27711 ( n18435 , n1628 , n25907 );
    and g27712 ( n12054 , n32258 , n15462 );
    and g27713 ( n2728 , n23496 , n15014 );
    or g27714 ( n26857 , n13717 , n25023 );
    or g27715 ( n28679 , n27291 , n8294 );
    or g27716 ( n26681 , n15403 , n2548 );
    or g27717 ( n12635 , n25702 , n15496 );
    xnor g27718 ( n18796 , n19668 , n11455 );
    not g27719 ( n25951 , n4960 );
    and g27720 ( n8913 , n21883 , n21356 );
    or g27721 ( n14062 , n35354 , n19336 );
    nor g27722 ( n26442 , n31672 , n23024 );
    or g27723 ( n16460 , n30125 , n31161 );
    or g27724 ( n3175 , n4758 , n5242 );
    or g27725 ( n28627 , n35615 , n24779 );
    or g27726 ( n24970 , n9842 , n27454 );
    or g27727 ( n18822 , n9524 , n24758 );
    and g27728 ( n19217 , n12291 , n10565 );
    and g27729 ( n26258 , n24804 , n22384 );
    or g27730 ( n8510 , n15330 , n6950 );
    xnor g27731 ( n1537 , n26234 , n12250 );
    xnor g27732 ( n10639 , n16539 , n11046 );
    or g27733 ( n29088 , n17240 , n10872 );
    and g27734 ( n18858 , n21573 , n11819 );
    xnor g27735 ( n11858 , n9417 , n13210 );
    not g27736 ( n22757 , n27069 );
    or g27737 ( n28724 , n1581 , n9592 );
    and g27738 ( n24746 , n28437 , n16036 );
    and g27739 ( n35792 , n5006 , n19308 );
    and g27740 ( n3568 , n34484 , n26810 );
    or g27741 ( n31530 , n11046 , n34664 );
    and g27742 ( n29699 , n11124 , n18910 );
    and g27743 ( n2501 , n29674 , n16147 );
    or g27744 ( n25153 , n21167 , n20377 );
    or g27745 ( n30273 , n13632 , n5470 );
    or g27746 ( n18693 , n7744 , n14887 );
    and g27747 ( n21970 , n28540 , n7611 );
    or g27748 ( n3621 , n23133 , n15256 );
    or g27749 ( n5246 , n16431 , n9202 );
    nor g27750 ( n13093 , n19768 , n18115 );
    xnor g27751 ( n3488 , n14786 , n35794 );
    not g27752 ( n28632 , n10527 );
    and g27753 ( n12951 , n27970 , n25364 );
    or g27754 ( n2530 , n7716 , n28324 );
    or g27755 ( n33972 , n16290 , n27043 );
    nor g27756 ( n26648 , n22790 , n833 );
    nor g27757 ( n15536 , n15097 , n23614 );
    or g27758 ( n22258 , n12043 , n26834 );
    or g27759 ( n34171 , n24322 , n29174 );
    or g27760 ( n17309 , n15209 , n17905 );
    and g27761 ( n29334 , n25593 , n32082 );
    or g27762 ( n15446 , n25066 , n3694 );
    or g27763 ( n10141 , n32857 , n22649 );
    xnor g27764 ( n2252 , n20256 , n18643 );
    xnor g27765 ( n19307 , n27289 , n29409 );
    or g27766 ( n24426 , n8931 , n10593 );
    nor g27767 ( n10701 , n31391 , n15809 );
    or g27768 ( n15384 , n22335 , n19892 );
    and g27769 ( n16696 , n26934 , n23975 );
    xnor g27770 ( n18022 , n28431 , n29839 );
    or g27771 ( n12818 , n32811 , n5868 );
    nor g27772 ( n28842 , n8357 , n12864 );
    xnor g27773 ( n29265 , n34152 , n31799 );
    or g27774 ( n30583 , n8121 , n23650 );
    xnor g27775 ( n35385 , n31693 , n6236 );
    or g27776 ( n27862 , n5600 , n23090 );
    or g27777 ( n11387 , n22311 , n7679 );
    and g27778 ( n15479 , n34015 , n22451 );
    and g27779 ( n18416 , n26075 , n6343 );
    or g27780 ( n25562 , n15736 , n6139 );
    xnor g27781 ( n13763 , n24331 , n16922 );
    and g27782 ( n25839 , n26231 , n10117 );
    xnor g27783 ( n473 , n17258 , n19551 );
    xnor g27784 ( n26854 , n25536 , n8376 );
    not g27785 ( n443 , n12428 );
    nor g27786 ( n26897 , n18934 , n31606 );
    or g27787 ( n14013 , n22939 , n20797 );
    xnor g27788 ( n11630 , n28151 , n29899 );
    and g27789 ( n13971 , n34230 , n26629 );
    not g27790 ( n36005 , n4962 );
    or g27791 ( n16496 , n8096 , n1476 );
    or g27792 ( n30641 , n164 , n2340 );
    xnor g27793 ( n9245 , n17899 , n22575 );
    or g27794 ( n33386 , n29242 , n585 );
    or g27795 ( n20102 , n25162 , n32507 );
    xnor g27796 ( n3305 , n7273 , n27325 );
    xnor g27797 ( n36040 , n10294 , n16620 );
    and g27798 ( n12142 , n19024 , n18187 );
    or g27799 ( n7456 , n31799 , n13601 );
    and g27800 ( n316 , n31613 , n32287 );
    xnor g27801 ( n5350 , n4807 , n19551 );
    or g27802 ( n13232 , n12928 , n32071 );
    not g27803 ( n463 , n14140 );
    or g27804 ( n29753 , n14571 , n3352 );
    nor g27805 ( n15445 , n27572 , n2912 );
    xnor g27806 ( n15449 , n9605 , n34011 );
    and g27807 ( n21941 , n25962 , n17369 );
    and g27808 ( n5039 , n4270 , n9492 );
    and g27809 ( n11058 , n35389 , n26741 );
    or g27810 ( n27173 , n32286 , n16464 );
    xnor g27811 ( n20662 , n7424 , n759 );
    and g27812 ( n29515 , n1675 , n4506 );
    or g27813 ( n28812 , n19650 , n21977 );
    or g27814 ( n6391 , n11455 , n35307 );
    or g27815 ( n13049 , n36009 , n29835 );
    xnor g27816 ( n22290 , n12544 , n4029 );
    or g27817 ( n31950 , n35951 , n23748 );
    or g27818 ( n35442 , n32715 , n20059 );
    not g27819 ( n23072 , n19952 );
    xnor g27820 ( n910 , n6367 , n8867 );
    or g27821 ( n18607 , n3162 , n10336 );
    nor g27822 ( n26051 , n3955 , n17657 );
    or g27823 ( n8626 , n2915 , n17675 );
    or g27824 ( n12313 , n12991 , n2955 );
    or g27825 ( n24436 , n9441 , n6374 );
    xnor g27826 ( n11330 , n33460 , n27291 );
    or g27827 ( n1835 , n32113 , n26730 );
    xnor g27828 ( n3955 , n16703 , n19984 );
    and g27829 ( n16884 , n487 , n17857 );
    buf g27830 ( n25940 , n17046 );
    or g27831 ( n5775 , n34444 , n5607 );
    and g27832 ( n29108 , n3655 , n13272 );
    and g27833 ( n33271 , n13535 , n8976 );
    and g27834 ( n16240 , n9473 , n16127 );
    or g27835 ( n22839 , n17548 , n31796 );
    and g27836 ( n32063 , n24367 , n21156 );
    or g27837 ( n18465 , n4918 , n12332 );
    not g27838 ( n11818 , n15597 );
    xnor g27839 ( n12934 , n13411 , n10894 );
    or g27840 ( n29721 , n3565 , n29366 );
    and g27841 ( n33476 , n23184 , n24203 );
    not g27842 ( n7087 , n17568 );
    xnor g27843 ( n22251 , n18875 , n27453 );
    nor g27844 ( n34046 , n11422 , n19834 );
    or g27845 ( n32652 , n1352 , n5538 );
    and g27846 ( n9882 , n34457 , n16430 );
    and g27847 ( n20194 , n25125 , n11895 );
    nor g27848 ( n9815 , n33717 , n13019 );
    not g27849 ( n828 , n10946 );
    xnor g27850 ( n12461 , n30124 , n3946 );
    not g27851 ( n21351 , n1950 );
    or g27852 ( n31798 , n16135 , n17250 );
    xnor g27853 ( n32267 , n14374 , n14949 );
    nor g27854 ( n32206 , n10199 , n6548 );
    or g27855 ( n5594 , n4288 , n24919 );
    or g27856 ( n11842 , n9793 , n27675 );
    or g27857 ( n7959 , n32857 , n33011 );
    nor g27858 ( n7228 , n9146 , n16934 );
    and g27859 ( n2047 , n23610 , n6585 );
    or g27860 ( n18792 , n23120 , n15577 );
    or g27861 ( n32488 , n28690 , n11518 );
    or g27862 ( n31346 , n29713 , n17736 );
    or g27863 ( n34465 , n5304 , n1642 );
    and g27864 ( n7346 , n27382 , n28884 );
    xnor g27865 ( n875 , n24161 , n3205 );
    or g27866 ( n14556 , n4288 , n18668 );
    and g27867 ( n31780 , n20737 , n2917 );
    and g27868 ( n32644 , n2672 , n5253 );
    or g27869 ( n6234 , n11455 , n12782 );
    not g27870 ( n3829 , n21737 );
    or g27871 ( n19037 , n31812 , n3694 );
    or g27872 ( n31814 , n11033 , n4508 );
    and g27873 ( n7079 , n22786 , n19948 );
    or g27874 ( n31891 , n25079 , n20139 );
    or g27875 ( n17595 , n10560 , n15178 );
    or g27876 ( n14092 , n18453 , n11351 );
    and g27877 ( n33397 , n34171 , n23398 );
    nor g27878 ( n32498 , n15464 , n25384 );
    and g27879 ( n32227 , n25641 , n28910 );
    or g27880 ( n33258 , n11455 , n36087 );
    or g27881 ( n29419 , n31215 , n16105 );
    or g27882 ( n1084 , n10983 , n31725 );
    or g27883 ( n19400 , n21355 , n22970 );
    nor g27884 ( n1314 , n34278 , n205 );
    and g27885 ( n34708 , n457 , n19620 );
    xnor g27886 ( n22665 , n22686 , n32857 );
    or g27887 ( n12831 , n19041 , n4664 );
    not g27888 ( n4069 , n7834 );
    or g27889 ( n31047 , n4905 , n25447 );
    or g27890 ( n4591 , n8470 , n19953 );
    or g27891 ( n21333 , n30064 , n28743 );
    or g27892 ( n4959 , n5476 , n34923 );
    or g27893 ( n21016 , n24941 , n31606 );
    or g27894 ( n13724 , n14461 , n4291 );
    and g27895 ( n11747 , n18526 , n7561 );
    or g27896 ( n27661 , n13922 , n16919 );
    and g27897 ( n26089 , n2382 , n16661 );
    nor g27898 ( n1405 , n24002 , n33917 );
    or g27899 ( n12361 , n9126 , n24489 );
    and g27900 ( n30144 , n26713 , n24724 );
    not g27901 ( n9706 , n16555 );
    xnor g27902 ( n8628 , n22340 , n33542 );
    or g27903 ( n19846 , n5263 , n8366 );
    or g27904 ( n17666 , n29839 , n27688 );
    and g27905 ( n9075 , n33215 , n8900 );
    nor g27906 ( n29939 , n16620 , n24892 );
    and g27907 ( n20284 , n30166 , n25498 );
    xnor g27908 ( n339 , n20334 , n15034 );
    or g27909 ( n6501 , n30442 , n24560 );
    or g27910 ( n15628 , n21296 , n31549 );
    xnor g27911 ( n6616 , n1343 , n32584 );
    or g27912 ( n6320 , n29839 , n27021 );
    nor g27913 ( n15135 , n18224 , n14224 );
    or g27914 ( n2321 , n9494 , n14554 );
    or g27915 ( n13989 , n29543 , n15109 );
    not g27916 ( n30615 , n22980 );
    and g27917 ( n4525 , n22833 , n32882 );
    or g27918 ( n28101 , n36035 , n6459 );
    and g27919 ( n2256 , n17090 , n26546 );
    or g27920 ( n1544 , n23960 , n5457 );
    and g27921 ( n17742 , n16498 , n11129 );
    xnor g27922 ( n4935 , n5423 , n31272 );
    and g27923 ( n16087 , n31353 , n17540 );
    or g27924 ( n2160 , n8285 , n5058 );
    xnor g27925 ( n35074 , n4194 , n11012 );
    xnor g27926 ( n33982 , n21121 , n19664 );
    or g27927 ( n11176 , n31492 , n21956 );
    or g27928 ( n27726 , n19645 , n15144 );
    and g27929 ( n12507 , n19655 , n2574 );
    and g27930 ( n29603 , n34163 , n20950 );
    or g27931 ( n9018 , n27208 , n31514 );
    or g27932 ( n4944 , n6252 , n12742 );
    xnor g27933 ( n112 , n35760 , n28362 );
    and g27934 ( n34707 , n32144 , n32222 );
    xnor g27935 ( n12736 , n15247 , n11409 );
    and g27936 ( n22953 , n6926 , n633 );
    nor g27937 ( n3721 , n25602 , n23098 );
    not g27938 ( n32194 , n35938 );
    or g27939 ( n17822 , n14809 , n9295 );
    xnor g27940 ( n7716 , n30746 , n27518 );
    and g27941 ( n19590 , n22450 , n19253 );
    or g27942 ( n22983 , n5802 , n34600 );
    and g27943 ( n27465 , n5817 , n22360 );
    or g27944 ( n29505 , n27783 , n28541 );
    or g27945 ( n14796 , n8778 , n11833 );
    and g27946 ( n16139 , n34653 , n18639 );
    xnor g27947 ( n4993 , n20418 , n17559 );
    xnor g27948 ( n3542 , n7906 , n5287 );
    not g27949 ( n17757 , n891 );
    and g27950 ( n22967 , n1395 , n34565 );
    or g27951 ( n31408 , n34844 , n13664 );
    and g27952 ( n5460 , n11563 , n8734 );
    or g27953 ( n1523 , n31289 , n14284 );
    or g27954 ( n7642 , n13683 , n9067 );
    nor g27955 ( n18380 , n11046 , n397 );
    not g27956 ( n11511 , n28273 );
    or g27957 ( n27618 , n16812 , n5252 );
    xnor g27958 ( n31943 , n22511 , n5455 );
    or g27959 ( n25517 , n1230 , n13408 );
    and g27960 ( n16671 , n1475 , n2951 );
    xnor g27961 ( n31634 , n15111 , n31595 );
    xnor g27962 ( n20793 , n19537 , n35927 );
    nor g27963 ( n20714 , n20079 , n23086 );
    buf g27964 ( n17974 , n34865 );
    xnor g27965 ( n14495 , n30415 , n32857 );
    and g27966 ( n20966 , n25654 , n18629 );
    xnor g27967 ( n16350 , n21072 , n21880 );
    and g27968 ( n16733 , n14764 , n5109 );
    and g27969 ( n18151 , n16345 , n1629 );
    or g27970 ( n21376 , n10466 , n25761 );
    and g27971 ( n11963 , n2972 , n21622 );
    nor g27972 ( n24365 , n4758 , n15498 );
    and g27973 ( n21851 , n15803 , n10502 );
    xnor g27974 ( n7150 , n23900 , n28846 );
    xnor g27975 ( n22541 , n33701 , n17568 );
    or g27976 ( n13373 , n25539 , n34272 );
    and g27977 ( n29441 , n5668 , n23581 );
    and g27978 ( n12385 , n5947 , n8032 );
    and g27979 ( n8586 , n20472 , n33160 );
    and g27980 ( n21753 , n6066 , n33432 );
    or g27981 ( n31529 , n29509 , n27728 );
    and g27982 ( n14298 , n22887 , n12795 );
    xnor g27983 ( n674 , n35349 , n33462 );
    or g27984 ( n33753 , n8330 , n13400 );
    or g27985 ( n6155 , n8771 , n27053 );
    or g27986 ( n17561 , n7540 , n27925 );
    nor g27987 ( n33503 , n32095 , n10149 );
    not g27988 ( n17559 , n16922 );
    xnor g27989 ( n34640 , n12257 , n26979 );
    and g27990 ( n13099 , n31444 , n5688 );
    or g27991 ( n311 , n18291 , n29106 );
    and g27992 ( n3100 , n20653 , n31454 );
    nor g27993 ( n22826 , n8332 , n9921 );
    and g27994 ( n29759 , n5809 , n30534 );
    or g27995 ( n10699 , n3212 , n16843 );
    xnor g27996 ( n11606 , n15649 , n4960 );
    or g27997 ( n30503 , n15855 , n17281 );
    buf g27998 ( n27447 , n22501 );
    or g27999 ( n7718 , n5818 , n30364 );
    or g28000 ( n29483 , n13089 , n33674 );
    and g28001 ( n14271 , n30060 , n11317 );
    or g28002 ( n25623 , n10710 , n10762 );
    or g28003 ( n30740 , n23334 , n30646 );
    not g28004 ( n19031 , n33428 );
    nor g28005 ( n11209 , n19483 , n31677 );
    xnor g28006 ( n10817 , n8715 , n934 );
    nor g28007 ( n9023 , n16922 , n5243 );
    and g28008 ( n15928 , n17428 , n32282 );
    nor g28009 ( n6104 , n25118 , n7454 );
    or g28010 ( n349 , n4960 , n7742 );
    or g28011 ( n28333 , n9789 , n21457 );
    not g28012 ( n23404 , n3819 );
    xnor g28013 ( n4389 , n30045 , n4962 );
    or g28014 ( n14549 , n18768 , n25019 );
    not g28015 ( n24345 , n2433 );
    or g28016 ( n27762 , n4758 , n35097 );
    xnor g28017 ( n17096 , n35772 , n4288 );
    xnor g28018 ( n1276 , n6848 , n528 );
    nor g28019 ( n24701 , n29504 , n33140 );
    xnor g28020 ( n15473 , n15804 , n4878 );
    and g28021 ( n32304 , n28303 , n26034 );
    and g28022 ( n33950 , n22032 , n15181 );
    not g28023 ( n5679 , n18955 );
    xnor g28024 ( n12467 , n24630 , n12566 );
    or g28025 ( n14048 , n22578 , n7417 );
    buf g28026 ( n16326 , n2791 );
    xnor g28027 ( n25430 , n9465 , n29228 );
    not g28028 ( n29256 , n34380 );
    nor g28029 ( n35315 , n10668 , n30444 );
    or g28030 ( n20753 , n4288 , n11415 );
    or g28031 ( n7278 , n25223 , n22322 );
    or g28032 ( n17371 , n31215 , n25742 );
    nor g28033 ( n1502 , n3205 , n2509 );
    or g28034 ( n8113 , n23008 , n14918 );
    not g28035 ( n21224 , n22980 );
    not g28036 ( n26590 , n20558 );
    not g28037 ( n33606 , n4960 );
    xnor g28038 ( n26758 , n9367 , n29713 );
    not g28039 ( n30098 , n30565 );
    or g28040 ( n5055 , n32695 , n6340 );
    or g28041 ( n19234 , n29713 , n9367 );
    and g28042 ( n22720 , n754 , n9215 );
    and g28043 ( n16547 , n12641 , n12623 );
    nor g28044 ( n27589 , n30742 , n22690 );
    and g28045 ( n32799 , n13774 , n756 );
    nor g28046 ( n33741 , n18462 , n2580 );
    and g28047 ( n8921 , n32942 , n32193 );
    or g28048 ( n23005 , n12011 , n24499 );
    xnor g28049 ( n34448 , n4629 , n22926 );
    xnor g28050 ( n30866 , n25862 , n14441 );
    xnor g28051 ( n31371 , n13097 , n11046 );
    and g28052 ( n33582 , n4012 , n11792 );
    and g28053 ( n32385 , n5574 , n20113 );
    or g28054 ( n12691 , n33898 , n4952 );
    nor g28055 ( n7407 , n4878 , n17526 );
    not g28056 ( n28926 , n35927 );
    or g28057 ( n16765 , n23406 , n31134 );
    and g28058 ( n5584 , n22706 , n29181 );
    or g28059 ( n33092 , n7263 , n16919 );
    not g28060 ( n18512 , n7726 );
    or g28061 ( n33659 , n23604 , n19791 );
    or g28062 ( n27331 , n15617 , n9072 );
    and g28063 ( n2994 , n15770 , n7294 );
    or g28064 ( n9369 , n28123 , n28668 );
    xnor g28065 ( n17972 , n16733 , n30742 );
    xnor g28066 ( n35489 , n26474 , n13113 );
    and g28067 ( n25764 , n33614 , n35499 );
    xnor g28068 ( n9060 , n26869 , n1917 );
    not g28069 ( n6511 , n13498 );
    or g28070 ( n26735 , n23604 , n17285 );
    or g28071 ( n29523 , n3931 , n9915 );
    and g28072 ( n13229 , n18951 , n4628 );
    and g28073 ( n22024 , n30284 , n30236 );
    not g28074 ( n13477 , n3205 );
    xnor g28075 ( n4634 , n19750 , n9793 );
    or g28076 ( n34133 , n21267 , n31549 );
    and g28077 ( n19581 , n12321 , n14117 );
    buf g28078 ( n11703 , n11712 );
    xnor g28079 ( n23857 , n17785 , n19551 );
    and g28080 ( n5117 , n12068 , n27837 );
    and g28081 ( n427 , n13722 , n19207 );
    xnor g28082 ( n27022 , n9416 , n4584 );
    or g28083 ( n32784 , n34172 , n25773 );
    xnor g28084 ( n18820 , n23237 , n18445 );
    xnor g28085 ( n35576 , n5301 , n21531 );
    and g28086 ( n30682 , n21833 , n18553 );
    not g28087 ( n22113 , n4542 );
    xnor g28088 ( n12181 , n1235 , n12419 );
    or g28089 ( n12571 , n9652 , n19403 );
    and g28090 ( n970 , n35106 , n31288 );
    xnor g28091 ( n5040 , n1277 , n31334 );
    xnor g28092 ( n33704 , n13629 , n1950 );
    and g28093 ( n32404 , n10015 , n4563 );
    or g28094 ( n2377 , n2516 , n17726 );
    or g28095 ( n34807 , n12855 , n7237 );
    xnor g28096 ( n28820 , n20511 , n15886 );
    not g28097 ( n34680 , n2471 );
    xnor g28098 ( n377 , n6616 , n34250 );
    or g28099 ( n537 , n32465 , n23209 );
    not g28100 ( n11461 , n19147 );
    not g28101 ( n5450 , n30457 );
    or g28102 ( n9188 , n23134 , n14076 );
    xnor g28103 ( n28372 , n29487 , n24129 );
    and g28104 ( n17415 , n185 , n24474 );
    or g28105 ( n10875 , n27751 , n6017 );
    or g28106 ( n24674 , n29032 , n10301 );
    or g28107 ( n14715 , n31289 , n5178 );
    nor g28108 ( n9080 , n17568 , n19395 );
    or g28109 ( n33980 , n12092 , n9864 );
    or g28110 ( n21194 , n33844 , n24025 );
    or g28111 ( n25434 , n32664 , n28364 );
    xnor g28112 ( n4220 , n21045 , n1950 );
    xnor g28113 ( n3939 , n35060 , n12876 );
    xnor g28114 ( n22287 , n27961 , n25471 );
    not g28115 ( n33368 , n19939 );
    or g28116 ( n2328 , n6368 , n3651 );
    or g28117 ( n35819 , n16922 , n3455 );
    nor g28118 ( n31548 , n4960 , n1525 );
    or g28119 ( n8727 , n34514 , n1826 );
    xnor g28120 ( n19669 , n7223 , n19971 );
    xnor g28121 ( n1803 , n23400 , n5532 );
    xnor g28122 ( n17146 , n4835 , n21459 );
    xnor g28123 ( n18920 , n12155 , n11046 );
    xnor g28124 ( n20250 , n6719 , n4057 );
    and g28125 ( n31863 , n9633 , n22852 );
    xnor g28126 ( n21666 , n4301 , n32095 );
    or g28127 ( n19299 , n26624 , n5403 );
    or g28128 ( n27676 , n5447 , n34097 );
    or g28129 ( n13599 , n34044 , n27355 );
    and g28130 ( n23850 , n14587 , n6379 );
    or g28131 ( n13405 , n1033 , n11772 );
    or g28132 ( n8318 , n27636 , n713 );
    and g28133 ( n14101 , n33664 , n26777 );
    or g28134 ( n17272 , n839 , n25306 );
    and g28135 ( n25612 , n26413 , n31132 );
    or g28136 ( n5244 , n35423 , n13425 );
    or g28137 ( n9719 , n13220 , n31148 );
    not g28138 ( n9260 , n29976 );
    xnor g28139 ( n10247 , n16176 , n151 );
    not g28140 ( n35800 , n15886 );
    or g28141 ( n30284 , n33156 , n17535 );
    or g28142 ( n27792 , n31650 , n7680 );
    nor g28143 ( n13720 , n33057 , n29294 );
    not g28144 ( n10207 , n30326 );
    or g28145 ( n9138 , n6054 , n17962 );
    and g28146 ( n16471 , n29182 , n6281 );
    or g28147 ( n8117 , n4960 , n34463 );
    or g28148 ( n17188 , n9411 , n12503 );
    nor g28149 ( n9074 , n26428 , n27511 );
    xnor g28150 ( n5693 , n23500 , n18283 );
    or g28151 ( n32172 , n23245 , n29393 );
    or g28152 ( n25824 , n14144 , n11897 );
    or g28153 ( n1294 , n22291 , n13537 );
    or g28154 ( n29154 , n13037 , n13305 );
    xnor g28155 ( n16253 , n11825 , n15886 );
    and g28156 ( n7763 , n7810 , n31157 );
    and g28157 ( n31492 , n16592 , n25947 );
    nor g28158 ( n4191 , n7540 , n17082 );
    xnor g28159 ( n33046 , n639 , n16922 );
    or g28160 ( n33203 , n35197 , n908 );
    or g28161 ( n28346 , n8439 , n16326 );
    xnor g28162 ( n25577 , n23091 , n3228 );
    and g28163 ( n7894 , n11622 , n28301 );
    xnor g28164 ( n23971 , n10306 , n5287 );
    buf g28165 ( n11295 , n9003 );
    or g28166 ( n31059 , n35000 , n32572 );
    xnor g28167 ( n8641 , n15720 , n7230 );
    or g28168 ( n20983 , n11906 , n20252 );
    nor g28169 ( n7381 , n5086 , n25701 );
    nor g28170 ( n29072 , n22356 , n7167 );
    or g28171 ( n790 , n28334 , n20364 );
    and g28172 ( n2572 , n4737 , n7012 );
    or g28173 ( n8394 , n25174 , n19972 );
    and g28174 ( n10181 , n31142 , n23293 );
    xnor g28175 ( n13069 , n20531 , n10573 );
    or g28176 ( n20433 , n25174 , n16490 );
    not g28177 ( n10548 , n25392 );
    and g28178 ( n34810 , n8189 , n1623 );
    xnor g28179 ( n21738 , n2352 , n25174 );
    or g28180 ( n20231 , n31056 , n27880 );
    or g28181 ( n11006 , n32095 , n7708 );
    and g28182 ( n33170 , n27042 , n26302 );
    not g28183 ( n5298 , n31665 );
    or g28184 ( n16003 , n16955 , n19261 );
    and g28185 ( n24529 , n26148 , n5007 );
    or g28186 ( n17656 , n10491 , n5005 );
    nor g28187 ( n32711 , n17568 , n26464 );
    not g28188 ( n24954 , n22980 );
    and g28189 ( n34767 , n2756 , n18031 );
    or g28190 ( n30823 , n5297 , n29411 );
    xnor g28191 ( n31146 , n6361 , n557 );
    or g28192 ( n33062 , n35546 , n12206 );
    and g28193 ( n28190 , n3361 , n35421 );
    nor g28194 ( n16889 , n9793 , n8513 );
    or g28195 ( n12576 , n15173 , n5900 );
    buf g28196 ( n27641 , n27144 );
    buf g28197 ( n3842 , n28497 );
    or g28198 ( n3620 , n24121 , n1404 );
    or g28199 ( n34917 , n425 , n20318 );
    or g28200 ( n16492 , n31799 , n6392 );
    or g28201 ( n29997 , n18908 , n27665 );
    xnor g28202 ( n16475 , n1905 , n20099 );
    or g28203 ( n18605 , n1448 , n2825 );
    and g28204 ( n35933 , n34182 , n15929 );
    and g28205 ( n29535 , n12849 , n17824 );
    xnor g28206 ( n6918 , n5243 , n17559 );
    or g28207 ( n18359 , n24332 , n29884 );
    and g28208 ( n20854 , n9732 , n27115 );
    nor g28209 ( n24714 , n1842 , n15144 );
    or g28210 ( n12579 , n3946 , n27742 );
    or g28211 ( n27071 , n11992 , n5189 );
    or g28212 ( n2557 , n5335 , n27552 );
    xnor g28213 ( n7777 , n1172 , n9658 );
    or g28214 ( n3264 , n32933 , n22954 );
    nor g28215 ( n1240 , n26027 , n2242 );
    or g28216 ( n30338 , n20671 , n2005 );
    and g28217 ( n32393 , n31892 , n2679 );
    or g28218 ( n20220 , n1428 , n22206 );
    and g28219 ( n9413 , n3208 , n14686 );
    nor g28220 ( n17648 , n5335 , n26751 );
    or g28221 ( n29245 , n15464 , n35324 );
    or g28222 ( n15879 , n18763 , n5779 );
    xnor g28223 ( n24768 , n27596 , n4962 );
    or g28224 ( n10546 , n13292 , n15497 );
    and g28225 ( n16959 , n13604 , n17688 );
    or g28226 ( n18842 , n20976 , n5602 );
    nor g28227 ( n33720 , n21814 , n3581 );
    not g28228 ( n6465 , n31722 );
    xnor g28229 ( n6003 , n10401 , n8913 );
    nor g28230 ( n20086 , n35879 , n18115 );
    not g28231 ( n7851 , n3205 );
    or g28232 ( n31510 , n7484 , n23209 );
    or g28233 ( n30639 , n15800 , n34634 );
    buf g28234 ( n3480 , n29437 );
    or g28235 ( n20505 , n5287 , n7906 );
    and g28236 ( n19972 , n28983 , n3439 );
    xnor g28237 ( n5481 , n15616 , n32669 );
    xnor g28238 ( n7036 , n3123 , n8765 );
    xnor g28239 ( n28966 , n30049 , n32584 );
    nor g28240 ( n8665 , n31054 , n22422 );
    and g28241 ( n20091 , n8590 , n19782 );
    or g28242 ( n31916 , n41 , n24869 );
    or g28243 ( n16932 , n549 , n28240 );
    or g28244 ( n9785 , n22453 , n27619 );
    and g28245 ( n10145 , n35272 , n23799 );
    xnor g28246 ( n35892 , n14782 , n3592 );
    xnor g28247 ( n26159 , n19178 , n5465 );
    xnor g28248 ( n30475 , n9926 , n10769 );
    or g28249 ( n8729 , n5248 , n35141 );
    and g28250 ( n30433 , n7617 , n716 );
    or g28251 ( n1223 , n6272 , n9488 );
    xnor g28252 ( n24834 , n27676 , n27291 );
    or g28253 ( n32547 , n32992 , n29241 );
    or g28254 ( n25599 , n20564 , n32063 );
    or g28255 ( n964 , n20987 , n11833 );
    xnor g28256 ( n12387 , n19829 , n4962 );
    xnor g28257 ( n1998 , n23126 , n15772 );
    and g28258 ( n19645 , n25092 , n29234 );
    or g28259 ( n13240 , n9658 , n16715 );
    and g28260 ( n23916 , n16226 , n6739 );
    xnor g28261 ( n9740 , n30501 , n33850 );
    and g28262 ( n8274 , n7394 , n7218 );
    nor g28263 ( n24485 , n21430 , n25343 );
    or g28264 ( n18179 , n13894 , n8105 );
    and g28265 ( n21923 , n27146 , n31448 );
    xnor g28266 ( n10664 , n9918 , n5335 );
    xnor g28267 ( n4018 , n8651 , n17664 );
    or g28268 ( n18556 , n31466 , n13635 );
    and g28269 ( n21974 , n35134 , n8395 );
    or g28270 ( n23073 , n5165 , n7734 );
    and g28271 ( n3009 , n5038 , n31836 );
    and g28272 ( n34205 , n25248 , n11052 );
    xnor g28273 ( n28810 , n27953 , n3192 );
    or g28274 ( n11948 , n17568 , n5552 );
    not g28275 ( n18972 , n12642 );
    and g28276 ( n23920 , n33637 , n13761 );
    not g28277 ( n5137 , n11046 );
    and g28278 ( n2918 , n2971 , n3578 );
    or g28279 ( n22136 , n31289 , n28835 );
    not g28280 ( n7744 , n26522 );
    xnor g28281 ( n30759 , n25798 , n25146 );
    xnor g28282 ( n5727 , n30705 , n13393 );
    or g28283 ( n17386 , n8357 , n8265 );
    not g28284 ( n19571 , n31217 );
    xnor g28285 ( n5559 , n29693 , n24332 );
    and g28286 ( n26439 , n8615 , n27595 );
    or g28287 ( n29087 , n14827 , n29592 );
    or g28288 ( n5330 , n26510 , n22192 );
    or g28289 ( n32583 , n24350 , n29998 );
    not g28290 ( n18638 , n15886 );
    xnor g28291 ( n16678 , n19948 , n35437 );
    or g28292 ( n1644 , n31694 , n17068 );
    and g28293 ( n4485 , n35412 , n19894 );
    not g28294 ( n21731 , n22980 );
    or g28295 ( n33939 , n20289 , n10487 );
    and g28296 ( n31467 , n31579 , n24975 );
    and g28297 ( n17002 , n12199 , n10513 );
    not g28298 ( n17560 , n35927 );
    not g28299 ( n24108 , n22856 );
    and g28300 ( n9816 , n18879 , n5734 );
    xnor g28301 ( n31932 , n32446 , n11046 );
    and g28302 ( n32067 , n18896 , n24239 );
    or g28303 ( n7681 , n7292 , n1414 );
    or g28304 ( n20003 , n13396 , n26199 );
    or g28305 ( n24445 , n32657 , n13328 );
    not g28306 ( n31472 , n25861 );
    and g28307 ( n11409 , n25890 , n32499 );
    or g28308 ( n32283 , n9325 , n26112 );
    not g28309 ( n5470 , n17068 );
    xnor g28310 ( n30713 , n15477 , n33767 );
    not g28311 ( n6383 , n4878 );
    xnor g28312 ( n36055 , n22114 , n19928 );
    xnor g28313 ( n13683 , n23494 , n11455 );
    or g28314 ( n25365 , n28661 , n26365 );
    xnor g28315 ( n35120 , n17194 , n18103 );
    and g28316 ( n10199 , n13800 , n26506 );
    nor g28317 ( n33561 , n23127 , n31699 );
    or g28318 ( n31474 , n32053 , n14732 );
    xnor g28319 ( n15631 , n33646 , n11577 );
    or g28320 ( n16795 , n10816 , n31451 );
    or g28321 ( n4891 , n3222 , n11315 );
    and g28322 ( n6627 , n27311 , n33526 );
    not g28323 ( n3581 , n13651 );
    xnor g28324 ( n25803 , n26317 , n23604 );
    and g28325 ( n9066 , n29344 , n30740 );
    xnor g28326 ( n20855 , n10396 , n4444 );
    xnor g28327 ( n11719 , n21454 , n965 );
    nor g28328 ( n19889 , n4288 , n12841 );
    nor g28329 ( n16610 , n21733 , n23089 );
    not g28330 ( n23655 , n11996 );
    or g28331 ( n30106 , n23604 , n32935 );
    not g28332 ( n25214 , n9005 );
    xnor g28333 ( n26013 , n1740 , n29713 );
    not g28334 ( n28730 , n15886 );
    xnor g28335 ( n12006 , n11276 , n3515 );
    or g28336 ( n31045 , n5286 , n6683 );
    nor g28337 ( n18929 , n20775 , n8981 );
    and g28338 ( n6463 , n8918 , n20421 );
    xnor g28339 ( n13773 , n8703 , n4962 );
    and g28340 ( n16310 , n20778 , n21979 );
    nor g28341 ( n5735 , n31799 , n8719 );
    or g28342 ( n9223 , n91 , n19336 );
    or g28343 ( n35439 , n32857 , n30415 );
    buf g28344 ( n27704 , n32434 );
    nor g28345 ( n14889 , n34713 , n12010 );
    not g28346 ( n1162 , n15095 );
    or g28347 ( n4567 , n29839 , n4176 );
    or g28348 ( n31623 , n33668 , n763 );
    buf g28349 ( n5168 , n17184 );
    xnor g28350 ( n30285 , n32967 , n4998 );
    or g28351 ( n5797 , n19587 , n7553 );
    xnor g28352 ( n5341 , n16310 , n35927 );
    buf g28353 ( n13900 , n21418 );
    or g28354 ( n20743 , n24187 , n1560 );
    or g28355 ( n6585 , n19692 , n26023 );
    not g28356 ( n309 , n26811 );
    xnor g28357 ( n31862 , n21040 , n17568 );
    and g28358 ( n1725 , n4802 , n13531 );
    and g28359 ( n25065 , n28380 , n8367 );
    or g28360 ( n31208 , n31375 , n35935 );
    not g28361 ( n36088 , n3025 );
    or g28362 ( n33686 , n5335 , n28901 );
    xnor g28363 ( n19679 , n25118 , n10758 );
    xnor g28364 ( n444 , n770 , n33353 );
    xnor g28365 ( n21171 , n6559 , n4960 );
    or g28366 ( n3549 , n6656 , n35422 );
    buf g28367 ( n2104 , n28675 );
    xnor g28368 ( n30722 , n19468 , n25976 );
    xnor g28369 ( n35112 , n13612 , n24679 );
    or g28370 ( n25260 , n22543 , n23086 );
    or g28371 ( n16131 , n16935 , n26512 );
    and g28372 ( n14299 , n33784 , n3494 );
    or g28373 ( n16823 , n6643 , n16457 );
    xnor g28374 ( n17942 , n31157 , n7810 );
    xnor g28375 ( n1507 , n7822 , n7961 );
    buf g28376 ( n25036 , n13343 );
    or g28377 ( n7927 , n34262 , n9316 );
    and g28378 ( n33803 , n28523 , n29263 );
    xnor g28379 ( n6762 , n4908 , n6825 );
    or g28380 ( n11398 , n11190 , n30130 );
    or g28381 ( n11909 , n27362 , n13015 );
    and g28382 ( n35699 , n27882 , n31319 );
    or g28383 ( n35548 , n10943 , n2104 );
    xnor g28384 ( n24016 , n1259 , n34347 );
    or g28385 ( n11316 , n27880 , n15256 );
    xnor g28386 ( n16880 , n33301 , n7540 );
    xnor g28387 ( n31841 , n10367 , n35927 );
    or g28388 ( n34304 , n19570 , n19553 );
    or g28389 ( n35688 , n3222 , n19606 );
    and g28390 ( n12703 , n14419 , n31817 );
    xnor g28391 ( n28811 , n25357 , n1465 );
    nor g28392 ( n5393 , n21218 , n25588 );
    or g28393 ( n33745 , n11639 , n16137 );
    or g28394 ( n14790 , n4962 , n1903 );
    or g28395 ( n8342 , n30637 , n1402 );
    or g28396 ( n11383 , n20727 , n28675 );
    xnor g28397 ( n16158 , n2625 , n11046 );
    or g28398 ( n28547 , n6332 , n4490 );
    nor g28399 ( n1558 , n309 , n4856 );
    xnor g28400 ( n14848 , n28608 , n19551 );
    or g28401 ( n35642 , n22871 , n17029 );
    or g28402 ( n32271 , n5049 , n4715 );
    or g28403 ( n32112 , n15923 , n18416 );
    xnor g28404 ( n19855 , n4212 , n7008 );
    not g28405 ( n18274 , n15799 );
    and g28406 ( n10267 , n7860 , n24637 );
    or g28407 ( n32630 , n14374 , n14949 );
    and g28408 ( n7853 , n26655 , n12917 );
    nor g28409 ( n5206 , n9789 , n22574 );
    or g28410 ( n28677 , n31843 , n11218 );
    and g28411 ( n3561 , n32435 , n17912 );
    and g28412 ( n5286 , n3412 , n11516 );
    or g28413 ( n8378 , n10971 , n1265 );
    and g28414 ( n26319 , n33984 , n35823 );
    xnor g28415 ( n6062 , n31686 , n23046 );
    nor g28416 ( n22147 , n16536 , n28507 );
    or g28417 ( n7627 , n14802 , n30769 );
    or g28418 ( n22304 , n4962 , n24934 );
    and g28419 ( n8704 , n15225 , n1390 );
    or g28420 ( n34857 , n553 , n6323 );
    or g28421 ( n18329 , n101 , n33034 );
    or g28422 ( n10019 , n30675 , n33034 );
    not g28423 ( n7543 , n9793 );
    and g28424 ( n9528 , n13458 , n1842 );
    and g28425 ( n10978 , n33628 , n22650 );
    and g28426 ( n6666 , n23389 , n18452 );
    not g28427 ( n6178 , n30459 );
    xnor g28428 ( n17995 , n3379 , n3205 );
    or g28429 ( n8017 , n29589 , n19464 );
    or g28430 ( n25516 , n16135 , n17267 );
    or g28431 ( n27354 , n19551 , n30139 );
    not g28432 ( n4526 , n24463 );
    and g28433 ( n11034 , n27988 , n30778 );
    nor g28434 ( n18378 , n6663 , n27770 );
    xnor g28435 ( n11452 , n31525 , n15732 );
    or g28436 ( n36012 , n17751 , n3776 );
    xnor g28437 ( n14019 , n16933 , n26652 );
    or g28438 ( n25092 , n8214 , n15496 );
    or g28439 ( n3777 , n8641 , n35630 );
    and g28440 ( n8748 , n32078 , n13169 );
    xnor g28441 ( n29512 , n5644 , n16135 );
    and g28442 ( n5602 , n5571 , n1434 );
    xnor g28443 ( n19833 , n4898 , n4878 );
    or g28444 ( n28506 , n32095 , n11925 );
    or g28445 ( n30145 , n22178 , n23790 );
    and g28446 ( n3382 , n1577 , n26717 );
    and g28447 ( n14788 , n1589 , n30880 );
    or g28448 ( n17403 , n17568 , n3653 );
    or g28449 ( n35305 , n8084 , n12082 );
    and g28450 ( n29559 , n3963 , n20648 );
    xnor g28451 ( n29338 , n26090 , n29713 );
    or g28452 ( n20916 , n29144 , n27580 );
    or g28453 ( n24087 , n5361 , n17990 );
    or g28454 ( n27697 , n22843 , n17962 );
    xnor g28455 ( n33133 , n18706 , n9155 );
    not g28456 ( n20335 , n21313 );
    xnor g28457 ( n13308 , n19606 , n3222 );
    and g28458 ( n28953 , n2724 , n24524 );
    and g28459 ( n35720 , n13828 , n12308 );
    and g28460 ( n13246 , n19233 , n33627 );
    xnor g28461 ( n7885 , n35256 , n18899 );
    not g28462 ( n5709 , n8865 );
    not g28463 ( n12626 , n29872 );
    or g28464 ( n15934 , n31056 , n21258 );
    or g28465 ( n27150 , n23875 , n16609 );
    or g28466 ( n3655 , n35508 , n23790 );
    and g28467 ( n3002 , n25007 , n6544 );
    and g28468 ( n18632 , n21561 , n6029 );
    or g28469 ( n12477 , n32647 , n25903 );
    or g28470 ( n9771 , n11455 , n24468 );
    xnor g28471 ( n35552 , n25558 , n1479 );
    xnor g28472 ( n15918 , n22786 , n3946 );
    or g28473 ( n30912 , n29597 , n29562 );
    or g28474 ( n20581 , n29692 , n20862 );
    or g28475 ( n28387 , n6991 , n29366 );
    or g28476 ( n20027 , n3111 , n10616 );
    or g28477 ( n14764 , n4978 , n28324 );
    and g28478 ( n29433 , n26796 , n23903 );
    xnor g28479 ( n7137 , n12645 , n26018 );
    or g28480 ( n30262 , n8302 , n31684 );
    xnor g28481 ( n6322 , n3876 , n7540 );
    or g28482 ( n25358 , n29536 , n23921 );
    xnor g28483 ( n20444 , n14296 , n33544 );
    or g28484 ( n3550 , n20598 , n2168 );
    xnor g28485 ( n18419 , n11797 , n5556 );
    or g28486 ( n8741 , n14296 , n33544 );
    and g28487 ( n18080 , n953 , n7707 );
    xnor g28488 ( n16829 , n33434 , n16037 );
    xnor g28489 ( n31276 , n19248 , n4288 );
    xnor g28490 ( n1235 , n11617 , n9793 );
    or g28491 ( n31358 , n11739 , n14736 );
    xnor g28492 ( n11626 , n22734 , n24371 );
    xnor g28493 ( n28581 , n23018 , n14973 );
    nor g28494 ( n12476 , n30742 , n33996 );
    and g28495 ( n11333 , n22151 , n18774 );
    or g28496 ( n1292 , n17748 , n12913 );
    or g28497 ( n14804 , n28171 , n17068 );
    nor g28498 ( n5748 , n8432 , n9126 );
    or g28499 ( n20814 , n6331 , n35960 );
    or g28500 ( n9742 , n3194 , n7553 );
    and g28501 ( n7664 , n4167 , n10877 );
    or g28502 ( n15242 , n27319 , n5507 );
    and g28503 ( n30989 , n14898 , n25044 );
    buf g28504 ( n34472 , n12275 );
    xnor g28505 ( n20536 , n21598 , n29713 );
    and g28506 ( n12544 , n4932 , n29073 );
    not g28507 ( n5993 , n13983 );
    not g28508 ( n11106 , n7150 );
    not g28509 ( n614 , n17661 );
    and g28510 ( n10489 , n23214 , n21850 );
    and g28511 ( n8041 , n28515 , n27598 );
    not g28512 ( n5726 , n17875 );
    or g28513 ( n9177 , n28472 , n10432 );
    not g28514 ( n18989 , n9229 );
    and g28515 ( n1115 , n12359 , n27926 );
    or g28516 ( n2773 , n21507 , n5450 );
    and g28517 ( n32359 , n13804 , n5474 );
    xnor g28518 ( n18237 , n32549 , n23355 );
    or g28519 ( n12730 , n27107 , n24730 );
    nor g28520 ( n27924 , n31215 , n28501 );
    xnor g28521 ( n22941 , n14396 , n15611 );
    xnor g28522 ( n12628 , n19948 , n18675 );
    and g28523 ( n22701 , n22278 , n7624 );
    and g28524 ( n16837 , n11641 , n14556 );
    or g28525 ( n14823 , n35747 , n7436 );
    or g28526 ( n8565 , n6076 , n15145 );
    or g28527 ( n1797 , n9658 , n12163 );
    or g28528 ( n16148 , n31357 , n26292 );
    and g28529 ( n3156 , n24282 , n15821 );
    not g28530 ( n1552 , n35917 );
    or g28531 ( n35959 , n9658 , n13889 );
    or g28532 ( n5576 , n29570 , n4490 );
    or g28533 ( n7391 , n16922 , n17744 );
    or g28534 ( n25059 , n23813 , n2119 );
    not g28535 ( n22036 , n20558 );
    xnor g28536 ( n27135 , n6685 , n19551 );
    xnor g28537 ( n9266 , n19796 , n25602 );
    nor g28538 ( n3643 , n31242 , n19657 );
    or g28539 ( n33171 , n19654 , n29453 );
    not g28540 ( n1949 , n14850 );
    or g28541 ( n23143 , n32248 , n24745 );
    and g28542 ( n19928 , n515 , n3743 );
    not g28543 ( n34501 , n1323 );
    xnor g28544 ( n15650 , n5090 , n10769 );
    not g28545 ( n30421 , n31799 );
    or g28546 ( n12199 , n12640 , n11977 );
    nor g28547 ( n10826 , n27188 , n31411 );
    not g28548 ( n24148 , n24865 );
    and g28549 ( n21712 , n5902 , n26528 );
    or g28550 ( n19724 , n33887 , n11977 );
    xnor g28551 ( n29255 , n32113 , n26730 );
    and g28552 ( n17642 , n3206 , n29745 );
    and g28553 ( n20375 , n19823 , n5594 );
    and g28554 ( n28751 , n14185 , n16630 );
    xnor g28555 ( n17570 , n11369 , n35277 );
    or g28556 ( n612 , n3225 , n3633 );
    and g28557 ( n8609 , n26961 , n21292 );
    or g28558 ( n32413 , n28155 , n11601 );
    xnor g28559 ( n14150 , n18353 , n11190 );
    or g28560 ( n13440 , n10532 , n15068 );
    or g28561 ( n10879 , n11263 , n32746 );
    or g28562 ( n27153 , n10068 , n34040 );
    or g28563 ( n21474 , n31675 , n17337 );
    and g28564 ( n29383 , n28454 , n27380 );
    or g28565 ( n30927 , n30775 , n28668 );
    or g28566 ( n25682 , n10360 , n4203 );
    and g28567 ( n31994 , n14126 , n14174 );
    or g28568 ( n31975 , n18246 , n1097 );
    xnor g28569 ( n7033 , n8713 , n814 );
    or g28570 ( n2672 , n19043 , n27707 );
    xnor g28571 ( n5915 , n33285 , n9793 );
    or g28572 ( n33836 , n4878 , n13940 );
    xnor g28573 ( n33132 , n4322 , n556 );
    and g28574 ( n20516 , n20459 , n9654 );
    or g28575 ( n27993 , n23913 , n4952 );
    and g28576 ( n32431 , n6410 , n33409 );
    and g28577 ( n14643 , n3024 , n6706 );
    xnor g28578 ( n24931 , n13121 , n2326 );
    nor g28579 ( n19331 , n3946 , n1845 );
    not g28580 ( n3196 , n17029 );
    not g28581 ( n12402 , n10894 );
    or g28582 ( n12195 , n28774 , n25648 );
    or g28583 ( n32888 , n32715 , n812 );
    xnor g28584 ( n31120 , n24897 , n1950 );
    and g28585 ( n1168 , n19673 , n18028 );
    and g28586 ( n29994 , n12805 , n15481 );
    and g28587 ( n23466 , n16193 , n9166 );
    and g28588 ( n15577 , n14881 , n2925 );
    or g28589 ( n32147 , n1463 , n21514 );
    xnor g28590 ( n20633 , n25690 , n31559 );
    or g28591 ( n374 , n1332 , n27630 );
    or g28592 ( n1882 , n31289 , n9853 );
    and g28593 ( n21124 , n2553 , n22894 );
    or g28594 ( n20047 , n4962 , n17344 );
    not g28595 ( n29434 , n17568 );
    xnor g28596 ( n14194 , n20912 , n10894 );
    xnor g28597 ( n27879 , n2750 , n13023 );
    or g28598 ( n12719 , n20470 , n33389 );
    not g28599 ( n1981 , n29032 );
    or g28600 ( n10934 , n19551 , n31546 );
    xnor g28601 ( n59 , n16988 , n13949 );
    or g28602 ( n8410 , n5451 , n2712 );
    xnor g28603 ( n4920 , n12073 , n22751 );
    and g28604 ( n13845 , n32204 , n4112 );
    and g28605 ( n20870 , n15220 , n35338 );
    not g28606 ( n27876 , n6970 );
    or g28607 ( n31254 , n32857 , n10437 );
    xnor g28608 ( n27267 , n31925 , n17341 );
    or g28609 ( n2046 , n12242 , n33098 );
    xnor g28610 ( n34278 , n7365 , n18379 );
    or g28611 ( n17614 , n5287 , n9944 );
    and g28612 ( n25281 , n25540 , n17717 );
    and g28613 ( n1740 , n23413 , n32846 );
    and g28614 ( n3876 , n13772 , n23928 );
    or g28615 ( n2904 , n12445 , n21977 );
    or g28616 ( n12906 , n28518 , n31514 );
    or g28617 ( n8499 , n9793 , n10311 );
    or g28618 ( n14080 , n17568 , n35722 );
    not g28619 ( n20877 , n16922 );
    or g28620 ( n4145 , n7566 , n7553 );
    xnor g28621 ( n477 , n12962 , n5193 );
    or g28622 ( n24218 , n14110 , n24757 );
    or g28623 ( n26274 , n18098 , n9764 );
    xnor g28624 ( n18084 , n4782 , n12425 );
    and g28625 ( n32529 , n13185 , n27909 );
    xnor g28626 ( n27755 , n21857 , n35294 );
    or g28627 ( n14560 , n9259 , n34084 );
    xnor g28628 ( n33395 , n27077 , n7540 );
    or g28629 ( n33429 , n16811 , n15981 );
    or g28630 ( n21260 , n3282 , n30287 );
    or g28631 ( n5038 , n24602 , n28240 );
    and g28632 ( n35574 , n6157 , n33857 );
    and g28633 ( n21514 , n28024 , n1125 );
    and g28634 ( n17395 , n11832 , n17143 );
    xnor g28635 ( n20325 , n561 , n7096 );
    xnor g28636 ( n24783 , n12137 , n8041 );
    xnor g28637 ( n15141 , n23380 , n14308 );
    not g28638 ( n13678 , n21576 );
    xnor g28639 ( n3255 , n6573 , n18379 );
    not g28640 ( n25583 , n10336 );
    or g28641 ( n23357 , n28658 , n19787 );
    or g28642 ( n23905 , n6286 , n27501 );
    and g28643 ( n21370 , n3400 , n27752 );
    and g28644 ( n2774 , n17074 , n16057 );
    or g28645 ( n9029 , n5287 , n34530 );
    and g28646 ( n28592 , n12945 , n12675 );
    or g28647 ( n23588 , n24371 , n9758 );
    xnor g28648 ( n8818 , n24350 , n29998 );
    or g28649 ( n12214 , n16922 , n25368 );
    or g28650 ( n19641 , n21405 , n35143 );
    xnor g28651 ( n24617 , n10168 , n9658 );
    or g28652 ( n16466 , n22390 , n15249 );
    or g28653 ( n3666 , n33735 , n2757 );
    or g28654 ( n5247 , n32663 , n29769 );
    and g28655 ( n25814 , n19332 , n30765 );
    and g28656 ( n14209 , n2031 , n23289 );
    or g28657 ( n23440 , n28403 , n15067 );
    xnor g28658 ( n23569 , n14500 , n3458 );
    not g28659 ( n14018 , n35225 );
    or g28660 ( n15478 , n29748 , n34484 );
    or g28661 ( n29147 , n3946 , n18258 );
    not g28662 ( n26911 , n27633 );
    nor g28663 ( n27558 , n27560 , n25605 );
    xnor g28664 ( n17479 , n22353 , n27291 );
    or g28665 ( n24012 , n10894 , n11120 );
    and g28666 ( n5527 , n16862 , n6274 );
    and g28667 ( n15552 , n35771 , n4625 );
    nor g28668 ( n19327 , n7540 , n1567 );
    and g28669 ( n7229 , n10131 , n33071 );
    or g28670 ( n10046 , n29952 , n35748 );
    nor g28671 ( n16283 , n7255 , n19834 );
    or g28672 ( n24782 , n32744 , n3756 );
    and g28673 ( n2794 , n12528 , n354 );
    or g28674 ( n12811 , n20111 , n27010 );
    xnor g28675 ( n2663 , n22055 , n19228 );
    and g28676 ( n12741 , n8991 , n22314 );
    nor g28677 ( n6454 , n32857 , n3995 );
    and g28678 ( n20816 , n29937 , n5768 );
    or g28679 ( n13764 , n33920 , n18544 );
    xnor g28680 ( n34262 , n12358 , n31289 );
    xnor g28681 ( n21344 , n14464 , n1950 );
    and g28682 ( n28890 , n22214 , n18004 );
    or g28683 ( n26452 , n21680 , n20762 );
    xnor g28684 ( n24948 , n33136 , n30742 );
    or g28685 ( n17290 , n22236 , n28574 );
    or g28686 ( n8020 , n5152 , n35111 );
    xnor g28687 ( n5388 , n32936 , n31409 );
    xnor g28688 ( n35558 , n6027 , n11308 );
    and g28689 ( n8580 , n32353 , n2840 );
    xnor g28690 ( n9120 , n5609 , n15886 );
    xnor g28691 ( n28721 , n16234 , n30076 );
    or g28692 ( n25316 , n3205 , n14623 );
    xnor g28693 ( n25854 , n30975 , n31289 );
    or g28694 ( n10096 , n19398 , n30519 );
    and g28695 ( n418 , n31916 , n4966 );
    nor g28696 ( n15705 , n835 , n11934 );
    or g28697 ( n574 , n8801 , n8671 );
    or g28698 ( n10200 , n13929 , n12453 );
    or g28699 ( n32228 , n26424 , n33310 );
    and g28700 ( n11590 , n9405 , n27986 );
    xnor g28701 ( n26541 , n34356 , n1950 );
    and g28702 ( n2468 , n16964 , n8482 );
    or g28703 ( n34409 , n16922 , n30434 );
    not g28704 ( n9609 , n29722 );
    or g28705 ( n29632 , n5940 , n26219 );
    or g28706 ( n3216 , n4962 , n19829 );
    and g28707 ( n22929 , n19180 , n17661 );
    or g28708 ( n17646 , n11479 , n25832 );
    or g28709 ( n9512 , n28063 , n13307 );
    or g28710 ( n18089 , n19646 , n3805 );
    or g28711 ( n28555 , n21863 , n1606 );
    xnor g28712 ( n1055 , n18336 , n14072 );
    or g28713 ( n4205 , n16249 , n15538 );
    and g28714 ( n20488 , n33237 , n17727 );
    not g28715 ( n4531 , n8432 );
    or g28716 ( n2283 , n26033 , n34627 );
    xnor g28717 ( n26291 , n18202 , n13011 );
    or g28718 ( n20718 , n878 , n3437 );
    or g28719 ( n35957 , n27051 , n13516 );
    xnor g28720 ( n3914 , n14941 , n9104 );
    xnor g28721 ( n12306 , n13595 , n31799 );
    and g28722 ( n12545 , n7222 , n23096 );
    or g28723 ( n15042 , n6358 , n34289 );
    or g28724 ( n20036 , n27949 , n703 );
    or g28725 ( n12917 , n31302 , n30292 );
    xnor g28726 ( n21411 , n3623 , n6958 );
    or g28727 ( n6197 , n7011 , n29872 );
    or g28728 ( n3211 , n26704 , n5208 );
    xnor g28729 ( n23902 , n2646 , n32857 );
    or g28730 ( n18589 , n10759 , n2119 );
    xnor g28731 ( n17955 , n12483 , n35473 );
    not g28732 ( n18194 , n33317 );
    xnor g28733 ( n13775 , n13252 , n28329 );
    or g28734 ( n15803 , n35446 , n16298 );
    and g28735 ( n21603 , n22615 , n26886 );
    xnor g28736 ( n8368 , n18326 , n655 );
    and g28737 ( n29330 , n20874 , n32501 );
    nor g28738 ( n15981 , n6540 , n106 );
    or g28739 ( n23527 , n13333 , n14805 );
    or g28740 ( n5922 , n34150 , n24489 );
    and g28741 ( n31881 , n1780 , n9959 );
    and g28742 ( n2063 , n32979 , n24521 );
    and g28743 ( n8379 , n3319 , n11271 );
    or g28744 ( n35110 , n10771 , n3634 );
    not g28745 ( n14389 , n11276 );
    or g28746 ( n16378 , n21799 , n28969 );
    and g28747 ( n365 , n23358 , n2552 );
    or g28748 ( n21253 , n3723 , n10430 );
    and g28749 ( n9126 , n7093 , n21726 );
    or g28750 ( n15246 , n3048 , n6950 );
    xnor g28751 ( n16920 , n30092 , n4892 );
    xnor g28752 ( n22364 , n28026 , n31626 );
    not g28753 ( n4161 , n22200 );
    or g28754 ( n25496 , n23604 , n2619 );
    and g28755 ( n21071 , n31542 , n32696 );
    and g28756 ( n24018 , n25093 , n22343 );
    xnor g28757 ( n26869 , n33752 , n13477 );
    or g28758 ( n7696 , n31056 , n7632 );
    buf g28759 ( n908 , n9449 );
    or g28760 ( n34127 , n1767 , n26626 );
    or g28761 ( n20060 , n33390 , n10762 );
    nor g28762 ( n3529 , n26299 , n9921 );
    or g28763 ( n14702 , n20519 , n22931 );
    not g28764 ( n14410 , n4878 );
    xnor g28765 ( n19990 , n35879 , n30553 );
    or g28766 ( n11973 , n4276 , n4744 );
    or g28767 ( n14362 , n19502 , n22961 );
    or g28768 ( n8610 , n4307 , n27966 );
    xnor g28769 ( n26702 , n27473 , n8844 );
    or g28770 ( n8573 , n24717 , n6947 );
    or g28771 ( n17085 , n32153 , n28434 );
    xnor g28772 ( n10751 , n30888 , n14626 );
    or g28773 ( n16273 , n5123 , n19939 );
    or g28774 ( n16289 , n32838 , n8723 );
    or g28775 ( n31108 , n9474 , n21042 );
    xnor g28776 ( n22358 , n27508 , n31056 );
    or g28777 ( n26311 , n7916 , n21862 );
    or g28778 ( n21940 , n543 , n18488 );
    or g28779 ( n30830 , n35999 , n544 );
    or g28780 ( n31123 , n12306 , n27242 );
    xnor g28781 ( n11647 , n31043 , n11361 );
    xnor g28782 ( n14531 , n5801 , n17078 );
    or g28783 ( n2867 , n15450 , n34092 );
    and g28784 ( n3455 , n18175 , n15859 );
    or g28785 ( n14538 , n21240 , n11024 );
    or g28786 ( n11762 , n12721 , n20300 );
    or g28787 ( n3826 , n4510 , n9930 );
    and g28788 ( n2957 , n35647 , n12769 );
    nor g28789 ( n19802 , n5335 , n17189 );
    xnor g28790 ( n16938 , n16370 , n33936 );
    buf g28791 ( n2712 , n3396 );
    not g28792 ( n7435 , n14766 );
    or g28793 ( n6490 , n25096 , n35825 );
    or g28794 ( n26835 , n10817 , n35998 );
    nor g28795 ( n21693 , n30858 , n28866 );
    and g28796 ( n3247 , n8421 , n31240 );
    or g28797 ( n9581 , n4086 , n31564 );
    or g28798 ( n19511 , n32095 , n33164 );
    xnor g28799 ( n4762 , n4118 , n27013 );
    xnor g28800 ( n22549 , n34494 , n33957 );
    xnor g28801 ( n2471 , n21088 , n2064 );
    and g28802 ( n22531 , n17534 , n3672 );
    nor g28803 ( n10953 , n33943 , n19189 );
    or g28804 ( n31826 , n8551 , n21084 );
    not g28805 ( n29513 , n22980 );
    or g28806 ( n14650 , n8898 , n12791 );
    and g28807 ( n13861 , n26113 , n9711 );
    or g28808 ( n31432 , n13805 , n3738 );
    and g28809 ( n10553 , n16963 , n28300 );
    or g28810 ( n28803 , n30799 , n19336 );
    or g28811 ( n31512 , n4659 , n14666 );
    or g28812 ( n19495 , n4960 , n29108 );
    or g28813 ( n14104 , n32612 , n27650 );
    and g28814 ( n6703 , n5579 , n11176 );
    and g28815 ( n30790 , n22760 , n1040 );
    xnor g28816 ( n30634 , n5127 , n9789 );
    or g28817 ( n33126 , n26312 , n26737 );
    and g28818 ( n24433 , n21471 , n7908 );
    or g28819 ( n12799 , n23333 , n30292 );
    xnor g28820 ( n21245 , n16840 , n24371 );
    and g28821 ( n29570 , n310 , n17383 );
    xnor g28822 ( n22354 , n26013 , n10694 );
    or g28823 ( n3861 , n5867 , n35200 );
    or g28824 ( n30510 , n3653 , n30299 );
    not g28825 ( n14170 , n27855 );
    nor g28826 ( n15020 , n11190 , n10498 );
    or g28827 ( n7290 , n28996 , n23717 );
    or g28828 ( n9799 , n8359 , n28191 );
    and g28829 ( n28865 , n21329 , n20510 );
    or g28830 ( n4415 , n13528 , n19421 );
    nor g28831 ( n22722 , n4758 , n5280 );
    xnor g28832 ( n2576 , n20273 , n9793 );
    xnor g28833 ( n6704 , n15301 , n25610 );
    xnor g28834 ( n17866 , n19611 , n6621 );
    or g28835 ( n4737 , n23697 , n18214 );
    or g28836 ( n24141 , n26124 , n27118 );
    or g28837 ( n9957 , n18221 , n6121 );
    and g28838 ( n21 , n21576 , n25849 );
    xnor g28839 ( n10233 , n3563 , n30604 );
    or g28840 ( n34144 , n12181 , n7553 );
    or g28841 ( n10077 , n23449 , n28668 );
    not g28842 ( n4532 , n7101 );
    or g28843 ( n11118 , n26090 , n35111 );
    or g28844 ( n29494 , n28640 , n9194 );
    or g28845 ( n6811 , n7388 , n24489 );
    or g28846 ( n14833 , n33598 , n6258 );
    xnor g28847 ( n30936 , n13367 , n32702 );
    or g28848 ( n9160 , n22211 , n18811 );
    and g28849 ( n6730 , n6461 , n20306 );
    xnor g28850 ( n12732 , n101 , n23604 );
    or g28851 ( n3554 , n10523 , n10374 );
    and g28852 ( n1864 , n35039 , n4360 );
    or g28853 ( n32364 , n17703 , n14141 );
    or g28854 ( n7753 , n2216 , n17337 );
    xnor g28855 ( n22044 , n27429 , n30669 );
    and g28856 ( n19552 , n15435 , n30085 );
    or g28857 ( n29834 , n23618 , n19490 );
    or g28858 ( n30945 , n29408 , n34472 );
    or g28859 ( n34428 , n21802 , n22316 );
    or g28860 ( n19292 , n18487 , n8490 );
    or g28861 ( n5893 , n16752 , n2814 );
    or g28862 ( n15428 , n13109 , n17402 );
    or g28863 ( n18948 , n9256 , n8970 );
    xnor g28864 ( n11195 , n20406 , n2799 );
    or g28865 ( n4872 , n1477 , n34481 );
    and g28866 ( n12899 , n1804 , n6448 );
    buf g28867 ( n20558 , n9554 );
    xnor g28868 ( n30147 , n34599 , n32715 );
    xnor g28869 ( n28154 , n16164 , n23504 );
    or g28870 ( n11345 , n21875 , n7309 );
    or g28871 ( n8596 , n13979 , n24497 );
    or g28872 ( n24113 , n19551 , n23435 );
    and g28873 ( n23651 , n35525 , n20234 );
    xnor g28874 ( n18618 , n16253 , n7703 );
    xnor g28875 ( n4463 , n26259 , n328 );
    xnor g28876 ( n182 , n22272 , n27291 );
    or g28877 ( n21979 , n16742 , n26002 );
    and g28878 ( n10901 , n10631 , n1290 );
    buf g28879 ( n29626 , n17009 );
    not g28880 ( n34431 , n30586 );
    and g28881 ( n23823 , n18579 , n12075 );
    xnor g28882 ( n15051 , n28658 , n19787 );
    and g28883 ( n31461 , n24712 , n22076 );
    or g28884 ( n17567 , n30045 , n9317 );
    xnor g28885 ( n21951 , n19142 , n12702 );
    or g28886 ( n16108 , n25527 , n18644 );
    xnor g28887 ( n33108 , n31423 , n33808 );
    and g28888 ( n30704 , n4729 , n11947 );
    xnor g28889 ( n14424 , n35022 , n30206 );
    xnor g28890 ( n6055 , n24048 , n7540 );
    not g28891 ( n5346 , n22088 );
    nor g28892 ( n30861 , n23910 , n5453 );
    xnor g28893 ( n3947 , n27632 , n18174 );
    or g28894 ( n25501 , n53 , n29174 );
    or g28895 ( n23408 , n32217 , n27895 );
    xnor g28896 ( n24407 , n35411 , n32693 );
    or g28897 ( n6037 , n20338 , n2633 );
    nor g28898 ( n2781 , n811 , n1041 );
    buf g28899 ( n27574 , n19058 );
    and g28900 ( n34918 , n11951 , n21031 );
    not g28901 ( n10560 , n34563 );
    or g28902 ( n18614 , n1319 , n17162 );
    and g28903 ( n10158 , n6922 , n18155 );
    or g28904 ( n22900 , n3127 , n20840 );
    and g28905 ( n2837 , n17440 , n18812 );
    xnor g28906 ( n1328 , n13630 , n31799 );
    xnor g28907 ( n33434 , n4668 , n22291 );
    or g28908 ( n243 , n32485 , n10432 );
    or g28909 ( n13256 , n7653 , n4438 );
    xnor g28910 ( n29400 , n987 , n32095 );
    and g28911 ( n8056 , n5510 , n22785 );
    and g28912 ( n13453 , n10296 , n21821 );
    or g28913 ( n32892 , n35927 , n33154 );
    or g28914 ( n2291 , n7428 , n8098 );
    xnor g28915 ( n6648 , n32421 , n2968 );
    xnor g28916 ( n23237 , n19449 , n35314 );
    or g28917 ( n17555 , n13127 , n11593 );
    or g28918 ( n19978 , n19259 , n4254 );
    xnor g28919 ( n11521 , n10087 , n29713 );
    and g28920 ( n31255 , n31493 , n20124 );
    and g28921 ( n4630 , n29775 , n21695 );
    xnor g28922 ( n24858 , n30270 , n20175 );
    or g28923 ( n11729 , n26055 , n29626 );
    xnor g28924 ( n15860 , n2191 , n32095 );
    nor g28925 ( n34226 , n3205 , n28571 );
    and g28926 ( n35241 , n35287 , n12463 );
    or g28927 ( n8287 , n29892 , n22318 );
    and g28928 ( n33853 , n4171 , n14939 );
    or g28929 ( n26961 , n8373 , n25592 );
    or g28930 ( n26397 , n4758 , n22494 );
    xnor g28931 ( n20222 , n25074 , n15895 );
    and g28932 ( n7507 , n19773 , n18254 );
    and g28933 ( n33467 , n32122 , n30945 );
    or g28934 ( n6298 , n20878 , n21547 );
    or g28935 ( n5722 , n35724 , n28675 );
    nor g28936 ( n10725 , n28637 , n7511 );
    or g28937 ( n32212 , n16914 , n35402 );
    or g28938 ( n29128 , n10407 , n11833 );
    and g28939 ( n6711 , n14181 , n33297 );
    nor g28940 ( n5721 , n13878 , n15002 );
    xnor g28941 ( n16432 , n17041 , n21983 );
    and g28942 ( n27722 , n2464 , n21264 );
    xnor g28943 ( n26912 , n2281 , n31062 );
    or g28944 ( n28790 , n31598 , n20094 );
    xnor g28945 ( n4811 , n7752 , n18926 );
    xnor g28946 ( n10595 , n2991 , n10894 );
    or g28947 ( n20236 , n36081 , n13217 );
    or g28948 ( n33451 , n6684 , n25392 );
    and g28949 ( n25788 , n23950 , n6169 );
    nor g28950 ( n15946 , n22497 , n27720 );
    and g28951 ( n27690 , n21387 , n12452 );
    or g28952 ( n8687 , n5287 , n32518 );
    or g28953 ( n19891 , n3416 , n9930 );
    or g28954 ( n4953 , n15684 , n20817 );
    or g28955 ( n22153 , n17006 , n13053 );
    xnor g28956 ( n6168 , n917 , n22224 );
    xnor g28957 ( n14953 , n35303 , n31799 );
    or g28958 ( n34928 , n32772 , n20579 );
    or g28959 ( n30148 , n882 , n30689 );
    or g28960 ( n22833 , n16563 , n18242 );
    and g28961 ( n7410 , n17825 , n25351 );
    xnor g28962 ( n17099 , n18303 , n20844 );
    and g28963 ( n13145 , n35904 , n9784 );
    nor g28964 ( n31605 , n32715 , n34604 );
    nor g28965 ( n2801 , n28947 , n2712 );
    or g28966 ( n19344 , n5045 , n23748 );
    and g28967 ( n242 , n16658 , n23526 );
    and g28968 ( n4670 , n3912 , n19396 );
    or g28969 ( n1070 , n6699 , n17612 );
    or g28970 ( n8086 , n22643 , n20576 );
    not g28971 ( n6939 , n26716 );
    xnor g28972 ( n12341 , n13291 , n6764 );
    xnor g28973 ( n23597 , n20987 , n11046 );
    and g28974 ( n5113 , n12415 , n16559 );
    nor g28975 ( n9306 , n10894 , n7355 );
    and g28976 ( n34864 , n27064 , n20947 );
    or g28977 ( n32771 , n988 , n31627 );
    nor g28978 ( n554 , n12934 , n16690 );
    not g28979 ( n33910 , n5335 );
    or g28980 ( n22911 , n18567 , n14918 );
    xnor g28981 ( n144 , n10454 , n5112 );
    or g28982 ( n20281 , n6416 , n12791 );
    xnor g28983 ( n18965 , n30164 , n18203 );
    not g28984 ( n15368 , n34512 );
    xnor g28985 ( n32836 , n14641 , n24018 );
    or g28986 ( n30931 , n25565 , n26220 );
    or g28987 ( n4160 , n22652 , n32059 );
    and g28988 ( n16992 , n7487 , n24588 );
    or g28989 ( n27561 , n26525 , n3382 );
    and g28990 ( n21560 , n31857 , n25229 );
    or g28991 ( n9905 , n22398 , n10611 );
    buf g28992 ( n9672 , n27561 );
    or g28993 ( n126 , n28639 , n5752 );
    and g28994 ( n12026 , n31568 , n25780 );
    or g28995 ( n25582 , n32148 , n15124 );
    and g28996 ( n2136 , n20369 , n3559 );
    nor g28997 ( n6358 , n32095 , n9499 );
    or g28998 ( n20446 , n17568 , n23418 );
    xnor g28999 ( n416 , n20191 , n32095 );
    or g29000 ( n2725 , n291 , n30519 );
    and g29001 ( n2786 , n24563 , n28930 );
    and g29002 ( n7669 , n6390 , n21829 );
    xnor g29003 ( n24932 , n13861 , n31559 );
    xnor g29004 ( n25328 , n4170 , n8432 );
    or g29005 ( n20653 , n14737 , n16710 );
    and g29006 ( n4033 , n35029 , n20996 );
    or g29007 ( n6221 , n31056 , n1365 );
    or g29008 ( n26658 , n8836 , n21579 );
    or g29009 ( n29095 , n762 , n21673 );
    or g29010 ( n17581 , n8219 , n28103 );
    or g29011 ( n30135 , n8703 , n1942 );
    or g29012 ( n14087 , n7064 , n31627 );
    or g29013 ( n6497 , n14767 , n27794 );
    not g29014 ( n2592 , n4977 );
    or g29015 ( n4808 , n7587 , n22501 );
    and g29016 ( n25789 , n9486 , n9585 );
    or g29017 ( n26309 , n4878 , n30600 );
    or g29018 ( n504 , n17331 , n31514 );
    and g29019 ( n965 , n16239 , n26598 );
    not g29020 ( n5106 , n25569 );
    not g29021 ( n13744 , n34785 );
    and g29022 ( n909 , n13915 , n34876 );
    nor g29023 ( n35319 , n15886 , n19376 );
    or g29024 ( n3903 , n5650 , n10960 );
    or g29025 ( n576 , n30772 , n27501 );
    xnor g29026 ( n22252 , n18835 , n17730 );
    not g29027 ( n25477 , n33613 );
    nor g29028 ( n24749 , n19551 , n15308 );
    or g29029 ( n13090 , n616 , n11874 );
    and g29030 ( n26760 , n3933 , n6809 );
    nor g29031 ( n5777 , n27291 , n22014 );
    and g29032 ( n25347 , n1987 , n5997 );
    nor g29033 ( n3339 , n991 , n21914 );
    nor g29034 ( n33917 , n26604 , n1595 );
    nor g29035 ( n17888 , n24437 , n23921 );
    or g29036 ( n7152 , n33112 , n17125 );
    and g29037 ( n3422 , n23391 , n3929 );
    or g29038 ( n7454 , n30230 , n31705 );
    or g29039 ( n29824 , n29513 , n18536 );
    or g29040 ( n6628 , n11187 , n13915 );
    or g29041 ( n18277 , n25740 , n19173 );
    or g29042 ( n3285 , n13429 , n7448 );
    or g29043 ( n18174 , n10903 , n21462 );
    or g29044 ( n20179 , n15403 , n19019 );
    xnor g29045 ( n14103 , n15683 , n19123 );
    buf g29046 ( n7553 , n17372 );
    or g29047 ( n5656 , n3471 , n31067 );
    xnor g29048 ( n31598 , n8294 , n27291 );
    and g29049 ( n23349 , n4600 , n24303 );
    or g29050 ( n35982 , n21479 , n1969 );
    and g29051 ( n30445 , n29632 , n4441 );
    nor g29052 ( n15654 , n4960 , n21022 );
    not g29053 ( n31382 , n22980 );
    or g29054 ( n2242 , n13416 , n18723 );
    or g29055 ( n9527 , n5335 , n6437 );
    or g29056 ( n20010 , n27163 , n12194 );
    xnor g29057 ( n6774 , n13140 , n10271 );
    and g29058 ( n12320 , n25891 , n26970 );
    or g29059 ( n6217 , n27589 , n14628 );
    xnor g29060 ( n14667 , n23087 , n16606 );
    and g29061 ( n27266 , n27531 , n20715 );
    or g29062 ( n32033 , n5719 , n2524 );
    xnor g29063 ( n23363 , n22665 , n22993 );
    and g29064 ( n2221 , n26650 , n31008 );
    or g29065 ( n12216 , n17736 , n17354 );
    and g29066 ( n2363 , n1490 , n29612 );
    or g29067 ( n7501 , n32584 , n33413 );
    or g29068 ( n185 , n7057 , n31067 );
    xnor g29069 ( n24580 , n31951 , n31474 );
    and g29070 ( n27456 , n5843 , n14058 );
    xnor g29071 ( n1916 , n23431 , n30582 );
    and g29072 ( n20205 , n17069 , n13147 );
    or g29073 ( n23995 , n16822 , n26468 );
    or g29074 ( n21161 , n17370 , n5457 );
    xnor g29075 ( n1369 , n13189 , n17118 );
    nor g29076 ( n13294 , n35312 , n29819 );
    or g29077 ( n12339 , n13718 , n25786 );
    xnor g29078 ( n22309 , n9980 , n10688 );
    xnor g29079 ( n34062 , n31061 , n27776 );
    or g29080 ( n26509 , n19415 , n6288 );
    nor g29081 ( n33854 , n33928 , n15422 );
    or g29082 ( n7729 , n11186 , n21210 );
    xnor g29083 ( n25852 , n34516 , n23604 );
    nor g29084 ( n20087 , n29460 , n4555 );
    not g29085 ( n27392 , n8366 );
    or g29086 ( n15857 , n5884 , n22946 );
    or g29087 ( n30886 , n3220 , n544 );
    or g29088 ( n21643 , n31215 , n26238 );
    and g29089 ( n31053 , n22375 , n23539 );
    and g29090 ( n22050 , n11173 , n10453 );
    or g29091 ( n12943 , n7540 , n11672 );
    not g29092 ( n9979 , n11659 );
    and g29093 ( n12566 , n34920 , n17723 );
    xnor g29094 ( n1601 , n20344 , n29839 );
    or g29095 ( n5504 , n25783 , n29393 );
    xnor g29096 ( n11181 , n19499 , n26647 );
    nor g29097 ( n13201 , n23604 , n34985 );
    xnor g29098 ( n10791 , n25115 , n9793 );
    not g29099 ( n13547 , n18441 );
    or g29100 ( n3494 , n34469 , n8203 );
    not g29101 ( n9175 , n9291 );
    nor g29102 ( n17028 , n16922 , n26398 );
    and g29103 ( n26047 , n35045 , n20883 );
    xor g29104 ( n27274 , n6775 , n10162 );
    or g29105 ( n27754 , n3222 , n897 );
    and g29106 ( n24069 , n12309 , n35624 );
    and g29107 ( n4291 , n30513 , n31569 );
    xnor g29108 ( n4884 , n7568 , n22291 );
    not g29109 ( n5501 , n6257 );
    and g29110 ( n8488 , n9311 , n29789 );
    or g29111 ( n8216 , n7540 , n12867 );
    xnor g29112 ( n18424 , n2786 , n15464 );
    xnor g29113 ( n18470 , n22123 , n7540 );
    not g29114 ( n11636 , n9064 );
    or g29115 ( n27506 , n26287 , n25255 );
    xnor g29116 ( n17605 , n33207 , n10801 );
    not g29117 ( n27384 , n13179 );
    xnor g29118 ( n1191 , n12482 , n35927 );
    xnor g29119 ( n17707 , n29160 , n29839 );
    not g29120 ( n34277 , n23126 );
    xnor g29121 ( n16522 , n11085 , n16922 );
    and g29122 ( n15341 , n26936 , n32556 );
    or g29123 ( n32994 , n4668 , n35111 );
    and g29124 ( n30368 , n3154 , n15122 );
    xnor g29125 ( n27606 , n16030 , n21251 );
    nor g29126 ( n26630 , n7021 , n6424 );
    nor g29127 ( n6855 , n16620 , n2726 );
    nor g29128 ( n18523 , n35283 , n9921 );
    or g29129 ( n12924 , n2191 , n4254 );
    and g29130 ( n19272 , n14572 , n34808 );
    or g29131 ( n20422 , n10894 , n26447 );
    or g29132 ( n9128 , n18183 , n4254 );
    xnor g29133 ( n10609 , n3822 , n29839 );
    and g29134 ( n12286 , n12745 , n34090 );
    not g29135 ( n16007 , n28273 );
    nor g29136 ( n132 , n15464 , n8045 );
    or g29137 ( n22131 , n28027 , n11295 );
    and g29138 ( n33088 , n28241 , n23188 );
    or g29139 ( n16269 , n22541 , n17576 );
    nor g29140 ( n32704 , n29884 , n35227 );
    and g29141 ( n32535 , n5273 , n19221 );
    not g29142 ( n29799 , n31447 );
    and g29143 ( n20934 , n5479 , n24915 );
    or g29144 ( n7007 , n21373 , n24108 );
    and g29145 ( n4377 , n5569 , n30844 );
    or g29146 ( n9012 , n16135 , n22082 );
    not g29147 ( n35156 , n4962 );
    and g29148 ( n10861 , n27578 , n35713 );
    xnor g29149 ( n644 , n519 , n5280 );
    nor g29150 ( n21522 , n1950 , n18066 );
    or g29151 ( n4306 , n1541 , n4490 );
    not g29152 ( n100 , n12537 );
    nor g29153 ( n21039 , n28632 , n14866 );
    or g29154 ( n1666 , n4193 , n4681 );
    or g29155 ( n4051 , n27067 , n14306 );
    and g29156 ( n20096 , n4968 , n17993 );
    xnor g29157 ( n34663 , n28214 , n28407 );
    or g29158 ( n17760 , n25232 , n3756 );
    xnor g29159 ( n33182 , n18231 , n19154 );
    xnor g29160 ( n6664 , n34029 , n1950 );
    or g29161 ( n4253 , n21178 , n8924 );
    or g29162 ( n25175 , n29713 , n35004 );
    xnor g29163 ( n28819 , n17805 , n35927 );
    xnor g29164 ( n27911 , n18247 , n33848 );
    xnor g29165 ( n15468 , n17063 , n22780 );
    or g29166 ( n6167 , n6667 , n10028 );
    or g29167 ( n275 , n22291 , n11744 );
    or g29168 ( n2645 , n14166 , n30037 );
    or g29169 ( n6499 , n10159 , n31583 );
    xnor g29170 ( n16966 , n27444 , n30742 );
    not g29171 ( n12838 , n15464 );
    nor g29172 ( n30327 , n22489 , n3340 );
    xnor g29173 ( n4345 , n21778 , n25174 );
    and g29174 ( n12752 , n31943 , n20487 );
    or g29175 ( n17516 , n27644 , n15499 );
    or g29176 ( n20384 , n33702 , n26116 );
    or g29177 ( n794 , n11407 , n1146 );
    or g29178 ( n35041 , n31433 , n19421 );
    or g29179 ( n25961 , n6211 , n23323 );
    xnor g29180 ( n10655 , n20961 , n31756 );
    xnor g29181 ( n10378 , n1122 , n9789 );
    xnor g29182 ( n23107 , n24168 , n5806 );
    xnor g29183 ( n7062 , n24990 , n18725 );
    or g29184 ( n27775 , n33395 , n26132 );
    or g29185 ( n26855 , n13629 , n12996 );
    xnor g29186 ( n17319 , n8414 , n17154 );
    xnor g29187 ( n11970 , n18442 , n8221 );
    and g29188 ( n15459 , n3699 , n20645 );
    or g29189 ( n32216 , n36019 , n6459 );
    xnor g29190 ( n32230 , n7793 , n32095 );
    nor g29191 ( n36008 , n30553 , n28305 );
    or g29192 ( n7983 , n35641 , n2293 );
    and g29193 ( n24528 , n25315 , n28782 );
    xnor g29194 ( n17996 , n27577 , n34362 );
    or g29195 ( n10055 , n10088 , n1763 );
    nor g29196 ( n6789 , n4878 , n33397 );
    xnor g29197 ( n16646 , n15594 , n25802 );
    or g29198 ( n13134 , n17853 , n28455 );
    nor g29199 ( n1961 , n30589 , n27322 );
    and g29200 ( n555 , n6457 , n2904 );
    xnor g29201 ( n11056 , n7220 , n32584 );
    and g29202 ( n26581 , n34958 , n35638 );
    and g29203 ( n19277 , n28050 , n11890 );
    and g29204 ( n15005 , n35102 , n1071 );
    and g29205 ( n30114 , n31983 , n21900 );
    and g29206 ( n32388 , n13380 , n20570 );
    xnor g29207 ( n20973 , n22134 , n31075 );
    or g29208 ( n23081 , n24666 , n22240 );
    nor g29209 ( n19639 , n6347 , n19137 );
    xnor g29210 ( n8459 , n25342 , n10894 );
    or g29211 ( n8327 , n10894 , n30290 );
    xnor g29212 ( n4250 , n2676 , n5067 );
    or g29213 ( n27142 , n21234 , n22501 );
    or g29214 ( n13722 , n21630 , n26737 );
    or g29215 ( n2574 , n15373 , n20558 );
    or g29216 ( n20974 , n12673 , n11258 );
    xnor g29217 ( n2545 , n19948 , n27397 );
    or g29218 ( n16691 , n6160 , n11005 );
    or g29219 ( n6728 , n2892 , n19034 );
    or g29220 ( n28386 , n27615 , n18542 );
    or g29221 ( n6989 , n7646 , n24025 );
    or g29222 ( n34507 , n15928 , n2117 );
    or g29223 ( n16210 , n16552 , n18944 );
    xnor g29224 ( n3598 , n11790 , n26884 );
    not g29225 ( n25834 , n8366 );
    or g29226 ( n11918 , n5324 , n12538 );
    or g29227 ( n27927 , n24048 , n19464 );
    and g29228 ( n11377 , n18902 , n7675 );
    xnor g29229 ( n25199 , n30675 , n18397 );
    and g29230 ( n28417 , n17211 , n2227 );
    or g29231 ( n963 , n13802 , n4416 );
    xnor g29232 ( n26206 , n1062 , n2249 );
    xnor g29233 ( n33288 , n7091 , n33649 );
    xnor g29234 ( n26084 , n21369 , n18240 );
    or g29235 ( n18550 , n32368 , n715 );
    or g29236 ( n25357 , n12022 , n23536 );
    and g29237 ( n1783 , n35551 , n15098 );
    not g29238 ( n14734 , n252 );
    and g29239 ( n32579 , n26446 , n12379 );
    or g29240 ( n29815 , n35180 , n23349 );
    xnor g29241 ( n25913 , n10119 , n15042 );
    or g29242 ( n11721 , n19984 , n4684 );
    xnor g29243 ( n18790 , n2546 , n11046 );
    xnor g29244 ( n20755 , n20101 , n9793 );
    xnor g29245 ( n23014 , n8595 , n10177 );
    nor g29246 ( n12521 , n25602 , n18981 );
    not g29247 ( n21135 , n28009 );
    or g29248 ( n36071 , n11190 , n31960 );
    nor g29249 ( n20137 , n35927 , n28888 );
    xnor g29250 ( n10 , n7504 , n32002 );
    or g29251 ( n30187 , n3114 , n35422 );
    nor g29252 ( n34540 , n17690 , n32059 );
    or g29253 ( n28667 , n3998 , n5692 );
    or g29254 ( n35031 , n31559 , n25998 );
    and g29255 ( n33523 , n6531 , n24063 );
    xnor g29256 ( n30501 , n18372 , n8432 );
    or g29257 ( n12564 , n25917 , n14102 );
    or g29258 ( n18969 , n14120 , n3479 );
    or g29259 ( n16189 , n1950 , n4379 );
    or g29260 ( n29524 , n32950 , n437 );
    and g29261 ( n33354 , n15246 , n32762 );
    or g29262 ( n29234 , n12743 , n28574 );
    or g29263 ( n32273 , n15655 , n35422 );
    or g29264 ( n19862 , n26362 , n25340 );
    not g29265 ( n33262 , n11240 );
    or g29266 ( n12378 , n12771 , n30395 );
    and g29267 ( n24279 , n18277 , n2285 );
    or g29268 ( n6744 , n28004 , n5868 );
    or g29269 ( n26839 , n17933 , n1402 );
    or g29270 ( n24056 , n19551 , n29599 );
    xnor g29271 ( n30243 , n3813 , n29959 );
    or g29272 ( n18775 , n11846 , n13480 );
    or g29273 ( n33856 , n33317 , n3221 );
    xnor g29274 ( n27899 , n28206 , n5287 );
    or g29275 ( n3641 , n32146 , n5833 );
    nor g29276 ( n25431 , n4288 , n21680 );
    and g29277 ( n35028 , n9223 , n17138 );
    and g29278 ( n2083 , n10543 , n13159 );
    or g29279 ( n9729 , n35242 , n4363 );
    xnor g29280 ( n10564 , n3176 , n30490 );
    xnor g29281 ( n12105 , n5523 , n22291 );
    xnor g29282 ( n8060 , n5341 , n32330 );
    buf g29283 ( n16456 , n4361 );
    and g29284 ( n9673 , n6476 , n11734 );
    and g29285 ( n3386 , n18556 , n20709 );
    xnor g29286 ( n32106 , n16632 , n4962 );
    or g29287 ( n27058 , n14230 , n2005 );
    or g29288 ( n34193 , n16620 , n27100 );
    xnor g29289 ( n23106 , n15085 , n32857 );
    or g29290 ( n1366 , n1839 , n2997 );
    or g29291 ( n19130 , n21822 , n22206 );
    or g29292 ( n1746 , n31289 , n21822 );
    or g29293 ( n7182 , n760 , n22302 );
    and g29294 ( n15732 , n29260 , n8605 );
    or g29295 ( n4754 , n3222 , n6915 );
    or g29296 ( n845 , n15464 , n8771 );
    xnor g29297 ( n5657 , n32603 , n4878 );
    or g29298 ( n11366 , n31969 , n20576 );
    or g29299 ( n19792 , n9789 , n17324 );
    nor g29300 ( n10659 , n30159 , n36059 );
    not g29301 ( n15053 , n22758 );
    or g29302 ( n32184 , n9360 , n20601 );
    xnor g29303 ( n6400 , n13601 , n31799 );
    or g29304 ( n3491 , n16420 , n20849 );
    or g29305 ( n17411 , n15406 , n9482 );
    xnor g29306 ( n10517 , n15001 , n12222 );
    xnor g29307 ( n27378 , n3977 , n8524 );
    or g29308 ( n33565 , n24082 , n12950 );
    or g29309 ( n21561 , n10076 , n22322 );
    or g29310 ( n14169 , n8387 , n26931 );
    xnor g29311 ( n3470 , n20837 , n33830 );
    nor g29312 ( n31912 , n30724 , n32203 );
    or g29313 ( n31266 , n34740 , n6075 );
    or g29314 ( n16208 , n4960 , n24790 );
    or g29315 ( n12868 , n18209 , n28866 );
    xnor g29316 ( n9752 , n4352 , n22138 );
    or g29317 ( n17538 , n6317 , n8090 );
    nor g29318 ( n31318 , n1795 , n27501 );
    not g29319 ( n16525 , n26365 );
    xnor g29320 ( n13713 , n52 , n4960 );
    and g29321 ( n13618 , n20382 , n16948 );
    or g29322 ( n33465 , n17105 , n18488 );
    and g29323 ( n8474 , n26652 , n16933 );
    and g29324 ( n13642 , n24388 , n32683 );
    or g29325 ( n34995 , n25354 , n29489 );
    or g29326 ( n7080 , n3205 , n22784 );
    not g29327 ( n2912 , n22471 );
    xnor g29328 ( n13269 , n31402 , n22945 );
    or g29329 ( n25720 , n18838 , n18255 );
    or g29330 ( n34713 , n33693 , n27342 );
    or g29331 ( n33091 , n9426 , n33149 );
    xnor g29332 ( n5071 , n19376 , n15886 );
    or g29333 ( n1079 , n29078 , n9275 );
    not g29334 ( n14523 , n21989 );
    or g29335 ( n9931 , n4837 , n16326 );
    or g29336 ( n8335 , n4878 , n16065 );
    or g29337 ( n1975 , n30553 , n32067 );
    and g29338 ( n2657 , n3459 , n30641 );
    or g29339 ( n29551 , n19534 , n4702 );
    xnor g29340 ( n15119 , n18009 , n3512 );
    xnor g29341 ( n20247 , n16527 , n20352 );
    or g29342 ( n27435 , n22114 , n19928 );
    not g29343 ( n13826 , n14259 );
    or g29344 ( n24536 , n3445 , n2168 );
    or g29345 ( n22517 , n7580 , n16598 );
    and g29346 ( n33001 , n3948 , n9390 );
    not g29347 ( n30756 , n14995 );
    or g29348 ( n27088 , n5746 , n20303 );
    or g29349 ( n5785 , n30742 , n28451 );
    and g29350 ( n25318 , n21016 , n28366 );
    not g29351 ( n6909 , n8432 );
    or g29352 ( n28619 , n22168 , n11258 );
    xnor g29353 ( n12643 , n4711 , n11455 );
    xnor g29354 ( n29422 , n3715 , n27291 );
    or g29355 ( n31706 , n6912 , n22316 );
    or g29356 ( n28061 , n30742 , n32350 );
    or g29357 ( n31031 , n13168 , n26184 );
    xnor g29358 ( n13447 , n27448 , n22940 );
    or g29359 ( n35091 , n11223 , n5168 );
    or g29360 ( n6673 , n21269 , n1041 );
    and g29361 ( n21782 , n33453 , n31852 );
    or g29362 ( n16312 , n15886 , n32110 );
    xnor g29363 ( n27332 , n26732 , n27124 );
    or g29364 ( n28580 , n34778 , n23642 );
    and g29365 ( n23828 , n9797 , n16091 );
    xnor g29366 ( n6681 , n9355 , n5287 );
    xnor g29367 ( n30512 , n14755 , n22004 );
    and g29368 ( n24412 , n19684 , n21289 );
    xnor g29369 ( n302 , n26428 , n5738 );
    not g29370 ( n17430 , n20480 );
    or g29371 ( n27350 , n23634 , n24837 );
    xnor g29372 ( n12012 , n9397 , n921 );
    or g29373 ( n5148 , n3485 , n6459 );
    and g29374 ( n12590 , n12635 , n28409 );
    or g29375 ( n22004 , n35084 , n32443 );
    or g29376 ( n19799 , n20161 , n20733 );
    nor g29377 ( n19078 , n27226 , n14281 );
    or g29378 ( n16104 , n11959 , n17162 );
    xnor g29379 ( n26822 , n10041 , n23266 );
    or g29380 ( n30346 , n18886 , n13035 );
    and g29381 ( n24628 , n32034 , n12192 );
    not g29382 ( n11543 , n31913 );
    xnor g29383 ( n4839 , n20565 , n28559 );
    or g29384 ( n1823 , n16350 , n15439 );
    xnor g29385 ( n15313 , n4072 , n10894 );
    and g29386 ( n34822 , n31903 , n24073 );
    xnor g29387 ( n3720 , n30960 , n35927 );
    or g29388 ( n15990 , n16620 , n4263 );
    or g29389 ( n149 , n1900 , n16543 );
    or g29390 ( n7846 , n580 , n11593 );
    xnor g29391 ( n12406 , n30814 , n20341 );
    not g29392 ( n29045 , n16223 );
    and g29393 ( n32913 , n15593 , n35902 );
    xnor g29394 ( n30536 , n13274 , n18878 );
    xnor g29395 ( n21424 , n29444 , n830 );
    not g29396 ( n1769 , n27732 );
    buf g29397 ( n23090 , n21398 );
    or g29398 ( n6987 , n13896 , n25550 );
    or g29399 ( n15036 , n25963 , n19314 );
    or g29400 ( n6169 , n21762 , n16345 );
    and g29401 ( n15834 , n5330 , n14914 );
    or g29402 ( n28008 , n19860 , n25392 );
    or g29403 ( n28481 , n18946 , n13305 );
    or g29404 ( n15433 , n8406 , n2005 );
    or g29405 ( n24325 , n5580 , n8392 );
    and g29406 ( n12515 , n4362 , n5418 );
    or g29407 ( n19823 , n31720 , n30057 );
    or g29408 ( n33881 , n9891 , n7598 );
    or g29409 ( n15035 , n11455 , n32 );
    xnor g29410 ( n15976 , n10640 , n3911 );
    nor g29411 ( n31230 , n17702 , n26769 );
    or g29412 ( n7445 , n10601 , n908 );
    or g29413 ( n27753 , n25662 , n35056 );
    or g29414 ( n17777 , n20946 , n3842 );
    not g29415 ( n28898 , n21075 );
    or g29416 ( n12484 , n29367 , n30708 );
    nor g29417 ( n17781 , n34558 , n17087 );
    or g29418 ( n31304 , n24371 , n409 );
    or g29419 ( n3558 , n19469 , n18477 );
    or g29420 ( n16074 , n14566 , n2104 );
    xnor g29421 ( n10429 , n14496 , n4965 );
    or g29422 ( n35210 , n1436 , n13015 );
    or g29423 ( n28090 , n22291 , n28938 );
    or g29424 ( n1390 , n31799 , n4113 );
    or g29425 ( n6483 , n14643 , n6459 );
    not g29426 ( n22422 , n18712 );
    or g29427 ( n33048 , n29839 , n24346 );
    and g29428 ( n19079 , n24145 , n13249 );
    or g29429 ( n9759 , n8487 , n27053 );
    buf g29430 ( n6257 , n18721 );
    or g29431 ( n25576 , n24337 , n21977 );
    nor g29432 ( n11968 , n11046 , n31531 );
    or g29433 ( n622 , n31799 , n35931 );
    or g29434 ( n20674 , n24371 , n11156 );
    and g29435 ( n11042 , n22910 , n1531 );
    or g29436 ( n17627 , n17759 , n1402 );
    nor g29437 ( n12450 , n12264 , n28787 );
    or g29438 ( n27233 , n11190 , n2176 );
    xnor g29439 ( n19518 , n30386 , n11455 );
    or g29440 ( n27247 , n8137 , n24696 );
    or g29441 ( n8664 , n14594 , n27580 );
    or g29442 ( n848 , n32263 , n1374 );
    and g29443 ( n27663 , n25083 , n4887 );
    xnor g29444 ( n10162 , n10076 , n4878 );
    or g29445 ( n27977 , n23049 , n31549 );
    and g29446 ( n27453 , n16183 , n16492 );
    or g29447 ( n12555 , n29631 , n12332 );
    or g29448 ( n25830 , n33740 , n16382 );
    or g29449 ( n8310 , n11894 , n12188 );
    or g29450 ( n936 , n31056 , n29552 );
    and g29451 ( n7163 , n10376 , n7331 );
    or g29452 ( n34890 , n11193 , n16259 );
    xnor g29453 ( n36051 , n27568 , n22616 );
    xnor g29454 ( n9323 , n5522 , n12288 );
    xnor g29455 ( n33459 , n32158 , n17862 );
    or g29456 ( n2937 , n19996 , n11258 );
    or g29457 ( n3827 , n10640 , n3911 );
    xnor g29458 ( n33010 , n24334 , n32468 );
    and g29459 ( n23328 , n30137 , n16857 );
    and g29460 ( n23045 , n22919 , n22671 );
    xnor g29461 ( n14807 , n20171 , n24093 );
    xnor g29462 ( n22409 , n1903 , n4962 );
    or g29463 ( n779 , n31215 , n16924 );
    or g29464 ( n8568 , n30485 , n31606 );
    or g29465 ( n28375 , n32535 , n8723 );
    xnor g29466 ( n23654 , n29208 , n22291 );
    and g29467 ( n8595 , n7034 , n7052 );
    or g29468 ( n60 , n17247 , n15805 );
    or g29469 ( n805 , n31155 , n24895 );
    or g29470 ( n30075 , n1447 , n29266 );
    or g29471 ( n18340 , n25174 , n9501 );
    nor g29472 ( n24310 , n30636 , n35472 );
    or g29473 ( n4312 , n26879 , n21862 );
    or g29474 ( n10059 , n30736 , n20601 );
    not g29475 ( n33673 , n27502 );
    or g29476 ( n12078 , n6847 , n15542 );
    or g29477 ( n29022 , n10894 , n33109 );
    xnor g29478 ( n22335 , n20977 , n8432 );
    xor g29479 ( n8895 , n2156 , n31958 );
    or g29480 ( n29809 , n11965 , n11996 );
    and g29481 ( n26924 , n12719 , n6889 );
    not g29482 ( n27892 , n1299 );
    not g29483 ( n32378 , n14653 );
    or g29484 ( n8939 , n8932 , n24333 );
    and g29485 ( n13767 , n6718 , n8971 );
    and g29486 ( n2556 , n1190 , n551 );
    xnor g29487 ( n11151 , n4880 , n4878 );
    xnor g29488 ( n33681 , n4995 , n19984 );
    or g29489 ( n6723 , n26908 , n240 );
    xnor g29490 ( n29792 , n9141 , n446 );
    and g29491 ( n15456 , n32245 , n6197 );
    and g29492 ( n30852 , n5946 , n26602 );
    and g29493 ( n25661 , n9719 , n8747 );
    xnor g29494 ( n3123 , n13338 , n34254 );
    or g29495 ( n10006 , n7921 , n24025 );
    or g29496 ( n3905 , n16004 , n14399 );
    or g29497 ( n31670 , n30888 , n14626 );
    and g29498 ( n17483 , n4126 , n8581 );
    or g29499 ( n25956 , n22645 , n27016 );
    or g29500 ( n18014 , n23604 , n2300 );
    xnor g29501 ( n3854 , n25878 , n8432 );
    nor g29502 ( n18810 , n1679 , n5387 );
    or g29503 ( n28075 , n14293 , n30519 );
    or g29504 ( n15229 , n25537 , n32572 );
    not g29505 ( n13222 , n17396 );
    xnor g29506 ( n31787 , n5182 , n3280 );
    xnor g29507 ( n12599 , n12968 , n4962 );
    not g29508 ( n24192 , n4960 );
    or g29509 ( n29335 , n911 , n8201 );
    or g29510 ( n30133 , n25220 , n18737 );
    and g29511 ( n9703 , n34389 , n15988 );
    nor g29512 ( n34735 , n8597 , n30242 );
    and g29513 ( n9668 , n33955 , n434 );
    or g29514 ( n2095 , n10346 , n33107 );
    or g29515 ( n30329 , n27584 , n34971 );
    or g29516 ( n21566 , n24768 , n3673 );
    or g29517 ( n22640 , n1612 , n30893 );
    and g29518 ( n32362 , n24123 , n25554 );
    xnor g29519 ( n16741 , n22843 , n5067 );
    or g29520 ( n26981 , n24404 , n18811 );
    xnor g29521 ( n24080 , n16672 , n18007 );
    and g29522 ( n8372 , n1607 , n16372 );
    and g29523 ( n9357 , n24683 , n11362 );
    or g29524 ( n30787 , n20155 , n24489 );
    not g29525 ( n22955 , n32558 );
    xnor g29526 ( n32277 , n6449 , n16191 );
    or g29527 ( n13004 , n25174 , n30704 );
    or g29528 ( n13313 , n22808 , n26008 );
    xnor g29529 ( n19650 , n14934 , n27659 );
    not g29530 ( n20341 , n9793 );
    not g29531 ( n13737 , n8266 );
    xnor g29532 ( n31913 , n16857 , n29276 );
    or g29533 ( n27286 , n27008 , n20318 );
    xnor g29534 ( n16742 , n1003 , n28252 );
    and g29535 ( n6913 , n1781 , n31254 );
    or g29536 ( n12060 , n27022 , n18264 );
    and g29537 ( n8438 , n21103 , n12421 );
    or g29538 ( n22566 , n17919 , n32738 );
    or g29539 ( n7622 , n31508 , n4337 );
    xnor g29540 ( n24731 , n25589 , n27294 );
    or g29541 ( n9224 , n8535 , n25314 );
    and g29542 ( n11039 , n5517 , n25016 );
    or g29543 ( n12430 , n11742 , n1474 );
    or g29544 ( n17865 , n7398 , n18268 );
    and g29545 ( n19044 , n14664 , n9771 );
    or g29546 ( n27922 , n411 , n4952 );
    or g29547 ( n34774 , n23688 , n20840 );
    or g29548 ( n12898 , n15659 , n1171 );
    xnor g29549 ( n14344 , n7666 , n22291 );
    or g29550 ( n4517 , n34269 , n21018 );
    and g29551 ( n12381 , n29110 , n13381 );
    or g29552 ( n3531 , n34356 , n21956 );
    xnor g29553 ( n14665 , n7380 , n31272 );
    or g29554 ( n31418 , n5614 , n27728 );
    not g29555 ( n16633 , n5019 );
    and g29556 ( n16582 , n30676 , n4259 );
    not g29557 ( n19649 , n828 );
    and g29558 ( n13250 , n14499 , n29982 );
    or g29559 ( n11443 , n8432 , n17562 );
    not g29560 ( n16894 , n1111 );
    xnor g29561 ( n25121 , n29161 , n21164 );
    nor g29562 ( n23586 , n31799 , n25645 );
    and g29563 ( n33605 , n17808 , n3971 );
    xnor g29564 ( n2562 , n30709 , n5701 );
    xnor g29565 ( n31070 , n14673 , n10787 );
    or g29566 ( n33028 , n12493 , n15344 );
    or g29567 ( n3269 , n19984 , n32725 );
    and g29568 ( n10737 , n28179 , n34630 );
    and g29569 ( n19584 , n6955 , n22199 );
    nor g29570 ( n17662 , n16857 , n3472 );
    and g29571 ( n5421 , n5159 , n19282 );
    and g29572 ( n14571 , n24487 , n32216 );
    xnor g29573 ( n13751 , n7623 , n33277 );
    xnor g29574 ( n35434 , n15450 , n34092 );
    nor g29575 ( n11403 , n5287 , n35292 );
    buf g29576 ( n20579 , n4367 );
    or g29577 ( n22872 , n16984 , n30826 );
    or g29578 ( n19943 , n26046 , n30708 );
    and g29579 ( n21142 , n13895 , n2407 );
    or g29580 ( n23061 , n18040 , n27276 );
    or g29581 ( n2007 , n34737 , n34537 );
    or g29582 ( n15566 , n26286 , n11601 );
    xnor g29583 ( n25474 , n33354 , n31799 );
    or g29584 ( n31636 , n20726 , n25594 );
    and g29585 ( n23015 , n25449 , n3260 );
    and g29586 ( n22264 , n7866 , n32902 );
    or g29587 ( n5043 , n16522 , n16729 );
    and g29588 ( n27443 , n3075 , n22167 );
    or g29589 ( n10711 , n14801 , n30013 );
    xnor g29590 ( n4487 , n17054 , n5200 );
    nor g29591 ( n29346 , n26498 , n9555 );
    xnor g29592 ( n32265 , n34517 , n31643 );
    not g29593 ( n7340 , n9905 );
    or g29594 ( n2052 , n30742 , n14350 );
    or g29595 ( n21170 , n25570 , n28668 );
    and g29596 ( n20268 , n10035 , n7541 );
    xnor g29597 ( n10222 , n8148 , n24120 );
    or g29598 ( n33691 , n3187 , n12560 );
    or g29599 ( n14016 , n19551 , n35746 );
    and g29600 ( n35586 , n10834 , n26565 );
    xnor g29601 ( n24598 , n19112 , n31696 );
    or g29602 ( n31360 , n3364 , n17354 );
    nor g29603 ( n27304 , n28574 , n30734 );
    xnor g29604 ( n7227 , n10227 , n35420 );
    and g29605 ( n17862 , n11602 , n9542 );
    or g29606 ( n15026 , n25292 , n32329 );
    and g29607 ( n29999 , n27798 , n642 );
    or g29608 ( n10047 , n14400 , n4478 );
    and g29609 ( n7708 , n30424 , n28951 );
    xnor g29610 ( n29184 , n12527 , n2537 );
    and g29611 ( n34075 , n4846 , n17937 );
    nor g29612 ( n14055 , n35883 , n4024 );
    or g29613 ( n18030 , n7785 , n2471 );
    nor g29614 ( n19808 , n8432 , n549 );
    xnor g29615 ( n18054 , n15017 , n9513 );
    nor g29616 ( n27905 , n835 , n12178 );
    and g29617 ( n6371 , n13596 , n32373 );
    not g29618 ( n18554 , n4288 );
    xnor g29619 ( n16986 , n21114 , n21616 );
    or g29620 ( n18060 , n17568 , n19038 );
    or g29621 ( n34019 , n13638 , n8412 );
    and g29622 ( n28351 , n28146 , n17176 );
    not g29623 ( n16502 , n11079 );
    and g29624 ( n27353 , n769 , n8947 );
    nor g29625 ( n11576 , n32095 , n18700 );
    and g29626 ( n15090 , n29806 , n32231 );
    or g29627 ( n16908 , n24744 , n26112 );
    and g29628 ( n11958 , n17706 , n10852 );
    xnor g29629 ( n1655 , n419 , n32095 );
    xnor g29630 ( n14230 , n16923 , n24843 );
    not g29631 ( n10923 , n11653 );
    not g29632 ( n32434 , n11712 );
    and g29633 ( n33112 , n30171 , n33239 );
    or g29634 ( n956 , n22416 , n13470 );
    or g29635 ( n32406 , n27896 , n35663 );
    not g29636 ( n26653 , n35938 );
    or g29637 ( n27668 , n10818 , n34971 );
    and g29638 ( n4937 , n14483 , n29027 );
    or g29639 ( n5524 , n32617 , n26002 );
    not g29640 ( n21641 , n18830 );
    and g29641 ( n4014 , n14713 , n412 );
    xnor g29642 ( n31694 , n7930 , n3338 );
    or g29643 ( n16036 , n17751 , n14605 );
    or g29644 ( n19706 , n31378 , n28248 );
    xnor g29645 ( n19723 , n29960 , n2828 );
    not g29646 ( n10669 , n13744 );
    or g29647 ( n13417 , n17532 , n949 );
    or g29648 ( n35430 , n11922 , n33416 );
    not g29649 ( n19702 , n33387 );
    or g29650 ( n13038 , n12911 , n33007 );
    or g29651 ( n11420 , n236 , n8476 );
    and g29652 ( n26001 , n20028 , n29325 );
    and g29653 ( n15507 , n6985 , n26079 );
    and g29654 ( n23572 , n33292 , n23055 );
    nor g29655 ( n2972 , n33514 , n7166 );
    not g29656 ( n1307 , n19194 );
    not g29657 ( n14274 , n29104 );
    xnor g29658 ( n8604 , n32394 , n13888 );
    nor g29659 ( n18038 , n15886 , n17194 );
    and g29660 ( n15678 , n33636 , n4516 );
    or g29661 ( n4027 , n21638 , n9601 );
    xnor g29662 ( n14767 , n24953 , n17568 );
    or g29663 ( n35195 , n27504 , n19952 );
    and g29664 ( n2091 , n31430 , n24096 );
    and g29665 ( n19810 , n36076 , n4415 );
    or g29666 ( n18696 , n32482 , n31055 );
    buf g29667 ( n5618 , n15967 );
    not g29668 ( n35840 , n5019 );
    or g29669 ( n34925 , n23632 , n32071 );
    or g29670 ( n8501 , n25438 , n12671 );
    xnor g29671 ( n30964 , n25008 , n31786 );
    or g29672 ( n19035 , n4288 , n28808 );
    and g29673 ( n31048 , n19329 , n21912 );
    and g29674 ( n3815 , n24903 , n18014 );
    and g29675 ( n28472 , n20290 , n16823 );
    xnor g29676 ( n4734 , n16924 , n31215 );
    and g29677 ( n8186 , n11868 , n19032 );
    or g29678 ( n24446 , n26733 , n17612 );
    or g29679 ( n29680 , n29981 , n31514 );
    or g29680 ( n22152 , n11455 , n20727 );
    or g29681 ( n5918 , n9942 , n16464 );
    xnor g29682 ( n24806 , n3376 , n18970 );
    or g29683 ( n25310 , n32857 , n30146 );
    and g29684 ( n16771 , n10106 , n14426 );
    not g29685 ( n20343 , n29732 );
    and g29686 ( n33892 , n31934 , n18352 );
    not g29687 ( n22464 , n22176 );
    or g29688 ( n31102 , n4758 , n16069 );
    or g29689 ( n29654 , n9446 , n17829 );
    and g29690 ( n3448 , n24658 , n19769 );
    xnor g29691 ( n18361 , n34969 , n1435 );
    or g29692 ( n17210 , n29908 , n22241 );
    or g29693 ( n26777 , n2753 , n28788 );
    nor g29694 ( n27317 , n14402 , n9921 );
    nor g29695 ( n3609 , n31559 , n4536 );
    xnor g29696 ( n12104 , n30961 , n18002 );
    or g29697 ( n2861 , n34018 , n21525 );
    xnor g29698 ( n9535 , n4630 , n18283 );
    or g29699 ( n5871 , n3747 , n16961 );
    xnor g29700 ( n17315 , n33274 , n33805 );
    and g29701 ( n34404 , n9462 , n29419 );
    and g29702 ( n17543 , n31764 , n34108 );
    not g29703 ( n13663 , n8767 );
    or g29704 ( n9496 , n29705 , n32853 );
    nor g29705 ( n11418 , n23328 , n16414 );
    not g29706 ( n26670 , n18555 );
    nor g29707 ( n12546 , n23453 , n7271 );
    xnor g29708 ( n25269 , n13565 , n5287 );
    xnor g29709 ( n17240 , n19280 , n35355 );
    or g29710 ( n13481 , n31559 , n31203 );
    xnor g29711 ( n9697 , n23098 , n29296 );
    and g29712 ( n25783 , n22584 , n25393 );
    nor g29713 ( n27544 , n9789 , n5488 );
    nor g29714 ( n13303 , n32857 , n6480 );
    or g29715 ( n9375 , n23508 , n35475 );
    nor g29716 ( n16084 , n29713 , n23722 );
    not g29717 ( n7151 , n28866 );
    xnor g29718 ( n3021 , n9357 , n16922 );
    or g29719 ( n36067 , n22947 , n26659 );
    or g29720 ( n4506 , n4104 , n1989 );
    or g29721 ( n23526 , n16722 , n29411 );
    or g29722 ( n21264 , n29888 , n28248 );
    nor g29723 ( n10690 , n11135 , n28974 );
    nor g29724 ( n23175 , n9515 , n29258 );
    xnor g29725 ( n21806 , n15503 , n35927 );
    or g29726 ( n35843 , n11254 , n4595 );
    or g29727 ( n20600 , n16954 , n32913 );
    nor g29728 ( n35969 , n33842 , n10962 );
    and g29729 ( n23163 , n8520 , n35284 );
    or g29730 ( n21858 , n4288 , n24744 );
    or g29731 ( n145 , n1055 , n24505 );
    and g29732 ( n14654 , n28216 , n6963 );
    or g29733 ( n31911 , n30679 , n475 );
    or g29734 ( n17432 , n16922 , n16075 );
    and g29735 ( n17794 , n24233 , n16121 );
    or g29736 ( n33350 , n34294 , n578 );
    and g29737 ( n16926 , n12522 , n24823 );
    not g29738 ( n8805 , n4960 );
    or g29739 ( n13621 , n11559 , n24696 );
    or g29740 ( n10880 , n11046 , n33633 );
    xnor g29741 ( n730 , n26574 , n5778 );
    and g29742 ( n26939 , n8733 , n26139 );
    or g29743 ( n34474 , n31269 , n16806 );
    and g29744 ( n17673 , n12005 , n29968 );
    xnor g29745 ( n33169 , n7637 , n9793 );
    xnor g29746 ( n15231 , n25118 , n30297 );
    or g29747 ( n34893 , n33376 , n13480 );
    and g29748 ( n23603 , n1933 , n8540 );
    and g29749 ( n5343 , n7431 , n11180 );
    nor g29750 ( n16965 , n805 , n33157 );
    or g29751 ( n14312 , n4960 , n505 );
    xnor g29752 ( n18094 , n23221 , n2082 );
    or g29753 ( n5105 , n30425 , n20308 );
    and g29754 ( n2129 , n3142 , n2190 );
    and g29755 ( n8975 , n1637 , n12854 );
    not g29756 ( n13051 , n9658 );
    and g29757 ( n18598 , n31042 , n26764 );
    xnor g29758 ( n8712 , n14662 , n32857 );
    nor g29759 ( n14272 , n25486 , n19025 );
    and g29760 ( n15503 , n23672 , n21915 );
    or g29761 ( n27338 , n24619 , n5618 );
    xnor g29762 ( n9052 , n10441 , n6002 );
    xnor g29763 ( n34054 , n20368 , n830 );
    or g29764 ( n5518 , n12736 , n5618 );
    nor g29765 ( n13012 , n20949 , n32526 );
    or g29766 ( n23837 , n16081 , n16553 );
    or g29767 ( n6068 , n36020 , n35196 );
    and g29768 ( n31072 , n15857 , n1308 );
    or g29769 ( n29958 , n31559 , n14179 );
    or g29770 ( n2809 , n11455 , n771 );
    nor g29771 ( n2341 , n35927 , n35649 );
    or g29772 ( n35893 , n3222 , n17027 );
    not g29773 ( n35475 , n33435 );
    not g29774 ( n19743 , n14756 );
    not g29775 ( n9440 , n20840 );
    or g29776 ( n31767 , n10894 , n33411 );
    or g29777 ( n18777 , n30796 , n7553 );
    nor g29778 ( n29741 , n24371 , n24985 );
    and g29779 ( n24121 , n10919 , n9977 );
    or g29780 ( n30172 , n8586 , n20308 );
    or g29781 ( n7924 , n1950 , n30772 );
    not g29782 ( n27665 , n2926 );
    xnor g29783 ( n30332 , n28358 , n14232 );
    and g29784 ( n6569 , n31130 , n4828 );
    xnor g29785 ( n9667 , n3002 , n32584 );
    xnor g29786 ( n8808 , n30695 , n29249 );
    or g29787 ( n29223 , n3205 , n12044 );
    nor g29788 ( n33915 , n15296 , n118 );
    and g29789 ( n8703 , n24917 , n16766 );
    or g29790 ( n31221 , n35344 , n5277 );
    buf g29791 ( n21691 , n3477 );
    and g29792 ( n17730 , n23505 , n14750 );
    not g29793 ( n4608 , n29137 );
    not g29794 ( n28648 , n19939 );
    and g29795 ( n18238 , n30639 , n10827 );
    xnor g29796 ( n8798 , n4407 , n21017 );
    xnor g29797 ( n3229 , n10855 , n9658 );
    nor g29798 ( n35762 , n14944 , n6414 );
    or g29799 ( n34190 , n22030 , n25255 );
    xnor g29800 ( n33777 , n33197 , n34909 );
    xnor g29801 ( n9201 , n31881 , n16571 );
    or g29802 ( n5401 , n10311 , n949 );
    or g29803 ( n4152 , n26242 , n25392 );
    nor g29804 ( n2522 , n34209 , n20148 );
    nor g29805 ( n23136 , n9793 , n25116 );
    or g29806 ( n2848 , n30212 , n17301 );
    xnor g29807 ( n13372 , n5719 , n31289 );
    or g29808 ( n15703 , n9789 , n26748 );
    or g29809 ( n28267 , n9359 , n4428 );
    or g29810 ( n6126 , n32921 , n32703 );
    or g29811 ( n25671 , n7188 , n20603 );
    or g29812 ( n33180 , n3205 , n36081 );
    or g29813 ( n29282 , n19833 , n16809 );
    xnor g29814 ( n14412 , n4131 , n25602 );
    and g29815 ( n35327 , n23162 , n12293 );
    and g29816 ( n32814 , n35423 , n22980 );
    or g29817 ( n26057 , n24749 , n20314 );
    buf g29818 ( n2955 , n2287 );
    or g29819 ( n7040 , n33132 , n35402 );
    xnor g29820 ( n8911 , n14150 , n8827 );
    or g29821 ( n8336 , n17271 , n6050 );
    not g29822 ( n15033 , n6075 );
    or g29823 ( n17449 , n7235 , n34973 );
    and g29824 ( n33674 , n31009 , n28464 );
    and g29825 ( n8317 , n36067 , n5025 );
    or g29826 ( n5143 , n32220 , n28574 );
    xnor g29827 ( n14649 , n24117 , n7982 );
    xnor g29828 ( n29304 , n30737 , n4878 );
    and g29829 ( n34150 , n30321 , n9130 );
    or g29830 ( n15171 , n31289 , n4710 );
    and g29831 ( n29077 , n23712 , n36058 );
    and g29832 ( n2548 , n22439 , n23326 );
    xnor g29833 ( n1033 , n17422 , n27226 );
    and g29834 ( n16711 , n26749 , n26603 );
    not g29835 ( n31233 , n18925 );
    nor g29836 ( n18924 , n16620 , n13027 );
    or g29837 ( n31860 , n4982 , n10872 );
    and g29838 ( n14137 , n19665 , n27861 );
    or g29839 ( n16279 , n704 , n2572 );
    or g29840 ( n26738 , n32584 , n12925 );
    xnor g29841 ( n21788 , n15399 , n27268 );
    and g29842 ( n3762 , n11299 , n13233 );
    or g29843 ( n165 , n34667 , n27437 );
    or g29844 ( n14074 , n32857 , n10504 );
    and g29845 ( n14950 , n22269 , n35254 );
    or g29846 ( n27302 , n29713 , n26090 );
    or g29847 ( n34177 , n10894 , n28822 );
    and g29848 ( n34234 , n13081 , n735 );
    and g29849 ( n25463 , n20607 , n33699 );
    not g29850 ( n33919 , n35407 );
    xnor g29851 ( n21942 , n13864 , n30194 );
    or g29852 ( n33509 , n29397 , n34484 );
    not g29853 ( n27186 , n3205 );
    not g29854 ( n14390 , n9496 );
    or g29855 ( n24659 , n29800 , n17233 );
    or g29856 ( n769 , n7832 , n585 );
    xnor g29857 ( n23470 , n846 , n5150 );
    or g29858 ( n27154 , n32077 , n2080 );
    xnor g29859 ( n27198 , n20708 , n13810 );
    buf g29860 ( n12465 , n21382 );
    or g29861 ( n19596 , n28568 , n1904 );
    or g29862 ( n3582 , n19447 , n22316 );
    not g29863 ( n841 , n35927 );
    xnor g29864 ( n5065 , n26049 , n3205 );
    and g29865 ( n34989 , n34474 , n19516 );
    or g29866 ( n19769 , n20101 , n35935 );
    xnor g29867 ( n24974 , n4951 , n31815 );
    not g29868 ( n1901 , n32721 );
    and g29869 ( n4422 , n31522 , n10996 );
    or g29870 ( n26140 , n34763 , n9317 );
    not g29871 ( n32412 , n17004 );
    and g29872 ( n3345 , n22928 , n3322 );
    nor g29873 ( n32120 , n32095 , n26529 );
    or g29874 ( n9007 , n10887 , n23748 );
    and g29875 ( n31750 , n32835 , n23158 );
    or g29876 ( n24480 , n29280 , n33956 );
    nor g29877 ( n31435 , n32363 , n14274 );
    nor g29878 ( n13712 , n27226 , n27815 );
    or g29879 ( n33264 , n33838 , n8465 );
    and g29880 ( n32073 , n5984 , n15077 );
    and g29881 ( n12466 , n13588 , n10231 );
    and g29882 ( n33254 , n2945 , n12427 );
    or g29883 ( n21009 , n7540 , n26146 );
    nor g29884 ( n19793 , n17109 , n1219 );
    xnor g29885 ( n10957 , n6100 , n4645 );
    or g29886 ( n18885 , n31799 , n21521 );
    or g29887 ( n20407 , n8028 , n30195 );
    or g29888 ( n22 , n17751 , n19341 );
    or g29889 ( n28310 , n9150 , n16216 );
    or g29890 ( n13576 , n3306 , n1010 );
    or g29891 ( n16418 , n22291 , n7568 );
    or g29892 ( n14051 , n10299 , n27962 );
    xnor g29893 ( n2525 , n25854 , n31487 );
    or g29894 ( n8747 , n17751 , n27259 );
    and g29895 ( n33229 , n29548 , n20889 );
    and g29896 ( n35791 , n6952 , n5846 );
    xnor g29897 ( n35753 , n25026 , n31215 );
    nor g29898 ( n29413 , n15886 , n33668 );
    or g29899 ( n16982 , n26825 , n26319 );
    or g29900 ( n20883 , n4901 , n1715 );
    nor g29901 ( n9054 , n4878 , n15079 );
    or g29902 ( n7687 , n1566 , n5972 );
    not g29903 ( n31225 , n5985 );
    and g29904 ( n6880 , n21526 , n10451 );
    not g29905 ( n32662 , n24434 );
    and g29906 ( n21653 , n2 , n8177 );
    and g29907 ( n35478 , n35370 , n34974 );
    not g29908 ( n28186 , n9789 );
    or g29909 ( n31281 , n19271 , n15538 );
    or g29910 ( n15672 , n30226 , n35141 );
    and g29911 ( n20964 , n35082 , n6213 );
    xnor g29912 ( n27430 , n16740 , n10181 );
    and g29913 ( n13492 , n14219 , n2616 );
    xnor g29914 ( n14741 , n10655 , n33987 );
    or g29915 ( n22969 , n17351 , n9478 );
    xnor g29916 ( n19570 , n6124 , n4758 );
    xnor g29917 ( n13296 , n33670 , n33302 );
    and g29918 ( n18357 , n35873 , n24206 );
    and g29919 ( n24713 , n21776 , n8113 );
    or g29920 ( n2924 , n13047 , n7553 );
    or g29921 ( n4235 , n28299 , n33177 );
    or g29922 ( n1400 , n3540 , n27574 );
    xnor g29923 ( n11318 , n8244 , n32095 );
    or g29924 ( n35016 , n18323 , n26806 );
    or g29925 ( n20990 , n5696 , n9930 );
    or g29926 ( n19411 , n31799 , n33354 );
    xnor g29927 ( n35886 , n6834 , n35146 );
    and g29928 ( n33205 , n25833 , n9535 );
    and g29929 ( n13933 , n6865 , n9408 );
    xnor g29930 ( n8470 , n29248 , n3222 );
    or g29931 ( n32291 , n2620 , n18654 );
    xnor g29932 ( n717 , n1377 , n25174 );
    not g29933 ( n20921 , n27685 );
    and g29934 ( n8752 , n7153 , n11542 );
    xnor g29935 ( n1965 , n7795 , n27786 );
    or g29936 ( n1213 , n11455 , n8965 );
    or g29937 ( n23641 , n8317 , n18936 );
    xnor g29938 ( n19828 , n31765 , n10894 );
    or g29939 ( n20975 , n23604 , n13548 );
    nor g29940 ( n22485 , n14320 , n32689 );
    and g29941 ( n15234 , n19096 , n32993 );
    nor g29942 ( n17845 , n23268 , n9480 );
    nor g29943 ( n23182 , n9789 , n8323 );
    or g29944 ( n16559 , n10894 , n35605 );
    and g29945 ( n9604 , n6152 , n19849 );
    or g29946 ( n23226 , n17471 , n15109 );
    xnor g29947 ( n9791 , n24457 , n11190 );
    xnor g29948 ( n8800 , n29561 , n26856 );
    xnor g29949 ( n664 , n11585 , n1499 );
    or g29950 ( n4483 , n4938 , n11312 );
    or g29951 ( n13699 , n2164 , n11039 );
    or g29952 ( n23376 , n15874 , n15256 );
    or g29953 ( n33273 , n31702 , n11593 );
    or g29954 ( n32145 , n18426 , n35618 );
    or g29955 ( n6691 , n11606 , n35078 );
    or g29956 ( n32979 , n11758 , n1734 );
    or g29957 ( n27640 , n25602 , n26773 );
    or g29958 ( n23767 , n32684 , n5459 );
    or g29959 ( n13353 , n7325 , n30445 );
    xnor g29960 ( n15182 , n31413 , n21189 );
    xnor g29961 ( n997 , n3900 , n14759 );
    or g29962 ( n20290 , n24372 , n25594 );
    and g29963 ( n3611 , n5246 , n33352 );
    and g29964 ( n4598 , n28677 , n29155 );
    or g29965 ( n28294 , n5335 , n30809 );
    xnor g29966 ( n1618 , n15469 , n12377 );
    or g29967 ( n22365 , n35259 , n18255 );
    or g29968 ( n15922 , n4916 , n24333 );
    or g29969 ( n11836 , n19551 , n20683 );
    not g29970 ( n3754 , n2029 );
    or g29971 ( n30681 , n21082 , n7914 );
    and g29972 ( n12100 , n22636 , n35675 );
    not g29973 ( n30056 , n33206 );
    not g29974 ( n30507 , n16326 );
    or g29975 ( n3715 , n9197 , n15610 );
    xnor g29976 ( n7432 , n30054 , n5335 );
    and g29977 ( n14533 , n15852 , n2919 );
    not g29978 ( n22101 , n30141 );
    and g29979 ( n10437 , n23982 , n5032 );
    or g29980 ( n2871 , n29326 , n27185 );
    xnor g29981 ( n19871 , n32770 , n22194 );
    xnor g29982 ( n3670 , n6851 , n2067 );
    and g29983 ( n33551 , n6142 , n17841 );
    xnor g29984 ( n8219 , n22693 , n5335 );
    or g29985 ( n21727 , n5623 , n31773 );
    xnor g29986 ( n34580 , n5092 , n24051 );
    or g29987 ( n6740 , n10528 , n10432 );
    and g29988 ( n4249 , n29636 , n27347 );
    or g29989 ( n10223 , n34096 , n23625 );
    or g29990 ( n24706 , n5977 , n29132 );
    xnor g29991 ( n536 , n9490 , n22105 );
    xnor g29992 ( n10091 , n30715 , n4288 );
    xnor g29993 ( n3003 , n13940 , n4878 );
    not g29994 ( n7274 , n10322 );
    or g29995 ( n13471 , n31649 , n32959 );
    or g29996 ( n12359 , n18027 , n27437 );
    or g29997 ( n11691 , n11671 , n11833 );
    xnor g29998 ( n28254 , n14364 , n32680 );
    xnor g29999 ( n7191 , n22799 , n34749 );
    and g30000 ( n3527 , n22120 , n12696 );
    xnor g30001 ( n3217 , n25376 , n581 );
    or g30002 ( n18254 , n8384 , n5208 );
    or g30003 ( n11146 , n30742 , n27169 );
    or g30004 ( n32427 , n3321 , n27558 );
    xnor g30005 ( n26224 , n293 , n25728 );
    and g30006 ( n1744 , n20365 , n24041 );
    or g30007 ( n13604 , n14899 , n12596 );
    xnor g30008 ( n27239 , n7479 , n15872 );
    or g30009 ( n12804 , n17578 , n28696 );
    or g30010 ( n7491 , n24371 , n22569 );
    and g30011 ( n7272 , n13984 , n30480 );
    and g30012 ( n20629 , n9748 , n3286 );
    or g30013 ( n25493 , n26757 , n25761 );
    or g30014 ( n2990 , n30286 , n5779 );
    or g30015 ( n11302 , n18862 , n30204 );
    nor g30016 ( n2561 , n32857 , n10601 );
    and g30017 ( n35204 , n17362 , n21609 );
    or g30018 ( n25901 , n9370 , n30732 );
    xnor g30019 ( n15807 , n24339 , n3205 );
    or g30020 ( n18019 , n1662 , n5116 );
    xnor g30021 ( n34496 , n8606 , n10067 );
    xnor g30022 ( n27723 , n2128 , n12764 );
    or g30023 ( n20005 , n28532 , n20576 );
    or g30024 ( n15776 , n14495 , n12663 );
    nor g30025 ( n5013 , n14826 , n9921 );
    or g30026 ( n13200 , n15886 , n12840 );
    or g30027 ( n25091 , n4758 , n29967 );
    not g30028 ( n26884 , n16620 );
    xnor g30029 ( n5655 , n9132 , n32958 );
    and g30030 ( n31953 , n23897 , n18616 );
    xnor g30031 ( n7957 , n8417 , n20922 );
    xnor g30032 ( n32571 , n8623 , n15707 );
    or g30033 ( n31427 , n4492 , n24345 );
    or g30034 ( n29814 , n11614 , n2832 );
    and g30035 ( n33615 , n5201 , n22709 );
    and g30036 ( n27309 , n24743 , n17059 );
    and g30037 ( n27962 , n4565 , n34243 );
    or g30038 ( n11795 , n29324 , n29643 );
    xnor g30039 ( n15923 , n20541 , n15464 );
    and g30040 ( n10425 , n35463 , n11917 );
    not g30041 ( n31734 , n9106 );
    xnor g30042 ( n26709 , n11870 , n3517 );
    xnor g30043 ( n30046 , n30003 , n35868 );
    or g30044 ( n34393 , n29713 , n21598 );
    and g30045 ( n12591 , n9767 , n26039 );
    xnor g30046 ( n13268 , n25435 , n31215 );
    or g30047 ( n27427 , n18956 , n34431 );
    and g30048 ( n8416 , n8333 , n1853 );
    or g30049 ( n21469 , n30289 , n2590 );
    not g30050 ( n24869 , n2092 );
    or g30051 ( n5571 , n23851 , n22757 );
    not g30052 ( n23337 , n34731 );
    or g30053 ( n32140 , n31932 , n33364 );
    or g30054 ( n26993 , n29490 , n25154 );
    or g30055 ( n24832 , n19963 , n30826 );
    buf g30056 ( n26192 , n22794 );
    or g30057 ( n10606 , n12820 , n4939 );
    or g30058 ( n22378 , n4726 , n8090 );
    or g30059 ( n34797 , n3222 , n24766 );
    not g30060 ( n33658 , n35682 );
    xnor g30061 ( n28175 , n18402 , n35927 );
    or g30062 ( n35905 , n20164 , n3756 );
    or g30063 ( n25971 , n19824 , n30804 );
    xnor g30064 ( n13109 , n28490 , n19551 );
    not g30065 ( n20439 , n17568 );
    xnor g30066 ( n34352 , n19256 , n27488 );
    not g30067 ( n22753 , n6288 );
    not g30068 ( n4657 , n22200 );
    xnor g30069 ( n3924 , n32417 , n9164 );
    or g30070 ( n23146 , n19551 , n30066 );
    not g30071 ( n22007 , n13715 );
    and g30072 ( n31451 , n16500 , n6290 );
    or g30073 ( n23928 , n21242 , n33581 );
    and g30074 ( n6756 , n18428 , n35469 );
    xnor g30075 ( n199 , n23914 , n8495 );
    or g30076 ( n13236 , n32497 , n33335 );
    or g30077 ( n2928 , n28958 , n19086 );
    xnor g30078 ( n6834 , n5949 , n1592 );
    or g30079 ( n8483 , n4088 , n2108 );
    or g30080 ( n31977 , n23953 , n28123 );
    xnor g30081 ( n12890 , n17923 , n27218 );
    or g30082 ( n22608 , n33825 , n19732 );
    nor g30083 ( n34782 , n7387 , n24259 );
    or g30084 ( n26593 , n24343 , n25594 );
    nor g30085 ( n24621 , n18379 , n10933 );
    and g30086 ( n33116 , n17330 , n2962 );
    or g30087 ( n34392 , n13623 , n23698 );
    xnor g30088 ( n20242 , n15341 , n3205 );
    or g30089 ( n14992 , n19413 , n15256 );
    nor g30090 ( n2819 , n23604 , n25606 );
    and g30091 ( n7990 , n32155 , n21476 );
    or g30092 ( n33349 , n13225 , n25019 );
    or g30093 ( n1724 , n31737 , n16456 );
    or g30094 ( n31234 , n31832 , n25773 );
    or g30095 ( n19481 , n6581 , n33471 );
    and g30096 ( n25411 , n3919 , n32374 );
    not g30097 ( n35190 , n27858 );
    xnor g30098 ( n31422 , n30034 , n9793 );
    xnor g30099 ( n28920 , n29010 , n10894 );
    and g30100 ( n19994 , n32339 , n18641 );
    xnor g30101 ( n383 , n11159 , n10894 );
    or g30102 ( n27140 , n23690 , n3805 );
    or g30103 ( n25556 , n22291 , n16168 );
    or g30104 ( n1333 , n18762 , n12465 );
    or g30105 ( n18085 , n5791 , n15256 );
    nor g30106 ( n26264 , n4267 , n29867 );
    nor g30107 ( n12767 , n3205 , n14029 );
    and g30108 ( n27929 , n11375 , n30030 );
    xnor g30109 ( n7284 , n10734 , n31068 );
    or g30110 ( n7920 , n28517 , n23819 );
    and g30111 ( n31832 , n34880 , n22049 );
    or g30112 ( n24571 , n12171 , n9731 );
    or g30113 ( n14314 , n23791 , n18348 );
    and g30114 ( n29368 , n17516 , n5764 );
    xnor g30115 ( n35614 , n196 , n9793 );
    or g30116 ( n31810 , n17856 , n8090 );
    not g30117 ( n25402 , n10894 );
    xnor g30118 ( n2264 , n17546 , n18122 );
    xnor g30119 ( n10017 , n25207 , n19455 );
    and g30120 ( n20084 , n15252 , n12906 );
    not g30121 ( n26782 , n9789 );
    or g30122 ( n20986 , n14489 , n4490 );
    or g30123 ( n11588 , n19028 , n25786 );
    and g30124 ( n11223 , n31995 , n34105 );
    and g30125 ( n30139 , n26544 , n9487 );
    xnor g30126 ( n10948 , n31492 , n25174 );
    or g30127 ( n19522 , n16135 , n1867 );
    or g30128 ( n29627 , n13667 , n15497 );
    and g30129 ( n35303 , n31537 , n3866 );
    or g30130 ( n4851 , n3622 , n35585 );
    nor g30131 ( n33731 , n16620 , n19881 );
    and g30132 ( n8824 , n20996 , n16620 );
    xnor g30133 ( n16584 , n11859 , n28989 );
    or g30134 ( n19270 , n35869 , n3298 );
    xnor g30135 ( n9351 , n13299 , n5287 );
    nor g30136 ( n21021 , n4878 , n7944 );
    or g30137 ( n1107 , n19907 , n18488 );
    or g30138 ( n32687 , n35467 , n22241 );
    or g30139 ( n33726 , n27151 , n32329 );
    or g30140 ( n26148 , n25954 , n8857 );
    or g30141 ( n318 , n33470 , n13785 );
    and g30142 ( n10484 , n32865 , n9830 );
    or g30143 ( n23053 , n12342 , n30287 );
    or g30144 ( n33293 , n6866 , n27284 );
    or g30145 ( n6836 , n922 , n6818 );
    and g30146 ( n34552 , n33437 , n21904 );
    and g30147 ( n7572 , n27321 , n295 );
    xnor g30148 ( n27513 , n15669 , n8432 );
    or g30149 ( n18016 , n3176 , n30490 );
    and g30150 ( n35923 , n220 , n29093 );
    or g30151 ( n31470 , n9793 , n13791 );
    not g30152 ( n24441 , n32574 );
    or g30153 ( n4350 , n5578 , n6940 );
    and g30154 ( n33018 , n21746 , n16578 );
    and g30155 ( n22396 , n34419 , n18679 );
    or g30156 ( n22314 , n20825 , n22732 );
    xnor g30157 ( n23195 , n2346 , n32537 );
    nor g30158 ( n31497 , n35048 , n33157 );
    and g30159 ( n2802 , n534 , n21669 );
    nor g30160 ( n35593 , n19850 , n22720 );
    xnor g30161 ( n27777 , n421 , n32857 );
    or g30162 ( n17632 , n4960 , n32224 );
    or g30163 ( n20802 , n17634 , n34891 );
    or g30164 ( n4730 , n32095 , n3931 );
    or g30165 ( n9839 , n21090 , n7553 );
    or g30166 ( n3982 , n28676 , n23090 );
    or g30167 ( n10018 , n18076 , n26919 );
    nor g30168 ( n31962 , n6160 , n25567 );
    xnor g30169 ( n31195 , n25375 , n16620 );
    or g30170 ( n12773 , n23312 , n35748 );
    nor g30171 ( n28558 , n24371 , n22334 );
    or g30172 ( n11122 , n4288 , n25448 );
    or g30173 ( n20970 , n23658 , n128 );
    not g30174 ( n4450 , n12622 );
    and g30175 ( n24873 , n7518 , n9138 );
    and g30176 ( n5490 , n35373 , n10705 );
    and g30177 ( n20500 , n34007 , n11842 );
    or g30178 ( n19598 , n24766 , n30365 );
    xnor g30179 ( n34264 , n30293 , n21819 );
    xnor g30180 ( n11991 , n9261 , n19091 );
    nor g30181 ( n31265 , n17568 , n30774 );
    not g30182 ( n14850 , n10828 );
    and g30183 ( n3362 , n29292 , n12518 );
    or g30184 ( n31876 , n3803 , n10336 );
    and g30185 ( n27253 , n14372 , n14569 );
    xnor g30186 ( n8417 , n4510 , n24371 );
    or g30187 ( n13809 , n4962 , n9238 );
    or g30188 ( n1186 , n31559 , n20490 );
    or g30189 ( n29193 , n6917 , n28859 );
    not g30190 ( n2237 , n16108 );
    not g30191 ( n16045 , n2568 );
    xnor g30192 ( n29342 , n31199 , n19514 );
    and g30193 ( n31960 , n31834 , n6084 );
    and g30194 ( n2338 , n11681 , n9586 );
    or g30195 ( n22694 , n6648 , n27580 );
    nor g30196 ( n33163 , n10057 , n1252 );
    nor g30197 ( n7500 , n18798 , n8134 );
    or g30198 ( n8066 , n1360 , n26613 );
    and g30199 ( n4695 , n30712 , n34950 );
    or g30200 ( n30002 , n9193 , n28574 );
    or g30201 ( n4692 , n31799 , n35303 );
    or g30202 ( n18485 , n18053 , n31549 );
    not g30203 ( n27178 , n24488 );
    or g30204 ( n23303 , n22291 , n30852 );
    not g30205 ( n32043 , n25602 );
    not g30206 ( n2211 , n20558 );
    or g30207 ( n34140 , n196 , n15919 );
    xnor g30208 ( n24290 , n20065 , n15444 );
    not g30209 ( n25381 , n4878 );
    or g30210 ( n31709 , n29311 , n20797 );
    xnor g30211 ( n7328 , n32585 , n11673 );
    or g30212 ( n8622 , n18379 , n33373 );
    xnor g30213 ( n8205 , n21165 , n26589 );
    xnor g30214 ( n30192 , n1365 , n31056 );
    xnor g30215 ( n13513 , n26680 , n1950 );
    and g30216 ( n30050 , n27676 , n6999 );
    and g30217 ( n34236 , n25142 , n20965 );
    not g30218 ( n2030 , n254 );
    xnor g30219 ( n32218 , n25460 , n9113 );
    and g30220 ( n33407 , n33314 , n27205 );
    and g30221 ( n2575 , n522 , n29779 );
    or g30222 ( n19595 , n4935 , n28873 );
    and g30223 ( n32972 , n16969 , n13128 );
    and g30224 ( n10557 , n24925 , n8659 );
    or g30225 ( n21809 , n3591 , n2168 );
    or g30226 ( n16287 , n32088 , n17829 );
    xnor g30227 ( n15979 , n15047 , n9658 );
    or g30228 ( n30509 , n330 , n34472 );
    and g30229 ( n29842 , n8144 , n8935 );
    or g30230 ( n10824 , n9978 , n12622 );
    xnor g30231 ( n28119 , n22531 , n31799 );
    not g30232 ( n1679 , n22980 );
    or g30233 ( n4575 , n11106 , n23871 );
    or g30234 ( n27684 , n1950 , n5566 );
    or g30235 ( n5938 , n30718 , n30419 );
    xnor g30236 ( n31478 , n11233 , n4878 );
    or g30237 ( n30051 , n9789 , n17729 );
    not g30238 ( n6442 , n2716 );
    and g30239 ( n3626 , n3230 , n16405 );
    or g30240 ( n18922 , n8313 , n3437 );
    or g30241 ( n27942 , n24332 , n16261 );
    xnor g30242 ( n6506 , n9064 , n10355 );
    and g30243 ( n7464 , n7562 , n12061 );
    and g30244 ( n9025 , n24201 , n21958 );
    and g30245 ( n25307 , n3133 , n11006 );
    or g30246 ( n27007 , n10510 , n15009 );
    or g30247 ( n35942 , n3785 , n32969 );
    and g30248 ( n14697 , n30551 , n12214 );
    nor g30249 ( n11871 , n34561 , n6806 );
    or g30250 ( n431 , n4469 , n34727 );
    and g30251 ( n2531 , n34605 , n24078 );
    xnor g30252 ( n8816 , n5961 , n27291 );
    or g30253 ( n26963 , n24371 , n3138 );
    and g30254 ( n5905 , n13856 , n9452 );
    or g30255 ( n14843 , n25373 , n30646 );
    xnor g30256 ( n27503 , n32493 , n25174 );
    or g30257 ( n1733 , n35411 , n32693 );
    and g30258 ( n30415 , n4412 , n3153 );
    or g30259 ( n17503 , n18289 , n6553 );
    and g30260 ( n18301 , n14087 , n22714 );
    and g30261 ( n23740 , n1194 , n25680 );
    or g30262 ( n35679 , n20232 , n6288 );
    not g30263 ( n34503 , n26261 );
    or g30264 ( n24469 , n35193 , n5208 );
    not g30265 ( n4214 , n5485 );
    and g30266 ( n10694 , n20802 , n24257 );
    nor g30267 ( n28200 , n15688 , n35538 );
    and g30268 ( n19550 , n6105 , n1834 );
    xnor g30269 ( n2512 , n9100 , n12020 );
    or g30270 ( n18788 , n30773 , n21037 );
    or g30271 ( n18594 , n5393 , n10386 );
    or g30272 ( n3857 , n5335 , n512 );
    xnor g30273 ( n27843 , n18837 , n8879 );
    xnor g30274 ( n10710 , n17972 , n28291 );
    or g30275 ( n17486 , n28642 , n13307 );
    nor g30276 ( n24895 , n30256 , n1419 );
    nor g30277 ( n25674 , n19551 , n8514 );
    or g30278 ( n8329 , n31799 , n6606 );
    nor g30279 ( n171 , n28249 , n31020 );
    or g30280 ( n31039 , n12245 , n32730 );
    or g30281 ( n31652 , n15886 , n13567 );
    or g30282 ( n15939 , n32857 , n34742 );
    or g30283 ( n28937 , n26156 , n19143 );
    and g30284 ( n34894 , n484 , n4589 );
    nor g30285 ( n23628 , n1950 , n18018 );
    xnor g30286 ( n30661 , n28374 , n19430 );
    xnor g30287 ( n7238 , n29639 , n3600 );
    nor g30288 ( n16580 , n17751 , n18204 );
    or g30289 ( n4949 , n699 , n3437 );
    and g30290 ( n36081 , n232 , n24126 );
    nor g30291 ( n19700 , n33925 , n1470 );
    and g30292 ( n12803 , n18627 , n10838 );
    or g30293 ( n33252 , n25612 , n25786 );
    xnor g30294 ( n8821 , n16206 , n15507 );
    and g30295 ( n24277 , n31028 , n12632 );
    xnor g30296 ( n27441 , n29165 , n2219 );
    or g30297 ( n12623 , n11478 , n24259 );
    or g30298 ( n33054 , n11268 , n18488 );
    or g30299 ( n32269 , n32752 , n3979 );
    and g30300 ( n26626 , n26399 , n1771 );
    or g30301 ( n24101 , n15574 , n28355 );
    or g30302 ( n18806 , n32584 , n33101 );
    nor g30303 ( n27808 , n25602 , n18562 );
    xnor g30304 ( n25079 , n20846 , n24371 );
    and g30305 ( n7270 , n35413 , n15306 );
    or g30306 ( n13460 , n21106 , n34472 );
    and g30307 ( n25419 , n34028 , n30000 );
    or g30308 ( n28116 , n17249 , n33275 );
    or g30309 ( n6863 , n9605 , n4772 );
    nor g30310 ( n23425 , n13639 , n25983 );
    not g30311 ( n33172 , n4874 );
    xnor g30312 ( n6412 , n22409 , n1934 );
    xnor g30313 ( n16923 , n4642 , n10115 );
    nor g30314 ( n28364 , n29400 , n4297 );
    or g30315 ( n31293 , n20107 , n2823 );
    or g30316 ( n26936 , n31985 , n11850 );
    and g30317 ( n3911 , n22532 , n7131 );
    or g30318 ( n18455 , n5275 , n30708 );
    and g30319 ( n2608 , n8321 , n452 );
    and g30320 ( n26794 , n4910 , n34513 );
    or g30321 ( n21373 , n10892 , n33661 );
    and g30322 ( n27815 , n27140 , n620 );
    or g30323 ( n28269 , n3766 , n25940 );
    and g30324 ( n20328 , n31938 , n7948 );
    xnor g30325 ( n259 , n25512 , n8283 );
    or g30326 ( n18805 , n1950 , n1340 );
    or g30327 ( n17534 , n14330 , n12596 );
    xnor g30328 ( n30777 , n32449 , n15403 );
    and g30329 ( n5249 , n9239 , n15448 );
    or g30330 ( n2475 , n25116 , n25831 );
    or g30331 ( n18530 , n32266 , n27574 );
    and g30332 ( n12968 , n3621 , n12608 );
    not g30333 ( n2085 , n31799 );
    or g30334 ( n26445 , n13497 , n18850 );
    and g30335 ( n7302 , n4393 , n3354 );
    and g30336 ( n1745 , n35006 , n32867 );
    or g30337 ( n29204 , n33604 , n13015 );
    nor g30338 ( n18291 , n3251 , n25370 );
    and g30339 ( n34599 , n31278 , n35991 );
    or g30340 ( n34642 , n16620 , n25357 );
    xnor g30341 ( n19534 , n18039 , n25602 );
    xnor g30342 ( n10054 , n33918 , n23604 );
    or g30343 ( n23320 , n12591 , n29376 );
    and g30344 ( n20529 , n21911 , n31642 );
    or g30345 ( n34498 , n17506 , n35630 );
    and g30346 ( n26883 , n16371 , n4652 );
    xnor g30347 ( n11152 , n4120 , n25602 );
    xnor g30348 ( n4881 , n7041 , n15303 );
    or g30349 ( n4420 , n27318 , n35891 );
    and g30350 ( n15393 , n19119 , n33660 );
    not g30351 ( n24581 , n9361 );
    or g30352 ( n29740 , n34846 , n16451 );
    or g30353 ( n661 , n18317 , n34600 );
    or g30354 ( n26080 , n11455 , n24035 );
    nor g30355 ( n23178 , n35927 , n17805 );
    nor g30356 ( n32581 , n13051 , n11596 );
    or g30357 ( n20080 , n5657 , n2651 );
    not g30358 ( n29730 , n17751 );
    or g30359 ( n26384 , n27646 , n27963 );
    buf g30360 ( n19403 , n2310 );
    or g30361 ( n20348 , n14300 , n7644 );
    and g30362 ( n20337 , n28267 , n34654 );
    or g30363 ( n4221 , n1399 , n29489 );
    nor g30364 ( n21268 , n29122 , n2996 );
    xnor g30365 ( n836 , n10653 , n4791 );
    not g30366 ( n27895 , n9361 );
    or g30367 ( n5159 , n5855 , n29592 );
    xnor g30368 ( n9552 , n3747 , n23604 );
    or g30369 ( n28482 , n21693 , n14777 );
    or g30370 ( n25538 , n31807 , n2253 );
    or g30371 ( n13852 , n14591 , n10960 );
    or g30372 ( n28629 , n3745 , n14748 );
    xnor g30373 ( n32670 , n26408 , n3167 );
    and g30374 ( n13300 , n7389 , n14007 );
    or g30375 ( n8485 , n22210 , n13307 );
    and g30376 ( n7670 , n11767 , n4521 );
    xnor g30377 ( n13163 , n12696 , n12487 );
    nor g30378 ( n16903 , n3570 , n28655 );
    or g30379 ( n17952 , n14467 , n11708 );
    not g30380 ( n11287 , n29921 );
    or g30381 ( n5776 , n27226 , n9852 );
    or g30382 ( n10232 , n17284 , n12596 );
    and g30383 ( n25116 , n34190 , n36050 );
    not g30384 ( n2812 , n8691 );
    xnor g30385 ( n15567 , n6322 , n9448 );
    and g30386 ( n21026 , n6642 , n7592 );
    xnor g30387 ( n30494 , n29983 , n26782 );
    and g30388 ( n1500 , n2228 , n31174 );
    or g30389 ( n28841 , n2429 , n5868 );
    or g30390 ( n32240 , n13389 , n9696 );
    or g30391 ( n20361 , n11808 , n34537 );
    xnor g30392 ( n17981 , n20556 , n22788 );
    and g30393 ( n417 , n11887 , n15706 );
    and g30394 ( n32449 , n3289 , n35621 );
    and g30395 ( n13344 , n17201 , n22759 );
    or g30396 ( n26925 , n25602 , n31949 );
    or g30397 ( n31645 , n26327 , n15145 );
    not g30398 ( n930 , n19727 );
    or g30399 ( n31646 , n35782 , n27437 );
    or g30400 ( n11545 , n29796 , n17337 );
    xnor g30401 ( n23373 , n4080 , n28159 );
    and g30402 ( n28647 , n27934 , n11694 );
    nor g30403 ( n35199 , n1950 , n22173 );
    not g30404 ( n3243 , n5784 );
    and g30405 ( n29519 , n10365 , n34715 );
    or g30406 ( n8837 , n7217 , n16919 );
    or g30407 ( n32706 , n31167 , n12879 );
    xnor g30408 ( n27515 , n17321 , n12296 );
    xnor g30409 ( n11885 , n31087 , n3940 );
    nor g30410 ( n30829 , n10389 , n33956 );
    or g30411 ( n14046 , n18923 , n17354 );
    or g30412 ( n21975 , n7540 , n12433 );
    xnor g30413 ( n6571 , n17033 , n16385 );
    or g30414 ( n33340 , n29265 , n21248 );
    not g30415 ( n13021 , n29839 );
    or g30416 ( n21387 , n8380 , n32329 );
    or g30417 ( n7362 , n23196 , n25392 );
    not g30418 ( n7348 , n31799 );
    xnor g30419 ( n22074 , n4262 , n17050 );
    and g30420 ( n30255 , n16774 , n29076 );
    or g30421 ( n3545 , n17485 , n25533 );
    and g30422 ( n34022 , n22917 , n10137 );
    and g30423 ( n25384 , n21101 , n24718 );
    xnor g30424 ( n15634 , n14073 , n20959 );
    or g30425 ( n13360 , n29839 , n32972 );
    or g30426 ( n28284 , n28990 , n20690 );
    and g30427 ( n11844 , n33867 , n626 );
    xnor g30428 ( n17394 , n33480 , n6166 );
    or g30429 ( n5496 , n15403 , n14101 );
    xnor g30430 ( n30557 , n21532 , n9789 );
    xnor g30431 ( n33047 , n764 , n27232 );
    and g30432 ( n742 , n14457 , n32999 );
    or g30433 ( n3044 , n4517 , n17068 );
    or g30434 ( n14972 , n27226 , n20887 );
    or g30435 ( n19640 , n1369 , n15344 );
    or g30436 ( n25529 , n33704 , n25789 );
    or g30437 ( n3120 , n20474 , n15144 );
    or g30438 ( n6312 , n34333 , n31627 );
    xnor g30439 ( n14241 , n651 , n4338 );
    xnor g30440 ( n3571 , n2169 , n12219 );
    not g30441 ( n16553 , n10455 );
    xnor g30442 ( n1958 , n5693 , n6068 );
    xnor g30443 ( n30061 , n5152 , n11046 );
    xnor g30444 ( n16391 , n12306 , n27242 );
    xnor g30445 ( n31258 , n8241 , n19984 );
    or g30446 ( n16268 , n27815 , n4844 );
    or g30447 ( n2517 , n11051 , n34862 );
    or g30448 ( n34125 , n29360 , n20576 );
    or g30449 ( n13185 , n16494 , n21042 );
    and g30450 ( n4570 , n29252 , n25461 );
    and g30451 ( n27552 , n7614 , n16786 );
    or g30452 ( n14875 , n1099 , n22737 );
    nor g30453 ( n34421 , n419 , n33956 );
    or g30454 ( n24010 , n33009 , n16676 );
    or g30455 ( n35592 , n24648 , n20300 );
    or g30456 ( n7545 , n4960 , n15752 );
    or g30457 ( n9912 , n11575 , n908 );
    buf g30458 ( n1511 , n3858 );
    and g30459 ( n28184 , n34570 , n1887 );
    not g30460 ( n22655 , n9039 );
    or g30461 ( n34630 , n27734 , n30431 );
    or g30462 ( n13072 , n9615 , n27443 );
    or g30463 ( n5302 , n8351 , n6442 );
    xnor g30464 ( n13831 , n18824 , n17357 );
    or g30465 ( n7946 , n31289 , n35579 );
    and g30466 ( n18183 , n8492 , n29753 );
    or g30467 ( n19329 , n8459 , n22102 );
    and g30468 ( n22377 , n25103 , n28671 );
    or g30469 ( n14926 , n8993 , n13204 );
    or g30470 ( n28552 , n26235 , n14218 );
    or g30471 ( n19253 , n27279 , n25761 );
    or g30472 ( n19701 , n2089 , n12973 );
    or g30473 ( n31018 , n12526 , n260 );
    and g30474 ( n2167 , n25501 , n22196 );
    not g30475 ( n25849 , n31559 );
    and g30476 ( n21251 , n15334 , n8536 );
    xnor g30477 ( n29981 , n11334 , n27171 );
    or g30478 ( n33912 , n4878 , n10529 );
    or g30479 ( n7933 , n4013 , n2814 );
    and g30480 ( n10537 , n29740 , n15171 );
    and g30481 ( n22649 , n32554 , n1775 );
    xnor g30482 ( n24796 , n20090 , n3928 );
    xnor g30483 ( n22327 , n15930 , n12057 );
    and g30484 ( n8587 , n9739 , n7323 );
    xnor g30485 ( n12488 , n7573 , n17483 );
    not g30486 ( n20350 , n22597 );
    buf g30487 ( n4508 , n6017 );
    or g30488 ( n5015 , n6804 , n4189 );
    nor g30489 ( n32764 , n24371 , n32520 );
    xnor g30490 ( n749 , n28693 , n32857 );
    or g30491 ( n13468 , n5730 , n6736 );
    or g30492 ( n4990 , n9897 , n10526 );
    not g30493 ( n33916 , n15918 );
    or g30494 ( n19868 , n15299 , n27885 );
    xnor g30495 ( n1843 , n15641 , n24651 );
    and g30496 ( n23115 , n4704 , n2507 );
    or g30497 ( n10732 , n21590 , n12499 );
    and g30498 ( n1293 , n6485 , n17830 );
    xnor g30499 ( n821 , n28965 , n28728 );
    and g30500 ( n34844 , n31256 , n29235 );
    or g30501 ( n24803 , n28736 , n16797 );
    or g30502 ( n28326 , n17751 , n18437 );
    or g30503 ( n34024 , n14683 , n17162 );
    or g30504 ( n28452 , n15631 , n21210 );
    xnor g30505 ( n24885 , n27098 , n5146 );
    nor g30506 ( n2975 , n9789 , n4204 );
    and g30507 ( n15896 , n979 , n11766 );
    or g30508 ( n20103 , n23 , n14824 );
    xnor g30509 ( n12150 , n7209 , n15464 );
    or g30510 ( n35399 , n4038 , n2798 );
    buf g30511 ( n15805 , n20140 );
    and g30512 ( n29963 , n16540 , n35003 );
    or g30513 ( n14004 , n1362 , n16456 );
    and g30514 ( n8564 , n24557 , n15591 );
    and g30515 ( n9033 , n27469 , n11130 );
    xnor g30516 ( n22383 , n13042 , n15221 );
    xnor g30517 ( n30523 , n22942 , n31559 );
    or g30518 ( n18133 , n4962 , n23466 );
    buf g30519 ( n3694 , n30406 );
    and g30520 ( n33389 , n2337 , n10851 );
    xnor g30521 ( n34166 , n12574 , n9033 );
    and g30522 ( n25219 , n29240 , n34895 );
    or g30523 ( n26042 , n11046 , n1436 );
    or g30524 ( n36083 , n16620 , n13226 );
    and g30525 ( n7388 , n1216 , n25286 );
    or g30526 ( n5510 , n30591 , n1511 );
    xnor g30527 ( n14995 , n23080 , n12652 );
    and g30528 ( n23594 , n26427 , n32895 );
    or g30529 ( n19795 , n31272 , n5423 );
    nor g30530 ( n35105 , n16922 , n19546 );
    and g30531 ( n17285 , n16278 , n15199 );
    xnor g30532 ( n1478 , n16314 , n11046 );
    or g30533 ( n1450 , n7751 , n20300 );
    and g30534 ( n32442 , n2012 , n13999 );
    and g30535 ( n6537 , n23527 , n3580 );
    or g30536 ( n27737 , n24136 , n31823 );
    nor g30537 ( n11163 , n20615 , n19617 );
    or g30538 ( n17443 , n3833 , n10752 );
    or g30539 ( n23058 , n29713 , n29531 );
    xnor g30540 ( n360 , n22163 , n20440 );
    and g30541 ( n11459 , n35872 , n4692 );
    or g30542 ( n29845 , n25606 , n26112 );
    or g30543 ( n5434 , n5683 , n8523 );
    or g30544 ( n2940 , n35719 , n35748 );
    xnor g30545 ( n14121 , n5899 , n20692 );
    or g30546 ( n6280 , n27037 , n24653 );
    nor g30547 ( n8688 , n25602 , n14619 );
    or g30548 ( n7490 , n2608 , n22946 );
    and g30549 ( n33889 , n8727 , n32833 );
    or g30550 ( n10130 , n11455 , n13863 );
    xnor g30551 ( n7880 , n878 , n31272 );
    not g30552 ( n27604 , n3475 );
    and g30553 ( n22737 , n30346 , n1729 );
    or g30554 ( n29695 , n17458 , n35748 );
    or g30555 ( n22355 , n14065 , n12465 );
    or g30556 ( n34629 , n28421 , n25019 );
    and g30557 ( n9205 , n33560 , n3903 );
    and g30558 ( n9657 , n27303 , n537 );
    not g30559 ( n21353 , n3675 );
    xnor g30560 ( n2596 , n10465 , n21342 );
    xnor g30561 ( n27036 , n26556 , n32095 );
    xnor g30562 ( n26784 , n5259 , n21712 );
    and g30563 ( n138 , n15933 , n22484 );
    or g30564 ( n31365 , n17606 , n32624 );
    and g30565 ( n2981 , n17064 , n18843 );
    not g30566 ( n1892 , n14911 );
    and g30567 ( n17181 , n18990 , n2036 );
    xnor g30568 ( n8823 , n3014 , n5546 );
    or g30569 ( n27372 , n21748 , n18219 );
    or g30570 ( n2181 , n32095 , n6867 );
    xnor g30571 ( n19100 , n15149 , n31714 );
    or g30572 ( n17282 , n9552 , n24836 );
    or g30573 ( n25135 , n8078 , n30698 );
    xnor g30574 ( n6015 , n16207 , n9658 );
    or g30575 ( n7952 , n11046 , n26973 );
    or g30576 ( n4082 , n27271 , n6191 );
    not g30577 ( n34534 , n13560 );
    buf g30578 ( n35938 , n20255 );
    or g30579 ( n7848 , n14584 , n18533 );
    xnor g30580 ( n18857 , n18802 , n16620 );
    and g30581 ( n24363 , n19270 , n9324 );
    or g30582 ( n30143 , n16922 , n31461 );
    or g30583 ( n24230 , n16612 , n29953 );
    nor g30584 ( n3109 , n9209 , n1215 );
    or g30585 ( n34419 , n22240 , n21037 );
    or g30586 ( n12676 , n4863 , n24868 );
    and g30587 ( n3821 , n11449 , n11451 );
    and g30588 ( n32515 , n5665 , n33247 );
    nor g30589 ( n26058 , n25436 , n13960 );
    and g30590 ( n615 , n4669 , n23582 );
    nor g30591 ( n16426 , n4519 , n19285 );
    and g30592 ( n101 , n29284 , n21340 );
    or g30593 ( n21552 , n18601 , n30708 );
    or g30594 ( n6239 , n7540 , n3628 );
    or g30595 ( n23474 , n15843 , n13307 );
    or g30596 ( n19175 , n14785 , n19421 );
    or g30597 ( n16193 , n3888 , n35244 );
    or g30598 ( n22072 , n26969 , n128 );
    xnor g30599 ( n5282 , n32508 , n18127 );
    or g30600 ( n2552 , n14437 , n5168 );
    not g30601 ( n21594 , n1554 );
    or g30602 ( n29738 , n7819 , n34084 );
    or g30603 ( n20112 , n35880 , n8210 );
    or g30604 ( n13363 , n1427 , n1922 );
    or g30605 ( n23137 , n28215 , n19895 );
    and g30606 ( n23840 , n10708 , n21934 );
    not g30607 ( n986 , n33856 );
    and g30608 ( n1996 , n23790 , n26543 );
    and g30609 ( n29835 , n32831 , n5181 );
    xnor g30610 ( n14296 , n1660 , n35927 );
    xnor g30611 ( n12352 , n11223 , n31272 );
    and g30612 ( n6473 , n8826 , n14951 );
    or g30613 ( n23144 , n16665 , n14076 );
    nor g30614 ( n25220 , n12734 , n33956 );
    xnor g30615 ( n16160 , n34059 , n24094 );
    and g30616 ( n19568 , n5918 , n11395 );
    or g30617 ( n29012 , n10357 , n9921 );
    or g30618 ( n4163 , n29985 , n202 );
    and g30619 ( n25664 , n9424 , n7575 );
    or g30620 ( n18866 , n20985 , n4779 );
    xnor g30621 ( n31206 , n17603 , n16125 );
    or g30622 ( n20351 , n23854 , n32697 );
    and g30623 ( n26556 , n21713 , n22284 );
    or g30624 ( n28071 , n13955 , n17162 );
    xnor g30625 ( n28063 , n17442 , n10861 );
    and g30626 ( n19425 , n30830 , n25815 );
    xnor g30627 ( n10788 , n2008 , n11665 );
    not g30628 ( n27209 , n19009 );
    or g30629 ( n16895 , n22885 , n4775 );
    xnor g30630 ( n6598 , n15695 , n24839 );
    or g30631 ( n18449 , n25742 , n27574 );
    xnor g30632 ( n15821 , n7925 , n28477 );
    or g30633 ( n4759 , n9793 , n7488 );
    or g30634 ( n6580 , n141 , n13307 );
    nor g30635 ( n1437 , n29756 , n26549 );
    or g30636 ( n12587 , n33424 , n6306 );
    not g30637 ( n34674 , n4232 );
    or g30638 ( n23458 , n15531 , n28574 );
    or g30639 ( n32849 , n7050 , n9915 );
    and g30640 ( n27850 , n11591 , n6304 );
    or g30641 ( n13195 , n2284 , n32425 );
    and g30642 ( n32537 , n22666 , n17080 );
    xnor g30643 ( n4876 , n20098 , n20272 );
    xnor g30644 ( n10073 , n35344 , n5277 );
    and g30645 ( n10409 , n8034 , n33214 );
    and g30646 ( n30354 , n24234 , n24461 );
    or g30647 ( n7549 , n28855 , n13305 );
    or g30648 ( n11845 , n22291 , n29208 );
    not g30649 ( n22751 , n31559 );
    nor g30650 ( n12692 , n16953 , n29366 );
    and g30651 ( n24349 , n7949 , n23515 );
    and g30652 ( n9316 , n6090 , n36082 );
    or g30653 ( n14860 , n25957 , n28248 );
    or g30654 ( n26959 , n25987 , n9317 );
    xnor g30655 ( n34021 , n5324 , n24371 );
    or g30656 ( n33671 , n25602 , n7385 );
    or g30657 ( n10057 , n27291 , n376 );
    or g30658 ( n23528 , n16027 , n35141 );
    xnor g30659 ( n27841 , n24698 , n2056 );
    or g30660 ( n28457 , n23606 , n19816 );
    or g30661 ( n8531 , n33473 , n29127 );
    and g30662 ( n14444 , n29200 , n16117 );
    xnor g30663 ( n34791 , n16381 , n27570 );
    or g30664 ( n15933 , n32970 , n8450 );
    xnor g30665 ( n18507 , n6481 , n22663 );
    nor g30666 ( n25920 , n29839 , n4624 );
    xnor g30667 ( n25294 , n33024 , n33168 );
    not g30668 ( n30221 , n21801 );
    and g30669 ( n15669 , n18804 , n31347 );
    or g30670 ( n24690 , n34830 , n6233 );
    or g30671 ( n26805 , n31399 , n11536 );
    and g30672 ( n28640 , n21988 , n17708 );
    or g30673 ( n11856 , n25602 , n25292 );
    buf g30674 ( n4203 , n8869 );
    xnor g30675 ( n30855 , n17075 , n4288 );
    xor g30676 ( n14871 , n1051 , n33641 );
    or g30677 ( n34504 , n17784 , n8802 );
    and g30678 ( n8423 , n10732 , n10667 );
    or g30679 ( n30761 , n29157 , n18126 );
    or g30680 ( n2787 , n15075 , n34549 );
    xnor g30681 ( n8893 , n14231 , n30461 );
    xor g30682 ( n35121 , n5129 , n16514 );
    or g30683 ( n1677 , n7363 , n1715 );
    buf g30684 ( n13664 , n13015 );
    nor g30685 ( n35813 , n35927 , n22089 );
    not g30686 ( n1273 , n31602 );
    and g30687 ( n10277 , n22380 , n23240 );
    or g30688 ( n9086 , n19663 , n21977 );
    or g30689 ( n31428 , n27395 , n538 );
    and g30690 ( n10003 , n15189 , n29924 );
    and g30691 ( n20157 , n27662 , n26937 );
    or g30692 ( n24154 , n33099 , n3858 );
    or g30693 ( n3941 , n15912 , n16762 );
    xnor g30694 ( n31875 , n4603 , n31272 );
    not g30695 ( n6436 , n25477 );
    and g30696 ( n30010 , n12099 , n20495 );
    or g30697 ( n26024 , n26474 , n15290 );
    or g30698 ( n27648 , n6915 , n30751 );
    xnor g30699 ( n20130 , n27235 , n3082 );
    or g30700 ( n2058 , n3525 , n1414 );
    or g30701 ( n25946 , n33774 , n2119 );
    xnor g30702 ( n35884 , n4624 , n11463 );
    and g30703 ( n29975 , n17817 , n25722 );
    xnor g30704 ( n31416 , n26447 , n10894 );
    or g30705 ( n14034 , n30745 , n29953 );
    and g30706 ( n10381 , n5647 , n31350 );
    not g30707 ( n23231 , n16366 );
    and g30708 ( n17716 , n10824 , n24090 );
    xnor g30709 ( n32402 , n1446 , n26937 );
    or g30710 ( n24854 , n10894 , n25523 );
    or g30711 ( n30436 , n28187 , n19336 );
    nor g30712 ( n7776 , n7418 , n25209 );
    xnor g30713 ( n31297 , n27505 , n25602 );
    or g30714 ( n27412 , n10843 , n22144 );
    xnor g30715 ( n12401 , n8238 , n29713 );
    and g30716 ( n22765 , n33050 , n15955 );
    or g30717 ( n2110 , n21366 , n15344 );
    nor g30718 ( n27118 , n3779 , n5779 );
    and g30719 ( n23020 , n131 , n32455 );
    and g30720 ( n19656 , n11168 , n35015 );
    or g30721 ( n6144 , n8229 , n24061 );
    and g30722 ( n9435 , n23753 , n6246 );
    or g30723 ( n31858 , n31056 , n17754 );
    xnor g30724 ( n34812 , n29058 , n15886 );
    or g30725 ( n24995 , n14165 , n885 );
    nor g30726 ( n23503 , n33493 , n10416 );
    and g30727 ( n22766 , n28162 , n24291 );
    not g30728 ( n23638 , n3317 );
    or g30729 ( n21886 , n36022 , n26480 );
    xnor g30730 ( n999 , n14827 , n4960 );
    xnor g30731 ( n29060 , n14592 , n3946 );
    and g30732 ( n16841 , n33404 , n2289 );
    or g30733 ( n30315 , n25552 , n16456 );
    and g30734 ( n18441 , n24771 , n6628 );
    or g30735 ( n4474 , n712 , n10960 );
    and g30736 ( n16760 , n6327 , n490 );
    or g30737 ( n602 , n4288 , n14108 );
    or g30738 ( n8177 , n32857 , n22939 );
    or g30739 ( n18945 , n11152 , n16471 );
    or g30740 ( n34158 , n33507 , n5717 );
    nor g30741 ( n15780 , n10298 , n33399 );
    xnor g30742 ( n24447 , n20490 , n31559 );
    or g30743 ( n15447 , n6627 , n30431 );
    or g30744 ( n8161 , n28747 , n10385 );
    or g30745 ( n29110 , n20670 , n22477 );
    not g30746 ( n29062 , n28273 );
    and g30747 ( n4311 , n23143 , n1263 );
    or g30748 ( n32654 , n18724 , n1996 );
    or g30749 ( n35799 , n23577 , n33152 );
    or g30750 ( n2766 , n20542 , n31055 );
    not g30751 ( n7712 , n32857 );
    xnor g30752 ( n35351 , n34907 , n15814 );
    or g30753 ( n11427 , n23604 , n9850 );
    and g30754 ( n31104 , n17969 , n14806 );
    or g30755 ( n15204 , n1066 , n7527 );
    or g30756 ( n30403 , n34938 , n16543 );
    and g30757 ( n21343 , n32240 , n34388 );
    and g30758 ( n7637 , n12561 , n18329 );
    or g30759 ( n6099 , n19731 , n35124 );
    or g30760 ( n15069 , n24281 , n10417 );
    xnor g30761 ( n20643 , n9288 , n4758 );
    xnor g30762 ( n32341 , n6402 , n9789 );
    and g30763 ( n10306 , n18145 , n15775 );
    and g30764 ( n35868 , n29483 , n3791 );
    or g30765 ( n34145 , n23604 , n31012 );
    xnor g30766 ( n15882 , n6206 , n30742 );
    or g30767 ( n30015 , n14445 , n128 );
    nor g30768 ( n22591 , n35537 , n33192 );
    and g30769 ( n27211 , n25734 , n21005 );
    xnor g30770 ( n33456 , n34691 , n15886 );
    not g30771 ( n11960 , n2540 );
    nor g30772 ( n4351 , n16620 , n33525 );
    xnor g30773 ( n5074 , n22264 , n24695 );
    or g30774 ( n5406 , n35739 , n19125 );
    or g30775 ( n11517 , n8081 , n21042 );
    and g30776 ( n6857 , n6411 , n23094 );
    and g30777 ( n31243 , n1614 , n18813 );
    and g30778 ( n19843 , n9987 , n35130 );
    or g30779 ( n29055 , n13529 , n31554 );
    or g30780 ( n10263 , n30659 , n19173 );
    and g30781 ( n24093 , n31473 , n26943 );
    xnor g30782 ( n26628 , n17222 , n460 );
    or g30783 ( n22171 , n2812 , n22616 );
    and g30784 ( n1678 , n35085 , n20439 );
    xnor g30785 ( n6145 , n19049 , n31049 );
    or g30786 ( n18284 , n31289 , n30326 );
    or g30787 ( n210 , n830 , n14610 );
    or g30788 ( n19872 , n6856 , n34379 );
    and g30789 ( n987 , n25059 , n29762 );
    and g30790 ( n20605 , n25643 , n22059 );
    xnor g30791 ( n18659 , n28968 , n12899 );
    xnor g30792 ( n9341 , n9885 , n564 );
    or g30793 ( n5131 , n14009 , n11833 );
    and g30794 ( n29622 , n6354 , n35477 );
    xnor g30795 ( n3578 , n14865 , n33457 );
    or g30796 ( n18960 , n15739 , n26292 );
    or g30797 ( n33938 , n17139 , n19464 );
    buf g30798 ( n24479 , n32071 );
    or g30799 ( n6389 , n35927 , n10367 );
    and g30800 ( n2619 , n8065 , n14860 );
    or g30801 ( n34550 , n25602 , n4609 );
    and g30802 ( n16616 , n4096 , n9485 );
    not g30803 ( n12778 , n22291 );
    or g30804 ( n32347 , n35927 , n13681 );
    or g30805 ( n17807 , n22364 , n25648 );
    or g30806 ( n35013 , n4962 , n3921 );
    or g30807 ( n1893 , n21539 , n34862 );
    or g30808 ( n2640 , n16384 , n8750 );
    xnor g30809 ( n335 , n22633 , n15952 );
    and g30810 ( n18925 , n9511 , n22980 );
    nor g30811 ( n12076 , n1981 , n10301 );
    and g30812 ( n23013 , n2004 , n18389 );
    buf g30813 ( n4490 , n6521 );
    nor g30814 ( n15610 , n836 , n10428 );
    or g30815 ( n1170 , n21057 , n16797 );
    xnor g30816 ( n19122 , n6480 , n21587 );
    or g30817 ( n19174 , n34035 , n28548 );
    or g30818 ( n12435 , n13843 , n4363 );
    nor g30819 ( n23536 , n8242 , n13757 );
    xnor g30820 ( n6140 , n10638 , n14152 );
    or g30821 ( n17088 , n5287 , n18918 );
    xor g30822 ( n29655 , n27803 , n31799 );
    xnor g30823 ( n8234 , n1087 , n4288 );
    or g30824 ( n2425 , n32095 , n16992 );
    or g30825 ( n22827 , n25877 , n29658 );
    or g30826 ( n4133 , n16620 , n30709 );
    xnor g30827 ( n33788 , n22080 , n25174 );
    or g30828 ( n17392 , n20173 , n3738 );
    and g30829 ( n1061 , n28885 , n9829 );
    or g30830 ( n34247 , n1972 , n31757 );
    or g30831 ( n32914 , n25602 , n4120 );
    and g30832 ( n21704 , n29126 , n30309 );
    xnor g30833 ( n11320 , n13340 , n17568 );
    or g30834 ( n1994 , n8178 , n2168 );
    not g30835 ( n29484 , n13659 );
    or g30836 ( n9678 , n2053 , n21839 );
    or g30837 ( n31831 , n347 , n17046 );
    xnor g30838 ( n7767 , n27149 , n11778 );
    or g30839 ( n11629 , n29713 , n4662 );
    buf g30840 ( n24696 , n14018 );
    and g30841 ( n20572 , n6601 , n12411 );
    or g30842 ( n2847 , n27761 , n20104 );
    xnor g30843 ( n16448 , n7663 , n33799 );
    or g30844 ( n7459 , n30154 , n11258 );
    not g30845 ( n5395 , n16223 );
    or g30846 ( n20861 , n33993 , n1557 );
    and g30847 ( n4801 , n9669 , n15083 );
    and g30848 ( n34665 , n35581 , n4153 );
    or g30849 ( n20630 , n8876 , n5707 );
    xnor g30850 ( n9310 , n32137 , n24548 );
    or g30851 ( n6971 , n4758 , n5921 );
    or g30852 ( n32582 , n6551 , n6677 );
    xnor g30853 ( n7281 , n7651 , n4962 );
    and g30854 ( n4757 , n24399 , n26031 );
    or g30855 ( n7037 , n8642 , n20762 );
    nor g30856 ( n18644 , n35163 , n25825 );
    or g30857 ( n4563 , n7572 , n25567 );
    not g30858 ( n21167 , n30158 );
    or g30859 ( n19220 , n23604 , n33918 );
    or g30860 ( n33470 , n6398 , n19543 );
    xnor g30861 ( n6852 , n11300 , n27631 );
    or g30862 ( n35098 , n26254 , n2823 );
    and g30863 ( n8745 , n20879 , n24711 );
    or g30864 ( n24625 , n26381 , n32124 );
    and g30865 ( n26483 , n32303 , n17136 );
    and g30866 ( n12044 , n29087 , n23144 );
    and g30867 ( n28830 , n21025 , n23216 );
    or g30868 ( n18736 , n18415 , n14076 );
    or g30869 ( n16099 , n20572 , n33416 );
    xnor g30870 ( n18370 , n35556 , n5067 );
    or g30871 ( n33453 , n10594 , n3388 );
    and g30872 ( n2078 , n27797 , n6858 );
    or g30873 ( n10259 , n10992 , n4464 );
    or g30874 ( n30480 , n22256 , n17337 );
    or g30875 ( n1595 , n33360 , n24696 );
    or g30876 ( n12772 , n35500 , n15248 );
    and g30877 ( n9051 , n1179 , n26526 );
    xor g30878 ( n29152 , n10992 , n4464 );
    xnor g30879 ( n35012 , n18531 , n29302 );
    and g30880 ( n28407 , n12629 , n18805 );
    and g30881 ( n22079 , n13339 , n14074 );
    nor g30882 ( n23901 , n5287 , n30716 );
    or g30883 ( n2551 , n12387 , n12470 );
    or g30884 ( n6977 , n21180 , n13267 );
    nor g30885 ( n33843 , n15515 , n27672 );
    xnor g30886 ( n30278 , n8901 , n17685 );
    not g30887 ( n14409 , n15042 );
    not g30888 ( n26245 , n5864 );
    or g30889 ( n24733 , n20235 , n23921 );
    or g30890 ( n27187 , n29225 , n19336 );
    and g30891 ( n33485 , n20102 , n16255 );
    and g30892 ( n26687 , n18226 , n34954 );
    or g30893 ( n28239 , n6310 , n14554 );
    and g30894 ( n5619 , n12863 , n4963 );
    and g30895 ( n5552 , n8193 , n18953 );
    or g30896 ( n3878 , n29287 , n26112 );
    and g30897 ( n16876 , n29992 , n36032 );
    not g30898 ( n11227 , n3742 );
    or g30899 ( n3153 , n21225 , n578 );
    xnor g30900 ( n12699 , n27763 , n752 );
    xnor g30901 ( n12726 , n9226 , n20228 );
    or g30902 ( n15897 , n28490 , n13305 );
    or g30903 ( n21698 , n30132 , n28675 );
    or g30904 ( n15801 , n29713 , n32083 );
    not g30905 ( n7858 , n22291 );
    and g30906 ( n16533 , n28324 , n3101 );
    or g30907 ( n20720 , n15697 , n20579 );
    and g30908 ( n35917 , n3757 , n22980 );
    xnor g30909 ( n34849 , n12713 , n5309 );
    or g30910 ( n13439 , n29839 , n26706 );
    and g30911 ( n7657 , n26836 , n17391 );
    or g30912 ( n10323 , n127 , n21914 );
    nor g30913 ( n2444 , n15299 , n17687 );
    xnor g30914 ( n27602 , n21285 , n14507 );
    or g30915 ( n32014 , n14194 , n18189 );
    or g30916 ( n19264 , n7917 , n15899 );
    and g30917 ( n18474 , n25513 , n28772 );
    not g30918 ( n30951 , n16315 );
    xnor g30919 ( n24037 , n29501 , n28113 );
    or g30920 ( n25950 , n23920 , n3858 );
    and g30921 ( n33460 , n21745 , n6155 );
    or g30922 ( n10646 , n25330 , n34727 );
    or g30923 ( n30198 , n7164 , n26690 );
    or g30924 ( n25143 , n15727 , n13305 );
    and g30925 ( n26443 , n12383 , n28411 );
    xnor g30926 ( n32183 , n28554 , n12228 );
    or g30927 ( n31201 , n7973 , n32929 );
    and g30928 ( n23292 , n3755 , n5861 );
    or g30929 ( n5191 , n7540 , n8435 );
    or g30930 ( n8670 , n24371 , n6912 );
    or g30931 ( n18401 , n32584 , n15991 );
    or g30932 ( n32318 , n29884 , n1741 );
    or g30933 ( n7617 , n6364 , n25647 );
    or g30934 ( n1157 , n4017 , n26365 );
    or g30935 ( n722 , n1785 , n14918 );
    and g30936 ( n18661 , n6243 , n27894 );
    xnor g30937 ( n18462 , n11225 , n17751 );
    or g30938 ( n31963 , n25065 , n19336 );
    xnor g30939 ( n33073 , n9326 , n3383 );
    and g30940 ( n3138 , n33790 , n21473 );
    or g30941 ( n5239 , n11190 , n21808 );
    or g30942 ( n24278 , n23604 , n32202 );
    or g30943 ( n13645 , n34341 , n13307 );
    and g30944 ( n30725 , n31248 , n31719 );
    not g30945 ( n35173 , n10600 );
    or g30946 ( n22849 , n4406 , n6340 );
    and g30947 ( n10707 , n3688 , n22038 );
    xnor g30948 ( n15353 , n34815 , n29713 );
    and g30949 ( n29790 , n18584 , n35927 );
    or g30950 ( n8918 , n34168 , n10499 );
    or g30951 ( n600 , n4304 , n21042 );
    or g30952 ( n35922 , n23518 , n8537 );
    or g30953 ( n17197 , n4288 , n19420 );
    and g30954 ( n20552 , n4163 , n13561 );
    and g30955 ( n35951 , n9996 , n6784 );
    or g30956 ( n13309 , n18034 , n12879 );
    or g30957 ( n27776 , n21891 , n10394 );
    or g30958 ( n29596 , n11046 , n24312 );
    or g30959 ( n5975 , n29698 , n25272 );
    or g30960 ( n14125 , n35927 , n8655 );
    xnor g30961 ( n32907 , n12845 , n24371 );
    or g30962 ( n7468 , n6512 , n16594 );
    or g30963 ( n25780 , n9789 , n27037 );
    and g30964 ( n24730 , n32783 , n15839 );
    and g30965 ( n142 , n30997 , n4092 );
    or g30966 ( n28241 , n680 , n14997 );
    xnor g30967 ( n7024 , n1655 , n34822 );
    or g30968 ( n25341 , n29137 , n9661 );
    and g30969 ( n10225 , n16496 , n34908 );
    and g30970 ( n35296 , n30482 , n17122 );
    or g30971 ( n17020 , n9658 , n15047 );
    xnor g30972 ( n33792 , n3542 , n19107 );
    or g30973 ( n17954 , n27649 , n17765 );
    or g30974 ( n944 , n6033 , n30646 );
    or g30975 ( n6163 , n35007 , n36079 );
    nor g30976 ( n13465 , n12547 , n35340 );
    and g30977 ( n1515 , n5885 , n23720 );
    and g30978 ( n5299 , n4148 , n25557 );
    or g30979 ( n28436 , n11190 , n13563 );
    or g30980 ( n6706 , n18309 , n35748 );
    and g30981 ( n34452 , n17728 , n1717 );
    and g30982 ( n30798 , n15471 , n27273 );
    and g30983 ( n1245 , n17838 , n33111 );
    or g30984 ( n27633 , n5840 , n28797 );
    not g30985 ( n32500 , n18366 );
    or g30986 ( n17143 , n168 , n20817 );
    not g30987 ( n25051 , n13651 );
    not g30988 ( n29071 , n12772 );
    or g30989 ( n34976 , n14940 , n11209 );
    xnor g30990 ( n5024 , n3628 , n7540 );
    not g30991 ( n29033 , n22501 );
    and g30992 ( n13518 , n16406 , n4003 );
    and g30993 ( n18046 , n20667 , n23779 );
    or g30994 ( n4012 , n14393 , n1402 );
    xnor g30995 ( n13485 , n34829 , n8432 );
    xnor g30996 ( n32008 , n23920 , n4288 );
    not g30997 ( n122 , n16223 );
    not g30998 ( n30457 , n25762 );
    or g30999 ( n1585 , n3222 , n34541 );
    and g31000 ( n5151 , n24846 , n16842 );
    or g31001 ( n24006 , n4587 , n23187 );
    nor g31002 ( n21466 , n4641 , n17893 );
    or g31003 ( n23159 , n22056 , n28934 );
    or g31004 ( n19739 , n20705 , n25725 );
    nor g31005 ( n10175 , n830 , n8186 );
    xnor g31006 ( n20076 , n16972 , n32715 );
    or g31007 ( n15761 , n3771 , n6366 );
    not g31008 ( n14035 , n32480 );
    or g31009 ( n27002 , n16678 , n21993 );
    not g31010 ( n32086 , n15936 );
    not g31011 ( n33455 , n33524 );
    and g31012 ( n18734 , n33059 , n9212 );
    not g31013 ( n29644 , n29713 );
    xnor g31014 ( n31588 , n16741 , n30433 );
    nor g31015 ( n30449 , n29427 , n5397 );
    not g31016 ( n20701 , n12666 );
    and g31017 ( n9091 , n10738 , n4650 );
    or g31018 ( n24464 , n31056 , n26621 );
    xnor g31019 ( n32643 , n6980 , n28186 );
    not g31020 ( n22330 , n11190 );
    or g31021 ( n21568 , n9418 , n2712 );
    xnor g31022 ( n28561 , n23760 , n13939 );
    and g31023 ( n10340 , n24894 , n10141 );
    and g31024 ( n16191 , n5605 , n22582 );
    and g31025 ( n20395 , n29615 , n4290 );
    or g31026 ( n10419 , n7301 , n30204 );
    and g31027 ( n27066 , n29922 , n25491 );
    or g31028 ( n30213 , n6247 , n24165 );
    or g31029 ( n21988 , n18814 , n30287 );
    xnor g31030 ( n25616 , n22287 , n29930 );
    and g31031 ( n18165 , n21945 , n9991 );
    or g31032 ( n23193 , n26348 , n26852 );
    xnor g31033 ( n25055 , n28110 , n25777 );
    and g31034 ( n28306 , n19355 , n30918 );
    and g31035 ( n19260 , n14729 , n21133 );
    or g31036 ( n24145 , n20527 , n2295 );
    and g31037 ( n5719 , n27129 , n5542 );
    or g31038 ( n15364 , n3375 , n28837 );
    or g31039 ( n26535 , n14967 , n9698 );
    or g31040 ( n31631 , n20871 , n10849 );
    and g31041 ( n18544 , n34729 , n23862 );
    xnor g31042 ( n525 , n30180 , n29214 );
    xnor g31043 ( n4002 , n17812 , n31289 );
    and g31044 ( n33326 , n5458 , n20935 );
    or g31045 ( n18869 , n27102 , n27447 );
    or g31046 ( n551 , n29839 , n11537 );
    xnor g31047 ( n5361 , n20832 , n32095 );
    or g31048 ( n32231 , n17751 , n6701 );
    and g31049 ( n35772 , n15500 , n8361 );
    not g31050 ( n35949 , n10427 );
    nor g31051 ( n28698 , n16620 , n14960 );
    not g31052 ( n18065 , n12622 );
    and g31053 ( n28291 , n15386 , n3899 );
    or g31054 ( n490 , n15886 , n11846 );
    or g31055 ( n30778 , n13870 , n29953 );
    and g31056 ( n4727 , n6150 , n13990 );
    and g31057 ( n29018 , n28575 , n1521 );
    or g31058 ( n23423 , n7385 , n559 );
    or g31059 ( n736 , n6472 , n17872 );
    or g31060 ( n5895 , n4962 , n6680 );
    and g31061 ( n12685 , n12430 , n4949 );
    and g31062 ( n33219 , n4138 , n23164 );
    or g31063 ( n10605 , n36013 , n2351 );
    or g31064 ( n23074 , n32714 , n24672 );
    or g31065 ( n26446 , n18442 , n8221 );
    or g31066 ( n35364 , n27291 , n36035 );
    and g31067 ( n31375 , n17013 , n15569 );
    or g31068 ( n12839 , n14624 , n20427 );
    xnor g31069 ( n15373 , n22362 , n178 );
    or g31070 ( n24253 , n8965 , n19058 );
    and g31071 ( n11772 , n20423 , n19453 );
    xnor g31072 ( n24754 , n9243 , n34417 );
    xnor g31073 ( n16407 , n5550 , n6061 );
    and g31074 ( n27996 , n24938 , n15061 );
    xnor g31075 ( n1902 , n2956 , n30753 );
    and g31076 ( n2108 , n5267 , n16408 );
    and g31077 ( n28502 , n2219 , n29165 );
    buf g31078 ( n32959 , n34084 );
    and g31079 ( n24300 , n22323 , n30398 );
    or g31080 ( n23186 , n35840 , n34540 );
    and g31081 ( n22198 , n1861 , n14602 );
    or g31082 ( n6458 , n24900 , n9915 );
    or g31083 ( n8447 , n11081 , n23163 );
    and g31084 ( n35944 , n15008 , n10547 );
    or g31085 ( n4331 , n8488 , n30646 );
    nor g31086 ( n12049 , n5981 , n29203 );
    or g31087 ( n7305 , n24371 , n6348 );
    or g31088 ( n2001 , n20086 , n29014 );
    or g31089 ( n16540 , n6393 , n16184 );
    xnor g31090 ( n27109 , n14709 , n9789 );
    or g31091 ( n21139 , n3299 , n24433 );
    and g31092 ( n33993 , n24217 , n15328 );
    xnor g31093 ( n24248 , n12263 , n2042 );
    or g31094 ( n35804 , n12394 , n21208 );
    and g31095 ( n19457 , n4253 , n15992 );
    or g31096 ( n28234 , n4758 , n20099 );
    nor g31097 ( n32030 , n17568 , n24315 );
    nor g31098 ( n31386 , n7540 , n28066 );
    and g31099 ( n34218 , n14815 , n3000 );
    or g31100 ( n23716 , n21522 , n27094 );
    and g31101 ( n12855 , n33213 , n9980 );
    not g31102 ( n19547 , n7726 );
    and g31103 ( n9734 , n14760 , n35510 );
    xnor g31104 ( n32752 , n24385 , n21518 );
    or g31105 ( n2038 , n34176 , n35757 );
    and g31106 ( n16834 , n18575 , n1070 );
    or g31107 ( n31759 , n31782 , n24259 );
    or g31108 ( n27711 , n14836 , n30499 );
    or g31109 ( n30120 , n9722 , n6374 );
    and g31110 ( n1282 , n27788 , n1709 );
    xnor g31111 ( n3723 , n26423 , n9658 );
    xnor g31112 ( n10743 , n3403 , n5291 );
    and g31113 ( n456 , n1914 , n32681 );
    xnor g31114 ( n8817 , n8705 , n14249 );
    or g31115 ( n16458 , n25173 , n30519 );
    or g31116 ( n3192 , n11165 , n1968 );
    or g31117 ( n18774 , n16771 , n23650 );
    and g31118 ( n35766 , n8526 , n22368 );
    or g31119 ( n18818 , n29117 , n32821 );
    xnor g31120 ( n11015 , n27470 , n15464 );
    not g31121 ( n12563 , n18121 );
    xnor g31122 ( n12686 , n32465 , n35927 );
    or g31123 ( n33414 , n4288 , n3949 );
    or g31124 ( n31602 , n9287 , n34505 );
    xnor g31125 ( n14332 , n23034 , n3893 );
    nor g31126 ( n9396 , n3205 , n11333 );
    not g31127 ( n19783 , n13362 );
    xnor g31128 ( n19466 , n28849 , n31695 );
    xnor g31129 ( n22818 , n12741 , n21587 );
    or g31130 ( n28761 , n21610 , n31936 );
    xnor g31131 ( n15822 , n19145 , n29884 );
    not g31132 ( n13705 , n27120 );
    or g31133 ( n32118 , n9031 , n25019 );
    xnor g31134 ( n6409 , n23238 , n10029 );
    not g31135 ( n28215 , n35497 );
    xnor g31136 ( n32400 , n22199 , n6955 );
    or g31137 ( n6594 , n33705 , n405 );
    nor g31138 ( n32396 , n20484 , n30289 );
    or g31139 ( n23664 , n32095 , n10839 );
    and g31140 ( n21162 , n26367 , n21211 );
    or g31141 ( n4425 , n11377 , n9896 );
    xnor g31142 ( n19162 , n6796 , n23604 );
    or g31143 ( n705 , n4544 , n29373 );
    or g31144 ( n32221 , n24342 , n35402 );
    nor g31145 ( n5274 , n36036 , n3799 );
    or g31146 ( n1899 , n11612 , n6366 );
    xnor g31147 ( n15655 , n12110 , n18435 );
    buf g31148 ( n11218 , n10600 );
    xnor g31149 ( n16674 , n18709 , n21732 );
    nor g31150 ( n1424 , n20913 , n916 );
    and g31151 ( n29995 , n35021 , n30789 );
    xnor g31152 ( n17919 , n575 , n7540 );
    or g31153 ( n21957 , n28030 , n3634 );
    or g31154 ( n21572 , n4960 , n35801 );
    and g31155 ( n17139 , n34655 , n17719 );
    and g31156 ( n16660 , n26803 , n21004 );
    and g31157 ( n16396 , n35231 , n10921 );
    xnor g31158 ( n13550 , n6872 , n1744 );
    or g31159 ( n28131 , n3638 , n34084 );
    or g31160 ( n11093 , n15464 , n3100 );
    or g31161 ( n8795 , n21791 , n18433 );
    and g31162 ( n8276 , n6625 , n13753 );
    and g31163 ( n9872 , n35539 , n2631 );
    xnor g31164 ( n32859 , n4776 , n18830 );
    or g31165 ( n9598 , n15234 , n2384 );
    or g31166 ( n13321 , n35796 , n4363 );
    or g31167 ( n11926 , n10253 , n9437 );
    or g31168 ( n24354 , n4889 , n29592 );
    or g31169 ( n23497 , n4418 , n9555 );
    or g31170 ( n15220 , n23756 , n28668 );
    xnor g31171 ( n33522 , n18439 , n21938 );
    or g31172 ( n32256 , n30319 , n33979 );
    or g31173 ( n18213 , n8432 , n7654 );
    or g31174 ( n6087 , n830 , n7063 );
    and g31175 ( n11896 , n19479 , n11146 );
    nor g31176 ( n2980 , n25587 , n6276 );
    and g31177 ( n28262 , n4537 , n34394 );
    or g31178 ( n28897 , n30311 , n22959 );
    xnor g31179 ( n21863 , n27472 , n32095 );
    and g31180 ( n19772 , n9365 , n32072 );
    or g31181 ( n20497 , n31289 , n34349 );
    not g31182 ( n13144 , n12659 );
    xnor g31183 ( n1259 , n30133 , n31289 );
    and g31184 ( n24013 , n11930 , n6070 );
    or g31185 ( n14573 , n532 , n29926 );
    xnor g31186 ( n3367 , n15858 , n27593 );
    and g31187 ( n21193 , n24167 , n5321 );
    xnor g31188 ( n6696 , n19102 , n20590 );
    or g31189 ( n8592 , n18261 , n25842 );
    and g31190 ( n35763 , n10712 , n23810 );
    or g31191 ( n35470 , n34845 , n16456 );
    and g31192 ( n23820 , n6526 , n12847 );
    xnor g31193 ( n11134 , n10676 , n31289 );
    or g31194 ( n1075 , n17194 , n35748 );
    nor g31195 ( n19523 , n27655 , n31411 );
    nor g31196 ( n28973 , n27559 , n11837 );
    and g31197 ( n24346 , n4190 , n2203 );
    or g31198 ( n11950 , n17513 , n31055 );
    and g31199 ( n33158 , n21388 , n25666 );
    xnor g31200 ( n21536 , n29733 , n4956 );
    or g31201 ( n15049 , n23604 , n4233 );
    and g31202 ( n26128 , n34868 , n20763 );
    or g31203 ( n21952 , n33223 , n20840 );
    or g31204 ( n6132 , n35542 , n13247 );
    not g31205 ( n14268 , n14226 );
    or g31206 ( n744 , n32584 , n29589 );
    or g31207 ( n15570 , n23486 , n27234 );
    nor g31208 ( n4098 , n4962 , n15197 );
    xnor g31209 ( n35546 , n31993 , n33141 );
    xnor g31210 ( n13243 , n17304 , n16571 );
    or g31211 ( n14829 , n19409 , n9074 );
    or g31212 ( n32894 , n15040 , n9675 );
    and g31213 ( n6275 , n24989 , n35695 );
    or g31214 ( n4864 , n10855 , n12996 );
    or g31215 ( n29017 , n34754 , n6288 );
    and g31216 ( n1132 , n31828 , n15840 );
    xnor g31217 ( n6368 , n4050 , n3222 );
    or g31218 ( n23036 , n7202 , n19952 );
    and g31219 ( n21502 , n27468 , n29702 );
    and g31220 ( n4682 , n3151 , n23816 );
    and g31221 ( n22685 , n3987 , n32024 );
    and g31222 ( n18974 , n32817 , n24284 );
    nor g31223 ( n24893 , n35169 , n23719 );
    or g31224 ( n30361 , n35707 , n12230 );
    or g31225 ( n17461 , n30146 , n16457 );
    or g31226 ( n16401 , n30034 , n9194 );
    nor g31227 ( n7947 , n4962 , n19283 );
    and g31228 ( n9936 , n1489 , n24269 );
    xnor g31229 ( n22638 , n11318 , n12221 );
    nor g31230 ( n32003 , n34649 , n8892 );
    xnor g31231 ( n10167 , n9039 , n26538 );
    or g31232 ( n8381 , n28123 , n6305 );
    nor g31233 ( n2312 , n25174 , n25312 );
    or g31234 ( n13688 , n28119 , n21071 );
    or g31235 ( n5586 , n10788 , n22682 );
    and g31236 ( n11027 , n12239 , n5198 );
    and g31237 ( n21585 , n32960 , n3355 );
    or g31238 ( n29922 , n6772 , n2005 );
    or g31239 ( n16071 , n20511 , n26737 );
    and g31240 ( n17451 , n22545 , n20741 );
    or g31241 ( n30208 , n20250 , n23921 );
    xnor g31242 ( n3245 , n549 , n4928 );
    or g31243 ( n35378 , n4962 , n11164 );
    or g31244 ( n9685 , n15915 , n15439 );
    or g31245 ( n17071 , n24200 , n7287 );
    and g31246 ( n21630 , n1329 , n23021 );
    and g31247 ( n8473 , n31117 , n28956 );
    and g31248 ( n26561 , n23724 , n35863 );
    and g31249 ( n8237 , n7053 , n5414 );
    xor g31250 ( n16015 , n8644 , n24413 );
    not g31251 ( n216 , n27437 );
    not g31252 ( n1513 , n22678 );
    and g31253 ( n24389 , n35658 , n21744 );
    or g31254 ( n11411 , n16922 , n3058 );
    or g31255 ( n35809 , n3222 , n913 );
    and g31256 ( n324 , n20641 , n4623 );
    or g31257 ( n13319 , n14784 , n19167 );
    or g31258 ( n24266 , n7733 , n16543 );
    or g31259 ( n28883 , n7540 , n20582 );
    or g31260 ( n6111 , n30734 , n13362 );
    xnor g31261 ( n10674 , n7112 , n26347 );
    and g31262 ( n2653 , n6041 , n11989 );
    or g31263 ( n29820 , n31215 , n18260 );
    or g31264 ( n6203 , n23411 , n17872 );
    or g31265 ( n8320 , n10894 , n30161 );
    xnor g31266 ( n22169 , n1963 , n29963 );
    or g31267 ( n11325 , n22394 , n1942 );
    or g31268 ( n34525 , n2387 , n2814 );
    or g31269 ( n11450 , n32641 , n33435 );
    and g31270 ( n1693 , n30926 , n2465 );
    xnor g31271 ( n34265 , n33743 , n621 );
    or g31272 ( n8721 , n24397 , n7649 );
    or g31273 ( n25939 , n26601 , n35475 );
    or g31274 ( n14776 , n11148 , n21002 );
    and g31275 ( n29881 , n24266 , n9160 );
    xnor g31276 ( n21485 , n25930 , n19155 );
    xnor g31277 ( n23872 , n27277 , n23440 );
    nor g31278 ( n32447 , n18372 , n16497 );
    not g31279 ( n13402 , n21676 );
    or g31280 ( n29948 , n28500 , n16659 );
    nor g31281 ( n16526 , n9789 , n19249 );
    xnor g31282 ( n6633 , n35280 , n24261 );
    and g31283 ( n29631 , n7871 , n7280 );
    nor g31284 ( n6107 , n13524 , n34139 );
    xnor g31285 ( n2973 , n7310 , n3946 );
    xnor g31286 ( n33052 , n2678 , n14382 );
    xnor g31287 ( n2141 , n19791 , n23604 );
    not g31288 ( n13335 , n9789 );
    xnor g31289 ( n6421 , n19810 , n15403 );
    and g31290 ( n35694 , n5629 , n13844 );
    or g31291 ( n18135 , n830 , n17839 );
    xnor g31292 ( n2483 , n24920 , n31799 );
    and g31293 ( n14141 , n26349 , n33165 );
    xnor g31294 ( n23380 , n28139 , n9658 );
    and g31295 ( n17755 , n17100 , n31033 );
    or g31296 ( n18157 , n775 , n10950 );
    not g31297 ( n13376 , n10119 );
    nor g31298 ( n14924 , n3468 , n12392 );
    or g31299 ( n21650 , n33524 , n26594 );
    or g31300 ( n33626 , n11046 , n30401 );
    xnor g31301 ( n23961 , n4734 , n10402 );
    xnor g31302 ( n16800 , n11317 , n30060 );
    or g31303 ( n33675 , n7540 , n13674 );
    and g31304 ( n35666 , n17903 , n24423 );
    xnor g31305 ( n34547 , n32577 , n33124 );
    or g31306 ( n22854 , n4288 , n15641 );
    and g31307 ( n28367 , n8173 , n1809 );
    xnor g31308 ( n34438 , n11505 , n22456 );
    or g31309 ( n17318 , n11521 , n15604 );
    or g31310 ( n17799 , n28035 , n33585 );
    or g31311 ( n30402 , n12277 , n16343 );
    xnor g31312 ( n14042 , n12164 , n24332 );
    not g31313 ( n33499 , n24265 );
    or g31314 ( n23785 , n33102 , n772 );
    and g31315 ( n11872 , n17694 , n3392 );
    xnor g31316 ( n25361 , n18502 , n29794 );
    or g31317 ( n1281 , n33488 , n9301 );
    not g31318 ( n23446 , n8104 );
    and g31319 ( n19741 , n24153 , n21395 );
    and g31320 ( n13902 , n20756 , n23436 );
    or g31321 ( n32407 , n5879 , n3323 );
    or g31322 ( n708 , n31630 , n19125 );
    xnor g31323 ( n4636 , n25065 , n3946 );
    or g31324 ( n21987 , n15886 , n29058 );
    xnor g31325 ( n26524 , n33199 , n23453 );
    or g31326 ( n21713 , n28921 , n17964 );
    and g31327 ( n30779 , n6691 , n2807 );
    buf g31328 ( n25594 , n19403 );
    not g31329 ( n10445 , n17478 );
    or g31330 ( n9622 , n10087 , n30646 );
    and g31331 ( n812 , n23752 , n15365 );
    and g31332 ( n219 , n34191 , n28347 );
    or g31333 ( n2348 , n26390 , n13449 );
    xnor g31334 ( n16327 , n3444 , n28699 );
    xnor g31335 ( n23343 , n1673 , n18332 );
    xnor g31336 ( n1353 , n16759 , n30779 );
    or g31337 ( n23051 , n17771 , n22946 );
    or g31338 ( n7360 , n26293 , n15381 );
    nor g31339 ( n5716 , n3946 , n9055 );
    nor g31340 ( n29841 , n23070 , n19710 );
    xnor g31341 ( n33507 , n33146 , n31559 );
    or g31342 ( n28303 , n4170 , n13015 );
    or g31343 ( n8571 , n23743 , n15439 );
    or g31344 ( n33963 , n15886 , n6556 );
    and g31345 ( n11831 , n25956 , n16478 );
    xor g31346 ( n23956 , n34952 , n34400 );
    or g31347 ( n29774 , n7888 , n4318 );
    xnor g31348 ( n5214 , n25384 , n15464 );
    or g31349 ( n29919 , n3222 , n22909 );
    xnor g31350 ( n33150 , n30488 , n30917 );
    or g31351 ( n23274 , n14983 , n16659 );
    not g31352 ( n34121 , n33588 );
    or g31353 ( n6922 , n8434 , n9832 );
    or g31354 ( n30477 , n19209 , n15144 );
    or g31355 ( n28662 , n31272 , n9779 );
    or g31356 ( n33998 , n30855 , n32943 );
    nor g31357 ( n7585 , n15886 , n7428 );
    xnor g31358 ( n19844 , n381 , n13647 );
    xnor g31359 ( n28091 , n6393 , n16184 );
    xnor g31360 ( n7458 , n17722 , n31799 );
    or g31361 ( n20850 , n10990 , n23685 );
    or g31362 ( n34859 , n5287 , n23761 );
    nor g31363 ( n17906 , n35990 , n13978 );
    xnor g31364 ( n29807 , n35869 , n32095 );
    not g31365 ( n34634 , n18121 );
    xnor g31366 ( n30077 , n11798 , n16620 );
    or g31367 ( n31494 , n9692 , n4912 );
    or g31368 ( n13190 , n29625 , n32969 );
    nor g31369 ( n12859 , n4288 , n32266 );
    or g31370 ( n18304 , n23258 , n11996 );
    xnor g31371 ( n21175 , n31533 , n25468 );
    and g31372 ( n22338 , n13950 , n36043 );
    or g31373 ( n28694 , n20334 , n15034 );
    and g31374 ( n10632 , n20795 , n35925 );
    xnor g31375 ( n31317 , n19341 , n17751 );
    or g31376 ( n11769 , n1089 , n2698 );
    and g31377 ( n18130 , n11909 , n352 );
    or g31378 ( n6827 , n16922 , n11085 );
    not g31379 ( n22876 , n35410 );
    or g31380 ( n22773 , n33067 , n32507 );
    or g31381 ( n7052 , n29883 , n26192 );
    or g31382 ( n29409 , n3135 , n12923 );
    not g31383 ( n30476 , n28969 );
    or g31384 ( n28906 , n30980 , n25617 );
    or g31385 ( n8557 , n15886 , n21452 );
    or g31386 ( n17894 , n13269 , n31067 );
    or g31387 ( n25649 , n12509 , n32507 );
    buf g31388 ( n6374 , n25369 );
    xnor g31389 ( n9688 , n30693 , n20283 );
    or g31390 ( n6029 , n27274 , n11518 );
    and g31391 ( n13940 , n34197 , n20048 );
    and g31392 ( n11925 , n35795 , n15718 );
    or g31393 ( n15186 , n28356 , n11977 );
    and g31394 ( n899 , n4656 , n21438 );
    and g31395 ( n20506 , n16687 , n10807 );
    xnor g31396 ( n6416 , n26991 , n23716 );
    or g31397 ( n6638 , n26545 , n10409 );
    xnor g31398 ( n17759 , n3322 , n22928 );
    or g31399 ( n34104 , n30006 , n27574 );
    and g31400 ( n4428 , n21166 , n35654 );
    or g31401 ( n4777 , n31189 , n2823 );
    or g31402 ( n25270 , n25753 , n34064 );
    or g31403 ( n3407 , n32857 , n10425 );
    xnor g31404 ( n30538 , n33133 , n34766 );
    or g31405 ( n18041 , n9453 , n27973 );
    or g31406 ( n18298 , n7219 , n31514 );
    nor g31407 ( n29540 , n22401 , n25051 );
    and g31408 ( n9551 , n15651 , n34180 );
    and g31409 ( n14382 , n29021 , n35236 );
    or g31410 ( n12849 , n34403 , n32481 );
    or g31411 ( n8207 , n26091 , n22118 );
    nor g31412 ( n26161 , n4878 , n3687 );
    xnor g31413 ( n22533 , n8708 , n406 );
    or g31414 ( n33580 , n11156 , n9601 );
    or g31415 ( n25846 , n24455 , n10417 );
    and g31416 ( n19694 , n27340 , n26216 );
    xnor g31417 ( n5650 , n28838 , n17882 );
    not g31418 ( n20015 , n4758 );
    xnor g31419 ( n1408 , n12151 , n2730 );
    xnor g31420 ( n22031 , n11444 , n29446 );
    nor g31421 ( n8640 , n11678 , n21525 );
    xnor g31422 ( n20652 , n17208 , n10894 );
    xnor g31423 ( n19605 , n23558 , n16922 );
    or g31424 ( n12232 , n22725 , n11850 );
    not g31425 ( n7038 , n10576 );
    and g31426 ( n22577 , n8385 , n30428 );
    or g31427 ( n25513 , n19188 , n3422 );
    nor g31428 ( n9213 , n35482 , n27359 );
    or g31429 ( n24766 , n31982 , n27691 );
    or g31430 ( n5823 , n13587 , n16974 );
    and g31431 ( n19887 , n20618 , n11213 );
    nor g31432 ( n34275 , n29850 , n12900 );
    or g31433 ( n35206 , n10279 , n4363 );
    xnor g31434 ( n21596 , n19629 , n5335 );
    or g31435 ( n3925 , n39 , n4175 );
    nor g31436 ( n5429 , n15403 , n7891 );
    or g31437 ( n18249 , n29839 , n6272 );
    or g31438 ( n25184 , n28106 , n17125 );
    or g31439 ( n29812 , n34924 , n34862 );
    or g31440 ( n34065 , n10629 , n194 );
    and g31441 ( n36003 , n35366 , n22986 );
    or g31442 ( n11132 , n35506 , n14706 );
    xnor g31443 ( n22684 , n18779 , n307 );
    or g31444 ( n33351 , n15464 , n2786 );
    xnor g31445 ( n27027 , n32419 , n24332 );
    not g31446 ( n34557 , n35422 );
    and g31447 ( n13632 , n25706 , n967 );
    or g31448 ( n3728 , n1869 , n578 );
    or g31449 ( n2178 , n35927 , n19537 );
    and g31450 ( n13630 , n15318 , n16813 );
    or g31451 ( n34943 , n5028 , n24017 );
    xnor g31452 ( n10624 , n33920 , n18544 );
    not g31453 ( n8540 , n27291 );
    or g31454 ( n26007 , n30237 , n35744 );
    or g31455 ( n30568 , n8685 , n19464 );
    or g31456 ( n16013 , n29480 , n21691 );
    xnor g31457 ( n23541 , n34319 , n14190 );
    and g31458 ( n27512 , n21537 , n11736 );
    xnor g31459 ( n7430 , n10268 , n35841 );
    or g31460 ( n21537 , n5156 , n20616 );
    nor g31461 ( n13973 , n30553 , n22003 );
    xnor g31462 ( n23684 , n30479 , n19843 );
    xnor g31463 ( n15616 , n22256 , n15886 );
    or g31464 ( n28918 , n2308 , n32572 );
    xnor g31465 ( n22554 , n34894 , n10067 );
    and g31466 ( n24411 , n23680 , n11552 );
    or g31467 ( n22516 , n9281 , n14184 );
    not g31468 ( n2909 , n31056 );
    or g31469 ( n19132 , n3222 , n21112 );
    and g31470 ( n8566 , n4109 , n7540 );
    and g31471 ( n24281 , n15160 , n4402 );
    or g31472 ( n15968 , n27291 , n7507 );
    nor g31473 ( n19731 , n35927 , n11014 );
    or g31474 ( n8347 , n30270 , n20175 );
    or g31475 ( n3908 , n24765 , n30292 );
    and g31476 ( n7043 , n4320 , n3718 );
    or g31477 ( n12863 , n25772 , n32621 );
    or g31478 ( n7643 , n21143 , n5900 );
    or g31479 ( n1860 , n2922 , n3979 );
    xnor g31480 ( n7382 , n30677 , n17560 );
    or g31481 ( n24721 , n11540 , n31998 );
    not g31482 ( n19487 , n31593 );
    or g31483 ( n8019 , n27715 , n35935 );
    nor g31484 ( n18221 , n4758 , n1541 );
    or g31485 ( n14994 , n22692 , n2821 );
    or g31486 ( n4674 , n10681 , n8722 );
    or g31487 ( n2028 , n26128 , n763 );
    or g31488 ( n7988 , n245 , n25761 );
    or g31489 ( n6491 , n17562 , n11712 );
    or g31490 ( n33904 , n28975 , n26220 );
    or g31491 ( n4768 , n22665 , n22993 );
    or g31492 ( n5072 , n3231 , n35402 );
    or g31493 ( n902 , n3802 , n1511 );
    nor g31494 ( n33729 , n5335 , n10943 );
    and g31495 ( n10943 , n28054 , n30011 );
    or g31496 ( n20333 , n1950 , n6937 );
    not g31497 ( n6713 , n14381 );
    and g31498 ( n17390 , n9545 , n14923 );
    or g31499 ( n6671 , n35801 , n29366 );
    nor g31500 ( n2637 , n31215 , n7074 );
    or g31501 ( n9963 , n13600 , n4478 );
    and g31502 ( n2513 , n27033 , n7168 );
    or g31503 ( n19921 , n32670 , n35757 );
    nor g31504 ( n5210 , n6644 , n18115 );
    or g31505 ( n1080 , n18327 , n6370 );
    and g31506 ( n12586 , n31235 , n8213 );
    nor g31507 ( n14621 , n4758 , n35716 );
    or g31508 ( n34910 , n17208 , n2104 );
    or g31509 ( n24748 , n16583 , n3352 );
    or g31510 ( n18394 , n11455 , n22013 );
    or g31511 ( n10035 , n22296 , n18887 );
    or g31512 ( n9362 , n4837 , n16979 );
    nor g31513 ( n6121 , n4257 , n5495 );
    or g31514 ( n16719 , n244 , n26292 );
    not g31515 ( n14809 , n15142 );
    and g31516 ( n28917 , n21655 , n35952 );
    nor g31517 ( n16172 , n5804 , n19128 );
    or g31518 ( n19349 , n34983 , n30384 );
    or g31519 ( n35146 , n17389 , n18399 );
    and g31520 ( n12514 , n6902 , n20720 );
    xnor g31521 ( n2053 , n9535 , n25833 );
    xnor g31522 ( n22199 , n28011 , n33530 );
    and g31523 ( n22340 , n2267 , n15723 );
    or g31524 ( n5025 , n3029 , n4203 );
    or g31525 ( n17021 , n33897 , n15497 );
    not g31526 ( n12089 , n16594 );
    or g31527 ( n10543 , n25415 , n4478 );
    or g31528 ( n29260 , n34456 , n1901 );
    xnor g31529 ( n33223 , n33016 , n25896 );
    nor g31530 ( n429 , n7022 , n1187 );
    and g31531 ( n3346 , n13503 , n34730 );
    and g31532 ( n15474 , n9219 , n19037 );
    or g31533 ( n16187 , n4960 , n23102 );
    xnor g31534 ( n25943 , n30998 , n32095 );
    and g31535 ( n363 , n24392 , n25379 );
    and g31536 ( n17984 , n3393 , n607 );
    or g31537 ( n732 , n32584 , n13872 );
    or g31538 ( n25012 , n8823 , n14554 );
    and g31539 ( n524 , n25937 , n24494 );
    and g31540 ( n11245 , n3198 , n33577 );
    or g31541 ( n896 , n25312 , n11703 );
    or g31542 ( n5142 , n14363 , n20812 );
    xnor g31543 ( n11595 , n35552 , n4417 );
    or g31544 ( n16123 , n32389 , n8882 );
    or g31545 ( n5000 , n33189 , n12996 );
    xnor g31546 ( n5667 , n16857 , n28219 );
    not g31547 ( n25883 , n12213 );
    or g31548 ( n11566 , n9789 , n17359 );
    and g31549 ( n16399 , n2804 , n1112 );
    or g31550 ( n26088 , n21536 , n25583 );
    or g31551 ( n30303 , n34062 , n19306 );
    or g31552 ( n20999 , n8662 , n15266 );
    nor g31553 ( n22564 , n35927 , n14912 );
    or g31554 ( n5861 , n35493 , n8366 );
    xnor g31555 ( n13779 , n825 , n12758 );
    xnor g31556 ( n5919 , n3212 , n16843 );
    and g31557 ( n26474 , n22143 , n14822 );
    or g31558 ( n314 , n14201 , n28995 );
    or g31559 ( n13842 , n34708 , n34971 );
    or g31560 ( n1209 , n12133 , n13480 );
    and g31561 ( n3730 , n28697 , n12690 );
    xnor g31562 ( n5520 , n31558 , n22291 );
    and g31563 ( n7104 , n9835 , n20394 );
    and g31564 ( n30033 , n28094 , n5332 );
    or g31565 ( n33717 , n25415 , n24271 );
    or g31566 ( n23637 , n25104 , n30646 );
    and g31567 ( n18855 , n8811 , n17023 );
    not g31568 ( n34027 , n210 );
    or g31569 ( n412 , n4962 , n8914 );
    or g31570 ( n2870 , n31799 , n35951 );
    not g31571 ( n8412 , n19952 );
    or g31572 ( n29074 , n22937 , n8312 );
    xnor g31573 ( n23018 , n27897 , n32095 );
    and g31574 ( n7568 , n13199 , n30834 );
    and g31575 ( n12984 , n157 , n33527 );
    and g31576 ( n25530 , n21637 , n13793 );
    nor g31577 ( n1688 , n12062 , n17758 );
    and g31578 ( n18371 , n22085 , n21975 );
    xnor g31579 ( n31879 , n34812 , n7364 );
    xnor g31580 ( n28956 , n17189 , n35631 );
    nor g31581 ( n18032 , n14182 , n2556 );
    not g31582 ( n32054 , n34094 );
    nor g31583 ( n1392 , n1979 , n19834 );
    xnor g31584 ( n24334 , n17249 , n24371 );
    and g31585 ( n8834 , n9400 , n26853 );
    xnor g31586 ( n9359 , n32101 , n9789 );
    or g31587 ( n35298 , n26154 , n20690 );
    or g31588 ( n14876 , n29822 , n29411 );
    xnor g31589 ( n29069 , n30199 , n29527 );
    or g31590 ( n19958 , n6334 , n18811 );
    or g31591 ( n2567 , n27254 , n35748 );
    and g31592 ( n16715 , n21446 , n20857 );
    and g31593 ( n33632 , n22880 , n16138 );
    xnor g31594 ( n30375 , n10369 , n8259 );
    or g31595 ( n22551 , n209 , n24587 );
    xnor g31596 ( n23235 , n16857 , n26608 );
    nor g31597 ( n304 , n14082 , n32379 );
    xnor g31598 ( n29670 , n13372 , n7422 );
    or g31599 ( n332 , n10820 , n35174 );
    and g31600 ( n19089 , n33216 , n26955 );
    or g31601 ( n2655 , n12172 , n763 );
    or g31602 ( n33682 , n31584 , n8203 );
    or g31603 ( n30083 , n9109 , n21902 );
    or g31604 ( n2504 , n4654 , n9030 );
    or g31605 ( n26305 , n8155 , n34397 );
    or g31606 ( n11581 , n11506 , n17612 );
    or g31607 ( n6932 , n34759 , n6340 );
    or g31608 ( n32372 , n5020 , n26931 );
    nor g31609 ( n7205 , n17621 , n18484 );
    or g31610 ( n21741 , n3315 , n28837 );
    or g31611 ( n18218 , n10894 , n7447 );
    or g31612 ( n1363 , n27353 , n27447 );
    nor g31613 ( n28203 , n4960 , n11575 );
    xnor g31614 ( n6291 , n5316 , n29156 );
    and g31615 ( n9428 , n30864 , n13671 );
    or g31616 ( n11185 , n22763 , n707 );
    buf g31617 ( n7673 , n32572 );
    or g31618 ( n22537 , n27865 , n20427 );
    or g31619 ( n26164 , n16044 , n1755 );
    or g31620 ( n8581 , n19551 , n23030 );
    xnor g31621 ( n17063 , n35108 , n3205 );
    and g31622 ( n20072 , n7401 , n22191 );
    or g31623 ( n2547 , n20901 , n13075 );
    nor g31624 ( n10346 , n3222 , n7835 );
    or g31625 ( n2720 , n2075 , n14726 );
    nor g31626 ( n7644 , n19010 , n22007 );
    nor g31627 ( n15265 , n34551 , n20758 );
    and g31628 ( n31619 , n24493 , n32228 );
    xnor g31629 ( n17076 , n30921 , n18171 );
    or g31630 ( n8386 , n18979 , n5220 );
    xnor g31631 ( n33480 , n25118 , n1564 );
    xnor g31632 ( n31406 , n14832 , n21370 );
    and g31633 ( n7192 , n32980 , n3234 );
    and g31634 ( n29782 , n22378 , n29845 );
    xnor g31635 ( n26254 , n4999 , n22077 );
    not g31636 ( n12206 , n8865 );
    xnor g31637 ( n10802 , n27582 , n29713 );
    or g31638 ( n24456 , n21014 , n13909 );
    or g31639 ( n5992 , n5466 , n11258 );
    or g31640 ( n18517 , n12360 , n8954 );
    or g31641 ( n24907 , n10149 , n19845 );
    or g31642 ( n8569 , n424 , n29626 );
    and g31643 ( n17314 , n1789 , n18496 );
    or g31644 ( n5097 , n28048 , n33750 );
    or g31645 ( n23240 , n23604 , n20651 );
    xnor g31646 ( n27082 , n16836 , n19933 );
    and g31647 ( n21361 , n28771 , n701 );
    and g31648 ( n33053 , n1530 , n400 );
    or g31649 ( n2415 , n6322 , n9448 );
    xnor g31650 ( n10405 , n2477 , n25174 );
    xnor g31651 ( n11667 , n12267 , n21653 );
    not g31652 ( n35609 , n3805 );
    xnor g31653 ( n34259 , n5593 , n35794 );
    not g31654 ( n8163 , n11960 );
    nor g31655 ( n7960 , n29177 , n3132 );
    xnor g31656 ( n14323 , n5892 , n13931 );
    nor g31657 ( n29226 , n5738 , n26656 );
    or g31658 ( n13934 , n7569 , n9989 );
    or g31659 ( n28880 , n4962 , n25514 );
    nor g31660 ( n29517 , n830 , n6714 );
    xnor g31661 ( n6386 , n4280 , n21585 );
    or g31662 ( n15902 , n35584 , n908 );
    or g31663 ( n26848 , n7432 , n12857 );
    not g31664 ( n11599 , n16620 );
    or g31665 ( n35502 , n32857 , n3178 );
    and g31666 ( n10572 , n17970 , n34751 );
    and g31667 ( n19210 , n29215 , n19339 );
    nor g31668 ( n4924 , n29713 , n23241 );
    xnor g31669 ( n32154 , n8343 , n2458 );
    or g31670 ( n7655 , n32559 , n20797 );
    and g31671 ( n23804 , n13183 , n30810 );
    not g31672 ( n28536 , n16922 );
    xnor g31673 ( n7772 , n32319 , n19625 );
    and g31674 ( n35928 , n9660 , n24288 );
    xnor g31675 ( n19504 , n9687 , n29438 );
    xnor g31676 ( n689 , n6184 , n20278 );
    nor g31677 ( n24046 , n20856 , n19834 );
    or g31678 ( n29019 , n11652 , n1796 );
    xnor g31679 ( n13647 , n25679 , n16620 );
    and g31680 ( n20465 , n18589 , n35487 );
    xnor g31681 ( n15558 , n24759 , n16922 );
    or g31682 ( n28847 , n23604 , n14744 );
    or g31683 ( n17047 , n24892 , n19845 );
    buf g31684 ( n24710 , n12956 );
    and g31685 ( n4379 , n33564 , n24092 );
    xnor g31686 ( n31525 , n9190 , n15464 );
    and g31687 ( n15717 , n22557 , n32643 );
    xnor g31688 ( n12485 , n11448 , n8075 );
    and g31689 ( n2700 , n6740 , n1727 );
    xnor g31690 ( n22513 , n3603 , n34807 );
    or g31691 ( n27170 , n2841 , n28240 );
    nor g31692 ( n5616 , n12235 , n35591 );
    xnor g31693 ( n31475 , n33887 , n10894 );
    and g31694 ( n18490 , n15221 , n13042 );
    xnor g31695 ( n30817 , n20882 , n32116 );
    or g31696 ( n29762 , n22334 , n19058 );
    not g31697 ( n16414 , n2630 );
    or g31698 ( n2480 , n14773 , n23790 );
    or g31699 ( n18154 , n15720 , n7230 );
    or g31700 ( n11476 , n18377 , n33677 );
    and g31701 ( n9398 , n26274 , n18339 );
    and g31702 ( n23233 , n35683 , n15948 );
    nor g31703 ( n2209 , n9789 , n22177 );
    xnor g31704 ( n35994 , n27874 , n25657 );
    and g31705 ( n21386 , n19007 , n19092 );
    and g31706 ( n9937 , n25716 , n24671 );
    xnor g31707 ( n13375 , n19368 , n29884 );
    xnor g31708 ( n32918 , n32921 , n32703 );
    and g31709 ( n4468 , n7330 , n22849 );
    and g31710 ( n14744 , n8874 , n1977 );
    or g31711 ( n21718 , n20786 , n10736 );
    xnor g31712 ( n29116 , n29546 , n14770 );
    or g31713 ( n27976 , n15464 , n7209 );
    xnor g31714 ( n8340 , n26843 , n33829 );
    or g31715 ( n27458 , n16620 , n6269 );
    and g31716 ( n11743 , n10045 , n227 );
    or g31717 ( n17176 , n1950 , n13287 );
    xnor g31718 ( n19880 , n26693 , n3205 );
    or g31719 ( n9886 , n31289 , n20768 );
    or g31720 ( n8768 , n10954 , n31403 );
    and g31721 ( n13567 , n4343 , n888 );
    or g31722 ( n30111 , n29956 , n35928 );
    or g31723 ( n27446 , n19712 , n3704 );
    xnor g31724 ( n34754 , n7499 , n11985 );
    xnor g31725 ( n14082 , n7981 , n6666 );
    or g31726 ( n6224 , n13205 , n35757 );
    or g31727 ( n21658 , n12546 , n31301 );
    or g31728 ( n6813 , n4878 , n4449 );
    or g31729 ( n18008 , n33944 , n23601 );
    and g31730 ( n29628 , n13916 , n7736 );
    or g31731 ( n9322 , n28920 , n1730 );
    nor g31732 ( n15989 , n32945 , n19834 );
    and g31733 ( n13560 , n4760 , n20520 );
    or g31734 ( n14713 , n26772 , n23605 );
    or g31735 ( n25258 , n3222 , n17151 );
    not g31736 ( n4209 , n17842 );
    buf g31737 ( n16762 , n20749 );
    and g31738 ( n29384 , n8073 , n29319 );
    xnor g31739 ( n18631 , n2674 , n23414 );
    and g31740 ( n20025 , n34703 , n21940 );
    and g31741 ( n29868 , n28018 , n14135 );
    or g31742 ( n16662 , n19982 , n20305 );
    not g31743 ( n20354 , n32857 );
    xnor g31744 ( n22337 , n771 , n11455 );
    or g31745 ( n17015 , n31289 , n10213 );
    xnor g31746 ( n19256 , n29278 , n31559 );
    or g31747 ( n1988 , n2170 , n14170 );
    and g31748 ( n26464 , n12718 , n3849 );
    or g31749 ( n5285 , n20823 , n19643 );
    or g31750 ( n10103 , n24468 , n27447 );
    and g31751 ( n20068 , n4486 , n33100 );
    xnor g31752 ( n27567 , n21830 , n27887 );
    xnor g31753 ( n34790 , n29952 , n27145 );
    or g31754 ( n8208 , n30136 , n7962 );
    not g31755 ( n13085 , n2875 );
    and g31756 ( n9467 , n27221 , n18869 );
    or g31757 ( n29085 , n20833 , n20817 );
    and g31758 ( n16377 , n34573 , n15200 );
    or g31759 ( n10116 , n35892 , n21579 );
    nor g31760 ( n28848 , n24371 , n22829 );
    nor g31761 ( n1675 , n14376 , n12103 );
    and g31762 ( n19474 , n8392 , n21039 );
    nor g31763 ( n17375 , n32584 , n16633 );
    or g31764 ( n3302 , n33019 , n36000 );
    or g31765 ( n15938 , n24371 , n16377 );
    xnor g31766 ( n19599 , n656 , n21318 );
    or g31767 ( n29416 , n16696 , n30700 );
    and g31768 ( n22859 , n5508 , n12190 );
    xnor g31769 ( n16176 , n1576 , n29713 );
    xnor g31770 ( n33127 , n31748 , n8477 );
    not g31771 ( n11974 , n4878 );
    xnor g31772 ( n6359 , n5408 , n3882 );
    xnor g31773 ( n42 , n17082 , n446 );
    or g31774 ( n7107 , n22074 , n22961 );
    or g31775 ( n25254 , n22354 , n19952 );
    or g31776 ( n26331 , n24332 , n6415 );
    or g31777 ( n35779 , n26849 , n19336 );
    nor g31778 ( n8155 , n19551 , n22264 );
    xnor g31779 ( n31322 , n13877 , n4878 );
    not g31780 ( n5424 , n22980 );
    and g31781 ( n4357 , n7276 , n9751 );
    or g31782 ( n29498 , n32335 , n24653 );
    xnor g31783 ( n15048 , n22505 , n25602 );
    nor g31784 ( n9477 , n9793 , n23420 );
    and g31785 ( n27746 , n29813 , n10980 );
    nor g31786 ( n16564 , n14807 , n7448 );
    or g31787 ( n35207 , n14907 , n22858 );
    xnor g31788 ( n737 , n13889 , n18711 );
    or g31789 ( n8908 , n14042 , n24004 );
    or g31790 ( n12260 , n28834 , n15144 );
    or g31791 ( n34188 , n17228 , n23921 );
    xnor g31792 ( n21709 , n13163 , n709 );
    or g31793 ( n14925 , n13445 , n23801 );
    or g31794 ( n15488 , n25055 , n29953 );
    not g31795 ( n34876 , n34503 );
    xnor g31796 ( n26158 , n26125 , n4878 );
    not g31797 ( n16056 , n33650 );
    not g31798 ( n7434 , n36045 );
    not g31799 ( n25539 , n24304 );
    xnor g31800 ( n30286 , n13660 , n10914 );
    not g31801 ( n20447 , n11838 );
    or g31802 ( n13589 , n1515 , n24653 );
    or g31803 ( n25467 , n27211 , n19058 );
    xnor g31804 ( n30899 , n27107 , n24730 );
    xnor g31805 ( n4457 , n22453 , n27619 );
    or g31806 ( n2021 , n13186 , n35111 );
    and g31807 ( n27827 , n1367 , n24708 );
    and g31808 ( n4587 , n9307 , n12825 );
    or g31809 ( n6222 , n18162 , n26023 );
    xnor g31810 ( n7149 , n19923 , n492 );
    or g31811 ( n27523 , n204 , n1414 );
    or g31812 ( n27938 , n22291 , n5299 );
    or g31813 ( n24232 , n2697 , n29562 );
    or g31814 ( n22576 , n32887 , n8271 );
    xnor g31815 ( n32541 , n20904 , n20022 );
    not g31816 ( n32422 , n31431 );
    and g31817 ( n21404 , n22893 , n25535 );
    or g31818 ( n387 , n14345 , n9953 );
    or g31819 ( n12543 , n10894 , n4072 );
    and g31820 ( n5588 , n12525 , n14338 );
    or g31821 ( n278 , n27249 , n22572 );
    or g31822 ( n8980 , n29923 , n4330 );
    and g31823 ( n5089 , n30257 , n21756 );
    or g31824 ( n18142 , n13854 , n35141 );
    not g31825 ( n20136 , n6658 );
    or g31826 ( n3871 , n15715 , n1061 );
    or g31827 ( n14263 , n5733 , n2820 );
    and g31828 ( n5830 , n12896 , n15395 );
    and g31829 ( n35392 , n2220 , n1208 );
    not g31830 ( n30734 , n28322 );
    not g31831 ( n35036 , n25547 );
    xnor g31832 ( n8359 , n6551 , n6677 );
    not g31833 ( n3314 , n18174 );
    or g31834 ( n1766 , n16804 , n16326 );
    or g31835 ( n16227 , n21286 , n33400 );
    or g31836 ( n30017 , n27231 , n23748 );
    xor g31837 ( n2106 , n5362 , n6372 );
    or g31838 ( n33106 , n11626 , n4929 );
    xnor g31839 ( n35989 , n28039 , n32909 );
    nor g31840 ( n27600 , n22255 , n20467 );
    nor g31841 ( n8774 , n830 , n20173 );
    nor g31842 ( n25137 , n16620 , n18271 );
    xnor g31843 ( n26888 , n11281 , n28660 );
    or g31844 ( n19455 , n417 , n17025 );
    xnor g31845 ( n1990 , n33777 , n6118 );
    and g31846 ( n18667 , n15632 , n35096 );
    or g31847 ( n1881 , n6645 , n17162 );
    nor g31848 ( n12025 , n16620 , n26335 );
    or g31849 ( n26954 , n34499 , n33098 );
    buf g31850 ( n18264 , n20798 );
    nor g31851 ( n4940 , n23604 , n34516 );
    or g31852 ( n18223 , n8960 , n21999 );
    not g31853 ( n14775 , n22980 );
    xnor g31854 ( n14782 , n35931 , n31799 );
    xnor g31855 ( n32663 , n14718 , n31289 );
    or g31856 ( n24103 , n16798 , n19919 );
    not g31857 ( n32968 , n1950 );
    xnor g31858 ( n10785 , n1601 , n8909 );
    or g31859 ( n32460 , n19528 , n14554 );
    or g31860 ( n20296 , n3222 , n35089 );
    and g31861 ( n20120 , n24268 , n16274 );
    or g31862 ( n24335 , n6980 , n20797 );
    and g31863 ( n24781 , n5651 , n29345 );
    or g31864 ( n3195 , n33843 , n18634 );
    and g31865 ( n29487 , n22773 , n1224 );
    xnor g31866 ( n25129 , n6870 , n6278 );
    or g31867 ( n21263 , n31056 , n33880 );
    or g31868 ( n18840 , n11470 , n25255 );
    xnor g31869 ( n17086 , n17487 , n31289 );
    or g31870 ( n12074 , n13126 , n17612 );
    or g31871 ( n20319 , n4878 , n20426 );
    or g31872 ( n31278 , n12925 , n1511 );
    xnor g31873 ( n2941 , n12171 , n10894 );
    or g31874 ( n35646 , n24450 , n19173 );
    and g31875 ( n8064 , n32134 , n30493 );
    xnor g31876 ( n14927 , n31508 , n4337 );
    and g31877 ( n21569 , n30571 , n31019 );
    or g31878 ( n20011 , n32466 , n23209 );
    or g31879 ( n21402 , n9658 , n18374 );
    or g31880 ( n9041 , n13386 , n11850 );
    not g31881 ( n14672 , n7588 );
    and g31882 ( n17202 , n28322 , n30048 );
    not g31883 ( n23297 , n23085 );
    buf g31884 ( n17125 , n18698 );
    not g31885 ( n6999 , n27291 );
    not g31886 ( n12926 , n23078 );
    xnor g31887 ( n14217 , n26703 , n1950 );
    or g31888 ( n17387 , n3222 , n2992 );
    or g31889 ( n5599 , n23551 , n8704 );
    not g31890 ( n22678 , n35859 );
    or g31891 ( n3347 , n2764 , n21731 );
    and g31892 ( n1652 , n19017 , n34485 );
    xnor g31893 ( n685 , n12078 , n13335 );
    nor g31894 ( n32077 , n34967 , n29366 );
    or g31895 ( n15421 , n25174 , n14059 );
    xnor g31896 ( n7235 , n31715 , n29884 );
    or g31897 ( n18476 , n28776 , n26023 );
    xnor g31898 ( n30059 , n29736 , n21332 );
    and g31899 ( n32517 , n2874 , n13253 );
    or g31900 ( n14928 , n30820 , n14746 );
    not g31901 ( n32983 , n13547 );
    or g31902 ( n2165 , n25216 , n6288 );
    and g31903 ( n28684 , n14347 , n7290 );
    xnor g31904 ( n23210 , n11322 , n9412 );
    and g31905 ( n22030 , n13506 , n8208 );
    not g31906 ( n20190 , n24623 );
    or g31907 ( n34669 , n3205 , n26049 );
    not g31908 ( n19848 , n27213 );
    or g31909 ( n3139 , n24275 , n26292 );
    xnor g31910 ( n31895 , n5093 , n22291 );
    or g31911 ( n12985 , n2758 , n31032 );
    xnor g31912 ( n5360 , n8624 , n19551 );
    xnor g31913 ( n25954 , n34737 , n23604 );
    and g31914 ( n27623 , n30178 , n5506 );
    or g31915 ( n24752 , n6715 , n14033 );
    and g31916 ( n20511 , n24935 , n24250 );
    and g31917 ( n28088 , n25348 , n25352 );
    and g31918 ( n20463 , n13150 , n24075 );
    or g31919 ( n6997 , n9789 , n4213 );
    or g31920 ( n22933 , n797 , n35216 );
    or g31921 ( n21541 , n21108 , n28240 );
    xnor g31922 ( n32433 , n498 , n30742 );
    xnor g31923 ( n29776 , n20604 , n16922 );
    xnor g31924 ( n15081 , n1113 , n3205 );
    or g31925 ( n15909 , n28228 , n33039 );
    or g31926 ( n33356 , n10398 , n16797 );
    and g31927 ( n2176 , n25622 , n7120 );
    or g31928 ( n21597 , n22008 , n12596 );
    xnor g31929 ( n26396 , n15170 , n22291 );
    or g31930 ( n24353 , n33986 , n31482 );
    and g31931 ( n2932 , n32592 , n27555 );
    or g31932 ( n9485 , n2462 , n7417 );
    or g31933 ( n29634 , n34899 , n25526 );
    or g31934 ( n17342 , n30049 , n31606 );
    or g31935 ( n5971 , n29382 , n15439 );
    or g31936 ( n1868 , n14284 , n10432 );
    or g31937 ( n4293 , n15735 , n25648 );
    and g31938 ( n27060 , n6892 , n24733 );
    or g31939 ( n29638 , n24859 , n20964 );
    xnor g31940 ( n9476 , n11320 , n34968 );
    or g31941 ( n26324 , n25523 , n28969 );
    or g31942 ( n3268 , n6034 , n19490 );
    or g31943 ( n17213 , n14600 , n9147 );
    and g31944 ( n8857 , n22342 , n34393 );
    or g31945 ( n30358 , n13677 , n2104 );
    and g31946 ( n18260 , n12313 , n23702 );
    not g31947 ( n35812 , n2889 );
    and g31948 ( n16621 , n26196 , n21877 );
    xnor g31949 ( n17457 , n5187 , n29713 );
    or g31950 ( n2474 , n32857 , n4258 );
    or g31951 ( n30647 , n12329 , n12763 );
    or g31952 ( n13354 , n2175 , n26192 );
    and g31953 ( n6528 , n1271 , n25892 );
    or g31954 ( n4358 , n32095 , n34590 );
    or g31955 ( n4549 , n8660 , n8153 );
    xnor g31956 ( n26573 , n4717 , n24829 );
    not g31957 ( n7557 , n3873 );
    or g31958 ( n23243 , n32250 , n28866 );
    nor g31959 ( n16796 , n16093 , n33956 );
    xnor g31960 ( n27298 , n3930 , n24826 );
    and g31961 ( n18651 , n9685 , n5294 );
    or g31962 ( n12187 , n5360 , n32716 );
    not g31963 ( n31205 , n29378 );
    or g31964 ( n22515 , n4988 , n7359 );
    or g31965 ( n10448 , n2361 , n4595 );
    and g31966 ( n30401 , n13917 , n32429 );
    xnor g31967 ( n22620 , n1872 , n31635 );
    xnor g31968 ( n10753 , n23115 , n7087 );
    not g31969 ( n27764 , n9427 );
    or g31970 ( n16890 , n5502 , n4478 );
    and g31971 ( n20364 , n32984 , n34243 );
    xnor g31972 ( n17495 , n7799 , n5121 );
    or g31973 ( n15748 , n17339 , n20812 );
    or g31974 ( n29307 , n24506 , n26480 );
    and g31975 ( n4540 , n137 , n24209 );
    nor g31976 ( n8877 , n34606 , n24673 );
    xnor g31977 ( n24964 , n29575 , n1810 );
    xnor g31978 ( n30727 , n17132 , n29447 );
    or g31979 ( n8825 , n33559 , n21042 );
    or g31980 ( n22493 , n33093 , n26112 );
    or g31981 ( n34870 , n13154 , n12340 );
    or g31982 ( n2406 , n23850 , n32425 );
    or g31983 ( n34095 , n21064 , n16473 );
    or g31984 ( n22423 , n31559 , n31039 );
    and g31985 ( n32822 , n2371 , n7791 );
    or g31986 ( n9774 , n20245 , n27580 );
    xnor g31987 ( n22317 , n6579 , n3946 );
    or g31988 ( n14155 , n3143 , n15256 );
    and g31989 ( n19244 , n26425 , n22145 );
    or g31990 ( n15487 , n17141 , n20601 );
    xnor g31991 ( n28814 , n26256 , n14410 );
    or g31992 ( n4248 , n20130 , n19403 );
    not g31993 ( n24851 , n915 );
    and g31994 ( n6124 , n2935 , n25462 );
    and g31995 ( n23418 , n18859 , n28928 );
    or g31996 ( n14235 , n24919 , n23626 );
    and g31997 ( n21297 , n7655 , n32413 );
    or g31998 ( n24268 , n16158 , n2360 );
    buf g31999 ( n26468 , n35410 );
    xnor g32000 ( n7968 , n12809 , n26174 );
    and g32001 ( n12809 , n15174 , n26721 );
    xnor g32002 ( n31976 , n2729 , n32584 );
    or g32003 ( n20390 , n13175 , n17068 );
    or g32004 ( n23649 , n3205 , n8358 );
    or g32005 ( n6330 , n30553 , n11648 );
    or g32006 ( n22635 , n4878 , n15804 );
    xnor g32007 ( n23120 , n25783 , n16135 );
    xnor g32008 ( n13557 , n15535 , n19614 );
    xnor g32009 ( n26038 , n25987 , n15464 );
    or g32010 ( n25626 , n27226 , n32841 );
    or g32011 ( n222 , n7666 , n2384 );
    or g32012 ( n28150 , n4288 , n30425 );
    and g32013 ( n35369 , n2529 , n31158 );
    or g32014 ( n25860 , n12729 , n15805 );
    or g32015 ( n26079 , n17568 , n20389 );
    buf g32016 ( n22501 , n26426 );
    or g32017 ( n15848 , n18379 , n15463 );
    or g32018 ( n6102 , n12494 , n25773 );
    and g32019 ( n733 , n6068 , n5693 );
    or g32020 ( n10755 , n31402 , n22945 );
    and g32021 ( n24811 , n34675 , n29428 );
    not g32022 ( n20024 , n1202 );
    and g32023 ( n10800 , n34326 , n28730 );
    xnor g32024 ( n6581 , n22947 , n32857 );
    xnor g32025 ( n4419 , n12150 , n30697 );
    or g32026 ( n22231 , n31040 , n34902 );
    and g32027 ( n10849 , n3659 , n15293 );
    or g32028 ( n4656 , n16018 , n19952 );
    not g32029 ( n9571 , n26153 );
    xnor g32030 ( n24421 , n16330 , n35927 );
    or g32031 ( n3969 , n23711 , n29626 );
    and g32032 ( n16409 , n11345 , n15880 );
    and g32033 ( n19452 , n650 , n20386 );
    xnor g32034 ( n22223 , n32778 , n7540 );
    and g32035 ( n18037 , n34931 , n25646 );
    xnor g32036 ( n14320 , n31412 , n4962 );
    or g32037 ( n32601 , n29272 , n24351 );
    xnor g32038 ( n22242 , n24298 , n3395 );
    or g32039 ( n27970 , n7663 , n33799 );
    or g32040 ( n2974 , n35722 , n5868 );
    and g32041 ( n19909 , n29299 , n21067 );
    xnor g32042 ( n33538 , n13287 , n1950 );
    buf g32043 ( n32425 , n34923 );
    xnor g32044 ( n6516 , n17022 , n14436 );
    or g32045 ( n24637 , n32584 , n7775 );
    xnor g32046 ( n32953 , n31702 , n25602 );
    nor g32047 ( n15165 , n15464 , n32682 );
    or g32048 ( n26248 , n28200 , n24841 );
    not g32049 ( n15919 , n10183 );
    not g32050 ( n27433 , n10009 );
    buf g32051 ( n15538 , n17793 );
    buf g32052 ( n21210 , n34458 );
    and g32053 ( n15878 , n16082 , n31095 );
    or g32054 ( n10527 , n8640 , n12268 );
    nor g32055 ( n9207 , n25426 , n24746 );
    xnor g32056 ( n11533 , n7708 , n32095 );
    and g32057 ( n19881 , n7494 , n2069 );
    or g32058 ( n23582 , n17054 , n4254 );
    or g32059 ( n1166 , n29903 , n14697 );
    and g32060 ( n29527 , n32555 , n21864 );
    xnor g32061 ( n8902 , n19328 , n21282 );
    and g32062 ( n24156 , n29294 , n31339 );
    or g32063 ( n32884 , n24371 , n25608 );
    nor g32064 ( n27075 , n21285 , n14507 );
    and g32065 ( n15197 , n18117 , n21718 );
    not g32066 ( n18393 , n31799 );
    nor g32067 ( n11676 , n17394 , n16112 );
    xnor g32068 ( n16906 , n13234 , n31727 );
    or g32069 ( n16839 , n23883 , n13480 );
    and g32070 ( n27405 , n28970 , n10258 );
    buf g32071 ( n1402 , n26110 );
    nor g32072 ( n13517 , n16620 , n9352 );
    or g32073 ( n2278 , n6629 , n19084 );
    or g32074 ( n27786 , n7051 , n17616 );
    xnor g32075 ( n11839 , n29570 , n830 );
    xnor g32076 ( n8227 , n18983 , n3989 );
    and g32077 ( n27046 , n36056 , n2321 );
    or g32078 ( n32852 , n27820 , n10400 );
    or g32079 ( n30986 , n28376 , n20954 );
    not g32080 ( n5124 , n28866 );
    or g32081 ( n32399 , n9655 , n2119 );
    xnor g32082 ( n28509 , n5242 , n4758 );
    and g32083 ( n703 , n14937 , n1816 );
    xnor g32084 ( n32119 , n26005 , n479 );
    xnor g32085 ( n35878 , n19425 , n19551 );
    or g32086 ( n2255 , n35327 , n34537 );
    xnor g32087 ( n15999 , n26330 , n2440 );
    or g32088 ( n3764 , n21062 , n27801 );
    and g32089 ( n13000 , n5434 , n34177 );
    or g32090 ( n27360 , n7939 , n10683 );
    or g32091 ( n1951 , n25908 , n2256 );
    or g32092 ( n6874 , n19741 , n1557 );
    and g32093 ( n17664 , n1710 , n5785 );
    or g32094 ( n17192 , n30218 , n9832 );
    or g32095 ( n21969 , n29699 , n6683 );
    and g32096 ( n2360 , n4680 , n29751 );
    xnor g32097 ( n29960 , n30096 , n16444 );
    or g32098 ( n25427 , n8118 , n26292 );
    or g32099 ( n9487 , n25808 , n17612 );
    not g32100 ( n3125 , n15403 );
    xnor g32101 ( n28598 , n30228 , n29288 );
    or g32102 ( n28369 , n32715 , n13714 );
    or g32103 ( n17900 , n31349 , n24489 );
    or g32104 ( n17216 , n11018 , n19260 );
    or g32105 ( n33749 , n20539 , n6950 );
    and g32106 ( n28659 , n22890 , n13626 );
    or g32107 ( n26544 , n20403 , n34484 );
    and g32108 ( n34977 , n21682 , n26880 );
    or g32109 ( n13027 , n10935 , n11464 );
    nor g32110 ( n30635 , n3557 , n9921 );
    xnor g32111 ( n21052 , n21171 , n29847 );
    xnor g32112 ( n4987 , n16275 , n23421 );
    or g32113 ( n25305 , n18271 , n20318 );
    xnor g32114 ( n7073 , n25238 , n32362 );
    or g32115 ( n28540 , n18110 , n9082 );
    and g32116 ( n19666 , n35016 , n28333 );
    xnor g32117 ( n245 , n30648 , n1168 );
    nor g32118 ( n32019 , n16620 , n20411 );
    and g32119 ( n35128 , n31728 , n6888 );
    and g32120 ( n10714 , n25339 , n24255 );
    not g32121 ( n20041 , n26098 );
    xnor g32122 ( n15062 , n13580 , n2661 );
    or g32123 ( n6160 , n28482 , n23390 );
    xnor g32124 ( n7560 , n7745 , n22291 );
    not g32125 ( n35393 , n18121 );
    or g32126 ( n30052 , n25425 , n4188 );
    or g32127 ( n29591 , n1340 , n4772 );
    xnor g32128 ( n28707 , n8313 , n10894 );
    xnor g32129 ( n1339 , n15409 , n5358 );
    and g32130 ( n29267 , n22712 , n4224 );
    or g32131 ( n14052 , n10492 , n16344 );
    or g32132 ( n32710 , n7809 , n17183 );
    or g32133 ( n24188 , n27385 , n10417 );
    xnor g32134 ( n32103 , n25118 , n29622 );
    and g32135 ( n11801 , n17787 , n25169 );
    xnor g32136 ( n7023 , n5684 , n31056 );
    and g32137 ( n30367 , n24711 , n31770 );
    and g32138 ( n30179 , n19114 , n5031 );
    not g32139 ( n5837 , n3205 );
    or g32140 ( n24003 , n26151 , n10276 );
    xnor g32141 ( n16508 , n33326 , n23604 );
    or g32142 ( n15613 , n31956 , n19999 );
    not g32143 ( n5077 , n6344 );
    not g32144 ( n19258 , n33172 );
    or g32145 ( n25348 , n20921 , n19036 );
    or g32146 ( n9264 , n19551 , n14696 );
    not g32147 ( n30973 , n27099 );
    or g32148 ( n33510 , n13368 , n34865 );
    and g32149 ( n11091 , n26451 , n34124 );
    xnor g32150 ( n18883 , n18160 , n2960 );
    nor g32151 ( n10612 , n25018 , n33859 );
    or g32152 ( n34335 , n4878 , n12601 );
    or g32153 ( n34638 , n7023 , n1021 );
    and g32154 ( n21465 , n17062 , n30706 );
    xnor g32155 ( n11999 , n12946 , n30044 );
    or g32156 ( n13876 , n35639 , n4952 );
    nor g32157 ( n12603 , n25174 , n34650 );
    nor g32158 ( n30954 , n13413 , n16896 );
    or g32159 ( n11405 , n8635 , n6553 );
    and g32160 ( n7102 , n6668 , n12699 );
    or g32161 ( n8182 , n16426 , n17257 );
    and g32162 ( n32929 , n32377 , n22884 );
    xnor g32163 ( n20435 , n6183 , n3946 );
    or g32164 ( n5540 , n11257 , n32917 );
    nor g32165 ( n28836 , n34850 , n16736 );
    xnor g32166 ( n6872 , n27158 , n19551 );
    and g32167 ( n35332 , n23246 , n7505 );
    or g32168 ( n32094 , n26843 , n33829 );
    or g32169 ( n17795 , n18883 , n5618 );
    or g32170 ( n7522 , n13513 , n9024 );
    xnor g32171 ( n20332 , n26687 , n4962 );
    nor g32172 ( n12082 , n35140 , n5537 );
    or g32173 ( n29729 , n4962 , n28593 );
    or g32174 ( n2872 , n11042 , n10417 );
    and g32175 ( n27710 , n13404 , n29308 );
    or g32176 ( n31818 , n18661 , n4912 );
    not g32177 ( n15967 , n4595 );
    or g32178 ( n23356 , n28546 , n5252 );
    or g32179 ( n29211 , n24371 , n5723 );
    nor g32180 ( n21064 , n4288 , n9792 );
    or g32181 ( n22894 , n1357 , n28191 );
    and g32182 ( n24560 , n30447 , n33208 );
    and g32183 ( n28242 , n9007 , n20916 );
    or g32184 ( n4622 , n31056 , n2753 );
    and g32185 ( n28099 , n16096 , n35382 );
    nor g32186 ( n31923 , n26584 , n11161 );
    and g32187 ( n34618 , n8194 , n2466 );
    xnor g32188 ( n11324 , n7347 , n32715 );
    or g32189 ( n629 , n16620 , n18802 );
    or g32190 ( n18611 , n16620 , n32568 );
    or g32191 ( n21746 , n29053 , n32176 );
    nor g32192 ( n12429 , n15886 , n7301 );
    not g32193 ( n8648 , n25761 );
    buf g32194 ( n17233 , n11127 );
    and g32195 ( n12118 , n4512 , n7378 );
    xnor g32196 ( n9490 , n13731 , n24371 );
    or g32197 ( n31489 , n6660 , n8648 );
    xnor g32198 ( n6185 , n11590 , n7913 );
    and g32199 ( n4204 , n18800 , n24321 );
    or g32200 ( n21580 , n4288 , n19210 );
    xnor g32201 ( n3311 , n11644 , n3205 );
    xnor g32202 ( n21096 , n17300 , n3205 );
    xnor g32203 ( n27955 , n16158 , n2360 );
    or g32204 ( n3354 , n5766 , n24696 );
    or g32205 ( n5531 , n34475 , n29461 );
    or g32206 ( n26491 , n31863 , n22206 );
    nor g32207 ( n13316 , n4273 , n6548 );
    not g32208 ( n3680 , n2092 );
    not g32209 ( n17232 , n26801 );
    or g32210 ( n8522 , n27111 , n22084 );
    or g32211 ( n20625 , n17592 , n33086 );
    nor g32212 ( n18834 , n19551 , n3371 );
    xnor g32213 ( n34034 , n31297 , n22010 );
    and g32214 ( n19791 , n5558 , n6954 );
    or g32215 ( n34523 , n9964 , n1018 );
    and g32216 ( n22686 , n22971 , n27914 );
    xnor g32217 ( n30040 , n22491 , n16888 );
    or g32218 ( n14247 , n25933 , n17553 );
    or g32219 ( n20555 , n12753 , n5168 );
    or g32220 ( n19762 , n15744 , n4989 );
    or g32221 ( n1831 , n24562 , n18621 );
    or g32222 ( n30733 , n20353 , n16326 );
    not g32223 ( n22432 , n10894 );
    or g32224 ( n7009 , n33010 , n7726 );
    nor g32225 ( n22658 , n4878 , n32549 );
    xnor g32226 ( n9124 , n21529 , n12927 );
    buf g32227 ( n5779 , n6288 );
    xnor g32228 ( n35060 , n21321 , n5335 );
    or g32229 ( n23412 , n7828 , n8366 );
    or g32230 ( n24318 , n33441 , n26911 );
    or g32231 ( n23568 , n1570 , n26939 );
    and g32232 ( n1165 , n33939 , n18548 );
    or g32233 ( n27278 , n25850 , n22691 );
    or g32234 ( n13227 , n21654 , n23748 );
    nor g32235 ( n16615 , n4960 , n10918 );
    and g32236 ( n25775 , n15792 , n30590 );
    or g32237 ( n8858 , n24371 , n13104 );
    or g32238 ( n15532 , n6293 , n13350 );
    and g32239 ( n15890 , n4411 , n2655 );
    xnor g32240 ( n10509 , n14494 , n837 );
    nor g32241 ( n27408 , n33057 , n7929 );
    and g32242 ( n13127 , n10558 , n27709 );
    or g32243 ( n18434 , n1950 , n22268 );
    xnor g32244 ( n19406 , n27231 , n29237 );
    nor g32245 ( n23691 , n830 , n12753 );
    or g32246 ( n3098 , n3613 , n28636 );
    or g32247 ( n26269 , n9612 , n17162 );
    and g32248 ( n8796 , n1817 , n10473 );
    or g32249 ( n16452 , n3594 , n13235 );
    or g32250 ( n15219 , n9760 , n908 );
    and g32251 ( n33924 , n35336 , n31657 );
    or g32252 ( n1602 , n28175 , n7845 );
    nor g32253 ( n19807 , n22418 , n7748 );
    not g32254 ( n33014 , n1950 );
    and g32255 ( n16904 , n6270 , n17632 );
    not g32256 ( n25564 , n12264 );
    and g32257 ( n33778 , n13988 , n34747 );
    nor g32258 ( n22661 , n25813 , n25307 );
    xnor g32259 ( n34908 , n15659 , n32649 );
    not g32260 ( n22807 , n9236 );
    or g32261 ( n28473 , n17751 , n23040 );
    xnor g32262 ( n23447 , n11396 , n9069 );
    and g32263 ( n30217 , n15944 , n34522 );
    not g32264 ( n18372 , n35514 );
    or g32265 ( n24849 , n1510 , n1103 );
    xnor g32266 ( n4149 , n32674 , n15886 );
    or g32267 ( n35731 , n31180 , n9832 );
    and g32268 ( n9097 , n28861 , n33546 );
    or g32269 ( n4167 , n11049 , n25226 );
    buf g32270 ( n22946 , n23748 );
    or g32271 ( n18630 , n30963 , n33712 );
    or g32272 ( n21150 , n19513 , n11867 );
    or g32273 ( n28600 , n11648 , n4490 );
    xnor g32274 ( n26320 , n27067 , n14306 );
    and g32275 ( n18691 , n7433 , n19290 );
    and g32276 ( n14854 , n24843 , n16923 );
    or g32277 ( n13141 , n19927 , n25940 );
    and g32278 ( n27385 , n8912 , n35729 );
    or g32279 ( n35053 , n11413 , n24549 );
    buf g32280 ( n27963 , n11350 );
    or g32281 ( n29803 , n19191 , n511 );
    and g32282 ( n20596 , n32751 , n26422 );
    xnor g32283 ( n541 , n27008 , n1151 );
    and g32284 ( n30715 , n1199 , n2691 );
    nor g32285 ( n8466 , n31741 , n32379 );
    or g32286 ( n32895 , n3626 , n35935 );
    xnor g32287 ( n35750 , n32497 , n33335 );
    xnor g32288 ( n34155 , n5688 , n31444 );
    or g32289 ( n12568 , n9637 , n17368 );
    or g32290 ( n5323 , n7425 , n14476 );
    and g32291 ( n5336 , n33745 , n26858 );
    xnor g32292 ( n20858 , n4652 , n16371 );
    and g32293 ( n27863 , n23560 , n23966 );
    not g32294 ( n7212 , n27437 );
    or g32295 ( n8444 , n33864 , n2104 );
    not g32296 ( n35062 , n27226 );
    not g32297 ( n26774 , n15339 );
    or g32298 ( n28756 , n20064 , n3643 );
    and g32299 ( n12679 , n16402 , n3913 );
    or g32300 ( n12072 , n4878 , n1768 );
    and g32301 ( n11456 , n22623 , n8679 );
    nor g32302 ( n5534 , n7379 , n5887 );
    and g32303 ( n247 , n24997 , n29343 );
    or g32304 ( n17789 , n13877 , n30708 );
    or g32305 ( n1044 , n10286 , n32071 );
    or g32306 ( n15514 , n20662 , n10872 );
    not g32307 ( n15676 , n1950 );
    or g32308 ( n24911 , n3222 , n32883 );
    or g32309 ( n6978 , n10241 , n3679 );
    and g32310 ( n28868 , n10794 , n25335 );
    and g32311 ( n18018 , n1647 , n14359 );
    and g32312 ( n7470 , n3433 , n19174 );
    or g32313 ( n11301 , n16356 , n31967 );
    xnor g32314 ( n21374 , n18826 , n30295 );
    or g32315 ( n14418 , n19293 , n22647 );
    and g32316 ( n1656 , n92 , n19784 );
    not g32317 ( n6521 , n6288 );
    and g32318 ( n16805 , n8426 , n25591 );
    xnor g32319 ( n15311 , n33432 , n6066 );
    nor g32320 ( n34189 , n27154 , n9071 );
    xnor g32321 ( n25367 , n4423 , n17751 );
    or g32322 ( n30690 , n29375 , n10617 );
    xnor g32323 ( n20542 , n30352 , n25470 );
    and g32324 ( n18063 , n34817 , n11691 );
    or g32325 ( n2233 , n7419 , n1459 );
    or g32326 ( n17727 , n6388 , n9317 );
    xnor g32327 ( n1732 , n17129 , n34135 );
    and g32328 ( n28073 , n31573 , n18736 );
    and g32329 ( n7173 , n11871 , n15750 );
    and g32330 ( n30667 , n26273 , n2097 );
    xnor g32331 ( n6361 , n14006 , n11455 );
    nor g32332 ( n14821 , n31799 , n20448 );
    xnor g32333 ( n7663 , n21700 , n8432 );
    buf g32334 ( n27728 , n20255 );
    or g32335 ( n13832 , n17083 , n24374 );
    buf g32336 ( n26365 , n24095 );
    or g32337 ( n17708 , n28678 , n28675 );
    or g32338 ( n9863 , n35865 , n17829 );
    not g32339 ( n30754 , n8077 );
    or g32340 ( n29040 , n5788 , n1856 );
    or g32341 ( n5567 , n18660 , n1926 );
    and g32342 ( n33256 , n33077 , n25089 );
    or g32343 ( n2455 , n29451 , n28046 );
    xnor g32344 ( n13969 , n9392 , n15013 );
    xnor g32345 ( n30796 , n223 , n2774 );
    not g32346 ( n17640 , n2092 );
    xnor g32347 ( n27328 , n34100 , n772 );
    xnor g32348 ( n25772 , n10001 , n19984 );
    and g32349 ( n12143 , n21967 , n22033 );
    nor g32350 ( n33730 , n9715 , n28757 );
    and g32351 ( n7345 , n31616 , n14508 );
    and g32352 ( n7068 , n10480 , n8676 );
    xnor g32353 ( n6622 , n7951 , n33171 );
    or g32354 ( n6117 , n34082 , n32740 );
    and g32355 ( n2454 , n2995 , n32790 );
    xnor g32356 ( n28312 , n30139 , n19551 );
    xnor g32357 ( n5987 , n35791 , n19551 );
    or g32358 ( n9541 , n17568 , n28096 );
    or g32359 ( n9736 , n6131 , n32262 );
    not g32360 ( n33177 , n22501 );
    not g32361 ( n4998 , n9789 );
    and g32362 ( n28261 , n14549 , n18021 );
    or g32363 ( n10438 , n23203 , n10289 );
    xnor g32364 ( n8406 , n10370 , n34990 );
    xnor g32365 ( n882 , n33803 , n31559 );
    or g32366 ( n4910 , n28141 , n14268 );
    or g32367 ( n7097 , n8432 , n14025 );
    nor g32368 ( n1859 , n12650 , n11050 );
    or g32369 ( n6805 , n21396 , n30431 );
    and g32370 ( n28500 , n5027 , n24370 );
    or g32371 ( n9681 , n4962 , n31392 );
    and g32372 ( n14064 , n7992 , n27239 );
    xnor g32373 ( n70 , n29508 , n5335 );
    or g32374 ( n21690 , n7863 , n10995 );
    or g32375 ( n34689 , n15139 , n4279 );
    xnor g32376 ( n6063 , n16989 , n32095 );
    nor g32377 ( n14120 , n31799 , n30695 );
    and g32378 ( n19789 , n14529 , n17977 );
    not g32379 ( n33656 , n20427 );
    xnor g32380 ( n9717 , n6769 , n12299 );
    nor g32381 ( n11834 , n4758 , n5313 );
    not g32382 ( n9165 , n17568 );
    or g32383 ( n35125 , n15464 , n16403 );
    or g32384 ( n19357 , n22291 , n2700 );
    or g32385 ( n10154 , n20953 , n18692 );
    or g32386 ( n19898 , n19551 , n687 );
    xnor g32387 ( n13140 , n28417 , n14265 );
    nor g32388 ( n1416 , n21272 , n474 );
    or g32389 ( n6078 , n6094 , n7647 );
    xnor g32390 ( n18448 , n22381 , n21631 );
    xnor g32391 ( n33695 , n28247 , n4962 );
    or g32392 ( n34108 , n31559 , n17902 );
    not g32393 ( n34312 , n15403 );
    not g32394 ( n6890 , n25401 );
    and g32395 ( n35825 , n34263 , n13351 );
    or g32396 ( n26723 , n1950 , n17339 );
    or g32397 ( n9783 , n26250 , n6553 );
    or g32398 ( n22754 , n22668 , n3437 );
    or g32399 ( n20019 , n31761 , n8153 );
    xnor g32400 ( n26761 , n23108 , n34575 );
    nor g32401 ( n5233 , n15886 , n19097 );
    xnor g32402 ( n29883 , n8183 , n17168 );
    or g32403 ( n2070 , n16479 , n2712 );
    or g32404 ( n3232 , n27031 , n19464 );
    and g32405 ( n27192 , n11231 , n2554 );
    xnor g32406 ( n22090 , n31679 , n16995 );
    and g32407 ( n25223 , n27922 , n1144 );
    and g32408 ( n19629 , n35069 , n11668 );
    or g32409 ( n6963 , n13995 , n5972 );
    or g32410 ( n34950 , n3205 , n11959 );
    or g32411 ( n11890 , n34622 , n17782 );
    nor g32412 ( n8468 , n35927 , n29868 );
    xnor g32413 ( n1180 , n18754 , n10161 );
    or g32414 ( n27299 , n12797 , n17337 );
    not g32415 ( n15951 , n28603 );
    and g32416 ( n32452 , n29210 , n21065 );
    and g32417 ( n36038 , n17327 , n23645 );
    buf g32418 ( n28248 , n22667 );
    and g32419 ( n9069 , n8944 , n15579 );
    xnor g32420 ( n18613 , n3723 , n10430 );
    and g32421 ( n34063 , n2202 , n1108 );
    or g32422 ( n14273 , n1707 , n31627 );
    or g32423 ( n25700 , n31289 , n15291 );
    or g32424 ( n20317 , n26176 , n24672 );
    not g32425 ( n23339 , n9386 );
    or g32426 ( n1008 , n17521 , n10872 );
    and g32427 ( n24810 , n19480 , n6426 );
    or g32428 ( n11930 , n28964 , n32116 );
    xnor g32429 ( n22999 , n10818 , n22291 );
    not g32430 ( n34749 , n17568 );
    xnor g32431 ( n33645 , n20468 , n11046 );
    and g32432 ( n14249 , n20339 , n29966 );
    or g32433 ( n25064 , n25602 , n27102 );
    and g32434 ( n10885 , n18024 , n26140 );
    or g32435 ( n4434 , n12376 , n5752 );
    or g32436 ( n10994 , n28931 , n11850 );
    or g32437 ( n5128 , n31603 , n568 );
    xnor g32438 ( n17187 , n6022 , n33174 );
    not g32439 ( n24032 , n2568 );
    xnor g32440 ( n3974 , n35555 , n29713 );
    xnor g32441 ( n29490 , n657 , n31559 );
    and g32442 ( n19546 , n22863 , n23637 );
    xnor g32443 ( n26315 , n10839 , n32095 );
    and g32444 ( n35468 , n4384 , n523 );
    or g32445 ( n13091 , n23516 , n2168 );
    and g32446 ( n35604 , n23193 , n19340 );
    or g32447 ( n29031 , n31230 , n2282 );
    or g32448 ( n17838 , n27886 , n4683 );
    or g32449 ( n17819 , n35575 , n23462 );
    not g32450 ( n19837 , n31820 );
    xnor g32451 ( n30276 , n16884 , n29713 );
    buf g32452 ( n13307 , n25834 );
    and g32453 ( n4510 , n2332 , n33709 );
    or g32454 ( n6841 , n20752 , n31887 );
    not g32455 ( n15580 , n31994 );
    xnor g32456 ( n496 , n5746 , n20303 );
    or g32457 ( n10503 , n1741 , n29393 );
    nor g32458 ( n17135 , n2579 , n23425 );
    buf g32459 ( n8203 , n17628 );
    or g32460 ( n4815 , n28766 , n17018 );
    or g32461 ( n13626 , n29539 , n10140 );
    xnor g32462 ( n7996 , n9980 , n1117 );
    or g32463 ( n31983 , n9684 , n32329 );
    buf g32464 ( n4363 , n28404 );
    or g32465 ( n13990 , n32095 , n27401 );
    or g32466 ( n2565 , n13427 , n32071 );
    or g32467 ( n2783 , n15003 , n21862 );
    and g32468 ( n12136 , n9854 , n31910 );
    not g32469 ( n35998 , n30459 );
    or g32470 ( n24073 , n24371 , n25569 );
    or g32471 ( n7768 , n13611 , n5779 );
    xnor g32472 ( n18791 , n7191 , n22021 );
    not g32473 ( n35837 , n22595 );
    and g32474 ( n8680 , n24058 , n20296 );
    xnor g32475 ( n10654 , n35846 , n17887 );
    nor g32476 ( n4875 , n22767 , n12900 );
    xnor g32477 ( n6098 , n16534 , n31581 );
    and g32478 ( n11665 , n31890 , n13851 );
    xnor g32479 ( n2620 , n19777 , n20546 );
    or g32480 ( n7856 , n10261 , n12908 );
    xnor g32481 ( n13263 , n22035 , n5287 );
    not g32482 ( n9689 , n20972 );
    or g32483 ( n11429 , n19235 , n13305 );
    xnor g32484 ( n12512 , n27 , n1073 );
    or g32485 ( n35821 , n30704 , n17337 );
    xnor g32486 ( n18622 , n11259 , n27853 );
    or g32487 ( n29553 , n26785 , n21691 );
    or g32488 ( n19965 , n35875 , n19241 );
    and g32489 ( n35561 , n16447 , n7275 );
    or g32490 ( n18730 , n25006 , n15402 );
    or g32491 ( n30803 , n33319 , n34738 );
    xnor g32492 ( n19065 , n28306 , n4288 );
    and g32493 ( n36042 , n35430 , n8451 );
    nor g32494 ( n20327 , n26066 , n12428 );
    and g32495 ( n15642 , n18227 , n1585 );
    or g32496 ( n26562 , n20859 , n21436 );
    and g32497 ( n1371 , n17280 , n2884 );
    not g32498 ( n29121 , n31734 );
    buf g32499 ( n2524 , n22445 );
    xnor g32500 ( n22228 , n10492 , n16344 );
    or g32501 ( n16550 , n25515 , n15052 );
    or g32502 ( n32339 , n24686 , n1253 );
    xnor g32503 ( n23552 , n19838 , n28331 );
    or g32504 ( n13310 , n1764 , n23209 );
    or g32505 ( n5664 , n14251 , n19121 );
    xnor g32506 ( n21529 , n22723 , n4960 );
    and g32507 ( n17575 , n1587 , n10773 );
    xnor g32508 ( n32287 , n17307 , n10607 );
    and g32509 ( n22676 , n35396 , n26814 );
    not g32510 ( n34826 , n16801 );
    or g32511 ( n30169 , n31272 , n27456 );
    xnor g32512 ( n24506 , n21460 , n13337 );
    or g32513 ( n32487 , n28809 , n35374 );
    or g32514 ( n13054 , n28556 , n10246 );
    and g32515 ( n14322 , n24656 , n34348 );
    not g32516 ( n9430 , n24689 );
    or g32517 ( n1853 , n4288 , n212 );
    xnor g32518 ( n27 , n11359 , n30703 );
    and g32519 ( n8004 , n21633 , n6655 );
    nor g32520 ( n7682 , n22291 , n6644 );
    xnor g32521 ( n24717 , n15827 , n35927 );
    and g32522 ( n6341 , n13543 , n11105 );
    and g32523 ( n16415 , n23088 , n179 );
    not g32524 ( n28548 , n30459 );
    not g32525 ( n15825 , n12328 );
    or g32526 ( n23392 , n7269 , n35422 );
    or g32527 ( n22076 , n22693 , n8366 );
    or g32528 ( n28264 , n26125 , n5868 );
    not g32529 ( n9488 , n6288 );
    and g32530 ( n21903 , n19463 , n6881 );
    and g32531 ( n32224 , n17541 , n34252 );
    or g32532 ( n9419 , n29069 , n34084 );
    xnor g32533 ( n15190 , n27358 , n6686 );
    xnor g32534 ( n21299 , n9122 , n11095 );
    xnor g32535 ( n22547 , n14412 , n8997 );
    xnor g32536 ( n5354 , n11414 , n31739 );
    or g32537 ( n31539 , n7947 , n442 );
    or g32538 ( n826 , n32857 , n11426 );
    or g32539 ( n25407 , n22055 , n19228 );
    xnor g32540 ( n9095 , n26100 , n3946 );
    and g32541 ( n13681 , n4764 , n9774 );
    and g32542 ( n21868 , n24473 , n27515 );
    or g32543 ( n11694 , n32042 , n14218 );
    nor g32544 ( n14588 , n7473 , n27667 );
    or g32545 ( n11553 , n3205 , n15609 );
    or g32546 ( n25921 , n31215 , n16073 );
    or g32547 ( n4210 , n26670 , n29294 );
    or g32548 ( n32346 , n19300 , n11518 );
    and g32549 ( n31968 , n34240 , n21917 );
    not g32550 ( n31829 , n31272 );
    and g32551 ( n34283 , n10530 , n4873 );
    xnor g32552 ( n35323 , n35955 , n10630 );
    and g32553 ( n19420 , n33813 , n21728 );
    or g32554 ( n29126 , n2250 , n23419 );
    nor g32555 ( n18126 , n6360 , n6081 );
    xnor g32556 ( n34972 , n33357 , n15886 );
    or g32557 ( n32605 , n7170 , n29045 );
    and g32558 ( n34794 , n34732 , n28371 );
    or g32559 ( n18910 , n75 , n22501 );
    not g32560 ( n10866 , n32571 );
    and g32561 ( n16385 , n32369 , n11856 );
    or g32562 ( n14898 , n21357 , n1232 );
    and g32563 ( n27925 , n24076 , n8350 );
    xnor g32564 ( n18956 , n29421 , n35858 );
    and g32565 ( n33210 , n11232 , n30349 );
    or g32566 ( n14602 , n11046 , n9105 );
    not g32567 ( n12462 , n9821 );
    and g32568 ( n11680 , n314 , n33449 );
    buf g32569 ( n22783 , n26860 );
    and g32570 ( n13824 , n7536 , n10104 );
    nor g32571 ( n20638 , n31397 , n8761 );
    xnor g32572 ( n5173 , n17218 , n17221 );
    or g32573 ( n7266 , n14917 , n24696 );
    and g32574 ( n9684 , n14272 , n12416 );
    nor g32575 ( n31930 , n2189 , n1130 );
    not g32576 ( n12146 , n17202 );
    or g32577 ( n21820 , n16927 , n18947 );
    or g32578 ( n6783 , n5740 , n13857 );
    or g32579 ( n32655 , n17568 , n35948 );
    or g32580 ( n21157 , n14685 , n34323 );
    xnor g32581 ( n35239 , n3055 , n19636 );
    and g32582 ( n8404 , n23148 , n25849 );
    or g32583 ( n30924 , n1451 , n23187 );
    or g32584 ( n3433 , n25888 , n908 );
    and g32585 ( n25041 , n32018 , n24887 );
    or g32586 ( n21444 , n3946 , n14780 );
    and g32587 ( n5612 , n31462 , n19230 );
    buf g32588 ( n20840 , n27509 );
    or g32589 ( n10803 , n5392 , n4363 );
    xnor g32590 ( n21079 , n5048 , n4288 );
    nor g32591 ( n8185 , n6207 , n26672 );
    or g32592 ( n25944 , n33518 , n25594 );
    nor g32593 ( n3493 , n29839 , n367 );
    or g32594 ( n884 , n12657 , n34607 );
    xnor g32595 ( n29421 , n25068 , n29713 );
    xnor g32596 ( n9150 , n1739 , n32095 );
    or g32597 ( n33662 , n4288 , n4366 );
    and g32598 ( n8607 , n1460 , n23199 );
    nor g32599 ( n26119 , n27291 , n25817 );
    or g32600 ( n28093 , n10826 , n5732 );
    or g32601 ( n30029 , n24371 , n7670 );
    xnor g32602 ( n14393 , n34220 , n26305 );
    or g32603 ( n1255 , n16129 , n5213 );
    or g32604 ( n33845 , n26146 , n16457 );
    xnor g32605 ( n33573 , n29507 , n30426 );
    and g32606 ( n26225 , n8132 , n32428 );
    and g32607 ( n33848 , n35485 , n21302 );
    xnor g32608 ( n27271 , n2636 , n3205 );
    and g32609 ( n3395 , n16929 , n29477 );
    xnor g32610 ( n11334 , n23013 , n32715 );
    or g32611 ( n29915 , n22134 , n31075 );
    nor g32612 ( n6868 , n35770 , n6693 );
    nor g32613 ( n1774 , n10894 , n13234 );
    not g32614 ( n22575 , n4960 );
    and g32615 ( n36014 , n32333 , n23412 );
    and g32616 ( n10523 , n27059 , n5335 );
    xnor g32617 ( n8698 , n14929 , n3091 );
    or g32618 ( n32081 , n6990 , n13886 );
    or g32619 ( n11321 , n33096 , n16463 );
    nor g32620 ( n29485 , n32857 , n2099 );
    nor g32621 ( n26899 , n29713 , n11855 );
    or g32622 ( n33862 , n35927 , n348 );
    or g32623 ( n20451 , n25717 , n28969 );
    xnor g32624 ( n17623 , n35246 , n10663 );
    or g32625 ( n1022 , n10966 , n13797 );
    not g32626 ( n14751 , n21 );
    or g32627 ( n26284 , n32519 , n18954 );
    or g32628 ( n36070 , n16185 , n14962 );
    xnor g32629 ( n14187 , n23929 , n12252 );
    and g32630 ( n3686 , n3391 , n3200 );
    or g32631 ( n28164 , n14991 , n26578 );
    not g32632 ( n12178 , n35845 );
    not g32633 ( n28072 , n29203 );
    and g32634 ( n30799 , n21127 , n13953 );
    and g32635 ( n15656 , n29933 , n23235 );
    and g32636 ( n17562 , n12967 , n8999 );
    or g32637 ( n16964 , n19881 , n23626 );
    xnor g32638 ( n9821 , n33676 , n5215 );
    or g32639 ( n21789 , n19628 , n17162 );
    xnor g32640 ( n8307 , n236 , n8476 );
    nor g32641 ( n14245 , n1950 , n26732 );
    or g32642 ( n7463 , n25627 , n11980 );
    and g32643 ( n11940 , n27449 , n20196 );
    and g32644 ( n25273 , n3280 , n5182 );
    not g32645 ( n1323 , n13610 );
    and g32646 ( n29009 , n17017 , n4124 );
    or g32647 ( n17079 , n27291 , n25318 );
    and g32648 ( n30867 , n19667 , n17020 );
    or g32649 ( n2017 , n17864 , n27040 );
    and g32650 ( n18268 , n34682 , n27549 );
    xnor g32651 ( n30369 , n25131 , n29707 );
    or g32652 ( n12952 , n12028 , n11996 );
    nor g32653 ( n5772 , n9789 , n5092 );
    nor g32654 ( n23109 , n3946 , n27584 );
    and g32655 ( n14997 , n7989 , n17225 );
    xnor g32656 ( n19888 , n6148 , n12036 );
    nor g32657 ( n26802 , n32584 , n2630 );
    nor g32658 ( n9472 , n20057 , n949 );
    xnor g32659 ( n13387 , n383 , n1480 );
    xnor g32660 ( n22126 , n14905 , n34744 );
    or g32661 ( n14430 , n1122 , n28705 );
    or g32662 ( n26882 , n31339 , n13720 );
    and g32663 ( n9103 , n6546 , n33446 );
    xnor g32664 ( n1287 , n9172 , n28601 );
    nor g32665 ( n17868 , n4288 , n22066 );
    xnor g32666 ( n23424 , n8464 , n25252 );
    and g32667 ( n34225 , n19615 , n23978 );
    or g32668 ( n9459 , n16248 , n17974 );
    xnor g32669 ( n13065 , n27074 , n15414 );
    and g32670 ( n20722 , n612 , n4927 );
    or g32671 ( n26045 , n34138 , n27745 );
    xnor g32672 ( n5892 , n9260 , n11455 );
    not g32673 ( n12763 , n19442 );
    not g32674 ( n19483 , n5315 );
    or g32675 ( n33784 , n29993 , n33435 );
    and g32676 ( n33618 , n1760 , n22835 );
    and g32677 ( n12315 , n2114 , n15146 );
    not g32678 ( n16006 , n13841 );
    or g32679 ( n7780 , n8180 , n33063 );
    xnor g32680 ( n12486 , n5086 , n25701 );
    or g32681 ( n27032 , n13340 , n10432 );
    xnor g32682 ( n32153 , n7250 , n11046 );
    or g32683 ( n29806 , n2762 , n4135 );
    and g32684 ( n30234 , n15909 , n8172 );
    or g32685 ( n28259 , n7540 , n9141 );
    not g32686 ( n31100 , n23748 );
    xnor g32687 ( n10858 , n19469 , n19551 );
    or g32688 ( n21195 , n15886 , n1393 );
    xnor g32689 ( n30873 , n16678 , n1874 );
    or g32690 ( n8436 , n20211 , n24710 );
    or g32691 ( n13324 , n12841 , n2479 );
    not g32692 ( n35794 , n25602 );
    or g32693 ( n5009 , n26380 , n12175 );
    xnor g32694 ( n22063 , n10512 , n17181 );
    nor g32695 ( n36059 , n33815 , n7464 );
    xnor g32696 ( n30705 , n19450 , n4758 );
    and g32697 ( n16192 , n22654 , n11524 );
    and g32698 ( n32526 , n31115 , n17406 );
    or g32699 ( n31076 , n20376 , n6374 );
    and g32700 ( n13674 , n29664 , n871 );
    and g32701 ( n33007 , n8252 , n12619 );
    or g32702 ( n28279 , n4878 , n2622 );
    not g32703 ( n1700 , n35927 );
    not g32704 ( n19317 , n9789 );
    or g32705 ( n24379 , n8344 , n20812 );
    or g32706 ( n34947 , n3278 , n26329 );
    or g32707 ( n28083 , n13187 , n14035 );
    or g32708 ( n18904 , n7540 , n25463 );
    or g32709 ( n28032 , n29974 , n32076 );
    or g32710 ( n15635 , n19977 , n19421 );
    and g32711 ( n4460 , n21516 , n24657 );
    and g32712 ( n20101 , n26181 , n15106 );
    and g32713 ( n13332 , n17329 , n2294 );
    or g32714 ( n4236 , n20586 , n5234 );
    and g32715 ( n17598 , n12831 , n6578 );
    or g32716 ( n14093 , n8191 , n23748 );
    and g32717 ( n21916 , n17049 , n33760 );
    and g32718 ( n16768 , n27417 , n25843 );
    nor g32719 ( n11177 , n33890 , n35269 );
    and g32720 ( n1232 , n34779 , n30390 );
    or g32721 ( n15334 , n12384 , n17804 );
    or g32722 ( n31940 , n1201 , n34537 );
    or g32723 ( n5783 , n6713 , n19601 );
    or g32724 ( n2065 , n17157 , n21192 );
    and g32725 ( n27990 , n7983 , n26135 );
    xnor g32726 ( n11975 , n7589 , n25602 );
    or g32727 ( n16082 , n13041 , n3072 );
    and g32728 ( n5317 , n20893 , n20391 );
    xnor g32729 ( n18438 , n25760 , n11891 );
    or g32730 ( n35412 , n30885 , n24140 );
    xnor g32731 ( n27280 , n6541 , n4520 );
    or g32732 ( n12990 , n16845 , n23696 );
    or g32733 ( n923 , n35281 , n1462 );
    not g32734 ( n20862 , n10423 );
    or g32735 ( n18639 , n24371 , n4037 );
    and g32736 ( n27488 , n30052 , n26994 );
    and g32737 ( n7598 , n23568 , n33075 );
    and g32738 ( n30558 , n5928 , n14590 );
    and g32739 ( n10465 , n34339 , n8572 );
    or g32740 ( n17626 , n33043 , n21644 );
    or g32741 ( n17034 , n6372 , n27626 );
    and g32742 ( n33927 , n25860 , n22754 );
    or g32743 ( n10280 , n23706 , n3426 );
    or g32744 ( n22639 , n8951 , n34727 );
    or g32745 ( n24615 , n24713 , n16961 );
    or g32746 ( n10180 , n24371 , n19042 );
    xnor g32747 ( n3750 , n11565 , n25123 );
    and g32748 ( n12502 , n19231 , n6983 );
    or g32749 ( n18185 , n32707 , n4069 );
    xnor g32750 ( n35769 , n2685 , n6916 );
    xnor g32751 ( n11585 , n35947 , n28286 );
    nor g32752 ( n5840 , n4878 , n22570 );
    xnor g32753 ( n483 , n29599 , n19551 );
    not g32754 ( n18986 , n7834 );
    or g32755 ( n3140 , n19800 , n28705 );
    xnor g32756 ( n33319 , n9944 , n5287 );
    or g32757 ( n5911 , n20602 , n4175 );
    xnor g32758 ( n14803 , n33490 , n23300 );
    or g32759 ( n13756 , n29546 , n14770 );
    xnor g32760 ( n30828 , n7652 , n8161 );
    or g32761 ( n14542 , n15343 , n31464 );
    xnor g32762 ( n23092 , n32641 , n19551 );
    xnor g32763 ( n19093 , n13587 , n16974 );
    or g32764 ( n5405 , n32908 , n19306 );
    and g32765 ( n30499 , n34017 , n4890 );
    and g32766 ( n28513 , n12807 , n32376 );
    xnor g32767 ( n5466 , n9432 , n31780 );
    and g32768 ( n25342 , n6580 , n28471 );
    or g32769 ( n32619 , n13043 , n21202 );
    xnor g32770 ( n17670 , n20463 , n9658 );
    xnor g32771 ( n25563 , n34846 , n16451 );
    or g32772 ( n33866 , n32385 , n9675 );
    xnor g32773 ( n12630 , n16105 , n31215 );
    buf g32774 ( n17068 , n32147 );
    and g32775 ( n17052 , n24019 , n34266 );
    xnor g32776 ( n25176 , n23156 , n33209 );
    xnor g32777 ( n10575 , n26398 , n28536 );
    or g32778 ( n643 , n7208 , n21091 );
    and g32779 ( n673 , n17034 , n4759 );
    and g32780 ( n31819 , n21319 , n28269 );
    nor g32781 ( n20040 , n35156 , n19691 );
    xnor g32782 ( n9586 , n34061 , n33302 );
    or g32783 ( n30472 , n18064 , n16392 );
    or g32784 ( n35851 , n12813 , n31683 );
    xnor g32785 ( n12151 , n20934 , n35927 );
    and g32786 ( n3746 , n26850 , n29554 );
    or g32787 ( n14162 , n13637 , n16456 );
    nor g32788 ( n13897 , n7062 , n16649 );
    or g32789 ( n30849 , n19524 , n28969 );
    not g32790 ( n15506 , n11660 );
    and g32791 ( n29253 , n23152 , n18753 );
    xnor g32792 ( n12237 , n10454 , n7823 );
    xnor g32793 ( n1 , n10454 , n852 );
    or g32794 ( n24066 , n8494 , n16445 );
    not g32795 ( n12179 , n32510 );
    nor g32796 ( n35816 , n30742 , n25948 );
    xnor g32797 ( n4407 , n1452 , n1225 );
    and g32798 ( n25068 , n13853 , n4644 );
    nor g32799 ( n22855 , n14323 , n24287 );
    buf g32800 ( n28191 , n31100 );
    and g32801 ( n22522 , n1346 , n8546 );
    xnor g32802 ( n27383 , n35491 , n6509 );
    or g32803 ( n34930 , n34530 , n1715 );
    or g32804 ( n25083 , n12748 , n20360 );
    xnor g32805 ( n23047 , n12443 , n2927 );
    xnor g32806 ( n16164 , n16248 , n31056 );
    or g32807 ( n24532 , n27525 , n30646 );
    not g32808 ( n29375 , n19679 );
    or g32809 ( n32829 , n35989 , n4478 );
    or g32810 ( n15944 , n35371 , n30947 );
    xnor g32811 ( n4978 , n30080 , n11756 );
    xnor g32812 ( n23648 , n33089 , n2789 );
    xnor g32813 ( n4616 , n20015 , n35048 );
    or g32814 ( n34123 , n5335 , n19656 );
    not g32815 ( n27562 , n21820 );
    and g32816 ( n3019 , n14180 , n28234 );
    or g32817 ( n731 , n9346 , n23823 );
    xnor g32818 ( n2258 , n16490 , n25174 );
    or g32819 ( n27282 , n1837 , n4912 );
    xnor g32820 ( n12780 , n29886 , n16768 );
    not g32821 ( n11912 , n671 );
    buf g32822 ( n10872 , n21691 );
    not g32823 ( n15742 , n915 );
    xnor g32824 ( n5182 , n25445 , n31756 );
    xnor g32825 ( n25136 , n14528 , n4305 );
    or g32826 ( n21095 , n25819 , n8937 );
    or g32827 ( n13641 , n6449 , n16191 );
    and g32828 ( n21652 , n10775 , n19122 );
    not g32829 ( n21983 , n4878 );
    or g32830 ( n2107 , n9523 , n8723 );
    or g32831 ( n34153 , n16407 , n17111 );
    xnor g32832 ( n6466 , n29776 , n31253 );
    and g32833 ( n26907 , n15855 , n3452 );
    not g32834 ( n1299 , n27902 );
    or g32835 ( n1608 , n14971 , n12879 );
    xnor g32836 ( n15247 , n27169 , n30742 );
    or g32837 ( n16101 , n33597 , n5779 );
    and g32838 ( n27635 , n22581 , n27535 );
    nor g32839 ( n11250 , n19104 , n29203 );
    or g32840 ( n8169 , n15162 , n12465 );
    or g32841 ( n35172 , n19551 , n17785 );
    and g32842 ( n35108 , n16360 , n12153 );
    xnor g32843 ( n18864 , n4088 , n2108 );
    xnor g32844 ( n1512 , n28596 , n3184 );
    xnor g32845 ( n8849 , n35837 , n26166 );
    or g32846 ( n25333 , n30244 , n23323 );
    not g32847 ( n24610 , n11046 );
    or g32848 ( n4320 , n27676 , n26590 );
    and g32849 ( n30318 , n18645 , n24434 );
    or g32850 ( n26970 , n23447 , n14746 );
    and g32851 ( n27151 , n907 , n1893 );
    or g32852 ( n22812 , n10894 , n130 );
    and g32853 ( n30776 , n4820 , n21506 );
    or g32854 ( n18217 , n31453 , n763 );
    or g32855 ( n27981 , n3205 , n25035 );
    or g32856 ( n35068 , n4134 , n29953 );
    and g32857 ( n16499 , n4626 , n31398 );
    or g32858 ( n33942 , n13974 , n30383 );
    and g32859 ( n18005 , n15523 , n17197 );
    or g32860 ( n15465 , n19574 , n16457 );
    or g32861 ( n31716 , n4551 , n24356 );
    or g32862 ( n33122 , n19512 , n22522 );
    xnor g32863 ( n31637 , n14643 , n7474 );
    nor g32864 ( n11178 , n1847 , n19834 );
    or g32865 ( n33575 , n36023 , n2798 );
    or g32866 ( n14707 , n22291 , n18487 );
    xnor g32867 ( n30921 , n10407 , n31799 );
    and g32868 ( n10965 , n23321 , n24446 );
    or g32869 ( n12634 , n33555 , n13902 );
    and g32870 ( n22789 , n35622 , n35308 );
    and g32871 ( n26504 , n18975 , n30081 );
    xnor g32872 ( n17038 , n22972 , n25174 );
    or g32873 ( n10131 , n13123 , n13664 );
    or g32874 ( n24904 , n15807 , n4047 );
    or g32875 ( n33802 , n8062 , n35143 );
    xnor g32876 ( n28727 , n22177 , n24394 );
    or g32877 ( n22890 , n19126 , n21042 );
    nor g32878 ( n31127 , n4960 , n24168 );
    and g32879 ( n19069 , n14492 , n25805 );
    or g32880 ( n32324 , n31920 , n23217 );
    and g32881 ( n34482 , n1561 , n17819 );
    xnor g32882 ( n23556 , n18323 , n26806 );
    and g32883 ( n11914 , n26469 , n12627 );
    xnor g32884 ( n18141 , n10521 , n35783 );
    xnor g32885 ( n31043 , n22303 , n25602 );
    not g32886 ( n21677 , n27226 );
    or g32887 ( n6395 , n16163 , n33545 );
    and g32888 ( n31173 , n32210 , n22651 );
    or g32889 ( n3214 , n4878 , n13877 );
    or g32890 ( n24348 , n6769 , n12299 );
    or g32891 ( n9110 , n5368 , n26112 );
    or g32892 ( n27840 , n27082 , n17046 );
    or g32893 ( n35828 , n12782 , n34537 );
    or g32894 ( n32789 , n35241 , n10336 );
    and g32895 ( n10841 , n9445 , n33236 );
    or g32896 ( n28755 , n6703 , n15290 );
    or g32897 ( n635 , n21827 , n12465 );
    or g32898 ( n2709 , n31799 , n34152 );
    or g32899 ( n25916 , n4463 , n12913 );
    or g32900 ( n24541 , n3850 , n19562 );
    or g32901 ( n21946 , n11046 , n7583 );
    and g32902 ( n11881 , n26450 , n5084 );
    or g32903 ( n34988 , n12821 , n18876 );
    or g32904 ( n23200 , n21703 , n35935 );
    or g32905 ( n6446 , n1289 , n35402 );
    or g32906 ( n666 , n30342 , n4269 );
    or g32907 ( n33431 , n32095 , n30985 );
    and g32908 ( n18518 , n31326 , n18298 );
    xnor g32909 ( n27361 , n1719 , n20096 );
    or g32910 ( n29388 , n5708 , n5527 );
    or g32911 ( n35203 , n1231 , n18962 );
    and g32912 ( n19143 , n13313 , n20446 );
    or g32913 ( n19674 , n10786 , n4129 );
    nor g32914 ( n35064 , n8100 , n32186 );
    xnor g32915 ( n2765 , n14421 , n30405 );
    or g32916 ( n26139 , n8432 , n7916 );
    or g32917 ( n21362 , n31559 , n4840 );
    not g32918 ( n18844 , n26610 );
    or g32919 ( n1564 , n11635 , n19947 );
    xnor g32920 ( n5867 , n11326 , n5335 );
    or g32921 ( n25103 , n32890 , n35253 );
    and g32922 ( n17278 , n10419 , n5948 );
    and g32923 ( n5095 , n6532 , n7383 );
    nor g32924 ( n11019 , n29839 , n18183 );
    xnor g32925 ( n11807 , n28906 , n19984 );
    nor g32926 ( n23787 , n22513 , n9921 );
    or g32927 ( n10558 , n26438 , n10289 );
    xnor g32928 ( n12817 , n34641 , n6913 );
    or g32929 ( n35335 , n31124 , n5252 );
    xnor g32930 ( n20888 , n13798 , n2611 );
    xnor g32931 ( n14793 , n32883 , n3222 );
    and g32932 ( n14680 , n4867 , n18217 );
    or g32933 ( n2020 , n31775 , n15743 );
    and g32934 ( n29287 , n10150 , n215 );
    buf g32935 ( n9675 , n14706 );
    or g32936 ( n16786 , n24974 , n6288 );
    xnor g32937 ( n25024 , n18943 , n13975 );
    xnor g32938 ( n24372 , n20803 , n4078 );
    xnor g32939 ( n8945 , n19192 , n1520 );
    and g32940 ( n2538 , n12605 , n8261 );
    and g32941 ( n14283 , n13423 , n18199 );
    and g32942 ( n10676 , n6493 , n10977 );
    and g32943 ( n22419 , n33342 , n5240 );
    and g32944 ( n10219 , n4899 , n11698 );
    or g32945 ( n12760 , n15678 , n19421 );
    and g32946 ( n4130 , n10936 , n3270 );
    or g32947 ( n34326 , n17237 , n6042 );
    or g32948 ( n6708 , n25636 , n19403 );
    or g32949 ( n7825 , n14389 , n27923 );
    and g32950 ( n10243 , n33584 , n32358 );
    or g32951 ( n32123 , n17174 , n5249 );
    or g32952 ( n26182 , n830 , n13033 );
    or g32953 ( n26328 , n15771 , n26468 );
    not g32954 ( n12061 , n11507 );
    and g32955 ( n4530 , n17198 , n3108 );
    xnor g32956 ( n35639 , n922 , n6818 );
    xnor g32957 ( n5473 , n1573 , n8593 );
    xnor g32958 ( n12115 , n20880 , n6742 );
    xnor g32959 ( n4088 , n3821 , n24371 );
    and g32960 ( n5351 , n35335 , n31 );
    or g32961 ( n28328 , n8613 , n31606 );
    and g32962 ( n10545 , n2603 , n8558 );
    or g32963 ( n17549 , n9181 , n21621 );
    nor g32964 ( n7668 , n13610 , n23187 );
    xnor g32965 ( n10784 , n12189 , n19786 );
    or g32966 ( n17391 , n9789 , n19550 );
    xnor g32967 ( n4631 , n14031 , n3088 );
    or g32968 ( n4375 , n26799 , n28191 );
    xnor g32969 ( n24196 , n20619 , n16196 );
    or g32970 ( n20122 , n31809 , n4478 );
    nor g32971 ( n3535 , n1950 , n29397 );
    xnor g32972 ( n35255 , n31330 , n33293 );
    and g32973 ( n4246 , n27165 , n24543 );
    xnor g32974 ( n8428 , n11454 , n12412 );
    and g32975 ( n1042 , n1646 , n26155 );
    or g32976 ( n778 , n4960 , n11501 );
    not g32977 ( n12821 , n11265 );
    nor g32978 ( n22434 , n19551 , n6880 );
    nor g32979 ( n18914 , n11455 , n29611 );
    xnor g32980 ( n10940 , n4204 , n33218 );
    nor g32981 ( n11906 , n11887 , n33956 );
    or g32982 ( n25161 , n8234 , n13492 );
    or g32983 ( n24609 , n29969 , n32198 );
    and g32984 ( n23744 , n11799 , n31623 );
    xnor g32985 ( n27800 , n4547 , n24965 );
    or g32986 ( n18170 , n21804 , n15754 );
    nor g32987 ( n30514 , n1327 , n4108 );
    xnor g32988 ( n28155 , n24684 , n32944 );
    or g32989 ( n23734 , n6031 , n35589 );
    or g32990 ( n10080 , n19380 , n28404 );
    and g32991 ( n9028 , n35203 , n23958 );
    xnor g32992 ( n20237 , n1726 , n19979 );
    or g32993 ( n248 , n13355 , n17294 );
    not g32994 ( n22357 , n29839 );
    xnor g32995 ( n30298 , n14600 , n9147 );
    or g32996 ( n31188 , n25749 , n8480 );
    nor g32997 ( n12680 , n2764 , n2607 );
    not g32998 ( n33387 , n15544 );
    or g32999 ( n1308 , n19677 , n28191 );
    not g33000 ( n18698 , n544 );
    xnor g33001 ( n3909 , n26267 , n22291 );
    xnor g33002 ( n14832 , n23052 , n4962 );
    xnor g33003 ( n31209 , n22994 , n33218 );
    or g33004 ( n8133 , n33164 , n11511 );
    or g33005 ( n17091 , n24714 , n25619 );
    xnor g33006 ( n18006 , n9418 , n30742 );
    xnor g33007 ( n32418 , n5117 , n8432 );
    or g33008 ( n10525 , n29140 , n30419 );
    xnor g33009 ( n21057 , n11152 , n16471 );
    and g33010 ( n18930 , n25087 , n21172 );
    or g33011 ( n16170 , n31106 , n10822 );
    or g33012 ( n28938 , n21961 , n29743 );
    and g33013 ( n31823 , n25042 , n20054 );
    xnor g33014 ( n20709 , n13082 , n1815 );
    nor g33015 ( n25006 , n15886 , n17524 );
    or g33016 ( n11094 , n24371 , n22734 );
    xnor g33017 ( n22056 , n14687 , n4288 );
    nor g33018 ( n30561 , n20332 , n26794 );
    or g33019 ( n816 , n25431 , n22661 );
    not g33020 ( n33457 , n17568 );
    and g33021 ( n17690 , n19153 , n16857 );
    and g33022 ( n27978 , n31816 , n31036 );
    xnor g33023 ( n20856 , n2893 , n4271 );
    not g33024 ( n23564 , n21976 );
    xnor g33025 ( n30186 , n7702 , n21944 );
    or g33026 ( n4317 , n4288 , n13037 );
    xnor g33027 ( n18551 , n31949 , n25602 );
    and g33028 ( n32570 , n27281 , n4622 );
    or g33029 ( n19651 , n3256 , n20300 );
    xnor g33030 ( n29362 , n16169 , n30742 );
    not g33031 ( n13909 , n20427 );
    and g33032 ( n10544 , n8700 , n13156 );
    or g33033 ( n22439 , n29552 , n1557 );
    xnor g33034 ( n34567 , n20487 , n31943 );
    or g33035 ( n31262 , n8042 , n7065 );
    xnor g33036 ( n13418 , n22914 , n24332 );
    or g33037 ( n20928 , n16922 , n2511 );
    or g33038 ( n29449 , n8711 , n21042 );
    or g33039 ( n2032 , n19404 , n30826 );
    xnor g33040 ( n5372 , n4149 , n1997 );
    and g33041 ( n23266 , n7207 , n24358 );
    or g33042 ( n3381 , n15596 , n15496 );
    buf g33043 ( n7153 , n25472 );
    or g33044 ( n35901 , n3504 , n34722 );
    and g33045 ( n20604 , n33022 , n32367 );
    and g33046 ( n27584 , n16118 , n12316 );
    and g33047 ( n14785 , n27639 , n24992 );
    and g33048 ( n25488 , n7258 , n34202 );
    xnor g33049 ( n13728 , n22209 , n16135 );
    nor g33050 ( n27234 , n30964 , n23378 );
    nor g33051 ( n25319 , n9793 , n27763 );
    or g33052 ( n18953 , n24822 , n1642 );
    or g33053 ( n28059 , n18432 , n28668 );
    or g33054 ( n6910 , n29363 , n4254 );
    or g33055 ( n26863 , n25750 , n21579 );
    or g33056 ( n35783 , n26699 , n21687 );
    xnor g33057 ( n1020 , n5334 , n34372 );
    or g33058 ( n6457 , n17002 , n13305 );
    or g33059 ( n30309 , n4758 , n27254 );
    xnor g33060 ( n18755 , n24583 , n25922 );
    or g33061 ( n11394 , n21606 , n13664 );
    and g33062 ( n5891 , n21938 , n18439 );
    or g33063 ( n20234 , n18808 , n3417 );
    or g33064 ( n21517 , n23604 , n4673 );
    or g33065 ( n18028 , n7540 , n33250 );
    not g33066 ( n29432 , n14033 );
    xnor g33067 ( n33555 , n26037 , n7540 );
    buf g33068 ( n22206 , n23348 );
    nor g33069 ( n25452 , n31289 , n35202 );
    xnor g33070 ( n14899 , n23590 , n10644 );
    xnor g33071 ( n17803 , n18180 , n13096 );
    or g33072 ( n14188 , n19210 , n27447 );
    xnor g33073 ( n12091 , n169 , n27291 );
    not g33074 ( n23421 , n4288 );
    not g33075 ( n14716 , n18296 );
    or g33076 ( n26223 , n12621 , n15290 );
    or g33077 ( n29734 , n9658 , n10887 );
    or g33078 ( n9638 , n11225 , n13217 );
    xnor g33079 ( n35363 , n22182 , n23099 );
    xnor g33080 ( n20646 , n11156 , n24371 );
    xnor g33081 ( n18082 , n28634 , n4687 );
    or g33082 ( n21491 , n10894 , n2991 );
    or g33083 ( n18117 , n22301 , n7153 );
    not g33084 ( n9463 , n11265 );
    xnor g33085 ( n21601 , n9816 , n35927 );
    xnor g33086 ( n34443 , n19934 , n25602 );
    xnor g33087 ( n4365 , n23466 , n4962 );
    xnor g33088 ( n29387 , n23102 , n4960 );
    nor g33089 ( n14967 , n19551 , n27008 );
    or g33090 ( n7394 , n3008 , n1856 );
    or g33091 ( n24282 , n28848 , n22448 );
    not g33092 ( n25456 , n3205 );
    xnor g33093 ( n34492 , n228 , n27705 );
    or g33094 ( n28197 , n15972 , n4363 );
    xnor g33095 ( n21504 , n24424 , n1019 );
    or g33096 ( n6493 , n11719 , n35306 );
    or g33097 ( n29973 , n9793 , n17788 );
    not g33098 ( n13224 , n11455 );
    or g33099 ( n21805 , n35533 , n6178 );
    xnor g33100 ( n33176 , n7826 , n35148 );
    not g33101 ( n12662 , n14148 );
    not g33102 ( n15744 , n22980 );
    or g33103 ( n36002 , n31440 , n35187 );
    xnor g33104 ( n18678 , n2451 , n9278 );
    or g33105 ( n16549 , n13719 , n14535 );
    or g33106 ( n31847 , n17851 , n8090 );
    xnor g33107 ( n12681 , n1088 , n14410 );
    or g33108 ( n6335 , n26010 , n34971 );
    and g33109 ( n22972 , n11394 , n21363 );
    or g33110 ( n23296 , n7110 , n10336 );
    and g33111 ( n12876 , n29797 , n30784 );
    xnor g33112 ( n10041 , n33112 , n29839 );
    not g33113 ( n28964 , n20882 );
    xnor g33114 ( n4322 , n7399 , n32095 );
    or g33115 ( n11062 , n152 , n3858 );
    and g33116 ( n33462 , n26914 , n706 );
    xnor g33117 ( n289 , n13226 , n22926 );
    and g33118 ( n32666 , n4581 , n11453 );
    and g33119 ( n14072 , n32948 , n9070 );
    or g33120 ( n5011 , n16922 , n20387 );
    and g33121 ( n13801 , n17883 , n30484 );
    or g33122 ( n16098 , n10294 , n33310 );
    xnor g33123 ( n9893 , n4037 , n24371 );
    and g33124 ( n3922 , n13118 , n28980 );
    not g33125 ( n6024 , n32608 );
    or g33126 ( n8863 , n14341 , n25895 );
    nor g33127 ( n24973 , n29787 , n8153 );
    xnor g33128 ( n19048 , n1120 , n12515 );
    or g33129 ( n7526 , n34224 , n24259 );
    xnor g33130 ( n9432 , n13368 , n19984 );
    not g33131 ( n2831 , n28853 );
    and g33132 ( n3510 , n4049 , n5363 );
    xnor g33133 ( n18225 , n4513 , n10142 );
    xnor g33134 ( n18422 , n20109 , n12764 );
    or g33135 ( n6090 , n19229 , n665 );
    not g33136 ( n9663 , n14646 );
    and g33137 ( n3742 , n3122 , n9659 );
    and g33138 ( n24867 , n9013 , n32269 );
    or g33139 ( n12200 , n27892 , n15620 );
    nor g33140 ( n31783 , n9658 , n20460 );
    and g33141 ( n24222 , n4111 , n20275 );
    and g33142 ( n30721 , n12577 , n26639 );
    not g33143 ( n8761 , n14136 );
    or g33144 ( n28177 , n29146 , n12834 );
    or g33145 ( n17163 , n26003 , n8101 );
    xnor g33146 ( n30854 , n20264 , n14984 );
    and g33147 ( n13718 , n33909 , n28704 );
    or g33148 ( n24481 , n17743 , n834 );
    xnor g33149 ( n22568 , n29298 , n17170 );
    not g33150 ( n7928 , n12659 );
    xnor g33151 ( n19054 , n2091 , n17568 );
    and g33152 ( n2494 , n11191 , n17880 );
    and g33153 ( n26823 , n11119 , n34882 );
    or g33154 ( n32475 , n30096 , n4318 );
    xnor g33155 ( n33019 , n13418 , n4095 );
    xnor g33156 ( n12617 , n7887 , n28360 );
    or g33157 ( n8333 , n10434 , n8886 );
    or g33158 ( n10224 , n24606 , n5618 );
    or g33159 ( n26297 , n3711 , n6288 );
    not g33160 ( n31339 , n35950 );
    not g33161 ( n27621 , n24010 );
    nor g33162 ( n32749 , n33650 , n25567 );
    or g33163 ( n23726 , n3343 , n20789 );
    and g33164 ( n19574 , n26040 , n13675 );
    not g33165 ( n33596 , n15096 );
    or g33166 ( n17583 , n29639 , n30431 );
    and g33167 ( n21164 , n5258 , n18068 );
    and g33168 ( n9831 , n23296 , n17792 );
    or g33169 ( n33085 , n1609 , n16262 );
    or g33170 ( n29826 , n31841 , n9079 );
    or g33171 ( n19805 , n14964 , n15250 );
    or g33172 ( n12572 , n35212 , n28675 );
    xnor g33173 ( n173 , n24796 , n5051 );
    xnor g33174 ( n4073 , n25066 , n4962 );
    not g33175 ( n35010 , n22305 );
    or g33176 ( n21686 , n26078 , n2005 );
    and g33177 ( n14842 , n3373 , n17567 );
    not g33178 ( n21622 , n32089 );
    xnor g33179 ( n33214 , n11995 , n5137 );
    or g33180 ( n9636 , n27025 , n7993 );
    xnor g33181 ( n17852 , n27100 , n16620 );
    or g33182 ( n6420 , n11228 , n4081 );
    or g33183 ( n35061 , n25893 , n2984 );
    and g33184 ( n35543 , n8949 , n32360 );
    not g33185 ( n27961 , n31056 );
    and g33186 ( n14765 , n11288 , n11695 );
    and g33187 ( n12217 , n11236 , n8089 );
    or g33188 ( n11696 , n18613 , n14716 );
    or g33189 ( n25494 , n11084 , n17964 );
    buf g33190 ( n17964 , n30940 );
    xnor g33191 ( n18418 , n13748 , n22577 );
    or g33192 ( n6809 , n21893 , n3437 );
    or g33193 ( n32205 , n9101 , n2262 );
    or g33194 ( n6799 , n35579 , n22322 );
    buf g33195 ( n21956 , n28816 );
    or g33196 ( n6788 , n8740 , n7726 );
    nor g33197 ( n26673 , n4288 , n15316 );
    or g33198 ( n20557 , n12398 , n1856 );
    nor g33199 ( n21765 , n21200 , n6548 );
    nor g33200 ( n9244 , n25602 , n18377 );
    or g33201 ( n2054 , n17754 , n17233 );
    or g33202 ( n7824 , n27291 , n31220 );
    or g33203 ( n11140 , n25858 , n9930 );
    or g33204 ( n372 , n27036 , n25459 );
    nor g33205 ( n16149 , n29902 , n9661 );
    and g33206 ( n3652 , n8204 , n431 );
    or g33207 ( n24467 , n25174 , n23840 );
    or g33208 ( n23247 , n2434 , n19241 );
    or g33209 ( n11832 , n10125 , n24489 );
    xnor g33210 ( n22755 , n32322 , n4960 );
    or g33211 ( n21850 , n8432 , n32739 );
    not g33212 ( n1142 , n30292 );
    nor g33213 ( n23934 , n30742 , n20531 );
    xnor g33214 ( n9836 , n4115 , n13519 );
    and g33215 ( n35294 , n4315 , n10964 );
    nor g33216 ( n24042 , n3946 , n5476 );
    or g33217 ( n20657 , n21201 , n1763 );
    xor g33218 ( n8094 , n34783 , n19513 );
    xnor g33219 ( n14613 , n13243 , n16108 );
    and g33220 ( n31782 , n86 , n5401 );
    xnor g33221 ( n386 , n4889 , n12806 );
    nor g33222 ( n25617 , n34717 , n35417 );
    or g33223 ( n15104 , n18379 , n10199 );
    and g33224 ( n8840 , n2087 , n4198 );
    nor g33225 ( n11616 , n4960 , n20687 );
    xnor g33226 ( n5018 , n9075 , n17115 );
    not g33227 ( n27671 , n11780 );
    and g33228 ( n2271 , n8809 , n35738 );
    and g33229 ( n18207 , n31738 , n6896 );
    xnor g33230 ( n5761 , n1723 , n23604 );
    and g33231 ( n14774 , n31695 , n28849 );
    and g33232 ( n25866 , n6687 , n7076 );
    not g33233 ( n17945 , n25191 );
    or g33234 ( n4146 , n4960 , n31107 );
    and g33235 ( n24979 , n29668 , n4474 );
    and g33236 ( n12663 , n22087 , n2869 );
    or g33237 ( n28912 , n6996 , n10933 );
    xnor g33238 ( n33082 , n5535 , n32281 );
    or g33239 ( n15126 , n13268 , n18047 );
    or g33240 ( n34647 , n31077 , n7086 );
    or g33241 ( n34734 , n8914 , n11833 );
    or g33242 ( n19108 , n24371 , n12502 );
    or g33243 ( n2968 , n26015 , n13290 );
    not g33244 ( n35894 , n4293 );
    xnor g33245 ( n26597 , n19785 , n30662 );
    and g33246 ( n14794 , n21899 , n9697 );
    or g33247 ( n35440 , n4028 , n23663 );
    or g33248 ( n17358 , n30747 , n32507 );
    or g33249 ( n21004 , n9789 , n25234 );
    not g33250 ( n33140 , n34865 );
    or g33251 ( n32986 , n22280 , n33896 );
    buf g33252 ( n16961 , n24022 );
    or g33253 ( n17808 , n5577 , n16461 );
    or g33254 ( n25453 , n7302 , n23187 );
    or g33255 ( n4741 , n3205 , n4594 );
    or g33256 ( n15080 , n17061 , n19105 );
    xnor g33257 ( n3735 , n29791 , n27855 );
    and g33258 ( n35741 , n24568 , n23827 );
    or g33259 ( n29179 , n15005 , n25831 );
    or g33260 ( n12031 , n14649 , n19732 );
    and g33261 ( n10529 , n23248 , n26710 );
    xnor g33262 ( n11206 , n9068 , n2446 );
    and g33263 ( n33964 , n32271 , n17666 );
    not g33264 ( n1227 , n30125 );
    xnor g33265 ( n25902 , n26436 , n29760 );
    xnor g33266 ( n14947 , n25426 , n24746 );
    not g33267 ( n10127 , n18296 );
    or g33268 ( n3334 , n20260 , n6950 );
    or g33269 ( n18325 , n31356 , n22316 );
    xnor g33270 ( n30531 , n15987 , n3222 );
    xnor g33271 ( n24337 , n24306 , n2722 );
    xnor g33272 ( n15108 , n35356 , n24371 );
    or g33273 ( n12243 , n30368 , n23626 );
    xnor g33274 ( n4837 , n8699 , n3329 );
    and g33275 ( n35197 , n34079 , n29944 );
    or g33276 ( n35213 , n29159 , n19265 );
    and g33277 ( n27355 , n28790 , n28679 );
    and g33278 ( n14910 , n9512 , n20381 );
    or g33279 ( n17320 , n27616 , n5615 );
    or g33280 ( n562 , n24760 , n22322 );
    xnor g33281 ( n29470 , n26615 , n25194 );
    or g33282 ( n16229 , n15457 , n21042 );
    or g33283 ( n29111 , n29068 , n33403 );
    or g33284 ( n8646 , n34706 , n5800 );
    not g33285 ( n5459 , n32427 );
    or g33286 ( n11619 , n35553 , n31854 );
    nor g33287 ( n21645 , n4758 , n1931 );
    and g33288 ( n34973 , n11352 , n5838 );
    or g33289 ( n9335 , n14444 , n16457 );
    xnor g33290 ( n27766 , n9076 , n14798 );
    or g33291 ( n1210 , n10894 , n31523 );
    or g33292 ( n24994 , n32095 , n19827 );
    and g33293 ( n5197 , n31944 , n35343 );
    xnor g33294 ( n10461 , n8191 , n16922 );
    xnor g33295 ( n15787 , n738 , n25904 );
    or g33296 ( n16009 , n19855 , n19732 );
    and g33297 ( n19589 , n4505 , n12957 );
    or g33298 ( n5632 , n22361 , n5626 );
    and g33299 ( n1297 , n14880 , n29695 );
    not g33300 ( n5547 , n3205 );
    and g33301 ( n12394 , n17335 , n10540 );
    or g33302 ( n23712 , n21236 , n6251 );
    and g33303 ( n6278 , n21876 , n21790 );
    or g33304 ( n34779 , n17783 , n35072 );
    and g33305 ( n4829 , n18200 , n4813 );
    and g33306 ( n2849 , n6778 , n8762 );
    xnor g33307 ( n15767 , n33250 , n7540 );
    xnor g33308 ( n3068 , n12213 , n23434 );
    and g33309 ( n3316 , n19962 , n8961 );
    or g33310 ( n12404 , n1950 , n6589 );
    xnor g33311 ( n1959 , n35327 , n25174 );
    xnor g33312 ( n23646 , n33334 , n23299 );
    and g33313 ( n22120 , n15917 , n10454 );
    not g33314 ( n10820 , n7504 );
    xnor g33315 ( n26180 , n4845 , n30255 );
    and g33316 ( n20352 , n2743 , n4741 );
    or g33317 ( n2203 , n26729 , n22501 );
    not g33318 ( n34359 , n25260 );
    xnor g33319 ( n29246 , n209 , n24587 );
    or g33320 ( n16587 , n25417 , n32593 );
    and g33321 ( n16357 , n15420 , n403 );
    or g33322 ( n20374 , n10660 , n31589 );
    and g33323 ( n3006 , n22813 , n30574 );
    and g33324 ( n4675 , n22171 , n19232 );
    and g33325 ( n21684 , n34164 , n34755 );
    buf g33326 ( n35043 , n25592 );
    or g33327 ( n29636 , n656 , n21318 );
    or g33328 ( n14608 , n12467 , n7726 );
    or g33329 ( n22525 , n21345 , n2005 );
    not g33330 ( n1941 , n3205 );
    and g33331 ( n14817 , n31908 , n21204 );
    xnor g33332 ( n11654 , n32739 , n8432 );
    and g33333 ( n17249 , n14385 , n34576 );
    or g33334 ( n15443 , n10321 , n23323 );
    and g33335 ( n2611 , n27047 , n14810 );
    xnor g33336 ( n23824 , n25267 , n23604 );
    nor g33337 ( n6767 , n830 , n29444 );
    or g33338 ( n31130 , n9421 , n31464 );
    and g33339 ( n22479 , n13314 , n21437 );
    and g33340 ( n21533 , n25718 , n27425 );
    xnor g33341 ( n20671 , n35645 , n11794 );
    xnor g33342 ( n18814 , n34662 , n19069 );
    nor g33343 ( n13808 , n30619 , n13823 );
    or g33344 ( n11431 , n34192 , n33310 );
    and g33345 ( n15169 , n19179 , n35245 );
    or g33346 ( n31010 , n31799 , n19789 );
    or g33347 ( n30341 , n7682 , n33776 );
    not g33348 ( n7830 , n31289 );
    or g33349 ( n28523 , n35847 , n3858 );
    or g33350 ( n33957 , n13486 , n12381 );
    or g33351 ( n28069 , n3205 , n7978 );
    xnor g33352 ( n11020 , n33433 , n17568 );
    or g33353 ( n19765 , n24251 , n21625 );
    nor g33354 ( n24921 , n32584 , n427 );
    or g33355 ( n10807 , n4468 , n30431 );
    buf g33356 ( n17204 , n24479 );
    nor g33357 ( n9744 , n12778 , n25910 );
    or g33358 ( n9701 , n21465 , n17337 );
    and g33359 ( n28451 , n18104 , n3969 );
    and g33360 ( n22495 , n35285 , n30249 );
    or g33361 ( n20580 , n10894 , n20829 );
    not g33362 ( n19104 , n20462 );
    xnor g33363 ( n19622 , n18626 , n29118 );
    or g33364 ( n32575 , n12229 , n31055 );
    and g33365 ( n30013 , n8545 , n6776 );
    not g33366 ( n24330 , n27859 );
    nor g33367 ( n2456 , n4960 , n26719 );
    or g33368 ( n35389 , n15509 , n25773 );
    or g33369 ( n29016 , n34697 , n5168 );
    and g33370 ( n11246 , n12862 , n13136 );
    or g33371 ( n17472 , n13508 , n34610 );
    and g33372 ( n13261 , n35240 , n14705 );
    and g33373 ( n16595 , n27993 , n25453 );
    and g33374 ( n13563 , n16013 , n30846 );
    and g33375 ( n28330 , n31385 , n27754 );
    or g33376 ( n10613 , n4960 , n5451 );
    or g33377 ( n35450 , n26099 , n7673 );
    and g33378 ( n17306 , n35090 , n3817 );
    or g33379 ( n19647 , n18585 , n5900 );
    and g33380 ( n11805 , n13040 , n13829 );
    not g33381 ( n20865 , n1433 );
    or g33382 ( n8194 , n23064 , n32697 );
    not g33383 ( n7671 , n1540 );
    or g33384 ( n7567 , n18573 , n4970 );
    nor g33385 ( n3431 , n11705 , n13511 );
    or g33386 ( n7010 , n1950 , n22676 );
    and g33387 ( n2729 , n22608 , n23616 );
    not g33388 ( n17297 , n6879 );
    nor g33389 ( n26787 , n30742 , n27352 );
    and g33390 ( n13544 , n25649 , n17584 );
    and g33391 ( n33685 , n10534 , n15192 );
    and g33392 ( n20344 , n35018 , n22441 );
    or g33393 ( n26553 , n20286 , n30150 );
    and g33394 ( n17413 , n22772 , n1004 );
    and g33395 ( n22416 , n1366 , n6263 );
    nor g33396 ( n13859 , n30742 , n8606 );
    or g33397 ( n31019 , n3222 , n21159 );
    nor g33398 ( n34711 , n18572 , n24827 );
    or g33399 ( n2426 , n2575 , n2117 );
    xnor g33400 ( n10244 , n13176 , n10862 );
    and g33401 ( n24553 , n25599 , n25626 );
    or g33402 ( n2695 , n31507 , n13664 );
    or g33403 ( n13569 , n32577 , n33124 );
    or g33404 ( n19149 , n1850 , n11128 );
    or g33405 ( n21575 , n18244 , n17068 );
    or g33406 ( n12204 , n26351 , n6288 );
    not g33407 ( n34470 , n18739 );
    or g33408 ( n22005 , n23925 , n27580 );
    xnor g33409 ( n22193 , n22317 , n21338 );
    not g33410 ( n16710 , n20840 );
    not g33411 ( n17120 , n29018 );
    and g33412 ( n32981 , n26006 , n17556 );
    or g33413 ( n2121 , n17751 , n31068 );
    and g33414 ( n5936 , n3328 , n21238 );
    or g33415 ( n24377 , n9658 , n20463 );
    and g33416 ( n10281 , n33254 , n34929 );
    and g33417 ( n11713 , n7738 , n11383 );
    xnor g33418 ( n24947 , n18475 , n324 );
    or g33419 ( n28495 , n29839 , n25775 );
    and g33420 ( n25448 , n11957 , n25403 );
    not g33421 ( n35423 , n30009 );
    and g33422 ( n27773 , n14195 , n7307 );
    and g33423 ( n33878 , n6577 , n22704 );
    or g33424 ( n31573 , n4830 , n29592 );
    xnor g33425 ( n25461 , n19394 , n2860 );
    or g33426 ( n28402 , n35936 , n28064 );
    and g33427 ( n34745 , n426 , n31499 );
    or g33428 ( n1800 , n13773 , n22604 );
    or g33429 ( n30414 , n8717 , n31621 );
    xnor g33430 ( n32319 , n24602 , n11463 );
    or g33431 ( n31908 , n25688 , n19403 );
    or g33432 ( n11994 , n21890 , n9317 );
    and g33433 ( n32694 , n24767 , n7279 );
    xnor g33434 ( n12661 , n18838 , n19551 );
    xnor g33435 ( n7213 , n23849 , n14328 );
    or g33436 ( n25481 , n35765 , n25940 );
    and g33437 ( n31757 , n8218 , n2102 );
    not g33438 ( n26826 , n22200 );
    and g33439 ( n9325 , n15137 , n19683 );
    or g33440 ( n33872 , n10821 , n12791 );
    xnor g33441 ( n25243 , n28707 , n19446 );
    or g33442 ( n29757 , n18562 , n24356 );
    buf g33443 ( n23209 , n24581 );
    or g33444 ( n28460 , n30298 , n23462 );
    or g33445 ( n22444 , n3765 , n27580 );
    or g33446 ( n13742 , n19682 , n27973 );
    xnor g33447 ( n25900 , n9792 , n16361 );
    xnor g33448 ( n27628 , n24410 , n4684 );
    and g33449 ( n9446 , n27026 , n5497 );
    xnor g33450 ( n26505 , n9937 , n9793 );
    not g33451 ( n19573 , n830 );
    or g33452 ( n16301 , n32171 , n16042 );
    or g33453 ( n13675 , n26614 , n18488 );
    or g33454 ( n18212 , n32095 , n1378 );
    or g33455 ( n24650 , n33250 , n21002 );
    or g33456 ( n18167 , n4288 , n23850 );
    or g33457 ( n5370 , n22684 , n19125 );
    or g33458 ( n27236 , n22618 , n4478 );
    xnor g33459 ( n29862 , n12944 , n31289 );
    and g33460 ( n20897 , n15549 , n8848 );
    or g33461 ( n6661 , n11574 , n31134 );
    xnor g33462 ( n33300 , n9639 , n32342 );
    xnor g33463 ( n10328 , n1451 , n17568 );
    xnor g33464 ( n31569 , n791 , n18495 );
    and g33465 ( n24777 , n23498 , n14870 );
    not g33466 ( n22041 , n18947 );
    and g33467 ( n21616 , n5132 , n399 );
    or g33468 ( n398 , n15886 , n6991 );
    nor g33469 ( n15124 , n28223 , n694 );
    nor g33470 ( n11479 , n32857 , n26584 );
    or g33471 ( n30632 , n11728 , n20812 );
    nor g33472 ( n21433 , n17568 , n1837 );
    xnor g33473 ( n31951 , n19821 , n2082 );
    or g33474 ( n16057 , n830 , n3050 );
    and g33475 ( n3071 , n21959 , n33895 );
    not g33476 ( n19295 , n8012 );
    xnor g33477 ( n5931 , n26312 , n830 );
    or g33478 ( n33926 , n13514 , n17612 );
    and g33479 ( n18760 , n28042 , n33350 );
    and g33480 ( n9380 , n11270 , n28714 );
    xnor g33481 ( n27644 , n176 , n15886 );
    xnor g33482 ( n35830 , n33220 , n15299 );
    or g33483 ( n5431 , n11282 , n13928 );
    or g33484 ( n20864 , n35162 , n5457 );
    or g33485 ( n2704 , n7540 , n33301 );
    and g33486 ( n34575 , n12492 , n23898 );
    or g33487 ( n22504 , n20418 , n35143 );
    xnor g33488 ( n20611 , n28137 , n24740 );
    nor g33489 ( n27400 , n147 , n13664 );
    and g33490 ( n20336 , n8297 , n19676 );
    or g33491 ( n23316 , n30833 , n6435 );
    not g33492 ( n20771 , n13019 );
    nor g33493 ( n27394 , n13473 , n28230 );
    and g33494 ( n15339 , n9577 , n31921 );
    or g33495 ( n15338 , n27969 , n32881 );
    and g33496 ( n18280 , n31358 , n25653 );
    or g33497 ( n27380 , n32584 , n32253 );
    nor g33498 ( n21092 , n30742 , n24442 );
    or g33499 ( n15937 , n28304 , n21034 );
    or g33500 ( n853 , n9793 , n12363 );
    or g33501 ( n6073 , n24600 , n4081 );
    xnor g33502 ( n31425 , n20572 , n24371 );
    not g33503 ( n9078 , n26907 );
    or g33504 ( n596 , n22555 , n22348 );
    xnor g33505 ( n28151 , n3917 , n32095 );
    nor g33506 ( n2174 , n956 , n21074 );
    or g33507 ( n31174 , n27933 , n32808 );
    and g33508 ( n28545 , n23501 , n14731 );
    xnor g33509 ( n10922 , n17117 , n17106 );
    and g33510 ( n23943 , n35133 , n30535 );
    not g33511 ( n25809 , n16247 );
    or g33512 ( n6798 , n5335 , n17304 );
    nor g33513 ( n21543 , n8980 , n18115 );
    or g33514 ( n8350 , n18159 , n35757 );
    xnor g33515 ( n16199 , n17083 , n24374 );
    or g33516 ( n24234 , n6125 , n30577 );
    and g33517 ( n31062 , n32044 , n27302 );
    or g33518 ( n2780 , n15793 , n30069 );
    and g33519 ( n14429 , n22576 , n33982 );
    or g33520 ( n31988 , n23044 , n31549 );
    xnor g33521 ( n16220 , n25084 , n15394 );
    and g33522 ( n7364 , n18866 , n24800 );
    or g33523 ( n7231 , n16001 , n17827 );
    or g33524 ( n27516 , n5477 , n33399 );
    not g33525 ( n11265 , n35949 );
    and g33526 ( n1370 , n22424 , n20236 );
    xnor g33527 ( n19838 , n10213 , n31289 );
    or g33528 ( n34410 , n13138 , n25927 );
    xnor g33529 ( n24235 , n34264 , n33294 );
    or g33530 ( n220 , n11893 , n23090 );
    or g33531 ( n6650 , n6072 , n33210 );
    not g33532 ( n842 , n18991 );
    or g33533 ( n31701 , n8432 , n6172 );
    or g33534 ( n12959 , n27487 , n9361 );
    or g33535 ( n6954 , n23212 , n11593 );
    or g33536 ( n12629 , n6539 , n10212 );
    or g33537 ( n716 , n15299 , n29666 );
    xnor g33538 ( n3918 , n23268 , n9480 );
    or g33539 ( n15387 , n34337 , n28191 );
    not g33540 ( n33746 , n4678 );
    not g33541 ( n20055 , n15377 );
    and g33542 ( n12987 , n3861 , n27219 );
    and g33543 ( n12724 , n31459 , n34436 );
    xnor g33544 ( n23508 , n15945 , n19576 );
    or g33545 ( n34093 , n35948 , n2955 );
    nor g33546 ( n7800 , n33439 , n16649 );
    xnor g33547 ( n8236 , n8697 , n16785 );
    nor g33548 ( n24670 , n1096 , n4697 );
    or g33549 ( n24084 , n35927 , n15066 );
    nor g33550 ( n31725 , n26063 , n27621 );
    or g33551 ( n1461 , n25020 , n12798 );
    xnor g33552 ( n6425 , n7325 , n30445 );
    or g33553 ( n32996 , n13315 , n32425 );
    and g33554 ( n28189 , n28327 , n16907 );
    or g33555 ( n23405 , n8776 , n9194 );
    or g33556 ( n4164 , n8377 , n35642 );
    or g33557 ( n27483 , n32336 , n19173 );
    or g33558 ( n35096 , n4749 , n17354 );
    or g33559 ( n3691 , n33298 , n23324 );
    nor g33560 ( n27537 , n26513 , n30755 );
    or g33561 ( n33672 , n7540 , n13672 );
    and g33562 ( n26747 , n13430 , n12004 );
    nor g33563 ( n4222 , n4962 , n7651 );
    or g33564 ( n32555 , n7623 , n33277 );
    xnor g33565 ( n32394 , n29363 , n23147 );
    or g33566 ( n254 , n10298 , n20526 );
    and g33567 ( n27980 , n4052 , n3478 );
    xnor g33568 ( n5535 , n23276 , n3222 );
    or g33569 ( n1517 , n27824 , n34865 );
    or g33570 ( n17550 , n14073 , n33416 );
    xnor g33571 ( n13885 , n18632 , n9195 );
    xnor g33572 ( n347 , n10876 , n15260 );
    and g33573 ( n28888 , n3061 , n35698 );
    or g33574 ( n5860 , n6124 , n7417 );
    and g33575 ( n35948 , n26373 , n32249 );
    xnor g33576 ( n856 , n1319 , n26740 );
    and g33577 ( n22519 , n21495 , n17649 );
    and g33578 ( n13425 , n30741 , n7905 );
    xnor g33579 ( n1691 , n22089 , n3004 );
    and g33580 ( n9015 , n2500 , n6716 );
    xnor g33581 ( n27039 , n35085 , n17568 );
    not g33582 ( n25778 , n29713 );
    or g33583 ( n3839 , n27978 , n22501 );
    xnor g33584 ( n14497 , n14597 , n32912 );
    and g33585 ( n32096 , n22520 , n32873 );
    and g33586 ( n24009 , n1449 , n25213 );
    or g33587 ( n10870 , n27771 , n28455 );
    xnor g33588 ( n24725 , n23574 , n9658 );
    xnor g33589 ( n25882 , n17563 , n816 );
    or g33590 ( n3697 , n27168 , n3805 );
    not g33591 ( n14277 , n11190 );
    or g33592 ( n34426 , n24371 , n20846 );
    not g33593 ( n7353 , n22471 );
    xnor g33594 ( n7658 , n34511 , n25411 );
    and g33595 ( n35978 , n24094 , n34059 );
    not g33596 ( n33885 , n28638 );
    or g33597 ( n16008 , n11481 , n10127 );
    xnor g33598 ( n14214 , n23822 , n5943 );
    not g33599 ( n3325 , n32209 );
    and g33600 ( n7944 , n33570 , n34787 );
    xnor g33601 ( n25429 , n8180 , n33063 );
    nor g33602 ( n35299 , n29713 , n24760 );
    xnor g33603 ( n19697 , n33643 , n8022 );
    or g33604 ( n4093 , n1827 , n8174 );
    and g33605 ( n31400 , n14130 , n6096 );
    nor g33606 ( n31482 , n13413 , n12367 );
    or g33607 ( n19798 , n15297 , n394 );
    xnor g33608 ( n35575 , n1052 , n6507 );
    or g33609 ( n34416 , n2048 , n16919 );
    xnor g33610 ( n9897 , n16731 , n3129 );
    or g33611 ( n15582 , n25105 , n30776 );
    and g33612 ( n688 , n16128 , n24870 );
    or g33613 ( n6218 , n6855 , n30489 );
    and g33614 ( n30130 , n15264 , n6904 );
    and g33615 ( n14379 , n11097 , n29169 );
    or g33616 ( n19361 , n4962 , n19874 );
    or g33617 ( n17334 , n18299 , n9015 );
    or g33618 ( n31915 , n31215 , n7867 );
    xnor g33619 ( n7704 , n8903 , n31272 );
    and g33620 ( n24840 , n7103 , n12576 );
    xnor g33621 ( n28337 , n7173 , n4878 );
    xnor g33622 ( n10638 , n19948 , n22859 );
    or g33623 ( n7659 , n22259 , n30024 );
    xnor g33624 ( n23359 , n16655 , n10744 );
    or g33625 ( n14088 , n30742 , n27070 );
    or g33626 ( n20923 , n8080 , n13305 );
    and g33627 ( n12088 , n27991 , n27413 );
    xnor g33628 ( n34855 , n1272 , n12602 );
    xnor g33629 ( n998 , n1150 , n13039 );
    and g33630 ( n35556 , n33754 , n12593 );
    not g33631 ( n2597 , n29203 );
    not g33632 ( n2693 , n23954 );
    xnor g33633 ( n14446 , n35024 , n21334 );
    xnor g33634 ( n31446 , n18414 , n12642 );
    and g33635 ( n11497 , n10848 , n21009 );
    and g33636 ( n20675 , n23576 , n13086 );
    and g33637 ( n2489 , n5319 , n20772 );
    or g33638 ( n6146 , n7583 , n11712 );
    and g33639 ( n35971 , n4082 , n21480 );
    xnor g33640 ( n31165 , n32625 , n31799 );
    not g33641 ( n33325 , n21434 );
    xnor g33642 ( n14381 , n20038 , n27177 );
    or g33643 ( n24418 , n25715 , n937 );
    or g33644 ( n18548 , n31272 , n1795 );
    and g33645 ( n1083 , n18292 , n32302 );
    or g33646 ( n19060 , n3946 , n12042 );
    xnor g33647 ( n28622 , n25575 , n31559 );
    or g33648 ( n33867 , n2628 , n16673 );
    and g33649 ( n22747 , n22596 , n34911 );
    or g33650 ( n29758 , n8943 , n28324 );
    or g33651 ( n33240 , n14423 , n26002 );
    and g33652 ( n16275 , n16680 , n11939 );
    or g33653 ( n21864 , n3205 , n35933 );
    xnor g33654 ( n31993 , n27746 , n23524 );
    not g33655 ( n32451 , n2030 );
    not g33656 ( n32932 , n11167 );
    or g33657 ( n35264 , n8150 , n21903 );
    xnor g33658 ( n28074 , n21304 , n28275 );
    or g33659 ( n17848 , n35703 , n31989 );
    and g33660 ( n31947 , n27348 , n30685 );
    and g33661 ( n24130 , n27079 , n33421 );
    or g33662 ( n30582 , n1492 , n26354 );
    and g33663 ( n32268 , n20018 , n1870 );
    xnor g33664 ( n1638 , n25766 , n18948 );
    xnor g33665 ( n4118 , n33198 , n96 );
    and g33666 ( n29185 , n25856 , n5957 );
    xnor g33667 ( n26585 , n10241 , n3679 );
    xnor g33668 ( n14233 , n28844 , n17876 );
    and g33669 ( n19786 , n27372 , n18729 );
    not g33670 ( n10581 , n17220 );
    or g33671 ( n29305 , n8070 , n2528 );
    xnor g33672 ( n10636 , n8438 , n24371 );
    or g33673 ( n6718 , n9430 , n35182 );
    xnor g33674 ( n4717 , n12840 , n15886 );
    or g33675 ( n18804 , n214 , n2384 );
    or g33676 ( n4323 , n35358 , n10336 );
    and g33677 ( n33473 , n9204 , n841 );
    or g33678 ( n9567 , n35672 , n19939 );
    or g33679 ( n9748 , n11546 , n13642 );
    or g33680 ( n2016 , n27876 , n29594 );
    and g33681 ( n25645 , n8859 , n33682 );
    or g33682 ( n26557 , n70 , n35900 );
    or g33683 ( n403 , n16620 , n34697 );
    xnor g33684 ( n30092 , n32567 , n32857 );
    nor g33685 ( n8096 , n4960 , n14584 );
    xnor g33686 ( n18943 , n8845 , n30742 );
    xnor g33687 ( n12111 , n1690 , n26562 );
    or g33688 ( n23616 , n30124 , n35143 );
    and g33689 ( n15754 , n10637 , n32876 );
    and g33690 ( n3548 , n5639 , n2602 );
    or g33691 ( n26160 , n10333 , n16893 );
    or g33692 ( n26781 , n23136 , n34518 );
    or g33693 ( n7126 , n755 , n17056 );
    xnor g33694 ( n380 , n18563 , n7421 );
    and g33695 ( n4523 , n7856 , n32640 );
    or g33696 ( n24575 , n3547 , n23790 );
    xnor g33697 ( n21143 , n32957 , n35440 );
    and g33698 ( n31786 , n16003 , n19885 );
    not g33699 ( n3298 , n10183 );
    or g33700 ( n2440 , n8031 , n26612 );
    or g33701 ( n6888 , n7944 , n2479 );
    not g33702 ( n32152 , n2734 );
    xnor g33703 ( n32627 , n1625 , n13608 );
    nor g33704 ( n6013 , n9793 , n25223 );
    or g33705 ( n20459 , n20659 , n8924 );
    not g33706 ( n10455 , n21146 );
    xnor g33707 ( n29955 , n29559 , n4288 );
    or g33708 ( n23693 , n24270 , n1756 );
    and g33709 ( n23245 , n26586 , n16856 );
    or g33710 ( n6000 , n33255 , n3144 );
    or g33711 ( n12539 , n23789 , n28248 );
    or g33712 ( n1329 , n4536 , n128 );
    xnor g33713 ( n32533 , n30314 , n28351 );
    or g33714 ( n14577 , n27675 , n2104 );
    not g33715 ( n14835 , n4962 );
    or g33716 ( n22476 , n329 , n35143 );
    and g33717 ( n15812 , n25371 , n29223 );
    or g33718 ( n28828 , n17938 , n13747 );
    or g33719 ( n23998 , n31558 , n13217 );
    and g33720 ( n34902 , n4420 , n13172 );
    or g33721 ( n26009 , n23091 , n3228 );
    and g33722 ( n18437 , n31234 , n21741 );
    not g33723 ( n26337 , n16620 );
    xnor g33724 ( n15292 , n13475 , n1133 );
    or g33725 ( n23096 , n20188 , n3694 );
    or g33726 ( n27914 , n11048 , n1642 );
    or g33727 ( n32358 , n25174 , n30967 );
    not g33728 ( n22350 , n33020 );
    or g33729 ( n15046 , n22892 , n20732 );
    or g33730 ( n10599 , n11501 , n6678 );
    and g33731 ( n4398 , n27154 , n9881 );
    or g33732 ( n19473 , n13562 , n17337 );
    xnor g33733 ( n12993 , n16194 , n7127 );
    or g33734 ( n28392 , n15996 , n2613 );
    nor g33735 ( n3092 , n16922 , n15150 );
    or g33736 ( n36066 , n7540 , n16107 );
    or g33737 ( n8249 , n14687 , n18193 );
    and g33738 ( n31190 , n2073 , n17780 );
    and g33739 ( n17877 , n31495 , n27706 );
    and g33740 ( n24150 , n31168 , n28436 );
    not g33741 ( n420 , n8299 );
    or g33742 ( n7606 , n13010 , n2104 );
    xnor g33743 ( n17856 , n32357 , n10643 );
    or g33744 ( n14690 , n28862 , n29148 );
    and g33745 ( n29194 , n5728 , n32233 );
    and g33746 ( n2138 , n23119 , n32238 );
    or g33747 ( n28281 , n26358 , n33475 );
    or g33748 ( n13986 , n9881 , n13649 );
    xnor g33749 ( n24521 , n5654 , n28926 );
    xnor g33750 ( n33540 , n2250 , n23419 );
    xnor g33751 ( n35701 , n27685 , n4350 );
    xnor g33752 ( n3907 , n6664 , n7192 );
    xnor g33753 ( n15842 , n8386 , n11190 );
    or g33754 ( n15765 , n20717 , n19336 );
    and g33755 ( n19836 , n17320 , n27364 );
    or g33756 ( n5462 , n24371 , n34618 );
    and g33757 ( n2128 , n8799 , n15974 );
    xnor g33758 ( n2055 , n6094 , n8432 );
    or g33759 ( n15401 , n30027 , n3437 );
    or g33760 ( n18997 , n27260 , n11850 );
    xnor g33761 ( n20219 , n20464 , n19 );
    or g33762 ( n4259 , n30297 , n31566 );
    xnor g33763 ( n23676 , n14067 , n11771 );
    or g33764 ( n19771 , n33586 , n10230 );
    or g33765 ( n15238 , n10706 , n5900 );
    nor g33766 ( n9911 , n29921 , n26157 );
    or g33767 ( n17913 , n27925 , n27625 );
    not g33768 ( n34231 , n21650 );
    nor g33769 ( n7000 , n9793 , n35493 );
    and g33770 ( n32468 , n7126 , n26798 );
    or g33771 ( n29857 , n4288 , n20395 );
    xnor g33772 ( n19471 , n1833 , n24371 );
    xnor g33773 ( n1355 , n27980 , n11455 );
    and g33774 ( n32898 , n20035 , n1513 );
    xnor g33775 ( n32375 , n19195 , n7270 );
    nor g33776 ( n11083 , n30767 , n6479 );
    and g33777 ( n20095 , n16368 , n11277 );
    and g33778 ( n11147 , n2206 , n11918 );
    or g33779 ( n14599 , n7584 , n24081 );
    or g33780 ( n24618 , n19551 , n32293 );
    xnor g33781 ( n25922 , n24892 , n16620 );
    or g33782 ( n21728 , n5157 , n17046 );
    or g33783 ( n26230 , n4783 , n36000 );
    xnor g33784 ( n7875 , n2034 , n31622 );
    or g33785 ( n2875 , n16337 , n28202 );
    nor g33786 ( n34561 , n18594 , n4254 );
    and g33787 ( n27308 , n14823 , n28128 );
    xnor g33788 ( n3249 , n30360 , n6308 );
    or g33789 ( n8862 , n21003 , n8924 );
    or g33790 ( n16204 , n29381 , n35935 );
    or g33791 ( n12812 , n24168 , n20579 );
    xnor g33792 ( n22803 , n27498 , n1317 );
    xnor g33793 ( n1288 , n12844 , n31559 );
    or g33794 ( n15174 , n24442 , n4912 );
    or g33795 ( n34090 , n24035 , n14918 );
    nor g33796 ( n31247 , n9658 , n3486 );
    or g33797 ( n25140 , n15066 , n27501 );
    and g33798 ( n13978 , n10084 , n29332 );
    or g33799 ( n13996 , n32859 , n19490 );
    or g33800 ( n30979 , n24037 , n17111 );
    or g33801 ( n2186 , n13863 , n24489 );
    xnor g33802 ( n20294 , n4447 , n10319 );
    and g33803 ( n31413 , n17245 , n19366 );
    and g33804 ( n26441 , n14568 , n7786 );
    not g33805 ( n1154 , n26262 );
    and g33806 ( n16750 , n24320 , n28293 );
    not g33807 ( n21146 , n30056 );
    and g33808 ( n13244 , n14443 , n2872 );
    or g33809 ( n30482 , n13875 , n9214 );
    and g33810 ( n27418 , n33547 , n17388 );
    and g33811 ( n8005 , n30075 , n17834 );
    or g33812 ( n6269 , n14858 , n12541 );
    xnor g33813 ( n5049 , n27688 , n29839 );
    not g33814 ( n24139 , n986 );
    xnor g33815 ( n5749 , n11862 , n20498 );
    xnor g33816 ( n23384 , n2608 , n29644 );
    not g33817 ( n9164 , n15886 );
    nor g33818 ( n3363 , n34853 , n8269 );
    xnor g33819 ( n33732 , n18436 , n929 );
    not g33820 ( n10983 , n3741 );
    or g33821 ( n32690 , n5612 , n949 );
    or g33822 ( n12454 , n26037 , n20601 );
    or g33823 ( n3904 , n21708 , n8891 );
    nor g33824 ( n1384 , n22330 , n2195 );
    and g33825 ( n8149 , n35554 , n4388 );
    or g33826 ( n11560 , n6406 , n13017 );
    or g33827 ( n19334 , n17961 , n13967 );
    or g33828 ( n11908 , n14782 , n3592 );
    xnor g33829 ( n25098 , n31682 , n15347 );
    or g33830 ( n20703 , n2061 , n9832 );
    or g33831 ( n35245 , n9793 , n20273 );
    or g33832 ( n35099 , n25274 , n20053 );
    or g33833 ( n31970 , n32133 , n14699 );
    or g33834 ( n27424 , n35767 , n12046 );
    or g33835 ( n11547 , n9588 , n10140 );
    xnor g33836 ( n24116 , n32520 , n30540 );
    or g33837 ( n28411 , n31559 , n19457 );
    and g33838 ( n9779 , n28573 , n11332 );
    and g33839 ( n3949 , n32723 , n29898 );
    nor g33840 ( n36026 , n30742 , n2690 );
    xnor g33841 ( n18908 , n13104 , n24371 );
    xnor g33842 ( n21866 , n23796 , n23930 );
    and g33843 ( n22788 , n16887 , n25413 );
    or g33844 ( n34932 , n30391 , n3842 );
    or g33845 ( n18900 , n345 , n13305 );
    xnor g33846 ( n23078 , n32804 , n23549 );
    and g33847 ( n26595 , n26284 , n27117 );
    and g33848 ( n17966 , n8266 , n17232 );
    or g33849 ( n24693 , n25602 , n31702 );
    xnor g33850 ( n12655 , n20689 , n29977 );
    xnor g33851 ( n30366 , n23070 , n19710 );
    or g33852 ( n32760 , n8311 , n2817 );
    xnor g33853 ( n12519 , n34510 , n33691 );
    buf g33854 ( n30204 , n34425 );
    or g33855 ( n15180 , n7971 , n34084 );
    and g33856 ( n12458 , n22949 , n18716 );
    or g33857 ( n21204 , n15827 , n16457 );
    xnor g33858 ( n17518 , n12312 , n31653 );
    and g33859 ( n548 , n11103 , n18704 );
    and g33860 ( n8244 , n29772 , n19713 );
    xnor g33861 ( n13351 , n15688 , n21450 );
    or g33862 ( n27188 , n27612 , n1437 );
    xnor g33863 ( n7379 , n35465 , n5287 );
    nor g33864 ( n30260 , n26862 , n4941 );
    nor g33865 ( n22885 , n20468 , n31411 );
    xnor g33866 ( n11186 , n21273 , n8833 );
    buf g33867 ( n9361 , n22761 );
    or g33868 ( n20249 , n20714 , n17430 );
    or g33869 ( n9932 , n4962 , n18632 );
    xnor g33870 ( n35455 , n2334 , n24517 );
    nor g33871 ( n31003 , n5335 , n31881 );
    or g33872 ( n6308 , n6289 , n34670 );
    xnor g33873 ( n9837 , n14281 , n27226 );
    xnor g33874 ( n31314 , n16761 , n26965 );
    nor g33875 ( n31578 , n18844 , n25444 );
    or g33876 ( n340 , n2393 , n11593 );
    xnor g33877 ( n1654 , n35362 , n31565 );
    nor g33878 ( n2275 , n14500 , n3458 );
    xnor g33879 ( n35408 , n19434 , n5587 );
    nor g33880 ( n5669 , n17751 , n29185 );
    xnor g33881 ( n24171 , n30064 , n28743 );
    or g33882 ( n5897 , n28211 , n1176 );
    nor g33883 ( n288 , n9873 , n25458 );
    or g33884 ( n24209 , n33015 , n4595 );
    or g33885 ( n24771 , n1862 , n5675 );
    nor g33886 ( n7882 , n16909 , n16649 );
    or g33887 ( n1822 , n35395 , n139 );
    and g33888 ( n10229 , n6903 , n23273 );
    or g33889 ( n34360 , n776 , n3634 );
    xnor g33890 ( n25002 , n28022 , n30109 );
    xnor g33891 ( n11528 , n11653 , n8104 );
    or g33892 ( n8289 , n31586 , n14918 );
    or g33893 ( n8673 , n26666 , n33140 );
    xnor g33894 ( n4698 , n18341 , n8197 );
    or g33895 ( n891 , n10800 , n5274 );
    or g33896 ( n29219 , n35363 , n26468 );
    or g33897 ( n28516 , n35239 , n11518 );
    or g33898 ( n20124 , n7540 , n28830 );
    and g33899 ( n31710 , n16506 , n9334 );
    xnor g33900 ( n988 , n1510 , n1103 );
    or g33901 ( n26886 , n30114 , n19421 );
    or g33902 ( n33409 , n23244 , n27801 );
    and g33903 ( n995 , n6597 , n27507 );
    or g33904 ( n28955 , n21570 , n24118 );
    nor g33905 ( n23335 , n16302 , n29203 );
    xnor g33906 ( n5702 , n7996 , n10781 );
    or g33907 ( n19780 , n119 , n12791 );
    or g33908 ( n8867 , n24889 , n29138 );
    or g33909 ( n4747 , n36086 , n28548 );
    or g33910 ( n7635 , n33301 , n25447 );
    xnor g33911 ( n8129 , n5623 , n4288 );
    or g33912 ( n34263 , n16521 , n20371 );
    or g33913 ( n7518 , n998 , n31464 );
    or g33914 ( n16150 , n1601 , n8909 );
    or g33915 ( n20545 , n27209 , n36088 );
    not g33916 ( n34714 , n21923 );
    or g33917 ( n30651 , n22169 , n9555 );
    or g33918 ( n32018 , n5841 , n25594 );
    xnor g33919 ( n27572 , n32463 , n20966 );
    or g33920 ( n31837 , n30467 , n16961 );
    or g33921 ( n4703 , n4975 , n1454 );
    or g33922 ( n21919 , n23751 , n17731 );
    or g33923 ( n3874 , n1725 , n24025 );
    and g33924 ( n25948 , n31396 , n2843 );
    nor g33925 ( n18707 , n26027 , n6160 );
    and g33926 ( n3583 , n19644 , n34077 );
    not g33927 ( n8567 , n6417 );
    xnor g33928 ( n3613 , n34463 , n4960 );
    not g33929 ( n2326 , n4960 );
    or g33930 ( n9968 , n21245 , n388 );
    not g33931 ( n4192 , n15222 );
    xnor g33932 ( n17800 , n10030 , n26371 );
    not g33933 ( n29476 , n2885 );
    or g33934 ( n18519 , n26423 , n27501 );
    and g33935 ( n3501 , n15205 , n17739 );
    or g33936 ( n14377 , n17950 , n2323 );
    not g33937 ( n20749 , n34923 );
    or g33938 ( n28476 , n29794 , n6837 );
    xnor g33939 ( n17580 , n8742 , n15756 );
    not g33940 ( n22561 , n34643 );
    xnor g33941 ( n7746 , n1598 , n9642 );
    nor g33942 ( n3350 , n16620 , n3157 );
    or g33943 ( n10963 , n20366 , n4675 );
    xnor g33944 ( n3137 , n8513 , n31397 );
    or g33945 ( n32308 , n18620 , n3185 );
    xnor g33946 ( n1928 , n18795 , n16620 );
    or g33947 ( n6105 , n18361 , n10289 );
    and g33948 ( n32235 , n7705 , n31272 );
    xnor g33949 ( n2308 , n20158 , n23157 );
    and g33950 ( n4972 , n20624 , n33900 );
    xnor g33951 ( n9544 , n12885 , n30462 );
    or g33952 ( n82 , n21716 , n5972 );
    or g33953 ( n26187 , n31091 , n25281 );
    nor g33954 ( n14981 , n25602 , n21029 );
    nor g33955 ( n30744 , n28889 , n18115 );
    and g33956 ( n34331 , n34000 , n3436 );
    or g33957 ( n23228 , n11905 , n35593 );
    or g33958 ( n35396 , n31193 , n25019 );
    and g33959 ( n29306 , n20281 , n19978 );
    and g33960 ( n29059 , n2783 , n35564 );
    or g33961 ( n31597 , n9789 , n24624 );
    or g33962 ( n6899 , n21404 , n32425 );
    or g33963 ( n21593 , n2040 , n15215 );
    or g33964 ( n21689 , n28908 , n10872 );
    or g33965 ( n29406 , n993 , n22499 );
    nor g33966 ( n25198 , n25897 , n1342 );
    or g33967 ( n17138 , n11206 , n34727 );
    and g33968 ( n23414 , n11298 , n2009 );
    and g33969 ( n17405 , n4671 , n29936 );
    and g33970 ( n15198 , n29846 , n30597 );
    xnor g33971 ( n8180 , n29967 , n4758 );
    and g33972 ( n34379 , n601 , n22735 );
    and g33973 ( n7184 , n27007 , n27001 );
    xnor g33974 ( n18216 , n13622 , n6292 );
    or g33975 ( n6023 , n2905 , n24008 );
    or g33976 ( n23598 , n22022 , n1474 );
    nor g33977 ( n15283 , n14275 , n33157 );
    xnor g33978 ( n22643 , n31141 , n5080 );
    or g33979 ( n9540 , n17766 , n27310 );
    or g33980 ( n31095 , n23169 , n25392 );
    xnor g33981 ( n12138 , n20299 , n10642 );
    nor g33982 ( n25945 , n18472 , n9921 );
    or g33983 ( n7574 , n25645 , n8392 );
    or g33984 ( n32786 , n4578 , n12913 );
    xnor g33985 ( n18345 , n18422 , n13669 );
    xnor g33986 ( n17971 , n1770 , n15423 );
    or g33987 ( n15346 , n15886 , n32997 );
    and g33988 ( n2099 , n19585 , n20968 );
    xnor g33989 ( n6781 , n12108 , n31733 );
    or g33990 ( n15815 , n14449 , n11295 );
    or g33991 ( n34655 , n575 , n10432 );
    xnor g33992 ( n20320 , n20015 , n35716 );
    not g33993 ( n12511 , n26365 );
    or g33994 ( n26836 , n23542 , n1050 );
    or g33995 ( n12970 , n35219 , n3842 );
    or g33996 ( n29380 , n32265 , n25761 );
    not g33997 ( n10577 , n2792 );
    or g33998 ( n7886 , n34690 , n16668 );
    xnor g33999 ( n14484 , n23817 , n6638 );
    or g34000 ( n13202 , n31215 , n34172 );
    or g34001 ( n34240 , n31027 , n22916 );
    xnor g34002 ( n4824 , n22274 , n19158 );
    or g34003 ( n960 , n7894 , n25392 );
    xnor g34004 ( n23038 , n8459 , n22102 );
    and g34005 ( n25918 , n10685 , n6382 );
    and g34006 ( n20418 , n6237 , n22930 );
    or g34007 ( n9248 , n30800 , n18264 );
    and g34008 ( n28887 , n2777 , n15366 );
    xnor g34009 ( n10604 , n16212 , n8432 );
    nor g34010 ( n18307 , n10669 , n23297 );
    xnor g34011 ( n23208 , n12934 , n16690 );
    or g34012 ( n7139 , n8783 , n27727 );
    or g34013 ( n13487 , n29495 , n10765 );
    or g34014 ( n29091 , n30130 , n9317 );
    xnor g34015 ( n4165 , n22735 , n601 );
    and g34016 ( n29050 , n4736 , n25004 );
    or g34017 ( n20632 , n25256 , n5779 );
    xnor g34018 ( n5942 , n9500 , n8432 );
    not g34019 ( n11678 , n16922 );
    or g34020 ( n4589 , n16528 , n20579 );
    xnor g34021 ( n20349 , n24715 , n4934 );
    and g34022 ( n2303 , n5367 , n15783 );
    or g34023 ( n4802 , n26168 , n31067 );
    or g34024 ( n32830 , n23604 , n33812 );
    or g34025 ( n11689 , n34921 , n25594 );
    xnor g34026 ( n17517 , n25606 , n16141 );
    or g34027 ( n21024 , n7183 , n21955 );
    xnor g34028 ( n35911 , n35075 , n7184 );
    or g34029 ( n21595 , n8110 , n19732 );
    and g34030 ( n26453 , n18091 , n779 );
    or g34031 ( n20868 , n21360 , n544 );
    or g34032 ( n20415 , n29839 , n12334 );
    not g34033 ( n28223 , n4542 );
    or g34034 ( n16783 , n33554 , n32257 );
    or g34035 ( n32181 , n21532 , n27447 );
    or g34036 ( n7044 , n6423 , n4175 );
    or g34037 ( n27475 , n3370 , n12961 );
    xnor g34038 ( n11300 , n8775 , n25602 );
    or g34039 ( n33393 , n19694 , n33416 );
    and g34040 ( n9923 , n21620 , n28418 );
    or g34041 ( n17850 , n16922 , n9380 );
    nor g34042 ( n13735 , n15580 , n24967 );
    and g34043 ( n11617 , n17287 , n7933 );
    not g34044 ( n11990 , n16620 );
    or g34045 ( n26310 , n18130 , n25786 );
    and g34046 ( n24118 , n29638 , n33394 );
    and g34047 ( n9899 , n11269 , n16293 );
    buf g34048 ( n31554 , n21785 );
    xnor g34049 ( n25779 , n8012 , n34943 );
    or g34050 ( n31877 , n3783 , n23790 );
    xnor g34051 ( n17588 , n23045 , n31799 );
    nor g34052 ( n3960 , n4960 , n19991 );
    xnor g34053 ( n36010 , n15537 , n9658 );
    or g34054 ( n19729 , n5335 , n15924 );
    xnor g34055 ( n24258 , n20453 , n17568 );
    xnor g34056 ( n20945 , n680 , n14997 );
    buf g34057 ( n34727 , n11773 );
    not g34058 ( n1382 , n9899 );
    and g34059 ( n6127 , n17165 , n17994 );
    and g34060 ( n1649 , n8460 , n34405 );
    xnor g34061 ( n13759 , n16538 , n18554 );
    xor g34062 ( n7652 , n26609 , n32857 );
    nor g34063 ( n8328 , n10989 , n32366 );
    not g34064 ( n30126 , n9789 );
    or g34065 ( n21249 , n17637 , n2168 );
    or g34066 ( n14490 , n5738 , n6992 );
    or g34067 ( n33057 , n1609 , n22470 );
    or g34068 ( n35426 , n9467 , n32425 );
    and g34069 ( n13454 , n17979 , n28992 );
    xnor g34070 ( n18538 , n19532 , n27291 );
    and g34071 ( n33670 , n9420 , n20367 );
    or g34072 ( n4289 , n13073 , n2950 );
    xnor g34073 ( n12417 , n1140 , n5588 );
    and g34074 ( n3167 , n162 , n24377 );
    or g34075 ( n1159 , n1634 , n6459 );
    xnor g34076 ( n25531 , n3463 , n17568 );
    or g34077 ( n17490 , n35746 , n22316 );
    nor g34078 ( n7324 , n3222 , n28554 );
    nor g34079 ( n29870 , n5424 , n9099 );
    not g34080 ( n1926 , n32812 );
    buf g34081 ( n25255 , n32167 );
    and g34082 ( n839 , n18592 , n33504 );
    or g34083 ( n34961 , n15752 , n35111 );
    or g34084 ( n12505 , n22291 , n18558 );
    or g34085 ( n22956 , n427 , n13900 );
    or g34086 ( n8986 , n16741 , n30433 );
    and g34087 ( n4995 , n32904 , n22307 );
    and g34088 ( n17951 , n2923 , n29005 );
    or g34089 ( n10518 , n10317 , n25255 );
    or g34090 ( n5293 , n24194 , n32697 );
    or g34091 ( n13079 , n25602 , n31675 );
    not g34092 ( n21252 , n32832 );
    or g34093 ( n10857 , n21636 , n12481 );
    or g34094 ( n11519 , n24909 , n16464 );
    xnor g34095 ( n4409 , n16626 , n35040 );
    and g34096 ( n22351 , n7469 , n18815 );
    and g34097 ( n32574 , n25564 , n22980 );
    not g34098 ( n26896 , n9658 );
    or g34099 ( n31348 , n16620 , n29595 );
    xnor g34100 ( n21242 , n36010 , n14938 );
    and g34101 ( n28206 , n33233 , n34357 );
    and g34102 ( n32589 , n16484 , n8280 );
    nor g34103 ( n2396 , n19551 , n18220 );
    or g34104 ( n23396 , n17468 , n17544 );
    not g34105 ( n18634 , n3450 );
    nor g34106 ( n19465 , n28563 , n27053 );
    nor g34107 ( n13083 , n26455 , n2706 );
    or g34108 ( n28249 , n16926 , n27678 );
    or g34109 ( n24883 , n11426 , n27447 );
    and g34110 ( n6402 , n8279 , n9282 );
    and g34111 ( n14009 , n7695 , n14544 );
    or g34112 ( n17649 , n29839 , n3822 );
    or g34113 ( n35192 , n9819 , n31566 );
    not g34114 ( n10185 , n30360 );
    or g34115 ( n7613 , n6616 , n34250 );
    or g34116 ( n19486 , n10328 , n2473 );
    or g34117 ( n32236 , n23189 , n4081 );
    nor g34118 ( n9197 , n560 , n33157 );
    and g34119 ( n11823 , n1249 , n26933 );
    or g34120 ( n6130 , n12817 , n5618 );
    nor g34121 ( n19600 , n8305 , n21434 );
    or g34122 ( n30166 , n30471 , n1264 );
    or g34123 ( n2602 , n19791 , n30646 );
    or g34124 ( n5714 , n6176 , n31549 );
    and g34125 ( n7032 , n9119 , n19937 );
    xnor g34126 ( n20543 , n14763 , n28592 );
    xnor g34127 ( n25938 , n26792 , n33764 );
    and g34128 ( n20977 , n27044 , n3084 );
    or g34129 ( n24827 , n17161 , n3188 );
    and g34130 ( n11648 , n8880 , n21111 );
    xnor g34131 ( n19822 , n19545 , n34591 );
    and g34132 ( n3604 , n20625 , n20391 );
    and g34133 ( n24422 , n15983 , n22660 );
    or g34134 ( n7431 , n31423 , n33808 );
    and g34135 ( n5478 , n25303 , n20679 );
    xnor g34136 ( n35522 , n1478 , n17223 );
    or g34137 ( n11119 , n15603 , n8392 );
    nor g34138 ( n31185 , n4962 , n31412 );
    not g34139 ( n7175 , n22200 );
    xnor g34140 ( n9810 , n5144 , n23633 );
    or g34141 ( n6575 , n5067 , n18525 );
    xnor g34142 ( n2093 , n26358 , n33475 );
    xnor g34143 ( n25731 , n15875 , n25174 );
    xnor g34144 ( n22937 , n22838 , n2932 );
    xnor g34145 ( n22447 , n7074 , n31215 );
    xnor g34146 ( n33613 , n33372 , n21508 );
    or g34147 ( n7723 , n25973 , n24479 );
    or g34148 ( n33339 , n17390 , n3736 );
    and g34149 ( n9862 , n12210 , n9169 );
    or g34150 ( n9595 , n32241 , n34437 );
    xnor g34151 ( n1169 , n16092 , n26057 );
    or g34152 ( n1361 , n32290 , n1942 );
    and g34153 ( n6212 , n28205 , n29714 );
    or g34154 ( n35842 , n32715 , n7587 );
    xnor g34155 ( n10353 , n30108 , n6737 );
    nor g34156 ( n4330 , n29152 , n20701 );
    or g34157 ( n28235 , n22261 , n28064 );
    and g34158 ( n18710 , n11462 , n8402 );
    and g34159 ( n10028 , n33264 , n9886 );
    xnor g34160 ( n11620 , n7888 , n32095 );
    and g34161 ( n6764 , n13682 , n35758 );
    and g34162 ( n13368 , n11380 , n3589 );
    xnor g34163 ( n6482 , n33728 , n32857 );
    and g34164 ( n25701 , n3051 , n8403 );
    nor g34165 ( n1628 , n25174 , n18534 );
    buf g34166 ( n11833 , n34963 );
    or g34167 ( n5176 , n8217 , n25594 );
    xnor g34168 ( n9524 , n21496 , n17751 );
    not g34169 ( n5200 , n24371 );
    or g34170 ( n4022 , n34769 , n29411 );
    nor g34171 ( n30065 , n22336 , n31411 );
    xnor g34172 ( n8140 , n32370 , n19551 );
    or g34173 ( n4994 , n18359 , n27276 );
    xnor g34174 ( n3765 , n29484 , n1928 );
    or g34175 ( n6071 , n10517 , n9591 );
    xnor g34176 ( n4923 , n30665 , n17568 );
    xor g34177 ( n25829 , n33428 , n13553 );
    or g34178 ( n29043 , n10791 , n25106 );
    xnor g34179 ( n750 , n21452 , n15886 );
    and g34180 ( n33443 , n22172 , n25222 );
    or g34181 ( n25261 , n22371 , n8924 );
    xnor g34182 ( n31985 , n27521 , n27735 );
    and g34183 ( n26745 , n552 , n28840 );
    xnor g34184 ( n6694 , n1563 , n33420 );
    not g34185 ( n13523 , n2433 );
    or g34186 ( n10672 , n1328 , n30504 );
    or g34187 ( n724 , n5748 , n15753 );
    xnor g34188 ( n3972 , n3548 , n9793 );
    xnor g34189 ( n19378 , n3974 , n669 );
    xnor g34190 ( n408 , n25839 , n15299 );
    and g34191 ( n23101 , n372 , n2617 );
    xnor g34192 ( n23979 , n25948 , n12787 );
    and g34193 ( n9543 , n33600 , n4953 );
    or g34194 ( n20133 , n1653 , n12853 );
    not g34195 ( n11699 , n34824 );
    xnor g34196 ( n32876 , n8187 , n24192 );
    or g34197 ( n8971 , n830 , n27870 );
    or g34198 ( n5966 , n20408 , n33489 );
    nor g34199 ( n31532 , n3294 , n13647 );
    xnor g34200 ( n34846 , n4710 , n31289 );
    or g34201 ( n4909 , n31821 , n4363 );
    and g34202 ( n16016 , n32172 , n26605 );
    and g34203 ( n834 , n5232 , n35684 );
    or g34204 ( n22181 , n23432 , n20854 );
    xnor g34205 ( n14450 , n7129 , n28672 );
    or g34206 ( n19854 , n13771 , n30476 );
    or g34207 ( n16983 , n3223 , n6683 );
    or g34208 ( n15845 , n21699 , n19421 );
    or g34209 ( n14852 , n10213 , n25023 );
    xnor g34210 ( n8239 , n24432 , n7544 );
    nor g34211 ( n35542 , n830 , n18923 );
    xnor g34212 ( n438 , n35202 , n18332 );
    or g34213 ( n16140 , n17258 , n25392 );
    or g34214 ( n24440 , n9658 , n2657 );
    not g34215 ( n15735 , n31599 );
    not g34216 ( n4267 , n6890 );
    or g34217 ( n9959 , n15398 , n29626 );
    xnor g34218 ( n28750 , n4141 , n16744 );
    xor g34219 ( n13386 , n8267 , n25991 );
    xnor g34220 ( n31450 , n25118 , n26879 );
    xnor g34221 ( n26377 , n26539 , n35832 );
    or g34222 ( n27507 , n32095 , n7793 );
    buf g34223 ( n30419 , n26962 );
    xnor g34224 ( n12407 , n35801 , n4960 );
    and g34225 ( n35157 , n12871 , n4458 );
    or g34226 ( n5928 , n34238 , n2977 );
    or g34227 ( n13841 , n32704 , n7776 );
    and g34228 ( n31577 , n33211 , n6924 );
    or g34229 ( n17846 , n19551 , n31781 );
    and g34230 ( n32351 , n27189 , n30491 );
    or g34231 ( n27272 , n6481 , n22663 );
    not g34232 ( n34888 , n9361 );
    and g34233 ( n7645 , n12959 , n9635 );
    or g34234 ( n33568 , n25629 , n26002 );
    or g34235 ( n366 , n5335 , n21232 );
    and g34236 ( n11683 , n33954 , n17084 );
    or g34237 ( n10446 , n32095 , n1524 );
    nor g34238 ( n33906 , n21424 , n13074 );
    xnor g34239 ( n34324 , n22814 , n27226 );
    or g34240 ( n25525 , n1086 , n24479 );
    and g34241 ( n33105 , n30454 , n22358 );
    or g34242 ( n30058 , n29442 , n12428 );
    nor g34243 ( n7444 , n14339 , n11666 );
    xnor g34244 ( n5154 , n33967 , n3489 );
    or g34245 ( n5500 , n1020 , n12879 );
    or g34246 ( n30712 , n19178 , n5465 );
    and g34247 ( n3537 , n8908 , n21140 );
    or g34248 ( n19254 , n31559 , n20592 );
    buf g34249 ( n20812 , n21971 );
    nor g34250 ( n1231 , n9793 , n33458 );
    and g34251 ( n15006 , n9729 , n16427 );
    not g34252 ( n26549 , n22471 );
    not g34253 ( n13245 , n20558 );
    or g34254 ( n5352 , n17643 , n20762 );
    xnor g34255 ( n28875 , n502 , n26458 );
    nor g34256 ( n5482 , n13159 , n29432 );
    or g34257 ( n10186 , n31799 , n17722 );
    or g34258 ( n33314 , n10839 , n10400 );
    and g34259 ( n11848 , n2200 , n34239 );
    or g34260 ( n23560 , n30139 , n24356 );
    xnor g34261 ( n28760 , n22042 , n30627 );
    nor g34262 ( n9063 , n23604 , n12400 );
    and g34263 ( n3228 , n35759 , n6138 );
    not g34264 ( n31924 , n16808 );
    or g34265 ( n20424 , n5287 , n9355 );
    or g34266 ( n5529 , n8714 , n18090 );
    not g34267 ( n1260 , n4288 );
    nor g34268 ( n11008 , n29839 , n22747 );
    and g34269 ( n33433 , n16322 , n32453 );
    xnor g34270 ( n7396 , n17901 , n24371 );
    and g34271 ( n25445 , n31379 , n11986 );
    nor g34272 ( n2096 , n3205 , n3992 );
    xnor g34273 ( n31017 , n4176 , n29839 );
    and g34274 ( n29692 , n26839 , n22912 );
    and g34275 ( n20958 , n22367 , n19877 );
    nor g34276 ( n22262 , n1836 , n6859 );
    or g34277 ( n3524 , n25088 , n11218 );
    xnor g34278 ( n11059 , n9339 , n30699 );
    and g34279 ( n10488 , n34095 , n29046 );
    and g34280 ( n24663 , n27593 , n15858 );
    nor g34281 ( n34583 , n25637 , n5637 );
    or g34282 ( n9203 , n28808 , n27501 );
    xnor g34283 ( n31238 , n12639 , n30010 );
    or g34284 ( n9089 , n27411 , n7553 );
    or g34285 ( n27702 , n20008 , n4792 );
    or g34286 ( n12779 , n14721 , n2782 );
    nor g34287 ( n3170 , n35927 , n23500 );
    xnor g34288 ( n12771 , n30132 , n32095 );
    or g34289 ( n12800 , n21488 , n34537 );
    and g34290 ( n16548 , n11053 , n30533 );
    or g34291 ( n32712 , n1619 , n13480 );
    or g34292 ( n981 , n24114 , n11823 );
    xnor g34293 ( n34866 , n10988 , n9443 );
    and g34294 ( n13777 , n18078 , n10092 );
    or g34295 ( n27579 , n28399 , n16751 );
    or g34296 ( n26130 , n3058 , n31541 );
    xnor g34297 ( n4115 , n27237 , n18301 );
    and g34298 ( n21902 , n8941 , n19709 );
    xnor g34299 ( n2189 , n28021 , n3205 );
    or g34300 ( n29105 , n10422 , n22350 );
    and g34301 ( n28143 , n21575 , n11118 );
    and g34302 ( n27169 , n645 , n22860 );
    or g34303 ( n19339 , n31762 , n2814 );
    or g34304 ( n27591 , n35927 , n26823 );
    or g34305 ( n3266 , n13366 , n17877 );
    and g34306 ( n1158 , n29803 , n20415 );
    xor g34307 ( n10070 , n27343 , n9994 );
    or g34308 ( n2285 , n13188 , n23462 );
    nor g34309 ( n10239 , n10894 , n25228 );
    xnor g34310 ( n34725 , n10945 , n4065 );
    xnor g34311 ( n32074 , n27594 , n33618 );
    and g34312 ( n29288 , n30684 , n26096 );
    or g34313 ( n34649 , n29143 , n27491 );
    xnor g34314 ( n5101 , n22922 , n4561 );
    nor g34315 ( n26172 , n4232 , n27484 );
    or g34316 ( n35243 , n16485 , n15344 );
    or g34317 ( n33045 , n29611 , n128 );
    or g34318 ( n16969 , n12835 , n36000 );
    or g34319 ( n25010 , n32433 , n28260 );
    or g34320 ( n30758 , n16788 , n11952 );
    xnor g34321 ( n5410 , n973 , n16724 );
    xnor g34322 ( n12242 , n2154 , n1569 );
    xnor g34323 ( n23945 , n6653 , n30193 );
    xnor g34324 ( n6351 , n11195 , n2095 );
    and g34325 ( n14592 , n6635 , n13555 );
    or g34326 ( n1548 , n35486 , n26292 );
    or g34327 ( n24288 , n24371 , n21108 );
    xnor g34328 ( n16530 , n15964 , n35185 );
    and g34329 ( n2335 , n4299 , n35686 );
    or g34330 ( n327 , n8525 , n28455 );
    or g34331 ( n27517 , n2103 , n34727 );
    xnor g34332 ( n35375 , n2379 , n5905 );
    and g34333 ( n28393 , n12682 , n14248 );
    or g34334 ( n16455 , n8583 , n31134 );
    nor g34335 ( n35359 , n15605 , n4508 );
    and g34336 ( n22002 , n15271 , n8509 );
    xnor g34337 ( n6656 , n11521 , n15604 );
    and g34338 ( n28550 , n28496 , n21300 );
    or g34339 ( n28910 , n15649 , n13217 );
    or g34340 ( n9119 , n17586 , n17681 );
    or g34341 ( n16683 , n20596 , n4318 );
    or g34342 ( n2315 , n18776 , n25678 );
    and g34343 ( n32354 , n27826 , n27233 );
    or g34344 ( n7705 , n16100 , n35427 );
    or g34345 ( n1121 , n14601 , n22328 );
    or g34346 ( n34147 , n21470 , n23921 );
    xnor g34347 ( n19760 , n17295 , n27108 );
    or g34348 ( n33215 , n24483 , n614 );
    and g34349 ( n6761 , n25571 , n24470 );
    or g34350 ( n2026 , n32109 , n22961 );
    or g34351 ( n33714 , n12363 , n11833 );
    not g34352 ( n27359 , n7588 );
    and g34353 ( n584 , n13752 , n15243 );
    and g34354 ( n7427 , n16196 , n20619 );
    xnor g34355 ( n29333 , n28337 , n27827 );
    and g34356 ( n11237 , n17848 , n10742 );
    or g34357 ( n21008 , n25289 , n1402 );
    nor g34358 ( n12298 , n18443 , n12879 );
    and g34359 ( n22691 , n14819 , n15041 );
    or g34360 ( n12239 , n33525 , n908 );
    nor g34361 ( n33871 , n20942 , n26282 );
    and g34362 ( n25343 , n8336 , n28718 );
    not g34363 ( n8057 , n34952 );
    xnor g34364 ( n3147 , n7301 , n23147 );
    or g34365 ( n3986 , n23092 , n16837 );
    and g34366 ( n8513 , n4048 , n271 );
    and g34367 ( n23419 , n29972 , n2699 );
    nor g34368 ( n15279 , n29492 , n15138 );
    or g34369 ( n3853 , n11644 , n34971 );
    and g34370 ( n23086 , n35402 , n32637 );
    or g34371 ( n30281 , n5287 , n35916 );
    or g34372 ( n35997 , n796 , n7726 );
    or g34373 ( n27659 , n35930 , n13564 );
    or g34374 ( n34684 , n2610 , n24333 );
    or g34375 ( n4873 , n13862 , n9675 );
    or g34376 ( n9739 , n20563 , n5634 );
    not g34377 ( n30624 , n16436 );
    or g34378 ( n2761 , n8307 , n27728 );
    xnor g34379 ( n32522 , n6031 , n35589 );
    or g34380 ( n17497 , n13603 , n14706 );
    not g34381 ( n19306 , n33435 );
    or g34382 ( n31907 , n33868 , n1350 );
    not g34383 ( n10944 , n1786 );
    not g34384 ( n22924 , n22667 );
    or g34385 ( n12609 , n23585 , n28952 );
    or g34386 ( n16625 , n1935 , n9553 );
    xnor g34387 ( n1254 , n1498 , n1156 );
    or g34388 ( n19110 , n7683 , n34084 );
    and g34389 ( n14224 , n33568 , n1178 );
    or g34390 ( n32374 , n3946 , n30124 );
    or g34391 ( n29679 , n9366 , n15169 );
    and g34392 ( n33652 , n14752 , n7405 );
    or g34393 ( n22490 , n23470 , n35043 );
    xnor g34394 ( n16879 , n22700 , n7540 );
    xnor g34395 ( n31807 , n19050 , n16922 );
    and g34396 ( n29302 , n16867 , n28786 );
    xnor g34397 ( n1658 , n16180 , n15403 );
    or g34398 ( n23479 , n30173 , n16543 );
    or g34399 ( n16106 , n22291 , n31433 );
    xnor g34400 ( n30440 , n31976 , n1069 );
    and g34401 ( n13745 , n32118 , n5202 );
    nor g34402 ( n14365 , n4345 , n26342 );
    or g34403 ( n34594 , n35261 , n16919 );
    and g34404 ( n33758 , n33620 , n7539 );
    or g34405 ( n20791 , n6652 , n33689 );
    or g34406 ( n32810 , n25511 , n26646 );
    not g34407 ( n16557 , n14742 );
    or g34408 ( n6343 , n31215 , n25984 );
    and g34409 ( n15143 , n24416 , n10443 );
    or g34410 ( n8397 , n7342 , n2712 );
    or g34411 ( n294 , n16316 , n14361 );
    nor g34412 ( n34709 , n31799 , n28717 );
    buf g34413 ( n1715 , n33469 );
    xnor g34414 ( n27632 , n9923 , n33353 );
    or g34415 ( n19431 , n13686 , n23921 );
    xnor g34416 ( n14735 , n22599 , n30418 );
    or g34417 ( n5903 , n3222 , n35057 );
    or g34418 ( n9299 , n9961 , n30646 );
    xnor g34419 ( n31612 , n25109 , n33344 );
    or g34420 ( n9788 , n31289 , n16016 );
    not g34421 ( n29296 , n25602 );
    or g34422 ( n32513 , n31571 , n30595 );
    or g34423 ( n34624 , n18965 , n25592 );
    or g34424 ( n14005 , n9789 , n14709 );
    or g34425 ( n14229 , n17652 , n27196 );
    not g34426 ( n8179 , n3946 );
    xnor g34427 ( n2762 , n6701 , n17751 );
    xnor g34428 ( n17536 , n1288 , n11749 );
    and g34429 ( n24862 , n17671 , n31559 );
    and g34430 ( n30604 , n18446 , n16916 );
    or g34431 ( n19773 , n34792 , n29393 );
    and g34432 ( n35789 , n12818 , n11 );
    and g34433 ( n6975 , n2065 , n19423 );
    or g34434 ( n24808 , n14682 , n28240 );
    xnor g34435 ( n16465 , n21921 , n6633 );
    and g34436 ( n18015 , n10493 , n17975 );
    and g34437 ( n14929 , n4221 , n18465 );
    or g34438 ( n15569 , n35899 , n21579 );
    or g34439 ( n4197 , n23604 , n6698 );
    and g34440 ( n10411 , n17328 , n32937 );
    and g34441 ( n2838 , n2733 , n29839 );
    xnor g34442 ( n30236 , n20717 , n12806 );
    or g34443 ( n9637 , n1392 , n13901 );
    or g34444 ( n33577 , n30332 , n7448 );
    or g34445 ( n17312 , n19743 , n17928 );
    and g34446 ( n4880 , n7116 , n31937 );
    and g34447 ( n3218 , n23988 , n14048 );
    buf g34448 ( n29643 , n15967 );
    not g34449 ( n16245 , n22599 );
    or g34450 ( n21901 , n15495 , n30431 );
    or g34451 ( n1646 , n15945 , n19576 );
    nor g34452 ( n13673 , n27291 , n35010 );
    xnor g34453 ( n15432 , n28479 , n8432 );
    and g34454 ( n17724 , n27072 , n33190 );
    or g34455 ( n300 , n26822 , n544 );
    or g34456 ( n24645 , n2936 , n22824 );
    not g34457 ( n24304 , n30711 );
    or g34458 ( n15546 , n27336 , n19581 );
    xnor g34459 ( n3342 , n31637 , n3134 );
    not g34460 ( n13495 , n2805 );
    or g34461 ( n3013 , n3946 , n1488 );
    and g34462 ( n29461 , n16523 , n15586 );
    xnor g34463 ( n3409 , n11992 , n5189 );
    or g34464 ( n25038 , n34646 , n11483 );
    and g34465 ( n27885 , n16453 , n14695 );
    nor g34466 ( n15667 , n18483 , n29810 );
    and g34467 ( n28260 , n21752 , n35049 );
    or g34468 ( n27081 , n22291 , n32331 );
    xnor g34469 ( n7084 , n12582 , n11827 );
    and g34470 ( n8259 , n16918 , n20333 );
    and g34471 ( n23346 , n35993 , n23861 );
    and g34472 ( n21147 , n1300 , n4025 );
    or g34473 ( n3037 , n31799 , n23045 );
    or g34474 ( n15521 , n11964 , n34381 );
    xnor g34475 ( n9997 , n4032 , n10415 );
    and g34476 ( n1866 , n31776 , n32103 );
    xnor g34477 ( n4728 , n17529 , n33113 );
    not g34478 ( n12956 , n30519 );
    and g34479 ( n29495 , n19743 , n30742 );
    or g34480 ( n12933 , n7136 , n18672 );
    and g34481 ( n20099 , n4781 , n31374 );
    or g34482 ( n32367 , n25577 , n15344 );
    and g34483 ( n1639 , n736 , n5755 );
    or g34484 ( n22125 , n34849 , n24672 );
    or g34485 ( n401 , n8044 , n23072 );
    and g34486 ( n34203 , n28373 , n33316 );
    and g34487 ( n13292 , n5153 , n29321 );
    not g34488 ( n30802 , n34225 );
    or g34489 ( n17214 , n4962 , n32816 );
    or g34490 ( n13727 , n1440 , n18255 );
    or g34491 ( n2846 , n3784 , n34472 );
    or g34492 ( n31852 , n32095 , n3956 );
    and g34493 ( n10498 , n9572 , n5718 );
    or g34494 ( n13835 , n590 , n24505 );
    xnor g34495 ( n35279 , n25167 , n11532 );
    xnor g34496 ( n8479 , n30224 , n9568 );
    or g34497 ( n27946 , n27226 , n26004 );
    or g34498 ( n31789 , n4960 , n14566 );
    and g34499 ( n12668 , n6023 , n22006 );
    and g34500 ( n13464 , n22095 , n13930 );
    or g34501 ( n29250 , n21611 , n17829 );
    nor g34502 ( n14467 , n7698 , n21739 );
    xnor g34503 ( n7171 , n6430 , n15788 );
    and g34504 ( n23490 , n14049 , n3365 );
    or g34505 ( n18373 , n34800 , n17612 );
    or g34506 ( n20280 , n27607 , n21954 );
    and g34507 ( n2539 , n3674 , n1238 );
    xnor g34508 ( n26878 , n14969 , n27785 );
    and g34509 ( n31743 , n22913 , n12555 );
    or g34510 ( n33235 , n24593 , n27740 );
    or g34511 ( n34750 , n4216 , n36039 );
    xnor g34512 ( n14494 , n25730 , n4960 );
    or g34513 ( n29404 , n1370 , n9675 );
    or g34514 ( n21287 , n1708 , n8181 );
    and g34515 ( n4017 , n35302 , n28270 );
    xnor g34516 ( n11139 , n29287 , n22455 );
    or g34517 ( n23738 , n10999 , n949 );
    not g34518 ( n1125 , n9437 );
    buf g34519 ( n22471 , n29203 );
    or g34520 ( n22596 , n9878 , n9194 );
    nor g34521 ( n19738 , n24371 , n5791 );
    or g34522 ( n31547 , n27240 , n36000 );
    and g34523 ( n34139 , n6603 , n32708 );
    or g34524 ( n22743 , n18498 , n34971 );
    nor g34525 ( n31937 , n5544 , n28685 );
    not g34526 ( n27816 , n20027 );
    xnor g34527 ( n10398 , n31077 , n7086 );
    or g34528 ( n17327 , n29357 , n24479 );
    and g34529 ( n14691 , n6079 , n32069 );
    and g34530 ( n19919 , n6408 , n35101 );
    xnor g34531 ( n18670 , n20320 , n14203 );
    xnor g34532 ( n16707 , n24098 , n31283 );
    not g34533 ( n25515 , n1694 );
    or g34534 ( n11423 , n31056 , n19028 );
    not g34535 ( n10897 , n14552 );
    or g34536 ( n9584 , n4288 , n11456 );
    or g34537 ( n4713 , n23173 , n34865 );
    and g34538 ( n9852 , n8162 , n8019 );
    or g34539 ( n10680 , n9658 , n16207 );
    or g34540 ( n23340 , n33913 , n26002 );
    or g34541 ( n3566 , n20460 , n11593 );
    xnor g34542 ( n23690 , n19954 , n7187 );
    or g34543 ( n29481 , n3205 , n14910 );
    xnor g34544 ( n27216 , n2803 , n9809 );
    or g34545 ( n22191 , n32218 , n32959 );
    xnor g34546 ( n35220 , n23006 , n15455 );
    buf g34547 ( n20300 , n12725 );
    nor g34548 ( n27642 , n19195 , n7270 );
    buf g34549 ( n21002 , n9006 );
    xnor g34550 ( n18412 , n6033 , n4878 );
    xnor g34551 ( n16612 , n9237 , n3832 );
    not g34552 ( n25021 , n13659 );
    xnor g34553 ( n29728 , n34883 , n4283 );
    or g34554 ( n30913 , n29991 , n25166 );
    and g34555 ( n22940 , n14783 , n21643 );
    or g34556 ( n19986 , n3768 , n10872 );
    or g34557 ( n15608 , n21722 , n34804 );
    or g34558 ( n26043 , n15168 , n19058 );
    or g34559 ( n26333 , n35235 , n8629 );
    and g34560 ( n11194 , n27791 , n10179 );
    xnor g34561 ( n21648 , n10372 , n13525 );
    not g34562 ( n860 , n22980 );
    or g34563 ( n11327 , n25136 , n17046 );
    not g34564 ( n3683 , n25347 );
    xnor g34565 ( n23403 , n2768 , n10354 );
    xnor g34566 ( n30974 , n25514 , n4962 );
    nor g34567 ( n29376 , n10675 , n14672 );
    xnor g34568 ( n24063 , n28385 , n22992 );
    and g34569 ( n32330 , n19797 , n13739 );
    xnor g34570 ( n24453 , n10290 , n11046 );
    nor g34571 ( n260 , n3859 , n19896 );
    and g34572 ( n10385 , n4925 , n7382 );
    and g34573 ( n10913 , n15493 , n33419 );
    or g34574 ( n6771 , n25727 , n100 );
    not g34575 ( n21382 , n27890 );
    not g34576 ( n9881 , n30553 );
    nor g34577 ( n23460 , n25602 , n29487 );
    or g34578 ( n18360 , n31750 , n11593 );
    and g34579 ( n8618 , n22271 , n18082 );
    or g34580 ( n8353 , n2317 , n10872 );
    or g34581 ( n30834 , n30393 , n17354 );
    or g34582 ( n22836 , n33782 , n171 );
    and g34583 ( n17675 , n25671 , n13846 );
    nor g34584 ( n22553 , n6025 , n24707 );
    and g34585 ( n17992 , n19445 , n22136 );
    nor g34586 ( n22886 , n6499 , n6538 );
    or g34587 ( n15789 , n4288 , n19720 );
    or g34588 ( n28967 , n25363 , n4952 );
    nor g34589 ( n23674 , n16620 , n25672 );
    or g34590 ( n7093 , n31830 , n12596 );
    nor g34591 ( n7991 , n15886 , n6730 );
    nor g34592 ( n16459 , n21317 , n6216 );
    xnor g34593 ( n2632 , n29145 , n33711 );
    and g34594 ( n19189 , n11932 , n16151 );
    or g34595 ( n35291 , n11791 , n35141 );
    not g34596 ( n28510 , n3222 );
    or g34597 ( n24845 , n35697 , n3736 );
    or g34598 ( n3318 , n3930 , n24826 );
    not g34599 ( n5079 , n7485 );
    not g34600 ( n26634 , n28273 );
    or g34601 ( n9603 , n16892 , n26480 );
    or g34602 ( n18178 , n4018 , n17068 );
    or g34603 ( n867 , n25174 , n14751 );
    and g34604 ( n13349 , n26599 , n26301 );
    nor g34605 ( n8542 , n5738 , n30575 );
    and g34606 ( n30185 , n3586 , n30509 );
    or g34607 ( n31520 , n13595 , n7293 );
    nor g34608 ( n971 , n29713 , n10164 );
    or g34609 ( n10763 , n27647 , n4175 );
    or g34610 ( n3472 , n5513 , n8601 );
    not g34611 ( n2436 , n16223 );
    and g34612 ( n12575 , n24039 , n10133 );
    or g34613 ( n5528 , n12300 , n5929 );
    xnor g34614 ( n27806 , n14363 , n32857 );
    xnor g34615 ( n26438 , n9201 , n6261 );
    xnor g34616 ( n7836 , n27513 , n2132 );
    and g34617 ( n351 , n1056 , n1743 );
    and g34618 ( n30037 , n10278 , n31348 );
    and g34619 ( n23880 , n17779 , n587 );
    or g34620 ( n28028 , n16573 , n19464 );
    or g34621 ( n31668 , n26005 , n479 );
    xnor g34622 ( n26176 , n15836 , n9613 );
    or g34623 ( n26273 , n26025 , n29178 );
    or g34624 ( n22727 , n34704 , n35852 );
    and g34625 ( n21540 , n8884 , n12009 );
    or g34626 ( n6702 , n4325 , n10960 );
    and g34627 ( n13011 , n11367 , n22265 );
    and g34628 ( n35171 , n2738 , n10220 );
    and g34629 ( n17468 , n22597 , n4878 );
    or g34630 ( n31952 , n5944 , n1402 );
    or g34631 ( n35515 , n23916 , n22206 );
    or g34632 ( n5832 , n4242 , n8153 );
    or g34633 ( n10641 , n25328 , n35561 );
    nor g34634 ( n25486 , n14537 , n17233 );
    xnor g34635 ( n49 , n19546 , n33630 );
    and g34636 ( n91 , n7082 , n11431 );
    or g34637 ( n13242 , n9779 , n4254 );
    xnor g34638 ( n35067 , n8683 , n29884 );
    or g34639 ( n21828 , n30742 , n4143 );
    nor g34640 ( n23826 , n9658 , n13615 );
    xnor g34641 ( n36075 , n3497 , n8432 );
    or g34642 ( n23498 , n12269 , n4260 );
    or g34643 ( n131 , n29764 , n3756 );
    xnor g34644 ( n15258 , n30953 , n32715 );
    or g34645 ( n23417 , n31799 , n13630 );
    xnor g34646 ( n25336 , n35925 , n20795 );
    or g34647 ( n5856 , n31862 , n6756 );
    xnor g34648 ( n21509 , n11078 , n1555 );
    or g34649 ( n27484 , n35824 , n7668 );
    or g34650 ( n6353 , n10290 , n17962 );
    or g34651 ( n12887 , n28927 , n10140 );
    nor g34652 ( n34777 , n31475 , n22111 );
    nor g34653 ( n32461 , n23604 , n14765 );
    xnor g34654 ( n13587 , n22891 , n31559 );
    xnor g34655 ( n11337 , n430 , n5271 );
    and g34656 ( n3191 , n10844 , n30168 );
    or g34657 ( n35086 , n4008 , n139 );
    or g34658 ( n11562 , n33023 , n20640 );
    xnor g34659 ( n30320 , n7662 , n4606 );
    or g34660 ( n24594 , n6852 , n8924 );
    xor g34661 ( n6047 , n20348 , n11151 );
    or g34662 ( n19141 , n3399 , n35979 );
    and g34663 ( n28734 , n18210 , n2788 );
    nor g34664 ( n34784 , n11455 , n1319 );
    xnor g34665 ( n15838 , n21394 , n32589 );
    or g34666 ( n18576 , n24371 , n4962 );
    or g34667 ( n8296 , n968 , n31067 );
    and g34668 ( n27849 , n20781 , n25480 );
    not g34669 ( n23791 , n8638 );
    xnor g34670 ( n18472 , n34824 , n256 );
    nor g34671 ( n29525 , n17250 , n6548 );
    and g34672 ( n13768 , n9643 , n4340 );
    and g34673 ( n12460 , n2129 , n14040 );
    or g34674 ( n23631 , n26910 , n21956 );
    or g34675 ( n15850 , n24276 , n33088 );
    and g34676 ( n34516 , n562 , n28352 );
    or g34677 ( n28400 , n18379 , n31953 );
    and g34678 ( n30838 , n26829 , n30550 );
    not g34679 ( n8958 , n22980 );
    or g34680 ( n4572 , n1950 , n22495 );
    or g34681 ( n7620 , n15267 , n16457 );
    or g34682 ( n25391 , n410 , n13900 );
    and g34683 ( n8121 , n4394 , n19788 );
    xnor g34684 ( n3045 , n12466 , n15886 );
    xnor g34685 ( n19907 , n24664 , n17152 );
    or g34686 ( n35674 , n18502 , n35394 );
    or g34687 ( n4505 , n35279 , n19403 );
    nor g34688 ( n7815 , n35415 , n16112 );
    not g34689 ( n15871 , n4772 );
    or g34690 ( n9211 , n7138 , n2119 );
    xnor g34691 ( n35988 , n25144 , n18033 );
    and g34692 ( n20050 , n6019 , n27464 );
    xnor g34693 ( n6225 , n25228 , n10894 );
    and g34694 ( n7578 , n7370 , n31176 );
    or g34695 ( n17720 , n2221 , n23625 );
    xnor g34696 ( n6832 , n969 , n1491 );
    xnor g34697 ( n23449 , n2345 , n27181 );
    or g34698 ( n10959 , n28791 , n19403 );
    xnor g34699 ( n34848 , n13018 , n23365 );
    not g34700 ( n6380 , n22279 );
    and g34701 ( n4901 , n23405 , n9741 );
    xnor g34702 ( n24462 , n13280 , n2127 );
    or g34703 ( n5902 , n2201 , n2813 );
    or g34704 ( n607 , n7347 , n22858 );
    or g34705 ( n14420 , n7094 , n25970 );
    and g34706 ( n32614 , n539 , n10886 );
    and g34707 ( n21105 , n463 , n518 );
    or g34708 ( n26610 , n16135 , n3990 );
    not g34709 ( n26346 , n16223 );
    xnor g34710 ( n15724 , n1356 , n22129 );
    xnor g34711 ( n23275 , n24346 , n29839 );
    not g34712 ( n19287 , n33795 );
    nor g34713 ( n4556 , n402 , n32731 );
    or g34714 ( n861 , n32715 , n14849 );
    or g34715 ( n31980 , n1950 , n21654 );
    xnor g34716 ( n4652 , n32157 , n961 );
    or g34717 ( n28884 , n20216 , n34537 );
    or g34718 ( n25472 , n2125 , n29077 );
    or g34719 ( n19033 , n27915 , n13948 );
    not g34720 ( n16497 , n20558 );
    not g34721 ( n5699 , n22471 );
    xnor g34722 ( n3793 , n3387 , n8844 );
    and g34723 ( n12419 , n19696 , n32880 );
    or g34724 ( n29337 , n23543 , n14473 );
    nor g34725 ( n24939 , n34834 , n6738 );
    or g34726 ( n7707 , n16620 , n11634 );
    xnor g34727 ( n16950 , n33182 , n34942 );
    or g34728 ( n8099 , n10884 , n545 );
    or g34729 ( n2036 , n32095 , n18334 );
    buf g34730 ( n30947 , n2712 );
    xnor g34731 ( n34747 , n30739 , n21735 );
    not g34732 ( n1463 , n21 );
    and g34733 ( n8716 , n32650 , n30931 );
    or g34734 ( n4251 , n4773 , n9951 );
    or g34735 ( n15462 , n28082 , n32484 );
    xnor g34736 ( n28892 , n4540 , n10894 );
    or g34737 ( n10024 , n29884 , n24791 );
    or g34738 ( n29619 , n8060 , n25761 );
    or g34739 ( n8822 , n33773 , n34862 );
    or g34740 ( n10712 , n22801 , n6077 );
    and g34741 ( n35808 , n20990 , n36061 );
    or g34742 ( n6242 , n30147 , n27990 );
    and g34743 ( n34883 , n3601 , n15224 );
    or g34744 ( n13052 , n29696 , n7964 );
    or g34745 ( n29875 , n32095 , n11468 );
    or g34746 ( n25087 , n8148 , n24120 );
    or g34747 ( n10165 , n17568 , n6645 );
    nor g34748 ( n17102 , n29824 , n11600 );
    xnor g34749 ( n8898 , n32232 , n10341 );
    and g34750 ( n21778 , n31327 , n10242 );
    nor g34751 ( n20314 , n11313 , n8423 );
    or g34752 ( n6345 , n16858 , n16594 );
    or g34753 ( n11783 , n16038 , n9832 );
    xnor g34754 ( n6373 , n34541 , n3222 );
    and g34755 ( n23933 , n31431 , n3778 );
    xnor g34756 ( n13696 , n24631 , n673 );
    xnor g34757 ( n25163 , n14038 , n20512 );
    or g34758 ( n7958 , n25520 , n34315 );
    not g34759 ( n21418 , n544 );
    and g34760 ( n32689 , n10854 , n15943 );
    and g34761 ( n20176 , n5797 , n5136 );
    and g34762 ( n18934 , n15344 , n5549 );
    or g34763 ( n3392 , n16209 , n23209 );
    xnor g34764 ( n177 , n11956 , n7254 );
    xnor g34765 ( n9890 , n17215 , n2292 );
    not g34766 ( n25521 , n648 );
    xnor g34767 ( n5944 , n2752 , n6897 );
    nor g34768 ( n23829 , n12701 , n10428 );
    or g34769 ( n7550 , n2770 , n2955 );
    and g34770 ( n5877 , n6413 , n2940 );
    or g34771 ( n23413 , n9544 , n4081 );
    or g34772 ( n10355 , n31997 , n10591 );
    xnor g34773 ( n25196 , n6624 , n19984 );
    or g34774 ( n8091 , n32715 , n5864 );
    xnor g34775 ( n5630 , n19205 , n33758 );
    or g34776 ( n27571 , n34885 , n30541 );
    xnor g34777 ( n877 , n14995 , n16292 );
    or g34778 ( n13542 , n28899 , n5209 );
    or g34779 ( n32635 , n22291 , n10818 );
    nor g34780 ( n3758 , n7540 , n22700 );
    nor g34781 ( n18524 , n3205 , n22590 );
    or g34782 ( n33628 , n21823 , n16554 );
    or g34783 ( n16726 , n10894 , n8658 );
    not g34784 ( n30310 , n4712 );
    or g34785 ( n23294 , n33701 , n16961 );
    not g34786 ( n26466 , n6307 );
    not g34787 ( n29959 , n23604 );
    not g34788 ( n13719 , n31421 );
    xnor g34789 ( n23432 , n25912 , n4962 );
    and g34790 ( n14827 , n1703 , n6186 );
    or g34791 ( n7489 , n31559 , n25575 );
    nor g34792 ( n34213 , n19551 , n18745 );
    xnor g34793 ( n27098 , n11470 , n5335 );
    and g34794 ( n33742 , n1599 , n3137 );
    xnor g34795 ( n9842 , n18801 , n10894 );
    xnor g34796 ( n7667 , n22119 , n11179 );
    nor g34797 ( n634 , n4803 , n30904 );
    not g34798 ( n18770 , n34098 );
    and g34799 ( n35258 , n26872 , n16433 );
    xnor g34800 ( n21153 , n14176 , n24169 );
    or g34801 ( n32867 , n20846 , n28675 );
    or g34802 ( n24535 , n24447 , n30825 );
    and g34803 ( n30813 , n24574 , n34582 );
    or g34804 ( n20915 , n1878 , n24944 );
    not g34805 ( n8515 , n16107 );
    not g34806 ( n29489 , n8977 );
    or g34807 ( n33703 , n22139 , n23323 );
    not g34808 ( n6216 , n22200 );
    xnor g34809 ( n33913 , n6422 , n34746 );
    or g34810 ( n30592 , n16733 , n30646 );
    or g34811 ( n21111 , n18525 , n17354 );
    xnor g34812 ( n35681 , n19819 , n30742 );
    not g34813 ( n12302 , n9789 );
    or g34814 ( n8588 , n22786 , n33956 );
    and g34815 ( n18045 , n32788 , n27976 );
    nor g34816 ( n23170 , n9246 , n13193 );
    or g34817 ( n35058 , n35927 , n29529 );
    xor g34818 ( n35520 , n2875 , n25231 );
    or g34819 ( n13631 , n10236 , n6950 );
    or g34820 ( n2407 , n16804 , n23028 );
    and g34821 ( n21015 , n30145 , n30640 );
    and g34822 ( n16102 , n18653 , n28296 );
    and g34823 ( n32281 , n22816 , n1213 );
    or g34824 ( n35025 , n6469 , n24489 );
    or g34825 ( n17030 , n12185 , n23211 );
    xnor g34826 ( n21030 , n35883 , n1950 );
    xnor g34827 ( n13491 , n8198 , n6975 );
    not g34828 ( n6908 , n29555 );
    not g34829 ( n26937 , n1950 );
    not g34830 ( n24410 , n19984 );
    and g34831 ( n32991 , n30939 , n1294 );
    and g34832 ( n4055 , n6010 , n5264 );
    or g34833 ( n17035 , n3045 , n31848 );
    or g34834 ( n1704 , n8658 , n34472 );
    or g34835 ( n25579 , n35311 , n3936 );
    xnor g34836 ( n23634 , n9501 , n25174 );
    xnor g34837 ( n14970 , n30304 , n5826 );
    and g34838 ( n27434 , n21686 , n11547 );
    nor g34839 ( n13377 , n4461 , n26466 );
    or g34840 ( n434 , n4288 , n16573 );
    xnor g34841 ( n430 , n18183 , n27121 );
    or g34842 ( n15377 , n31961 , n17651 );
    or g34843 ( n24526 , n10509 , n21210 );
    and g34844 ( n23864 , n21943 , n27365 );
    and g34845 ( n32580 , n6146 , n21992 );
    not g34846 ( n10316 , n2666 );
    xnor g34847 ( n25271 , n29665 , n11878 );
    or g34848 ( n15014 , n9789 , n7350 );
    or g34849 ( n9258 , n9919 , n31740 );
    not g34850 ( n16247 , n35877 );
    or g34851 ( n2478 , n11046 , n34119 );
    buf g34852 ( n35422 , n21100 );
    or g34853 ( n1647 , n13107 , n6554 );
    or g34854 ( n33589 , n16048 , n22206 );
    or g34855 ( n5796 , n22202 , n1642 );
    xnor g34856 ( n35 , n22117 , n13306 );
    xnor g34857 ( n77 , n610 , n23604 );
    and g34858 ( n4917 , n5323 , n20724 );
    and g34859 ( n31643 , n8768 , n9541 );
    xnor g34860 ( n12556 , n7921 , n8432 );
    and g34861 ( n35228 , n20473 , n4473 );
    or g34862 ( n21790 , n11046 , n10290 );
    xnor g34863 ( n11889 , n25128 , n18170 );
    or g34864 ( n32724 , n23185 , n14918 );
    or g34865 ( n20935 , n28587 , n18488 );
    or g34866 ( n17584 , n34918 , n35748 );
    or g34867 ( n10179 , n5287 , n13299 );
    or g34868 ( n11486 , n6605 , n34970 );
    and g34869 ( n13743 , n17987 , n3446 );
    and g34870 ( n29081 , n12063 , n31640 );
    or g34871 ( n18570 , n11320 , n34968 );
    not g34872 ( n18803 , n10336 );
    and g34873 ( n11468 , n5815 , n777 );
    and g34874 ( n21490 , n5486 , n27520 );
    and g34875 ( n32437 , n24309 , n22094 );
    and g34876 ( n23052 , n30596 , n29798 );
    and g34877 ( n30159 , n34420 , n22796 );
    or g34878 ( n25479 , n9673 , n9731 );
    nor g34879 ( n5691 , n3205 , n14037 );
    and g34880 ( n241 , n14644 , n17561 );
    or g34881 ( n9452 , n23604 , n24537 );
    xnor g34882 ( n16050 , n7502 , n22898 );
    buf g34883 ( n6340 , n7214 );
    or g34884 ( n5371 , n22815 , n22377 );
    not g34885 ( n18711 , n9658 );
    and g34886 ( n8914 , n29247 , n35376 );
    xnor g34887 ( n10512 , n16841 , n4288 );
    nor g34888 ( n22708 , n4960 , n13121 );
    or g34889 ( n24123 , n3197 , n15766 );
    nor g34890 ( n16163 , n1950 , n13292 );
    and g34891 ( n4301 , n26679 , n31171 );
    and g34892 ( n35659 , n21028 , n15971 );
    or g34893 ( n2350 , n17944 , n6532 );
    or g34894 ( n33934 , n31215 , n10829 );
    and g34895 ( n23565 , n18 , n804 );
    and g34896 ( n296 , n33617 , n7640 );
    or g34897 ( n5003 , n22865 , n3619 );
    and g34898 ( n10479 , n18239 , n16106 );
    or g34899 ( n14974 , n34134 , n19521 );
    xnor g34900 ( n12083 , n2610 , n31289 );
    nor g34901 ( n21681 , n72 , n35468 );
    xnor g34902 ( n16702 , n35004 , n29713 );
    not g34903 ( n35643 , n7588 );
    xnor g34904 ( n3557 , n9808 , n27201 );
    or g34905 ( n5035 , n8432 , n20977 );
    and g34906 ( n34039 , n19882 , n5217 );
    not g34907 ( n4496 , n28273 );
    and g34908 ( n10457 , n28256 , n8515 );
    and g34909 ( n13045 , n2773 , n8246 );
    or g34910 ( n16066 , n11346 , n4653 );
    or g34911 ( n31251 , n15349 , n29493 );
    or g34912 ( n33684 , n35022 , n30206 );
    or g34913 ( n34343 , n34004 , n21210 );
    not g34914 ( n542 , n18296 );
    or g34915 ( n22656 , n10353 , n12428 );
    xnor g34916 ( n22254 , n34847 , n19955 );
    and g34917 ( n14579 , n24010 , n30652 );
    or g34918 ( n28829 , n1752 , n2119 );
    xnor g34919 ( n24648 , n386 , n2736 );
    nor g34920 ( n28376 , n7139 , n31411 );
    xnor g34921 ( n11141 , n3626 , n23604 );
    not g34922 ( n1327 , n17998 );
    and g34923 ( n655 , n17956 , n24215 );
    and g34924 ( n30967 , n1735 , n26658 );
    and g34925 ( n30282 , n11517 , n1486 );
    or g34926 ( n2388 , n19926 , n30983 );
    and g34927 ( n34676 , n16386 , n27068 );
    and g34928 ( n28839 , n19899 , n17283 );
    and g34929 ( n6106 , n11012 , n4194 );
    and g34930 ( n11798 , n26000 , n7311 );
    and g34931 ( n6091 , n18582 , n34149 );
    and g34932 ( n5996 , n19369 , n3705 );
    or g34933 ( n19505 , n4288 , n28306 );
    and g34934 ( n29911 , n16932 , n4549 );
    not g34935 ( n15795 , n30713 );
    and g34936 ( n30132 , n22648 , n12799 );
    or g34937 ( n26715 , n26967 , n30156 );
    or g34938 ( n9694 , n8713 , n814 );
    or g34939 ( n25279 , n687 , n29393 );
    xnor g34940 ( n15876 , n29452 , n2495 );
    xnor g34941 ( n31084 , n30173 , n4960 );
    not g34942 ( n26578 , n12428 );
    or g34943 ( n19567 , n4758 , n25612 );
    xnor g34944 ( n27049 , n33101 , n32584 );
    xnor g34945 ( n27646 , n9791 , n3583 );
    and g34946 ( n19544 , n30623 , n26372 );
    and g34947 ( n20582 , n32628 , n18733 );
    or g34948 ( n31121 , n16620 , n22153 );
    or g34949 ( n30138 , n6848 , n528 );
    or g34950 ( n5463 , n32095 , n18862 );
    not g34951 ( n35113 , n4288 );
    nor g34952 ( n23043 , n35704 , n19169 );
    and g34953 ( n25841 , n32310 , n15208 );
    or g34954 ( n25660 , n20262 , n33654 );
    not g34955 ( n35541 , n16620 );
    xnor g34956 ( n22922 , n6645 , n17568 );
    not g34957 ( n28157 , n15464 );
    xnor g34958 ( n31591 , n9267 , n16922 );
    or g34959 ( n33419 , n11455 , n19821 );
    not g34960 ( n29510 , n35927 );
    or g34961 ( n7986 , n33370 , n31140 );
    or g34962 ( n17519 , n36077 , n30183 );
    or g34963 ( n35848 , n23475 , n4649 );
    or g34964 ( n35991 , n20894 , n35757 );
    nor g34965 ( n29914 , n8165 , n22535 );
    xnor g34966 ( n22771 , n21200 , n29884 );
    not g34967 ( n9590 , n3071 );
    xnor g34968 ( n695 , n5178 , n31289 );
    xnor g34969 ( n31183 , n30144 , n32715 );
    or g34970 ( n6271 , n31799 , n23843 );
    and g34971 ( n30660 , n3410 , n30857 );
    xnor g34972 ( n11396 , n31948 , n29839 );
    not g34973 ( n6293 , n14394 );
    xnor g34974 ( n5945 , n24258 , n6339 );
    and g34975 ( n12127 , n9907 , n25493 );
    or g34976 ( n11561 , n2333 , n8983 );
    xnor g34977 ( n2784 , n17171 , n11737 );
    xnor g34978 ( n21255 , n16209 , n11046 );
    or g34979 ( n65 , n32965 , n20257 );
    and g34980 ( n28187 , n22490 , n5769 );
    xnor g34981 ( n27459 , n26194 , n33444 );
    xnor g34982 ( n17012 , n26910 , n31753 );
    or g34983 ( n15243 , n24332 , n29693 );
    or g34984 ( n17540 , n8784 , n32425 );
    and g34985 ( n4896 , n4686 , n1742 );
    buf g34986 ( n15109 , n4852 );
    or g34987 ( n6644 , n32758 , n3267 );
    or g34988 ( n25451 , n24162 , n32718 );
    nor g34989 ( n16676 , n18787 , n21294 );
    and g34990 ( n3610 , n14132 , n17768 );
    and g34991 ( n7254 , n6342 , n826 );
    xnor g34992 ( n27339 , n33046 , n5850 );
    xnor g34993 ( n30645 , n23570 , n33221 );
    not g34994 ( n16996 , n15299 );
    xnor g34995 ( n27565 , n27188 , n9568 );
    or g34996 ( n34222 , n13859 , n29602 );
    not g34997 ( n27626 , n5362 );
    not g34998 ( n26467 , n20650 );
    or g34999 ( n27303 , n33347 , n17111 );
    or g35000 ( n29717 , n1012 , n31067 );
    not g35001 ( n19218 , n16223 );
    or g35002 ( n23739 , n1268 , n16519 );
    xnor g35003 ( n35533 , n18648 , n24561 );
    not g35004 ( n8070 , n36074 );
    or g35005 ( n3740 , n31861 , n20318 );
    xnor g35006 ( n35486 , n23857 , n20375 );
    xnor g35007 ( n31629 , n26859 , n7976 );
    or g35008 ( n24099 , n12931 , n15602 );
    or g35009 ( n31139 , n6707 , n29872 );
    nor g35010 ( n24824 , n16922 , n9878 );
    xnor g35011 ( n34554 , n2758 , n31032 );
    or g35012 ( n12720 , n26304 , n2903 );
    or g35013 ( n17686 , n18905 , n26002 );
    or g35014 ( n33238 , n17134 , n12596 );
    or g35015 ( n5927 , n25174 , n24286 );
    not g35016 ( n5795 , n25602 );
    not g35017 ( n10568 , n12550 );
    not g35018 ( n1438 , n32857 );
    or g35019 ( n1637 , n10698 , n32572 );
    not g35020 ( n18484 , n18194 );
    xnor g35021 ( n520 , n17445 , n30354 );
    xnor g35022 ( n35888 , n10674 , n11185 );
    not g35023 ( n15745 , n15886 );
    xnor g35024 ( n4401 , n34830 , n6233 );
    xnor g35025 ( n27767 , n880 , n13246 );
    or g35026 ( n35336 , n16342 , n6721 );
    or g35027 ( n25396 , n19150 , n15439 );
    xnor g35028 ( n16319 , n15191 , n5335 );
    or g35029 ( n26114 , n16377 , n35143 );
    or g35030 ( n30031 , n8927 , n32959 );
    and g35031 ( n12498 , n26061 , n5832 );
    or g35032 ( n16613 , n13392 , n20762 );
    nor g35033 ( n11038 , n31559 , n2387 );
    or g35034 ( n14403 , n13830 , n5900 );
    not g35035 ( n15877 , n9789 );
    nor g35036 ( n17985 , n16135 , n22932 );
    and g35037 ( n5005 , n7190 , n33659 );
    nor g35038 ( n22440 , n5345 , n28778 );
    xnor g35039 ( n33222 , n30588 , n13760 );
    or g35040 ( n15891 , n31272 , n34283 );
    and g35041 ( n7877 , n26248 , n25845 );
    and g35042 ( n28139 , n29473 , n9871 );
    nor g35043 ( n8500 , n5067 , n34967 );
    or g35044 ( n582 , n23183 , n34557 );
    or g35045 ( n11026 , n30742 , n313 );
    xnor g35046 ( n19858 , n36078 , n4878 );
    and g35047 ( n10313 , n5291 , n3403 );
    and g35048 ( n17986 , n9865 , n24089 );
    and g35049 ( n28247 , n19964 , n10189 );
    and g35050 ( n14652 , n16859 , n199 );
    or g35051 ( n14675 , n28767 , n15490 );
    and g35052 ( n30190 , n13741 , n35023 );
    and g35053 ( n15369 , n24242 , n34193 );
    not g35054 ( n10428 , n29560 );
    or g35055 ( n10337 , n3463 , n2524 );
    or g35056 ( n32699 , n1842 , n28123 );
    and g35057 ( n441 , n28773 , n11290 );
    or g35058 ( n8112 , n1865 , n14886 );
    xnor g35059 ( n25642 , n32021 , n30079 );
    and g35060 ( n13646 , n16221 , n35910 );
    or g35061 ( n18571 , n20016 , n15496 );
    or g35062 ( n35063 , n16620 , n19209 );
    or g35063 ( n31842 , n21280 , n2823 );
    or g35064 ( n33546 , n23604 , n3626 );
    nor g35065 ( n21985 , n22982 , n24864 );
    nor g35066 ( n24200 , n16636 , n18151 );
    xnor g35067 ( n34535 , n19948 , n27584 );
    nor g35068 ( n16602 , n12064 , n28666 );
    and g35069 ( n10801 , n25210 , n16434 );
    xnor g35070 ( n1962 , n1127 , n15834 );
    or g35071 ( n32373 , n6880 , n21673 );
    and g35072 ( n7443 , n2265 , n34520 );
    buf g35073 ( n28455 , n266 );
    and g35074 ( n9309 , n3447 , n23408 );
    not g35075 ( n10895 , n30372 );
    buf g35076 ( n13015 , n29928 );
    and g35077 ( n10591 , n22315 , n35034 );
    and g35078 ( n1407 , n12523 , n22126 );
    nor g35079 ( n16688 , n21664 , n30335 );
    and g35080 ( n18398 , n28085 , n33030 );
    xnor g35081 ( n10629 , n365 , n31272 );
    xnor g35082 ( n20586 , n15727 , n4962 );
    nor g35083 ( n22664 , n31215 , n4492 );
    or g35084 ( n14729 , n24117 , n7982 );
    or g35085 ( n3478 , n12155 , n7647 );
    or g35086 ( n6006 , n13580 , n2661 );
    not g35087 ( n11571 , n2006 );
    xnor g35088 ( n29158 , n199 , n16859 );
    xnor g35089 ( n10567 , n28735 , n5094 );
    nor g35090 ( n34292 , n830 , n852 );
    or g35091 ( n22212 , n17751 , n17505 );
    or g35092 ( n29175 , n35927 , n31535 );
    xnor g35093 ( n35322 , n13545 , n25171 );
    not g35094 ( n33295 , n21030 );
    xnor g35095 ( n19142 , n1297 , n35927 );
    or g35096 ( n5756 , n19438 , n27854 );
    or g35097 ( n24576 , n23373 , n4478 );
    xnor g35098 ( n1268 , n32856 , n30742 );
    or g35099 ( n34257 , n14373 , n10420 );
    or g35100 ( n1816 , n32095 , n18426 );
    or g35101 ( n16866 , n20565 , n28559 );
    and g35102 ( n34315 , n29869 , n4705 );
    and g35103 ( n30716 , n21581 , n15302 );
    or g35104 ( n26945 , n35292 , n5252 );
    or g35105 ( n28597 , n18375 , n5008 );
    or g35106 ( n11402 , n31559 , n17755 );
    and g35107 ( n16395 , n3028 , n32095 );
    and g35108 ( n30337 , n22148 , n21805 );
    or g35109 ( n22565 , n4288 , n23322 );
    or g35110 ( n33946 , n3946 , n25065 );
    xnor g35111 ( n18683 , n19009 , n3025 );
    or g35112 ( n31476 , n1422 , n1856 );
    or g35113 ( n1814 , n1408 , n11850 );
    or g35114 ( n1607 , n3812 , n3738 );
    xnor g35115 ( n15156 , n13177 , n9658 );
    and g35116 ( n20371 , n10695 , n12904 );
    or g35117 ( n29664 , n8498 , n34912 );
    nor g35118 ( n7629 , n24371 , n35282 );
    nor g35119 ( n4860 , n20631 , n5602 );
    and g35120 ( n32091 , n31805 , n22435 );
    or g35121 ( n8709 , n23604 , n25267 );
    xnor g35122 ( n36065 , n31400 , n16079 );
    or g35123 ( n8718 , n34650 , n14699 );
    or g35124 ( n18337 , n7902 , n743 );
    or g35125 ( n23802 , n31317 , n33647 );
    or g35126 ( n20121 , n24596 , n7657 );
    or g35127 ( n17882 , n18245 , n32679 );
    or g35128 ( n25335 , n17568 , n8804 );
    xnor g35129 ( n19047 , n16422 , n9826 );
    or g35130 ( n18351 , n28509 , n15501 );
    xnor g35131 ( n9042 , n17349 , n2890 );
    or g35132 ( n14054 , n11455 , n13805 );
    or g35133 ( n15598 , n14239 , n1715 );
    or g35134 ( n31732 , n18612 , n10634 );
    or g35135 ( n29169 , n8798 , n16326 );
    xnor g35136 ( n12258 , n11391 , n7371 );
    and g35137 ( n10761 , n23056 , n15484 );
    or g35138 ( n9868 , n7887 , n28360 );
    and g35139 ( n13898 , n1481 , n27106 );
    or g35140 ( n31063 , n9793 , n19718 );
    and g35141 ( n27739 , n11291 , n33451 );
    or g35142 ( n16183 , n33104 , n23828 );
    or g35143 ( n6886 , n4091 , n18274 );
    or g35144 ( n24158 , n15601 , n13106 );
    or g35145 ( n21403 , n27950 , n18477 );
    and g35146 ( n20453 , n24154 , n11828 );
    buf g35147 ( n13480 , n32194 );
    not g35148 ( n14861 , n15997 );
    buf g35149 ( n1642 , n30877 );
    xnor g35150 ( n4355 , n2470 , n30742 );
    and g35151 ( n31112 , n15307 , n8006 );
    or g35152 ( n28722 , n20685 , n30089 );
    xnor g35153 ( n31027 , n34162 , n32857 );
    and g35154 ( n7166 , n1227 , n21913 );
    and g35155 ( n11704 , n27711 , n19535 );
    not g35156 ( n28236 , n11455 );
    xnor g35157 ( n686 , n29083 , n16922 );
    not g35158 ( n30317 , n23651 );
    or g35159 ( n526 , n999 , n10721 );
    xnor g35160 ( n34608 , n28889 , n15706 );
    or g35161 ( n157 , n35886 , n31055 );
    xnor g35162 ( n17180 , n7611 , n28540 );
    and g35163 ( n9811 , n33307 , n36047 );
    xnor g35164 ( n26967 , n34667 , n24371 );
    nor g35165 ( n10610 , n1010 , n23790 );
    xnor g35166 ( n14200 , n9690 , n31289 );
    nor g35167 ( n19947 , n35974 , n1603 );
    or g35168 ( n35771 , n15409 , n5358 );
    xnor g35169 ( n24599 , n29122 , n2996 );
    or g35170 ( n31614 , n31203 , n14706 );
    or g35171 ( n27913 , n3205 , n1619 );
    not g35172 ( n20925 , n20548 );
    or g35173 ( n31542 , n16740 , n10181 );
    or g35174 ( n22331 , n3946 , n8056 );
    and g35175 ( n4443 , n15438 , n29659 );
    not g35176 ( n30950 , n19562 );
    xnor g35177 ( n19294 , n29617 , n23066 );
    not g35178 ( n17355 , n6992 );
    or g35179 ( n20114 , n16135 , n17379 );
    or g35180 ( n85 , n4288 , n35506 );
    nor g35181 ( n21859 , n35140 , n27732 );
    and g35182 ( n17189 , n26024 , n23215 );
    or g35183 ( n12215 , n21324 , n17705 );
    not g35184 ( n20139 , n15769 );
    not g35185 ( n24191 , n10366 );
    not g35186 ( n29336 , n35740 );
    or g35187 ( n18895 , n15017 , n9513 );
    and g35188 ( n13708 , n1995 , n28194 );
    or g35189 ( n355 , n31060 , n3864 );
    not g35190 ( n7865 , n14977 );
    nor g35191 ( n4100 , n7697 , n25877 );
    or g35192 ( n16830 , n1944 , n12823 );
    xnor g35193 ( n14555 , n30974 , n22002 );
    xnor g35194 ( n27585 , n6976 , n11455 );
    xnor g35195 ( n16028 , n9199 , n24481 );
    not g35196 ( n11867 , n34783 );
    not g35197 ( n27080 , n16620 );
    xnor g35198 ( n12 , n25105 , n30776 );
    not g35199 ( n29907 , n35570 );
    and g35200 ( n6596 , n3829 , n22980 );
    not g35201 ( n4437 , n15107 );
    xnor g35202 ( n15187 , n12075 , n18579 );
    xnor g35203 ( n4472 , n25711 , n14101 );
    or g35204 ( n35536 , n23902 , n7711 );
    or g35205 ( n17780 , n22676 , n35143 );
    or g35206 ( n19386 , n4066 , n32026 );
    or g35207 ( n22986 , n9789 , n17128 );
    nor g35208 ( n22950 , n33201 , n26023 );
    xnor g35209 ( n10318 , n8489 , n19551 );
    xnor g35210 ( n18831 , n22771 , n7758 );
    or g35211 ( n20397 , n28593 , n8253 );
    or g35212 ( n28316 , n13713 , n29425 );
    or g35213 ( n26789 , n6148 , n12036 );
    not g35214 ( n30451 , n5335 );
    and g35215 ( n5277 , n11679 , n18131 );
    xnor g35216 ( n22405 , n21635 , n3763 );
    or g35217 ( n32254 , n31362 , n22858 );
    or g35218 ( n8790 , n21397 , n30221 );
    xnor g35219 ( n25828 , n29478 , n7540 );
    xnor g35220 ( n30948 , n33213 , n32715 );
    or g35221 ( n30628 , n18238 , n9930 );
    or g35222 ( n2598 , n7018 , n20897 );
    and g35223 ( n10213 , n9765 , n31270 );
    and g35224 ( n4157 , n18571 , n31207 );
    not g35225 ( n29124 , n22980 );
    nor g35226 ( n21432 , n5287 , n8784 );
    xnor g35227 ( n8455 , n7496 , n7118 );
    not g35228 ( n376 , n33977 );
    nor g35229 ( n12101 , n21991 , n16649 );
    xnor g35230 ( n12231 , n10753 , n13687 );
    or g35231 ( n23989 , n10894 , n2506 );
    or g35232 ( n22087 , n20904 , n20022 );
    or g35233 ( n4985 , n9793 , n18726 );
    or g35234 ( n29257 , n3603 , n22026 );
    not g35235 ( n10883 , n22291 );
    and g35236 ( n17406 , n6267 , n10722 );
    or g35237 ( n18809 , n33976 , n21644 );
    xnor g35238 ( n1827 , n14059 , n25174 );
    and g35239 ( n33557 , n22253 , n35116 );
    or g35240 ( n9044 , n18635 , n32912 );
    and g35241 ( n28182 , n22372 , n35524 );
    xnor g35242 ( n5753 , n21075 , n35453 );
    or g35243 ( n29616 , n15658 , n4260 );
    or g35244 ( n13966 , n9023 , n28623 );
    and g35245 ( n11671 , n11526 , n18717 );
    or g35246 ( n25142 , n1259 , n34347 );
    and g35247 ( n4284 , n33179 , n25288 );
    xnor g35248 ( n10702 , n32561 , n12873 );
    not g35249 ( n27687 , n17646 );
    or g35250 ( n28992 , n1204 , n2814 );
    nor g35251 ( n12349 , n4288 , n5623 );
    xnor g35252 ( n23443 , n18946 , n8866 );
    and g35253 ( n14684 , n13039 , n1150 );
    or g35254 ( n27686 , n16237 , n24479 );
    xnor g35255 ( n940 , n13617 , n9345 );
    and g35256 ( n7888 , n31404 , n662 );
    and g35257 ( n20739 , n8240 , n14294 );
    or g35258 ( n8695 , n25153 , n32126 );
    or g35259 ( n7047 , n30742 , n24822 );
    and g35260 ( n8619 , n26882 , n14622 );
    xnor g35261 ( n17672 , n31523 , n10894 );
    or g35262 ( n15098 , n11190 , n31832 );
    nor g35263 ( n15963 , n25174 , n24341 );
    and g35264 ( n29103 , n27460 , n13585 );
    or g35265 ( n34775 , n4233 , n22206 );
    and g35266 ( n23068 , n34858 , n2873 );
    or g35267 ( n25034 , n32814 , n7528 );
    xnor g35268 ( n3877 , n15291 , n31289 );
    or g35269 ( n31521 , n21502 , n2117 );
    xnor g35270 ( n20366 , n2622 , n4878 );
    or g35271 ( n5443 , n30722 , n6288 );
    and g35272 ( n15826 , n33684 , n13484 );
    and g35273 ( n5348 , n5345 , n4983 );
    or g35274 ( n1930 , n27796 , n35143 );
    and g35275 ( n6251 , n16376 , n9993 );
    or g35276 ( n34079 , n17901 , n31773 );
    or g35277 ( n3719 , n26084 , n28668 );
    nor g35278 ( n14940 , n17485 , n11712 );
    or g35279 ( n16306 , n12440 , n9951 );
    xnor g35280 ( n2648 , n15230 , n35113 );
    or g35281 ( n34239 , n5067 , n1083 );
    or g35282 ( n27480 , n7220 , n26112 );
    not g35283 ( n19895 , n274 );
    and g35284 ( n545 , n33091 , n5545 );
    and g35285 ( n34541 , n30928 , n6727 );
    or g35286 ( n1071 , n14761 , n29953 );
    and g35287 ( n2131 , n18895 , n20162 );
    or g35288 ( n25723 , n17751 , n21496 );
    and g35289 ( n34742 , n10002 , n19428 );
    or g35290 ( n4888 , n19984 , n5794 );
    or g35291 ( n11552 , n130 , n13480 );
    xnor g35292 ( n25289 , n5018 , n27285 );
    or g35293 ( n13892 , n26350 , n9030 );
    xnor g35294 ( n12768 , n12749 , n27291 );
    or g35295 ( n8395 , n32857 , n30799 );
    xnor g35296 ( n23853 , n6262 , n21308 );
    nor g35297 ( n26127 , n15886 , n20596 );
    xnor g35298 ( n30648 , n10714 , n31289 );
    and g35299 ( n10730 , n20263 , n24641 );
    or g35300 ( n29746 , n28318 , n14699 );
    and g35301 ( n19657 , n13444 , n1716 );
    or g35302 ( n8842 , n23946 , n6498 );
    or g35303 ( n12310 , n17751 , n5627 );
    nor g35304 ( n3733 , n33663 , n19957 );
    or g35305 ( n3313 , n13348 , n12996 );
    not g35306 ( n31285 , n26717 );
    xnor g35307 ( n10252 , n29715 , n4962 );
    and g35308 ( n14375 , n8354 , n2204 );
    or g35309 ( n5834 , n31906 , n18686 );
    nor g35310 ( n29491 , n18514 , n29203 );
    or g35311 ( n25624 , n9658 , n8948 );
    or g35312 ( n19498 , n28210 , n20817 );
    or g35313 ( n13116 , n23466 , n33435 );
    or g35314 ( n23050 , n25337 , n5338 );
    or g35315 ( n7376 , n23275 , n2834 );
    and g35316 ( n8022 , n32710 , n14525 );
    not g35317 ( n35883 , n22495 );
    xnor g35318 ( n502 , n4757 , n35927 );
    nor g35319 ( n6113 , n17568 , n10197 );
    not g35320 ( n27695 , n7726 );
    or g35321 ( n29137 , n31181 , n31312 );
    xnor g35322 ( n34118 , n22932 , n16135 );
    or g35323 ( n20740 , n22975 , n763 );
    and g35324 ( n3371 , n9567 , n30891 );
    xnor g35325 ( n6274 , n18309 , n382 );
    and g35326 ( n28198 , n21685 , n14753 );
    nor g35327 ( n14276 , n4962 , n20044 );
    nor g35328 ( n17811 , n3205 , n6054 );
    and g35329 ( n7256 , n9203 , n32097 );
    and g35330 ( n24360 , n33323 , n33083 );
    or g35331 ( n19625 , n18382 , n14516 );
    xnor g35332 ( n4541 , n29269 , n10900 );
    nor g35333 ( n30748 , n32584 , n16692 );
    or g35334 ( n137 , n10349 , n29643 );
    and g35335 ( n14873 , n2731 , n13574 );
    or g35336 ( n4 , n4758 , n9288 );
    or g35337 ( n24484 , n16537 , n32354 );
    xnor g35338 ( n24350 , n687 , n19551 );
    or g35339 ( n35725 , n17404 , n17150 );
    and g35340 ( n31417 , n20259 , n25344 );
    xnor g35341 ( n2815 , n4044 , n30742 );
    and g35342 ( n33697 , n30267 , n12757 );
    or g35343 ( n8209 , n24514 , n8541 );
    and g35344 ( n12813 , n11399 , n27427 );
    or g35345 ( n30601 , n2589 , n18264 );
    and g35346 ( n9612 , n27371 , n27547 );
    not g35347 ( n27542 , n29079 );
    or g35348 ( n23911 , n34030 , n4254 );
    and g35349 ( n17446 , n802 , n30914 );
    not g35350 ( n11891 , n23604 );
    xnor g35351 ( n9901 , n11001 , n32095 );
    or g35352 ( n23329 , n28145 , n34413 );
    not g35353 ( n17926 , n20837 );
    xnor g35354 ( n16740 , n20155 , n17568 );
    or g35355 ( n18716 , n14609 , n17046 );
    or g35356 ( n26575 , n5735 , n19552 );
    and g35357 ( n22882 , n24993 , n15576 );
    or g35358 ( n13665 , n27169 , n4595 );
    or g35359 ( n27189 , n34324 , n24069 );
    or g35360 ( n26178 , n24371 , n36090 );
    and g35361 ( n33044 , n26645 , n3646 );
    or g35362 ( n16928 , n8432 , n25835 );
    xnor g35363 ( n17918 , n28070 , n17568 );
    buf g35364 ( n34862 , n25648 );
    or g35365 ( n14919 , n13329 , n21042 );
    or g35366 ( n11393 , n32907 , n239 );
    or g35367 ( n12762 , n8821 , n25940 );
    nor g35368 ( n32758 , n30814 , n33157 );
    and g35369 ( n22236 , n13839 , n15522 );
    or g35370 ( n9898 , n2618 , n8959 );
    or g35371 ( n7387 , n34275 , n17810 );
    nor g35372 ( n4853 , n2172 , n9336 );
    xnor g35373 ( n26035 , n23824 , n34816 );
    or g35374 ( n8391 , n23507 , n27895 );
    xnor g35375 ( n9518 , n25684 , n9658 );
    and g35376 ( n22270 , n33377 , n7952 );
    not g35377 ( n13196 , n21906 );
    xnor g35378 ( n11592 , n22810 , n370 );
    nor g35379 ( n32356 , n32325 , n19336 );
    xor g35380 ( n29316 , n13265 , n10998 );
    not g35381 ( n14636 , n2067 );
    not g35382 ( n13203 , n30459 );
    or g35383 ( n20093 , n12101 , n15216 );
    xnor g35384 ( n2459 , n35171 , n32095 );
    and g35385 ( n24928 , n1166 , n13360 );
    or g35386 ( n3159 , n20435 , n20654 );
    xnor g35387 ( n24863 , n20032 , n25602 );
    nor g35388 ( n5708 , n9789 , n18309 );
    nor g35389 ( n18933 , n34231 , n36040 );
    or g35390 ( n33813 , n26515 , n12950 );
    xnor g35391 ( n18279 , n14789 , n1950 );
    and g35392 ( n9760 , n14853 , n30203 );
    or g35393 ( n15786 , n17022 , n14436 );
    and g35394 ( n27242 , n17874 , n1696 );
    or g35395 ( n24993 , n3959 , n24505 );
    or g35396 ( n6329 , n7618 , n13305 );
    and g35397 ( n34842 , n3941 , n6208 );
    or g35398 ( n13155 , n22594 , n2438 );
    not g35399 ( n31397 , n9793 );
    or g35400 ( n12981 , n5660 , n17612 );
    or g35401 ( n17843 , n25384 , n1942 );
    and g35402 ( n34064 , n26054 , n25829 );
    nor g35403 ( n11244 , n32095 , n13046 );
    buf g35404 ( n30732 , n2866 );
    or g35405 ( n14302 , n33167 , n34923 );
    or g35406 ( n19676 , n894 , n11295 );
    or g35407 ( n10810 , n31289 , n17487 );
    or g35408 ( n31292 , n4288 , n1718 );
    or g35409 ( n10106 , n23068 , n10634 );
    and g35410 ( n31680 , n23561 , n10414 );
    or g35411 ( n15726 , n10485 , n24025 );
    and g35412 ( n13872 , n18818 , n23298 );
    or g35413 ( n17266 , n31973 , n25648 );
    or g35414 ( n9935 , n34661 , n15109 );
    not g35415 ( n35321 , n22980 );
    xnor g35416 ( n31460 , n34853 , n32715 );
    or g35417 ( n4326 , n5335 , n23485 );
    and g35418 ( n17915 , n24323 , n17836 );
    or g35419 ( n11385 , n28744 , n2119 );
    or g35420 ( n22204 , n17066 , n8004 );
    or g35421 ( n13169 , n6571 , n11258 );
    and g35422 ( n15884 , n29710 , n34101 );
    not g35423 ( n5923 , n16808 );
    or g35424 ( n3203 , n2948 , n16543 );
    or g35425 ( n35466 , n35754 , n22591 );
    or g35426 ( n3161 , n35687 , n14407 );
    and g35427 ( n20067 , n1947 , n3453 );
    not g35428 ( n9071 , n2029 );
    and g35429 ( n31850 , n5620 , n14023 );
    xnor g35430 ( n30952 , n13759 , n3605 );
    xnor g35431 ( n6626 , n14201 , n28995 );
    or g35432 ( n633 , n16002 , n9921 );
    xnor g35433 ( n11432 , n33173 , n4878 );
    or g35434 ( n20678 , n15283 , n15445 );
    nor g35435 ( n17425 , n32095 , n33632 );
    or g35436 ( n2339 , n21882 , n10309 );
    not g35437 ( n21914 , n26112 );
    xnor g35438 ( n21845 , n9842 , n27454 );
    and g35439 ( n21037 , n31228 , n21412 );
    or g35440 ( n20057 , n4327 , n34216 );
    not g35441 ( n19992 , n3222 );
    not g35442 ( n28584 , n5180 );
    or g35443 ( n22433 , n9102 , n901 );
    not g35444 ( n2666 , n35981 );
    or g35445 ( n16869 , n4878 , n6033 );
    or g35446 ( n5734 , n24858 , n32608 );
    xnor g35447 ( n17419 , n34083 , n31491 );
    and g35448 ( n33357 , n26533 , n2038 );
    and g35449 ( n17379 , n1631 , n31035 );
    xnor g35450 ( n25871 , n2161 , n8453 );
    or g35451 ( n24077 , n5335 , n17699 );
    or g35452 ( n28287 , n4075 , n2536 );
    and g35453 ( n24341 , n19598 , n18640 );
    buf g35454 ( n27580 , n31100 );
    or g35455 ( n34055 , n1960 , n23090 );
    or g35456 ( n12954 , n7807 , n32634 );
    not g35457 ( n28102 , n31300 );
    and g35458 ( n31310 , n28724 , n12878 );
    or g35459 ( n22205 , n11336 , n1414 );
    or g35460 ( n20839 , n11910 , n33098 );
    or g35461 ( n19912 , n16666 , n2524 );
    and g35462 ( n5243 , n23842 , n27731 );
    or g35463 ( n4315 , n14641 , n24018 );
    or g35464 ( n1825 , n5487 , n36027 );
    or g35465 ( n22600 , n21816 , n26468 );
    xnor g35466 ( n13329 , n21350 , n26081 );
    or g35467 ( n13039 , n34860 , n12529 );
    or g35468 ( n26607 , n4962 , n770 );
    and g35469 ( n15740 , n6057 , n17 );
    xnor g35470 ( n11949 , n31101 , n29448 );
    or g35471 ( n30643 , n22502 , n18899 );
    or g35472 ( n28080 , n7199 , n10537 );
    or g35473 ( n28876 , n33792 , n8724 );
    and g35474 ( n19796 , n9863 , n30339 );
    or g35475 ( n1776 , n1229 , n1176 );
    xnor g35476 ( n11285 , n32822 , n29713 );
    or g35477 ( n23370 , n33459 , n139 );
    not g35478 ( n33759 , n7141 );
    xnor g35479 ( n19695 , n35827 , n3222 );
    or g35480 ( n18726 , n24512 , n3568 );
    and g35481 ( n4185 , n17954 , n35013 );
    or g35482 ( n29971 , n26137 , n1763 );
    or g35483 ( n24425 , n14694 , n6064 );
    xnor g35484 ( n15342 , n34109 , n35913 );
    or g35485 ( n30063 , n33875 , n25773 );
    not g35486 ( n6479 , n2910 );
    or g35487 ( n343 , n6405 , n33098 );
    or g35488 ( n2550 , n29150 , n11357 );
    xnor g35489 ( n19624 , n23597 , n23566 );
    and g35490 ( n23064 , n25321 , n22098 );
    or g35491 ( n5141 , n3050 , n27447 );
    nor g35492 ( n4756 , n9789 , n23612 );
    nor g35493 ( n6618 , n26888 , n19957 );
    or g35494 ( n10026 , n30923 , n11996 );
    or g35495 ( n32044 , n29338 , n29368 );
    and g35496 ( n33036 , n32112 , n6058 );
    and g35497 ( n25189 , n18206 , n8433 );
    or g35498 ( n14511 , n24371 , n17901 );
    or g35499 ( n3648 , n9789 , n9467 );
    or g35500 ( n31218 , n16711 , n17354 );
    or g35501 ( n13199 , n17219 , n8924 );
    and g35502 ( n22951 , n6637 , n22473 );
    xnor g35503 ( n25047 , n4954 , n9146 );
    or g35504 ( n31483 , n10288 , n14699 );
    or g35505 ( n33930 , n11455 , n27980 );
    xnor g35506 ( n35002 , n12095 , n11896 );
    or g35507 ( n13118 , n15165 , n34103 );
    or g35508 ( n6803 , n27104 , n8203 );
    and g35509 ( n850 , n25769 , n21784 );
    nor g35510 ( n30219 , n11314 , n31411 );
    xnor g35511 ( n17247 , n21357 , n1232 );
    and g35512 ( n5145 , n6846 , n19868 );
    or g35513 ( n7541 , n22291 , n12498 );
    or g35514 ( n3902 , n30985 , n28969 );
    and g35515 ( n8215 , n2054 , n35544 );
    xnor g35516 ( n24328 , n28932 , n35296 );
    and g35517 ( n27966 , n28657 , n26665 );
    or g35518 ( n34028 , n14081 , n18598 );
    or g35519 ( n30220 , n14993 , n14361 );
    or g35520 ( n35047 , n17171 , n11737 );
    or g35521 ( n3189 , n30960 , n17354 );
    and g35522 ( n621 , n17697 , n4067 );
    nor g35523 ( n34375 , n24191 , n32666 );
    or g35524 ( n283 , n34760 , n16621 );
    or g35525 ( n35600 , n4642 , n34472 );
    xnor g35526 ( n34371 , n22574 , n9789 );
    and g35527 ( n17754 , n6112 , n29550 );
    or g35528 ( n2901 , n7285 , n8063 );
    xnor g35529 ( n17890 , n23916 , n15464 );
    and g35530 ( n4016 , n4768 , n218 );
    and g35531 ( n7232 , n15937 , n34492 );
    or g35532 ( n21320 , n27673 , n14365 );
    xnor g35533 ( n11919 , n681 , n31056 );
    not g35534 ( n1247 , n4235 );
    or g35535 ( n265 , n10334 , n4422 );
    or g35536 ( n16368 , n29209 , n9394 );
    or g35537 ( n6850 , n33207 , n10801 );
    and g35538 ( n4335 , n12390 , n12614 );
    or g35539 ( n27576 , n3816 , n18921 );
    or g35540 ( n26241 , n17952 , n914 );
    or g35541 ( n23668 , n8797 , n12431 );
    and g35542 ( n11771 , n21139 , n6574 );
    and g35543 ( n12850 , n14480 , n13173 );
    or g35544 ( n659 , n33788 , n25990 );
    or g35545 ( n19262 , n25174 , n27615 );
    or g35546 ( n35617 , n10894 , n16959 );
    and g35547 ( n6370 , n16998 , n2086 );
    and g35548 ( n18636 , n8067 , n3010 );
    or g35549 ( n34357 , n11914 , n8723 );
    or g35550 ( n21838 , n19568 , n1942 );
    not g35551 ( n15226 , n4609 );
    and g35552 ( n17054 , n18086 , n23814 );
    or g35553 ( n22709 , n19984 , n4995 );
    and g35554 ( n7666 , n7244 , n13026 );
    or g35555 ( n14587 , n2564 , n31627 );
    or g35556 ( n20116 , n1950 , n20206 );
    xnor g35557 ( n15155 , n15559 , n7540 );
    xnor g35558 ( n8699 , n19163 , n3091 );
    and g35559 ( n13482 , n26718 , n21861 );
    xnor g35560 ( n3250 , n23727 , n6326 );
    or g35561 ( n26850 , n14658 , n17951 );
    and g35562 ( n21010 , n34757 , n25069 );
    or g35563 ( n16363 , n19518 , n3096 );
    and g35564 ( n863 , n22983 , n1400 );
    xnor g35565 ( n28133 , n19875 , n24371 );
    or g35566 ( n34389 , n30576 , n35043 );
    nor g35567 ( n23258 , n26067 , n28680 );
    or g35568 ( n5673 , n3976 , n29953 );
    xnor g35569 ( n29625 , n5793 , n5674 );
    xnor g35570 ( n19751 , n782 , n1689 );
    not g35571 ( n10063 , n3527 );
    and g35572 ( n13667 , n3309 , n13324 );
    or g35573 ( n22699 , n353 , n11690 );
    or g35574 ( n8547 , n25108 , n13540 );
    and g35575 ( n15110 , n22231 , n19729 );
    xnor g35576 ( n24326 , n4997 , n17568 );
    xnor g35577 ( n26846 , n8440 , n32715 );
    or g35578 ( n18024 , n7248 , n13301 );
    xnor g35579 ( n10771 , n22999 , n34075 );
    or g35580 ( n7482 , n22291 , n27989 );
    xnor g35581 ( n3635 , n23519 , n10380 );
    xnor g35582 ( n3900 , n10485 , n24371 );
    or g35583 ( n34882 , n12548 , n28248 );
    or g35584 ( n20728 , n22186 , n4700 );
    or g35585 ( n25303 , n32442 , n25255 );
    and g35586 ( n449 , n18614 , n5622 );
    or g35587 ( n19941 , n2113 , n21453 );
    not g35588 ( n11243 , n35570 );
    not g35589 ( n33206 , n21398 );
    xnor g35590 ( n3456 , n7597 , n28789 );
    or g35591 ( n3775 , n17267 , n31554 );
    nor g35592 ( n1630 , n31371 , n13824 );
    or g35593 ( n23966 , n26551 , n27973 );
    not g35594 ( n30982 , n1178 );
    xnor g35595 ( n13496 , n737 , n8066 );
    xnor g35596 ( n5307 , n3578 , n2971 );
    or g35597 ( n28253 , n21588 , n14689 );
    or g35598 ( n26218 , n29912 , n18265 );
    or g35599 ( n13582 , n11047 , n3936 );
    or g35600 ( n30000 , n9658 , n684 );
    and g35601 ( n5670 , n9466 , n6600 );
    not g35602 ( n33793 , n33890 );
    xnor g35603 ( n16494 , n17072 , n803 );
    not g35604 ( n11040 , n27269 );
    not g35605 ( n14824 , n11200 );
    or g35606 ( n22319 , n7155 , n31632 );
    nor g35607 ( n24512 , n18151 , n34484 );
    nor g35608 ( n10016 , n13224 , n16557 );
    or g35609 ( n7372 , n14912 , n31773 );
    nor g35610 ( n31312 , n3830 , n32484 );
    and g35611 ( n24897 , n28803 , n10515 );
    or g35612 ( n33748 , n15654 , n9398 );
    xnor g35613 ( n18695 , n30188 , n3262 );
    or g35614 ( n27744 , n31760 , n6473 );
    not g35615 ( n17220 , n30589 );
    and g35616 ( n17227 , n27901 , n18671 );
    xnor g35617 ( n10192 , n4179 , n4878 );
    or g35618 ( n4274 , n6960 , n4175 );
    xnor g35619 ( n32823 , n2544 , n50 );
    or g35620 ( n32343 , n5738 , n32229 );
    nor g35621 ( n18650 , n3778 , n32422 );
    or g35622 ( n24632 , n27657 , n35748 );
    not g35623 ( n3639 , n12348 );
    and g35624 ( n23500 , n22762 , n12339 );
    xnor g35625 ( n22453 , n9387 , n10894 );
    not g35626 ( n9003 , n30586 );
    or g35627 ( n8828 , n30742 , n21802 );
    and g35628 ( n19499 , n4986 , n12405 );
    xnor g35629 ( n18336 , n1229 , n30553 );
    and g35630 ( n18399 , n34479 , n19390 );
    buf g35631 ( n12428 , n16814 );
    or g35632 ( n26964 , n8774 , n667 );
    or g35633 ( n34998 , n13338 , n19058 );
    xnor g35634 ( n22735 , n33897 , n17408 );
    not g35635 ( n21959 , n12852 );
    and g35636 ( n34373 , n29446 , n11444 );
    xnor g35637 ( n34068 , n2055 , n30763 );
    or g35638 ( n17374 , n7884 , n27704 );
    or g35639 ( n20672 , n8368 , n20817 );
    xnor g35640 ( n25992 , n25523 , n25524 );
    xnor g35641 ( n1068 , n23848 , n24329 );
    xnor g35642 ( n18504 , n27910 , n30140 );
    or g35643 ( n13997 , n25561 , n26393 );
    or g35644 ( n33617 , n9816 , n10336 );
    and g35645 ( n5116 , n18290 , n35161 );
    xnor g35646 ( n30018 , n5263 , n1950 );
    not g35647 ( n19508 , n28719 );
    or g35648 ( n23617 , n35921 , n11472 );
    xnor g35649 ( n13636 , n12657 , n34607 );
    not g35650 ( n12261 , n30181 );
    and g35651 ( n23521 , n24561 , n18648 );
    or g35652 ( n6566 , n1950 , n33412 );
    and g35653 ( n15756 , n28435 , n325 );
    xnor g35654 ( n29671 , n22066 , n35909 );
    and g35655 ( n22749 , n13399 , n22710 );
    and g35656 ( n7309 , n34633 , n14922 );
    xnor g35657 ( n14166 , n9684 , n4878 );
    and g35658 ( n5189 , n14543 , n3796 );
    and g35659 ( n34938 , n21244 , n15494 );
    and g35660 ( n16738 , n20998 , n18288 );
    xnor g35661 ( n5102 , n19059 , n27590 );
    or g35662 ( n32047 , n11455 , n7990 );
    and g35663 ( n25035 , n32962 , n13120 );
    and g35664 ( n7919 , n13214 , n21737 );
    xnor g35665 ( n19405 , n22285 , n6929 );
    and g35666 ( n151 , n748 , n21987 );
    or g35667 ( n24925 , n10441 , n6002 );
    xnor g35668 ( n5316 , n3174 , n11190 );
    or g35669 ( n14061 , n17566 , n26220 );
    or g35670 ( n33756 , n4638 , n16579 );
    or g35671 ( n26576 , n32437 , n1557 );
    and g35672 ( n9241 , n23709 , n18611 );
    or g35673 ( n25856 , n18520 , n3239 );
    or g35674 ( n28928 , n22791 , n6683 );
    nor g35675 ( n15653 , n13861 , n18113 );
    and g35676 ( n19353 , n2787 , n6016 );
    or g35677 ( n10297 , n27729 , n27689 );
    or g35678 ( n21241 , n7367 , n32808 );
    xnor g35679 ( n9371 , n31720 , n30057 );
    or g35680 ( n32411 , n8500 , n29587 );
    and g35681 ( n7215 , n13707 , n21973 );
    or g35682 ( n24203 , n27226 , n29080 );
    not g35683 ( n35498 , n35941 );
    or g35684 ( n1444 , n17926 , n34546 );
    or g35685 ( n26240 , n27226 , n1645 );
    xnor g35686 ( n17159 , n4247 , n6470 );
    and g35687 ( n4269 , n8853 , n31304 );
    or g35688 ( n18568 , n12993 , n544 );
    nor g35689 ( n26980 , n19551 , n19425 );
    or g35690 ( n8448 , n19236 , n8600 );
    xnor g35691 ( n16935 , n12554 , n27226 );
    xnor g35692 ( n21896 , n32519 , n18954 );
    and g35693 ( n1706 , n27898 , n2238 );
    and g35694 ( n35722 , n27733 , n18362 );
    or g35695 ( n32311 , n4785 , n2479 );
    or g35696 ( n34903 , n30744 , n27394 );
    and g35697 ( n4710 , n29040 , n33339 );
    or g35698 ( n10684 , n35916 , n14699 );
    and g35699 ( n24646 , n35226 , n1828 );
    or g35700 ( n29299 , n26060 , n9875 );
    or g35701 ( n12182 , n7540 , n9862 );
    xnor g35702 ( n26093 , n24873 , n21130 );
    xnor g35703 ( n6870 , n7990 , n11455 );
    or g35704 ( n16118 , n23648 , n29562 );
    or g35705 ( n14498 , n26158 , n21560 );
    or g35706 ( n30020 , n860 , n13652 );
    or g35707 ( n28832 , n22425 , n5900 );
    and g35708 ( n1451 , n16440 , n13432 );
    or g35709 ( n28723 , n2991 , n10432 );
    or g35710 ( n15484 , n6907 , n2524 );
    xnor g35711 ( n7999 , n15037 , n4288 );
    or g35712 ( n21640 , n22784 , n17337 );
    nor g35713 ( n25917 , n10894 , n11159 );
    xnor g35714 ( n16991 , n22514 , n29713 );
    or g35715 ( n14526 , n10894 , n16696 );
    or g35716 ( n16629 , n24332 , n34676 );
    and g35717 ( n31704 , n13155 , n9695 );
    xnor g35718 ( n27062 , n6123 , n24412 );
    and g35719 ( n24779 , n731 , n13078 );
    or g35720 ( n30446 , n4878 , n9549 );
    xnor g35721 ( n7519 , n24764 , n16388 );
    or g35722 ( n34964 , n27077 , n34923 );
    xnor g35723 ( n292 , n28917 , n3946 );
    xnor g35724 ( n11603 , n10639 , n20340 );
    and g35725 ( n18891 , n21041 , n7768 );
    or g35726 ( n9880 , n12346 , n3308 );
    or g35727 ( n13001 , n23121 , n35757 );
    and g35728 ( n31124 , n14645 , n16276 );
    or g35729 ( n3499 , n4728 , n21579 );
    or g35730 ( n17073 , n4147 , n24928 );
    and g35731 ( n23254 , n9945 , n18907 );
    not g35732 ( n2492 , n22291 );
    or g35733 ( n12550 , n10928 , n5061 );
    or g35734 ( n22927 , n21464 , n28064 );
    and g35735 ( n27793 , n11370 , n26334 );
    xnor g35736 ( n35999 , n15166 , n11029 );
    xnor g35737 ( n7027 , n29367 , n29959 );
    xnor g35738 ( n12639 , n31782 , n22291 );
    or g35739 ( n9497 , n246 , n21579 );
    or g35740 ( n24910 , n23233 , n26659 );
    or g35741 ( n6385 , n8978 , n5618 );
    or g35742 ( n28786 , n11190 , n24457 );
    and g35743 ( n7909 , n7058 , n31448 );
    not g35744 ( n19566 , n31990 );
    not g35745 ( n23524 , n4878 );
    xnor g35746 ( n13512 , n12735 , n30780 );
    or g35747 ( n30956 , n32584 , n15474 );
    xnor g35748 ( n32158 , n25368 , n16922 );
    xnor g35749 ( n22406 , n22777 , n24051 );
    xnor g35750 ( n18546 , n34671 , n3465 );
    or g35751 ( n30550 , n28984 , n26220 );
    xnor g35752 ( n21927 , n10829 , n31215 );
    or g35753 ( n6152 , n35459 , n16747 );
    or g35754 ( n33623 , n3946 , n2770 );
    xnor g35755 ( n6137 , n12102 , n9947 );
    xnor g35756 ( n10500 , n35743 , n24003 );
    and g35757 ( n16777 , n29019 , n9866 );
    and g35758 ( n10149 , n11804 , n20168 );
    xnor g35759 ( n21279 , n25416 , n3501 );
    xnor g35760 ( n31570 , n143 , n28475 );
    or g35761 ( n33937 , n17942 , n19125 );
    nor g35762 ( n25108 , n4878 , n32707 );
    and g35763 ( n20616 , n19689 , n8320 );
    nor g35764 ( n6844 , n4758 , n14000 );
    or g35765 ( n10874 , n6371 , n21644 );
    not g35766 ( n29166 , n23622 );
    xnor g35767 ( n10371 , n29311 , n7540 );
    nor g35768 ( n4244 , n27839 , n14274 );
    or g35769 ( n11376 , n30742 , n25465 );
    not g35770 ( n14068 , n7437 );
    and g35771 ( n7925 , n497 , n17277 );
    xnor g35772 ( n27005 , n22402 , n1950 );
    and g35773 ( n10540 , n19641 , n32798 );
    and g35774 ( n14907 , n19913 , n15401 );
    not g35775 ( n16179 , n28032 );
    not g35776 ( n6306 , n3858 );
    nor g35777 ( n11735 , n1833 , n6548 );
    or g35778 ( n7942 , n27550 , n19353 );
    or g35779 ( n5526 , n33676 , n25392 );
    or g35780 ( n21270 , n10098 , n26220 );
    xnor g35781 ( n9940 , n110 , n20676 );
    or g35782 ( n34906 , n13121 , n26659 );
    nor g35783 ( n7580 , n10894 , n15429 );
    or g35784 ( n33337 , n18180 , n25786 );
    xnor g35785 ( n2334 , n1228 , n24371 );
    or g35786 ( n24169 , n5228 , n25080 );
    xnor g35787 ( n6262 , n34650 , n31370 );
    not g35788 ( n1198 , n22471 );
    and g35789 ( n16330 , n9171 , n6989 );
    or g35790 ( n21329 , n34664 , n27501 );
    and g35791 ( n4753 , n28650 , n17459 );
    xnor g35792 ( n21115 , n34118 , n3537 );
    xnor g35793 ( n35641 , n17642 , n32584 );
    and g35794 ( n27742 , n13510 , n25117 );
    or g35795 ( n27421 , n31501 , n27086 );
    not g35796 ( n28852 , n31799 );
    and g35797 ( n28490 , n726 , n8251 );
    or g35798 ( n17849 , n9255 , n8203 );
    and g35799 ( n1060 , n7718 , n14614 );
    or g35800 ( n35577 , n161 , n31243 );
    and g35801 ( n33448 , n29199 , n11662 );
    or g35802 ( n3868 , n32822 , n33310 );
    and g35803 ( n5565 , n33872 , n7551 );
    and g35804 ( n24929 , n809 , n30494 );
    or g35805 ( n8990 , n30899 , n4203 );
    and g35806 ( n28440 , n23329 , n17380 );
    or g35807 ( n30428 , n4758 , n29188 );
    or g35808 ( n27141 , n34878 , n9921 );
    nor g35809 ( n20991 , n27100 , n18115 );
    not g35810 ( n1274 , n8432 );
    and g35811 ( n772 , n9270 , n21854 );
    or g35812 ( n33809 , n28929 , n11752 );
    and g35813 ( n24868 , n5037 , n17930 );
    not g35814 ( n8724 , n18296 );
    xnor g35815 ( n6662 , n11049 , n25226 );
    xnor g35816 ( n12212 , n10437 , n32857 );
    and g35817 ( n19614 , n18996 , n34752 );
    xnor g35818 ( n3511 , n36077 , n30183 );
    xnor g35819 ( n14755 , n9193 , n23769 );
    and g35820 ( n7075 , n13926 , n20847 );
    xnor g35821 ( n29736 , n11338 , n16922 );
    or g35822 ( n23048 , n26608 , n25355 );
    and g35823 ( n23801 , n23639 , n17371 );
    and g35824 ( n4997 , n20665 , n4431 );
    and g35825 ( n20059 , n24831 , n29598 );
    or g35826 ( n17003 , n20858 , n32634 );
    xnor g35827 ( n16238 , n22154 , n32857 );
    and g35828 ( n31231 , n12710 , n2596 );
    xnor g35829 ( n2587 , n28770 , n4288 );
    and g35830 ( n8221 , n26923 , n5776 );
    or g35831 ( n14893 , n28325 , n4203 );
    not g35832 ( n16723 , n4776 );
    and g35833 ( n20177 , n12287 , n25168 );
    or g35834 ( n3507 , n13139 , n14950 );
    or g35835 ( n25844 , n15986 , n12791 );
    nor g35836 ( n33738 , n19268 , n3958 );
    xnor g35837 ( n14658 , n15890 , n16922 );
    and g35838 ( n11224 , n24904 , n27287 );
    and g35839 ( n28695 , n5329 , n22694 );
    or g35840 ( n29314 , n4002 , n32278 );
    or g35841 ( n7665 , n18367 , n33698 );
    xnor g35842 ( n5604 , n33533 , n31799 );
    or g35843 ( n20639 , n31436 , n21002 );
    or g35844 ( n7415 , n35432 , n22316 );
    and g35845 ( n22632 , n10874 , n23226 );
    or g35846 ( n1110 , n32190 , n28064 );
    or g35847 ( n28595 , n823 , n19125 );
    or g35848 ( n25598 , n15829 , n25355 );
    or g35849 ( n10496 , n17798 , n6374 );
    and g35850 ( n7014 , n26338 , n13001 );
    or g35851 ( n20673 , n32055 , n21328 );
    or g35852 ( n32620 , n10377 , n23282 );
    xnor g35853 ( n29784 , n13489 , n3356 );
    or g35854 ( n27788 , n8834 , n22322 );
    or g35855 ( n20695 , n15580 , n9709 );
    or g35856 ( n34256 , n15886 , n1079 );
    and g35857 ( n24905 , n18134 , n4891 );
    xnor g35858 ( n8793 , n21234 , n22291 );
    and g35859 ( n31363 , n3247 , n14538 );
    or g35860 ( n19479 , n15247 , n11409 );
    or g35861 ( n5254 , n27688 , n27447 );
    or g35862 ( n14026 , n24171 , n1763 );
    or g35863 ( n4828 , n2998 , n4318 );
    or g35864 ( n32499 , n1950 , n31149 );
    not g35865 ( n29359 , n31893 );
    or g35866 ( n21929 , n1403 , n35935 );
    or g35867 ( n2244 , n4480 , n36085 );
    nor g35868 ( n32313 , n3630 , n4912 );
    and g35869 ( n19643 , n13304 , n35054 );
    or g35870 ( n29354 , n19572 , n15439 );
    or g35871 ( n13279 , n13708 , n25786 );
    and g35872 ( n28465 , n11651 , n25011 );
    not g35873 ( n21785 , n3842 );
    and g35874 ( n24419 , n8645 , n19110 );
    xnor g35875 ( n25216 , n33104 , n23828 );
    or g35876 ( n16754 , n20768 , n32329 );
    or g35877 ( n2631 , n29713 , n35150 );
    and g35878 ( n12413 , n5645 , n7449 );
    and g35879 ( n23325 , n31373 , n35946 );
    or g35880 ( n29477 , n25602 , n19796 );
    or g35881 ( n6920 , n17772 , n26292 );
    not g35882 ( n32203 , n17131 );
    or g35883 ( n27417 , n8505 , n30721 );
    and g35884 ( n6561 , n22155 , n30048 );
    not g35885 ( n30978 , n18296 );
    or g35886 ( n9708 , n26664 , n30252 );
    or g35887 ( n11030 , n7632 , n17893 );
    xnor g35888 ( n27937 , n19536 , n15513 );
    or g35889 ( n29070 , n3158 , n4053 );
    nor g35890 ( n21804 , n4960 , n8187 );
    and g35891 ( n15024 , n23657 , n2050 );
    or g35892 ( n30892 , n7296 , n966 );
    xnor g35893 ( n4447 , n34529 , n13553 );
    and g35894 ( n31535 , n21689 , n6039 );
    not g35895 ( n30229 , n34209 );
    and g35896 ( n25106 , n18223 , n20975 );
    and g35897 ( n34229 , n9540 , n21098 );
    or g35898 ( n26520 , n34383 , n27437 );
    or g35899 ( n3447 , n12115 , n15145 );
    and g35900 ( n24819 , n11883 , n8759 );
    xnor g35901 ( n26348 , n22578 , n9789 );
    or g35902 ( n7556 , n23768 , n21223 );
    or g35903 ( n22902 , n29160 , n29592 );
    or g35904 ( n33724 , n11190 , n10885 );
    or g35905 ( n10746 , n16234 , n30076 );
    or g35906 ( n4548 , n4960 , n26001 );
    and g35907 ( n31758 , n6549 , n133 );
    not g35908 ( n19163 , n32861 );
    not g35909 ( n10952 , n12301 );
    or g35910 ( n17792 , n15824 , n3979 );
    not g35911 ( n27568 , n8691 );
    or g35912 ( n27789 , n20682 , n24538 );
    buf g35913 ( n28324 , n33464 );
    and g35914 ( n26419 , n14370 , n7600 );
    xnor g35915 ( n24098 , n23711 , n1950 );
    nor g35916 ( n28742 , n18349 , n32875 );
    or g35917 ( n15687 , n19984 , n15128 );
    not g35918 ( n18407 , n12428 );
    and g35919 ( n33887 , n27845 , n31129 );
    or g35920 ( n8126 , n2911 , n11372 );
    or g35921 ( n23775 , n33411 , n13664 );
    xnor g35922 ( n21830 , n23315 , n4288 );
    nor g35923 ( n34945 , n13204 , n14727 );
    xnor g35924 ( n15702 , n27806 , n28440 );
    and g35925 ( n9450 , n485 , n10446 );
    xnor g35926 ( n7100 , n8960 , n21999 );
    or g35927 ( n30929 , n10302 , n21839 );
    or g35928 ( n24065 , n3205 , n29038 );
    not g35929 ( n27912 , n16620 );
    nor g35930 ( n15112 , n30615 , n19501 );
    or g35931 ( n7133 , n6240 , n34583 );
    not g35932 ( n4844 , n25648 );
    and g35933 ( n225 , n31631 , n605 );
    and g35934 ( n253 , n30135 , n4200 );
    or g35935 ( n21316 , n33497 , n32634 );
    or g35936 ( n35403 , n24590 , n22142 );
    nor g35937 ( n26143 , n20633 , n4522 );
    xnor g35938 ( n30212 , n8498 , n9658 );
    and g35939 ( n32088 , n1923 , n29646 );
    or g35940 ( n11088 , n23030 , n27447 );
    xnor g35941 ( n20419 , n26258 , n32584 );
    or g35942 ( n5636 , n21982 , n12791 );
    or g35943 ( n15674 , n1423 , n20300 );
    or g35944 ( n25754 , n1950 , n22402 );
    xnor g35945 ( n22163 , n26175 , n3222 );
    xnor g35946 ( n20985 , n8167 , n9789 );
    and g35947 ( n14789 , n12970 , n14416 );
    and g35948 ( n20571 , n29499 , n6153 );
    or g35949 ( n24401 , n4960 , n35392 );
    or g35950 ( n7595 , n11675 , n32608 );
    or g35951 ( n8301 , n29652 , n139 );
    or g35952 ( n20684 , n18625 , n27728 );
    or g35953 ( n6923 , n23985 , n12428 );
    not g35954 ( n1102 , n8725 );
    or g35955 ( n35562 , n15690 , n32808 );
    or g35956 ( n34752 , n4960 , n17746 );
    xnor g35957 ( n13572 , n32407 , n27226 );
    xnor g35958 ( n4553 , n24853 , n32095 );
    and g35959 ( n15713 , n1022 , n15211 );
    xnor g35960 ( n28166 , n10054 , n27663 );
    or g35961 ( n15646 , n647 , n19084 );
    or g35962 ( n7954 , n17953 , n16456 );
    nor g35963 ( n14376 , n14960 , n25952 );
endmodule
