module top( n0 , n2 , n17 , n18 , n23 , n24 , n26 , n27 , n29 , 
n37 , n43 , n58 , n59 , n61 , n66 , n70 , n73 , n75 , n80 , 
n81 , n84 , n86 , n88 , n89 , n90 , n91 , n94 , n98 , n104 , 
n107 , n123 , n129 , n130 , n133 , n137 , n145 , n151 , n160 , n164 , 
n168 , n169 , n174 , n179 , n187 , n194 , n196 , n199 , n210 , n211 , 
n212 , n213 , n214 , n217 , n221 , n226 , n234 , n237 , n238 , n246 , 
n249 , n253 , n256 , n260 , n261 , n265 , n272 , n278 , n281 , n286 , 
n289 , n292 , n304 , n310 );
    input n0 , n2 , n17 , n18 , n23 , n27 , n29 , n37 , n43 , 
n58 , n59 , n70 , n75 , n84 , n90 , n91 , n107 , n130 , n133 , 
n137 , n169 , n174 , n179 , n187 , n194 , n196 , n210 , n211 , n214 , 
n226 , n234 , n237 , n238 , n249 , n256 , n260 , n272 , n278 , n281 , 
n289 , n292 ;
    output n24 , n26 , n61 , n66 , n73 , n80 , n81 , n86 , n88 , 
n89 , n94 , n98 , n104 , n123 , n129 , n145 , n151 , n160 , n164 , 
n168 , n199 , n212 , n213 , n217 , n221 , n246 , n253 , n261 , n265 , 
n286 , n304 , n310 ;
    wire n1 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
n11 , n12 , n13 , n14 , n15 , n16 , n19 , n20 , n21 , n22 , 
n25 , n28 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n38 , 
n39 , n40 , n41 , n42 , n44 , n45 , n46 , n47 , n48 , n49 , 
n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n60 , n62 , 
n63 , n64 , n65 , n67 , n68 , n69 , n71 , n72 , n74 , n76 , 
n77 , n78 , n79 , n82 , n83 , n85 , n87 , n92 , n93 , n95 , 
n96 , n97 , n99 , n100 , n101 , n102 , n103 , n105 , n106 , n108 , 
n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , 
n119 , n120 , n121 , n122 , n124 , n125 , n126 , n127 , n128 , n131 , 
n132 , n134 , n135 , n136 , n138 , n139 , n140 , n141 , n142 , n143 , 
n144 , n146 , n147 , n148 , n149 , n150 , n152 , n153 , n154 , n155 , 
n156 , n157 , n158 , n159 , n161 , n162 , n163 , n165 , n166 , n167 , 
n170 , n171 , n172 , n173 , n175 , n176 , n177 , n178 , n180 , n181 , 
n182 , n183 , n184 , n185 , n186 , n188 , n189 , n190 , n191 , n192 , 
n193 , n195 , n197 , n198 , n200 , n201 , n202 , n203 , n204 , n205 , 
n206 , n207 , n208 , n209 , n215 , n216 , n218 , n219 , n220 , n222 , 
n223 , n224 , n225 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , 
n235 , n236 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n247 , 
n248 , n250 , n251 , n252 , n254 , n255 , n257 , n258 , n259 , n262 , 
n263 , n264 , n266 , n267 , n268 , n269 , n270 , n271 , n273 , n274 , 
n275 , n276 , n277 , n279 , n280 , n282 , n283 , n284 , n285 , n287 , 
n288 , n290 , n291 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
n300 , n301 , n302 , n303 , n305 , n306 , n307 , n308 , n309 , n311 ;
    xnor g0 ( n163 , n174 , n169 );
    xnor g1 ( n129 , n153 , n210 );
    or g2 ( n53 , n205 , n155 );
    or g3 ( n28 , n279 , n298 );
    xnor g4 ( n14 , n124 , n126 );
    xnor g5 ( n66 , n30 , n29 );
    or g6 ( n143 , n140 , n216 );
    or g7 ( n38 , n301 , n72 );
    xnor g8 ( n262 , n238 , n29 );
    not g9 ( n259 , n180 );
    or g10 ( n251 , n96 , n51 );
    xnor g11 ( n45 , n43 , n214 );
    xnor g12 ( n60 , n8 , n114 );
    or g13 ( n19 , n273 , n297 );
    xnor g14 ( n34 , n70 , n174 );
    or g15 ( n209 , n140 , n175 );
    or g16 ( n275 , n53 , n276 );
    xnor g17 ( n239 , n14 , n288 );
    xnor g18 ( n308 , n70 , n2 );
    or g19 ( n255 , n251 , n172 );
    or g20 ( n166 , n305 , n181 );
    or g21 ( n198 , n252 , n173 );
    xnor g22 ( n86 , n200 , n196 );
    or g23 ( n223 , n250 , n46 );
    or g24 ( n5 , n62 , n85 );
    or g25 ( n161 , n178 , n64 );
    not g26 ( n204 , n58 );
    xnor g27 ( n1 , n189 , n296 );
    not g28 ( n301 , n119 );
    or g29 ( n9 , n283 , n291 );
    xnor g30 ( n304 , n224 , n214 );
    xnor g31 ( n208 , n225 , n83 );
    or g32 ( n21 , n110 , n82 );
    xnor g33 ( n57 , n135 , n197 );
    xnor g34 ( n296 , n179 , n0 );
    or g35 ( n203 , n171 , n103 );
    or g36 ( n243 , n205 , n155 );
    xnor g37 ( n303 , n237 , n210 );
    xnor g38 ( n191 , n278 , n272 );
    not g39 ( n171 , n226 );
    xor g40 ( n233 , n149 , n309 );
    not g41 ( n140 , n78 );
    not g42 ( n279 , n119 );
    xnor g43 ( n63 , n130 , n107 );
    or g44 ( n220 , n235 , n274 );
    or g45 ( n65 , n128 , n68 );
    not g46 ( n103 , n281 );
    buf g47 ( n150 , n60 );
    xnor g48 ( n149 , n32 , n141 );
    or g49 ( n270 , n112 , n190 );
    or g50 ( n41 , n155 , n230 );
    xnor g51 ( n248 , n17 , n75 );
    or g52 ( n267 , n56 , n273 );
    or g53 ( n294 , n204 , n103 );
    or g54 ( n85 , n152 , n276 );
    or g55 ( n62 , n140 , n216 );
    or g56 ( n274 , n95 , n76 );
    xnor g57 ( n311 , n130 , n256 );
    xnor g58 ( n114 , n294 , n87 );
    xnor g59 ( n222 , n77 , n191 );
    or g60 ( n69 , n156 , n76 );
    or g61 ( n263 , n162 , n51 );
    xnor g62 ( n221 , n219 , n179 );
    or g63 ( n36 , n258 , n33 );
    xnor g64 ( n254 , n23 , n249 );
    xnor g65 ( n306 , n290 , n10 );
    not g66 ( n297 , n279 );
    xnor g67 ( n286 , n49 , n238 );
    xnor g68 ( n141 , n256 , n289 );
    or g69 ( n67 , n167 , n159 );
    xnor g70 ( n104 , n142 , n289 );
    xnor g71 ( n26 , n115 , n169 );
    or g72 ( n92 , n127 , n113 );
    or g73 ( n244 , n243 , n232 );
    or g74 ( n269 , n56 , n72 );
    or g75 ( n142 , n209 , n9 );
    xnor g76 ( n10 , n234 , n196 );
    or g77 ( n215 , n15 , n33 );
    not g78 ( n216 , n134 );
    or g79 ( n154 , n263 , n198 );
    or g80 ( n113 , n183 , n230 );
    or g81 ( n186 , n184 , n103 );
    or g82 ( n68 , n206 , n255 );
    not g83 ( n93 , n74 );
    xnor g84 ( n52 , n238 , n17 );
    or g85 ( n49 , n28 , n159 );
    or g86 ( n188 , n162 , n106 );
    or g87 ( n250 , n301 , n298 );
    or g88 ( n115 , n105 , n64 );
    xnor g89 ( n240 , n229 , n303 );
    or g90 ( n33 , n267 , n173 );
    xnor g91 ( n197 , n285 , n42 );
    xnor g92 ( n87 , n278 , n234 );
    xnor g93 ( n88 , n299 , n107 );
    xnor g94 ( n117 , n194 , n27 );
    xnor g95 ( n227 , n242 , n240 );
    xnor g96 ( n89 , n271 , n43 );
    xnor g97 ( n290 , n260 , n27 );
    or g98 ( n202 , n101 , n9 );
    or g99 ( n280 , n177 , n297 );
    not g100 ( n155 , n60 );
    or g101 ( n46 , n7 , n181 );
    or g102 ( n258 , n301 , n138 );
    xnor g103 ( n126 , n249 , n214 );
    not g104 ( n190 , n100 );
    or g105 ( n158 , n112 , n190 );
    not g106 ( n177 , n233 );
    or g107 ( n30 , n13 , n274 );
    not g108 ( n175 , n134 );
    or g109 ( n232 , n301 , n25 );
    or g110 ( n252 , n96 , n93 );
    or g111 ( n156 , n96 , n93 );
    xnor g112 ( n160 , n16 , n70 );
    or g113 ( n167 , n177 , n51 );
    or g114 ( n159 , n266 , n92 );
    or g115 ( n152 , n150 , n230 );
    or g116 ( n172 , n298 , n93 );
    xnor g117 ( n287 , n83 , n222 );
    or g118 ( n101 , n112 , n231 );
    or g119 ( n235 , n177 , n259 );
    xnor g120 ( n94 , n223 , n137 );
    xnor g121 ( n310 , n65 , n237 );
    or g122 ( n25 , n138 , n106 );
    or g123 ( n299 , n144 , n244 );
    or g124 ( n31 , n38 , n69 );
    xnor g125 ( n81 , n132 , n90 );
    or g126 ( n39 , n301 , n298 );
    not g127 ( n72 , n50 );
    not g128 ( n134 , n71 );
    xnor g129 ( n246 , n277 , n249 );
    xnor g130 ( n245 , n136 , n108 );
    or g131 ( n11 , n39 , n201 );
    not g132 ( n183 , n110 );
    not g133 ( n298 , n50 );
    not g134 ( n162 , n233 );
    xnor g135 ( n213 , n220 , n75 );
    or g136 ( n305 , n56 , n273 );
    not g137 ( n82 , n241 );
    xnor g138 ( n164 , n161 , n2 );
    xnor g139 ( n131 , n102 , n120 );
    xnor g140 ( n122 , n208 , n45 );
    or g141 ( n132 , n158 , n85 );
    or g142 ( n293 , n157 , n103 );
    or g143 ( n95 , n56 , n273 );
    buf g144 ( n205 , n57 );
    not g145 ( n257 , n91 );
    or g146 ( n148 , n112 , n41 );
    xnor g147 ( n120 , n187 , n211 );
    or g148 ( n283 , n205 , n155 );
    or g149 ( n99 , n307 , n147 );
    or g150 ( n284 , n55 , n46 );
    xnor g151 ( n6 , n306 , n222 );
    xnor g152 ( n73 , n284 , n260 );
    or g153 ( n178 , n112 , n231 );
    xor g154 ( n78 , n131 , n44 );
    or g155 ( n173 , n140 , n3 );
    xnor g156 ( n125 , n287 , n63 );
    xnor g157 ( n136 , n163 , n195 );
    xnor g158 ( n195 , n210 , n59 );
    or g159 ( n105 , n110 , n175 );
    or g160 ( n7 , n96 , n93 );
    xnor g161 ( n199 , n36 , n187 );
    or g162 ( n277 , n21 , n147 );
    xnor g163 ( n118 , n293 , n34 );
    xnor g164 ( n145 , n11 , n278 );
    xnor g165 ( n218 , n97 , n268 );
    or g166 ( n291 , n297 , n188 );
    xnor g167 ( n32 , n225 , n306 );
    xnor g168 ( n121 , n137 , n260 );
    or g169 ( n48 , n279 , n138 );
    or g170 ( n153 , n143 , n68 );
    xnor g171 ( n80 , n116 , n174 );
    or g172 ( n229 , n257 , n103 );
    xnor g173 ( n61 , n67 , n17 );
    xnor g174 ( n54 , n2 , n169 );
    or g175 ( n200 , n236 , n69 );
    buf g176 ( n96 , n227 );
    or g177 ( n193 , n150 , n230 );
    or g178 ( n176 , n280 , n166 );
    or g179 ( n185 , n162 , n297 );
    or g180 ( n128 , n112 , n183 );
    not g181 ( n100 , n78 );
    xnor g182 ( n24 , n5 , n59 );
    xnor g183 ( n77 , n137 , n194 );
    xnor g184 ( n207 , n29 , n75 );
    or g185 ( n276 , n269 , n19 );
    or g186 ( n139 , n96 , n93 );
    xnor g187 ( n212 , n99 , n23 );
    xnor g188 ( n217 , n202 , n256 );
    or g189 ( n302 , n185 , n201 );
    xnor g190 ( n146 , n179 , n187 );
    xnor g191 ( n268 , n90 , n59 );
    or g192 ( n206 , n150 , n230 );
    not g193 ( n230 , n57 );
    or g194 ( n12 , n241 , n183 );
    or g195 ( n3 , n82 , n41 );
    or g196 ( n109 , n47 , n232 );
    or g197 ( n236 , n162 , n259 );
    xnor g198 ( n135 , n239 , n207 );
    or g199 ( n47 , n150 , n230 );
    or g200 ( n64 , n193 , n291 );
    or g201 ( n4 , n35 , n198 );
    buf g202 ( n56 , n74 );
    or g203 ( n264 , n12 , n244 );
    xnor g204 ( n74 , n122 , n218 );
    xnor g205 ( n168 , n264 , n130 );
    not g206 ( n112 , n71 );
    xnor g207 ( n189 , n288 , n108 );
    xnor g208 ( n102 , n14 , n136 );
    xnor g209 ( n8 , n245 , n52 );
    xor g210 ( n71 , n1 , n182 );
    or g211 ( n300 , n155 , n82 );
    xnor g212 ( n242 , n6 , n254 );
    not g213 ( n79 , n84 );
    xnor g214 ( n123 , n215 , n211 );
    xnor g215 ( n151 , n302 , n234 );
    or g216 ( n127 , n150 , n175 );
    or g217 ( n266 , n56 , n273 );
    not g218 ( n50 , n233 );
    xnor g219 ( n295 , n23 , n43 );
    or g220 ( n22 , n247 , n103 );
    or g221 ( n16 , n270 , n109 );
    xnor g222 ( n42 , n272 , n196 );
    or g223 ( n116 , n20 , n109 );
    or g224 ( n147 , n165 , n255 );
    or g225 ( n181 , n183 , n148 );
    or g226 ( n170 , n241 , n231 );
    or g227 ( n165 , n205 , n155 );
    xnor g228 ( n225 , n111 , n248 );
    not g229 ( n241 , n71 );
    xnor g230 ( n265 , n4 , n194 );
    or g231 ( n35 , n301 , n138 );
    not g232 ( n157 , n37 );
    not g233 ( n192 , n292 );
    or g234 ( n285 , n79 , n103 );
    not g235 ( n184 , n18 );
    or g236 ( n55 , n162 , n259 );
    xnor g237 ( n309 , n186 , n54 );
    xor g238 ( n119 , n125 , n118 );
    or g239 ( n97 , n192 , n103 );
    or g240 ( n13 , n279 , n72 );
    or g241 ( n106 , n273 , n93 );
    not g242 ( n273 , n227 );
    or g243 ( n307 , n241 , n190 );
    not g244 ( n231 , n100 );
    not g245 ( n51 , n180 );
    or g246 ( n76 , n282 , n300 );
    or g247 ( n224 , n228 , n275 );
    not g248 ( n247 , n133 );
    xnor g249 ( n83 , n146 , n262 );
    or g250 ( n201 , n139 , n92 );
    or g251 ( n228 , n140 , n82 );
    xnor g252 ( n182 , n203 , n121 );
    xnor g253 ( n124 , n107 , n289 );
    or g254 ( n15 , n162 , n51 );
    or g255 ( n219 , n48 , n166 );
    xnor g256 ( n253 , n31 , n272 );
    not g257 ( n180 , n119 );
    not g258 ( n138 , n177 );
    xnor g259 ( n108 , n308 , n40 );
    not g260 ( n110 , n78 );
    or g261 ( n271 , n170 , n275 );
    or g262 ( n20 , n140 , n175 );
    xnor g263 ( n98 , n154 , n27 );
    xnor g264 ( n44 , n22 , n117 );
    xnor g265 ( n111 , n0 , n211 );
    or g266 ( n282 , n205 , n231 );
    xnor g267 ( n288 , n311 , n295 );
    xnor g268 ( n40 , n237 , n90 );
    xnor g269 ( n261 , n176 , n0 );
    or g270 ( n144 , n110 , n216 );
endmodule
