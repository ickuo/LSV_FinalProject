// Benchmark "top" written by ABC on Sun Dec 21 18:12:26 2025

module top ( 
    n0, n21, n36, n38, n45, n49, n77, n95, n98, n104, n107, n108, n116,
    n122, n127, n128, n138, n153, n192, n196, n200, n208, n221, n231, n236,
    n244, n245, n246, n252, n258, n260, n262, n267, n268, n281, n284, n288,
    n301, n305, n310, n319, n323, n324, n332, n336, n359, n360, n364, n366,
    n381, n384, n393, n398, n421, n423, n431, n433, n438, n439, n441, n444,
    n448, n449, n475, n491, n500, n505, n507, n510, n519, n532, n536, n540,
    n571, n577, n589, n599, n610, n631, n635, n640, n644, n650, n657, n667,
    n685, n688, n695, n714, n716, n741, n745, n749, n766, n767, n771, n774,
    n787, n802, n804, n806, n818, n819, n823, n825, n826, n833, n839, n841,
    n845, n851, n857, n862, n863, n866, n870, n879, n893, n896, n901, n928,
    n929, n936, n944, n952, n955, n961, n975, n976, n986, n997, n1005,
    n1022, n1029, n1035, n1036, n1041, n1044, n1045, n1048, n1064, n1067,
    n1069, n1072, n1073, n1077, n1080, n1081, n1089, n1091, n1097, n1098,
    n1120, n1131, n1132, n1140, n1141, n1143, n1146, n1151, n1163, n1164,
    n1180, n1191, n1198, n1219, n1226, n1229, n1231, n1236, n1257, n1269,
    n1273, n1277, n1279, n1298, n1308, n1311, n1321, n1326, n1342, n1344,
    n1352,
    n29, n34, n60, n81, n82, n88, n90, n91, n112, n129, n130, n135, n150,
    n159, n167, n168, n175, n185, n190, n193, n204, n206, n207, n218, n223,
    n227, n228, n229, n240, n275, n299, n307, n342, n347, n374, n383, n389,
    n408, n409, n410, n415, n432, n452, n456, n492, n516, n554, n580, n592,
    n598, n607, n608, n613, n617, n621, n623, n627, n638, n651, n653, n662,
    n679, n683, n707, n710, n718, n723, n733, n734, n747, n779, n785, n801,
    n807, n808, n817, n835, n842, n853, n854, n877, n905, n908, n927, n962,
    n966, n973, n999, n1023, n1027, n1057, n1059, n1061, n1085, n1099,
    n1150, n1153, n1178, n1184, n1194, n1202, n1206, n1232, n1239, n1259,
    n1264, n1288, n1301  );
  input  n0, n21, n36, n38, n45, n49, n77, n95, n98, n104, n107, n108,
    n116, n122, n127, n128, n138, n153, n192, n196, n200, n208, n221, n231,
    n236, n244, n245, n246, n252, n258, n260, n262, n267, n268, n281, n284,
    n288, n301, n305, n310, n319, n323, n324, n332, n336, n359, n360, n364,
    n366, n381, n384, n393, n398, n421, n423, n431, n433, n438, n439, n441,
    n444, n448, n449, n475, n491, n500, n505, n507, n510, n519, n532, n536,
    n540, n571, n577, n589, n599, n610, n631, n635, n640, n644, n650, n657,
    n667, n685, n688, n695, n714, n716, n741, n745, n749, n766, n767, n771,
    n774, n787, n802, n804, n806, n818, n819, n823, n825, n826, n833, n839,
    n841, n845, n851, n857, n862, n863, n866, n870, n879, n893, n896, n901,
    n928, n929, n936, n944, n952, n955, n961, n975, n976, n986, n997,
    n1005, n1022, n1029, n1035, n1036, n1041, n1044, n1045, n1048, n1064,
    n1067, n1069, n1072, n1073, n1077, n1080, n1081, n1089, n1091, n1097,
    n1098, n1120, n1131, n1132, n1140, n1141, n1143, n1146, n1151, n1163,
    n1164, n1180, n1191, n1198, n1219, n1226, n1229, n1231, n1236, n1257,
    n1269, n1273, n1277, n1279, n1298, n1308, n1311, n1321, n1326, n1342,
    n1344, n1352;
  output n29, n34, n60, n81, n82, n88, n90, n91, n112, n129, n130, n135, n150,
    n159, n167, n168, n175, n185, n190, n193, n204, n206, n207, n218, n223,
    n227, n228, n229, n240, n275, n299, n307, n342, n347, n374, n383, n389,
    n408, n409, n410, n415, n432, n452, n456, n492, n516, n554, n580, n592,
    n598, n607, n608, n613, n617, n621, n623, n627, n638, n651, n653, n662,
    n679, n683, n707, n710, n718, n723, n733, n734, n747, n779, n785, n801,
    n807, n808, n817, n835, n842, n853, n854, n877, n905, n908, n927, n962,
    n966, n973, n999, n1023, n1027, n1057, n1059, n1061, n1085, n1099,
    n1150, n1153, n1178, n1184, n1194, n1202, n1206, n1232, n1239, n1259,
    n1264, n1288, n1301;
  wire new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299_1, new_n300, new_n301_1, new_n302, new_n303, new_n304,
    new_n305_1, new_n306, new_n307_1, new_n308, new_n309, new_n310_1,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319_1, new_n320, new_n321, new_n322, new_n323_1,
    new_n324_1, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n331, new_n332_1, new_n333, new_n334, new_n335, new_n336_1,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342_1, new_n343,
    new_n344, new_n345, new_n346, new_n347_1, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359_1, new_n360_1, new_n361, new_n362, new_n363,
    new_n364_1, new_n365, new_n366_1, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374_1, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381_1, new_n382,
    new_n383_1, new_n384_1, new_n385, new_n386, new_n387, new_n388,
    new_n389_1, new_n390, new_n391, new_n392, new_n393_1, new_n394,
    new_n395, new_n396, new_n397, new_n398_1, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408_1,
    new_n409_1, new_n410_1, new_n411, new_n412, new_n413, new_n414,
    new_n415_1, new_n416, new_n417, new_n418, new_n419, new_n420,
    new_n421_1, new_n422, new_n423_1, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n430, new_n431_1, new_n432_1,
    new_n433_1, new_n434, new_n435, new_n436, new_n437, new_n438_1,
    new_n439_1, new_n440, new_n441_1, new_n442, new_n443, new_n444_1,
    new_n445, new_n446, new_n447, new_n448_1, new_n449_1, new_n450,
    new_n451, new_n452_1, new_n453, new_n454, new_n455, new_n456_1,
    new_n457, new_n458, new_n459, new_n460, new_n461, new_n462, new_n463,
    new_n464, new_n465, new_n466, new_n467, new_n468, new_n469, new_n470,
    new_n471, new_n472, new_n473, new_n474, new_n475_1, new_n476, new_n477,
    new_n478, new_n479, new_n480, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491_1,
    new_n492_1, new_n493, new_n494, new_n495, new_n496, new_n497, new_n498,
    new_n499, new_n500_1, new_n501, new_n502, new_n503, new_n504,
    new_n505_1, new_n506, new_n507_1, new_n508, new_n509, new_n510_1,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516_1, new_n517,
    new_n518, new_n519_1, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532_1, new_n533, new_n534, new_n535, new_n536_1, new_n537,
    new_n538, new_n539, new_n540_1, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554_1, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571_1, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577_1, new_n578, new_n579,
    new_n580_1, new_n581, new_n582, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589_1, new_n590, new_n591, new_n592_1, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598_1, new_n599_1,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607_1, new_n608_1, new_n609, new_n610_1, new_n611, new_n612,
    new_n613_1, new_n614, new_n615, new_n616, new_n617_1, new_n618,
    new_n619, new_n620, new_n621_1, new_n622, new_n623_1, new_n624,
    new_n625, new_n626, new_n627_1, new_n628, new_n629, new_n630,
    new_n631_1, new_n632, new_n633, new_n634, new_n635_1, new_n636,
    new_n637, new_n638_1, new_n639, new_n640_1, new_n641, new_n642,
    new_n643, new_n644_1, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650_1, new_n651_1, new_n652, new_n653_1, new_n654, new_n655,
    new_n656, new_n657_1, new_n658, new_n659, new_n660, new_n661,
    new_n662_1, new_n663, new_n664, new_n665, new_n666, new_n667_1,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679_1, new_n680, new_n681,
    new_n682, new_n683_1, new_n684, new_n685_1, new_n686, new_n687,
    new_n688_1, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695_1, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707_1, new_n708,
    new_n709, new_n710_1, new_n711, new_n712, new_n713, new_n714_1,
    new_n715, new_n716_1, new_n717, new_n718_1, new_n719, new_n720,
    new_n721, new_n722, new_n723_1, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734_1, new_n735,
    new_n738, new_n739, new_n740, new_n741_1, new_n742, new_n743, new_n744,
    new_n745_1, new_n746, new_n747_1, new_n748, new_n749_1, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766_1,
    new_n767_1, new_n768, new_n769, new_n770, new_n771_1, new_n772,
    new_n774_1, new_n775, new_n776, new_n778, new_n779_1, new_n781,
    new_n782, new_n783, new_n784, new_n785_1, new_n786, new_n787_1,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801_1,
    new_n802_1, new_n803, new_n804_1, new_n805, new_n806_1, new_n807_1,
    new_n808_1, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817_1, new_n818_1, new_n819_1, new_n820,
    new_n821, new_n822, new_n823_1, new_n824, new_n825_1, new_n826_1,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833_1,
    new_n834, new_n835_1, new_n836, new_n837, new_n838, new_n839_1,
    new_n840, new_n841_1, new_n842_1, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n851_1, new_n852, new_n853_1,
    new_n854_1, new_n855, new_n856, new_n857_1, new_n858, new_n859,
    new_n860, new_n861, new_n862_1, new_n863_1, new_n864, new_n866_1,
    new_n868, new_n871, new_n873, new_n874, new_n875, new_n876, new_n877_1,
    new_n878, new_n879_1, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893_1, new_n894, new_n895, new_n896_1, new_n897,
    new_n898, new_n899, new_n900, new_n901_1, new_n902, new_n903, new_n904,
    new_n905_1, new_n906, new_n907, new_n908_1, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927_1, new_n928_1, new_n929_1, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936_1, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944_1,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952_1, new_n953, new_n954, new_n955_1, new_n956, new_n957,
    new_n959, new_n960, new_n962_1, new_n963, new_n964, new_n965,
    new_n966_1, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973_1, new_n974, new_n975_1, new_n976_1, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986_1, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997_1, new_n998,
    new_n999_1, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005_1, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022_1,
    new_n1023_1, new_n1024, new_n1025, new_n1026, new_n1027_1, new_n1028,
    new_n1029_1, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035_1, new_n1036_1, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041_1, new_n1042, new_n1043, new_n1044_1, new_n1045_1, new_n1046,
    new_n1047, new_n1048_1, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057_1, new_n1058,
    new_n1059_1, new_n1060, new_n1061_1, new_n1062, new_n1063, new_n1064_1,
    new_n1065, new_n1067_1, new_n1068, new_n1069_1, new_n1070, new_n1071,
    new_n1072_1, new_n1073_1, new_n1074, new_n1075, new_n1076, new_n1077_1,
    new_n1078, new_n1079, new_n1080_1, new_n1081_1, new_n1082, new_n1083,
    new_n1084, new_n1085_1, new_n1086, new_n1087, new_n1091_1, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097_1, new_n1099_1, new_n1101,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120_1,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131_1, new_n1132_1,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140_1, new_n1141_1, new_n1142, new_n1143_1, new_n1144,
    new_n1145, new_n1146_1, new_n1147, new_n1148, new_n1149, new_n1150_1,
    new_n1151_1, new_n1152, new_n1153_1, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163_1, new_n1164_1, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178_1, new_n1179, new_n1180_1,
    new_n1181, new_n1182, new_n1183, new_n1184_1, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191_1, new_n1192,
    new_n1193, new_n1194_1, new_n1195, new_n1196, new_n1197, new_n1198_1,
    new_n1200, new_n1201, new_n1202_1, new_n1203, new_n1206_1, new_n1208,
    new_n1210, new_n1211, new_n1212, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219_1, new_n1221, new_n1222, new_n1224, new_n1225,
    new_n1226_1, new_n1227, new_n1228, new_n1229_1, new_n1230, new_n1231_1,
    new_n1232_1, new_n1233, new_n1234, new_n1235, new_n1236_1, new_n1237,
    new_n1238, new_n1239_1, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257_1, new_n1258, new_n1259_1, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264_1, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269_1, new_n1270, new_n1271, new_n1272, new_n1273_1,
    new_n1274, new_n1275, new_n1276, new_n1277_1, new_n1278, new_n1279_1,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288_1, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298_1, new_n1299, new_n1300, new_n1301_1, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308_1, new_n1309,
    new_n1310, new_n1311_1, new_n1312, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1320, new_n1321_1,
    new_n1322, new_n1323, new_n1324, new_n1325, new_n1326_1, new_n1327,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1339, new_n1341, new_n1342_1, new_n1343,
    new_n1345, new_n1346, new_n1347, new_n1349, new_n1350, new_n1351,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1363, new_n1365, new_n1367, new_n1369,
    new_n1370, new_n1371, new_n1372, new_n1373, new_n1374, new_n1375,
    new_n1376, new_n1377, new_n1378, new_n1379, new_n1380, new_n1381,
    new_n1382, new_n1383, new_n1384, new_n1385, new_n1386, new_n1387,
    new_n1388, new_n1389, new_n1390, new_n1391, new_n1392, new_n1393,
    new_n1394, new_n1395, new_n1396, new_n1397, new_n1398, new_n1399,
    new_n1400, new_n1401, new_n1402, new_n1403, new_n1404, new_n1405,
    new_n1406, new_n1407, new_n1408, new_n1409, new_n1410, new_n1411,
    new_n1412, new_n1413, new_n1414, new_n1415, new_n1416, new_n1417,
    new_n1418, new_n1419, new_n1420, new_n1421, new_n1422, new_n1423,
    new_n1424, new_n1425, new_n1426, new_n1427, new_n1428, new_n1429,
    new_n1430, new_n1431, new_n1432, new_n1433, new_n1434, new_n1435,
    new_n1436, new_n1437, new_n1438, new_n1439, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1444, new_n1445, new_n1447, new_n1448,
    new_n1449, new_n1451, new_n1453, new_n1454, new_n1455, new_n1456,
    new_n1458, new_n1459, new_n1460;
  assign new_n293 = ~n839 & ~n1022;
  assign new_n294 = n975 & new_n293;
  assign new_n295 = n1352 & ~new_n294;
  assign new_n296 = ~n688 & ~n1229;
  assign new_n297 = n688 & ~n1098;
  assign new_n298 = ~new_n296 & ~new_n297;
  assign new_n299_1 = n208 & ~n688;
  assign new_n300 = ~n107 & n688;
  assign new_n301_1 = ~new_n299_1 & ~new_n300;
  assign new_n302 = new_n298 & ~new_n301_1;
  assign new_n303 = n688 & n823;
  assign new_n304 = n631 & ~n688;
  assign new_n305_1 = ~new_n303 & ~new_n304;
  assign new_n306 = n77 & ~n688;
  assign new_n307_1 = ~n589 & n688;
  assign new_n308 = ~new_n306 & ~new_n307_1;
  assign new_n309 = ~new_n305_1 & ~new_n308;
  assign new_n310_1 = ~new_n302 & ~new_n309;
  assign new_n311 = new_n305_1 & new_n308;
  assign new_n312 = ~new_n310_1 & ~new_n311;
  assign new_n313 = ~new_n298 & new_n301_1;
  assign new_n314 = n657 & n688;
  assign new_n315 = ~n688 & n1132;
  assign new_n316 = ~new_n314 & ~new_n315;
  assign new_n317 = n260 & ~n688;
  assign new_n318 = ~n360 & n688;
  assign new_n319_1 = ~new_n317 & ~new_n318;
  assign new_n320 = new_n316 & new_n319_1;
  assign new_n321 = n366 & n688;
  assign new_n322 = ~n688 & n879;
  assign new_n323_1 = ~new_n321 & ~new_n322;
  assign new_n324_1 = ~n688 & n1005;
  assign new_n325 = ~n301 & n688;
  assign new_n326 = ~new_n324_1 & ~new_n325;
  assign new_n327 = ~new_n323_1 & ~new_n326;
  assign new_n328 = ~n688 & n1069;
  assign new_n329 = n650 & n688;
  assign new_n330 = ~new_n328 & ~new_n329;
  assign new_n331 = ~n688 & n1279;
  assign new_n332_1 = n688 & ~n1321;
  assign new_n333 = ~new_n331 & ~new_n332_1;
  assign new_n334 = ~new_n330 & ~new_n333;
  assign new_n335 = ~new_n327 & ~new_n334;
  assign new_n336_1 = new_n323_1 & new_n326;
  assign new_n337 = n688 & n1097;
  assign new_n338 = n200 & ~n688;
  assign new_n339 = ~new_n337 & ~new_n338;
  assign new_n340 = ~n688 & n1131;
  assign new_n341 = ~n571 & n688;
  assign new_n342_1 = ~new_n340 & ~new_n341;
  assign new_n343 = ~new_n339 & ~new_n342_1;
  assign new_n344 = n323 & ~n688;
  assign new_n345 = n98 & n688;
  assign new_n346 = ~new_n344 & ~new_n345;
  assign new_n347_1 = n262 & ~n688;
  assign new_n348 = n688 & ~n1198;
  assign new_n349 = ~new_n347_1 & ~new_n348;
  assign new_n350 = ~new_n346 & ~new_n349;
  assign new_n351 = ~new_n343 & ~new_n350;
  assign new_n352 = new_n339 & new_n342_1;
  assign new_n353 = ~new_n351 & ~new_n352;
  assign new_n354 = ~new_n336_1 & new_n353;
  assign new_n355 = new_n335 & ~new_n354;
  assign new_n356 = new_n330 & new_n333;
  assign new_n357 = n688 & n1064;
  assign new_n358 = n536 & ~n688;
  assign new_n359_1 = ~new_n357 & ~new_n358;
  assign new_n360_1 = n441 & ~n688;
  assign new_n361 = ~n104 & n688;
  assign new_n362 = ~new_n360_1 & ~new_n361;
  assign new_n363 = new_n359_1 & new_n362;
  assign new_n364_1 = ~new_n356 & ~new_n363;
  assign new_n365 = ~new_n355 & new_n364_1;
  assign new_n366_1 = ~new_n359_1 & ~new_n362;
  assign new_n367 = ~new_n316 & ~new_n319_1;
  assign new_n368 = ~new_n366_1 & ~new_n367;
  assign new_n369 = ~new_n365 & new_n368;
  assign new_n370 = ~new_n320 & ~new_n369;
  assign new_n371 = n500 & ~n688;
  assign new_n372 = n688 & n1073;
  assign new_n373 = ~new_n371 & ~new_n372;
  assign new_n374_1 = n258 & ~n688;
  assign new_n375 = n688 & ~n1311;
  assign new_n376 = ~new_n374_1 & ~new_n375;
  assign new_n377 = ~new_n373 & ~new_n376;
  assign new_n378 = n688 & n1219;
  assign new_n379 = ~n688 & n1072;
  assign new_n380 = ~new_n378 & ~new_n379;
  assign new_n381_1 = ~n688 & n929;
  assign new_n382 = n688 & ~n1035;
  assign new_n383_1 = ~new_n381_1 & ~new_n382;
  assign new_n384_1 = new_n380 & new_n383_1;
  assign new_n385 = n688 & n714;
  assign new_n386 = ~n688 & n1151;
  assign new_n387 = ~new_n385 & ~new_n386;
  assign new_n388 = ~n688 & n1141;
  assign new_n389_1 = n688 & ~n1081;
  assign new_n390 = ~new_n388 & ~new_n389_1;
  assign new_n391 = new_n387 & new_n390;
  assign new_n392 = n364 & n688;
  assign new_n393_1 = n221 & ~n688;
  assign new_n394 = ~new_n392 & ~new_n393_1;
  assign new_n395 = n510 & ~n688;
  assign new_n396 = ~n45 & n688;
  assign new_n397 = ~new_n395 & ~new_n396;
  assign new_n398_1 = new_n394 & new_n397;
  assign new_n399 = n305 & n688;
  assign new_n400 = ~n688 & n845;
  assign new_n401 = ~new_n399 & ~new_n400;
  assign new_n402 = ~n688 & n1120;
  assign new_n403 = ~n138 & n688;
  assign new_n404 = ~new_n402 & ~new_n403;
  assign new_n405 = ~new_n401 & ~new_n404;
  assign new_n406 = ~new_n387 & ~new_n390;
  assign new_n407 = ~new_n405 & ~new_n406;
  assign new_n408_1 = n688 & n1146;
  assign new_n409_1 = ~n688 & n863;
  assign new_n410_1 = ~new_n408_1 & ~new_n409_1;
  assign new_n411 = ~n688 & n774;
  assign new_n412 = n688 & ~n997;
  assign new_n413 = ~new_n411 & ~new_n412;
  assign new_n414 = ~new_n410_1 & ~new_n413;
  assign new_n415_1 = n688 & n1140;
  assign new_n416 = ~n688 & n893;
  assign new_n417 = ~new_n415_1 & ~new_n416;
  assign new_n418 = ~n688 & n833;
  assign new_n419 = n688 & ~n1308;
  assign new_n420 = ~new_n418 & ~new_n419;
  assign new_n421_1 = new_n417 & new_n420;
  assign new_n422 = n431 & n688;
  assign new_n423_1 = ~n688 & n741;
  assign new_n424 = ~new_n422 & ~new_n423_1;
  assign new_n425 = n540 & ~n688;
  assign new_n426 = ~n36 & n688;
  assign new_n427 = ~new_n425 & ~new_n426;
  assign new_n428 = new_n424 & new_n427;
  assign new_n429 = ~n532 & n685;
  assign new_n430 = ~n688 & ~n857;
  assign new_n431_1 = n685 & ~n688;
  assign new_n432_1 = n532 & ~new_n431_1;
  assign new_n433_1 = ~new_n430 & ~new_n432_1;
  assign new_n434 = ~new_n429 & ~new_n433_1;
  assign new_n435 = ~new_n428 & ~new_n434;
  assign new_n436 = n688 & n1080;
  assign new_n437 = ~n688 & n1077;
  assign new_n438_1 = ~new_n436 & ~new_n437;
  assign new_n439_1 = ~n688 & n1164;
  assign new_n440 = ~n38 & n688;
  assign new_n441_1 = ~new_n439_1 & ~new_n440;
  assign new_n442 = ~new_n438_1 & ~new_n441_1;
  assign new_n443 = ~new_n424 & ~new_n427;
  assign new_n444_1 = ~new_n442 & ~new_n443;
  assign new_n445 = ~new_n435 & new_n444_1;
  assign new_n446 = new_n438_1 & new_n441_1;
  assign new_n447 = ~new_n445 & ~new_n446;
  assign new_n448_1 = ~new_n421_1 & new_n447;
  assign new_n449_1 = ~new_n417 & ~new_n420;
  assign new_n450 = ~new_n448_1 & ~new_n449_1;
  assign new_n451 = ~new_n414 & new_n450;
  assign new_n452_1 = new_n410_1 & new_n413;
  assign new_n453 = new_n401 & new_n404;
  assign new_n454 = ~new_n452_1 & ~new_n453;
  assign new_n455 = ~new_n451 & new_n454;
  assign new_n456_1 = new_n407 & ~new_n455;
  assign new_n457 = ~new_n398_1 & ~new_n456_1;
  assign new_n458 = ~new_n391 & new_n457;
  assign new_n459 = ~new_n380 & ~new_n383_1;
  assign new_n460 = ~new_n394 & ~new_n397;
  assign new_n461 = ~new_n459 & ~new_n460;
  assign new_n462 = ~new_n458 & new_n461;
  assign new_n463 = ~new_n384_1 & ~new_n462;
  assign new_n464 = ~new_n377 & ~new_n463;
  assign new_n465 = new_n373 & new_n376;
  assign new_n466 = ~new_n363 & ~new_n465;
  assign new_n467 = new_n335 & new_n466;
  assign new_n468 = ~new_n320 & ~new_n356;
  assign new_n469 = new_n467 & new_n468;
  assign new_n470 = new_n346 & new_n349;
  assign new_n471 = ~new_n366_1 & ~new_n470;
  assign new_n472 = ~new_n336_1 & ~new_n352;
  assign new_n473 = new_n471 & new_n472;
  assign new_n474 = new_n469 & new_n473;
  assign new_n475_1 = ~new_n464 & new_n474;
  assign new_n476 = new_n351 & new_n475_1;
  assign new_n477 = ~new_n370 & ~new_n476;
  assign new_n478 = new_n310_1 & ~new_n311;
  assign new_n479 = ~new_n477 & new_n478;
  assign new_n480 = ~new_n313 & new_n479;
  assign n456 = new_n312 | new_n480;
  assign new_n482 = n839 & n1022;
  assign new_n483 = n975 & ~new_n482;
  assign new_n484 = ~n1352 & new_n483;
  assign new_n485 = n95 & n866;
  assign new_n486 = n336 & n384;
  assign new_n487 = ~n688 & new_n486;
  assign new_n488 = ~new_n485 & new_n487;
  assign new_n489 = ~new_n484 & ~new_n488;
  assign new_n490 = ~n688 & ~n804;
  assign new_n491_1 = ~n688 & ~new_n486;
  assign new_n492_1 = n936 & ~new_n486;
  assign new_n493 = ~new_n491_1 & ~new_n492_1;
  assign new_n494 = ~new_n490 & ~new_n493;
  assign new_n495 = ~n519 & ~n688;
  assign new_n496 = n284 & ~new_n486;
  assign new_n497 = ~new_n491_1 & ~new_n496;
  assign new_n498 = ~new_n495 & ~new_n497;
  assign new_n499 = ~n667 & ~n688;
  assign new_n500_1 = n688 & ~n928;
  assign new_n501 = ~new_n486 & ~new_n500_1;
  assign new_n502 = ~new_n499 & new_n501;
  assign new_n503 = ~new_n498 & ~new_n502;
  assign new_n504 = ~n281 & n688;
  assign new_n505_1 = ~new_n486 & ~new_n504;
  assign new_n506 = n640 & ~n688;
  assign new_n507_1 = ~n393 & n688;
  assign new_n508 = ~new_n506 & ~new_n507_1;
  assign new_n509 = new_n505_1 & ~new_n508;
  assign new_n510_1 = new_n503 & ~new_n509;
  assign new_n511 = ~new_n494 & new_n510_1;
  assign new_n512 = n688 & n1044;
  assign new_n513 = ~n688 & n695;
  assign new_n514 = ~new_n512 & ~new_n513;
  assign new_n515 = ~n688 & n1326;
  assign new_n516_1 = ~n644 & n688;
  assign new_n517 = ~new_n515 & ~new_n516_1;
  assign new_n518 = ~new_n514 & ~new_n517;
  assign new_n519_1 = ~new_n490 & ~new_n495;
  assign new_n520 = ~new_n499 & new_n519_1;
  assign new_n521 = ~new_n508 & new_n520;
  assign new_n522 = ~new_n505_1 & ~new_n521;
  assign new_n523 = n196 & ~n688;
  assign new_n524 = n688 & n806;
  assign new_n525 = ~new_n523 & ~new_n524;
  assign new_n526 = ~n688 & n1091;
  assign new_n527 = ~n332 & n688;
  assign new_n528 = ~new_n526 & ~new_n527;
  assign new_n529 = ~new_n525 & ~new_n528;
  assign new_n530 = n688 & n745;
  assign new_n531 = ~n688 & n825;
  assign new_n532_1 = ~new_n530 & ~new_n531;
  assign new_n533 = n245 & ~n688;
  assign new_n534 = n688 & ~n716;
  assign new_n535 = ~new_n533 & ~new_n534;
  assign new_n536_1 = ~new_n532_1 & ~new_n535;
  assign new_n537 = ~new_n529 & ~new_n536_1;
  assign new_n538 = n610 & n688;
  assign new_n539 = ~n688 & n841;
  assign new_n540_1 = ~new_n538 & ~new_n539;
  assign new_n541 = n423 & ~n688;
  assign new_n542 = ~n449 & n688;
  assign new_n543 = ~new_n541 & ~new_n542;
  assign new_n544 = new_n540_1 & new_n543;
  assign new_n545 = new_n537 & ~new_n544;
  assign new_n546 = ~new_n522 & new_n545;
  assign new_n547 = ~new_n518 & new_n546;
  assign new_n548 = new_n511 & new_n547;
  assign new_n549 = n688 & ~n771;
  assign new_n550 = ~new_n486 & ~new_n549;
  assign new_n551 = n246 & ~n688;
  assign new_n552 = ~n231 & n688;
  assign new_n553 = ~new_n551 & ~new_n552;
  assign new_n554_1 = new_n550 & ~new_n553;
  assign new_n555 = new_n532_1 & new_n535;
  assign new_n556 = ~new_n554_1 & ~new_n555;
  assign new_n557 = new_n525 & new_n528;
  assign new_n558 = new_n514 & new_n517;
  assign new_n559 = ~new_n550 & new_n553;
  assign new_n560 = ~new_n558 & ~new_n559;
  assign new_n561 = ~new_n557 & new_n560;
  assign new_n562 = new_n556 & new_n561;
  assign new_n563 = new_n548 & new_n562;
  assign new_n564 = new_n489 & new_n563;
  assign new_n565 = n456 & new_n564;
  assign new_n566 = ~new_n295 & ~new_n565;
  assign new_n567 = ~new_n540_1 & ~new_n543;
  assign new_n568 = ~new_n518 & ~new_n567;
  assign new_n569 = ~new_n558 & ~new_n568;
  assign new_n570 = ~new_n555 & new_n569;
  assign new_n571_1 = new_n537 & ~new_n570;
  assign new_n572 = ~new_n557 & ~new_n571_1;
  assign new_n573 = ~new_n554_1 & ~new_n572;
  assign new_n574 = ~new_n522 & ~new_n559;
  assign new_n575 = ~new_n573 & new_n574;
  assign new_n576 = new_n511 & ~new_n575;
  assign new_n577_1 = new_n489 & ~new_n576;
  assign new_n578 = ~n95 & ~n866;
  assign new_n579 = ~n688 & new_n578;
  assign new_n580_1 = ~new_n486 & ~new_n579;
  assign new_n581 = ~new_n484 & new_n580_1;
  assign new_n582 = ~new_n577_1 & ~new_n581;
  assign n29 = ~new_n566 | ~new_n582;
  assign new_n584 = n310 & n688;
  assign new_n585 = ~new_n531 & ~new_n584;
  assign new_n586 = n716 & new_n585;
  assign new_n587 = ~n716 & ~new_n585;
  assign new_n588 = ~new_n586 & ~new_n587;
  assign new_n589_1 = n688 & n1180;
  assign new_n590 = ~new_n304 & ~new_n589_1;
  assign new_n591 = ~n589 & ~new_n590;
  assign new_n592_1 = n589 & new_n590;
  assign new_n593 = ~new_n591 & ~new_n592_1;
  assign new_n594 = ~n421 & n688;
  assign new_n595 = ~new_n296 & ~new_n594;
  assign new_n596 = ~n107 & new_n595;
  assign new_n597 = n107 & ~new_n595;
  assign new_n598_1 = n0 & n688;
  assign new_n599_1 = ~new_n315 & ~new_n598_1;
  assign new_n600 = ~n360 & ~new_n599_1;
  assign new_n601 = n360 & new_n599_1;
  assign new_n602 = n688 & n1273;
  assign new_n603 = ~new_n358 & ~new_n602;
  assign new_n604 = ~n104 & ~new_n603;
  assign new_n605 = ~new_n601 & new_n604;
  assign new_n606 = ~new_n600 & ~new_n605;
  assign new_n607_1 = ~new_n597 & ~new_n606;
  assign new_n608_1 = ~new_n596 & ~new_n607_1;
  assign new_n609 = ~new_n596 & ~new_n597;
  assign new_n610_1 = ~new_n600 & ~new_n601;
  assign new_n611 = n104 & new_n603;
  assign new_n612 = ~new_n604 & ~new_n611;
  assign new_n613_1 = new_n610_1 & new_n612;
  assign new_n614 = new_n609 & new_n613_1;
  assign new_n615 = n688 & n826;
  assign new_n616 = ~new_n328 & ~new_n615;
  assign new_n617_1 = ~n1321 & ~new_n616;
  assign new_n618 = n1321 & new_n616;
  assign new_n619 = ~new_n617_1 & ~new_n618;
  assign new_n620 = n688 & n1045;
  assign new_n621_1 = ~new_n322 & ~new_n620;
  assign new_n622 = n301 & new_n621_1;
  assign new_n623_1 = n688 & n1089;
  assign new_n624 = ~new_n379 & ~new_n623_1;
  assign new_n625 = ~n1035 & ~new_n624;
  assign new_n626 = n1035 & new_n624;
  assign new_n627_1 = ~new_n625 & ~new_n626;
  assign new_n628 = n688 & n1191;
  assign new_n629 = ~new_n393_1 & ~new_n628;
  assign new_n630 = ~n45 & ~new_n629;
  assign new_n631_1 = n45 & new_n629;
  assign new_n632 = n688 & n961;
  assign new_n633 = ~new_n386 & ~new_n632;
  assign new_n634 = n1081 & new_n633;
  assign new_n635_1 = ~n1081 & ~new_n633;
  assign new_n636 = n122 & n688;
  assign new_n637 = ~new_n400 & ~new_n636;
  assign new_n638_1 = ~n138 & ~new_n637;
  assign new_n639 = ~new_n635_1 & ~new_n638_1;
  assign new_n640_1 = ~new_n634 & ~new_n639;
  assign new_n641 = ~new_n631_1 & new_n640_1;
  assign new_n642 = ~new_n630 & ~new_n641;
  assign new_n643 = ~new_n630 & ~new_n631_1;
  assign new_n644_1 = n138 & new_n637;
  assign new_n645 = ~new_n634 & ~new_n644_1;
  assign new_n646 = new_n639 & new_n645;
  assign new_n647 = new_n643 & new_n646;
  assign new_n648 = ~new_n409_1 & ~new_n636;
  assign new_n649 = ~n997 & ~new_n648;
  assign new_n650_1 = n997 & new_n648;
  assign new_n651_1 = ~new_n649 & ~new_n650_1;
  assign new_n652 = ~new_n416 & ~new_n636;
  assign new_n653_1 = ~n1308 & ~new_n652;
  assign new_n654 = n1308 & new_n652;
  assign new_n655 = ~new_n653_1 & ~new_n654;
  assign new_n656 = n108 & n688;
  assign new_n657_1 = ~new_n437 & ~new_n656;
  assign new_n658 = ~n38 & ~new_n657_1;
  assign new_n659 = n38 & new_n657_1;
  assign new_n660 = ~new_n658 & ~new_n659;
  assign new_n661 = n444 & n688;
  assign new_n662_1 = ~new_n423_1 & ~new_n661;
  assign new_n663 = ~n36 & ~new_n662_1;
  assign new_n664 = n36 & new_n662_1;
  assign new_n665 = ~new_n663 & ~new_n664;
  assign new_n666 = new_n660 & new_n665;
  assign new_n667_1 = ~n268 & new_n431_1;
  assign new_n668 = ~new_n664 & new_n667_1;
  assign new_n669 = ~new_n663 & ~new_n668;
  assign new_n670 = ~new_n659 & ~new_n669;
  assign new_n671 = ~new_n658 & ~new_n670;
  assign new_n672 = ~new_n666 & new_n671;
  assign new_n673 = ~n685 & ~n688;
  assign new_n674 = n268 & new_n673;
  assign new_n675 = ~new_n667_1 & ~new_n674;
  assign new_n676 = ~n944 & new_n675;
  assign new_n677 = new_n671 & ~new_n676;
  assign new_n678 = ~new_n672 & ~new_n677;
  assign new_n679_1 = new_n655 & new_n678;
  assign new_n680 = ~new_n653_1 & ~new_n679_1;
  assign new_n681 = new_n651_1 & ~new_n680;
  assign new_n682 = ~new_n649 & ~new_n681;
  assign new_n683_1 = new_n647 & ~new_n682;
  assign new_n684 = new_n642 & ~new_n683_1;
  assign new_n685_1 = new_n627_1 & ~new_n684;
  assign new_n686 = ~new_n625 & ~new_n685_1;
  assign new_n687 = n688 & n1036;
  assign new_n688_1 = ~new_n338 & ~new_n687;
  assign new_n689 = ~n571 & ~new_n688_1;
  assign new_n690 = n571 & new_n688_1;
  assign new_n691 = ~new_n689 & ~new_n690;
  assign new_n692 = n236 & n688;
  assign new_n693 = ~new_n344 & ~new_n692;
  assign new_n694 = ~n1198 & ~new_n693;
  assign new_n695_1 = n1198 & new_n693;
  assign new_n696 = ~new_n694 & ~new_n695_1;
  assign new_n697 = new_n691 & new_n696;
  assign new_n698 = n688 & n901;
  assign new_n699 = ~new_n371 & ~new_n698;
  assign new_n700 = ~n1311 & ~new_n699;
  assign new_n701 = n1311 & new_n699;
  assign new_n702 = ~new_n700 & ~new_n701;
  assign new_n703 = new_n697 & new_n702;
  assign new_n704 = ~new_n686 & new_n703;
  assign new_n705 = ~n301 & ~new_n621_1;
  assign new_n706 = ~new_n695_1 & new_n700;
  assign new_n707_1 = ~new_n694 & ~new_n706;
  assign new_n708 = ~new_n690 & ~new_n707_1;
  assign new_n709 = ~new_n689 & ~new_n708;
  assign new_n710_1 = ~new_n705 & new_n709;
  assign new_n711 = ~new_n704 & new_n710_1;
  assign new_n712 = ~new_n622 & ~new_n711;
  assign new_n713 = new_n619 & new_n712;
  assign new_n714_1 = ~new_n617_1 & ~new_n713;
  assign new_n715 = new_n614 & ~new_n714_1;
  assign new_n716_1 = new_n608_1 & ~new_n715;
  assign new_n717 = new_n593 & ~new_n716_1;
  assign new_n718_1 = ~new_n591 & ~new_n717;
  assign new_n719 = ~new_n513 & ~new_n584;
  assign new_n720 = ~n644 & ~new_n719;
  assign new_n721 = n644 & new_n719;
  assign new_n722 = ~new_n539 & ~new_n584;
  assign new_n723_1 = ~n449 & ~new_n722;
  assign new_n724 = ~new_n721 & new_n723_1;
  assign new_n725 = ~new_n720 & ~new_n724;
  assign new_n726 = new_n718_1 & new_n725;
  assign new_n727 = n449 & new_n722;
  assign new_n728 = ~new_n721 & ~new_n727;
  assign new_n729 = ~new_n720 & ~new_n728;
  assign new_n730 = ~new_n726 & ~new_n729;
  assign new_n731 = ~new_n588 & new_n730;
  assign new_n732 = new_n588 & ~new_n730;
  assign n81 = new_n731 | new_n732;
  assign new_n734_1 = new_n612 & new_n714_1;
  assign new_n735 = ~new_n612 & ~new_n714_1;
  assign n90 = new_n734_1 | new_n735;
  assign n112 = n116 & n1257;
  assign new_n738 = ~new_n523 & ~new_n584;
  assign new_n739 = n332 & new_n738;
  assign new_n740 = ~n332 & ~new_n738;
  assign new_n741_1 = ~new_n739 & ~new_n740;
  assign new_n742 = ~new_n586 & ~new_n725;
  assign new_n743 = ~new_n587 & ~new_n742;
  assign new_n744 = new_n741_1 & ~new_n743;
  assign new_n745_1 = ~new_n741_1 & new_n743;
  assign new_n746 = ~new_n744 & ~new_n745_1;
  assign new_n747_1 = ~new_n723_1 & ~new_n727;
  assign new_n748 = ~new_n718_1 & new_n747_1;
  assign new_n749_1 = ~new_n720 & ~new_n721;
  assign new_n750 = new_n588 & new_n749_1;
  assign new_n751 = new_n748 & new_n750;
  assign new_n752 = ~new_n746 & ~new_n751;
  assign new_n753 = new_n741_1 & new_n751;
  assign n129 = ~new_n752 & ~new_n753;
  assign new_n755 = new_n686 & new_n702;
  assign new_n756 = ~new_n686 & ~new_n702;
  assign n135 = new_n755 | new_n756;
  assign new_n758 = n599 & ~new_n486;
  assign new_n759 = ~new_n491_1 & ~new_n758;
  assign new_n760 = ~n310 & n688;
  assign new_n761 = ~new_n486 & ~new_n760;
  assign new_n762 = ~n231 & new_n761;
  assign new_n763 = ~new_n740 & ~new_n744;
  assign new_n764 = ~new_n753 & new_n763;
  assign new_n765 = n231 & ~new_n761;
  assign new_n766_1 = ~new_n762 & ~new_n765;
  assign new_n767_1 = ~new_n764 & new_n766_1;
  assign new_n768 = ~new_n762 & ~new_n767_1;
  assign new_n769 = ~n393 & ~new_n768;
  assign new_n770 = ~new_n761 & ~new_n769;
  assign new_n771_1 = ~new_n759 & ~new_n770;
  assign new_n772 = ~new_n758 & new_n770;
  assign n150 = new_n771_1 | new_n772;
  assign new_n774_1 = ~new_n723_1 & ~new_n748;
  assign new_n775 = ~new_n749_1 & new_n774_1;
  assign new_n776 = new_n749_1 & ~new_n774_1;
  assign n167 = ~new_n775 & ~new_n776;
  assign new_n778 = n802 & n1344;
  assign new_n779_1 = n288 & n359;
  assign n168 = new_n778 & new_n779_1;
  assign new_n781 = n393 & new_n768;
  assign new_n782 = ~new_n758 & new_n781;
  assign new_n783 = ~new_n761 & ~new_n782;
  assign new_n784 = new_n758 & ~new_n781;
  assign new_n785_1 = new_n783 & ~new_n784;
  assign new_n786 = ~new_n769 & ~new_n785_1;
  assign new_n787_1 = n1298 & ~new_n486;
  assign new_n788 = ~new_n491_1 & ~new_n787_1;
  assign new_n789 = new_n758 & new_n788;
  assign new_n790 = new_n759 & new_n787_1;
  assign new_n791 = ~new_n789 & ~new_n790;
  assign new_n792 = new_n747_1 & new_n750;
  assign new_n793 = new_n741_1 & new_n792;
  assign new_n794 = ~new_n747_1 & ~new_n763;
  assign new_n795 = new_n747_1 & new_n763;
  assign new_n796 = ~new_n794 & ~new_n795;
  assign new_n797 = ~new_n793 & ~new_n796;
  assign new_n798 = ~new_n588 & ~new_n766_1;
  assign new_n799 = new_n588 & new_n766_1;
  assign new_n800 = ~new_n798 & ~new_n799;
  assign new_n801_1 = new_n741_1 & new_n749_1;
  assign new_n802_1 = ~new_n741_1 & ~new_n749_1;
  assign new_n803 = ~new_n801_1 & ~new_n802_1;
  assign new_n804_1 = new_n729 & ~new_n803;
  assign new_n805 = ~new_n729 & new_n803;
  assign new_n806_1 = ~new_n804_1 & ~new_n805;
  assign new_n807_1 = ~new_n800 & ~new_n806_1;
  assign new_n808_1 = new_n800 & new_n806_1;
  assign new_n809 = ~new_n807_1 & ~new_n808_1;
  assign new_n810 = ~new_n727 & ~new_n743;
  assign new_n811 = new_n727 & new_n743;
  assign new_n812 = ~new_n810 & ~new_n811;
  assign new_n813 = ~new_n792 & new_n812;
  assign new_n814 = ~new_n809 & new_n813;
  assign new_n815 = new_n809 & ~new_n813;
  assign new_n816 = ~new_n814 & ~new_n815;
  assign new_n817_1 = new_n797 & new_n816;
  assign new_n818_1 = ~new_n797 & ~new_n816;
  assign new_n819_1 = ~new_n817_1 & ~new_n818_1;
  assign new_n820 = ~new_n718_1 & ~new_n819_1;
  assign new_n821 = new_n723_1 & new_n746;
  assign new_n822 = ~new_n723_1 & ~new_n746;
  assign new_n823_1 = ~new_n821 & ~new_n822;
  assign new_n824 = ~new_n588 & ~new_n749_1;
  assign new_n825_1 = ~new_n750 & ~new_n824;
  assign new_n826_1 = new_n725 & ~new_n766_1;
  assign new_n827 = ~new_n725 & new_n766_1;
  assign new_n828 = ~new_n826_1 & ~new_n827;
  assign new_n829 = ~new_n825_1 & new_n828;
  assign new_n830 = new_n825_1 & ~new_n828;
  assign new_n831 = ~new_n829 & ~new_n830;
  assign new_n832 = new_n823_1 & ~new_n831;
  assign new_n833_1 = ~new_n823_1 & new_n831;
  assign new_n834 = ~new_n832 & ~new_n833_1;
  assign new_n835_1 = ~new_n796 & new_n834;
  assign new_n836 = new_n796 & ~new_n834;
  assign new_n837 = ~new_n835_1 & ~new_n836;
  assign new_n838 = new_n718_1 & ~new_n837;
  assign new_n839_1 = ~new_n820 & ~new_n838;
  assign new_n840 = ~new_n791 & new_n839_1;
  assign new_n841_1 = new_n791 & ~new_n839_1;
  assign new_n842_1 = ~new_n840 & ~new_n841_1;
  assign new_n843 = new_n786 & new_n842_1;
  assign new_n844 = ~new_n786 & ~new_n842_1;
  assign n190 = ~new_n843 & ~new_n844;
  assign new_n846 = ~n393 & ~new_n761;
  assign new_n847 = ~new_n768 & ~new_n846;
  assign new_n848 = n393 & new_n761;
  assign new_n849 = ~new_n767_1 & ~new_n848;
  assign n204 = new_n847 | new_n849;
  assign new_n851_1 = n749 & ~new_n486;
  assign new_n852 = ~new_n491_1 & ~new_n851_1;
  assign new_n853_1 = n896 & ~new_n486;
  assign new_n854_1 = n986 & ~new_n486;
  assign new_n855 = new_n772 & new_n788;
  assign new_n856 = n505 & ~new_n486;
  assign new_n857_1 = new_n855 & ~new_n856;
  assign new_n858 = ~n398 & n688;
  assign new_n859 = ~new_n486 & ~new_n858;
  assign new_n860 = new_n857_1 & ~new_n859;
  assign new_n861 = ~new_n854_1 & new_n860;
  assign new_n862_1 = ~new_n853_1 & new_n861;
  assign new_n863_1 = ~new_n852 & ~new_n862_1;
  assign new_n864 = new_n852 & new_n862_1;
  assign n206 = new_n863_1 | new_n864;
  assign new_n866_1 = ~new_n857_1 & new_n859;
  assign n218 = new_n860 | new_n866_1;
  assign new_n868 = n944 & ~new_n675;
  assign n228 = ~new_n676 & ~new_n868;
  assign n299 = n1352 | new_n864;
  assign new_n871 = n1352 & new_n864;
  assign n229 = n299 & ~new_n871;
  assign new_n873 = ~new_n667_1 & ~new_n671;
  assign new_n874 = new_n667_1 & new_n671;
  assign new_n875 = ~new_n873 & ~new_n874;
  assign new_n876 = new_n651_1 & new_n655;
  assign new_n877_1 = ~new_n651_1 & ~new_n655;
  assign new_n878 = ~new_n876 & ~new_n877_1;
  assign new_n879_1 = new_n669 & ~new_n878;
  assign new_n880 = ~new_n669 & new_n878;
  assign new_n881 = ~new_n879_1 & ~new_n880;
  assign new_n882 = ~new_n875 & ~new_n881;
  assign new_n883 = new_n875 & new_n881;
  assign new_n884 = ~new_n882 & ~new_n883;
  assign new_n885 = ~new_n665 & ~new_n675;
  assign new_n886 = new_n665 & new_n675;
  assign new_n887 = ~new_n885 & ~new_n886;
  assign new_n888 = new_n660 & ~new_n887;
  assign new_n889 = ~new_n660 & new_n887;
  assign new_n890 = ~new_n888 & ~new_n889;
  assign new_n891 = ~new_n654 & ~new_n671;
  assign new_n892 = ~new_n653_1 & ~new_n891;
  assign new_n893_1 = ~new_n890 & ~new_n892;
  assign new_n894 = new_n890 & new_n892;
  assign new_n895 = ~new_n893_1 & ~new_n894;
  assign new_n896_1 = ~new_n884 & new_n895;
  assign new_n897 = new_n884 & ~new_n895;
  assign new_n898 = n944 & ~new_n897;
  assign new_n899 = ~new_n896_1 & new_n898;
  assign new_n900 = new_n675 & ~new_n892;
  assign new_n901_1 = new_n655 & new_n666;
  assign new_n902 = new_n675 & ~new_n901_1;
  assign new_n903 = new_n892 & ~new_n902;
  assign new_n904 = ~new_n900 & ~new_n903;
  assign new_n905_1 = new_n672 & new_n675;
  assign new_n906 = ~new_n675 & ~new_n875;
  assign new_n907 = ~new_n905_1 & ~new_n906;
  assign new_n908_1 = new_n904 & ~new_n907;
  assign new_n909 = ~new_n904 & new_n907;
  assign new_n910 = ~new_n908_1 & ~new_n909;
  assign new_n911 = new_n669 & ~new_n886;
  assign new_n912 = new_n655 & new_n665;
  assign new_n913 = ~new_n655 & ~new_n665;
  assign new_n914 = ~new_n912 & ~new_n913;
  assign new_n915 = new_n911 & ~new_n914;
  assign new_n916 = ~new_n911 & new_n914;
  assign new_n917 = ~new_n915 & ~new_n916;
  assign new_n918 = new_n651_1 & new_n660;
  assign new_n919 = ~new_n651_1 & ~new_n660;
  assign new_n920 = ~new_n918 & ~new_n919;
  assign new_n921 = new_n917 & ~new_n920;
  assign new_n922 = ~new_n917 & new_n920;
  assign new_n923 = ~new_n921 & ~new_n922;
  assign new_n924 = ~new_n910 & ~new_n923;
  assign new_n925 = new_n910 & new_n923;
  assign new_n926 = ~new_n924 & ~new_n925;
  assign new_n927_1 = ~n944 & new_n926;
  assign new_n928_1 = ~new_n899 & ~new_n927_1;
  assign new_n929_1 = ~new_n634 & ~new_n635_1;
  assign new_n930 = ~new_n638_1 & ~new_n644_1;
  assign new_n931 = ~new_n929_1 & ~new_n930;
  assign new_n932 = ~new_n646 & ~new_n931;
  assign new_n933 = new_n642 & ~new_n932;
  assign new_n934 = ~new_n642 & new_n932;
  assign new_n935 = ~new_n933 & ~new_n934;
  assign new_n936_1 = ~new_n647 & ~new_n935;
  assign new_n937 = ~new_n635_1 & new_n644_1;
  assign new_n938 = ~new_n645 & ~new_n937;
  assign new_n939 = new_n936_1 & new_n938;
  assign new_n940 = ~new_n936_1 & ~new_n938;
  assign new_n941 = ~new_n939 & ~new_n940;
  assign new_n942 = ~new_n682 & new_n941;
  assign new_n943 = ~new_n634 & new_n638_1;
  assign new_n944_1 = ~new_n639 & ~new_n943;
  assign new_n945 = new_n935 & new_n944_1;
  assign new_n946 = ~new_n935 & ~new_n944_1;
  assign new_n947 = ~new_n945 & ~new_n946;
  assign new_n948 = new_n682 & new_n947;
  assign new_n949 = ~new_n942 & ~new_n948;
  assign new_n950 = new_n627_1 & new_n643;
  assign new_n951 = ~new_n627_1 & ~new_n643;
  assign new_n952_1 = ~new_n950 & ~new_n951;
  assign new_n953 = new_n949 & ~new_n952_1;
  assign new_n954 = ~new_n949 & new_n952_1;
  assign new_n955_1 = ~new_n953 & ~new_n954;
  assign new_n956 = ~new_n928_1 & ~new_n955_1;
  assign new_n957 = new_n928_1 & new_n955_1;
  assign n240 = new_n956 | new_n957;
  assign new_n959 = ~new_n491_1 & ~new_n854_1;
  assign new_n960 = ~new_n860 & ~new_n959;
  assign n389 = new_n861 | new_n960;
  assign new_n962_1 = ~n688 & ~new_n293;
  assign new_n963 = ~new_n482 & new_n962_1;
  assign new_n964 = ~n475 & n688;
  assign new_n965 = n866 & n1231;
  assign new_n966_1 = ~n866 & ~n1231;
  assign new_n967 = ~new_n965 & ~new_n966_1;
  assign new_n968 = ~n688 & ~new_n967;
  assign new_n969 = ~new_n964 & ~new_n968;
  assign new_n970 = ~new_n963 & new_n969;
  assign new_n971 = new_n963 & ~new_n969;
  assign new_n972 = ~new_n970 & ~new_n971;
  assign new_n973_1 = ~new_n499 & new_n535;
  assign new_n974 = n245 & new_n499;
  assign new_n975_1 = ~new_n973_1 & ~new_n974;
  assign new_n976_1 = n688 & n819;
  assign new_n977 = ~n688 & ~n818;
  assign new_n978 = ~new_n976_1 & ~new_n977;
  assign new_n979 = new_n975_1 & new_n978;
  assign new_n980 = ~new_n975_1 & ~new_n978;
  assign new_n981 = ~new_n979 & ~new_n980;
  assign new_n982 = ~n519 & ~n804;
  assign new_n983 = ~new_n519_1 & ~new_n982;
  assign new_n984 = ~new_n517 & new_n983;
  assign new_n985 = new_n517 & ~new_n983;
  assign new_n986_1 = ~new_n984 & ~new_n985;
  assign new_n987 = ~new_n528 & new_n543;
  assign new_n988 = new_n528 & ~new_n543;
  assign new_n989 = ~new_n987 & ~new_n988;
  assign new_n990 = new_n508 & new_n553;
  assign new_n991 = ~new_n508 & ~new_n553;
  assign new_n992 = ~new_n990 & ~new_n991;
  assign new_n993 = new_n989 & ~new_n992;
  assign new_n994 = ~new_n989 & new_n992;
  assign new_n995 = ~new_n993 & ~new_n994;
  assign new_n996 = ~new_n986_1 & new_n995;
  assign new_n997_1 = new_n986_1 & ~new_n995;
  assign new_n998 = ~new_n996 & ~new_n997_1;
  assign new_n999_1 = new_n981 & ~new_n998;
  assign new_n1000 = ~new_n981 & new_n998;
  assign new_n1001 = ~new_n999_1 & ~new_n1000;
  assign new_n1002 = ~new_n972 & ~new_n1001;
  assign new_n1003 = n267 & ~n688;
  assign new_n1004 = n688 & ~n1342;
  assign new_n1005_1 = ~new_n1003 & ~new_n1004;
  assign new_n1006 = ~new_n349 & new_n1005_1;
  assign new_n1007 = new_n349 & ~new_n1005_1;
  assign new_n1008 = ~new_n1006 & ~new_n1007;
  assign new_n1009 = ~new_n342_1 & new_n376;
  assign new_n1010 = new_n342_1 & ~new_n376;
  assign new_n1011 = ~new_n1009 & ~new_n1010;
  assign new_n1012 = new_n326 & new_n333;
  assign new_n1013 = ~new_n326 & ~new_n333;
  assign new_n1014 = ~new_n1012 & ~new_n1013;
  assign new_n1015 = new_n1011 & new_n1014;
  assign new_n1016 = ~new_n1011 & ~new_n1014;
  assign new_n1017 = ~new_n1015 & ~new_n1016;
  assign new_n1018 = ~new_n319_1 & new_n362;
  assign new_n1019 = new_n319_1 & ~new_n362;
  assign new_n1020 = ~new_n1018 & ~new_n1019;
  assign new_n1021 = new_n301_1 & new_n308;
  assign new_n1022_1 = ~new_n301_1 & ~new_n308;
  assign new_n1023_1 = ~new_n1021 & ~new_n1022_1;
  assign new_n1024 = new_n1020 & new_n1023_1;
  assign new_n1025 = ~new_n1020 & ~new_n1023_1;
  assign new_n1026 = ~new_n1024 & ~new_n1025;
  assign new_n1027_1 = new_n1017 & new_n1026;
  assign new_n1028 = ~new_n1017 & ~new_n1026;
  assign new_n1029_1 = ~new_n1027_1 & ~new_n1028;
  assign new_n1030 = ~new_n1008 & new_n1029_1;
  assign new_n1031 = new_n1008 & ~new_n1029_1;
  assign new_n1032 = ~new_n1030 & ~new_n1031;
  assign new_n1033 = ~new_n390 & new_n404;
  assign new_n1034 = new_n390 & ~new_n404;
  assign new_n1035_1 = ~new_n1033 & ~new_n1034;
  assign new_n1036_1 = new_n383_1 & new_n397;
  assign new_n1037 = ~new_n383_1 & ~new_n397;
  assign new_n1038 = ~new_n1036_1 & ~new_n1037;
  assign new_n1039 = new_n1035_1 & new_n1038;
  assign new_n1040 = ~new_n1035_1 & ~new_n1038;
  assign new_n1041_1 = ~new_n1039 & ~new_n1040;
  assign new_n1042 = new_n413 & new_n1041_1;
  assign new_n1043 = ~new_n413 & ~new_n1041_1;
  assign new_n1044_1 = ~new_n1042 & ~new_n1043;
  assign new_n1045_1 = n381 & n688;
  assign new_n1046 = ~n688 & ~n1269;
  assign new_n1047 = ~new_n1045_1 & ~new_n1046;
  assign new_n1048_1 = n268 & n688;
  assign new_n1049 = ~new_n430 & ~new_n1048_1;
  assign new_n1050 = new_n441_1 & new_n1049;
  assign new_n1051 = ~new_n441_1 & ~new_n1049;
  assign new_n1052 = ~new_n1050 & ~new_n1051;
  assign new_n1053 = new_n420 & new_n427;
  assign new_n1054 = ~new_n420 & ~new_n427;
  assign new_n1055 = ~new_n1053 & ~new_n1054;
  assign new_n1056 = new_n1052 & ~new_n1055;
  assign new_n1057_1 = ~new_n1052 & new_n1055;
  assign new_n1058 = ~new_n1056 & ~new_n1057_1;
  assign new_n1059_1 = new_n1047 & new_n1058;
  assign new_n1060 = ~new_n1047 & ~new_n1058;
  assign new_n1061_1 = ~new_n1059_1 & ~new_n1060;
  assign new_n1062 = new_n1044_1 & ~new_n1061_1;
  assign new_n1063 = ~new_n1044_1 & new_n1061_1;
  assign new_n1064_1 = ~new_n1062 & ~new_n1063;
  assign new_n1065 = new_n1032 & ~new_n1064_1;
  assign n408 = new_n1002 & new_n1065;
  assign new_n1067_1 = new_n852 & new_n853_1;
  assign new_n1068 = ~new_n491_1 & ~new_n853_1;
  assign new_n1069_1 = new_n851_1 & new_n1068;
  assign new_n1070 = ~new_n1067_1 & ~new_n1069_1;
  assign new_n1071 = ~new_n491_1 & ~new_n856;
  assign new_n1072_1 = ~n398 & new_n854_1;
  assign new_n1073_1 = new_n1071 & ~new_n1072_1;
  assign new_n1074 = new_n855 & ~new_n1073_1;
  assign new_n1075 = new_n854_1 & ~new_n859;
  assign new_n1076 = new_n859 & new_n959;
  assign new_n1077_1 = ~new_n1075 & ~new_n1076;
  assign new_n1078 = ~new_n1071 & ~new_n1077_1;
  assign new_n1079 = new_n1071 & new_n1077_1;
  assign new_n1080_1 = ~new_n1078 & ~new_n1079;
  assign new_n1081_1 = ~new_n1074 & new_n1080_1;
  assign new_n1082 = new_n1074 & ~new_n1080_1;
  assign new_n1083 = ~new_n1081_1 & ~new_n1082;
  assign new_n1084 = ~new_n862_1 & new_n1083;
  assign new_n1085_1 = new_n1070 & new_n1084;
  assign new_n1086 = ~new_n1070 & ~new_n1084;
  assign new_n1087 = ~new_n1085_1 & ~new_n1086;
  assign n409 = ~new_n871 & new_n1087;
  assign n432 = n127 | n976;
  assign n592 = n127 | ~n1041;
  assign new_n1091_1 = n491 & n787;
  assign n598 = n127 | ~new_n1091_1;
  assign new_n1093 = new_n606 & ~new_n613_1;
  assign new_n1094 = new_n606 & new_n714_1;
  assign new_n1095 = ~new_n1093 & ~new_n1094;
  assign new_n1096 = ~new_n609 & new_n1095;
  assign new_n1097_1 = new_n609 & ~new_n1095;
  assign n607 = new_n1096 | new_n1097_1;
  assign new_n1099_1 = ~new_n655 & ~new_n678;
  assign n621 = ~new_n679_1 & ~new_n1099_1;
  assign new_n1101 = new_n718_1 & ~new_n747_1;
  assign n627 = ~new_n748 & ~new_n1101;
  assign new_n1103 = n439 & n507;
  assign new_n1104 = ~n439 & ~n507;
  assign new_n1105 = n688 & ~new_n1104;
  assign new_n1106 = ~new_n1103 & new_n1105;
  assign new_n1107 = ~new_n486 & ~new_n1106;
  assign new_n1108 = ~new_n1070 & new_n1107;
  assign new_n1109 = new_n1070 & ~new_n1107;
  assign new_n1110 = ~new_n1108 & ~new_n1109;
  assign new_n1111 = new_n1080_1 & ~new_n1110;
  assign new_n1112 = ~new_n1080_1 & new_n1110;
  assign new_n1113 = ~new_n1111 & ~new_n1112;
  assign new_n1114 = n688 & n1163;
  assign new_n1115 = ~n688 & n1143;
  assign new_n1116 = ~new_n1114 & ~new_n1115;
  assign new_n1117 = new_n719 & ~new_n1116;
  assign new_n1118 = ~new_n719 & new_n1116;
  assign new_n1119 = ~new_n1117 & ~new_n1118;
  assign new_n1120_1 = new_n523 & new_n722;
  assign new_n1121 = ~new_n722 & new_n738;
  assign new_n1122 = ~new_n1120_1 & ~new_n1121;
  assign new_n1123 = ~new_n1119 & new_n1122;
  assign new_n1124 = new_n1119 & ~new_n1122;
  assign new_n1125 = ~new_n1123 & ~new_n1124;
  assign new_n1126 = new_n585 & new_n1125;
  assign new_n1127 = ~new_n585 & ~new_n1125;
  assign new_n1128 = ~new_n1126 & ~new_n1127;
  assign new_n1129 = new_n761 & ~new_n791;
  assign new_n1130 = ~new_n761 & new_n791;
  assign new_n1131_1 = ~new_n1129 & ~new_n1130;
  assign new_n1132_1 = new_n1128 & ~new_n1131_1;
  assign new_n1133 = ~new_n1128 & new_n1131_1;
  assign new_n1134 = ~new_n1132_1 & ~new_n1133;
  assign new_n1135 = ~n252 & n688;
  assign new_n1136 = ~new_n673 & ~new_n1135;
  assign new_n1137 = ~new_n409_1 & ~new_n416;
  assign new_n1138 = n863 & new_n416;
  assign new_n1139 = ~new_n1137 & ~new_n1138;
  assign new_n1140_1 = ~new_n1136 & new_n1139;
  assign new_n1141_1 = new_n1136 & ~new_n1139;
  assign new_n1142 = ~new_n1140_1 & ~new_n1141_1;
  assign new_n1143_1 = new_n662_1 & ~new_n1142;
  assign new_n1144 = ~new_n662_1 & new_n1142;
  assign new_n1145 = ~new_n1143_1 & ~new_n1144;
  assign new_n1146_1 = new_n624 & new_n629;
  assign new_n1147 = ~new_n624 & ~new_n629;
  assign new_n1148 = ~new_n1146_1 & ~new_n1147;
  assign new_n1149 = ~n153 & ~n688;
  assign new_n1150_1 = ~n128 & n688;
  assign new_n1151_1 = ~new_n1149 & ~new_n1150_1;
  assign new_n1152 = ~new_n657_1 & new_n1151_1;
  assign new_n1153_1 = new_n657_1 & ~new_n1151_1;
  assign new_n1154 = ~new_n1152 & ~new_n1153_1;
  assign new_n1155 = new_n633 & new_n637;
  assign new_n1156 = ~new_n633 & ~new_n637;
  assign new_n1157 = ~new_n1155 & ~new_n1156;
  assign new_n1158 = new_n1154 & ~new_n1157;
  assign new_n1159 = ~new_n1154 & new_n1157;
  assign new_n1160 = ~new_n1158 & ~new_n1159;
  assign new_n1161 = ~new_n1148 & new_n1160;
  assign new_n1162 = new_n1148 & ~new_n1160;
  assign new_n1163_1 = ~new_n1161 & ~new_n1162;
  assign new_n1164_1 = ~new_n1145 & new_n1163_1;
  assign new_n1165 = new_n1145 & ~new_n1163_1;
  assign new_n1166 = ~new_n1164_1 & ~new_n1165;
  assign new_n1167 = ~new_n1134 & new_n1166;
  assign new_n1168 = new_n599_1 & ~new_n603;
  assign new_n1169 = ~new_n599_1 & new_n603;
  assign new_n1170 = ~new_n1168 & ~new_n1169;
  assign new_n1171 = new_n590 & new_n595;
  assign new_n1172 = ~new_n590 & ~new_n595;
  assign new_n1173 = ~new_n1171 & ~new_n1172;
  assign new_n1174 = new_n1170 & ~new_n1173;
  assign new_n1175 = ~new_n1170 & new_n1173;
  assign new_n1176 = ~new_n1174 & ~new_n1175;
  assign new_n1177 = new_n621_1 & new_n688_1;
  assign new_n1178_1 = ~new_n621_1 & ~new_n688_1;
  assign new_n1179 = ~new_n1177 & ~new_n1178_1;
  assign new_n1180_1 = n688 & n767;
  assign new_n1181 = n192 & ~n688;
  assign new_n1182 = ~new_n1180_1 & ~new_n1181;
  assign new_n1183 = ~new_n699 & new_n1182;
  assign new_n1184_1 = new_n699 & ~new_n1182;
  assign new_n1185 = ~new_n1183 & ~new_n1184_1;
  assign new_n1186 = new_n1179 & new_n1185;
  assign new_n1187 = ~new_n1179 & ~new_n1185;
  assign new_n1188 = ~new_n1186 & ~new_n1187;
  assign new_n1189 = new_n616 & new_n693;
  assign new_n1190 = ~new_n616 & ~new_n693;
  assign new_n1191_1 = ~new_n1189 & ~new_n1190;
  assign new_n1192 = new_n1188 & ~new_n1191_1;
  assign new_n1193 = ~new_n1188 & new_n1191_1;
  assign new_n1194_1 = ~new_n1192 & ~new_n1193;
  assign new_n1195 = ~new_n1176 & new_n1194_1;
  assign new_n1196 = new_n1176 & ~new_n1194_1;
  assign new_n1197 = ~new_n1195 & ~new_n1196;
  assign new_n1198_1 = new_n1167 & new_n1197;
  assign n653 = new_n1113 & new_n1198_1;
  assign new_n1200 = new_n646 & ~new_n682;
  assign new_n1201 = ~new_n640_1 & ~new_n1200;
  assign new_n1202_1 = ~new_n643 & new_n1201;
  assign new_n1203 = new_n643 & ~new_n1201;
  assign n662 = ~new_n1202_1 & ~new_n1203;
  assign n679 = n1352 | ~new_n864;
  assign new_n1206_1 = new_n764 & ~new_n766_1;
  assign n707 = ~new_n767_1 & ~new_n1206_1;
  assign new_n1208 = ~new_n627_1 & new_n684;
  assign n723 = ~new_n685_1 & ~new_n1208;
  assign new_n1210 = ~new_n846 & ~new_n848;
  assign new_n1211 = new_n768 & ~new_n1210;
  assign new_n1212 = ~new_n768 & new_n1210;
  assign n733 = new_n1211 | new_n1212;
  assign new_n1214 = ~new_n611 & ~new_n714_1;
  assign new_n1215 = ~new_n604 & ~new_n1214;
  assign new_n1216 = ~new_n610_1 & new_n1215;
  assign new_n1217 = new_n610_1 & ~new_n1215;
  assign n747 = ~new_n1216 & ~new_n1217;
  assign new_n1219_1 = ~new_n772 & ~new_n788;
  assign n779 = new_n855 | new_n1219_1;
  assign new_n1221 = ~new_n682 & ~new_n930;
  assign new_n1222 = new_n682 & new_n930;
  assign n808 = new_n1221 | new_n1222;
  assign new_n1224 = ~new_n316 & new_n359_1;
  assign new_n1225 = new_n316 & ~new_n359_1;
  assign new_n1226_1 = ~new_n1224 & ~new_n1225;
  assign new_n1227 = new_n298 & new_n305_1;
  assign new_n1228 = ~new_n298 & ~new_n305_1;
  assign new_n1229_1 = ~new_n1227 & ~new_n1228;
  assign new_n1230 = new_n1226_1 & new_n1229_1;
  assign new_n1231_1 = ~new_n1226_1 & ~new_n1229_1;
  assign new_n1232_1 = ~new_n1230 & ~new_n1231_1;
  assign new_n1233 = new_n346 & new_n1232_1;
  assign new_n1234 = ~new_n346 & ~new_n1232_1;
  assign new_n1235 = ~new_n1233 & ~new_n1234;
  assign new_n1236_1 = n688 & ~n1067;
  assign new_n1237 = ~new_n1181 & ~new_n1236_1;
  assign new_n1238 = ~new_n339 & new_n1237;
  assign new_n1239_1 = new_n339 & ~new_n1237;
  assign new_n1240 = ~new_n1238 & ~new_n1239_1;
  assign new_n1241 = new_n323_1 & new_n330;
  assign new_n1242 = ~new_n323_1 & ~new_n330;
  assign new_n1243 = ~new_n1241 & ~new_n1242;
  assign new_n1244 = new_n373 & ~new_n1243;
  assign new_n1245 = ~new_n373 & new_n1243;
  assign new_n1246 = ~new_n1244 & ~new_n1245;
  assign new_n1247 = ~new_n1240 & ~new_n1246;
  assign new_n1248 = new_n1240 & new_n1246;
  assign new_n1249 = ~new_n1247 & ~new_n1248;
  assign new_n1250 = ~new_n1235 & ~new_n1249;
  assign new_n1251 = new_n438_1 & ~new_n673;
  assign new_n1252 = n1077 & new_n673;
  assign new_n1253 = ~new_n1251 & ~new_n1252;
  assign new_n1254 = n893 & new_n1149;
  assign new_n1255 = new_n417 & ~new_n1149;
  assign new_n1256 = ~new_n1254 & ~new_n1255;
  assign new_n1257_1 = ~new_n1253 & new_n1256;
  assign new_n1258 = new_n1253 & ~new_n1256;
  assign new_n1259_1 = ~new_n1257_1 & ~new_n1258;
  assign new_n1260 = ~new_n387 & new_n401;
  assign new_n1261 = new_n387 & ~new_n401;
  assign new_n1262 = ~new_n1260 & ~new_n1261;
  assign new_n1263 = new_n380 & new_n394;
  assign new_n1264_1 = ~new_n380 & ~new_n394;
  assign new_n1265 = ~new_n1263 & ~new_n1264_1;
  assign new_n1266 = new_n1262 & new_n1265;
  assign new_n1267 = ~new_n1262 & ~new_n1265;
  assign new_n1268 = ~new_n1266 & ~new_n1267;
  assign new_n1269_1 = new_n410_1 & new_n424;
  assign new_n1270 = ~new_n410_1 & ~new_n424;
  assign new_n1271 = ~new_n1269_1 & ~new_n1270;
  assign new_n1272 = new_n1268 & ~new_n1271;
  assign new_n1273_1 = ~new_n1268 & new_n1271;
  assign new_n1274 = ~new_n1272 & ~new_n1273_1;
  assign new_n1275 = ~new_n1259_1 & new_n1274;
  assign new_n1276 = new_n1259_1 & ~new_n1274;
  assign new_n1277_1 = ~new_n1275 & ~new_n1276;
  assign new_n1278 = ~new_n1250 & new_n1277_1;
  assign new_n1279_1 = new_n492_1 & new_n497;
  assign new_n1280 = new_n493 & new_n496;
  assign new_n1281 = ~new_n1279_1 & ~new_n1280;
  assign new_n1282 = new_n532_1 & new_n540_1;
  assign new_n1283 = ~new_n532_1 & ~new_n540_1;
  assign new_n1284 = ~new_n1282 & ~new_n1283;
  assign new_n1285 = ~new_n1281 & new_n1284;
  assign new_n1286 = new_n1281 & ~new_n1284;
  assign new_n1287 = ~new_n1285 & ~new_n1286;
  assign new_n1288_1 = ~n433 & n688;
  assign new_n1289 = ~new_n1115 & ~new_n1288_1;
  assign new_n1290 = new_n550 & ~new_n1289;
  assign new_n1291 = ~new_n550 & new_n1289;
  assign new_n1292 = ~new_n1290 & ~new_n1291;
  assign new_n1293 = new_n514 & new_n525;
  assign new_n1294 = ~new_n514 & ~new_n525;
  assign new_n1295 = ~new_n1293 & ~new_n1294;
  assign new_n1296 = new_n1292 & ~new_n1295;
  assign new_n1297 = ~new_n1292 & new_n1295;
  assign new_n1298_1 = ~new_n1296 & ~new_n1297;
  assign new_n1299 = new_n500_1 & new_n505_1;
  assign new_n1300 = new_n501 & ~new_n505_1;
  assign new_n1301_1 = ~new_n1299 & ~new_n1300;
  assign new_n1302 = ~new_n1298_1 & new_n1301_1;
  assign new_n1303 = new_n1298_1 & ~new_n1301_1;
  assign new_n1304 = ~new_n1302 & ~new_n1303;
  assign new_n1305 = ~new_n1287 & ~new_n1304;
  assign new_n1306 = new_n1287 & new_n1304;
  assign new_n1307 = ~new_n1305 & ~new_n1306;
  assign new_n1308_1 = new_n1235 & new_n1249;
  assign new_n1309 = ~n955 & n1048;
  assign new_n1310 = n955 & ~n1048;
  assign new_n1311_1 = ~new_n1309 & ~new_n1310;
  assign new_n1312 = n438 & n851;
  assign new_n1313 = ~n438 & ~n851;
  assign new_n1314 = ~new_n1312 & ~new_n1313;
  assign new_n1315 = new_n1311_1 & new_n1314;
  assign new_n1316 = ~new_n1311_1 & ~new_n1314;
  assign new_n1317 = ~new_n1315 & ~new_n1316;
  assign new_n1318 = n49 & ~n244;
  assign new_n1319 = ~n49 & n244;
  assign new_n1320 = ~new_n1318 & ~new_n1319;
  assign new_n1321_1 = new_n1317 & ~new_n1320;
  assign new_n1322 = ~new_n1317 & new_n1320;
  assign new_n1323 = ~new_n486 & ~new_n1322;
  assign new_n1324 = n688 & new_n1323;
  assign new_n1325 = ~new_n1321_1 & new_n1324;
  assign new_n1326_1 = ~new_n1308_1 & ~new_n1325;
  assign new_n1327 = ~new_n1307 & new_n1326_1;
  assign n817 = new_n1278 & new_n1327;
  assign new_n1329 = new_n686 & new_n707_1;
  assign new_n1330 = ~new_n694 & new_n701;
  assign new_n1331 = ~new_n695_1 & ~new_n1330;
  assign new_n1332 = ~new_n1329 & new_n1331;
  assign new_n1333 = ~new_n691 & new_n1332;
  assign new_n1334 = new_n691 & ~new_n1332;
  assign n835 = new_n1333 | new_n1334;
  assign new_n1336 = n577 & n870;
  assign new_n1337 = n324 & n448;
  assign n854 = new_n1336 & new_n1337;
  assign new_n1339 = ~new_n855 & ~new_n1071;
  assign n905 = new_n857_1 | new_n1339;
  assign new_n1341 = n408 & n817;
  assign new_n1342_1 = n1029 & n1236;
  assign new_n1343 = n319 & n952;
  assign n1027 = new_n1342_1 & new_n1343;
  assign new_n1345 = n854 & n1027;
  assign new_n1346 = n766 & n1226;
  assign new_n1347 = n21 & n635;
  assign n999 = new_n1346 & new_n1347;
  assign new_n1349 = new_n1345 & n999;
  assign new_n1350 = new_n1341 & new_n1349;
  assign new_n1351 = n168 & n653;
  assign n927 = new_n1350 & new_n1351;
  assign new_n1353 = ~new_n638_1 & new_n682;
  assign new_n1354 = ~new_n644_1 & ~new_n1353;
  assign new_n1355 = new_n929_1 & new_n1354;
  assign new_n1356 = ~new_n929_1 & ~new_n1354;
  assign n962 = ~new_n1355 & ~new_n1356;
  assign new_n1358 = ~new_n622 & ~new_n705;
  assign new_n1359 = ~new_n704 & new_n709;
  assign new_n1360 = ~new_n1358 & new_n1359;
  assign new_n1361 = new_n1358 & ~new_n1359;
  assign n1059 = ~new_n1360 & ~new_n1361;
  assign new_n1363 = ~new_n619 & ~new_n712;
  assign n1061 = ~new_n713 & ~new_n1363;
  assign new_n1365 = ~new_n651_1 & new_n680;
  assign n1085 = ~new_n681 & ~new_n1365;
  assign new_n1367 = ~new_n861 & ~new_n1068;
  assign n1099 = new_n862_1 | new_n1367;
  assign new_n1369 = ~new_n610_1 & ~new_n612;
  assign new_n1370 = ~new_n613_1 & ~new_n1369;
  assign new_n1371 = ~new_n608_1 & new_n1370;
  assign new_n1372 = new_n608_1 & ~new_n1370;
  assign new_n1373 = ~new_n1371 & ~new_n1372;
  assign new_n1374 = ~new_n614 & ~new_n1373;
  assign new_n1375 = new_n600 & new_n611;
  assign new_n1376 = new_n601 & ~new_n611;
  assign new_n1377 = ~new_n1375 & ~new_n1376;
  assign new_n1378 = new_n593 & ~new_n609;
  assign new_n1379 = ~new_n593 & new_n609;
  assign new_n1380 = ~new_n1378 & ~new_n1379;
  assign new_n1381 = new_n1377 & ~new_n1380;
  assign new_n1382 = ~new_n1377 & new_n1380;
  assign new_n1383 = ~new_n1381 & ~new_n1382;
  assign new_n1384 = new_n1374 & new_n1383;
  assign new_n1385 = ~new_n1374 & ~new_n1383;
  assign new_n1386 = ~new_n1384 & ~new_n1385;
  assign new_n1387 = ~new_n714_1 & ~new_n1386;
  assign new_n1388 = ~new_n600 & ~new_n604;
  assign new_n1389 = ~new_n605 & ~new_n1388;
  assign new_n1390 = ~new_n1380 & new_n1389;
  assign new_n1391 = new_n1380 & ~new_n1389;
  assign new_n1392 = ~new_n1390 & ~new_n1391;
  assign new_n1393 = new_n1373 & new_n1392;
  assign new_n1394 = ~new_n1373 & ~new_n1392;
  assign new_n1395 = ~new_n1393 & ~new_n1394;
  assign new_n1396 = new_n714_1 & new_n1395;
  assign new_n1397 = ~new_n1387 & ~new_n1396;
  assign new_n1398 = ~new_n622 & ~new_n710_1;
  assign new_n1399 = ~new_n702 & new_n1398;
  assign new_n1400 = new_n702 & ~new_n1398;
  assign new_n1401 = ~new_n1399 & ~new_n1400;
  assign new_n1402 = ~new_n694 & ~new_n700;
  assign new_n1403 = ~new_n706 & ~new_n1402;
  assign new_n1404 = new_n619 & new_n1358;
  assign new_n1405 = ~new_n619 & ~new_n1358;
  assign new_n1406 = ~new_n1404 & ~new_n1405;
  assign new_n1407 = new_n1403 & ~new_n1406;
  assign new_n1408 = ~new_n1403 & new_n1406;
  assign new_n1409 = ~new_n1407 & ~new_n1408;
  assign new_n1410 = ~new_n691 & ~new_n696;
  assign new_n1411 = ~new_n697 & ~new_n1410;
  assign new_n1412 = new_n709 & new_n1411;
  assign new_n1413 = ~new_n709 & ~new_n1411;
  assign new_n1414 = ~new_n1412 & ~new_n1413;
  assign new_n1415 = new_n1409 & ~new_n1414;
  assign new_n1416 = ~new_n1409 & new_n1414;
  assign new_n1417 = ~new_n1415 & ~new_n1416;
  assign new_n1418 = ~new_n1401 & new_n1417;
  assign new_n1419 = new_n1401 & ~new_n1417;
  assign new_n1420 = ~new_n1418 & ~new_n1419;
  assign new_n1421 = new_n686 & ~new_n1420;
  assign new_n1422 = ~new_n701 & ~new_n703;
  assign new_n1423 = new_n709 & new_n1422;
  assign new_n1424 = new_n701 & ~new_n709;
  assign new_n1425 = ~new_n1423 & ~new_n1424;
  assign new_n1426 = new_n1358 & new_n1401;
  assign new_n1427 = ~new_n703 & new_n1358;
  assign new_n1428 = ~new_n1401 & ~new_n1427;
  assign new_n1429 = ~new_n1426 & ~new_n1428;
  assign new_n1430 = ~new_n619 & new_n1331;
  assign new_n1431 = new_n619 & ~new_n1331;
  assign new_n1432 = ~new_n1430 & ~new_n1431;
  assign new_n1433 = ~new_n1411 & new_n1432;
  assign new_n1434 = new_n1411 & ~new_n1432;
  assign new_n1435 = ~new_n1433 & ~new_n1434;
  assign new_n1436 = new_n1429 & new_n1435;
  assign new_n1437 = ~new_n1429 & ~new_n1435;
  assign new_n1438 = ~new_n1436 & ~new_n1437;
  assign new_n1439 = new_n1425 & new_n1438;
  assign new_n1440 = ~new_n1425 & ~new_n1438;
  assign new_n1441 = ~new_n1439 & ~new_n1440;
  assign new_n1442 = ~new_n686 & ~new_n1441;
  assign new_n1443 = ~new_n1421 & ~new_n1442;
  assign new_n1444 = new_n1397 & ~new_n1443;
  assign new_n1445 = ~new_n1397 & new_n1443;
  assign n1150 = new_n1444 | new_n1445;
  assign new_n1447 = ~new_n667_1 & ~new_n676;
  assign new_n1448 = ~new_n665 & new_n1447;
  assign new_n1449 = new_n665 & ~new_n1447;
  assign n1178 = ~new_n1448 & ~new_n1449;
  assign new_n1451 = ~new_n593 & new_n716_1;
  assign n1202 = ~new_n717 & ~new_n1451;
  assign new_n1453 = new_n686 & ~new_n700;
  assign new_n1454 = ~new_n701 & ~new_n1453;
  assign new_n1455 = new_n696 & new_n1454;
  assign new_n1456 = ~new_n696 & ~new_n1454;
  assign n1239 = ~new_n1455 & ~new_n1456;
  assign new_n1458 = ~new_n663 & ~new_n1449;
  assign new_n1459 = ~new_n660 & new_n1458;
  assign new_n1460 = new_n660 & ~new_n1458;
  assign n1301 = ~new_n1459 & ~new_n1460;
  assign n88 = 1'b0;
  assign n159 = 1'b0;
  assign n223 = 1'b0;
  assign n227 = 1'b0;
  assign n374 = 1'b0;
  assign n410 = 1'b0;
  assign n492 = 1'b0;
  assign n608 = 1'b0;
  assign n623 = 1'b0;
  assign n1206 = 1'b0;
  assign n651 = ~n862;
  assign n34 = n116;
  assign n60 = n1081;
  assign n82 = n104;
  assign n91 = n29;
  assign n130 = n716;
  assign n175 = n138;
  assign n185 = n571;
  assign n193 = n644;
  assign n207 = n1198;
  assign n275 = n1277;
  assign n307 = n1308;
  assign n342 = n299;
  assign n347 = n1342;
  assign n383 = n1321;
  assign n415 = n997;
  assign n452 = n393;
  assign n516 = n301;
  assign n554 = n360;
  assign n580 = n449;
  assign n613 = n592;
  assign n617 = n598;
  assign n638 = n1311;
  assign n683 = n381;
  assign n710 = n36;
  assign n718 = n116;
  assign n734 = n475;
  assign n785 = n229;
  assign n801 = n679;
  assign n807 = n45;
  assign n842 = n651;
  assign n853 = n589;
  assign n877 = n679;
  assign n908 = n679;
  assign n966 = n107;
  assign n973 = n819;
  assign n1023 = n38;
  assign n1057 = n332;
  assign n1153 = n231;
  assign n1184 = n651;
  assign n1194 = n116;
  assign n1232 = n268;
  assign n1259 = n29;
  assign n1264 = n116;
  assign n1288 = n1035;
endmodule


