module top( n7 , n18 , n21 , n50 , n55 , n108 , n142 , n175 , n196 , 
n235 , n242 , n243 , n248 , n266 , n268 , n298 , n317 , n329 , n332 , 
n337 , n342 , n357 , n376 , n422 , n431 , n442 , n457 , n463 , n468 , 
n491 , n496 , n498 , n521 , n548 , n554 , n567 , n583 , n588 , n597 , 
n604 , n626 , n637 , n646 , n647 , n655 , n696 , n723 , n735 , n752 , 
n767 , n779 , n809 , n819 , n829 , n849 , n858 , n873 , n879 , n887 , 
n904 , n919 , n932 , n948 , n957 , n980 , n982 , n984 , n987 , n1005 , 
n1016 , n1020 , n1040 , n1044 , n1060 , n1069 , n1099 , n1111 , n1112 , n1118 , 
n1119 , n1120 , n1136 , n1152 , n1163 , n1196 , n1204 , n1222 , n1237 , n1239 , 
n1255 , n1269 , n1279 , n1288 , n1293 , n1302 , n1314 , n1320 , n1332 , n1357 , 
n1371 , n1385 , n1432 , n1437 , n1451 , n1483 , n1498 , n1501 , n1518 , n1525 , 
n1527 , n1536 , n1558 , n1580 , n1586 , n1590 , n1602 , n1611 , n1630 , n1634 , 
n1636 , n1639 , n1654 , n1662 , n1667 , n1681 , n1682 , n1684 , n1689 , n1701 , 
n1703 , n1721 , n1738 , n1742 , n1752 , n1760 , n1777 , n1791 , n1808 , n1821 , 
n1831 , n1832 , n1859 , n1860 , n1861 , n1881 , n1891 , n1925 , n1942 , n1949 , 
n1972 , n1981 , n1999 , n2004 , n2007 , n2013 , n2035 , n2061 , n2088 , n2092 , 
n2095 , n2102 , n2105 , n2113 , n2117 , n2122 , n2145 , n2146 , n2147 , n2160 , 
n2175 , n2184 , n2209 , n2210 , n2214 , n2238 , n2272 , n2289 , n2327 , n2328 , 
n2331 , n2343 , n2355 , n2361 , n2363 , n2374 , n2387 , n2388 , n2409 , n2416 , 
n2420 , n2421 , n2440 , n2444 , n2479 , n2513 , n2515 , n2533 , n2535 , n2537 , 
n2547 , n2553 , n2555 , n2560 , n2561 , n2570 , n2573 , n2578 , n2582 , n2602 , 
n2619 , n2646 , n2659 , n2661 , n2680 , n2693 , n2703 , n2706 , n2711 , n2731 , 
n2743 , n2761 , n2774 , n2779 , n2783 , n2809 , n2816 , n2826 , n2853 , n2858 , 
n2860 , n2886 , n2887 , n2929 , n2944 , n2948 , n2961 , n2971 , n2978 , n2979 , 
n2985 , n2999 , n3010 , n3017 , n3018 , n3020 , n3030 , n3067 , n3076 , n3089 , 
n3125 , n3126 , n3136 , n3161 , n3164 , n3208 , n3219 , n3228 , n3235 , n3244 , 
n3253 , n3260 , n3263 , n3279 , n3289 , n3301 , n3306 , n3316 , n3320 , n3324 , 
n3332 , n3340 , n3343 , n3349 , n3366 , n3390 , n3425 , n3426 , n3451 , n3459 , 
n3460 , n3468 , n3480 , n3502 , n3506 , n3516 , n3528 , n3541 , n3555 , n3561 , 
n3563 , n3570 , n3582 , n3617 , n3618 , n3642 , n3649 , n3665 , n3679 , n3710 , 
n3725 , n3733 , n3740 , n3755 , n3758 , n3760 , n3781 , n3785 , n3794 , n3795 , 
n3828 , n3842 , n3850 , n3869 , n3871 , n3891 , n3909 , n3918 , n3925 , n3932 , 
n3934 , n3945 , n3952 , n3959 , n3962 , n3971 , n3983 , n3984 , n4000 , n4010 , 
n4014 , n4071 , n4085 , n4088 , n4089 , n4100 , n4103 , n4119 , n4123 , n4134 , 
n4146 , n4150 , n4151 , n4152 , n4153 , n4165 , n4172 , n4173 , n4176 , n4186 , 
n4204 , n4205 , n4215 , n4221 , n4224 , n4231 , n4256 , n4266 , n4272 , n4306 , 
n4319 , n4325 , n4326 , n4340 , n4374 , n4376 , n4401 , n4409 , n4424 , n4426 , 
n4432 , n4441 , n4451 , n4476 , n4478 , n4514 , n4529 , n4552 , n4588 , n4590 , 
n4595 , n4624 , n4646 , n4665 , n4674 , n4693 , n4722 , n4731 , n4745 , n4747 , 
n4766 , n4770 , n4777 , n4785 , n4804 , n4810 , n4812 , n4814 , n4850 , n4858 , 
n4891 , n4913 , n4925 , n4939 , n4947 , n4952 , n4957 , n4964 , n4966 , n4967 , 
n4972 , n5011 , n5020 , n5024 , n5025 , n5026 , n5031 , n5046 , n5060 , n5062 , 
n5064 , n5077 , n5082 , n5098 , n5101 , n5115 , n5120 , n5128 , n5131 , n5140 , 
n5158 , n5168 , n5184 , n5211 , n5213 , n5226 , n5228 , n5255 , n5256 , n5265 , 
n5273 , n5274 , n5300 , n5302 , n5325 , n5330 , n5337 , n5351 , n5353 , n5376 , 
n5386 , n5399 , n5400 , n5403 , n5430 , n5438 , n5439 , n5443 , n5451 , n5472 , 
n5485 , n5517 , n5521 , n5524 , n5532 , n5564 , n5579 , n5593 , n5603 , n5605 , 
n5609 , n5634 , n5643 , n5680 , n5687 , n5696 , n5700 , n5704 , n5732 , n5742 , 
n5752 , n5765 , n5776 , n5782 , n5822 , n5833 , n5834 , n5840 , n5841 , n5842 , 
n5850 , n5882 , n5903 , n5904 , n5911 , n5936 , n5943 , n5964 , n5980 , n6012 , 
n6022 , n6031 , n6044 , n6046 , n6084 , n6104 , n6105 , n6160 , n6171 , n6183 , 
n6189 , n6204 , n6218 , n6223 , n6233 , n6245 , n6248 , n6256 , n6271 , n6276 , 
n6308 , n6311 , n6323 , n6330 , n6339 , n6354 , n6356 , n6369 , n6375 , n6379 , 
n6381 , n6383 , n6385 , n6397 , n6407 , n6427 , n6431 , n6437 , n6456 , n6457 , 
n6465 , n6470 , n6476 , n6485 , n6502 , n6506 , n6513 , n6514 , n6542 , n6556 , 
n6558 , n6560 , n6567 , n6576 , n6587 , n6590 , n6596 , n6611 , n6612 , n6628 , 
n6630 , n6631 , n6634 , n6652 , n6655 , n6659 , n6669 , n6671 , n6673 , n6674 , 
n6684 , n6691 , n6706 , n6707 , n6729 , n6736 , n6773 , n6775 , n6785 , n6790 , 
n6791 , n6794 , n6802 , n6814 , n6826 , n6835 , n6853 , n6861 , n6862 , n6863 , 
n6867 , n6965 , n6967 , n6971 , n6975 , n6983 , n6985 , n6998 , n7026 , n7032 , 
n7038 , n7057 , n7079 , n7099 , n7139 , n7149 , n7190 , n7229 , n7230 , n7233 , 
n7236 , n7253 , n7256 , n7268 , n7277 , n7280 , n7298 , n7305 , n7308 , n7313 , 
n7330 , n7335 , n7339 , n7346 , n7349 , n7363 , n7377 , n7390 , n7403 , n7408 , 
n7421 , n7428 , n7432 , n7437 , n7460 , n7475 , n7477 , n7507 , n7514 , n7524 , 
n7558 , n7566 , n7569 , n7572 , n7575 , n7585 , n7588 , n7593 , n7598 , n7607 , 
n7610 , n7616 , n7630 , n7643 , n7647 , n7657 , n7670 , n7674 , n7678 , n7679 , 
n7686 , n7692 , n7693 , n7698 , n7708 , n7721 , n7731 , n7751 , n7759 , n7769 , 
n7773 , n7780 , n7788 , n7794 , n7811 , n7830 , n7834 , n7841 , n7876 , n7884 , 
n7917 , n7937 , n7943 , n7949 , n7950 , n7959 , n7963 , n7968 , n7992 , n7999 , 
n8006 , n8027 , n8031 , n8042 , n8052 , n8067 , n8095 , n8103 , n8109 , n8127 , 
n8130 , n8135 , n8139 , n8148 , n8149 , n8159 , n8179 , n8194 , n8215 , n8244 , 
n8255 , n8256 , n8259 , n8267 , n8276 , n8285 , n8288 , n8305 , n8306 , n8309 , 
n8320 , n8321 , n8324 , n8339 , n8363 , n8376 , n8381 , n8399 , n8405 , n8408 , 
n8417 , n8432 , n8439 , n8453 , n8480 , n8489 , n8505 , n8510 , n8519 , n8526 , 
n8535 , n8550 , n8563 , n8581 , n8594 , n8608 , n8614 , n8620 , n8637 , n8638 , 
n8656 , n8662 , n8678 , n8687 , n8694 , n8716 , n8721 , n8744 , n8745 , n8782 , 
n8803 , n8806 , n8809 , n8821 , n8824 , n8827 , n8849 , n8856 , n8861 , n8862 , 
n8869 , n8884 , n8909 , n8911 , n8920 , n8943 , n8964 , n8971 , n8982 , n8993 , 
n9003 , n9012 , n9032 , n9042 , n9046 , n9047 , n9090 , n9104 , n9129 , n9146 , 
n9164 , n9166 , n9172 , n9182 , n9191 , n9217 , n9220 , n9246 , n9251 , n9259 , 
n9261 , n9287 , n9308 , n9318 , n9323 , n9344 , n9364 , n9371 , n9372 , n9380 , 
n9382 , n9396 , n9399 , n9403 , n9419 , n9423 , n9430 , n9435 , n9445 , n9451 , 
n9458 , n9459 , n9460 , n9493 , n9507 , n9508 , n9512 , n9552 , n9554 , n9556 , 
n9557 , n9558 , n9598 , n9616 , n9622 , n9626 , n9633 , n9635 , n9646 , n9648 , 
n9655 , n9689 , n9695 , n9699 , n9726 , n9753 , n9761 , n9763 , n9767 , n9771 , 
n9778 , n9783 , n9803 , n9832 , n9833 , n9838 , n9867 , n9872 , n9890 , n9917 , 
n9919 , n9926 , n9934 , n9938 , n9942 , n9946 , n9967 , n9968 , n10009 , n10010 , 
n10017 , n10018 , n10019 , n10021 , n10053 , n10055 , n10057 , n10096 , n10101 , n10111 , 
n10117 , n10125 , n10158 , n10165 , n10201 , n10236 , n10239 , n10244 , n10250 , n10261 , 
n10262 , n10275 , n10287 , n10295 , n10321 , n10326 , n10327 , n10330 , n10340 , n10345 , 
n10356 , n10372 , n10385 , n10387 , n10388 , n10390 , n10404 , n10405 , n10409 , n10411 , 
n10420 , n10432 , n10484 , n10489 , n10514 , n10525 , n10540 , n10561 , n10564 , n10577 , 
n10588 , n10593 , n10595 , n10611 , n10614 , n10617 , n10628 , n10647 , n10650 , n10653 , 
n10692 , n10694 , n10701 , n10710 , n10712 , n10739 , n10756 , n10763 , n10775 , n10780 , 
n10792 , n10817 , n10834 , n10851 , n10874 , n10924 , n10943 , n10961 , n11005 , n11011 , 
n11023 , n11025 , n11044 , n11056 , n11063 , n11078 , n11080 , n11094 , n11101 , n11103 , 
n11120 , n11121 , n11127 , n11132 , n11134 , n11138 , n11182 , n11184 , n11192 , n11201 , 
n11220 , n11223 , n11234 , n11245 , n11261 , n11266 , n11273 , n11275 , n11290 , n11302 , 
n11313 , n11325 , n11326 , n11330 , n11347 , n11348 , n11352 , n11356 , n11375 , n11379 , 
n11386 , n11391 , n11398 , n11403 , n11419 , n11424 , n11439 , n11455 , n11462 , n11470 , 
n11472 , n11473 , n11479 , n11481 , n11486 , n11496 , n11503 , n11506 , n11515 , n11538 , 
n11548 , n11564 , n11566 , n11579 , n11580 , n11591 , n11607 , n11615 , n11630 , n11647 , 
n11667 , n11674 , n11682 , n11710 , n11712 , n11724 , n11736 , n11741 , n11749 , n11770 , 
n11771 , n11775 , n11818 , n11837 , n11841 , n11842 , n11843 , n11898 , n11905 , n11926 , 
n11965 , n11980 , n12000 , n12003 , n12011 , n12072 , n12113 , n12121 , n12131 , n12146 , 
n12152 , n12153 , n12157 , n12158 , n12161 , n12179 , n12192 , n12209 , n12223 , n12225 , 
n12228 , n12235 , n12302 , n12304 , n12315 , n12324 , n12325 , n12329 , n12330 , n12341 , 
n12346 , n12349 , n12364 , n12380 , n12383 , n12384 , n12397 , n12398 , n12408 , n12446 , 
n12449 , n12461 , n12462 , n12467 , n12469 , n12495 , n12507 , n12515 , n12516 , n12540 , 
n12545 , n12546 , n12552 , n12562 , n12566 , n12569 , n12587 , n12593 , n12607 , n12620 , 
n12621 , n12626 , n12650 , n12654 , n12657 , n12665 , n12670 , n12702 , n12707 , n12725 , 
n12727 , n12740 , n12742 , n12746 , n12756 , n12783 , n12801 , n12811 , n12812 , n12816 , 
n12821 , n12843 , n12861 , n12864 , n12865 , n12870 , n12871 , n12873 , n12875 , n12892 , 
n12900 , n12904 , n12917 , n12941 , n12942 , n12956 , n12978 , n12980 , n12985 , n12987 , 
n12992 , n13005 , n13026 , n13043 , n13044 , n13048 , n13054 , n13074 , n13082 , n13096 , 
n13110 , n13116 , n13122 , n13137 , n13141 , n13144 , n13168 , n13190 , n13198 , n13199 , 
n13204 , n13209 , n13263 , n13270 , n13273 , n13285 , n13319 , n13333 , n13338 , n13367 , 
n13407 , n13409 , n13419 , n13424 , n13453 , n13456 , n13457 , n13460 , n13477 , n13484 , 
n13486 , n13487 , n13490 , n13494 , n13500 , n13501 , n13506 , n13548 , n13549 , n13551 , 
n13602 , n13626 , n13668 , n13677 , n13683 , n13708 , n13710 , n13714 , n13719 , n13722 , 
n13754 , n13764 , n13775 , n13781 , n13783 , n13798 , n13835 , n13850 , n13851 , n13912 , 
n13914 , n13922 , n13923 , n13951 , n14004 , n14036 , n14059 , n14071 , n14081 , n14090 , 
n14095 , n14107 , n14121 , n14126 , n14130 , n14136 , n14147 , n14148 , n14174 , n14190 , 
n14211 , n14222 , n14230 , n14267 , n14271 , n14275 , n14277 , n14294 , n14310 , n14323 , 
n14326 , n14342 , n14345 , n14353 , n14364 , n14375 , n14412 , n14414 , n14440 , n14457 , 
n14464 , n14471 , n14475 , n14510 , n14541 , n14546 , n14547 , n14570 , n14575 , n14576 , 
n14593 , n14603 , n14633 , n14636 , n14680 , n14684 , n14692 , n14701 , n14702 , n14704 , 
n14734 , n14746 , n14763 , n14772 , n14790 , n14801 , n14819 , n14826 , n14827 , n14839 , 
n14849 , n14891 , n14899 , n14931 , n14944 , n14954 , n14977 , n14989 , n15002 , n15004 , 
n15011 , n15019 , n15031 , n15033 , n15052 , n15053 , n15077 , n15082 , n15094 , n15118 , 
n15128 , n15139 , n15145 , n15146 , n15165 , n15167 , n15176 , n15180 , n15182 , n15205 , 
n15230 , n15241 , n15255 , n15258 , n15271 , n15275 , n15289 , n15300 , n15307 , n15327 , 
n15332 , n15345 , n15353 , n15366 , n15378 , n15382 , n15407 , n15424 , n15428 , n15435 , 
n15438 , n15465 , n15467 , n15470 , n15477 , n15481 , n15490 , n15496 , n15501 , n15506 , 
n15508 , n15539 , n15546 , n15555 , n15558 , n15559 , n15570 , n15573 , n15588 , n15590 , 
n15598 , n15602 , n15614 , n15636 , n15652 , n15662 , n15716 , n15743 , n15749 , n15761 , 
n15762 , n15766 , n15780 , n15793 , n15812 , n15815 , n15816 , n15831 , n15846 , n15859 , 
n15869 , n15884 , n15885 , n15889 , n15917 , n15918 , n15922 , n15936 , n15947 , n15956 , 
n15958 , n15967 , n15979 , n15986 , n16013 , n16029 , n16060 , n16062 , n16068 , n16080 , 
n16098 , n16110 , n16142 , n16158 , n16167 , n16185 , n16196 , n16206 , n16215 , n16217 , 
n16218 , n16219 , n16223 , n16230 , n16243 , n16247 , n16275 , n16279 , n16322 , n16327 , 
n16350 , n16367 , n16376 , n16379 , n16396 , n16398 , n16406 , n16407 , n16419 , n16424 , 
n16428 , n16433 , n16439 , n16440 , n16445 , n16460 , n16476 , n16481 , n16482 , n16493 , 
n16502 , n16506 , n16507 , n16516 , n16517 , n16521 , n16524 , n16527 , n16544 , n16554 , 
n16583 , n16584 , n16589 , n16596 , n16608 , n16617 , n16630 , n16640 , n16656 , n16674 , 
n16682 , n16684 , n16688 , n16722 , n16733 , n16743 , n16798 , n16812 , n16818 , n16824 , 
n16834 , n16837 , n16841 , n16885 , n16905 , n16911 , n16951 , n16954 , n16968 , n16971 , 
n16988 , n16989 , n16994 , n17006 , n17035 , n17037 , n17068 , n17069 , n17070 , n17075 , 
n17077 , n17084 , n17090 , n17095 , n17104 , n17106 , n17119 , n17130 , n17138 , n17163 , 
n17168 , n17202 , n17219 , n17232 , n17236 , n17243 , n17250 , n17251 , n17263 , n17285 , 
n17302 , n17320 , n17337 , n17344 , n17351 , n17359 , n17387 , n17391 , n17392 , n17421 , 
n17432 , n17436 , n17440 , n17450 , n17458 , n17461 , n17466 , n17493 , n17500 , n17524 , 
n17529 , n17557 , n17583 , n17592 , n17638 , n17664 , n17687 , n17721 , n17735 , n17738 , 
n17746 , n17749 , n17784 , n17820 , n17855 , n17877 , n17889 , n17911 , n17912 , n17927 , 
n17931 , n17948 , n17954 , n17956 , n17959 , n17963 , n17968 , n17976 , n17998 , n18025 , 
n18035 , n18043 , n18045 , n18059 , n18061 , n18071 , n18105 , n18143 , n18145 , n18151 , 
n18152 , n18157 , n18171 , n18193 , n18227 , n18232 , n18238 , n18241 , n18254 , n18274 , 
n18288 , n18290 , n18295 , n18301 , n18304 , n18310 , n18311 , n18323 , n18332 , n18343 , 
n18345 , n18350 , n18362 , n18377 , n18405 , n18409 , n18414 , n18418 , n18437 , n18439 , 
n18444 , n18445 , n18452 , n18467 , n18482 , n18483 , n18496 , n18509 , n18513 , n18515 , 
n18537 , n18558 , n18572 , n18574 , n18576 , n18578 , n18582 , n18583 , n18584 , n18610 , 
n18635 , n18649 , n18653 , n18679 , n18690 , n18693 , n18708 , n18721 , n18725 , n18737 , 
n18745 , n18751 , n18780 , n18782 , n18802 , n18830 , n18831 , n18843 , n18858 , n18859 , 
n18864 , n18865 , n18880 , n18886 , n18887 , n18901 , n18907 , n18919 , n18926 , n18940 , 
n18945 , n18962 , n18970 , n18977 , n18982 , n18999 , n19005 , n19033 , n19042 , n19044 , 
n19081 , n19107 , n19116 , n19125 , n19141 , n19144 , n19163 , n19164 , n19174 , n19176 , 
n19196 , n19202 , n19220 , n19221 , n19223 , n19224 , n19228 , n19233 , n19234 , n19244 , 
n19270 , n19282 , n19314 , n19315 , n19323 , n19327 , n19333 , n19348 , n19354 , n19357 , 
n19361 , n19367 , n19385 , n19389 , n19401 , n19414 , n19424 , n19450 , n19454 , n19458 , 
n19467 , n19472 , n19477 , n19494 , n19496 , n19514 , n19515 , n19523 , n19531 , n19539 , 
n19570 , n19575 , n19584 , n19602 , n19608 , n19617 , n19618 , n19623 , n19641 , n19648 , 
n19652 , n19664 , n19680 , n19701 , n19736 , n19749 , n19756 , n19767 , n19770 , n19780 , 
n19789 , n19792 , n19798 , n19803 , n19873 , n19905 , n19909 , n19911 , n19916 , n19922 , 
n19923 , n19930 , n19941 , n19968 , n19988 , n20004 , n20013 , n20017 , n20033 , n20036 , 
n20040 , n20061 , n20069 , n20077 , n20086 , n20096 , n20103 , n20126 , n20138 , n20149 , 
n20151 , n20169 , n20179 , n20187 , n20213 , n20235 , n20250 , n20259 , n20279 , n20287 , 
n20301 , n20330 , n20333 , n20349 , n20355 , n20359 , n20366 , n20385 , n20388 , n20402 , 
n20403 , n20409 , n20411 , n20424 , n20429 , n20436 , n20441 , n20445 , n20450 , n20455 , 
n20470 , n20478 , n20489 , n20490 , n20495 , n20515 , n20533 , n20582 , n20590 , n20602 , 
n20604 , n20609 , n20623 , n20629 , n20658 , n20661 , n20673 , n20678 , n20680 , n20685 , 
n20691 , n20696 , n20700 , n20704 , n20705 , n20709 , n20713 , n20722 , n20723 , n20748 , 
n20761 , n20774 , n20788 , n20794 , n20795 , n20803 , n20826 , n20869 , n20879 , n20915 , 
n20923 , n20929 , n20935 , n20936 , n20946 , n20986 , n21008 , n21017 , n21034 , n21046 , 
n21062 , n21078 , n21093 , n21094 , n21095 , n21123 , n21134 , n21138 , n21154 , n21157 , 
n21168 , n21173 , n21176 , n21182 , n21193 , n21203 , n21222 , n21225 , n21226 , n21238 , 
n21254 , n21276 , n21287 , n21298 , n21302 , n21317 , n21349 , n21365 , n21367 , n21396 , 
n21398 , n21399 , n21404 , n21446 , n21471 , n21472 , n21489 , n21525 , n21538 , n21549 , 
n21599 , n21615 , n21628 , n21637 , n21645 , n21649 , n21654 , n21665 , n21674 , n21680 , 
n21685 , n21687 , n21717 , n21719 , n21735 , n21749 , n21750 , n21753 , n21765 , n21779 , 
n21784 , n21800 , n21820 , n21832 , n21839 , n21874 , n21898 , n21905 , n21915 , n21934 , 
n21943 , n21957 , n21960 , n21976 , n21981 , n21986 , n21993 , n21997 , n22016 , n22027 , 
n22043 , n22050 , n22063 , n22068 , n22072 , n22076 , n22090 , n22107 , n22113 , n22124 , 
n22126 , n22130 , n22144 , n22150 , n22157 , n22173 , n22198 , n22201 , n22213 , n22253 , 
n22270 , n22274 , n22283 , n22290 , n22309 , n22311 , n22317 , n22332 , n22335 , n22341 , 
n22353 , n22358 , n22359 , n22379 , n22433 , n22442 , n22444 , n22467 , n22470 , n22484 , 
n22489 , n22492 , n22494 , n22533 , n22554 , n22584 , n22588 , n22589 , n22591 , n22597 , 
n22619 , n22620 , n22623 , n22626 , n22631 , n22660 , n22697 , n22714 , n22761 , n22764 , 
n22779 , n22787 , n22793 , n22819 , n22843 , n22858 , n22870 , n22871 , n22879 , n22891 , 
n22897 , n22903 , n22907 , n22910 , n22914 , n22918 , n22939 , n22998 , n23006 , n23007 , 
n23009 , n23014 , n23035 , n23039 , n23047 , n23058 , n23065 , n23066 , n23067 , n23068 , 
n23120 , n23146 , n23160 , n23166 , n23200 , n23238 , n23247 , n23248 , n23250 , n23270 , 
n23272 , n23289 , n23304 , n23305 , n23333 , n23341 , n23342 , n23355 , n23369 , n23371 , 
n23401 , n23414 , n23429 , n23430 , n23433 , n23434 , n23450 , n23463 , n23471 , n23480 , 
n23493 , n23513 , n23529 , n23541 , n23546 , n23550 , n23585 , n23586 , n23588 , n23619 , 
n23624 , n23628 , n23637 , n23657 , n23663 , n23669 , n23684 , n23690 , n23697 , n23714 , 
n23717 , n23719 , n23748 , n23755 , n23775 , n23831 , n23842 , n23849 , n23856 , n23883 , 
n23888 , n23895 , n23899 , n23903 , n23912 , n23913 , n23923 , n23924 , n23935 , n23942 , 
n23954 , n23958 , n23974 , n23986 , n24002 , n24004 , n24032 , n24039 , n24048 , n24052 , 
n24085 , n24092 , n24093 , n24096 , n24097 , n24105 , n24119 , n24129 , n24133 , n24141 , 
n24145 , n24146 , n24150 , n24155 , n24160 , n24167 , n24170 , n24172 , n24177 , n24196 , 
n24228 , n24258 , n24260 , n24278 , n24289 , n24297 , n24307 , n24319 , n24323 , n24327 , 
n24342 , n24345 , n24347 , n24373 , n24374 , n24406 , n24415 , n24421 , n24431 , n24472 , 
n24476 , n24483 , n24485 , n24501 , n24512 , n24558 , n24576 , n24579 , n24602 , n24604 , 
n24618 , n24620 , n24626 , n24629 , n24636 , n24638 , n24715 , n24723 , n24732 , n24749 , 
n24758 , n24768 , n24784 , n24786 , n24807 , n24826 , n24840 , n24841 , n24853 , n24857 , 
n24879 , n24887 , n24934 , n24937 , n24998 , n25006 , n25023 , n25032 , n25062 , n25068 , 
n25073 , n25074 , n25083 , n25094 , n25097 , n25119 , n25120 , n25126 , n25133 , n25155 , 
n25168 , n25181 , n25200 , n25209 , n25215 , n25240 , n25244 , n25254 , n25256 , n25293 , 
n25296 , n25316 , n25328 , n25331 , n25332 , n25336 , n25337 , n25345 , n25356 , n25362 , 
n25365 , n25370 , n25381 , n25412 , n25435 , n25460 , n25464 , n25468 , n25471 , n25475 , 
n25494 , n25499 , n25513 , n25518 , n25523 , n25532 , n25539 , n25550 , n25565 , n25586 , 
n25611 , n25614 , n25619 , n25629 , n25643 , n25665 , n25694 , n25706 , n25719 , n25738 , 
n25749 , n25751 , n25756 , n25758 , n25773 , n25784 , n25792 , n25797 , n25816 , n25826 , 
n25839 , n25840 , n25872 , n25873 , n25877 , n25923 , n25926 , n25934 , n25938 , n25972 , 
n25974 , n25985 , n25994 , n26036 , n26053 , n26054 , n26084 , n26096 , n26107 , n26111 , 
n26113 , n26156 , n26159 , n26167 , n26179 , n26180 , n26191 , n26220 , n26224 , n26229 , 
n26237 , n26250 , n26264 , n26274 , n26287 , n26317 , n26318 , n26353 , n26375 , n26396 , 
n26408 , n26429 , n26431 , n26439 , n26443 , n26452 , n26483 , n26492 , n26510 , n26512 , 
n26515 , n26538 , n26553 , n26565 , n26572 , n26590 , n26598 , n26605 , n26625 , n26656 , 
n26660 , n26674 , n26675 , n26681 , n26696 , n26698 , n26707 , n26719 , n26725 , n26727 , 
n26729 , n26744 , n26745 , n26748 , n26752 , n26775 , n26780 , n26794 , n26795 , n26797 , 
n26801 , n26808 , n26815 , n26823 , n26847 , n26882 , n26900 , n26902 , n26905 , n26913 , 
n26921 , n26923 , n26929 , n26930 , n26943 , n26970 , n26979 , n26986 , n27004 , n27011 , 
n27019 , n27031 , n27037 , n27051 , n27072 , n27079 , n27089 , n27096 , n27104 , n27110 , 
n27112 , n27120 , n27130 , n27134 , n27145 , n27158 , n27163 , n27188 , n27194 );
    input n18 , n21 , n196 , n268 , n329 , n337 , n342 , n376 , n442 , 
n468 , n583 , n604 , n626 , n647 , n655 , n752 , n767 , n919 , n932 , 
n987 , n1040 , n1099 , n1112 , n1118 , n1136 , n1152 , n1163 , n1204 , n1222 , 
n1255 , n1269 , n1279 , n1288 , n1293 , n1314 , n1320 , n1432 , n1437 , n1451 , 
n1483 , n1525 , n1536 , n1558 , n1611 , n1630 , n1639 , n1654 , n1662 , n1667 , 
n1681 , n1682 , n1689 , n1738 , n1742 , n1752 , n1777 , n1831 , n1881 , n1949 , 
n1999 , n2013 , n2035 , n2088 , n2102 , n2113 , n2117 , n2145 , n2146 , n2160 , 
n2175 , n2184 , n2210 , n2272 , n2289 , n2328 , n2331 , n2355 , n2387 , n2409 , 
n2416 , n2420 , n2421 , n2479 , n2547 , n2570 , n2646 , n2659 , n2680 , n2731 , 
n2743 , n2783 , n2809 , n2816 , n2858 , n2886 , n2944 , n2978 , n2979 , n2985 , 
n2999 , n3018 , n3030 , n3136 , n3161 , n3164 , n3228 , n3253 , n3260 , n3279 , 
n3306 , n3320 , n3324 , n3349 , n3366 , n3425 , n3460 , n3468 , n3480 , n3506 , 
n3541 , n3570 , n3582 , n3618 , n3710 , n3740 , n3785 , n3795 , n3828 , n3909 , 
n3918 , n3925 , n3945 , n3952 , n3959 , n3962 , n3984 , n4085 , n4100 , n4119 , 
n4256 , n4272 , n4306 , n4319 , n4325 , n4326 , n4376 , n4409 , n4426 , n4514 , 
n4588 , n4590 , n4665 , n4722 , n4812 , n4858 , n4913 , n4939 , n4957 , n4964 , 
n4967 , n5025 , n5026 , n5031 , n5060 , n5077 , n5098 , n5101 , n5115 , n5128 , 
n5131 , n5140 , n5211 , n5213 , n5226 , n5255 , n5302 , n5330 , n5337 , n5376 , 
n5386 , n5400 , n5438 , n5443 , n5451 , n5517 , n5521 , n5532 , n5579 , n5605 , 
n5696 , n5704 , n5752 , n5822 , n5834 , n5842 , n5882 , n6104 , n6105 , n6204 , 
n6218 , n6356 , n6369 , n6379 , n6381 , n6385 , n6397 , n6427 , n6456 , n6485 , 
n6502 , n6513 , n6556 , n6590 , n6596 , n6611 , n6631 , n6659 , n6691 , n6729 , 
n6773 , n6775 , n6785 , n6790 , n6794 , n6814 , n6861 , n6971 , n7026 , n7057 , 
n7099 , n7139 , n7149 , n7305 , n7330 , n7335 , n7339 , n7377 , n7421 , n7428 , 
n7437 , n7460 , n7524 , n7566 , n7569 , n7593 , n7657 , n7670 , n7674 , n7678 , 
n7692 , n7693 , n7721 , n7731 , n7751 , n7759 , n7769 , n7773 , n7788 , n7841 , 
n7876 , n7917 , n7949 , n7963 , n8006 , n8052 , n8067 , n8194 , n8244 , n8255 , 
n8256 , n8259 , n8285 , n8305 , n8309 , n8324 , n8363 , n8381 , n8399 , n8405 , 
n8439 , n8526 , n8581 , n8614 , n8638 , n8656 , n8678 , n8687 , n8694 , n8721 , 
n8745 , n8782 , n8806 , n8827 , n8856 , n8869 , n8920 , n8943 , n8964 , n9003 , 
n9090 , n9172 , n9246 , n9251 , n9259 , n9318 , n9323 , n9372 , n9380 , n9396 , 
n9399 , n9445 , n9460 , n9493 , n9507 , n9512 , n9554 , n9557 , n9598 , n9646 , 
n9655 , n9832 , n9872 , n9926 , n9934 , n9942 , n9967 , n10017 , n10018 , n10053 , 
n10057 , n10096 , n10117 , n10125 , n10158 , n10201 , n10250 , n10275 , n10372 , n10405 , 
n10411 , n10514 , n10577 , n10593 , n10611 , n10614 , n10650 , n10710 , n10712 , n10739 , 
n10763 , n10792 , n11011 , n11044 , n11056 , n11121 , n11184 , n11192 , n11201 , n11220 , 
n11223 , n11266 , n11273 , n11302 , n11356 , n11424 , n11455 , n11473 , n11479 , n11481 , 
n11486 , n11503 , n11566 , n11579 , n11580 , n11615 , n11630 , n11667 , n11736 , n11749 , 
n11775 , n11841 , n11898 , n11926 , n11980 , n12113 , n12121 , n12152 , n12153 , n12161 , 
n12209 , n12315 , n12341 , n12380 , n12384 , n12398 , n12446 , n12495 , n12507 , n12546 , 
n12562 , n12587 , n12593 , n12626 , n12650 , n12657 , n12702 , n12811 , n12821 , n12861 , 
n12871 , n12875 , n12892 , n12900 , n12917 , n12956 , n13026 , n13044 , n13074 , n13110 , 
n13137 , n13190 , n13263 , n13319 , n13333 , n13367 , n13419 , n13424 , n13453 , n13460 , 
n13490 , n13494 , n13549 , n13668 , n13677 , n13708 , n13714 , n13719 , n13775 , n13781 , 
n13783 , n13851 , n13912 , n13914 , n13951 , n14071 , n14090 , n14130 , n14148 , n14230 , 
n14275 , n14323 , n14345 , n14440 , n14510 , n14570 , n14575 , n14576 , n14603 , n14633 , 
n14680 , n14684 , n14692 , n14702 , n14704 , n14790 , n14826 , n14899 , n14954 , n15053 , 
n15077 , n15146 , n15167 , n15182 , n15241 , n15258 , n15271 , n15289 , n15332 , n15378 , 
n15424 , n15490 , n15506 , n15508 , n15539 , n15546 , n15602 , n15636 , n15652 , n15743 , 
n15761 , n15766 , n15780 , n15884 , n15918 , n15936 , n15967 , n15979 , n16029 , n16158 , 
n16167 , n16217 , n16223 , n16247 , n16376 , n16396 , n16439 , n16476 , n16482 , n16502 , 
n16507 , n16521 , n16524 , n16544 , n16608 , n16722 , n16743 , n16812 , n16818 , n16824 , 
n16911 , n16968 , n16971 , n16988 , n16994 , n17035 , n17037 , n17069 , n17077 , n17090 , 
n17095 , n17250 , n17251 , n17302 , n17351 , n17458 , n17664 , n17784 , n17911 , n17954 , 
n17959 , n17968 , n18035 , n18105 , n18145 , n18151 , n18157 , n18171 , n18227 , n18274 , 
n18290 , n18295 , n18345 , n18409 , n18444 , n18452 , n18483 , n18496 , n18537 , n18558 , 
n18578 , n18584 , n18649 , n18690 , n18737 , n18745 , n18880 , n18901 , n18907 , n18926 , 
n18962 , n19005 , n19033 , n19042 , n19081 , n19107 , n19116 , n19144 , n19163 , n19196 , 
n19228 , n19234 , n19270 , n19282 , n19327 , n19357 , n19361 , n19454 , n19472 , n19477 , 
n19494 , n19514 , n19515 , n19531 , n19539 , n19575 , n19584 , n19608 , n19618 , n19652 , 
n19680 , n19701 , n19770 , n19789 , n19803 , n19905 , n19911 , n19922 , n19941 , n20013 , 
n20036 , n20040 , n20077 , n20138 , n20151 , n20169 , n20179 , n20213 , n20235 , n20250 , 
n20259 , n20349 , n20359 , n20385 , n20409 , n20411 , n20429 , n20455 , n20470 , n20478 , 
n20489 , n20604 , n20658 , n20700 , n20794 , n20826 , n20923 , n20929 , n20946 , n20986 , 
n21078 , n21095 , n21134 , n21138 , n21222 , n21226 , n21276 , n21287 , n21317 , n21398 , 
n21471 , n21489 , n21538 , n21599 , n21649 , n21654 , n21674 , n21687 , n21735 , n21749 , 
n21753 , n21779 , n21784 , n21832 , n21839 , n21898 , n21905 , n21915 , n21934 , n21957 , 
n21981 , n21993 , n21997 , n22043 , n22068 , n22072 , n22173 , n22198 , n22201 , n22253 , 
n22270 , n22274 , n22290 , n22309 , n22332 , n22335 , n22358 , n22359 , n22379 , n22433 , 
n22442 , n22470 , n22492 , n22554 , n22588 , n22591 , n22597 , n22619 , n22626 , n22631 , 
n22660 , n22764 , n22793 , n22843 , n22871 , n22879 , n22918 , n23035 , n23039 , n23065 , 
n23068 , n23120 , n23146 , n23160 , n23166 , n23200 , n23250 , n23272 , n23304 , n23333 , 
n23369 , n23430 , n23463 , n23493 , n23513 , n23529 , n23541 , n23586 , n23657 , n23697 , 
n23717 , n23755 , n23775 , n23831 , n23842 , n23849 , n23895 , n23912 , n23913 , n23923 , 
n23974 , n24004 , n24032 , n24048 , n24085 , n24093 , n24129 , n24150 , n24170 , n24196 , 
n24278 , n24319 , n24323 , n24327 , n24374 , n24485 , n24618 , n24620 , n24638 , n24732 , 
n24768 , n24786 , n24879 , n24937 , n25023 , n25068 , n25073 , n25074 , n25094 , n25119 , 
n25120 , n25126 , n25168 , n25240 , n25296 , n25316 , n25331 , n25336 , n25345 , n25365 , 
n25370 , n25381 , n25435 , n25464 , n25471 , n25475 , n25494 , n25523 , n25565 , n25586 , 
n25629 , n25643 , n25694 , n25738 , n25749 , n25751 , n25797 , n25872 , n25877 , n25923 , 
n25926 , n25972 , n25974 , n26036 , n26053 , n26054 , n26107 , n26167 , n26180 , n26191 , 
n26224 , n26264 , n26318 , n26408 , n26443 , n26452 , n26483 , n26510 , n26512 , n26553 , 
n26565 , n26572 , n26625 , n26660 , n26725 , n26744 , n26748 , n26752 , n26797 , n26808 , 
n26823 , n26882 , n26913 , n26979 , n26986 , n27037 , n27089 , n27104 , n27120 , n27134 , 
n27188 ;
    output n7 , n50 , n55 , n108 , n142 , n175 , n235 , n242 , n243 , 
n248 , n266 , n298 , n317 , n332 , n357 , n422 , n431 , n457 , n463 , 
n491 , n496 , n498 , n521 , n548 , n554 , n567 , n588 , n597 , n637 , 
n646 , n696 , n723 , n735 , n779 , n809 , n819 , n829 , n849 , n858 , 
n873 , n879 , n887 , n904 , n948 , n957 , n980 , n982 , n984 , n1005 , 
n1016 , n1020 , n1044 , n1060 , n1069 , n1111 , n1119 , n1120 , n1196 , n1237 , 
n1239 , n1302 , n1332 , n1357 , n1371 , n1385 , n1498 , n1501 , n1518 , n1527 , 
n1580 , n1586 , n1590 , n1602 , n1634 , n1636 , n1684 , n1701 , n1703 , n1721 , 
n1760 , n1791 , n1808 , n1821 , n1832 , n1859 , n1860 , n1861 , n1891 , n1925 , 
n1942 , n1972 , n1981 , n2004 , n2007 , n2061 , n2092 , n2095 , n2105 , n2122 , 
n2147 , n2209 , n2214 , n2238 , n2327 , n2343 , n2361 , n2363 , n2374 , n2388 , 
n2440 , n2444 , n2513 , n2515 , n2533 , n2535 , n2537 , n2553 , n2555 , n2560 , 
n2561 , n2573 , n2578 , n2582 , n2602 , n2619 , n2661 , n2693 , n2703 , n2706 , 
n2711 , n2761 , n2774 , n2779 , n2826 , n2853 , n2860 , n2887 , n2929 , n2948 , 
n2961 , n2971 , n3010 , n3017 , n3020 , n3067 , n3076 , n3089 , n3125 , n3126 , 
n3208 , n3219 , n3235 , n3244 , n3263 , n3289 , n3301 , n3316 , n3332 , n3340 , 
n3343 , n3390 , n3426 , n3451 , n3459 , n3502 , n3516 , n3528 , n3555 , n3561 , 
n3563 , n3617 , n3642 , n3649 , n3665 , n3679 , n3725 , n3733 , n3755 , n3758 , 
n3760 , n3781 , n3794 , n3842 , n3850 , n3869 , n3871 , n3891 , n3932 , n3934 , 
n3971 , n3983 , n4000 , n4010 , n4014 , n4071 , n4088 , n4089 , n4103 , n4123 , 
n4134 , n4146 , n4150 , n4151 , n4152 , n4153 , n4165 , n4172 , n4173 , n4176 , 
n4186 , n4204 , n4205 , n4215 , n4221 , n4224 , n4231 , n4266 , n4340 , n4374 , 
n4401 , n4424 , n4432 , n4441 , n4451 , n4476 , n4478 , n4529 , n4552 , n4595 , 
n4624 , n4646 , n4674 , n4693 , n4731 , n4745 , n4747 , n4766 , n4770 , n4777 , 
n4785 , n4804 , n4810 , n4814 , n4850 , n4891 , n4925 , n4947 , n4952 , n4966 , 
n4972 , n5011 , n5020 , n5024 , n5046 , n5062 , n5064 , n5082 , n5120 , n5158 , 
n5168 , n5184 , n5228 , n5256 , n5265 , n5273 , n5274 , n5300 , n5325 , n5351 , 
n5353 , n5399 , n5403 , n5430 , n5439 , n5472 , n5485 , n5524 , n5564 , n5593 , 
n5603 , n5609 , n5634 , n5643 , n5680 , n5687 , n5700 , n5732 , n5742 , n5765 , 
n5776 , n5782 , n5833 , n5840 , n5841 , n5850 , n5903 , n5904 , n5911 , n5936 , 
n5943 , n5964 , n5980 , n6012 , n6022 , n6031 , n6044 , n6046 , n6084 , n6160 , 
n6171 , n6183 , n6189 , n6223 , n6233 , n6245 , n6248 , n6256 , n6271 , n6276 , 
n6308 , n6311 , n6323 , n6330 , n6339 , n6354 , n6375 , n6383 , n6407 , n6431 , 
n6437 , n6457 , n6465 , n6470 , n6476 , n6506 , n6514 , n6542 , n6558 , n6560 , 
n6567 , n6576 , n6587 , n6612 , n6628 , n6630 , n6634 , n6652 , n6655 , n6669 , 
n6671 , n6673 , n6674 , n6684 , n6706 , n6707 , n6736 , n6791 , n6802 , n6826 , 
n6835 , n6853 , n6862 , n6863 , n6867 , n6965 , n6967 , n6975 , n6983 , n6985 , 
n6998 , n7032 , n7038 , n7079 , n7190 , n7229 , n7230 , n7233 , n7236 , n7253 , 
n7256 , n7268 , n7277 , n7280 , n7298 , n7308 , n7313 , n7346 , n7349 , n7363 , 
n7390 , n7403 , n7408 , n7432 , n7475 , n7477 , n7507 , n7514 , n7558 , n7572 , 
n7575 , n7585 , n7588 , n7598 , n7607 , n7610 , n7616 , n7630 , n7643 , n7647 , 
n7679 , n7686 , n7698 , n7708 , n7780 , n7794 , n7811 , n7830 , n7834 , n7884 , 
n7937 , n7943 , n7950 , n7959 , n7968 , n7992 , n7999 , n8027 , n8031 , n8042 , 
n8095 , n8103 , n8109 , n8127 , n8130 , n8135 , n8139 , n8148 , n8149 , n8159 , 
n8179 , n8215 , n8267 , n8276 , n8288 , n8306 , n8320 , n8321 , n8339 , n8376 , 
n8408 , n8417 , n8432 , n8453 , n8480 , n8489 , n8505 , n8510 , n8519 , n8535 , 
n8550 , n8563 , n8594 , n8608 , n8620 , n8637 , n8662 , n8716 , n8744 , n8803 , 
n8809 , n8821 , n8824 , n8849 , n8861 , n8862 , n8884 , n8909 , n8911 , n8971 , 
n8982 , n8993 , n9012 , n9032 , n9042 , n9046 , n9047 , n9104 , n9129 , n9146 , 
n9164 , n9166 , n9182 , n9191 , n9217 , n9220 , n9261 , n9287 , n9308 , n9344 , 
n9364 , n9371 , n9382 , n9403 , n9419 , n9423 , n9430 , n9435 , n9451 , n9458 , 
n9459 , n9508 , n9552 , n9556 , n9558 , n9616 , n9622 , n9626 , n9633 , n9635 , 
n9648 , n9689 , n9695 , n9699 , n9726 , n9753 , n9761 , n9763 , n9767 , n9771 , 
n9778 , n9783 , n9803 , n9833 , n9838 , n9867 , n9890 , n9917 , n9919 , n9938 , 
n9946 , n9968 , n10009 , n10010 , n10019 , n10021 , n10055 , n10101 , n10111 , n10165 , 
n10236 , n10239 , n10244 , n10261 , n10262 , n10287 , n10295 , n10321 , n10326 , n10327 , 
n10330 , n10340 , n10345 , n10356 , n10385 , n10387 , n10388 , n10390 , n10404 , n10409 , 
n10420 , n10432 , n10484 , n10489 , n10525 , n10540 , n10561 , n10564 , n10588 , n10595 , 
n10617 , n10628 , n10647 , n10653 , n10692 , n10694 , n10701 , n10756 , n10775 , n10780 , 
n10817 , n10834 , n10851 , n10874 , n10924 , n10943 , n10961 , n11005 , n11023 , n11025 , 
n11063 , n11078 , n11080 , n11094 , n11101 , n11103 , n11120 , n11127 , n11132 , n11134 , 
n11138 , n11182 , n11234 , n11245 , n11261 , n11275 , n11290 , n11313 , n11325 , n11326 , 
n11330 , n11347 , n11348 , n11352 , n11375 , n11379 , n11386 , n11391 , n11398 , n11403 , 
n11419 , n11439 , n11462 , n11470 , n11472 , n11496 , n11506 , n11515 , n11538 , n11548 , 
n11564 , n11591 , n11607 , n11647 , n11674 , n11682 , n11710 , n11712 , n11724 , n11741 , 
n11770 , n11771 , n11818 , n11837 , n11842 , n11843 , n11905 , n11965 , n12000 , n12003 , 
n12011 , n12072 , n12131 , n12146 , n12157 , n12158 , n12179 , n12192 , n12223 , n12225 , 
n12228 , n12235 , n12302 , n12304 , n12324 , n12325 , n12329 , n12330 , n12346 , n12349 , 
n12364 , n12383 , n12397 , n12408 , n12449 , n12461 , n12462 , n12467 , n12469 , n12515 , 
n12516 , n12540 , n12545 , n12552 , n12566 , n12569 , n12607 , n12620 , n12621 , n12654 , 
n12665 , n12670 , n12707 , n12725 , n12727 , n12740 , n12742 , n12746 , n12756 , n12783 , 
n12801 , n12812 , n12816 , n12843 , n12864 , n12865 , n12870 , n12873 , n12904 , n12941 , 
n12942 , n12978 , n12980 , n12985 , n12987 , n12992 , n13005 , n13043 , n13048 , n13054 , 
n13082 , n13096 , n13116 , n13122 , n13141 , n13144 , n13168 , n13198 , n13199 , n13204 , 
n13209 , n13270 , n13273 , n13285 , n13338 , n13407 , n13409 , n13456 , n13457 , n13477 , 
n13484 , n13486 , n13487 , n13500 , n13501 , n13506 , n13548 , n13551 , n13602 , n13626 , 
n13683 , n13710 , n13722 , n13754 , n13764 , n13798 , n13835 , n13850 , n13922 , n13923 , 
n14004 , n14036 , n14059 , n14081 , n14095 , n14107 , n14121 , n14126 , n14136 , n14147 , 
n14174 , n14190 , n14211 , n14222 , n14267 , n14271 , n14277 , n14294 , n14310 , n14326 , 
n14342 , n14353 , n14364 , n14375 , n14412 , n14414 , n14457 , n14464 , n14471 , n14475 , 
n14541 , n14546 , n14547 , n14593 , n14636 , n14701 , n14734 , n14746 , n14763 , n14772 , 
n14801 , n14819 , n14827 , n14839 , n14849 , n14891 , n14931 , n14944 , n14977 , n14989 , 
n15002 , n15004 , n15011 , n15019 , n15031 , n15033 , n15052 , n15082 , n15094 , n15118 , 
n15128 , n15139 , n15145 , n15165 , n15176 , n15180 , n15205 , n15230 , n15255 , n15275 , 
n15300 , n15307 , n15327 , n15345 , n15353 , n15366 , n15382 , n15407 , n15428 , n15435 , 
n15438 , n15465 , n15467 , n15470 , n15477 , n15481 , n15496 , n15501 , n15555 , n15558 , 
n15559 , n15570 , n15573 , n15588 , n15590 , n15598 , n15614 , n15662 , n15716 , n15749 , 
n15762 , n15793 , n15812 , n15815 , n15816 , n15831 , n15846 , n15859 , n15869 , n15885 , 
n15889 , n15917 , n15922 , n15947 , n15956 , n15958 , n15986 , n16013 , n16060 , n16062 , 
n16068 , n16080 , n16098 , n16110 , n16142 , n16185 , n16196 , n16206 , n16215 , n16218 , 
n16219 , n16230 , n16243 , n16275 , n16279 , n16322 , n16327 , n16350 , n16367 , n16379 , 
n16398 , n16406 , n16407 , n16419 , n16424 , n16428 , n16433 , n16440 , n16445 , n16460 , 
n16481 , n16493 , n16506 , n16516 , n16517 , n16527 , n16554 , n16583 , n16584 , n16589 , 
n16596 , n16617 , n16630 , n16640 , n16656 , n16674 , n16682 , n16684 , n16688 , n16733 , 
n16798 , n16834 , n16837 , n16841 , n16885 , n16905 , n16951 , n16954 , n16989 , n17006 , 
n17068 , n17070 , n17075 , n17084 , n17104 , n17106 , n17119 , n17130 , n17138 , n17163 , 
n17168 , n17202 , n17219 , n17232 , n17236 , n17243 , n17263 , n17285 , n17320 , n17337 , 
n17344 , n17359 , n17387 , n17391 , n17392 , n17421 , n17432 , n17436 , n17440 , n17450 , 
n17461 , n17466 , n17493 , n17500 , n17524 , n17529 , n17557 , n17583 , n17592 , n17638 , 
n17687 , n17721 , n17735 , n17738 , n17746 , n17749 , n17820 , n17855 , n17877 , n17889 , 
n17912 , n17927 , n17931 , n17948 , n17956 , n17963 , n17976 , n17998 , n18025 , n18043 , 
n18045 , n18059 , n18061 , n18071 , n18143 , n18152 , n18193 , n18232 , n18238 , n18241 , 
n18254 , n18288 , n18301 , n18304 , n18310 , n18311 , n18323 , n18332 , n18343 , n18350 , 
n18362 , n18377 , n18405 , n18414 , n18418 , n18437 , n18439 , n18445 , n18467 , n18482 , 
n18509 , n18513 , n18515 , n18572 , n18574 , n18576 , n18582 , n18583 , n18610 , n18635 , 
n18653 , n18679 , n18693 , n18708 , n18721 , n18725 , n18751 , n18780 , n18782 , n18802 , 
n18830 , n18831 , n18843 , n18858 , n18859 , n18864 , n18865 , n18886 , n18887 , n18919 , 
n18940 , n18945 , n18970 , n18977 , n18982 , n18999 , n19044 , n19125 , n19141 , n19164 , 
n19174 , n19176 , n19202 , n19220 , n19221 , n19223 , n19224 , n19233 , n19244 , n19314 , 
n19315 , n19323 , n19333 , n19348 , n19354 , n19367 , n19385 , n19389 , n19401 , n19414 , 
n19424 , n19450 , n19458 , n19467 , n19496 , n19523 , n19570 , n19602 , n19617 , n19623 , 
n19641 , n19648 , n19664 , n19736 , n19749 , n19756 , n19767 , n19780 , n19792 , n19798 , 
n19873 , n19909 , n19916 , n19923 , n19930 , n19968 , n19988 , n20004 , n20017 , n20033 , 
n20061 , n20069 , n20086 , n20096 , n20103 , n20126 , n20149 , n20187 , n20279 , n20287 , 
n20301 , n20330 , n20333 , n20355 , n20366 , n20388 , n20402 , n20403 , n20424 , n20436 , 
n20441 , n20445 , n20450 , n20490 , n20495 , n20515 , n20533 , n20582 , n20590 , n20602 , 
n20609 , n20623 , n20629 , n20661 , n20673 , n20678 , n20680 , n20685 , n20691 , n20696 , 
n20704 , n20705 , n20709 , n20713 , n20722 , n20723 , n20748 , n20761 , n20774 , n20788 , 
n20795 , n20803 , n20869 , n20879 , n20915 , n20935 , n20936 , n21008 , n21017 , n21034 , 
n21046 , n21062 , n21093 , n21094 , n21123 , n21154 , n21157 , n21168 , n21173 , n21176 , 
n21182 , n21193 , n21203 , n21225 , n21238 , n21254 , n21298 , n21302 , n21349 , n21365 , 
n21367 , n21396 , n21399 , n21404 , n21446 , n21472 , n21525 , n21549 , n21615 , n21628 , 
n21637 , n21645 , n21665 , n21680 , n21685 , n21717 , n21719 , n21750 , n21765 , n21800 , 
n21820 , n21874 , n21943 , n21960 , n21976 , n21986 , n22016 , n22027 , n22050 , n22063 , 
n22076 , n22090 , n22107 , n22113 , n22124 , n22126 , n22130 , n22144 , n22150 , n22157 , 
n22213 , n22283 , n22311 , n22317 , n22341 , n22353 , n22444 , n22467 , n22484 , n22489 , 
n22494 , n22533 , n22584 , n22589 , n22620 , n22623 , n22697 , n22714 , n22761 , n22779 , 
n22787 , n22819 , n22858 , n22870 , n22891 , n22897 , n22903 , n22907 , n22910 , n22914 , 
n22939 , n22998 , n23006 , n23007 , n23009 , n23014 , n23047 , n23058 , n23066 , n23067 , 
n23238 , n23247 , n23248 , n23270 , n23289 , n23305 , n23341 , n23342 , n23355 , n23371 , 
n23401 , n23414 , n23429 , n23433 , n23434 , n23450 , n23471 , n23480 , n23546 , n23550 , 
n23585 , n23588 , n23619 , n23624 , n23628 , n23637 , n23663 , n23669 , n23684 , n23690 , 
n23714 , n23719 , n23748 , n23856 , n23883 , n23888 , n23899 , n23903 , n23924 , n23935 , 
n23942 , n23954 , n23958 , n23986 , n24002 , n24039 , n24052 , n24092 , n24096 , n24097 , 
n24105 , n24119 , n24133 , n24141 , n24145 , n24146 , n24155 , n24160 , n24167 , n24172 , 
n24177 , n24228 , n24258 , n24260 , n24289 , n24297 , n24307 , n24342 , n24345 , n24347 , 
n24373 , n24406 , n24415 , n24421 , n24431 , n24472 , n24476 , n24483 , n24501 , n24512 , 
n24558 , n24576 , n24579 , n24602 , n24604 , n24626 , n24629 , n24636 , n24715 , n24723 , 
n24749 , n24758 , n24784 , n24807 , n24826 , n24840 , n24841 , n24853 , n24857 , n24887 , 
n24934 , n24998 , n25006 , n25032 , n25062 , n25083 , n25097 , n25133 , n25155 , n25181 , 
n25200 , n25209 , n25215 , n25244 , n25254 , n25256 , n25293 , n25328 , n25332 , n25337 , 
n25356 , n25362 , n25412 , n25460 , n25468 , n25499 , n25513 , n25518 , n25532 , n25539 , 
n25550 , n25611 , n25614 , n25619 , n25665 , n25706 , n25719 , n25756 , n25758 , n25773 , 
n25784 , n25792 , n25816 , n25826 , n25839 , n25840 , n25873 , n25934 , n25938 , n25985 , 
n25994 , n26084 , n26096 , n26111 , n26113 , n26156 , n26159 , n26179 , n26220 , n26229 , 
n26237 , n26250 , n26274 , n26287 , n26317 , n26353 , n26375 , n26396 , n26429 , n26431 , 
n26439 , n26492 , n26515 , n26538 , n26590 , n26598 , n26605 , n26656 , n26674 , n26675 , 
n26681 , n26696 , n26698 , n26707 , n26719 , n26727 , n26729 , n26745 , n26775 , n26780 , 
n26794 , n26795 , n26801 , n26815 , n26847 , n26900 , n26902 , n26905 , n26921 , n26923 , 
n26929 , n26930 , n26943 , n26970 , n27004 , n27011 , n27019 , n27031 , n27051 , n27072 , 
n27079 , n27096 , n27110 , n27112 , n27130 , n27145 , n27158 , n27163 , n27194 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n8 , n9 , 
n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n19 , n20 , 
n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , 
n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , 
n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n51 , n52 , 
n53 , n54 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , 
n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , 
n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , 
n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , 
n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , 
n104 , n105 , n106 , n107 , n109 , n110 , n111 , n112 , n113 , n114 , 
n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , 
n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , 
n135 , n136 , n137 , n138 , n139 , n140 , n141 , n143 , n144 , n145 , 
n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , 
n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , 
n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n176 , 
n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , 
n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n197 , 
n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , 
n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , 
n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , 
n228 , n229 , n230 , n231 , n232 , n233 , n234 , n236 , n237 , n238 , 
n239 , n240 , n241 , n244 , n245 , n246 , n247 , n249 , n250 , n251 , 
n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , 
n262 , n263 , n264 , n265 , n267 , n269 , n270 , n271 , n272 , n273 , 
n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , 
n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , 
n294 , n295 , n296 , n297 , n299 , n300 , n301 , n302 , n303 , n304 , 
n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , 
n315 , n316 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , 
n326 , n327 , n328 , n330 , n331 , n333 , n334 , n335 , n336 , n338 , 
n339 , n340 , n341 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
n350 , n351 , n352 , n353 , n354 , n355 , n356 , n358 , n359 , n360 , 
n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , 
n371 , n372 , n373 , n374 , n375 , n377 , n378 , n379 , n380 , n381 , 
n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , 
n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , 
n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , 
n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , 
n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n432 , n433 , 
n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n443 , n444 , 
n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , 
n455 , n456 , n458 , n459 , n460 , n461 , n462 , n464 , n465 , n466 , 
n467 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , 
n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , 
n488 , n489 , n490 , n492 , n493 , n494 , n495 , n497 , n499 , n500 , 
n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , 
n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , 
n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , 
n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , 
n542 , n543 , n544 , n545 , n546 , n547 , n549 , n550 , n551 , n552 , 
n553 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , 
n564 , n565 , n566 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n584 , n585 , 
n586 , n587 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , 
n598 , n599 , n600 , n601 , n602 , n603 , n605 , n606 , n607 , n608 , 
n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , 
n619 , n620 , n621 , n622 , n623 , n624 , n625 , n627 , n628 , n629 , 
n630 , n631 , n632 , n633 , n634 , n635 , n636 , n638 , n639 , n640 , 
n641 , n642 , n643 , n644 , n645 , n648 , n649 , n650 , n651 , n652 , 
n653 , n654 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , 
n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , 
n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , 
n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , 
n694 , n695 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , 
n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , 
n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n724 , n725 , 
n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n736 , 
n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , 
n747 , n748 , n749 , n750 , n751 , n753 , n754 , n755 , n756 , n757 , 
n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n768 , 
n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , 
n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n810 , 
n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n820 , n821 , 
n822 , n823 , n824 , n825 , n826 , n827 , n828 , n830 , n831 , n832 , 
n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , 
n843 , n844 , n845 , n846 , n847 , n848 , n850 , n851 , n852 , n853 , 
n854 , n855 , n856 , n857 , n859 , n860 , n861 , n862 , n863 , n864 , 
n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n874 , n875 , 
n876 , n877 , n878 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , 
n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , 
n898 , n899 , n900 , n901 , n902 , n903 , n905 , n906 , n907 , n908 , 
n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , 
n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
n930 , n931 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , 
n941 , n942 , n943 , n944 , n945 , n946 , n947 , n949 , n950 , n951 , 
n952 , n953 , n954 , n955 , n956 , n958 , n959 , n960 , n961 , n962 , 
n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , 
n973 , n974 , n975 , n976 , n977 , n978 , n979 , n981 , n983 , n985 , 
n986 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , 
n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1006 , n1007 , 
n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1017 , n1018 , 
n1019 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
n1041 , n1042 , n1043 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , 
n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1061 , n1062 , 
n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1070 , n1071 , n1072 , n1073 , 
n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , 
n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , 
n1094 , n1095 , n1096 , n1097 , n1098 , n1100 , n1101 , n1102 , n1103 , n1104 , 
n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1113 , n1114 , n1115 , n1116 , 
n1117 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1137 , n1138 , n1139 , n1140 , 
n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , 
n1151 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , 
n1162 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , 
n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , 
n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , 
n1193 , n1194 , n1195 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , 
n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , 
n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1223 , n1224 , n1225 , 
n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , 
n1236 , n1238 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , 
n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1256 , n1257 , n1258 , 
n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , 
n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1280 , 
n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1289 , n1290 , n1291 , 
n1292 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1303 , 
n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , 
n1315 , n1316 , n1317 , n1318 , n1319 , n1321 , n1322 , n1323 , n1324 , n1325 , 
n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1333 , n1334 , n1335 , n1336 , 
n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , 
n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , 
n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , 
n1368 , n1369 , n1370 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , 
n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1386 , n1387 , n1388 , n1389 , 
n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
n1430 , n1431 , n1433 , n1434 , n1435 , n1436 , n1438 , n1439 , n1440 , n1441 , 
n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1452 , 
n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , 
n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , 
n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , 
n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , 
n1494 , n1495 , n1496 , n1497 , n1499 , n1500 , n1502 , n1503 , n1504 , n1505 , 
n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , 
n1516 , n1517 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1526 , n1528 , 
n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1537 , n1538 , n1539 , 
n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1559 , n1560 , 
n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , 
n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1581 , 
n1582 , n1583 , n1584 , n1585 , n1587 , n1588 , n1589 , n1591 , n1592 , n1593 , 
n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1603 , n1604 , 
n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1612 , n1613 , n1614 , n1615 , 
n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , 
n1626 , n1627 , n1628 , n1629 , n1631 , n1632 , n1633 , n1635 , n1637 , n1638 , 
n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
n1650 , n1651 , n1652 , n1653 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , 
n1661 , n1663 , n1664 , n1665 , n1666 , n1668 , n1669 , n1670 , n1671 , n1672 , 
n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1683 , n1685 , 
n1686 , n1687 , n1688 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , 
n1697 , n1698 , n1699 , n1700 , n1702 , n1704 , n1705 , n1706 , n1707 , n1708 , 
n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , 
n1719 , n1720 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1739 , n1740 , 
n1741 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , 
n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1761 , n1762 , n1763 , 
n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , 
n1774 , n1775 , n1776 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , 
n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1792 , n1793 , n1794 , n1795 , 
n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , 
n1806 , n1807 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , 
n1817 , n1818 , n1819 , n1820 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , 
n1828 , n1829 , n1830 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1862 , 
n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , 
n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1882 , n1883 , 
n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1892 , n1893 , n1894 , 
n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , 
n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , 
n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , 
n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , 
n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1943 , n1944 , n1945 , n1946 , 
n1947 , n1948 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , 
n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , 
n1968 , n1969 , n1970 , n1971 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , 
n1979 , n1980 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n2000 , 
n2001 , n2002 , n2003 , n2005 , n2006 , n2008 , n2009 , n2010 , n2011 , n2012 , 
n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , 
n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , 
n2034 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , 
n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , 
n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2062 , n2063 , n2064 , n2065 , 
n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , 
n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , 
n2086 , n2087 , n2089 , n2090 , n2091 , n2093 , n2094 , n2096 , n2097 , n2098 , 
n2099 , n2100 , n2101 , n2103 , n2104 , n2106 , n2107 , n2108 , n2109 , n2110 , 
n2111 , n2112 , n2114 , n2115 , n2116 , n2118 , n2119 , n2120 , n2121 , n2123 , 
n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , 
n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , 
n2144 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , 
n2157 , n2158 , n2159 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , 
n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2176 , n2177 , n2178 , 
n2179 , n2180 , n2181 , n2182 , n2183 , n2185 , n2186 , n2187 , n2188 , n2189 , 
n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2211 , 
n2212 , n2213 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , 
n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , 
n2233 , n2234 , n2235 , n2236 , n2237 , n2239 , n2240 , n2241 , n2242 , n2243 , 
n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , 
n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , 
n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2273 , n2274 , 
n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , 
n2285 , n2286 , n2287 , n2288 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , 
n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , 
n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , 
n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , 
n2326 , n2329 , n2330 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , 
n2339 , n2340 , n2341 , n2342 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
n2350 , n2351 , n2352 , n2353 , n2354 , n2356 , n2357 , n2358 , n2359 , n2360 , 
n2362 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , 
n2373 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , 
n2384 , n2385 , n2386 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , 
n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , 
n2406 , n2407 , n2408 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2417 , 
n2418 , n2419 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
n2441 , n2442 , n2443 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , 
n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , 
n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , 
n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2480 , n2481 , n2482 , 
n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , 
n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , 
n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , 
n2514 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , 
n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2534 , n2536 , 
n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2548 , 
n2549 , n2550 , n2551 , n2552 , n2554 , n2556 , n2557 , n2558 , n2559 , n2562 , 
n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2571 , n2572 , n2574 , 
n2575 , n2576 , n2577 , n2579 , n2580 , n2581 , n2583 , n2584 , n2585 , n2586 , 
n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , 
n2597 , n2598 , n2599 , n2600 , n2601 , n2603 , n2604 , n2605 , n2606 , n2607 , 
n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , 
n2618 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , 
n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , 
n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2647 , n2648 , n2649 , 
n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2660 , 
n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , 
n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2681 , n2682 , 
n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , 
n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2704 , 
n2705 , n2707 , n2708 , n2709 , n2710 , n2712 , n2713 , n2714 , n2715 , n2716 , 
n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , 
n2727 , n2728 , n2729 , n2730 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , 
n2738 , n2739 , n2740 , n2741 , n2742 , n2744 , n2745 , n2746 , n2747 , n2748 , 
n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , 
n2759 , n2760 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
n2770 , n2771 , n2772 , n2773 , n2775 , n2776 , n2777 , n2778 , n2780 , n2781 , 
n2782 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , 
n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , 
n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2810 , n2811 , n2812 , n2813 , 
n2814 , n2815 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , 
n2825 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , 
n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , 
n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2854 , n2855 , n2856 , 
n2857 , n2859 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , 
n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , 
n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2888 , n2889 , n2890 , 
n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , 
n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , 
n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , 
n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2930 , n2931 , 
n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , 
n2942 , n2943 , n2945 , n2946 , n2947 , n2949 , n2950 , n2951 , n2952 , n2953 , 
n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2962 , n2963 , n2964 , 
n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2972 , n2973 , n2974 , n2975 , 
n2976 , n2977 , n2980 , n2981 , n2982 , n2983 , n2984 , n2986 , n2987 , n2988 , 
n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , 
n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3019 , n3021 , n3022 , n3023 , 
n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3031 , n3032 , n3033 , n3034 , 
n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , 
n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , 
n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , 
n3065 , n3066 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , 
n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , 
n3087 , n3088 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , 
n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , 
n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , 
n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3127 , n3128 , n3129 , 
n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3137 , n3138 , n3139 , n3140 , 
n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , 
n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , 
n3162 , n3163 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , 
n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , 
n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , 
n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , 
n3203 , n3204 , n3205 , n3206 , n3207 , n3209 , n3210 , n3211 , n3212 , n3213 , 
n3214 , n3215 , n3216 , n3217 , n3218 , n3220 , n3221 , n3222 , n3223 , n3224 , 
n3225 , n3226 , n3227 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3236 , 
n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3245 , n3246 , n3247 , 
n3248 , n3249 , n3250 , n3251 , n3252 , n3254 , n3255 , n3256 , n3257 , n3258 , 
n3259 , n3261 , n3262 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , 
n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3280 , n3281 , 
n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3290 , n3291 , n3292 , 
n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3302 , n3303 , 
n3304 , n3305 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , 
n3315 , n3317 , n3318 , n3319 , n3321 , n3322 , n3323 , n3325 , n3326 , n3327 , 
n3328 , n3329 , n3330 , n3331 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , 
n3339 , n3341 , n3342 , n3344 , n3345 , n3346 , n3347 , n3348 , n3350 , n3351 , 
n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , 
n3362 , n3363 , n3364 , n3365 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , 
n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , 
n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3391 , n3392 , n3393 , 
n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , 
n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , 
n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , 
n3424 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , 
n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , 
n3446 , n3447 , n3448 , n3449 , n3450 , n3452 , n3453 , n3454 , n3455 , n3456 , 
n3457 , n3458 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3469 , 
n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
n3501 , n3503 , n3504 , n3505 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , 
n3513 , n3514 , n3515 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , 
n3524 , n3525 , n3526 , n3527 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , 
n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3542 , n3543 , n3544 , n3545 , 
n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3556 , 
n3557 , n3558 , n3559 , n3560 , n3562 , n3564 , n3565 , n3566 , n3567 , n3568 , 
n3569 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
n3580 , n3581 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , 
n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , 
n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , 
n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3619 , n3620 , n3621 , n3622 , 
n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , 
n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3643 , 
n3644 , n3645 , n3646 , n3647 , n3648 , n3650 , n3651 , n3652 , n3653 , n3654 , 
n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , 
n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , 
n3676 , n3677 , n3678 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , 
n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , 
n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , 
n3707 , n3708 , n3709 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , 
n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3726 , n3727 , n3728 , 
n3729 , n3730 , n3731 , n3732 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , 
n3751 , n3752 , n3753 , n3754 , n3756 , n3757 , n3759 , n3761 , n3762 , n3763 , 
n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , 
n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3782 , n3783 , n3784 , 
n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3796 , n3797 , 
n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , 
n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , 
n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , 
n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , 
n3839 , n3840 , n3841 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , 
n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , 
n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3870 , n3872 , 
n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , 
n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3892 , n3893 , 
n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , 
n3904 , n3905 , n3906 , n3907 , n3908 , n3910 , n3911 , n3912 , n3913 , n3914 , 
n3915 , n3916 , n3917 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3926 , 
n3927 , n3928 , n3929 , n3930 , n3931 , n3933 , n3935 , n3936 , n3937 , n3938 , 
n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3946 , n3947 , n3948 , n3949 , 
n3950 , n3951 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3960 , n3961 , 
n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3972 , n3973 , 
n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3985 , 
n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , 
n3996 , n3997 , n3998 , n3999 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , 
n4007 , n4008 , n4009 , n4011 , n4012 , n4013 , n4015 , n4016 , n4017 , n4018 , 
n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , 
n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , 
n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , 
n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , 
n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , 
n4069 , n4070 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , 
n4080 , n4081 , n4082 , n4083 , n4084 , n4086 , n4087 , n4090 , n4091 , n4092 , 
n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4101 , n4102 , n4104 , 
n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , 
n4115 , n4116 , n4117 , n4118 , n4120 , n4121 , n4122 , n4124 , n4125 , n4126 , 
n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4135 , n4136 , n4137 , 
n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4147 , n4148 , 
n4149 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , 
n4163 , n4164 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4174 , n4175 , 
n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4187 , 
n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , 
n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4206 , n4207 , n4208 , n4209 , 
n4210 , n4211 , n4212 , n4213 , n4214 , n4216 , n4217 , n4218 , n4219 , n4220 , 
n4222 , n4223 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4232 , n4233 , 
n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , 
n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , 
n4254 , n4255 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , 
n4265 , n4267 , n4268 , n4269 , n4270 , n4271 , n4273 , n4274 , n4275 , n4276 , 
n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , 
n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , 
n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4307 , 
n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , 
n4318 , n4320 , n4321 , n4322 , n4323 , n4324 , n4327 , n4328 , n4329 , n4330 , 
n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4341 , 
n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , 
n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , 
n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , 
n4372 , n4373 , n4375 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , 
n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , 
n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4402 , n4403 , n4404 , 
n4405 , n4406 , n4407 , n4408 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , 
n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4425 , n4427 , 
n4428 , n4429 , n4430 , n4431 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , 
n4439 , n4440 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , 
n4450 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
n4471 , n4472 , n4473 , n4474 , n4475 , n4477 , n4479 , n4480 , n4481 , n4482 , 
n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , 
n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , 
n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , 
n4513 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , 
n4524 , n4525 , n4526 , n4527 , n4528 , n4530 , n4531 , n4532 , n4533 , n4534 , 
n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , 
n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4553 , n4554 , n4555 , 
n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , 
n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , 
n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , 
n4586 , n4587 , n4589 , n4591 , n4592 , n4593 , n4594 , n4596 , n4597 , n4598 , 
n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , 
n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , 
n4619 , n4620 , n4621 , n4622 , n4623 , n4625 , n4626 , n4627 , n4628 , n4629 , 
n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , 
n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4647 , n4648 , n4649 , n4650 , 
n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
n4661 , n4662 , n4663 , n4664 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , 
n4672 , n4673 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , 
n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , 
n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , 
n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , 
n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4723 , n4724 , 
n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4732 , n4733 , n4734 , n4735 , 
n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4746 , 
n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , 
n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4767 , n4768 , 
n4769 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4778 , n4779 , n4780 , 
n4781 , n4782 , n4783 , n4784 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , 
n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , 
n4802 , n4803 , n4805 , n4806 , n4807 , n4808 , n4809 , n4811 , n4813 , n4815 , 
n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , 
n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , 
n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , 
n4846 , n4847 , n4848 , n4849 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , 
n4857 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , 
n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , 
n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , 
n4888 , n4889 , n4890 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , 
n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , 
n4909 , n4910 , n4911 , n4912 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , 
n4920 , n4921 , n4922 , n4923 , n4924 , n4926 , n4927 , n4928 , n4929 , n4930 , 
n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4940 , n4941 , 
n4942 , n4943 , n4944 , n4945 , n4946 , n4948 , n4949 , n4950 , n4951 , n4953 , 
n4954 , n4955 , n4956 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4965 , 
n4968 , n4969 , n4970 , n4971 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , 
n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , 
n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , 
n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , 
n5009 , n5010 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , 
n5021 , n5022 , n5023 , n5027 , n5028 , n5029 , n5030 , n5032 , n5033 , n5034 , 
n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , 
n5045 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , 
n5056 , n5057 , n5058 , n5059 , n5061 , n5063 , n5065 , n5066 , n5067 , n5068 , 
n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5078 , n5079 , 
n5080 , n5081 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5099 , n5100 , n5102 , 
n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , 
n5113 , n5114 , n5116 , n5117 , n5118 , n5119 , n5121 , n5122 , n5123 , n5124 , 
n5125 , n5126 , n5127 , n5129 , n5130 , n5132 , n5133 , n5134 , n5135 , n5136 , 
n5137 , n5138 , n5139 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , 
n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , 
n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5169 , 
n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , 
n5180 , n5181 , n5182 , n5183 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
n5212 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , 
n5223 , n5224 , n5225 , n5227 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , 
n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , 
n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , 
n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5266 , n5267 , 
n5268 , n5269 , n5270 , n5271 , n5272 , n5275 , n5276 , n5277 , n5278 , n5279 , 
n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , 
n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , 
n5301 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , 
n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , 
n5322 , n5323 , n5324 , n5326 , n5327 , n5328 , n5329 , n5331 , n5332 , n5333 , 
n5334 , n5335 , n5336 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , 
n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5352 , n5354 , n5355 , n5356 , 
n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , 
n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5377 , 
n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5387 , n5388 , 
n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , 
n5401 , n5402 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , 
n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , 
n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5431 , n5432 , 
n5433 , n5434 , n5435 , n5436 , n5437 , n5440 , n5441 , n5442 , n5444 , n5445 , 
n5446 , n5447 , n5448 , n5449 , n5450 , n5452 , n5453 , n5454 , n5455 , n5456 , 
n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , 
n5467 , n5468 , n5469 , n5470 , n5471 , n5473 , n5474 , n5475 , n5476 , n5477 , 
n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5486 , n5487 , n5488 , 
n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , 
n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , 
n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5518 , n5519 , 
n5520 , n5522 , n5523 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , 
n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , 
n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , 
n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , 
n5563 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , 
n5574 , n5575 , n5576 , n5577 , n5578 , n5580 , n5581 , n5582 , n5583 , n5584 , 
n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5594 , n5595 , 
n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5604 , n5606 , n5607 , 
n5608 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , 
n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , 
n5629 , n5630 , n5631 , n5632 , n5633 , n5635 , n5636 , n5637 , n5638 , n5639 , 
n5640 , n5641 , n5642 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , 
n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , 
n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , 
n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5681 , 
n5682 , n5683 , n5684 , n5685 , n5686 , n5688 , n5689 , n5690 , n5691 , n5692 , 
n5693 , n5694 , n5695 , n5697 , n5698 , n5699 , n5701 , n5702 , n5703 , n5705 , 
n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , 
n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , 
n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5733 , n5734 , n5735 , n5736 , 
n5737 , n5738 , n5739 , n5740 , n5741 , n5743 , n5744 , n5745 , n5746 , n5747 , 
n5748 , n5749 , n5750 , n5751 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , 
n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5766 , n5767 , n5768 , n5769 , 
n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5777 , n5778 , n5779 , n5780 , 
n5781 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , 
n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , 
n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , 
n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , 
n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , 
n5835 , n5836 , n5837 , n5838 , n5839 , n5843 , n5844 , n5845 , n5846 , n5847 , 
n5848 , n5849 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , 
n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , 
n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , 
n5879 , n5880 , n5881 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , 
n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , 
n5900 , n5901 , n5902 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5912 , 
n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , 
n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , 
n5933 , n5934 , n5935 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5944 , 
n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , 
n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5965 , 
n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , 
n5976 , n5977 , n5978 , n5979 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , 
n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , 
n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , 
n6007 , n6008 , n6009 , n6010 , n6011 , n6013 , n6014 , n6015 , n6016 , n6017 , 
n6018 , n6019 , n6020 , n6021 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , 
n6029 , n6030 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , 
n6040 , n6041 , n6042 , n6043 , n6045 , n6047 , n6048 , n6049 , n6050 , n6051 , 
n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , 
n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , 
n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , 
n6082 , n6083 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , 
n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , 
n6103 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , 
n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , 
n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , 
n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , 
n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , 
n6155 , n6156 , n6157 , n6158 , n6159 , n6161 , n6162 , n6163 , n6164 , n6165 , 
n6166 , n6167 , n6168 , n6169 , n6170 , n6172 , n6173 , n6174 , n6175 , n6176 , 
n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6184 , n6185 , n6186 , n6187 , 
n6188 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , 
n6199 , n6200 , n6201 , n6202 , n6203 , n6205 , n6206 , n6207 , n6208 , n6209 , 
n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6219 , n6220 , 
n6221 , n6222 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , 
n6232 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , 
n6243 , n6244 , n6246 , n6247 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , 
n6255 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , 
n6266 , n6267 , n6268 , n6269 , n6270 , n6272 , n6273 , n6274 , n6275 , n6277 , 
n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , 
n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , 
n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , 
n6309 , n6310 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , 
n6320 , n6321 , n6322 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6331 , 
n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6340 , n6341 , n6342 , 
n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , 
n6353 , n6355 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , 
n6365 , n6366 , n6367 , n6368 , n6370 , n6371 , n6372 , n6373 , n6374 , n6376 , 
n6377 , n6378 , n6380 , n6382 , n6384 , n6386 , n6387 , n6388 , n6389 , n6390 , 
n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6398 , n6399 , n6400 , n6401 , 
n6402 , n6403 , n6404 , n6405 , n6406 , n6408 , n6409 , n6410 , n6411 , n6412 , 
n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , 
n6423 , n6424 , n6425 , n6426 , n6428 , n6429 , n6430 , n6432 , n6433 , n6434 , 
n6435 , n6436 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , 
n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , 
n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6466 , n6467 , n6468 , 
n6469 , n6471 , n6472 , n6473 , n6474 , n6475 , n6477 , n6478 , n6479 , n6480 , 
n6481 , n6482 , n6483 , n6484 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , 
n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , 
n6503 , n6504 , n6505 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6515 , 
n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , 
n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , 
n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6543 , n6544 , n6545 , n6546 , 
n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6557 , 
n6559 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6568 , n6569 , n6570 , 
n6571 , n6572 , n6573 , n6574 , n6575 , n6577 , n6578 , n6579 , n6580 , n6581 , 
n6582 , n6583 , n6584 , n6585 , n6586 , n6588 , n6589 , n6591 , n6592 , n6593 , 
n6594 , n6595 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , 
n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6613 , n6614 , n6615 , n6616 , 
n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , 
n6627 , n6629 , n6632 , n6633 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , 
n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , 
n6651 , n6653 , n6654 , n6656 , n6657 , n6658 , n6660 , n6661 , n6662 , n6663 , 
n6664 , n6665 , n6666 , n6667 , n6668 , n6670 , n6672 , n6675 , n6676 , n6677 , 
n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6685 , n6686 , n6687 , n6688 , 
n6689 , n6690 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , 
n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6708 , n6709 , n6710 , n6711 , 
n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , 
n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6730 , n6731 , n6732 , 
n6733 , n6734 , n6735 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , 
n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , 
n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , 
n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6774 , 
n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6786 , 
n6787 , n6788 , n6789 , n6792 , n6793 , n6795 , n6796 , n6797 , n6798 , n6799 , 
n6800 , n6801 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , 
n6811 , n6812 , n6813 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , 
n6822 , n6823 , n6824 , n6825 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , 
n6833 , n6834 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , 
n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6854 , 
n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6864 , n6865 , n6866 , n6868 , 
n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , 
n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , 
n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , 
n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , 
n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , 
n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , 
n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , 
n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , 
n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , 
n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6966 , n6968 , n6969 , n6970 , 
n6972 , n6973 , n6974 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , 
n6984 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , 
n6995 , n6996 , n6997 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , 
n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , 
n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , 
n7027 , n7028 , n7029 , n7030 , n7031 , n7033 , n7034 , n7035 , n7036 , n7037 , 
n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , 
n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7058 , n7059 , 
n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , 
n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7080 , 
n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , 
n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7100 , n7101 , 
n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , 
n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , 
n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , 
n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7140 , n7141 , n7142 , 
n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7150 , n7151 , n7152 , n7153 , 
n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , 
n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , 
n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , 
n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7191 , n7192 , n7193 , n7194 , 
n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , 
n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , 
n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , 
n7225 , n7226 , n7227 , n7228 , n7231 , n7232 , n7234 , n7235 , n7237 , n7238 , 
n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , 
n7249 , n7250 , n7251 , n7252 , n7254 , n7255 , n7257 , n7258 , n7259 , n7260 , 
n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7269 , n7270 , n7271 , 
n7272 , n7273 , n7274 , n7275 , n7276 , n7278 , n7279 , n7281 , n7282 , n7283 , 
n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , 
n7294 , n7295 , n7296 , n7297 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , 
n7306 , n7307 , n7309 , n7310 , n7311 , n7312 , n7314 , n7315 , n7316 , n7317 , 
n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , 
n7328 , n7329 , n7331 , n7332 , n7333 , n7334 , n7336 , n7337 , n7338 , n7340 , 
n7341 , n7342 , n7343 , n7344 , n7345 , n7347 , n7348 , n7350 , n7351 , n7352 , 
n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , 
n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , 
n7374 , n7375 , n7376 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , 
n7385 , n7386 , n7387 , n7388 , n7389 , n7391 , n7392 , n7393 , n7394 , n7395 , 
n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7404 , n7405 , n7406 , 
n7407 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , 
n7418 , n7419 , n7420 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7429 , 
n7430 , n7431 , n7433 , n7434 , n7435 , n7436 , n7438 , n7439 , n7440 , n7441 , 
n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , 
n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7461 , n7462 , 
n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , 
n7473 , n7474 , n7476 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , 
n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , 
n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , 
n7505 , n7506 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7515 , n7516 , 
n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7525 , n7526 , n7527 , 
n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , 
n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , 
n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , 
n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7567 , n7568 , n7570 , 
n7571 , n7573 , n7574 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , 
n7583 , n7584 , n7586 , n7587 , n7589 , n7590 , n7591 , n7592 , n7594 , n7595 , 
n7596 , n7597 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , 
n7608 , n7609 , n7611 , n7612 , n7613 , n7614 , n7615 , n7617 , n7618 , n7619 , 
n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , 
n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , 
n7641 , n7642 , n7644 , n7645 , n7646 , n7648 , n7649 , n7650 , n7651 , n7652 , 
n7653 , n7654 , n7655 , n7656 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , 
n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7671 , n7672 , n7673 , n7675 , 
n7676 , n7677 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7687 , n7688 , 
n7689 , n7690 , n7691 , n7694 , n7695 , n7696 , n7697 , n7699 , n7700 , n7701 , 
n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7709 , n7710 , n7711 , n7712 , 
n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7722 , n7723 , 
n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7732 , n7733 , n7734 , 
n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , 
n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7752 , n7753 , n7754 , n7755 , 
n7756 , n7757 , n7758 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , 
n7767 , n7768 , n7770 , n7771 , n7772 , n7774 , n7775 , n7776 , n7777 , n7778 , 
n7779 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7789 , n7790 , 
n7791 , n7792 , n7793 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , 
n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7812 , 
n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , 
n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7831 , n7832 , n7833 , 
n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7842 , n7843 , n7844 , n7845 , 
n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , 
n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , 
n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , 
n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7885 , n7886 , n7887 , 
n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , 
n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , 
n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7918 , 
n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , 
n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7938 , n7939 , 
n7940 , n7941 , n7942 , n7944 , n7945 , n7946 , n7947 , n7948 , n7951 , n7952 , 
n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7960 , n7961 , n7962 , n7964 , 
n7965 , n7966 , n7967 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , 
n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , 
n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7993 , n7994 , n7995 , n7996 , 
n7997 , n7998 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8007 , n8008 , 
n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , 
n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8028 , n8029 , 
n8030 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , 
n8041 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , 
n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , 
n8063 , n8064 , n8065 , n8066 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , 
n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , 
n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , 
n8094 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8104 , n8105 , 
n8106 , n8107 , n8108 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , 
n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , 
n8128 , n8129 , n8131 , n8132 , n8133 , n8134 , n8136 , n8137 , n8138 , n8140 , 
n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8150 , n8151 , n8152 , 
n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8160 , n8161 , n8162 , n8163 , 
n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , 
n8174 , n8175 , n8176 , n8177 , n8178 , n8180 , n8181 , n8182 , n8183 , n8184 , 
n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8195 , 
n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , 
n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8216 , 
n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , 
n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , 
n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8245 , n8246 , n8247 , 
n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8257 , n8258 , n8260 , 
n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8268 , n8269 , n8270 , n8271 , 
n8272 , n8273 , n8274 , n8275 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , 
n8283 , n8284 , n8286 , n8287 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , 
n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , 
n8307 , n8308 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , 
n8318 , n8319 , n8322 , n8323 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , 
n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8340 , n8341 , 
n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , 
n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , 
n8362 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , 
n8373 , n8374 , n8375 , n8377 , n8378 , n8379 , n8380 , n8382 , n8383 , n8384 , 
n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , 
n8395 , n8396 , n8397 , n8398 , n8400 , n8401 , n8402 , n8403 , n8404 , n8406 , 
n8407 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8418 , 
n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , 
n8429 , n8430 , n8431 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8440 , 
n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , 
n8451 , n8452 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , 
n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , 
n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8481 , n8482 , 
n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8490 , n8491 , n8492 , n8493 , 
n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , 
n8504 , n8506 , n8507 , n8508 , n8509 , n8511 , n8512 , n8513 , n8514 , n8515 , 
n8516 , n8517 , n8518 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8527 , 
n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8536 , n8537 , n8538 , 
n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , 
n8549 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , 
n8560 , n8561 , n8562 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , 
n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , 
n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , 
n8592 , n8593 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , 
n8603 , n8604 , n8605 , n8606 , n8607 , n8609 , n8610 , n8611 , n8612 , n8613 , 
n8615 , n8616 , n8617 , n8618 , n8619 , n8621 , n8622 , n8623 , n8624 , n8625 , 
n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , 
n8636 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , 
n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8657 , n8658 , 
n8659 , n8660 , n8661 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , 
n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8679 , n8680 , 
n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8688 , n8689 , n8690 , n8691 , 
n8692 , n8693 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , 
n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , 
n8713 , n8714 , n8715 , n8717 , n8718 , n8719 , n8720 , n8722 , n8723 , n8724 , 
n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , 
n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8746 , 
n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , 
n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , 
n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , 
n8777 , n8778 , n8779 , n8780 , n8781 , n8783 , n8784 , n8785 , n8786 , n8787 , 
n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , 
n8798 , n8799 , n8800 , n8801 , n8802 , n8804 , n8805 , n8807 , n8808 , n8810 , 
n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , 
n8822 , n8823 , n8825 , n8826 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , 
n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , 
n8844 , n8845 , n8846 , n8847 , n8848 , n8850 , n8851 , n8852 , n8853 , n8854 , 
n8855 , n8857 , n8858 , n8859 , n8860 , n8863 , n8864 , n8865 , n8866 , n8867 , 
n8868 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , 
n8879 , n8880 , n8881 , n8882 , n8883 , n8885 , n8886 , n8887 , n8888 , n8889 , 
n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , 
n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8910 , 
n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8921 , n8922 , 
n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , 
n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , 
n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , 
n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , 
n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8972 , n8973 , n8974 , n8975 , 
n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8983 , n8984 , n8985 , n8986 , 
n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8994 , n8995 , n8996 , n8997 , 
n8998 , n8999 , n9000 , n9001 , n9002 , n9004 , n9005 , n9006 , n9007 , n9008 , 
n9009 , n9010 , n9011 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , 
n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , 
n9030 , n9031 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , 
n9041 , n9043 , n9044 , n9045 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , 
n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , 
n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , 
n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , 
n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9091 , n9092 , n9093 , n9094 , 
n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9105 , 
n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , 
n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , 
n9126 , n9127 , n9128 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , 
n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9147 , 
n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , 
n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9165 , n9167 , n9168 , n9169 , 
n9170 , n9171 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , 
n9181 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9192 , 
n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , 
n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , 
n9213 , n9214 , n9215 , n9216 , n9218 , n9219 , n9221 , n9222 , n9223 , n9224 , 
n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , 
n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , 
n9245 , n9247 , n9248 , n9249 , n9250 , n9252 , n9253 , n9254 , n9255 , n9256 , 
n9257 , n9258 , n9260 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , 
n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , 
n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9288 , n9289 , 
n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , 
n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9309 , n9310 , 
n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9319 , n9320 , n9321 , 
n9322 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , 
n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , 
n9343 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , 
n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , 
n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9373 , n9374 , n9375 , n9376 , 
n9377 , n9378 , n9379 , n9381 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , 
n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9397 , n9398 , n9400 , 
n9401 , n9402 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , 
n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9420 , n9421 , n9422 , 
n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9431 , n9432 , n9433 , n9434 , 
n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9446 , 
n9447 , n9448 , n9449 , n9450 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , 
n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , 
n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , 
n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , 
n9491 , n9492 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , 
n9502 , n9503 , n9504 , n9505 , n9506 , n9509 , n9510 , n9511 , n9513 , n9514 , 
n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , 
n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , 
n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , 
n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9553 , n9555 , n9559 , 
n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , 
n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , 
n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , 
n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9599 , n9600 , 
n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , 
n9611 , n9612 , n9613 , n9614 , n9615 , n9617 , n9618 , n9619 , n9620 , n9621 , 
n9623 , n9624 , n9625 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9634 , 
n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , 
n9647 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9656 , n9657 , n9658 , 
n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , 
n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , 
n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , 
n9690 , n9691 , n9692 , n9693 , n9694 , n9696 , n9697 , n9698 , n9700 , n9701 , 
n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , 
n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , 
n9722 , n9723 , n9724 , n9725 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , 
n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , 
n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , 
n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9762 , n9764 , n9765 , 
n9766 , n9768 , n9769 , n9770 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , 
n9779 , n9780 , n9781 , n9782 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , 
n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , 
n9800 , n9801 , n9802 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , 
n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , 
n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , 
n9831 , n9834 , n9835 , n9836 , n9837 , n9839 , n9840 , n9841 , n9842 , n9843 , 
n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , 
n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , 
n9864 , n9865 , n9866 , n9868 , n9869 , n9870 , n9871 , n9873 , n9874 , n9875 , 
n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , 
n9886 , n9887 , n9888 , n9889 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , 
n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , 
n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , 
n9918 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9927 , n9928 , n9929 , 
n9930 , n9931 , n9932 , n9933 , n9935 , n9936 , n9937 , n9939 , n9940 , n9941 , 
n9943 , n9944 , n9945 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , 
n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , 
n9964 , n9965 , n9966 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , 
n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , 
n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , 
n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , 
n10006 , n10007 , n10008 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10020 , 
n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , 
n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , 
n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , 
n10052 , n10054 , n10056 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , 
n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , 
n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , 
n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , 
n10095 , n10097 , n10098 , n10099 , n10100 , n10102 , n10103 , n10104 , n10105 , n10106 , 
n10107 , n10108 , n10109 , n10110 , n10112 , n10113 , n10114 , n10115 , n10116 , n10118 , 
n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10126 , n10127 , n10128 , n10129 , 
n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , 
n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , 
n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10159 , n10160 , 
n10161 , n10162 , n10163 , n10164 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , 
n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , 
n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , 
n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10202 , 
n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , 
n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , 
n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , 
n10233 , n10234 , n10235 , n10237 , n10238 , n10240 , n10241 , n10242 , n10243 , n10245 , 
n10246 , n10247 , n10248 , n10249 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , 
n10257 , n10258 , n10259 , n10260 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , 
n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10276 , n10277 , n10278 , n10279 , 
n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10288 , n10289 , n10290 , 
n10291 , n10292 , n10293 , n10294 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , 
n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , 
n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10322 , 
n10323 , n10324 , n10325 , n10328 , n10329 , n10331 , n10332 , n10333 , n10334 , n10335 , 
n10336 , n10337 , n10338 , n10339 , n10341 , n10342 , n10343 , n10344 , n10346 , n10347 , 
n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10357 , n10358 , 
n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , 
n10369 , n10370 , n10371 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , 
n10380 , n10381 , n10382 , n10383 , n10384 , n10386 , n10389 , n10391 , n10392 , n10393 , 
n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , 
n10406 , n10407 , n10408 , n10410 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , 
n10418 , n10419 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , 
n10429 , n10430 , n10431 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , 
n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , 
n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , 
n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , 
n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , 
n10480 , n10481 , n10482 , n10483 , n10485 , n10486 , n10487 , n10488 , n10490 , n10491 , 
n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , 
n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , 
n10512 , n10513 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , 
n10523 , n10524 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , 
n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10541 , n10542 , n10543 , n10544 , 
n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , 
n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10562 , n10563 , n10565 , n10566 , 
n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , 
n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , 
n10589 , n10590 , n10591 , n10592 , n10594 , n10596 , n10597 , n10598 , n10599 , n10600 , 
n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , 
n10612 , n10613 , n10615 , n10616 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , 
n10624 , n10625 , n10626 , n10627 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , 
n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , 
n10645 , n10646 , n10648 , n10649 , n10651 , n10652 , n10654 , n10655 , n10656 , n10657 , 
n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , 
n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , 
n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , 
n10688 , n10689 , n10690 , n10691 , n10693 , n10695 , n10696 , n10697 , n10698 , n10699 , 
n10700 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10711 , 
n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , 
n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , 
n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10740 , n10741 , n10742 , n10743 , 
n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , 
n10754 , n10755 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10764 , n10765 , 
n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10776 , 
n10777 , n10778 , n10779 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , 
n10788 , n10789 , n10790 , n10791 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , 
n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , 
n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10818 , n10819 , 
n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , 
n10830 , n10831 , n10832 , n10833 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , 
n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , 
n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , 
n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , 
n10872 , n10873 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , 
n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , 
n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , 
n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , 
n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , 
n10923 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , 
n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10944 , 
n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , 
n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10962 , n10963 , n10964 , n10965 , 
n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , 
n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , 
n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , 
n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11006 , 
n11007 , n11008 , n11009 , n11010 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , 
n11018 , n11019 , n11020 , n11021 , n11022 , n11024 , n11026 , n11027 , n11028 , n11029 , 
n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , 
n11040 , n11041 , n11042 , n11043 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , 
n11051 , n11052 , n11053 , n11054 , n11055 , n11057 , n11058 , n11059 , n11060 , n11061 , 
n11062 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , 
n11073 , n11074 , n11075 , n11076 , n11077 , n11079 , n11081 , n11082 , n11083 , n11084 , 
n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11095 , 
n11096 , n11097 , n11098 , n11099 , n11100 , n11102 , n11104 , n11105 , n11106 , n11107 , 
n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , 
n11118 , n11119 , n11122 , n11123 , n11124 , n11125 , n11126 , n11128 , n11129 , n11130 , 
n11131 , n11133 , n11135 , n11136 , n11137 , n11139 , n11140 , n11141 , n11142 , n11143 , 
n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , 
n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , 
n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , 
n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11183 , n11185 , 
n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11193 , n11194 , n11195 , n11196 , 
n11197 , n11198 , n11199 , n11200 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , 
n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , 
n11218 , n11219 , n11221 , n11222 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , 
n11230 , n11231 , n11232 , n11233 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , 
n11241 , n11242 , n11243 , n11244 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , 
n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11262 , 
n11263 , n11264 , n11265 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11274 , 
n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , 
n11286 , n11287 , n11288 , n11289 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , 
n11297 , n11298 , n11299 , n11300 , n11301 , n11303 , n11304 , n11305 , n11306 , n11307 , 
n11308 , n11309 , n11310 , n11311 , n11312 , n11314 , n11315 , n11316 , n11317 , n11318 , 
n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11327 , n11328 , n11329 , n11331 , 
n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , 
n11342 , n11343 , n11344 , n11345 , n11346 , n11349 , n11350 , n11351 , n11353 , n11354 , 
n11355 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , 
n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11376 , 
n11377 , n11378 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11387 , n11388 , 
n11389 , n11390 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11399 , n11400 , 
n11401 , n11402 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , 
n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11420 , n11421 , n11422 , 
n11423 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , 
n11434 , n11435 , n11436 , n11437 , n11438 , n11440 , n11441 , n11442 , n11443 , n11444 , 
n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , 
n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11463 , n11464 , n11465 , n11466 , 
n11467 , n11468 , n11469 , n11471 , n11474 , n11475 , n11476 , n11477 , n11478 , n11480 , 
n11482 , n11483 , n11484 , n11485 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , 
n11493 , n11494 , n11495 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11504 , 
n11505 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11516 , 
n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , 
n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , 
n11537 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , 
n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , 
n11559 , n11560 , n11561 , n11562 , n11563 , n11565 , n11567 , n11568 , n11569 , n11570 , 
n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11581 , n11582 , 
n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11592 , n11593 , 
n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , 
n11604 , n11605 , n11606 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , 
n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , 
n11626 , n11627 , n11628 , n11629 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , 
n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , 
n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , 
n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11668 , 
n11669 , n11670 , n11671 , n11672 , n11673 , n11675 , n11676 , n11677 , n11678 , n11679 , 
n11680 , n11681 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , 
n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , 
n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11711 , 
n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , 
n11723 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , 
n11734 , n11735 , n11737 , n11738 , n11739 , n11740 , n11742 , n11743 , n11744 , n11745 , 
n11746 , n11747 , n11748 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , 
n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , 
n11767 , n11768 , n11769 , n11772 , n11773 , n11774 , n11776 , n11777 , n11778 , n11779 , 
n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , 
n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , 
n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , 
n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11819 , n11820 , 
n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , 
n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11838 , n11839 , n11840 , n11844 , 
n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , 
n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , 
n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , 
n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , 
n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , 
n11895 , n11896 , n11897 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11906 , 
n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , 
n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11927 , 
n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , 
n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , 
n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , 
n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11966 , n11967 , n11968 , 
n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , 
n11979 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , 
n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , 
n12001 , n12002 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12012 , 
n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , 
n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , 
n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , 
n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , 
n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , 
n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12073 , 
n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , 
n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , 
n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , 
n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12114 , 
n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12122 , n12123 , n12124 , n12125 , 
n12126 , n12127 , n12128 , n12129 , n12130 , n12132 , n12133 , n12134 , n12135 , n12136 , 
n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12147 , 
n12148 , n12149 , n12150 , n12151 , n12154 , n12155 , n12156 , n12159 , n12160 , n12162 , 
n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , 
n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12180 , n12181 , n12182 , n12183 , 
n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12193 , n12194 , 
n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , 
n12205 , n12206 , n12207 , n12208 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , 
n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12224 , n12226 , n12227 , 
n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12236 , n12237 , n12238 , n12239 , 
n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , 
n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , 
n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , 
n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , 
n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , 
n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , 
n12300 , n12301 , n12303 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , 
n12312 , n12313 , n12314 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , 
n12323 , n12326 , n12327 , n12328 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , 
n12337 , n12338 , n12339 , n12340 , n12342 , n12343 , n12344 , n12345 , n12347 , n12348 , 
n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , 
n12360 , n12361 , n12362 , n12363 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , 
n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12381 , 
n12382 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , 
n12394 , n12395 , n12396 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , 
n12406 , n12407 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , 
n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , 
n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , 
n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12447 , 
n12448 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , 
n12459 , n12460 , n12463 , n12464 , n12465 , n12466 , n12468 , n12470 , n12471 , n12472 , 
n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , 
n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , 
n12493 , n12494 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , 
n12504 , n12505 , n12506 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , 
n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , 
n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , 
n12537 , n12538 , n12539 , n12541 , n12542 , n12543 , n12544 , n12547 , n12548 , n12549 , 
n12550 , n12551 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , 
n12561 , n12563 , n12564 , n12565 , n12567 , n12568 , n12570 , n12571 , n12572 , n12573 , 
n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , 
n12584 , n12585 , n12586 , n12588 , n12589 , n12590 , n12591 , n12592 , n12594 , n12595 , 
n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , 
n12606 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , 
n12617 , n12618 , n12619 , n12622 , n12623 , n12624 , n12625 , n12627 , n12628 , n12629 , 
n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , 
n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , 
n12651 , n12652 , n12653 , n12655 , n12656 , n12658 , n12659 , n12660 , n12661 , n12662 , 
n12663 , n12664 , n12666 , n12667 , n12668 , n12669 , n12671 , n12672 , n12673 , n12674 , 
n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , 
n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , 
n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12703 , n12704 , n12705 , 
n12706 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , 
n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12726 , n12728 , 
n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , 
n12739 , n12741 , n12743 , n12744 , n12745 , n12747 , n12748 , n12749 , n12750 , n12751 , 
n12752 , n12753 , n12754 , n12755 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , 
n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , 
n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , 
n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , 
n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12802 , n12803 , n12804 , 
n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12813 , n12814 , n12815 , n12817 , 
n12818 , n12819 , n12820 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , 
n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , 
n12839 , n12840 , n12841 , n12842 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , 
n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , 
n12860 , n12862 , n12863 , n12866 , n12867 , n12868 , n12869 , n12872 , n12874 , n12876 , 
n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , 
n12887 , n12888 , n12889 , n12890 , n12891 , n12893 , n12894 , n12895 , n12896 , n12897 , 
n12898 , n12899 , n12901 , n12902 , n12903 , n12905 , n12906 , n12907 , n12908 , n12909 , 
n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12918 , n12919 , n12920 , 
n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , 
n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , 
n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , 
n12953 , n12954 , n12955 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , 
n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , 
n12974 , n12975 , n12976 , n12977 , n12979 , n12981 , n12982 , n12983 , n12984 , n12986 , 
n12988 , n12989 , n12990 , n12991 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , 
n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13006 , n13007 , n13008 , n13009 , 
n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , 
n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13027 , n13028 , n13029 , n13030 , 
n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , 
n13041 , n13042 , n13045 , n13046 , n13047 , n13049 , n13050 , n13051 , n13052 , n13053 , 
n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , 
n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13075 , 
n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13083 , n13084 , n13085 , n13086 , 
n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13097 , 
n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , 
n13108 , n13109 , n13111 , n13112 , n13113 , n13114 , n13115 , n13117 , n13118 , n13119 , 
n13120 , n13121 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , 
n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13138 , n13139 , n13140 , n13142 , 
n13143 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , 
n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , 
n13164 , n13165 , n13166 , n13167 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , 
n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , 
n13185 , n13186 , n13187 , n13188 , n13189 , n13191 , n13192 , n13193 , n13194 , n13195 , 
n13196 , n13197 , n13200 , n13201 , n13202 , n13203 , n13205 , n13206 , n13207 , n13208 , 
n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , 
n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , 
n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , 
n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , 
n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , 
n13260 , n13261 , n13262 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13271 , 
n13272 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , 
n13283 , n13284 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , 
n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , 
n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , 
n13314 , n13315 , n13316 , n13317 , n13318 , n13320 , n13321 , n13322 , n13323 , n13324 , 
n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13334 , n13335 , 
n13336 , n13337 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , 
n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , 
n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , 
n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , 
n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , 
n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , 
n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13408 , 
n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13420 , 
n13421 , n13422 , n13423 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , 
n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , 
n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , 
n13452 , n13454 , n13455 , n13458 , n13459 , n13461 , n13462 , n13463 , n13464 , n13465 , 
n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , 
n13476 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13485 , n13488 , n13489 , 
n13491 , n13492 , n13493 , n13495 , n13496 , n13497 , n13498 , n13499 , n13502 , n13503 , 
n13504 , n13505 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , 
n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , 
n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , 
n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , 
n13545 , n13546 , n13547 , n13550 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , 
n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , 
n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , 
n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , 
n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , 
n13598 , n13599 , n13600 , n13601 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , 
n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , 
n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13627 , n13628 , n13629 , 
n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , 
n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , 
n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , 
n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13669 , n13670 , 
n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13678 , n13679 , n13680 , n13681 , 
n13682 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , 
n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , 
n13703 , n13704 , n13705 , n13706 , n13707 , n13709 , n13711 , n13712 , n13713 , n13715 , 
n13716 , n13717 , n13718 , n13720 , n13721 , n13723 , n13724 , n13725 , n13726 , n13727 , 
n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , 
n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , 
n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13755 , n13756 , n13757 , n13758 , 
n13759 , n13760 , n13761 , n13762 , n13763 , n13765 , n13766 , n13767 , n13768 , n13769 , 
n13770 , n13771 , n13772 , n13773 , n13774 , n13776 , n13777 , n13778 , n13779 , n13780 , 
n13782 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , 
n13793 , n13794 , n13795 , n13796 , n13797 , n13799 , n13800 , n13801 , n13802 , n13803 , 
n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , 
n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , 
n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , 
n13834 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , 
n13845 , n13846 , n13847 , n13848 , n13849 , n13852 , n13853 , n13854 , n13855 , n13856 , 
n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , 
n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , 
n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , 
n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , 
n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , 
n13907 , n13908 , n13909 , n13910 , n13911 , n13913 , n13915 , n13916 , n13917 , n13918 , 
n13919 , n13920 , n13921 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , 
n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , 
n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , 
n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , 
n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , 
n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , 
n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , 
n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , 
n14002 , n14003 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , 
n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , 
n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , 
n14033 , n14034 , n14035 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , 
n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , 
n14054 , n14055 , n14056 , n14057 , n14058 , n14060 , n14061 , n14062 , n14063 , n14064 , 
n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14072 , n14073 , n14074 , n14075 , 
n14076 , n14077 , n14078 , n14079 , n14080 , n14082 , n14083 , n14084 , n14085 , n14086 , 
n14087 , n14088 , n14089 , n14091 , n14092 , n14093 , n14094 , n14096 , n14097 , n14098 , 
n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14108 , n14109 , 
n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , 
n14120 , n14122 , n14123 , n14124 , n14125 , n14127 , n14128 , n14129 , n14131 , n14132 , 
n14133 , n14134 , n14135 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , 
n14144 , n14145 , n14146 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , 
n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , 
n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14175 , n14176 , 
n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , 
n14187 , n14188 , n14189 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , 
n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , 
n14208 , n14209 , n14210 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , 
n14219 , n14220 , n14221 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , 
n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , 
n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , 
n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , 
n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14268 , n14269 , n14270 , n14272 , 
n14273 , n14274 , n14276 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , 
n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14295 , 
n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , 
n14306 , n14307 , n14308 , n14309 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , 
n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14324 , n14325 , n14327 , n14328 , 
n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , 
n14339 , n14340 , n14341 , n14343 , n14344 , n14346 , n14347 , n14348 , n14349 , n14350 , 
n14351 , n14352 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , 
n14362 , n14363 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , 
n14373 , n14374 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , 
n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , 
n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , 
n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14413 , n14415 , 
n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , 
n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , 
n14436 , n14437 , n14438 , n14439 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , 
n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , 
n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14465 , n14466 , n14467 , n14468 , 
n14469 , n14470 , n14472 , n14473 , n14474 , n14476 , n14477 , n14478 , n14479 , n14480 , 
n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , 
n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , 
n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14511 , 
n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , 
n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , 
n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14542 , 
n14543 , n14544 , n14545 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , 
n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , 
n14565 , n14566 , n14567 , n14568 , n14569 , n14571 , n14572 , n14573 , n14574 , n14577 , 
n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , 
n14588 , n14589 , n14590 , n14591 , n14592 , n14594 , n14595 , n14596 , n14597 , n14598 , 
n14599 , n14600 , n14601 , n14602 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , 
n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , 
n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , 
n14630 , n14631 , n14632 , n14634 , n14635 , n14637 , n14638 , n14639 , n14640 , n14641 , 
n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , 
n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , 
n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , 
n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14681 , n14682 , 
n14683 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14693 , n14694 , 
n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14703 , n14705 , n14706 , n14707 , 
n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , 
n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , 
n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14735 , n14736 , n14737 , n14738 , 
n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14747 , n14748 , n14749 , 
n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , 
n14760 , n14761 , n14762 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , 
n14771 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , 
n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14791 , n14792 , 
n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14802 , n14803 , 
n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , 
n14814 , n14815 , n14816 , n14817 , n14818 , n14820 , n14821 , n14822 , n14823 , n14824 , 
n14825 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , 
n14837 , n14838 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , 
n14848 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , 
n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , 
n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , 
n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , 
n14889 , n14890 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14900 , 
n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , 
n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , 
n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , 
n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , 
n14942 , n14943 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , 
n14953 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , 
n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , 
n14974 , n14975 , n14976 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , 
n14985 , n14986 , n14987 , n14988 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , 
n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15003 , n15005 , n15006 , n15007 , 
n15008 , n15009 , n15010 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , 
n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , 
n15030 , n15032 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , 
n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , 
n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , 
n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , 
n15074 , n15075 , n15076 , n15078 , n15079 , n15080 , n15081 , n15083 , n15084 , n15085 , 
n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15095 , n15096 , 
n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , 
n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , 
n15117 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , 
n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , 
n15140 , n15141 , n15142 , n15143 , n15144 , n15147 , n15148 , n15149 , n15150 , n15151 , 
n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , 
n15162 , n15163 , n15164 , n15166 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , 
n15174 , n15175 , n15177 , n15178 , n15179 , n15181 , n15183 , n15184 , n15185 , n15186 , 
n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , 
n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15206 , n15207 , 
n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , 
n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , 
n15228 , n15229 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , 
n15239 , n15240 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , 
n15250 , n15251 , n15252 , n15253 , n15254 , n15256 , n15257 , n15259 , n15260 , n15261 , 
n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15272 , 
n15273 , n15274 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , 
n15284 , n15285 , n15286 , n15287 , n15288 , n15290 , n15291 , n15292 , n15293 , n15294 , 
n15295 , n15296 , n15297 , n15298 , n15299 , n15301 , n15302 , n15303 , n15304 , n15305 , 
n15306 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , 
n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , 
n15328 , n15329 , n15330 , n15331 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , 
n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15346 , n15347 , n15348 , n15349 , 
n15350 , n15351 , n15352 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , 
n15361 , n15362 , n15363 , n15364 , n15365 , n15367 , n15368 , n15369 , n15370 , n15371 , 
n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15379 , n15380 , n15381 , n15383 , 
n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , 
n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , 
n15404 , n15405 , n15406 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , 
n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15425 , 
n15426 , n15427 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15436 , n15437 , 
n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , 
n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , 
n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15466 , n15468 , n15469 , n15471 , 
n15472 , n15473 , n15474 , n15475 , n15476 , n15478 , n15479 , n15480 , n15482 , n15483 , 
n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15491 , n15492 , n15493 , n15494 , 
n15495 , n15497 , n15498 , n15499 , n15500 , n15502 , n15503 , n15504 , n15505 , n15507 , 
n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , 
n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , 
n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , 
n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15547 , n15548 , n15549 , n15550 , 
n15551 , n15552 , n15553 , n15554 , n15556 , n15557 , n15560 , n15561 , n15562 , n15563 , 
n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15571 , n15572 , n15574 , n15575 , 
n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , 
n15586 , n15587 , n15589 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , 
n15599 , n15600 , n15601 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , 
n15610 , n15611 , n15612 , n15613 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , 
n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , 
n15631 , n15632 , n15633 , n15634 , n15635 , n15637 , n15638 , n15639 , n15640 , n15641 , 
n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , 
n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15663 , 
n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , 
n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , 
n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , 
n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , 
n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , 
n15714 , n15715 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , 
n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , 
n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15744 , n15745 , 
n15746 , n15747 , n15748 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , 
n15757 , n15758 , n15759 , n15760 , n15763 , n15764 , n15765 , n15767 , n15768 , n15769 , 
n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , 
n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , 
n15791 , n15792 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , 
n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , 
n15813 , n15814 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , 
n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15832 , n15833 , n15834 , n15835 , 
n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , 
n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , 
n15857 , n15858 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , 
n15868 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , 
n15879 , n15880 , n15881 , n15882 , n15883 , n15886 , n15887 , n15888 , n15890 , n15891 , 
n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , 
n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , 
n15912 , n15913 , n15914 , n15915 , n15916 , n15919 , n15920 , n15921 , n15923 , n15924 , 
n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , 
n15935 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , 
n15946 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15957 , 
n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15968 , n15969 , 
n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15980 , 
n15981 , n15982 , n15983 , n15984 , n15985 , n15987 , n15988 , n15989 , n15990 , n15991 , 
n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , 
n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , 
n16012 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , 
n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16030 , n16031 , n16032 , n16033 , 
n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , 
n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , 
n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16061 , n16063 , n16064 , n16065 , 
n16066 , n16067 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , 
n16077 , n16078 , n16079 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , 
n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , 
n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , 
n16109 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , 
n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , 
n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , 
n16140 , n16141 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , 
n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16159 , n16160 , n16161 , 
n16162 , n16163 , n16164 , n16165 , n16166 , n16168 , n16169 , n16170 , n16171 , n16172 , 
n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , 
n16183 , n16184 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , 
n16194 , n16195 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , 
n16205 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16216 , 
n16220 , n16221 , n16222 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16231 , 
n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , 
n16242 , n16244 , n16245 , n16246 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , 
n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , 
n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , 
n16274 , n16276 , n16277 , n16278 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , 
n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , 
n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , 
n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , 
n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16323 , n16324 , n16325 , n16326 , 
n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , 
n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , 
n16348 , n16349 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , 
n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16368 , n16369 , 
n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16377 , n16378 , n16380 , n16381 , 
n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , 
n16392 , n16393 , n16394 , n16395 , n16397 , n16399 , n16400 , n16401 , n16402 , n16403 , 
n16404 , n16405 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , 
n16416 , n16417 , n16418 , n16420 , n16421 , n16422 , n16423 , n16425 , n16426 , n16427 , 
n16429 , n16430 , n16431 , n16432 , n16434 , n16435 , n16436 , n16437 , n16438 , n16441 , 
n16442 , n16443 , n16444 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , 
n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16461 , n16462 , n16463 , 
n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , 
n16474 , n16475 , n16477 , n16478 , n16479 , n16480 , n16483 , n16484 , n16485 , n16486 , 
n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16494 , n16495 , n16496 , n16497 , 
n16498 , n16499 , n16500 , n16501 , n16503 , n16504 , n16505 , n16508 , n16509 , n16510 , 
n16511 , n16512 , n16513 , n16514 , n16515 , n16518 , n16519 , n16520 , n16522 , n16523 , 
n16525 , n16526 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , 
n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16545 , n16546 , 
n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16555 , n16556 , n16557 , 
n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , 
n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , 
n16578 , n16579 , n16580 , n16581 , n16582 , n16585 , n16586 , n16587 , n16588 , n16590 , 
n16591 , n16592 , n16593 , n16594 , n16595 , n16597 , n16598 , n16599 , n16600 , n16601 , 
n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16609 , n16610 , n16611 , n16612 , 
n16613 , n16614 , n16615 , n16616 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , 
n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16631 , n16632 , n16633 , n16634 , 
n16635 , n16636 , n16637 , n16638 , n16639 , n16641 , n16642 , n16643 , n16644 , n16645 , 
n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , 
n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , 
n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16675 , n16676 , n16677 , 
n16678 , n16679 , n16680 , n16681 , n16683 , n16685 , n16686 , n16687 , n16689 , n16690 , 
n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , 
n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , 
n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , 
n16721 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , 
n16732 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , 
n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , 
n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , 
n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , 
n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , 
n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , 
n16794 , n16795 , n16796 , n16797 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , 
n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16813 , n16814 , n16815 , 
n16816 , n16817 , n16819 , n16820 , n16821 , n16822 , n16823 , n16825 , n16826 , n16827 , 
n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16835 , n16836 , n16838 , n16839 , 
n16840 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , 
n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , 
n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , 
n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , 
n16881 , n16882 , n16883 , n16884 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , 
n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , 
n16902 , n16903 , n16904 , n16906 , n16907 , n16908 , n16909 , n16910 , n16912 , n16913 , 
n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , 
n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , 
n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , 
n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16952 , n16953 , n16955 , 
n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , 
n16966 , n16967 , n16969 , n16970 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , 
n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , 
n16990 , n16991 , n16992 , n16993 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , 
n17001 , n17002 , n17003 , n17004 , n17005 , n17007 , n17008 , n17009 , n17010 , n17011 , 
n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , 
n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , 
n17032 , n17033 , n17034 , n17036 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , 
n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , 
n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , 
n17064 , n17065 , n17066 , n17067 , n17071 , n17072 , n17073 , n17074 , n17076 , n17078 , 
n17079 , n17080 , n17081 , n17082 , n17083 , n17085 , n17086 , n17087 , n17088 , n17089 , 
n17091 , n17092 , n17093 , n17094 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , 
n17102 , n17103 , n17105 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , 
n17114 , n17115 , n17116 , n17117 , n17118 , n17120 , n17121 , n17122 , n17123 , n17124 , 
n17125 , n17126 , n17127 , n17128 , n17129 , n17131 , n17132 , n17133 , n17134 , n17135 , 
n17136 , n17137 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , 
n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , 
n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17164 , n17165 , n17166 , n17167 , 
n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , 
n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , 
n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , 
n17199 , n17200 , n17201 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , 
n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17220 , 
n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , 
n17231 , n17233 , n17234 , n17235 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , 
n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17252 , n17253 , n17254 , n17255 , 
n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17264 , n17265 , n17266 , 
n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , 
n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17286 , n17287 , 
n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , 
n17298 , n17299 , n17300 , n17301 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , 
n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , 
n17319 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , 
n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17338 , n17339 , n17340 , 
n17341 , n17342 , n17343 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17352 , 
n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17360 , n17361 , n17362 , n17363 , 
n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , 
n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , 
n17384 , n17385 , n17386 , n17388 , n17389 , n17390 , n17393 , n17394 , n17395 , n17396 , 
n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , 
n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , 
n17417 , n17418 , n17419 , n17420 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , 
n17428 , n17429 , n17430 , n17431 , n17433 , n17434 , n17435 , n17437 , n17438 , n17439 , 
n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17451 , 
n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17459 , n17460 , n17462 , n17463 , 
n17464 , n17465 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , 
n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , 
n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17494 , n17495 , 
n17496 , n17497 , n17498 , n17499 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , 
n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , 
n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17525 , n17526 , n17527 , 
n17528 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , 
n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , 
n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17558 , n17559 , 
n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , 
n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , 
n17580 , n17581 , n17582 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , 
n17591 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , 
n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , 
n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , 
n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , 
n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17639 , n17640 , n17641 , n17642 , 
n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , 
n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , 
n17663 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , 
n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , 
n17684 , n17685 , n17686 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , 
n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , 
n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , 
n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17722 , n17723 , n17724 , n17725 , 
n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17736 , 
n17737 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17747 , n17748 , 
n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , 
n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , 
n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , 
n17780 , n17781 , n17782 , n17783 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , 
n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , 
n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , 
n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17821 , 
n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , 
n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , 
n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , 
n17852 , n17853 , n17854 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , 
n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , 
n17873 , n17874 , n17875 , n17876 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , 
n17884 , n17885 , n17886 , n17887 , n17888 , n17890 , n17891 , n17892 , n17893 , n17894 , 
n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , 
n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17913 , n17914 , n17915 , n17916 , 
n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , 
n17928 , n17929 , n17930 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , 
n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17949 , 
n17950 , n17951 , n17952 , n17953 , n17955 , n17957 , n17958 , n17960 , n17961 , n17962 , 
n17964 , n17965 , n17966 , n17967 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , 
n17975 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , 
n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , 
n17996 , n17997 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , 
n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , 
n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18026 , n18027 , 
n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18036 , n18037 , n18038 , 
n18039 , n18040 , n18041 , n18042 , n18044 , n18046 , n18047 , n18048 , n18049 , n18050 , 
n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18060 , n18062 , 
n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18072 , n18073 , 
n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , 
n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , 
n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , 
n18104 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , 
n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , 
n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , 
n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18144 , n18146 , 
n18147 , n18148 , n18149 , n18150 , n18153 , n18154 , n18155 , n18156 , n18158 , n18159 , 
n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , 
n18170 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , 
n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , 
n18191 , n18192 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , 
n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , 
n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , 
n18222 , n18223 , n18224 , n18225 , n18226 , n18228 , n18229 , n18230 , n18231 , n18233 , 
n18234 , n18235 , n18236 , n18237 , n18239 , n18240 , n18242 , n18243 , n18244 , n18245 , 
n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18255 , n18256 , 
n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , 
n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18275 , n18276 , n18277 , 
n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , 
n18289 , n18291 , n18292 , n18293 , n18294 , n18296 , n18297 , n18298 , n18299 , n18300 , 
n18302 , n18303 , n18305 , n18306 , n18307 , n18308 , n18309 , n18312 , n18313 , n18314 , 
n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18324 , n18325 , 
n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18333 , n18334 , n18335 , n18336 , 
n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18344 , n18346 , n18347 , n18348 , 
n18349 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , 
n18360 , n18361 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , 
n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18378 , n18379 , n18380 , n18381 , 
n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , 
n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , 
n18402 , n18403 , n18404 , n18406 , n18407 , n18408 , n18410 , n18411 , n18412 , n18413 , 
n18415 , n18416 , n18417 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , 
n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , 
n18436 , n18438 , n18440 , n18441 , n18442 , n18443 , n18446 , n18447 , n18448 , n18449 , 
n18450 , n18451 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , 
n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18468 , n18469 , n18470 , n18471 , 
n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , 
n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , 
n18494 , n18495 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , 
n18505 , n18506 , n18507 , n18508 , n18510 , n18511 , n18512 , n18514 , n18516 , n18517 , 
n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , 
n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18538 , 
n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , 
n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18559 , 
n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , 
n18570 , n18571 , n18573 , n18575 , n18577 , n18579 , n18580 , n18581 , n18585 , n18586 , 
n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , 
n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , 
n18607 , n18608 , n18609 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , 
n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , 
n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18636 , n18637 , n18638 , 
n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , 
n18650 , n18651 , n18652 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , 
n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , 
n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18680 , n18681 , 
n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18691 , n18692 , 
n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , 
n18704 , n18705 , n18706 , n18707 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , 
n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18722 , n18723 , n18724 , n18726 , 
n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , 
n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18746 , n18747 , n18748 , 
n18749 , n18750 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , 
n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , 
n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , 
n18781 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , 
n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , 
n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , 
n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , 
n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18832 , n18833 , n18834 , 
n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18844 , n18845 , 
n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , 
n18856 , n18857 , n18860 , n18861 , n18862 , n18863 , n18866 , n18867 , n18868 , n18869 , 
n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , 
n18881 , n18882 , n18883 , n18884 , n18885 , n18888 , n18889 , n18890 , n18891 , n18892 , 
n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18902 , n18903 , 
n18904 , n18905 , n18906 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , 
n18915 , n18916 , n18917 , n18918 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , 
n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , 
n18937 , n18938 , n18939 , n18941 , n18942 , n18943 , n18944 , n18946 , n18947 , n18948 , 
n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , 
n18959 , n18960 , n18961 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , 
n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18978 , n18979 , n18980 , n18981 , 
n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , 
n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n19000 , n19001 , n19002 , n19003 , 
n19004 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , 
n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , 
n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19034 , n19035 , 
n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19043 , n19045 , n19046 , n19047 , 
n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , 
n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , 
n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , 
n19078 , n19079 , n19080 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , 
n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , 
n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19108 , n19109 , 
n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19117 , n19118 , n19119 , n19120 , 
n19121 , n19122 , n19123 , n19124 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , 
n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19142 , 
n19143 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , 
n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19165 , 
n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19175 , n19177 , 
n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , 
n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19197 , n19198 , 
n19199 , n19200 , n19201 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , 
n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , 
n19222 , n19225 , n19226 , n19227 , n19229 , n19230 , n19231 , n19232 , n19235 , n19236 , 
n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19245 , n19246 , n19247 , 
n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , 
n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , 
n19268 , n19269 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , 
n19279 , n19280 , n19281 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , 
n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , 
n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , 
n19310 , n19311 , n19312 , n19313 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , 
n19322 , n19324 , n19325 , n19326 , n19328 , n19329 , n19330 , n19331 , n19332 , n19334 , 
n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , 
n19345 , n19346 , n19347 , n19349 , n19350 , n19351 , n19352 , n19353 , n19355 , n19356 , 
n19358 , n19359 , n19360 , n19362 , n19363 , n19364 , n19365 , n19366 , n19368 , n19369 , 
n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , 
n19380 , n19381 , n19382 , n19383 , n19384 , n19386 , n19387 , n19388 , n19390 , n19391 , 
n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19402 , 
n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , 
n19413 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , 
n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , 
n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , 
n19445 , n19446 , n19447 , n19448 , n19449 , n19451 , n19452 , n19453 , n19455 , n19456 , 
n19457 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19468 , 
n19469 , n19470 , n19471 , n19473 , n19474 , n19475 , n19476 , n19478 , n19479 , n19480 , 
n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , 
n19491 , n19492 , n19493 , n19495 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , 
n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , 
n19513 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19524 , n19525 , 
n19526 , n19527 , n19528 , n19529 , n19530 , n19532 , n19533 , n19534 , n19535 , n19536 , 
n19537 , n19538 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , 
n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , 
n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , 
n19568 , n19569 , n19571 , n19572 , n19573 , n19574 , n19576 , n19577 , n19578 , n19579 , 
n19580 , n19581 , n19582 , n19583 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , 
n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , 
n19601 , n19603 , n19604 , n19605 , n19606 , n19607 , n19609 , n19610 , n19611 , n19612 , 
n19613 , n19614 , n19615 , n19616 , n19619 , n19620 , n19621 , n19622 , n19624 , n19625 , 
n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , 
n19636 , n19637 , n19638 , n19639 , n19640 , n19642 , n19643 , n19644 , n19645 , n19646 , 
n19647 , n19649 , n19650 , n19651 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , 
n19659 , n19660 , n19661 , n19662 , n19663 , n19665 , n19666 , n19667 , n19668 , n19669 , 
n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , 
n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , 
n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , 
n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , 
n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , 
n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , 
n19732 , n19733 , n19734 , n19735 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , 
n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19750 , n19751 , n19752 , n19753 , 
n19754 , n19755 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , 
n19765 , n19766 , n19768 , n19769 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , 
n19777 , n19778 , n19779 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , 
n19788 , n19790 , n19791 , n19793 , n19794 , n19795 , n19796 , n19797 , n19799 , n19800 , 
n19801 , n19802 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , 
n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , 
n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , 
n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , 
n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , 
n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , 
n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , 
n19872 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , 
n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , 
n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , 
n19903 , n19904 , n19906 , n19907 , n19908 , n19910 , n19912 , n19913 , n19914 , n19915 , 
n19917 , n19918 , n19919 , n19920 , n19921 , n19924 , n19925 , n19926 , n19927 , n19928 , 
n19929 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , 
n19940 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , 
n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , 
n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19969 , n19970 , n19971 , 
n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , 
n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19989 , n19990 , n19991 , n19992 , 
n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , 
n20003 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20014 , 
n20015 , n20016 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , 
n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20034 , n20035 , n20037 , 
n20038 , n20039 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , 
n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , 
n20059 , n20060 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20070 , 
n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20078 , n20079 , n20080 , n20081 , 
n20082 , n20083 , n20084 , n20085 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , 
n20093 , n20094 , n20095 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20104 , 
n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , 
n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , 
n20125 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , 
n20136 , n20137 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , 
n20147 , n20148 , n20150 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , 
n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , 
n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20180 , 
n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20188 , n20189 , n20190 , n20191 , 
n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , 
n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , 
n20212 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , 
n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , 
n20233 , n20234 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , 
n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20251 , n20252 , n20253 , n20254 , 
n20255 , n20256 , n20257 , n20258 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , 
n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , 
n20276 , n20277 , n20278 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , 
n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , 
n20298 , n20299 , n20300 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , 
n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , 
n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , 
n20329 , n20331 , n20332 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , 
n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20350 , n20351 , 
n20352 , n20353 , n20354 , n20356 , n20357 , n20358 , n20360 , n20361 , n20362 , n20363 , 
n20364 , n20365 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , 
n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , 
n20386 , n20387 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , 
n20397 , n20398 , n20399 , n20400 , n20401 , n20404 , n20405 , n20406 , n20407 , n20408 , 
n20410 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , 
n20421 , n20422 , n20423 , n20425 , n20426 , n20427 , n20428 , n20430 , n20431 , n20432 , 
n20433 , n20434 , n20435 , n20437 , n20438 , n20439 , n20440 , n20442 , n20443 , n20444 , 
n20446 , n20447 , n20448 , n20449 , n20451 , n20452 , n20453 , n20454 , n20456 , n20457 , 
n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , 
n20468 , n20469 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20479 , 
n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20491 , 
n20492 , n20493 , n20494 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , 
n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , 
n20513 , n20514 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , 
n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20534 , 
n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , 
n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , 
n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , 
n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , 
n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20583 , n20584 , n20585 , 
n20586 , n20587 , n20588 , n20589 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , 
n20597 , n20598 , n20599 , n20600 , n20601 , n20603 , n20605 , n20606 , n20607 , n20608 , 
n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , 
n20620 , n20621 , n20622 , n20624 , n20625 , n20626 , n20627 , n20628 , n20630 , n20631 , 
n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , 
n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , 
n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20659 , n20660 , n20662 , n20663 , 
n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20674 , 
n20675 , n20676 , n20677 , n20679 , n20681 , n20682 , n20683 , n20684 , n20686 , n20687 , 
n20688 , n20689 , n20690 , n20692 , n20693 , n20694 , n20695 , n20697 , n20698 , n20699 , 
n20701 , n20702 , n20703 , n20706 , n20707 , n20708 , n20710 , n20711 , n20712 , n20714 , 
n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20724 , n20725 , n20726 , 
n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , 
n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , 
n20747 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , 
n20758 , n20759 , n20760 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , 
n20769 , n20770 , n20771 , n20772 , n20773 , n20775 , n20776 , n20777 , n20778 , n20779 , 
n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20789 , n20790 , 
n20791 , n20792 , n20793 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , 
n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , 
n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , 
n20824 , n20825 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , 
n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , 
n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , 
n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , 
n20865 , n20866 , n20867 , n20868 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , 
n20876 , n20877 , n20878 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , 
n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , 
n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , 
n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20916 , n20917 , 
n20918 , n20919 , n20920 , n20921 , n20922 , n20924 , n20925 , n20926 , n20927 , n20928 , 
n20930 , n20931 , n20932 , n20933 , n20934 , n20937 , n20938 , n20939 , n20940 , n20941 , 
n20942 , n20943 , n20944 , n20945 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , 
n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , 
n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , 
n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , 
n20983 , n20984 , n20985 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , 
n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , 
n21004 , n21005 , n21006 , n21007 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , 
n21015 , n21016 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , 
n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21035 , n21036 , 
n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21047 , 
n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , 
n21058 , n21059 , n21060 , n21061 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , 
n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21079 , 
n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , 
n21090 , n21091 , n21092 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , 
n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , 
n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , 
n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , 
n21135 , n21136 , n21137 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , 
n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21155 , n21156 , 
n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , 
n21169 , n21170 , n21171 , n21172 , n21174 , n21175 , n21177 , n21178 , n21179 , n21180 , 
n21181 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , 
n21192 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , 
n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , 
n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21223 , n21224 , 
n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , 
n21237 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , 
n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21255 , n21256 , n21257 , n21258 , 
n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , 
n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21277 , n21278 , n21279 , 
n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21288 , n21289 , n21290 , 
n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21299 , n21300 , n21301 , 
n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , 
n21313 , n21314 , n21315 , n21316 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , 
n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , 
n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , 
n21344 , n21345 , n21346 , n21347 , n21348 , n21350 , n21351 , n21352 , n21353 , n21354 , 
n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , 
n21366 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , 
n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , 
n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21397 , 
n21400 , n21401 , n21402 , n21403 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , 
n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , 
n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , 
n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , 
n21441 , n21442 , n21443 , n21444 , n21445 , n21447 , n21448 , n21449 , n21450 , n21451 , 
n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , 
n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21473 , 
n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , 
n21484 , n21485 , n21486 , n21487 , n21488 , n21490 , n21491 , n21492 , n21493 , n21494 , 
n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , 
n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , 
n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , 
n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , 
n21536 , n21537 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , 
n21547 , n21548 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , 
n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , 
n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , 
n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , 
n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , 
n21598 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , 
n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21616 , n21617 , n21618 , n21619 , 
n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21629 , n21630 , 
n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21638 , n21639 , n21640 , n21641 , 
n21642 , n21643 , n21644 , n21646 , n21647 , n21648 , n21650 , n21651 , n21652 , n21653 , 
n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , 
n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21675 , n21676 , 
n21677 , n21678 , n21679 , n21681 , n21682 , n21683 , n21684 , n21686 , n21688 , n21689 , 
n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , 
n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , 
n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21718 , n21720 , n21721 , 
n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , 
n21732 , n21733 , n21734 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , 
n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21751 , n21752 , n21754 , n21755 , 
n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21766 , 
n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , 
n21777 , n21778 , n21780 , n21781 , n21782 , n21783 , n21785 , n21786 , n21787 , n21788 , 
n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , 
n21799 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , 
n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , 
n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , 
n21831 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21840 , n21841 , n21842 , 
n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , 
n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , 
n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , 
n21873 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , 
n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , 
n21894 , n21895 , n21896 , n21897 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , 
n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21916 , 
n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , 
n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21935 , n21936 , n21937 , 
n21938 , n21939 , n21940 , n21941 , n21942 , n21944 , n21945 , n21946 , n21947 , n21948 , 
n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21958 , n21959 , 
n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , 
n21971 , n21972 , n21973 , n21974 , n21975 , n21977 , n21978 , n21979 , n21980 , n21982 , 
n21983 , n21984 , n21985 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21994 , 
n21995 , n21996 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , 
n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , 
n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , 
n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , 
n22038 , n22039 , n22040 , n22041 , n22042 , n22044 , n22045 , n22046 , n22047 , n22048 , 
n22049 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , 
n22060 , n22061 , n22062 , n22064 , n22065 , n22066 , n22067 , n22069 , n22070 , n22071 , 
n22073 , n22074 , n22075 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , 
n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22091 , n22092 , n22093 , n22094 , 
n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , 
n22105 , n22106 , n22108 , n22109 , n22110 , n22111 , n22112 , n22114 , n22115 , n22116 , 
n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22125 , n22127 , n22128 , 
n22129 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , 
n22140 , n22141 , n22142 , n22143 , n22145 , n22146 , n22147 , n22148 , n22149 , n22151 , 
n22152 , n22153 , n22154 , n22155 , n22156 , n22158 , n22159 , n22160 , n22161 , n22162 , 
n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , 
n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , 
n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , 
n22194 , n22195 , n22196 , n22197 , n22199 , n22200 , n22202 , n22203 , n22204 , n22205 , 
n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22214 , n22215 , n22216 , 
n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , 
n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , 
n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , 
n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22254 , n22255 , n22256 , n22257 , 
n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , 
n22268 , n22269 , n22271 , n22272 , n22273 , n22275 , n22276 , n22277 , n22278 , n22279 , 
n22280 , n22281 , n22282 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22291 , 
n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , 
n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22310 , n22312 , n22313 , 
n22314 , n22315 , n22316 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , 
n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22333 , n22334 , n22336 , 
n22337 , n22338 , n22339 , n22340 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , 
n22348 , n22349 , n22350 , n22351 , n22352 , n22354 , n22355 , n22356 , n22357 , n22360 , 
n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , 
n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22380 , n22381 , 
n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , 
n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , 
n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , 
n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , 
n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , 
n22432 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22443 , 
n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , 
n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , 
n22465 , n22466 , n22468 , n22469 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , 
n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22485 , n22486 , n22487 , 
n22488 , n22490 , n22491 , n22493 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , 
n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , 
n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , 
n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , 
n22531 , n22532 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , 
n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , 
n22552 , n22553 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , 
n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , 
n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , 
n22583 , n22585 , n22586 , n22587 , n22590 , n22592 , n22593 , n22594 , n22595 , n22596 , 
n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , 
n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , 
n22618 , n22621 , n22622 , n22624 , n22625 , n22627 , n22628 , n22629 , n22630 , n22632 , 
n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , 
n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , 
n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22661 , n22662 , n22663 , 
n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , 
n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , 
n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , 
n22694 , n22695 , n22696 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , 
n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22715 , 
n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , 
n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , 
n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , 
n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , 
n22756 , n22757 , n22758 , n22759 , n22760 , n22762 , n22763 , n22765 , n22766 , n22767 , 
n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , 
n22778 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22788 , n22789 , 
n22790 , n22791 , n22792 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , 
n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , 
n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22820 , n22821 , 
n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , 
n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , 
n22842 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , 
n22853 , n22854 , n22855 , n22856 , n22857 , n22859 , n22860 , n22861 , n22862 , n22863 , 
n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22872 , n22873 , n22874 , n22875 , 
n22876 , n22877 , n22878 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , 
n22887 , n22888 , n22889 , n22890 , n22892 , n22893 , n22894 , n22895 , n22896 , n22898 , 
n22899 , n22900 , n22901 , n22902 , n22904 , n22905 , n22906 , n22908 , n22909 , n22911 , 
n22912 , n22913 , n22915 , n22916 , n22917 , n22919 , n22920 , n22921 , n22922 , n22923 , 
n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , 
n22934 , n22935 , n22936 , n22937 , n22938 , n22940 , n22941 , n22942 , n22943 , n22944 , 
n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , 
n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , 
n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , 
n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , 
n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , 
n22995 , n22996 , n22997 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , 
n23008 , n23010 , n23011 , n23012 , n23013 , n23015 , n23016 , n23017 , n23018 , n23019 , 
n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , 
n23030 , n23031 , n23032 , n23033 , n23034 , n23036 , n23037 , n23038 , n23040 , n23041 , 
n23042 , n23043 , n23044 , n23045 , n23046 , n23048 , n23049 , n23050 , n23051 , n23052 , 
n23053 , n23054 , n23055 , n23056 , n23057 , n23059 , n23060 , n23061 , n23062 , n23063 , 
n23064 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , 
n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , 
n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , 
n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , 
n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , 
n23118 , n23119 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , 
n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , 
n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23147 , n23148 , n23149 , 
n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , 
n23161 , n23162 , n23163 , n23164 , n23165 , n23167 , n23168 , n23169 , n23170 , n23171 , 
n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , 
n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , 
n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23201 , n23202 , 
n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , 
n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , 
n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , 
n23233 , n23234 , n23235 , n23236 , n23237 , n23239 , n23240 , n23241 , n23242 , n23243 , 
n23244 , n23245 , n23246 , n23249 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , 
n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , 
n23267 , n23268 , n23269 , n23271 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , 
n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , 
n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , 
n23300 , n23301 , n23302 , n23303 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , 
n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , 
n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , 
n23332 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23343 , n23344 , 
n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , 
n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , 
n23366 , n23367 , n23368 , n23370 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , 
n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , 
n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , 
n23398 , n23399 , n23400 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , 
n23409 , n23410 , n23411 , n23412 , n23413 , n23415 , n23416 , n23417 , n23418 , n23419 , 
n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23431 , 
n23432 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , 
n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23451 , n23452 , n23453 , n23454 , 
n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23464 , n23465 , 
n23466 , n23467 , n23468 , n23469 , n23470 , n23472 , n23473 , n23474 , n23475 , n23476 , 
n23477 , n23478 , n23479 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , 
n23488 , n23489 , n23490 , n23491 , n23492 , n23494 , n23495 , n23496 , n23497 , n23498 , 
n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , 
n23509 , n23510 , n23511 , n23512 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , 
n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23530 , 
n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , 
n23542 , n23543 , n23544 , n23545 , n23547 , n23548 , n23549 , n23551 , n23552 , n23553 , 
n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , 
n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , 
n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , 
n23584 , n23587 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , 
n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , 
n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , 
n23617 , n23618 , n23620 , n23621 , n23622 , n23623 , n23625 , n23626 , n23627 , n23629 , 
n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23638 , n23639 , n23640 , 
n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , 
n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23658 , n23659 , n23660 , n23661 , 
n23662 , n23664 , n23665 , n23666 , n23667 , n23668 , n23670 , n23671 , n23672 , n23673 , 
n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , 
n23685 , n23686 , n23687 , n23688 , n23689 , n23691 , n23692 , n23693 , n23694 , n23695 , 
n23696 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , 
n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23715 , n23716 , n23718 , 
n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , 
n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , 
n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23749 , n23750 , 
n23751 , n23752 , n23753 , n23754 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , 
n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , 
n23772 , n23773 , n23774 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , 
n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , 
n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , 
n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , 
n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , 
n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23832 , n23833 , 
n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23843 , n23844 , 
n23845 , n23846 , n23847 , n23848 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , 
n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , 
n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , 
n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23884 , n23885 , n23886 , n23887 , 
n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23896 , n23897 , n23898 , n23900 , 
n23901 , n23902 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , 
n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23925 , 
n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23936 , 
n23937 , n23938 , n23939 , n23940 , n23941 , n23943 , n23944 , n23945 , n23946 , n23947 , 
n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23955 , n23956 , n23957 , n23959 , 
n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , 
n23970 , n23971 , n23972 , n23973 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , 
n23981 , n23982 , n23983 , n23984 , n23985 , n23987 , n23988 , n23989 , n23990 , n23991 , 
n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , 
n24003 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , 
n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , 
n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24033 , n24034 , 
n24035 , n24036 , n24037 , n24038 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , 
n24046 , n24047 , n24049 , n24050 , n24051 , n24053 , n24054 , n24055 , n24056 , n24057 , 
n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , 
n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , 
n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24086 , n24087 , n24088 , 
n24089 , n24090 , n24091 , n24094 , n24095 , n24098 , n24099 , n24100 , n24101 , n24102 , 
n24103 , n24104 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , 
n24114 , n24115 , n24116 , n24117 , n24118 , n24120 , n24121 , n24122 , n24123 , n24124 , 
n24125 , n24126 , n24127 , n24128 , n24130 , n24131 , n24132 , n24134 , n24135 , n24136 , 
n24137 , n24138 , n24139 , n24140 , n24142 , n24143 , n24144 , n24147 , n24148 , n24149 , 
n24151 , n24152 , n24153 , n24154 , n24156 , n24157 , n24158 , n24159 , n24161 , n24162 , 
n24163 , n24164 , n24165 , n24166 , n24168 , n24169 , n24171 , n24173 , n24174 , n24175 , 
n24176 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , 
n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24197 , 
n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , 
n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , 
n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , 
n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , 
n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , 
n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24259 , 
n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , 
n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24279 , n24280 , n24281 , 
n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24290 , n24291 , n24292 , 
n24293 , n24294 , n24295 , n24296 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , 
n24304 , n24305 , n24306 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , 
n24315 , n24316 , n24317 , n24318 , n24320 , n24321 , n24322 , n24324 , n24325 , n24326 , 
n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , 
n24338 , n24339 , n24340 , n24341 , n24343 , n24344 , n24346 , n24348 , n24349 , n24350 , 
n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , 
n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , 
n24371 , n24372 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , 
n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , 
n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , 
n24403 , n24404 , n24405 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , 
n24414 , n24416 , n24417 , n24418 , n24419 , n24420 , n24422 , n24423 , n24424 , n24425 , 
n24426 , n24427 , n24428 , n24429 , n24430 , n24432 , n24433 , n24434 , n24435 , n24436 , 
n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , 
n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , 
n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , 
n24467 , n24468 , n24469 , n24470 , n24471 , n24473 , n24474 , n24475 , n24477 , n24478 , 
n24479 , n24480 , n24481 , n24482 , n24484 , n24486 , n24487 , n24488 , n24489 , n24490 , 
n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , 
n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , 
n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , 
n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , 
n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , 
n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , 
n24553 , n24554 , n24555 , n24556 , n24557 , n24559 , n24560 , n24561 , n24562 , n24563 , 
n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , 
n24574 , n24575 , n24577 , n24578 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , 
n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , 
n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24603 , n24605 , n24606 , n24607 , 
n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , 
n24619 , n24621 , n24622 , n24623 , n24624 , n24625 , n24627 , n24628 , n24630 , n24631 , 
n24632 , n24633 , n24634 , n24635 , n24637 , n24639 , n24640 , n24641 , n24642 , n24643 , 
n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , 
n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , 
n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , 
n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , 
n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , 
n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , 
n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , 
n24714 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24724 , n24725 , 
n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24733 , n24734 , n24735 , n24736 , 
n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , 
n24747 , n24748 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , 
n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24769 , 
n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , 
n24780 , n24781 , n24782 , n24783 , n24785 , n24787 , n24788 , n24789 , n24790 , n24791 , 
n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , 
n24802 , n24803 , n24804 , n24805 , n24806 , n24808 , n24809 , n24810 , n24811 , n24812 , 
n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , 
n24823 , n24824 , n24825 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , 
n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24842 , n24843 , n24844 , n24845 , 
n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24854 , n24855 , n24856 , 
n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , 
n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , 
n24878 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24888 , n24889 , 
n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , 
n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , 
n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , 
n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , 
n24930 , n24931 , n24932 , n24933 , n24935 , n24936 , n24938 , n24939 , n24940 , n24941 , 
n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , 
n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , 
n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , 
n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , 
n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , 
n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24999 , n25000 , n25001 , n25002 , 
n25003 , n25004 , n25005 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , 
n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25024 , 
n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25033 , n25034 , n25035 , 
n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , 
n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , 
n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25063 , n25064 , n25065 , n25066 , 
n25067 , n25069 , n25070 , n25071 , n25072 , n25075 , n25076 , n25077 , n25078 , n25079 , 
n25080 , n25081 , n25082 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , 
n25091 , n25092 , n25093 , n25095 , n25096 , n25098 , n25099 , n25100 , n25101 , n25102 , 
n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , 
n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25121 , n25122 , n25123 , n25124 , 
n25125 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25134 , n25135 , n25136 , 
n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , 
n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25156 , n25157 , 
n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , 
n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , 
n25179 , n25180 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , 
n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , 
n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25210 , n25211 , 
n25212 , n25213 , n25214 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , 
n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , 
n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25241 , n25242 , n25243 , 
n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25255 , 
n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , 
n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , 
n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , 
n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25294 , n25295 , n25297 , n25298 , 
n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , 
n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25317 , n25318 , n25319 , 
n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25329 , n25330 , 
n25333 , n25334 , n25335 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , 
n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , 
n25357 , n25358 , n25359 , n25360 , n25361 , n25363 , n25364 , n25366 , n25367 , n25368 , 
n25369 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , 
n25380 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , 
n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , 
n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , 
n25411 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , 
n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , 
n25432 , n25433 , n25434 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , 
n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , 
n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25461 , n25462 , n25463 , 
n25465 , n25466 , n25467 , n25469 , n25470 , n25472 , n25473 , n25474 , n25476 , n25477 , 
n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , 
n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25495 , n25496 , n25497 , n25498 , 
n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , 
n25510 , n25511 , n25512 , n25514 , n25515 , n25516 , n25517 , n25519 , n25520 , n25521 , 
n25522 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25533 , 
n25534 , n25535 , n25536 , n25537 , n25538 , n25540 , n25541 , n25542 , n25543 , n25544 , 
n25545 , n25546 , n25547 , n25548 , n25549 , n25551 , n25552 , n25553 , n25554 , n25555 , 
n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25566 , 
n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , 
n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25587 , 
n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , 
n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , 
n25608 , n25609 , n25610 , n25612 , n25613 , n25615 , n25616 , n25617 , n25618 , n25620 , 
n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25630 , n25631 , 
n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , 
n25642 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , 
n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , 
n25663 , n25664 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , 
n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , 
n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , 
n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , 
n25705 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , 
n25716 , n25717 , n25718 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , 
n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , 
n25737 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , 
n25748 , n25750 , n25752 , n25753 , n25754 , n25755 , n25757 , n25759 , n25760 , n25761 , 
n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , 
n25772 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , 
n25783 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25793 , n25794 , 
n25795 , n25796 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , 
n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , 
n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25827 , 
n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , 
n25838 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , 
n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , 
n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , 
n25870 , n25871 , n25874 , n25875 , n25876 , n25878 , n25879 , n25880 , n25881 , n25882 , 
n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , 
n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , 
n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , 
n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , 
n25924 , n25925 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25935 , 
n25936 , n25937 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , 
n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , 
n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , 
n25967 , n25968 , n25969 , n25970 , n25971 , n25973 , n25975 , n25976 , n25977 , n25978 , 
n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25986 , n25987 , n25988 , n25989 , 
n25990 , n25991 , n25992 , n25993 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , 
n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , 
n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , 
n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , 
n26031 , n26032 , n26033 , n26034 , n26035 , n26037 , n26038 , n26039 , n26040 , n26041 , 
n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , 
n26052 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , 
n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , 
n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , 
n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , 
n26095 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , 
n26106 , n26108 , n26109 , n26110 , n26112 , n26114 , n26115 , n26116 , n26117 , n26118 , 
n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , 
n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , 
n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , 
n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26157 , n26158 , n26160 , 
n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26168 , n26169 , n26170 , n26171 , 
n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26181 , n26182 , n26183 , 
n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26192 , n26193 , n26194 , 
n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , 
n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , 
n26215 , n26216 , n26217 , n26218 , n26219 , n26221 , n26222 , n26223 , n26225 , n26226 , 
n26227 , n26228 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26238 , 
n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , 
n26249 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , 
n26260 , n26261 , n26262 , n26263 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , 
n26271 , n26272 , n26273 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , 
n26282 , n26283 , n26284 , n26285 , n26286 , n26288 , n26289 , n26290 , n26291 , n26292 , 
n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , 
n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , 
n26313 , n26314 , n26315 , n26316 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , 
n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , 
n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , 
n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26354 , n26355 , 
n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , 
n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26376 , 
n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , 
n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26397 , 
n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , 
n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , 
n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , 
n26430 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26440 , n26441 , 
n26442 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26453 , 
n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , 
n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , 
n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26484 , 
n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26493 , n26494 , n26495 , 
n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , 
n26506 , n26507 , n26508 , n26509 , n26511 , n26513 , n26514 , n26516 , n26517 , n26518 , 
n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , 
n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26539 , 
n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , 
n26550 , n26551 , n26552 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , 
n26561 , n26562 , n26563 , n26564 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , 
n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , 
n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26591 , n26592 , n26593 , 
n26594 , n26595 , n26596 , n26597 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , 
n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , 
n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26626 , 
n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , 
n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , 
n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26657 , 
n26658 , n26659 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , 
n26669 , n26670 , n26671 , n26672 , n26673 , n26676 , n26677 , n26678 , n26679 , n26680 , 
n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , 
n26692 , n26693 , n26694 , n26695 , n26697 , n26699 , n26700 , n26701 , n26702 , n26703 , 
n26704 , n26705 , n26706 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , 
n26715 , n26716 , n26717 , n26718 , n26720 , n26721 , n26722 , n26723 , n26724 , n26726 , 
n26728 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , 
n26739 , n26740 , n26741 , n26742 , n26743 , n26746 , n26747 , n26749 , n26750 , n26751 , 
n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , 
n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , 
n26773 , n26774 , n26776 , n26777 , n26778 , n26779 , n26781 , n26782 , n26783 , n26784 , 
n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26796 , 
n26798 , n26799 , n26800 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26809 , 
n26810 , n26811 , n26812 , n26813 , n26814 , n26816 , n26817 , n26818 , n26819 , n26820 , 
n26821 , n26822 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , 
n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , 
n26842 , n26843 , n26844 , n26845 , n26846 , n26848 , n26849 , n26850 , n26851 , n26852 , 
n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , 
n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , 
n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26883 , 
n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , 
n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26901 , n26903 , n26904 , n26906 , 
n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26914 , n26915 , n26916 , n26917 , 
n26918 , n26919 , n26920 , n26922 , n26924 , n26925 , n26926 , n26927 , n26928 , n26931 , 
n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , 
n26942 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , 
n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , 
n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26971 , n26972 , n26973 , 
n26974 , n26975 , n26976 , n26977 , n26978 , n26980 , n26981 , n26982 , n26983 , n26984 , 
n26985 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , 
n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27005 , n27006 , 
n27007 , n27008 , n27009 , n27010 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , 
n27018 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , 
n27029 , n27030 , n27032 , n27033 , n27034 , n27035 , n27036 , n27038 , n27039 , n27040 , 
n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , 
n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , 
n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , 
n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27080 , n27081 , n27082 , n27083 , 
n27084 , n27085 , n27086 , n27087 , n27088 , n27090 , n27091 , n27092 , n27093 , n27094 , 
n27095 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27105 , n27106 , 
n27107 , n27108 , n27109 , n27111 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , 
n27119 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , 
n27131 , n27132 , n27133 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , 
n27142 , n27143 , n27144 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , 
n27153 , n27154 , n27155 , n27156 , n27157 , n27159 , n27160 , n27161 , n27162 , n27164 , 
n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , 
n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , 
n27185 , n27186 , n27187 , n27189 , n27190 , n27191 , n27192 , n27193 , n27195 , n27196 , 
n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 ;
    or g0 ( n25456 , n12222 , n17800 );
    not g1 ( n4950 , n24186 );
    and g2 ( n12724 , n24693 , n14425 );
    or g3 ( n5884 , n17333 , n19247 );
    not g4 ( n13231 , n1735 );
    or g5 ( n363 , n15446 , n2417 );
    or g6 ( n12601 , n3124 , n3018 );
    not g7 ( n54 , n21300 );
    xnor g8 ( n21820 , n20820 , n14706 );
    not g9 ( n22318 , n12713 );
    not g10 ( n21745 , n21544 );
    not g11 ( n15177 , n13572 );
    or g12 ( n26507 , n22220 , n14118 );
    or g13 ( n11793 , n1963 , n21122 );
    xnor g14 ( n17152 , n3747 , n21909 );
    xnor g15 ( n7943 , n20710 , n21590 );
    or g16 ( n6658 , n22626 , n8583 );
    or g17 ( n7064 , n17471 , n6429 );
    and g18 ( n27148 , n11024 , n25179 );
    or g19 ( n20223 , n23276 , n5847 );
    or g20 ( n21320 , n16928 , n25210 );
    not g21 ( n5572 , n14089 );
    or g22 ( n21011 , n14363 , n1476 );
    xnor g23 ( n8578 , n10709 , n18924 );
    not g24 ( n8495 , n20410 );
    not g25 ( n18595 , n12969 );
    not g26 ( n17670 , n4879 );
    or g27 ( n14512 , n9502 , n15705 );
    nor g28 ( n3873 , n24313 , n26728 );
    xnor g29 ( n11734 , n3824 , n7395 );
    xnor g30 ( n3299 , n23618 , n8329 );
    xnor g31 ( n17003 , n21347 , n15280 );
    and g32 ( n2679 , n24317 , n6516 );
    not g33 ( n13649 , n3590 );
    nor g34 ( n8887 , n623 , n11195 );
    nor g35 ( n25052 , n18717 , n15155 );
    or g36 ( n24531 , n10568 , n18558 );
    xnor g37 ( n15082 , n26753 , n7886 );
    and g38 ( n20173 , n2268 , n22417 );
    and g39 ( n12897 , n22856 , n10163 );
    xnor g40 ( n11091 , n11016 , n9883 );
    or g41 ( n14307 , n9910 , n23272 );
    not g42 ( n22644 , n5060 );
    xnor g43 ( n21615 , n7998 , n12883 );
    not g44 ( n23233 , n25902 );
    or g45 ( n8928 , n20833 , n9536 );
    or g46 ( n865 , n20401 , n2489 );
    xnor g47 ( n23890 , n5059 , n14583 );
    not g48 ( n25890 , n1314 );
    and g49 ( n13709 , n8186 , n20797 );
    and g50 ( n12843 , n10218 , n4788 );
    and g51 ( n23844 , n5290 , n11851 );
    or g52 ( n16048 , n21071 , n2110 );
    xnor g53 ( n14394 , n27148 , n18538 );
    nor g54 ( n12328 , n9594 , n8285 );
    or g55 ( n26628 , n17013 , n10611 );
    not g56 ( n21340 , n10493 );
    or g57 ( n23817 , n8105 , n14522 );
    and g58 ( n17139 , n8123 , n10975 );
    xnor g59 ( n18341 , n3637 , n2783 );
    or g60 ( n5543 , n1522 , n14138 );
    or g61 ( n14935 , n20837 , n13470 );
    not g62 ( n1565 , n10660 );
    or g63 ( n20724 , n655 , n26253 );
    not g64 ( n21434 , n5196 );
    and g65 ( n4768 , n17860 , n16055 );
    or g66 ( n7011 , n1959 , n14473 );
    or g67 ( n756 , n21327 , n22876 );
    or g68 ( n18475 , n12342 , n16519 );
    or g69 ( n14183 , n14331 , n23294 );
    and g70 ( n15724 , n4638 , n49 );
    xnor g71 ( n4632 , n1509 , n16521 );
    xnor g72 ( n16576 , n20830 , n18596 );
    xnor g73 ( n4854 , n19259 , n5749 );
    or g74 ( n14775 , n1176 , n3480 );
    nor g75 ( n23867 , n22278 , n7465 );
    not g76 ( n8044 , n11095 );
    and g77 ( n10635 , n15870 , n5748 );
    nor g78 ( n24477 , n6232 , n13472 );
    or g79 ( n14912 , n4494 , n19986 );
    nor g80 ( n14542 , n16065 , n26413 );
    xnor g81 ( n515 , n575 , n3570 );
    and g82 ( n25252 , n22235 , n18699 );
    and g83 ( n10089 , n18505 , n8369 );
    and g84 ( n25395 , n8678 , n16500 );
    and g85 ( n21195 , n1041 , n13744 );
    nor g86 ( n22762 , n27037 , n20099 );
    xnor g87 ( n7811 , n17890 , n18231 );
    and g88 ( n1933 , n10763 , n18799 );
    and g89 ( n19474 , n14744 , n17936 );
    and g90 ( n7927 , n13762 , n10110 );
    and g91 ( n9079 , n15575 , n14072 );
    xnor g92 ( n20192 , n1084 , n21832 );
    or g93 ( n5519 , n2331 , n12546 );
    or g94 ( n21186 , n9493 , n15507 );
    xnor g95 ( n3755 , n15690 , n14252 );
    and g96 ( n20468 , n9401 , n25042 );
    xnor g97 ( n13095 , n12232 , n8526 );
    nor g98 ( n23133 , n26211 , n15583 );
    or g99 ( n1372 , n8309 , n24203 );
    nor g100 ( n2668 , n13137 , n7674 );
    or g101 ( n24057 , n161 , n24154 );
    or g102 ( n3922 , n22265 , n18194 );
    nor g103 ( n2669 , n7437 , n13367 );
    xnor g104 ( n2703 , n11983 , n18667 );
    and g105 ( n16256 , n6341 , n23512 );
    xnor g106 ( n10723 , n14032 , n14651 );
    not g107 ( n17620 , n1386 );
    or g108 ( n7046 , n18274 , n24202 );
    xnor g109 ( n16829 , n17629 , n8317 );
    or g110 ( n14470 , n20566 , n18211 );
    or g111 ( n11876 , n4957 , n5034 );
    and g112 ( n14443 , n2435 , n11984 );
    xnor g113 ( n2431 , n7107 , n5183 );
    or g114 ( n15706 , n23316 , n9122 );
    or g115 ( n5705 , n10620 , n17142 );
    xnor g116 ( n19749 , n93 , n12777 );
    xnor g117 ( n13300 , n5611 , n20600 );
    xnor g118 ( n5374 , n26758 , n13026 );
    xnor g119 ( n8315 , n813 , n19294 );
    xnor g120 ( n18433 , n21479 , n22435 );
    not g121 ( n25431 , n25353 );
    xnor g122 ( n11971 , n25146 , n13444 );
    xnor g123 ( n24147 , n20595 , n2322 );
    not g124 ( n3882 , n461 );
    or g125 ( n10007 , n3862 , n10392 );
    not g126 ( n19603 , n4660 );
    or g127 ( n25904 , n21860 , n1513 );
    or g128 ( n7266 , n6442 , n8959 );
    xnor g129 ( n2551 , n763 , n5222 );
    or g130 ( n16817 , n14465 , n23230 );
    xnor g131 ( n8805 , n106 , n22516 );
    xnor g132 ( n10240 , n21451 , n4893 );
    or g133 ( n1193 , n6054 , n16114 );
    nor g134 ( n12210 , n10113 , n11006 );
    and g135 ( n11367 , n9964 , n4880 );
    xnor g136 ( n3148 , n14733 , n13453 );
    and g137 ( n25666 , n1363 , n13692 );
    xnor g138 ( n25180 , n3349 , n25464 );
    or g139 ( n13307 , n6734 , n3 );
    xnor g140 ( n14050 , n7149 , n16971 );
    xnor g141 ( n17242 , n5160 , n5652 );
    or g142 ( n25351 , n18115 , n10837 );
    or g143 ( n14322 , n10557 , n8070 );
    not g144 ( n6900 , n20039 );
    and g145 ( n7028 , n8500 , n23716 );
    xnor g146 ( n23229 , n12869 , n17277 );
    or g147 ( n9097 , n27185 , n4660 );
    and g148 ( n7665 , n11446 , n8831 );
    nor g149 ( n5432 , n16573 , n788 );
    not g150 ( n19127 , n7180 );
    and g151 ( n16090 , n11041 , n7112 );
    xnor g152 ( n13296 , n12880 , n24684 );
    xnor g153 ( n19164 , n18845 , n6021 );
    xnor g154 ( n14832 , n6554 , n26205 );
    or g155 ( n4327 , n13590 , n1765 );
    or g156 ( n10396 , n23973 , n6738 );
    or g157 ( n22728 , n26642 , n3569 );
    and g158 ( n25020 , n2497 , n25695 );
    or g159 ( n5953 , n4760 , n24711 );
    xnor g160 ( n20039 , n14219 , n12529 );
    xnor g161 ( n6290 , n15519 , n5924 );
    or g162 ( n3398 , n17098 , n11510 );
    xnor g163 ( n23613 , n11056 , n20250 );
    nor g164 ( n21191 , n23474 , n12333 );
    xnor g165 ( n21760 , n4490 , n13167 );
    xnor g166 ( n948 , n9641 , n11267 );
    xnor g167 ( n20705 , n18839 , n22632 );
    and g168 ( n11480 , n24539 , n11709 );
    and g169 ( n3527 , n18851 , n5606 );
    xnor g170 ( n22908 , n22139 , n19472 );
    and g171 ( n5001 , n17173 , n1906 );
    xnor g172 ( n7592 , n22190 , n9243 );
    nor g173 ( n17403 , n8309 , n13158 );
    xnor g174 ( n20445 , n26203 , n24681 );
    and g175 ( n14640 , n6872 , n16559 );
    or g176 ( n7897 , n4098 , n13323 );
    or g177 ( n20679 , n4218 , n26981 );
    not g178 ( n9531 , n13034 );
    or g179 ( n16875 , n15258 , n4588 );
    xnor g180 ( n4886 , n19298 , n6611 );
    and g181 ( n11517 , n19939 , n26624 );
    or g182 ( n12118 , n18677 , n19416 );
    nor g183 ( n7712 , n10882 , n10760 );
    or g184 ( n13130 , n1796 , n21748 );
    xnor g185 ( n4765 , n24460 , n23261 );
    nor g186 ( n19631 , n24364 , n21280 );
    nor g187 ( n26458 , n25622 , n11945 );
    and g188 ( n19423 , n11452 , n14689 );
    nor g189 ( n5155 , n11161 , n8281 );
    and g190 ( n15747 , n23039 , n12734 );
    not g191 ( n21163 , n25168 );
    or g192 ( n5754 , n1402 , n24675 );
    not g193 ( n4667 , n16502 );
    and g194 ( n4472 , n13314 , n15099 );
    and g195 ( n20715 , n8773 , n10610 );
    xnor g196 ( n15624 , n17077 , n2289 );
    xnor g197 ( n4851 , n26702 , n1172 );
    xnor g198 ( n20595 , n11345 , n7045 );
    xnor g199 ( n21081 , n13233 , n8944 );
    and g200 ( n6340 , n7084 , n15381 );
    xnor g201 ( n1981 , n2765 , n15981 );
    xnor g202 ( n18154 , n16697 , n20293 );
    not g203 ( n18047 , n11185 );
    not g204 ( n7317 , n22014 );
    or g205 ( n18727 , n2659 , n16619 );
    and g206 ( n5368 , n3062 , n18047 );
    nor g207 ( n4347 , n25872 , n20196 );
    not g208 ( n21838 , n7329 );
    and g209 ( n7302 , n4078 , n25281 );
    xnor g210 ( n22353 , n4751 , n15406 );
    nor g211 ( n11827 , n19157 , n22379 );
    or g212 ( n15264 , n24610 , n8900 );
    and g213 ( n19781 , n13780 , n21949 );
    not g214 ( n11533 , n24609 );
    xnor g215 ( n22679 , n11841 , n2479 );
    nor g216 ( n9670 , n1777 , n26724 );
    or g217 ( n8390 , n5712 , n16701 );
    or g218 ( n4145 , n22764 , n14448 );
    or g219 ( n3747 , n6395 , n1335 );
    and g220 ( n17073 , n6739 , n25488 );
    not g221 ( n11535 , n61 );
    nor g222 ( n17782 , n2268 , n11503 );
    xnor g223 ( n14931 , n8901 , n14919 );
    xnor g224 ( n10150 , n16366 , n3018 );
    and g225 ( n26798 , n1750 , n21321 );
    and g226 ( n21172 , n14979 , n14317 );
    not g227 ( n8454 , n2481 );
    and g228 ( n19713 , n16773 , n4219 );
    or g229 ( n716 , n4892 , n21466 );
    and g230 ( n3084 , n22312 , n3762 );
    or g231 ( n8790 , n7861 , n16401 );
    xnor g232 ( n22973 , n19789 , n15424 );
    or g233 ( n22573 , n15809 , n4721 );
    and g234 ( n10803 , n18813 , n7219 );
    nor g235 ( n16509 , n23408 , n25643 );
    xnor g236 ( n7407 , n12653 , n18965 );
    nor g237 ( n9060 , n21114 , n17814 );
    or g238 ( n14476 , n14149 , n2397 );
    and g239 ( n6291 , n21905 , n24481 );
    not g240 ( n12475 , n12920 );
    not g241 ( n12105 , n9731 );
    xnor g242 ( n21131 , n19529 , n4049 );
    xnor g243 ( n23383 , n20487 , n2968 );
    nor g244 ( n7606 , n8155 , n10763 );
    and g245 ( n21938 , n22479 , n18618 );
    xnor g246 ( n20221 , n20235 , n6502 );
    nor g247 ( n57 , n5231 , n14048 );
    or g248 ( n20143 , n11891 , n18985 );
    or g249 ( n15550 , n2156 , n18931 );
    xnor g250 ( n26248 , n18985 , n26931 );
    not g251 ( n1587 , n3785 );
    not g252 ( n7948 , n22043 );
    not g253 ( n21208 , n10899 );
    xnor g254 ( n20919 , n7437 , n17077 );
    or g255 ( n4126 , n20801 , n6363 );
    or g256 ( n14123 , n20898 , n5110 );
    or g257 ( n16494 , n20658 , n6307 );
    xnor g258 ( n527 , n13828 , n19905 );
    xnor g259 ( n2706 , n18949 , n15725 );
    and g260 ( n11654 , n23487 , n18542 );
    or g261 ( n7595 , n4845 , n24624 );
    and g262 ( n16415 , n15041 , n13224 );
    xnor g263 ( n16276 , n19067 , n17643 );
    not g264 ( n26105 , n9043 );
    or g265 ( n21053 , n20583 , n3298 );
    not g266 ( n10499 , n13333 );
    nor g267 ( n3022 , n856 , n11365 );
    or g268 ( n14956 , n3293 , n25189 );
    nor g269 ( n24457 , n7057 , n14570 );
    xnor g270 ( n16788 , n15282 , n9859 );
    or g271 ( n12294 , n13106 , n21028 );
    xnor g272 ( n25063 , n25066 , n8827 );
    not g273 ( n5963 , n14580 );
    or g274 ( n13726 , n10120 , n22629 );
    and g275 ( n11858 , n13712 , n6945 );
    or g276 ( n15324 , n10885 , n19276 );
    or g277 ( n9816 , n5255 , n25289 );
    xnor g278 ( n15325 , n2436 , n11714 );
    and g279 ( n24407 , n1867 , n14308 );
    xnor g280 ( n9499 , n7099 , n6691 );
    and g281 ( n1328 , n11634 , n3437 );
    xnor g282 ( n13504 , n3840 , n24908 );
    xnor g283 ( n26668 , n17141 , n494 );
    or g284 ( n4863 , n7974 , n24618 );
    xnor g285 ( n9086 , n12050 , n19982 );
    and g286 ( n22543 , n12589 , n22979 );
    or g287 ( n11487 , n26312 , n13873 );
    or g288 ( n1966 , n6406 , n12100 );
    xnor g289 ( n13157 , n14440 , n14130 );
    or g290 ( n12779 , n25890 , n25494 );
    xnor g291 ( n13836 , n10951 , n13895 );
    xnor g292 ( n11275 , n24719 , n26343 );
    xnor g293 ( n10284 , n18724 , n6891 );
    not g294 ( n13539 , n7416 );
    nor g295 ( n25658 , n13459 , n15167 );
    and g296 ( n20563 , n342 , n26789 );
    or g297 ( n22920 , n4687 , n19245 );
    not g298 ( n13898 , n9399 );
    or g299 ( n1271 , n22459 , n9662 );
    xnor g300 ( n20838 , n12341 , n15053 );
    xnor g301 ( n17975 , n7112 , n20919 );
    xnor g302 ( n6683 , n26499 , n25604 );
    nor g303 ( n7757 , n6173 , n12917 );
    xnor g304 ( n19576 , n9557 , n16158 );
    xnor g305 ( n6412 , n4469 , n25071 );
    xnor g306 ( n8569 , n16377 , n4269 );
    xnor g307 ( n25816 , n16538 , n4506 );
    not g308 ( n7005 , n24557 );
    and g309 ( n1377 , n18980 , n22096 );
    and g310 ( n16007 , n2342 , n12984 );
    and g311 ( n10161 , n4419 , n8291 );
    or g312 ( n7063 , n13563 , n26889 );
    xnor g313 ( n4764 , n18286 , n1884 );
    xor g314 ( n12884 , n10995 , n6397 );
    xnor g315 ( n25784 , n17067 , n2946 );
    nor g316 ( n6744 , n6698 , n20556 );
    nor g317 ( n17836 , n10169 , n7133 );
    xnor g318 ( n24561 , n10188 , n25738 );
    xnor g319 ( n13660 , n6794 , n14090 );
    and g320 ( n35 , n24337 , n11954 );
    and g321 ( n12736 , n3988 , n8686 );
    xnor g322 ( n25985 , n2475 , n1419 );
    not g323 ( n6568 , n1710 );
    not g324 ( n17409 , n12137 );
    xnor g325 ( n13119 , n5741 , n15081 );
    or g326 ( n3031 , n120 , n21687 );
    xnor g327 ( n22493 , n6731 , n5066 );
    or g328 ( n18996 , n17826 , n23878 );
    or g329 ( n8137 , n13786 , n10242 );
    xnor g330 ( n14675 , n14400 , n6857 );
    xnor g331 ( n972 , n18178 , n18840 );
    and g332 ( n27090 , n7300 , n6793 );
    xnor g333 ( n24135 , n27081 , n1622 );
    xnor g334 ( n6620 , n7871 , n5696 );
    or g335 ( n9790 , n15944 , n2783 );
    not g336 ( n15845 , n6719 );
    or g337 ( n24339 , n15651 , n3613 );
    nor g338 ( n25571 , n1835 , n2645 );
    nor g339 ( n83 , n3009 , n1288 );
    not g340 ( n15405 , n2868 );
    not g341 ( n20630 , n11941 );
    or g342 ( n13085 , n8518 , n231 );
    xnor g343 ( n26538 , n3658 , n23325 );
    not g344 ( n21224 , n21291 );
    xnor g345 ( n25867 , n8609 , n9584 );
    nor g346 ( n6067 , n746 , n27078 );
    and g347 ( n11805 , n12446 , n966 );
    xnor g348 ( n24508 , n23876 , n14477 );
    or g349 ( n24891 , n20667 , n14151 );
    xnor g350 ( n19204 , n56 , n17590 );
    or g351 ( n3494 , n11989 , n2981 );
    or g352 ( n7513 , n5364 , n22653 );
    or g353 ( n20318 , n17110 , n17502 );
    or g354 ( n21806 , n1848 , n5421 );
    xnor g355 ( n5980 , n21920 , n6210 );
    xnor g356 ( n15458 , n9504 , n26524 );
    xnor g357 ( n6756 , n20210 , n19144 );
    or g358 ( n1600 , n23793 , n12004 );
    not g359 ( n6946 , n25947 );
    or g360 ( n18713 , n24126 , n18359 );
    not g361 ( n17626 , n13621 );
    xnor g362 ( n10442 , n12423 , n9259 );
    xnor g363 ( n18123 , n3128 , n4566 );
    xnor g364 ( n14973 , n19446 , n3931 );
    xnor g365 ( n15408 , n5858 , n10127 );
    xnor g366 ( n12950 , n2333 , n5161 );
    or g367 ( n7087 , n4920 , n26664 );
    or g368 ( n3768 , n3654 , n23601 );
    and g369 ( n15544 , n23267 , n25005 );
    or g370 ( n11914 , n13186 , n11611 );
    xnor g371 ( n12440 , n9251 , n2387 );
    nor g372 ( n17092 , n17184 , n18587 );
    or g373 ( n7482 , n24304 , n7425 );
    or g374 ( n16546 , n11731 , n16991 );
    and g375 ( n16539 , n3395 , n11939 );
    and g376 ( n21077 , n12963 , n6797 );
    xor g377 ( n12548 , n17409 , n26000 );
    xnor g378 ( n21540 , n1256 , n11281 );
    or g379 ( n19621 , n5140 , n14158 );
    and g380 ( n4099 , n1432 , n2852 );
    or g381 ( n9518 , n23000 , n24908 );
    or g382 ( n838 , n21593 , n7787 );
    xnor g383 ( n6999 , n17647 , n20146 );
    and g384 ( n14815 , n20922 , n17950 );
    or g385 ( n4354 , n26129 , n22292 );
    nor g386 ( n11856 , n21969 , n5949 );
    or g387 ( n27198 , n913 , n6390 );
    xnor g388 ( n16206 , n13191 , n12913 );
    or g389 ( n21009 , n19272 , n25541 );
    xnor g390 ( n16517 , n17914 , n4596 );
    and g391 ( n26581 , n397 , n5177 );
    not g392 ( n18861 , n22511 );
    and g393 ( n26762 , n6551 , n5527 );
    or g394 ( n24673 , n17812 , n4675 );
    or g395 ( n4421 , n5575 , n13019 );
    and g396 ( n16813 , n14440 , n7523 );
    or g397 ( n6439 , n21174 , n4065 );
    xnor g398 ( n16938 , n6658 , n1980 );
    or g399 ( n15148 , n7953 , n6397 );
    and g400 ( n22181 , n23178 , n3418 );
    nor g401 ( n25444 , n5547 , n3241 );
    or g402 ( n20481 , n14963 , n12379 );
    xnor g403 ( n25873 , n5008 , n24433 );
    or g404 ( n11434 , n1176 , n26913 );
    and g405 ( n16334 , n17645 , n10945 );
    or g406 ( n7564 , n3681 , n18510 );
    nor g407 ( n4676 , n19163 , n13945 );
    xnor g408 ( n13098 , n4212 , n15679 );
    and g409 ( n10079 , n21314 , n23051 );
    or g410 ( n15029 , n15935 , n22738 );
    nor g411 ( n3252 , n16183 , n5283 );
    xnor g412 ( n20936 , n15811 , n1943 );
    or g413 ( n11594 , n19386 , n6561 );
    not g414 ( n24130 , n10514 );
    or g415 ( n1871 , n22558 , n5733 );
    nor g416 ( n24229 , n16524 , n13668 );
    nor g417 ( n21341 , n24969 , n13124 );
    xnor g418 ( n4540 , n23688 , n12697 );
    xnor g419 ( n15284 , n1756 , n4464 );
    and g420 ( n13147 , n18239 , n11541 );
    or g421 ( n19595 , n16812 , n21688 );
    xnor g422 ( n6506 , n7239 , n4064 );
    nor g423 ( n25463 , n21222 , n26752 );
    nor g424 ( n10700 , n9244 , n6303 );
    xnor g425 ( n3440 , n8356 , n5853 );
    xnor g426 ( n18183 , n15810 , n17306 );
    and g427 ( n5542 , n20186 , n15844 );
    xnor g428 ( n18569 , n25484 , n22586 );
    xnor g429 ( n18445 , n16306 , n1857 );
    or g430 ( n14962 , n2336 , n6842 );
    and g431 ( n1606 , n103 , n16388 );
    or g432 ( n3079 , n11152 , n22880 );
    not g433 ( n20542 , n10403 );
    or g434 ( n18161 , n20020 , n448 );
    xnor g435 ( n11587 , n7494 , n19483 );
    and g436 ( n14780 , n17030 , n20547 );
    xnor g437 ( n16427 , n3375 , n8033 );
    nor g438 ( n15136 , n3603 , n455 );
    not g439 ( n23400 , n5648 );
    xnor g440 ( n10970 , n8043 , n26699 );
    xnor g441 ( n18213 , n24506 , n1681 );
    xnor g442 ( n3880 , n5767 , n22440 );
    and g443 ( n25111 , n1474 , n3032 );
    xnor g444 ( n17131 , n19674 , n5131 );
    xnor g445 ( n16456 , n22820 , n8244 );
    or g446 ( n24544 , n25564 , n25390 );
    nor g447 ( n11338 , n20826 , n835 );
    nor g448 ( n8949 , n2559 , n26255 );
    xnor g449 ( n10910 , n7351 , n6464 );
    or g450 ( n25894 , n24680 , n4931 );
    or g451 ( n5395 , n7597 , n17156 );
    or g452 ( n19587 , n21035 , n9696 );
    or g453 ( n14169 , n9439 , n24624 );
    and g454 ( n22303 , n16708 , n10518 );
    and g455 ( n4928 , n774 , n25145 );
    xnor g456 ( n17305 , n23966 , n18770 );
    and g457 ( n7191 , n23312 , n18920 );
    or g458 ( n23574 , n12522 , n12674 );
    or g459 ( n22163 , n6565 , n12310 );
    nor g460 ( n23479 , n24890 , n19150 );
    or g461 ( n20448 , n22675 , n15810 );
    not g462 ( n2168 , n6911 );
    or g463 ( n21360 , n3009 , n24031 );
    and g464 ( n17018 , n9988 , n21667 );
    or g465 ( n1740 , n18598 , n20946 );
    and g466 ( n10444 , n17230 , n26747 );
    xnor g467 ( n7118 , n3556 , n21434 );
    or g468 ( n7148 , n26224 , n8672 );
    xnor g469 ( n3935 , n11486 , n20138 );
    not g470 ( n1646 , n12380 );
    or g471 ( n20003 , n3458 , n2001 );
    and g472 ( n13362 , n13730 , n18019 );
    xnor g473 ( n2238 , n2925 , n5810 );
    or g474 ( n16322 , n201 , n15877 );
    or g475 ( n9444 , n1269 , n18416 );
    and g476 ( n18774 , n17846 , n12488 );
    or g477 ( n1101 , n1979 , n16245 );
    xnor g478 ( n21509 , n8942 , n15516 );
    and g479 ( n19038 , n10379 , n13772 );
    or g480 ( n17925 , n11228 , n10821 );
    not g481 ( n19464 , n12767 );
    or g482 ( n12403 , n1216 , n26887 );
    and g483 ( n25257 , n10092 , n11477 );
    nor g484 ( n7747 , n8285 , n20036 );
    not g485 ( n7325 , n477 );
    xnor g486 ( n18924 , n22587 , n16681 );
    or g487 ( n1514 , n1151 , n16111 );
    not g488 ( n13156 , n17108 );
    and g489 ( n232 , n26859 , n8590 );
    nor g490 ( n6936 , n1252 , n6204 );
    xnor g491 ( n23454 , n17552 , n7337 );
    or g492 ( n11500 , n26188 , n10652 );
    or g493 ( n20237 , n26508 , n20945 );
    not g494 ( n4896 , n22455 );
    and g495 ( n26846 , n19052 , n16826 );
    nor g496 ( n3096 , n19616 , n18558 );
    nor g497 ( n12162 , n747 , n20164 );
    or g498 ( n10363 , n24089 , n1233 );
    or g499 ( n9482 , n15408 , n19158 );
    or g500 ( n5859 , n20291 , n27027 );
    xnor g501 ( n3739 , n7853 , n22407 );
    or g502 ( n14253 , n26778 , n22520 );
    nor g503 ( n225 , n15519 , n5924 );
    and g504 ( n4113 , n18975 , n8411 );
    or g505 ( n19800 , n13741 , n3841 );
    xnor g506 ( n21602 , n23304 , n17069 );
    or g507 ( n25207 , n5557 , n23013 );
    xnor g508 ( n3850 , n6410 , n17651 );
    or g509 ( n5464 , n13591 , n24156 );
    nor g510 ( n26704 , n21974 , n20437 );
    xnor g511 ( n15737 , n11898 , n23166 );
    or g512 ( n25725 , n15338 , n20280 );
    xnor g513 ( n17119 , n397 , n26076 );
    or g514 ( n6801 , n12055 , n25855 );
    and g515 ( n14122 , n19243 , n9776 );
    and g516 ( n26138 , n16582 , n8945 );
    not g517 ( n18262 , n13112 );
    xnor g518 ( n9274 , n11202 , n15304 );
    xnor g519 ( n2785 , n1831 , n10250 );
    or g520 ( n16188 , n2724 , n9399 );
    not g521 ( n11215 , n2898 );
    xnor g522 ( n2240 , n2908 , n17771 );
    xnor g523 ( n7857 , n9825 , n133 );
    xnor g524 ( n6799 , n23254 , n6204 );
    and g525 ( n5666 , n19682 , n7041 );
    xnor g526 ( n15521 , n532 , n18272 );
    nor g527 ( n20666 , n2980 , n4781 );
    not g528 ( n26807 , n8518 );
    or g529 ( n24657 , n14510 , n8994 );
    or g530 ( n22100 , n22554 , n1414 );
    or g531 ( n18392 , n1424 , n6810 );
    not g532 ( n18539 , n13133 );
    and g533 ( n3667 , n25013 , n25965 );
    not g534 ( n14085 , n13538 );
    or g535 ( n6110 , n17447 , n22380 );
    and g536 ( n21752 , n20520 , n2859 );
    not g537 ( n3034 , n1947 );
    nor g538 ( n7382 , n21235 , n19241 );
    nor g539 ( n9956 , n11393 , n19875 );
    and g540 ( n15913 , n7593 , n17415 );
    or g541 ( n8708 , n3206 , n21931 );
    and g542 ( n19240 , n20698 , n3157 );
    xnor g543 ( n20611 , n11308 , n26205 );
    nor g544 ( n14714 , n22660 , n26823 );
    xnor g545 ( n16834 , n3250 , n22831 );
    or g546 ( n5459 , n24942 , n8789 );
    or g547 ( n4030 , n18290 , n26888 );
    or g548 ( n25477 , n13381 , n10063 );
    xnor g549 ( n1603 , n22322 , n468 );
    and g550 ( n6488 , n23974 , n26085 );
    and g551 ( n2806 , n14328 , n5720 );
    or g552 ( n24689 , n9091 , n1607 );
    nor g553 ( n26833 , n17250 , n10125 );
    or g554 ( n9203 , n5484 , n18484 );
    and g555 ( n26152 , n8273 , n3292 );
    nor g556 ( n19650 , n27074 , n19391 );
    nor g557 ( n25800 , n17660 , n1704 );
    not g558 ( n7691 , n2612 );
    or g559 ( n3688 , n19002 , n18340 );
    or g560 ( n9614 , n1319 , n3769 );
    and g561 ( n26039 , n11816 , n24954 );
    and g562 ( n17332 , n2449 , n19470 );
    xnor g563 ( n16274 , n18426 , n25168 );
    and g564 ( n15806 , n15167 , n20948 );
    nor g565 ( n22389 , n4718 , n16715 );
    or g566 ( n8412 , n23076 , n18950 );
    or g567 ( n6997 , n11732 , n13219 );
    not g568 ( n26673 , n24278 );
    xnor g569 ( n26193 , n10676 , n5556 );
    not g570 ( n2525 , n7426 );
    or g571 ( n17375 , n3975 , n22303 );
    or g572 ( n3657 , n14409 , n7806 );
    xnor g573 ( n21627 , n4466 , n15346 );
    and g574 ( n18904 , n2576 , n1325 );
    and g575 ( n10510 , n14571 , n26818 );
    or g576 ( n5118 , n16623 , n26060 );
    xnor g577 ( n13581 , n25043 , n25612 );
    or g578 ( n25828 , n3811 , n17139 );
    or g579 ( n6424 , n26036 , n1505 );
    or g580 ( n3129 , n22585 , n8680 );
    xnor g581 ( n4202 , n1466 , n7996 );
    xnor g582 ( n14243 , n23089 , n12877 );
    or g583 ( n10310 , n26506 , n26248 );
    and g584 ( n1476 , n13598 , n3467 );
    xnor g585 ( n19386 , n11003 , n22721 );
    and g586 ( n25874 , n9158 , n10223 );
    not g587 ( n18258 , n462 );
    xnor g588 ( n11632 , n23591 , n24690 );
    xnor g589 ( n6741 , n21839 , n19282 );
    and g590 ( n14247 , n21761 , n26083 );
    nor g591 ( n14099 , n5145 , n25486 );
    not g592 ( n19841 , n1986 );
    nor g593 ( n22877 , n11321 , n8933 );
    nor g594 ( n6243 , n20937 , n13435 );
    nor g595 ( n2746 , n23529 , n20700 );
    xnor g596 ( n3199 , n17090 , n6773 );
    xnor g597 ( n18446 , n701 , n23960 );
    xnor g598 ( n24554 , n1220 , n13573 );
    not g599 ( n1675 , n4768 );
    xnor g600 ( n12630 , n15073 , n15827 );
    or g601 ( n20091 , n21846 , n22861 );
    and g602 ( n2293 , n13978 , n21332 );
    not g603 ( n14155 , n15490 );
    or g604 ( n5198 , n1811 , n13994 );
    or g605 ( n27035 , n921 , n10590 );
    xnor g606 ( n15481 , n5116 , n15617 );
    or g607 ( n13127 , n21485 , n6445 );
    xnor g608 ( n16295 , n19606 , n13735 );
    xnor g609 ( n18683 , n17430 , n23852 );
    xnor g610 ( n560 , n16502 , n21654 );
    or g611 ( n4027 , n14860 , n7030 );
    not g612 ( n2281 , n8084 );
    xnor g613 ( n17372 , n8773 , n11476 );
    or g614 ( n12389 , n24990 , n22321 );
    xnor g615 ( n24155 , n21220 , n11987 );
    or g616 ( n74 , n729 , n25813 );
    not g617 ( n3681 , n25738 );
    or g618 ( n20753 , n21828 , n7177 );
    xnor g619 ( n9175 , n1405 , n9067 );
    xnor g620 ( n12556 , n21915 , n7674 );
    nor g621 ( n18625 , n3485 , n24070 );
    nor g622 ( n19205 , n6369 , n3164 );
    or g623 ( n1668 , n5809 , n25176 );
    or g624 ( n15211 , n10944 , n720 );
    not g625 ( n4844 , n24618 );
    not g626 ( n20506 , n4375 );
    buf g627 ( n27008 , n11070 );
    not g628 ( n9671 , n23586 );
    nor g629 ( n23830 , n1181 , n5708 );
    not g630 ( n16420 , n21693 );
    xnor g631 ( n16612 , n3587 , n15766 );
    and g632 ( n7819 , n16745 , n12828 );
    not g633 ( n8268 , n9506 );
    or g634 ( n17673 , n3345 , n10375 );
    or g635 ( n8284 , n7057 , n16729 );
    xnor g636 ( n23763 , n23531 , n8036 );
    or g637 ( n11661 , n24437 , n21738 );
    or g638 ( n13254 , n17542 , n6185 );
    xnor g639 ( n2349 , n19911 , n24278 );
    xnor g640 ( n18489 , n12513 , n14106 );
    xnor g641 ( n6465 , n12803 , n807 );
    and g642 ( n20847 , n3079 , n20143 );
    not g643 ( n8097 , n14600 );
    nor g644 ( n25682 , n2899 , n24731 );
    or g645 ( n27040 , n5831 , n3181 );
    and g646 ( n572 , n11011 , n1019 );
    not g647 ( n8328 , n16993 );
    not g648 ( n12770 , n15808 );
    xnor g649 ( n25499 , n24871 , n7867 );
    nor g650 ( n22411 , n8675 , n26541 );
    and g651 ( n21215 , n10535 , n10172 );
    or g652 ( n24633 , n23102 , n11677 );
    or g653 ( n17169 , n22926 , n23866 );
    and g654 ( n3826 , n10402 , n22570 );
    xnor g655 ( n851 , n368 , n19925 );
    xnor g656 ( n24188 , n3003 , n17172 );
    or g657 ( n13006 , n16168 , n11757 );
    and g658 ( n24391 , n15613 , n8157 );
    and g659 ( n9675 , n17091 , n9711 );
    nor g660 ( n6800 , n20667 , n19616 );
    or g661 ( n11660 , n487 , n1919 );
    xnor g662 ( n25203 , n12871 , n20411 );
    or g663 ( n22044 , n8904 , n25978 );
    xnor g664 ( n20033 , n21445 , n10829 );
    or g665 ( n14771 , n11679 , n24509 );
    nor g666 ( n12986 , n6595 , n23681 );
    xnor g667 ( n18502 , n24897 , n24040 );
    or g668 ( n2037 , n13709 , n3302 );
    or g669 ( n17512 , n22370 , n22332 );
    or g670 ( n2671 , n24403 , n8850 );
    or g671 ( n9652 , n4722 , n6403 );
    or g672 ( n14873 , n22919 , n8794 );
    not g673 ( n11597 , n26528 );
    xnor g674 ( n13569 , n13319 , n25435 );
    nor g675 ( n22319 , n19057 , n26292 );
    and g676 ( n1931 , n20081 , n20846 );
    or g677 ( n12989 , n328 , n22173 );
    xnor g678 ( n8563 , n1494 , n13235 );
    not g679 ( n25160 , n3220 );
    not g680 ( n20284 , n6444 );
    and g681 ( n18303 , n16937 , n5488 );
    not g682 ( n22425 , n17954 );
    nor g683 ( n3052 , n25330 , n13518 );
    or g684 ( n6715 , n24992 , n22139 );
    and g685 ( n17391 , n3958 , n18354 );
    xnor g686 ( n23879 , n6561 , n19386 );
    or g687 ( n7945 , n10459 , n13243 );
    xnor g688 ( n2952 , n20138 , n9251 );
    or g689 ( n4916 , n4900 , n10215 );
    or g690 ( n19897 , n6435 , n9245 );
    not g691 ( n14671 , n1065 );
    or g692 ( n12643 , n1164 , n4388 );
    xnor g693 ( n20714 , n17536 , n11201 );
    or g694 ( n18033 , n3096 , n17775 );
    and g695 ( n1187 , n6404 , n23349 );
    and g696 ( n6905 , n17580 , n11008 );
    xnor g697 ( n17140 , n9770 , n25054 );
    and g698 ( n6033 , n8307 , n18616 );
    and g699 ( n19839 , n14341 , n10398 );
    not g700 ( n23555 , n25877 );
    xnor g701 ( n25044 , n17077 , n4256 );
    nor g702 ( n16179 , n8013 , n27147 );
    xnor g703 ( n17862 , n3338 , n20647 );
    and g704 ( n8641 , n7102 , n280 );
    nor g705 ( n26770 , n21687 , n6606 );
    and g706 ( n711 , n639 , n16132 );
    or g707 ( n8780 , n19527 , n7808 );
    or g708 ( n24124 , n23768 , n8353 );
    and g709 ( n17348 , n6104 , n19985 );
    or g710 ( n17126 , n16679 , n7341 );
    not g711 ( n9779 , n26224 );
    xnor g712 ( n15883 , n8864 , n6334 );
    xnor g713 ( n25204 , n25573 , n18592 );
    or g714 ( n25459 , n12002 , n11382 );
    xnor g715 ( n19740 , n1562 , n2422 );
    xnor g716 ( n21622 , n9611 , n24834 );
    xnor g717 ( n12967 , n199 , n8587 );
    and g718 ( n21946 , n15030 , n17231 );
    or g719 ( n2195 , n570 , n19701 );
    xnor g720 ( n14984 , n22469 , n12358 );
    or g721 ( n16123 , n11856 , n2070 );
    or g722 ( n458 , n26810 , n12797 );
    not g723 ( n16903 , n21378 );
    or g724 ( n12028 , n21063 , n7164 );
    xnor g725 ( n6727 , n2165 , n664 );
    xnor g726 ( n5795 , n1296 , n16758 );
    or g727 ( n3192 , n24974 , n7460 );
    and g728 ( n1478 , n20565 , n14644 );
    nor g729 ( n18837 , n18921 , n17926 );
    xnor g730 ( n23942 , n16578 , n3897 );
    or g731 ( n15878 , n6916 , n7160 );
    xnor g732 ( n6019 , n21793 , n3352 );
    nor g733 ( n13638 , n13443 , n6580 );
    xnor g734 ( n5246 , n19446 , n11980 );
    not g735 ( n20976 , n14484 );
    and g736 ( n25899 , n5309 , n15523 );
    xnor g737 ( n11335 , n4980 , n6436 );
    or g738 ( n17459 , n14528 , n3552 );
    or g739 ( n21110 , n5838 , n13399 );
    not g740 ( n9561 , n15242 );
    or g741 ( n24771 , n14728 , n8570 );
    nor g742 ( n6995 , n19711 , n11697 );
    or g743 ( n20195 , n24389 , n3650 );
    xnor g744 ( n18725 , n20386 , n13001 );
    xnor g745 ( n1028 , n14908 , n23405 );
    and g746 ( n12101 , n24149 , n9933 );
    or g747 ( n19846 , n2487 , n15834 );
    and g748 ( n21338 , n991 , n1659 );
    nor g749 ( n5157 , n11410 , n18706 );
    not g750 ( n1532 , n1484 );
    xnor g751 ( n6364 , n6814 , n23463 );
    or g752 ( n5909 , n12988 , n24854 );
    or g753 ( n20026 , n796 , n24197 );
    not g754 ( n24134 , n15277 );
    xnor g755 ( n25706 , n6415 , n23060 );
    nor g756 ( n10334 , n1467 , n18113 );
    nor g757 ( n22540 , n8964 , n18539 );
    or g758 ( n21086 , n2469 , n21946 );
    not g759 ( n12673 , n5768 );
    and g760 ( n24954 , n16561 , n23596 );
    nor g761 ( n6509 , n11901 , n27089 );
    or g762 ( n17480 , n2178 , n16329 );
    or g763 ( n899 , n2332 , n19532 );
    and g764 ( n14549 , n2516 , n25638 );
    not g765 ( n25989 , n11693 );
    xnor g766 ( n22225 , n4534 , n13522 );
    or g767 ( n16312 , n7026 , n21165 );
    not g768 ( n24402 , n18326 );
    xnor g769 ( n19683 , n10281 , n24638 );
    xnor g770 ( n27098 , n11481 , n23493 );
    or g771 ( n16970 , n21512 , n23988 );
    or g772 ( n11016 , n4534 , n13522 );
    or g773 ( n1546 , n8709 , n17787 );
    xnor g774 ( n16406 , n462 , n23495 );
    xnor g775 ( n2148 , n1403 , n12898 );
    or g776 ( n13241 , n4683 , n23926 );
    xnor g777 ( n7038 , n11925 , n25964 );
    xor g778 ( n11995 , n18451 , n12278 );
    xnor g779 ( n18092 , n20425 , n15170 );
    xnor g780 ( n22064 , n21073 , n3472 );
    or g781 ( n7960 , n18869 , n22548 );
    not g782 ( n5683 , n24452 );
    not g783 ( n13990 , n10133 );
    xnor g784 ( n4656 , n16722 , n8381 );
    xnor g785 ( n25225 , n17360 , n19680 );
    nor g786 ( n14051 , n2146 , n19144 );
    xnor g787 ( n4331 , n11533 , n11095 );
    or g788 ( n4084 , n2174 , n11455 );
    not g789 ( n9125 , n24121 );
    and g790 ( n23395 , n12220 , n14553 );
    and g791 ( n3854 , n6806 , n18722 );
    xnor g792 ( n19225 , n24728 , n24161 );
    or g793 ( n19329 , n5437 , n3205 );
    and g794 ( n22725 , n12644 , n18314 );
    not g795 ( n17718 , n22480 );
    xnor g796 ( n7486 , n1408 , n23643 );
    not g797 ( n9026 , n19378 );
    or g798 ( n3712 , n6936 , n19182 );
    xnor g799 ( n5636 , n23923 , n16608 );
    xnor g800 ( n107 , n11670 , n7281 );
    or g801 ( n25183 , n5185 , n18444 );
    not g802 ( n11100 , n9646 );
    and g803 ( n3180 , n4834 , n23823 );
    and g804 ( n23919 , n26687 , n25830 );
    nor g805 ( n21035 , n14680 , n20359 );
    or g806 ( n24981 , n11193 , n9135 );
    and g807 ( n8676 , n11270 , n11976 );
    and g808 ( n8645 , n20089 , n21216 );
    xnor g809 ( n23481 , n8302 , n16840 );
    not g810 ( n21071 , n16582 );
    and g811 ( n4724 , n26257 , n9205 );
    or g812 ( n8069 , n10112 , n21849 );
    or g813 ( n13966 , n10138 , n10105 );
    xor g814 ( n17553 , n8161 , n4232 );
    and g815 ( n12949 , n2685 , n26426 );
    xnor g816 ( n15662 , n13609 , n5597 );
    nor g817 ( n15601 , n22101 , n17553 );
    xnor g818 ( n10094 , n9770 , n24612 );
    xnor g819 ( n22156 , n17982 , n8028 );
    or g820 ( n14922 , n3909 , n17045 );
    not g821 ( n15380 , n10642 );
    not g822 ( n4061 , n3018 );
    or g823 ( n12077 , n3664 , n21830 );
    not g824 ( n20749 , n12658 );
    xnor g825 ( n25670 , n744 , n13714 );
    xnor g826 ( n15547 , n15834 , n22433 );
    or g827 ( n11279 , n1151 , n20536 );
    xnor g828 ( n5273 , n7789 , n8871 );
    nor g829 ( n23159 , n5440 , n11503 );
    xnor g830 ( n6671 , n10724 , n24965 );
    not g831 ( n20862 , n17640 );
    xnor g832 ( n14949 , n4652 , n1573 );
    or g833 ( n15699 , n14153 , n21894 );
    not g834 ( n16727 , n21850 );
    and g835 ( n22963 , n987 , n11871 );
    not g836 ( n12789 , n18690 );
    and g837 ( n13470 , n25295 , n25774 );
    or g838 ( n6114 , n4339 , n6286 );
    and g839 ( n8892 , n8917 , n24753 );
    or g840 ( n2702 , n4733 , n7497 );
    or g841 ( n26976 , n11877 , n21824 );
    and g842 ( n21903 , n15886 , n5459 );
    and g843 ( n16568 , n21822 , n2462 );
    nor g844 ( n4942 , n7134 , n9830 );
    or g845 ( n5995 , n8218 , n3854 );
    xnor g846 ( n20932 , n14899 , n7026 );
    or g847 ( n4110 , n10659 , n23586 );
    xnor g848 ( n25869 , n17028 , n18444 );
    xnor g849 ( n4647 , n10760 , n801 );
    not g850 ( n17368 , n1279 );
    and g851 ( n22246 , n6282 , n15387 );
    or g852 ( n21033 , n7286 , n12030 );
    or g853 ( n4291 , n9294 , n4319 );
    or g854 ( n5390 , n4159 , n14776 );
    xnor g855 ( n10943 , n17882 , n10456 );
    xnor g856 ( n12801 , n24380 , n17476 );
    nor g857 ( n26592 , n23581 , n4572 );
    or g858 ( n9389 , n10768 , n17821 );
    xnor g859 ( n7010 , n14911 , n20494 );
    or g860 ( n24522 , n15905 , n14996 );
    xnor g861 ( n5840 , n1210 , n21579 );
    xnor g862 ( n17244 , n19608 , n4426 );
    or g863 ( n17396 , n1845 , n7169 );
    or g864 ( n11334 , n15902 , n23605 );
    xnor g865 ( n20361 , n6680 , n7667 );
    and g866 ( n6353 , n18141 , n8870 );
    xnor g867 ( n6210 , n21740 , n12547 );
    xnor g868 ( n15607 , n11533 , n4100 );
    not g869 ( n22919 , n1681 );
    xnor g870 ( n21030 , n26414 , n3506 );
    not g871 ( n26758 , n13369 );
    xnor g872 ( n17833 , n9125 , n22472 );
    and g873 ( n239 , n19829 , n18441 );
    xnor g874 ( n10035 , n14040 , n8477 );
    not g875 ( n24734 , n5944 );
    and g876 ( n16181 , n14962 , n26308 );
    xnor g877 ( n9748 , n4817 , n25605 );
    not g878 ( n21260 , n22472 );
    or g879 ( n21461 , n24299 , n630 );
    not g880 ( n19852 , n23657 );
    and g881 ( n14697 , n7522 , n18824 );
    and g882 ( n287 , n4460 , n25217 );
    or g883 ( n17377 , n3545 , n25889 );
    not g884 ( n15257 , n13318 );
    and g885 ( n10744 , n8455 , n24835 );
    or g886 ( n19964 , n2287 , n26176 );
    xnor g887 ( n22106 , n25565 , n24374 );
    and g888 ( n13246 , n1463 , n17053 );
    xnor g889 ( n20023 , n2539 , n1279 );
    and g890 ( n14535 , n7294 , n8171 );
    or g891 ( n15354 , n12996 , n19196 );
    xnor g892 ( n18462 , n14440 , n17911 );
    or g893 ( n453 , n13653 , n25051 );
    not g894 ( n15017 , n20633 );
    not g895 ( n17310 , n281 );
    xnor g896 ( n3792 , n7841 , n9445 );
    not g897 ( n9462 , n7473 );
    not g898 ( n17816 , n790 );
    or g899 ( n5083 , n6096 , n278 );
    not g900 ( n5113 , n3097 );
    or g901 ( n6454 , n10025 , n24456 );
    not g902 ( n22527 , n22173 );
    not g903 ( n24839 , n5178 );
    not g904 ( n23528 , n8721 );
    xnor g905 ( n20308 , n11764 , n26946 );
    xor g906 ( n8402 , n1583 , n1648 );
    xnor g907 ( n23624 , n7016 , n7729 );
    xnor g908 ( n14872 , n12052 , n19590 );
    xnor g909 ( n9454 , n20138 , n19494 );
    and g910 ( n23362 , n12513 , n8395 );
    xnor g911 ( n2850 , n27064 , n25850 );
    and g912 ( n8407 , n25108 , n7064 );
    or g913 ( n10933 , n13695 , n26056 );
    or g914 ( n22141 , n23004 , n14913 );
    xnor g915 ( n18068 , n6377 , n987 );
    or g916 ( n20232 , n8071 , n26851 );
    and g917 ( n18159 , n136 , n15982 );
    nor g918 ( n19535 , n10167 , n24104 );
    or g919 ( n7329 , n9979 , n1227 );
    or g920 ( n18026 , n18705 , n8083 );
    xnor g921 ( n8589 , n7375 , n5454 );
    and g922 ( n18472 , n12732 , n15250 );
    xnor g923 ( n11647 , n22543 , n4540 );
    and g924 ( n20820 , n9289 , n17309 );
    xnor g925 ( n2565 , n13930 , n6105 );
    not g926 ( n26661 , n24732 );
    or g927 ( n1736 , n13278 , n23372 );
    and g928 ( n12513 , n24249 , n3058 );
    xnor g929 ( n17078 , n15490 , n7339 );
    or g930 ( n6332 , n26892 , n11623 );
    xnor g931 ( n25144 , n3952 , n12315 );
    or g932 ( n14079 , n9964 , n5067 );
    and g933 ( n18849 , n25324 , n5951 );
    nor g934 ( n12893 , n10763 , n5696 );
    xnor g935 ( n17865 , n6726 , n22934 );
    or g936 ( n19023 , n26661 , n19371 );
    nor g937 ( n5825 , n9180 , n8006 );
    nor g938 ( n1242 , n23692 , n15236 );
    xnor g939 ( n280 , n2855 , n2002 );
    not g940 ( n10804 , n7284 );
    and g941 ( n17297 , n21641 , n7383 );
    not g942 ( n25389 , n12562 );
    or g943 ( n4638 , n17162 , n868 );
    or g944 ( n15485 , n5371 , n22539 );
    xnor g945 ( n5561 , n13328 , n16439 );
    or g946 ( n8183 , n4210 , n17628 );
    xnor g947 ( n11379 , n24584 , n6873 );
    not g948 ( n7347 , n8858 );
    or g949 ( n7508 , n2098 , n606 );
    nor g950 ( n12682 , n3540 , n10885 );
    nor g951 ( n22781 , n8520 , n18338 );
    nor g952 ( n8606 , n11201 , n14366 );
    xnor g953 ( n18726 , n11575 , n16703 );
    and g954 ( n25901 , n25163 , n9354 );
    nor g955 ( n12447 , n18947 , n10331 );
    xnor g956 ( n4333 , n21638 , n7567 );
    or g957 ( n24564 , n3827 , n5055 );
    nor g958 ( n18228 , n16261 , n24188 );
    or g959 ( n16043 , n2348 , n25064 );
    or g960 ( n18470 , n23527 , n18275 );
    or g961 ( n900 , n1866 , n17656 );
    xnor g962 ( n16654 , n13441 , n13094 );
    not g963 ( n14251 , n2429 );
    nor g964 ( n22366 , n7319 , n17458 );
    not g965 ( n6400 , n21138 );
    xnor g966 ( n23251 , n25119 , n21934 );
    or g967 ( n13185 , n13674 , n14316 );
    and g968 ( n16799 , n8146 , n5285 );
    not g969 ( n26495 , n2829 );
    and g970 ( n26027 , n12811 , n11822 );
    and g971 ( n4773 , n14831 , n21415 );
    xnor g972 ( n6802 , n7140 , n26934 );
    nor g973 ( n20243 , n387 , n9300 );
    or g974 ( n6797 , n26607 , n13840 );
    xnor g975 ( n8401 , n12436 , n24937 );
    or g976 ( n13225 , n18058 , n3828 );
    or g977 ( n2641 , n18527 , n1991 );
    not g978 ( n16331 , n1320 );
    xnor g979 ( n849 , n2221 , n26917 );
    and g980 ( n19735 , n13430 , n1056 );
    or g981 ( n24534 , n8134 , n27005 );
    and g982 ( n22846 , n10195 , n14889 );
    nor g983 ( n16591 , n19474 , n151 );
    or g984 ( n1814 , n6686 , n2163 );
    xnor g985 ( n4051 , n25068 , n6790 );
    or g986 ( n11288 , n4586 , n3381 );
    or g987 ( n18244 , n21841 , n14110 );
    and g988 ( n14357 , n20167 , n19826 );
    nor g989 ( n15439 , n19110 , n5467 );
    or g990 ( n26690 , n4398 , n12694 );
    nor g991 ( n3652 , n2424 , n84 );
    not g992 ( n17835 , n31 );
    or g993 ( n22466 , n20918 , n7874 );
    or g994 ( n6825 , n13731 , n6195 );
    and g995 ( n5078 , n2762 , n17868 );
    not g996 ( n5585 , n837 );
    not g997 ( n8835 , n1878 );
    xnor g998 ( n17519 , n20671 , n26963 );
    or g999 ( n26401 , n19260 , n8830 );
    nor g1000 ( n777 , n5498 , n12928 );
    not g1001 ( n172 , n6988 );
    not g1002 ( n20552 , n22918 );
    xnor g1003 ( n22828 , n23186 , n24047 );
    xnor g1004 ( n20215 , n6389 , n14350 );
    not g1005 ( n15773 , n18569 );
    or g1006 ( n2874 , n10710 , n26510 );
    and g1007 ( n1707 , n23922 , n2843 );
    nor g1008 ( n13017 , n19094 , n1197 );
    not g1009 ( n12464 , n26823 );
    or g1010 ( n1856 , n15329 , n7528 );
    not g1011 ( n12888 , n25017 );
    or g1012 ( n12590 , n19568 , n162 );
    xnor g1013 ( n5048 , n7383 , n19576 );
    nor g1014 ( n22566 , n12573 , n19312 );
    xnor g1015 ( n23534 , n18035 , n3279 );
    not g1016 ( n27142 , n6230 );
    and g1017 ( n18230 , n3874 , n1485 );
    not g1018 ( n20094 , n21567 );
    or g1019 ( n18803 , n2812 , n18812 );
    nor g1020 ( n16128 , n658 , n27120 );
    nor g1021 ( n25615 , n6744 , n18568 );
    xnor g1022 ( n14883 , n16856 , n21081 );
    xnor g1023 ( n26219 , n22378 , n5026 );
    not g1024 ( n17015 , n23765 );
    xnor g1025 ( n24335 , n24511 , n10096 );
    and g1026 ( n19400 , n5303 , n7508 );
    xnor g1027 ( n4935 , n23832 , n3161 );
    or g1028 ( n12312 , n11270 , n11976 );
    xnor g1029 ( n4861 , n1426 , n12419 );
    not g1030 ( n166 , n19080 );
    nor g1031 ( n8196 , n2979 , n9554 );
    xnor g1032 ( n6044 , n1564 , n2050 );
    xnor g1033 ( n6550 , n12422 , n1780 );
    or g1034 ( n27097 , n3021 , n16308 );
    xnor g1035 ( n26174 , n24668 , n23671 );
    xnor g1036 ( n1885 , n15090 , n12209 );
    xnor g1037 ( n4693 , n4907 , n1012 );
    xnor g1038 ( n6914 , n10405 , n25370 );
    xnor g1039 ( n6662 , n22153 , n3984 );
    or g1040 ( n19397 , n13058 , n7749 );
    or g1041 ( n24492 , n7195 , n12861 );
    nor g1042 ( n7683 , n9498 , n12494 );
    not g1043 ( n10331 , n21444 );
    and g1044 ( n4700 , n21730 , n18464 );
    xnor g1045 ( n25181 , n12450 , n5876 );
    and g1046 ( n24334 , n24885 , n20381 );
    or g1047 ( n8129 , n19444 , n20689 );
    not g1048 ( n5923 , n10735 );
    nor g1049 ( n18929 , n12475 , n18263 );
    xnor g1050 ( n20959 , n1365 , n10158 );
    and g1051 ( n24064 , n23703 , n2344 );
    and g1052 ( n11270 , n8436 , n4886 );
    xnor g1053 ( n2711 , n2375 , n6453 );
    and g1054 ( n7856 , n14307 , n6629 );
    and g1055 ( n23275 , n17486 , n25662 );
    nor g1056 ( n22030 , n12112 , n20444 );
    and g1057 ( n3168 , n5137 , n9762 );
    and g1058 ( n798 , n25090 , n3182 );
    and g1059 ( n7431 , n27006 , n7197 );
    or g1060 ( n26938 , n14559 , n4290 );
    xnor g1061 ( n9388 , n18398 , n1605 );
    or g1062 ( n10528 , n9857 , n27148 );
    and g1063 ( n24436 , n21153 , n11907 );
    xnor g1064 ( n17667 , n13490 , n7751 );
    not g1065 ( n598 , n25360 );
    xnor g1066 ( n12449 , n11969 , n25279 );
    or g1067 ( n13750 , n7191 , n25697 );
    or g1068 ( n1256 , n16049 , n18199 );
    not g1069 ( n7615 , n20183 );
    xnor g1070 ( n26856 , n12861 , n1255 );
    and g1071 ( n13661 , n25354 , n16936 );
    and g1072 ( n15552 , n36 , n23127 );
    xnor g1073 ( n15314 , n14774 , n23200 );
    not g1074 ( n6011 , n3274 );
    nor g1075 ( n15192 , n8230 , n10454 );
    and g1076 ( n17134 , n6880 , n775 );
    and g1077 ( n15631 , n329 , n6541 );
    and g1078 ( n13527 , n23852 , n17430 );
    or g1079 ( n16442 , n3043 , n3861 );
    and g1080 ( n3900 , n15734 , n18664 );
    xnor g1081 ( n19762 , n556 , n26348 );
    or g1082 ( n6009 , n19804 , n14311 );
    and g1083 ( n194 , n14775 , n14925 );
    nor g1084 ( n4301 , n8739 , n23655 );
    nor g1085 ( n20300 , n15942 , n17499 );
    xnor g1086 ( n8406 , n27128 , n12275 );
    xnor g1087 ( n21963 , n7330 , n2479 );
    and g1088 ( n14340 , n25722 , n16004 );
    xnor g1089 ( n11325 , n8341 , n4443 );
    xnor g1090 ( n2481 , n5130 , n24419 );
    nor g1091 ( n13903 , n23459 , n10603 );
    xnor g1092 ( n11512 , n26875 , n5530 );
    or g1093 ( n17860 , n12143 , n20215 );
    or g1094 ( n10907 , n5501 , n23824 );
    or g1095 ( n9884 , n2453 , n26318 );
    or g1096 ( n14188 , n22167 , n11373 );
    not g1097 ( n25238 , n13774 );
    xnor g1098 ( n26552 , n16653 , n16558 );
    xnor g1099 ( n8242 , n7439 , n15182 );
    or g1100 ( n9868 , n12822 , n10231 );
    or g1101 ( n3073 , n12368 , n14670 );
    or g1102 ( n62 , n14542 , n23147 );
    or g1103 ( n16438 , n19097 , n5333 );
    xnor g1104 ( n21210 , n2085 , n21361 );
    xnor g1105 ( n5082 , n25807 , n9388 );
    not g1106 ( n9335 , n19544 );
    nor g1107 ( n20684 , n337 , n17902 );
    xnor g1108 ( n12281 , n25056 , n23192 );
    not g1109 ( n11193 , n9940 );
    or g1110 ( n993 , n16152 , n1377 );
    and g1111 ( n1530 , n22072 , n7529 );
    or g1112 ( n11727 , n18218 , n7430 );
    or g1113 ( n26398 , n4119 , n24746 );
    not g1114 ( n21668 , n9575 );
    not g1115 ( n9310 , n1525 );
    xnor g1116 ( n15985 , n5124 , n14675 );
    or g1117 ( n15384 , n752 , n4105 );
    xnor g1118 ( n20144 , n10191 , n23279 );
    or g1119 ( n26242 , n1179 , n6579 );
    and g1120 ( n13121 , n15347 , n1774 );
    and g1121 ( n10892 , n22236 , n3399 );
    nor g1122 ( n22420 , n494 , n17141 );
    xnor g1123 ( n6001 , n20777 , n13848 );
    nor g1124 ( n3155 , n9586 , n24196 );
    or g1125 ( n22757 , n1771 , n17033 );
    not g1126 ( n2423 , n161 );
    or g1127 ( n18835 , n5206 , n2937 );
    xnor g1128 ( n12484 , n16091 , n16602 );
    xnor g1129 ( n22496 , n17536 , n19060 );
    xnor g1130 ( n26835 , n24473 , n19472 );
    and g1131 ( n426 , n4514 , n21162 );
    or g1132 ( n10297 , n1870 , n18701 );
    xnor g1133 ( n21497 , n12379 , n1434 );
    and g1134 ( n1323 , n2414 , n5754 );
    xnor g1135 ( n10699 , n4724 , n6418 );
    nor g1136 ( n20142 , n18639 , n20771 );
    or g1137 ( n2012 , n3018 , n16366 );
    or g1138 ( n11310 , n786 , n24281 );
    xnor g1139 ( n16026 , n7619 , n16446 );
    xnor g1140 ( n6575 , n18754 , n5211 );
    not g1141 ( n16333 , n1601 );
    xnor g1142 ( n9160 , n19507 , n17798 );
    and g1143 ( n25760 , n3403 , n3271 );
    not g1144 ( n26023 , n8164 );
    xnor g1145 ( n7387 , n14741 , n25454 );
    nor g1146 ( n6120 , n1525 , n11018 );
    or g1147 ( n10957 , n7523 , n8385 );
    not g1148 ( n18205 , n10963 );
    and g1149 ( n21864 , n5174 , n24336 );
    and g1150 ( n10153 , n15290 , n25734 );
    or g1151 ( n23945 , n23144 , n10306 );
    and g1152 ( n8151 , n4939 , n120 );
    not g1153 ( n26999 , n5206 );
    xnor g1154 ( n12907 , n24493 , n22198 );
    and g1155 ( n686 , n9905 , n20174 );
    or g1156 ( n8586 , n22964 , n19924 );
    and g1157 ( n11672 , n12017 , n8169 );
    xnor g1158 ( n16393 , n10523 , n25203 );
    nor g1159 ( n7141 , n1896 , n27104 );
    or g1160 ( n2496 , n15911 , n26939 );
    xnor g1161 ( n11593 , n11840 , n15423 );
    or g1162 ( n6075 , n26450 , n22958 );
    or g1163 ( n5928 , n6268 , n1218 );
    and g1164 ( n16702 , n7322 , n15689 );
    or g1165 ( n16754 , n19432 , n11337 );
    or g1166 ( n2865 , n13274 , n8524 );
    xnor g1167 ( n18177 , n2035 , n26054 );
    xnor g1168 ( n16752 , n26974 , n10305 );
    or g1169 ( n19855 , n19018 , n20910 );
    or g1170 ( n15263 , n20303 , n14598 );
    or g1171 ( n24438 , n4539 , n368 );
    xnor g1172 ( n23698 , n4963 , n24796 );
    or g1173 ( n19942 , n15989 , n7665 );
    xnor g1174 ( n22881 , n6122 , n678 );
    xnor g1175 ( n1302 , n10891 , n10367 );
    nor g1176 ( n22959 , n16163 , n15932 );
    nor g1177 ( n25752 , n24902 , n25572 );
    and g1178 ( n17289 , n4164 , n9865 );
    xnor g1179 ( n22852 , n9615 , n21055 );
    not g1180 ( n17210 , n563 );
    and g1181 ( n19180 , n27088 , n10031 );
    or g1182 ( n22965 , n23490 , n15048 );
    or g1183 ( n10132 , n751 , n14788 );
    or g1184 ( n21546 , n22534 , n12577 );
    or g1185 ( n22893 , n3769 , n4485 );
    xnor g1186 ( n5732 , n8346 , n6344 );
    xnor g1187 ( n6142 , n24480 , n14634 );
    and g1188 ( n20121 , n11246 , n14974 );
    or g1189 ( n18391 , n13709 , n15696 );
    nor g1190 ( n26766 , n1398 , n20548 );
    xnor g1191 ( n10878 , n8679 , n14516 );
    or g1192 ( n3597 , n25470 , n3307 );
    and g1193 ( n9632 , n3849 , n10750 );
    not g1194 ( n10207 , n16197 );
    or g1195 ( n20514 , n15326 , n21875 );
    nor g1196 ( n7462 , n18537 , n4376 );
    not g1197 ( n5506 , n5288 );
    not g1198 ( n1798 , n23337 );
    nor g1199 ( n3648 , n22795 , n2100 );
    or g1200 ( n25633 , n25428 , n22412 );
    and g1201 ( n19370 , n10290 , n3824 );
    or g1202 ( n20511 , n14415 , n8032 );
    xnor g1203 ( n10644 , n3967 , n27054 );
    and g1204 ( n8438 , n14764 , n13836 );
    and g1205 ( n1608 , n4344 , n13849 );
    xnor g1206 ( n18736 , n14795 , n14189 );
    nor g1207 ( n24709 , n19454 , n15042 );
    nor g1208 ( n26042 , n1192 , n5743 );
    not g1209 ( n22977 , n21 );
    xnor g1210 ( n26784 , n12944 , n6864 );
    xnor g1211 ( n20269 , n18444 , n13719 );
    and g1212 ( n15738 , n26299 , n25208 );
    or g1213 ( n9613 , n3648 , n5405 );
    and g1214 ( n1285 , n667 , n15372 );
    xnor g1215 ( n8821 , n25583 , n15286 );
    xnor g1216 ( n3979 , n2783 , n1667 );
    not g1217 ( n17156 , n24009 );
    xnor g1218 ( n7476 , n16330 , n14597 );
    and g1219 ( n18286 , n27080 , n24515 );
    or g1220 ( n1985 , n12024 , n18622 );
    and g1221 ( n10082 , n23945 , n21411 );
    nor g1222 ( n22589 , n14829 , n21889 );
    not g1223 ( n22349 , n3143 );
    and g1224 ( n9976 , n4733 , n7497 );
    and g1225 ( n12165 , n16869 , n14908 );
    or g1226 ( n1317 , n23873 , n21726 );
    or g1227 ( n10395 , n25038 , n12639 );
    and g1228 ( n14066 , n13795 , n17404 );
    not g1229 ( n2566 , n24072 );
    or g1230 ( n9836 , n15766 , n3587 );
    nor g1231 ( n22179 , n21226 , n2906 );
    and g1232 ( n25019 , n7166 , n9271 );
    xnor g1233 ( n8383 , n21134 , n11356 );
    xnor g1234 ( n7638 , n7170 , n24606 );
    or g1235 ( n13160 , n22942 , n712 );
    xnor g1236 ( n3492 , n17369 , n26512 );
    xnor g1237 ( n11905 , n3913 , n8140 );
    or g1238 ( n26732 , n23089 , n9830 );
    not g1239 ( n24031 , n7674 );
    xnor g1240 ( n22467 , n3631 , n14493 );
    or g1241 ( n14918 , n25434 , n22086 );
    xnor g1242 ( n1446 , n9542 , n12773 );
    and g1243 ( n5217 , n15493 , n21345 );
    and g1244 ( n4493 , n25923 , n24184 );
    nor g1245 ( n25326 , n21134 , n11356 );
    and g1246 ( n12344 , n14813 , n16863 );
    or g1247 ( n13942 , n7012 , n24830 );
    xnor g1248 ( n6747 , n10486 , n19584 );
    not g1249 ( n1554 , n23523 );
    xnor g1250 ( n13387 , n20957 , n21897 );
    and g1251 ( n15219 , n12284 , n363 );
    xnor g1252 ( n17084 , n9304 , n6345 );
    and g1253 ( n26662 , n5783 , n11432 );
    or g1254 ( n14012 , n22743 , n2346 );
    not g1255 ( n26022 , n14031 );
    xnor g1256 ( n13934 , n3770 , n24801 );
    or g1257 ( n27176 , n26211 , n15333 );
    or g1258 ( n19405 , n8285 , n14480 );
    xnor g1259 ( n794 , n11235 , n10352 );
    and g1260 ( n25723 , n21805 , n13937 );
    xnor g1261 ( n21402 , n19005 , n19144 );
    nor g1262 ( n20918 , n10629 , n6660 );
    and g1263 ( n2206 , n1948 , n16250 );
    not g1264 ( n24379 , n15141 );
    or g1265 ( n26041 , n15625 , n2049 );
    not g1266 ( n18431 , n17663 );
    not g1267 ( n14336 , n22433 );
    xnor g1268 ( n2515 , n5027 , n21335 );
    not g1269 ( n2782 , n4520 );
    or g1270 ( n12260 , n24903 , n26466 );
    nor g1271 ( n19611 , n19594 , n6235 );
    or g1272 ( n11464 , n16784 , n15500 );
    not g1273 ( n26894 , n20171 );
    or g1274 ( n250 , n27062 , n12805 );
    not g1275 ( n21465 , n18809 );
    not g1276 ( n2003 , n13291 );
    xnor g1277 ( n9468 , n22875 , n5813 );
    xnor g1278 ( n21180 , n23264 , n27120 );
    nor g1279 ( n4500 , n4031 , n24560 );
    not g1280 ( n9599 , n22780 );
    not g1281 ( n17062 , n25483 );
    xnor g1282 ( n6436 , n8241 , n11566 );
    xnor g1283 ( n22136 , n9748 , n6915 );
    and g1284 ( n9874 , n11464 , n16425 );
    or g1285 ( n24915 , n8999 , n1122 );
    xnor g1286 ( n1859 , n14112 , n22639 );
    nor g1287 ( n5772 , n15294 , n15270 );
    and g1288 ( n23654 , n6651 , n12037 );
    or g1289 ( n4390 , n8186 , n3425 );
    xnor g1290 ( n6567 , n22551 , n6020 );
    and g1291 ( n9305 , n22860 , n21494 );
    and g1292 ( n19384 , n7237 , n2813 );
    or g1293 ( n12948 , n26309 , n11726 );
    not g1294 ( n3985 , n1610 );
    nor g1295 ( n17678 , n14048 , n4467 );
    or g1296 ( n23011 , n16302 , n2489 );
    xnor g1297 ( n24151 , n26249 , n4129 );
    xnor g1298 ( n22633 , n21849 , n5954 );
    or g1299 ( n7307 , n6411 , n5649 );
    xnor g1300 ( n75 , n10702 , n12776 );
    xnor g1301 ( n14211 , n6188 , n17117 );
    xnor g1302 ( n11048 , n25560 , n13914 );
    xnor g1303 ( n10467 , n7673 , n3176 );
    xnor g1304 ( n14196 , n19797 , n4559 );
    or g1305 ( n10670 , n1405 , n27181 );
    and g1306 ( n1084 , n15426 , n22521 );
    xnor g1307 ( n20607 , n16874 , n530 );
    and g1308 ( n11534 , n5025 , n12771 );
    not g1309 ( n25795 , n11008 );
    and g1310 ( n17257 , n26844 , n18964 );
    and g1311 ( n1216 , n23150 , n2183 );
    xnor g1312 ( n6640 , n2809 , n15508 );
    not g1313 ( n16204 , n12885 );
    and g1314 ( n23201 , n17871 , n15067 );
    or g1315 ( n20893 , n6750 , n13328 );
    and g1316 ( n26967 , n26627 , n6577 );
    and g1317 ( n2413 , n23901 , n16038 );
    or g1318 ( n8075 , n14939 , n25449 );
    and g1319 ( n7024 , n3192 , n15388 );
    xnor g1320 ( n24723 , n21553 , n7660 );
    not g1321 ( n16982 , n6003 );
    and g1322 ( n10291 , n24263 , n3608 );
    or g1323 ( n15123 , n14198 , n12902 );
    or g1324 ( n10195 , n10018 , n513 );
    and g1325 ( n5693 , n4998 , n4888 );
    and g1326 ( n26392 , n17540 , n14987 );
    or g1327 ( n10657 , n25355 , n5110 );
    nor g1328 ( n25570 , n9211 , n24394 );
    and g1329 ( n25482 , n2227 , n24079 );
    or g1330 ( n16031 , n21474 , n19865 );
    or g1331 ( n219 , n1447 , n22482 );
    or g1332 ( n2933 , n5696 , n23463 );
    not g1333 ( n16551 , n7609 );
    and g1334 ( n19807 , n13203 , n2430 );
    not g1335 ( n5790 , n24609 );
    not g1336 ( n16590 , n21509 );
    xnor g1337 ( n21352 , n12428 , n18215 );
    not g1338 ( n3687 , n18674 );
    nor g1339 ( n22462 , n1587 , n22977 );
    or g1340 ( n4637 , n20467 , n13615 );
    and g1341 ( n18314 , n11090 , n26267 );
    not g1342 ( n24601 , n3829 );
    or g1343 ( n12150 , n9906 , n22349 );
    not g1344 ( n4781 , n26403 );
    or g1345 ( n19600 , n19195 , n177 );
    not g1346 ( n11177 , n1288 );
    or g1347 ( n14062 , n25022 , n7441 );
    xnor g1348 ( n23399 , n25318 , n3955 );
    nor g1349 ( n6355 , n19839 , n6518 );
    xnor g1350 ( n3202 , n2145 , n5521 );
    xnor g1351 ( n20161 , n6032 , n13623 );
    xnor g1352 ( n20532 , n149 , n15243 );
    or g1353 ( n13624 , n9850 , n1162 );
    or g1354 ( n1496 , n14523 , n19419 );
    and g1355 ( n23571 , n23367 , n1856 );
    or g1356 ( n19212 , n2084 , n17135 );
    xnor g1357 ( n20564 , n1801 , n18906 );
    and g1358 ( n15615 , n22373 , n5009 );
    or g1359 ( n15429 , n15894 , n10560 );
    xnor g1360 ( n6560 , n7385 , n11493 );
    or g1361 ( n18979 , n6962 , n5119 );
    nor g1362 ( n10619 , n15204 , n14122 );
    nor g1363 ( n6416 , n2939 , n6366 );
    or g1364 ( n23858 , n25888 , n19149 );
    and g1365 ( n1077 , n22197 , n5927 );
    or g1366 ( n21507 , n17173 , n21644 );
    and g1367 ( n24719 , n8923 , n26175 );
    or g1368 ( n8248 , n15454 , n2171 );
    not g1369 ( n24625 , n252 );
    or g1370 ( n18602 , n10763 , n18799 );
    nor g1371 ( n7065 , n7099 , n6691 );
    or g1372 ( n17999 , n218 , n25327 );
    and g1373 ( n7985 , n5375 , n18267 );
    xnor g1374 ( n4877 , n11198 , n4391 );
    xnor g1375 ( n8637 , n3866 , n7491 );
    not g1376 ( n13033 , n18901 );
    or g1377 ( n16363 , n17676 , n25404 );
    xnor g1378 ( n16811 , n17846 , n12488 );
    nor g1379 ( n3439 , n21380 , n11592 );
    not g1380 ( n11028 , n17652 );
    xnor g1381 ( n10261 , n25145 , n14423 );
    and g1382 ( n18594 , n23234 , n1688 );
    or g1383 ( n26214 , n14920 , n8591 );
    not g1384 ( n729 , n15339 );
    xnor g1385 ( n14484 , n23493 , n8405 );
    not g1386 ( n7107 , n4448 );
    xnor g1387 ( n26729 , n9984 , n25526 );
    xnor g1388 ( n19283 , n2979 , n11898 );
    xnor g1389 ( n24872 , n23352 , n25659 );
    or g1390 ( n15040 , n6702 , n14893 );
    and g1391 ( n6056 , n6368 , n8879 );
    and g1392 ( n6058 , n21438 , n2291 );
    and g1393 ( n26550 , n20777 , n2461 );
    and g1394 ( n23625 , n21828 , n7177 );
    xnor g1395 ( n17971 , n14411 , n16983 );
    and g1396 ( n14160 , n5438 , n9964 );
    xnor g1397 ( n825 , n24908 , n23000 );
    xnor g1398 ( n24106 , n44 , n26290 );
    xnor g1399 ( n26128 , n3097 , n3764 );
    or g1400 ( n17308 , n23804 , n21422 );
    buf g1401 ( n1553 , n24440 );
    or g1402 ( n16269 , n5582 , n24842 );
    and g1403 ( n20492 , n1372 , n16414 );
    not g1404 ( n26961 , n5128 );
    xnor g1405 ( n12615 , n13367 , n13074 );
    or g1406 ( n6198 , n6946 , n11136 );
    and g1407 ( n16412 , n4802 , n25725 );
    xnor g1408 ( n9591 , n11603 , n16399 );
    and g1409 ( n2025 , n19346 , n1985 );
    xnor g1410 ( n26119 , n15264 , n19720 );
    or g1411 ( n24288 , n10700 , n23468 );
    nor g1412 ( n20875 , n6704 , n21878 );
    xnor g1413 ( n20290 , n6832 , n11898 );
    xnor g1414 ( n15972 , n20627 , n12036 );
    xnor g1415 ( n25883 , n4858 , n26752 );
    xnor g1416 ( n783 , n12622 , n26289 );
    not g1417 ( n21972 , n13783 );
    not g1418 ( n11110 , n6224 );
    or g1419 ( n1836 , n9712 , n9214 );
    xnor g1420 ( n18515 , n24507 , n12809 );
    and g1421 ( n14659 , n27116 , n10170 );
    xnor g1422 ( n18260 , n8827 , n4306 );
    or g1423 ( n3469 , n20472 , n2181 );
    not g1424 ( n5 , n5625 );
    nor g1425 ( n12459 , n10131 , n8507 );
    xnor g1426 ( n24990 , n14376 , n9608 );
    not g1427 ( n15755 , n11823 );
    xnor g1428 ( n12342 , n23395 , n8950 );
    or g1429 ( n8885 , n1403 , n16176 );
    and g1430 ( n8310 , n20290 , n21577 );
    xnor g1431 ( n15062 , n9367 , n12353 );
    xnor g1432 ( n11296 , n456 , n24479 );
    or g1433 ( n13097 , n7141 , n7654 );
    nor g1434 ( n24866 , n11229 , n17195 );
    and g1435 ( n17683 , n18604 , n4912 );
    xnor g1436 ( n11771 , n938 , n4524 );
    not g1437 ( n18196 , n4068 );
    nor g1438 ( n889 , n15217 , n14695 );
    or g1439 ( n14884 , n26918 , n18827 );
    xnor g1440 ( n27193 , n19408 , n6879 );
    nor g1441 ( n22767 , n27111 , n25265 );
    not g1442 ( n1876 , n11482 );
    and g1443 ( n4636 , n14053 , n12253 );
    not g1444 ( n4203 , n5051 );
    or g1445 ( n15987 , n13360 , n16392 );
    or g1446 ( n5799 , n2903 , n4570 );
    nor g1447 ( n17300 , n7731 , n13109 );
    and g1448 ( n14481 , n15903 , n10802 );
    and g1449 ( n21418 , n11334 , n8696 );
    xnor g1450 ( n13161 , n14695 , n15473 );
    nor g1451 ( n25510 , n23234 , n20235 );
    and g1452 ( n15172 , n19663 , n8025 );
    not g1453 ( n26134 , n10932 );
    not g1454 ( n9365 , n19234 );
    or g1455 ( n24185 , n23555 , n26443 );
    or g1456 ( n7855 , n10026 , n18432 );
    nor g1457 ( n5186 , n15409 , n1145 );
    and g1458 ( n19630 , n22729 , n18744 );
    xnor g1459 ( n3906 , n7826 , n26600 );
    xnor g1460 ( n12234 , n14723 , n24560 );
    not g1461 ( n20120 , n10908 );
    xnor g1462 ( n15902 , n12025 , n21198 );
    or g1463 ( n25011 , n19619 , n2625 );
    xnor g1464 ( n1114 , n15261 , n16902 );
    or g1465 ( n9762 , n955 , n13509 );
    or g1466 ( n4884 , n4143 , n19184 );
    not g1467 ( n21456 , n11382 );
    xnor g1468 ( n18668 , n6283 , n19081 );
    and g1469 ( n10098 , n14139 , n14838 );
    xnor g1470 ( n18006 , n5893 , n22488 );
    and g1471 ( n18417 , n7618 , n22560 );
    and g1472 ( n8340 , n17578 , n8653 );
    xnor g1473 ( n12231 , n21114 , n14477 );
    xnor g1474 ( n19836 , n3144 , n1683 );
    nor g1475 ( n6923 , n5355 , n19094 );
    xnor g1476 ( n26111 , n7656 , n24176 );
    and g1477 ( n7668 , n8468 , n24026 );
    or g1478 ( n15694 , n17602 , n8644 );
    xnor g1479 ( n19333 , n18211 , n8674 );
    nor g1480 ( n3551 , n2666 , n14739 );
    or g1481 ( n99 , n12236 , n11589 );
    or g1482 ( n5814 , n25036 , n18498 );
    xnor g1483 ( n5981 , n1267 , n12507 );
    xnor g1484 ( n10728 , n18650 , n17206 );
    not g1485 ( n9453 , n25069 );
    xnor g1486 ( n19080 , n374 , n10483 );
    nor g1487 ( n9875 , n23083 , n17858 );
    xnor g1488 ( n15058 , n7626 , n13691 );
    and g1489 ( n7772 , n19790 , n19151 );
    or g1490 ( n18507 , n3161 , n16888 );
    xnor g1491 ( n26169 , n6353 , n8434 );
    xnor g1492 ( n822 , n14743 , n2990 );
    and g1493 ( n14850 , n15789 , n261 );
    not g1494 ( n23261 , n25490 );
    not g1495 ( n663 , n26102 );
    or g1496 ( n4439 , n25759 , n25224 );
    or g1497 ( n13655 , n14840 , n12489 );
    not g1498 ( n18547 , n25594 );
    xnor g1499 ( n4618 , n10890 , n14157 );
    or g1500 ( n17570 , n26644 , n15403 );
    xnor g1501 ( n14972 , n12335 , n11148 );
    or g1502 ( n866 , n23912 , n25601 );
    and g1503 ( n10844 , n24241 , n23713 );
    or g1504 ( n3444 , n18268 , n15526 );
    xnor g1505 ( n19524 , n7397 , n14196 );
    xnor g1506 ( n21786 , n25291 , n7061 );
    xnor g1507 ( n13060 , n6164 , n22850 );
    xnor g1508 ( n25256 , n15247 , n19403 );
    nor g1509 ( n123 , n12281 , n15007 );
    not g1510 ( n26654 , n5682 );
    or g1511 ( n26779 , n3120 , n14361 );
    nor g1512 ( n27091 , n12291 , n25689 );
    or g1513 ( n11946 , n16234 , n25069 );
    not g1514 ( n6580 , n2210 );
    xnor g1515 ( n19294 , n2919 , n27037 );
    or g1516 ( n4979 , n15895 , n16222 );
    xnor g1517 ( n21424 , n9589 , n18427 );
    nor g1518 ( n4633 , n26472 , n7359 );
    and g1519 ( n16357 , n4145 , n20725 );
    or g1520 ( n1901 , n11052 , n21691 );
    and g1521 ( n14432 , n21669 , n11836 );
    or g1522 ( n17962 , n12444 , n25048 );
    or g1523 ( n416 , n17212 , n16627 );
    or g1524 ( n5489 , n17549 , n1657 );
    and g1525 ( n17552 , n15344 , n4264 );
    xnor g1526 ( n7859 , n14899 , n18496 );
    and g1527 ( n24466 , n16587 , n9501 );
    and g1528 ( n21869 , n25877 , n6393 );
    not g1529 ( n8816 , n11543 );
    nor g1530 ( n8525 , n16576 , n10581 );
    and g1531 ( n3538 , n12900 , n16547 );
    xnor g1532 ( n9451 , n22611 , n16979 );
    nor g1533 ( n11569 , n20470 , n4590 );
    xnor g1534 ( n23757 , n5413 , n2185 );
    xnor g1535 ( n227 , n22964 , n19907 );
    and g1536 ( n3242 , n3430 , n12994 );
    not g1537 ( n26316 , n19765 );
    or g1538 ( n13107 , n17981 , n7125 );
    and g1539 ( n12437 , n16022 , n1519 );
    or g1540 ( n7315 , n5432 , n12092 );
    not g1541 ( n19371 , n26808 );
    xnor g1542 ( n23861 , n12734 , n23039 );
    xnor g1543 ( n1060 , n877 , n13202 );
    nor g1544 ( n26231 , n21070 , n27078 );
    and g1545 ( n23562 , n3198 , n18766 );
    or g1546 ( n16225 , n21896 , n12494 );
    xnor g1547 ( n20579 , n15636 , n11615 );
    and g1548 ( n21183 , n19242 , n3215 );
    nor g1549 ( n14632 , n4181 , n2194 );
    and g1550 ( n3413 , n14336 , n18149 );
    and g1551 ( n14240 , n15819 , n3763 );
    or g1552 ( n22423 , n9692 , n6761 );
    nor g1553 ( n11392 , n3843 , n1336 );
    and g1554 ( n12715 , n14818 , n26491 );
    or g1555 ( n23557 , n3828 , n10392 );
    not g1556 ( n6222 , n11273 );
    nor g1557 ( n11968 , n23996 , n5685 );
    xnor g1558 ( n12099 , n19110 , n5467 );
    or g1559 ( n24869 , n867 , n21430 );
    and g1560 ( n4474 , n20180 , n26616 );
    or g1561 ( n1382 , n25070 , n20637 );
    and g1562 ( n7140 , n24223 , n14259 );
    or g1563 ( n10825 , n23901 , n16038 );
    or g1564 ( n6347 , n25846 , n5874 );
    or g1565 ( n18030 , n2235 , n3556 );
    not g1566 ( n25271 , n19357 );
    nor g1567 ( n27191 , n8402 , n10987 );
    or g1568 ( n14623 , n27131 , n473 );
    xnor g1569 ( n9151 , n20175 , n4514 );
    and g1570 ( n2800 , n10530 , n21500 );
    xnor g1571 ( n21818 , n14016 , n22282 );
    or g1572 ( n12240 , n20777 , n4712 );
    xnor g1573 ( n16519 , n18196 , n25380 );
    xnor g1574 ( n2454 , n12229 , n442 );
    not g1575 ( n151 , n11971 );
    not g1576 ( n15905 , n7678 );
    nor g1577 ( n15503 , n3959 , n5855 );
    not g1578 ( n17433 , n9997 );
    and g1579 ( n10215 , n20097 , n11934 );
    or g1580 ( n7153 , n20864 , n25262 );
    xnor g1581 ( n1883 , n21577 , n20290 );
    not g1582 ( n13305 , n1160 );
    nor g1583 ( n9027 , n2453 , n23095 );
    nor g1584 ( n5619 , n24018 , n10499 );
    xnor g1585 ( n5608 , n9493 , n4426 );
    and g1586 ( n16437 , n27061 , n8617 );
    and g1587 ( n284 , n11590 , n21690 );
    nor g1588 ( n5690 , n20259 , n22043 );
    or g1589 ( n22001 , n24014 , n12728 );
    not g1590 ( n19862 , n6385 );
    xnor g1591 ( n10685 , n13945 , n19163 );
    xnor g1592 ( n11494 , n25688 , n27104 );
    xnor g1593 ( n154 , n2982 , n21120 );
    or g1594 ( n25544 , n987 , n11871 );
    and g1595 ( n13192 , n20522 , n17007 );
    nor g1596 ( n22418 , n24879 , n3687 );
    xnor g1597 ( n20060 , n17886 , n20219 );
    xnor g1598 ( n10468 , n20374 , n1266 );
    or g1599 ( n14802 , n7119 , n25171 );
    or g1600 ( n25035 , n15276 , n21659 );
    xnor g1601 ( n26699 , n10995 , n13894 );
    xnor g1602 ( n2948 , n19343 , n7958 );
    or g1603 ( n7411 , n16417 , n2924 );
    and g1604 ( n12571 , n13514 , n5492 );
    not g1605 ( n19956 , n16833 );
    xnor g1606 ( n22458 , n20754 , n24786 );
    not g1607 ( n23321 , n22909 );
    nor g1608 ( n3422 , n20036 , n23537 );
    or g1609 ( n16741 , n14909 , n2601 );
    or g1610 ( n4708 , n18554 , n4497 );
    or g1611 ( n14604 , n20489 , n26913 );
    nor g1612 ( n7733 , n25015 , n1850 );
    or g1613 ( n21709 , n3160 , n9414 );
    nor g1614 ( n12831 , n446 , n12650 );
    not g1615 ( n642 , n17780 );
    and g1616 ( n21616 , n4584 , n11916 );
    xnor g1617 ( n25102 , n24561 , n8782 );
    xnor g1618 ( n18277 , n2601 , n10304 );
    nor g1619 ( n22523 , n23114 , n3454 );
    or g1620 ( n12331 , n15620 , n7977 );
    not g1621 ( n21608 , n376 );
    xnor g1622 ( n15004 , n23201 , n23151 );
    and g1623 ( n7903 , n10648 , n18392 );
    or g1624 ( n8876 , n12169 , n6414 );
    not g1625 ( n19543 , n9376 );
    or g1626 ( n21279 , n15217 , n17542 );
    and g1627 ( n16955 , n22424 , n25417 );
    nor g1628 ( n12524 , n16543 , n22862 );
    and g1629 ( n25022 , n23913 , n8144 );
    xnor g1630 ( n26044 , n6848 , n23920 );
    not g1631 ( n14016 , n25436 );
    nor g1632 ( n2296 , n16536 , n13492 );
    or g1633 ( n23765 , n592 , n3347 );
    and g1634 ( n15245 , n21138 , n23804 );
    nor g1635 ( n10738 , n25021 , n21997 );
    xnor g1636 ( n8965 , n14635 , n15773 );
    or g1637 ( n11984 , n27001 , n12263 );
    not g1638 ( n5108 , n1658 );
    xnor g1639 ( n19646 , n13077 , n7702 );
    not g1640 ( n25953 , n25490 );
    and g1641 ( n23730 , n17240 , n4355 );
    or g1642 ( n11887 , n6995 , n8452 );
    or g1643 ( n5966 , n1819 , n19709 );
    or g1644 ( n19458 , n7501 , n14717 );
    or g1645 ( n668 , n19887 , n22246 );
    or g1646 ( n15098 , n7382 , n20018 );
    or g1647 ( n5686 , n26830 , n19707 );
    nor g1648 ( n16326 , n18123 , n4569 );
    and g1649 ( n21445 , n18185 , n19801 );
    or g1650 ( n15348 , n22480 , n17703 );
    xnor g1651 ( n17353 , n26124 , n6379 );
    nor g1652 ( n3737 , n4859 , n25972 );
    or g1653 ( n25311 , n8735 , n2055 );
    or g1654 ( n21019 , n11337 , n12430 );
    nor g1655 ( n24571 , n27113 , n16704 );
    xor g1656 ( n5164 , n25249 , n25795 );
    and g1657 ( n17952 , n9690 , n24036 );
    or g1658 ( n21145 , n18382 , n24216 );
    or g1659 ( n5017 , n18101 , n12550 );
    xnor g1660 ( n13005 , n2074 , n2390 );
    or g1661 ( n26430 , n26266 , n22785 );
    or g1662 ( n13063 , n9138 , n10896 );
    not g1663 ( n173 , n24129 );
    or g1664 ( n6384 , n20617 , n26977 );
    or g1665 ( n3212 , n3142 , n12937 );
    nor g1666 ( n3561 , n16776 , n25386 );
    or g1667 ( n164 , n3473 , n20580 );
    or g1668 ( n15953 , n26592 , n21932 );
    or g1669 ( n9181 , n5295 , n9812 );
    not g1670 ( n12693 , n14110 );
    and g1671 ( n17602 , n26636 , n19661 );
    not g1672 ( n24936 , n18833 );
    xnor g1673 ( n5770 , n17350 , n8784 );
    not g1674 ( n2049 , n16896 );
    or g1675 ( n20856 , n18916 , n1974 );
    nor g1676 ( n24181 , n22191 , n265 );
    and g1677 ( n364 , n1118 , n6477 );
    xnor g1678 ( n25043 , n8708 , n21047 );
    xnor g1679 ( n450 , n14337 , n7876 );
    and g1680 ( n8504 , n6659 , n12991 );
    not g1681 ( n20558 , n13743 );
    xnor g1682 ( n14008 , n928 , n21384 );
    nor g1683 ( n18669 , n16029 , n19228 );
    nor g1684 ( n15622 , n12405 , n19489 );
    or g1685 ( n2795 , n2371 , n19255 );
    or g1686 ( n8499 , n19867 , n27191 );
    or g1687 ( n22205 , n15066 , n6970 );
    not g1688 ( n16200 , n16312 );
    or g1689 ( n981 , n7049 , n18877 );
    or g1690 ( n21277 , n13944 , n23871 );
    not g1691 ( n17428 , n18281 );
    nor g1692 ( n15942 , n15167 , n23921 );
    and g1693 ( n13552 , n18138 , n14743 );
    and g1694 ( n22784 , n7129 , n8211 );
    xnor g1695 ( n21044 , n12658 , n26618 );
    or g1696 ( n20762 , n24867 , n5310 );
    xnor g1697 ( n10233 , n26748 , n12161 );
    and g1698 ( n1544 , n12866 , n24713 );
    nor g1699 ( n12976 , n11669 , n11366 );
    not g1700 ( n10683 , n3161 );
    xnor g1701 ( n24629 , n11240 , n24271 );
    and g1702 ( n18918 , n16580 , n19587 );
    xnor g1703 ( n21005 , n13282 , n14685 );
    not g1704 ( n24890 , n18558 );
    or g1705 ( n3605 , n15167 , n25330 );
    nor g1706 ( n22220 , n17979 , n11158 );
    nor g1707 ( n6959 , n27100 , n25637 );
    nor g1708 ( n17794 , n7817 , n23036 );
    xnor g1709 ( n6129 , n16474 , n15491 );
    and g1710 ( n17054 , n20040 , n23983 );
    or g1711 ( n2907 , n25409 , n23154 );
    not g1712 ( n19844 , n4296 );
    xnor g1713 ( n15220 , n18049 , n2365 );
    and g1714 ( n9236 , n26263 , n77 );
    or g1715 ( n5534 , n14163 , n921 );
    not g1716 ( n19914 , n4446 );
    nor g1717 ( n3452 , n23168 , n13028 );
    xnor g1718 ( n17075 , n2687 , n6346 );
    nor g1719 ( n20486 , n2141 , n23851 );
    xnor g1720 ( n12776 , n106 , n26882 );
    or g1721 ( n26175 , n15665 , n1033 );
    nor g1722 ( n19827 , n3124 , n5516 );
    xnor g1723 ( n7894 , n10303 , n1136 );
    xnor g1724 ( n24700 , n21415 , n924 );
    or g1725 ( n12899 , n22918 , n20719 );
    and g1726 ( n4504 , n13781 , n24358 );
    nor g1727 ( n13887 , n10051 , n3526 );
    not g1728 ( n19181 , n26936 );
    xnor g1729 ( n5419 , n10981 , n6517 );
    not g1730 ( n8623 , n23181 );
    and g1731 ( n3323 , n18442 , n12611 );
    nor g1732 ( n1804 , n25021 , n19025 );
    and g1733 ( n19339 , n11159 , n10186 );
    and g1734 ( n20815 , n26779 , n5588 );
    or g1735 ( n14219 , n1825 , n15095 );
    not g1736 ( n26680 , n3846 );
    xnor g1737 ( n13826 , n18707 , n19618 );
    xnor g1738 ( n21525 , n25780 , n26969 );
    or g1739 ( n7655 , n17300 , n12466 );
    xnor g1740 ( n4813 , n1398 , n1552 );
    or g1741 ( n16112 , n18857 , n5242 );
    and g1742 ( n4080 , n18080 , n24398 );
    and g1743 ( n23907 , n13385 , n8618 );
    or g1744 ( n20870 , n26571 , n21791 );
    nor g1745 ( n19088 , n11425 , n12657 );
    and g1746 ( n39 , n9193 , n12854 );
    not g1747 ( n1151 , n6218 );
    xnor g1748 ( n9463 , n11062 , n21489 );
    nor g1749 ( n15186 , n18814 , n8645 );
    and g1750 ( n25075 , n8685 , n21283 );
    xnor g1751 ( n16617 , n18359 , n1052 );
    xnor g1752 ( n16077 , n5570 , n17667 );
    and g1753 ( n13896 , n17523 , n5671 );
    or g1754 ( n19559 , n5885 , n17686 );
    or g1755 ( n8450 , n9011 , n19143 );
    xnor g1756 ( n4424 , n18706 , n11744 );
    or g1757 ( n18884 , n9679 , n4319 );
    or g1758 ( n19073 , n744 , n18630 );
    not g1759 ( n23921 , n3786 );
    xnor g1760 ( n14176 , n16743 , n5882 );
    or g1761 ( n25481 , n25291 , n13743 );
    and g1762 ( n7179 , n22039 , n1520 );
    xnor g1763 ( n23498 , n5165 , n6834 );
    or g1764 ( n14660 , n23990 , n14184 );
    or g1765 ( n24249 , n8827 , n26142 );
    xnor g1766 ( n26343 , n11390 , n26705 );
    or g1767 ( n26253 , n18145 , n12168 );
    or g1768 ( n25105 , n20411 , n17212 );
    xnor g1769 ( n20609 , n378 , n23743 );
    or g1770 ( n11490 , n5624 , n21632 );
    not g1771 ( n14557 , n17152 );
    xnor g1772 ( n6467 , n26584 , n14830 );
    nor g1773 ( n9805 , n12446 , n6553 );
    and g1774 ( n6582 , n15070 , n25672 );
    not g1775 ( n10885 , n24292 );
    xnor g1776 ( n11539 , n21121 , n22692 );
    or g1777 ( n25287 , n27183 , n2150 );
    and g1778 ( n8301 , n25218 , n5527 );
    or g1779 ( n8350 , n5491 , n4664 );
    or g1780 ( n17260 , n3791 , n24301 );
    nor g1781 ( n12444 , n22425 , n4461 );
    xnor g1782 ( n21736 , n14758 , n25636 );
    xnor g1783 ( n16068 , n22648 , n8530 );
    not g1784 ( n20358 , n23104 );
    and g1785 ( n13742 , n24639 , n7663 );
    xnor g1786 ( n13142 , n2289 , n20946 );
    xnor g1787 ( n5617 , n9236 , n17157 );
    or g1788 ( n20903 , n20532 , n7416 );
    or g1789 ( n21650 , n24402 , n13123 );
    and g1790 ( n25646 , n15882 , n25039 );
    xnor g1791 ( n2723 , n1846 , n22502 );
    not g1792 ( n25237 , n5669 );
    and g1793 ( n22528 , n16020 , n10907 );
    and g1794 ( n5431 , n16476 , n19146 );
    or g1795 ( n662 , n10721 , n7845 );
    or g1796 ( n1748 , n22186 , n11657 );
    nor g1797 ( n23314 , n23864 , n17994 );
    nor g1798 ( n3408 , n1262 , n1777 );
    xnor g1799 ( n3343 , n18298 , n14952 );
    and g1800 ( n334 , n6984 , n3954 );
    and g1801 ( n6927 , n8244 , n22820 );
    and g1802 ( n11084 , n19764 , n8114 );
    xnor g1803 ( n20364 , n4299 , n10843 );
    or g1804 ( n25028 , n12217 , n5701 );
    xnor g1805 ( n21120 , n4870 , n2857 );
    xnor g1806 ( n26073 , n3783 , n11630 );
    not g1807 ( n8851 , n20794 );
    xnor g1808 ( n6407 , n2554 , n14949 );
    not g1809 ( n15695 , n22843 );
    not g1810 ( n7143 , n400 );
    and g1811 ( n3214 , n13859 , n26276 );
    xnor g1812 ( n7660 , n12217 , n23798 );
    xnor g1813 ( n13877 , n8107 , n18363 );
    xnor g1814 ( n23279 , n26983 , n24076 );
    not g1815 ( n8735 , n23559 );
    or g1816 ( n18184 , n9705 , n12448 );
    or g1817 ( n6588 , n16464 , n16223 );
    not g1818 ( n13172 , n8827 );
    xnor g1819 ( n26287 , n18757 , n5162 );
    and g1820 ( n715 , n23494 , n14812 );
    not g1821 ( n26993 , n18805 );
    and g1822 ( n4837 , n6442 , n8959 );
    or g1823 ( n9951 , n8101 , n3019 );
    and g1824 ( n26684 , n12624 , n15735 );
    xnor g1825 ( n7162 , n14815 , n18958 );
    or g1826 ( n17825 , n24264 , n7178 );
    not g1827 ( n11835 , n10651 );
    or g1828 ( n18292 , n18765 , n21975 );
    or g1829 ( n8325 , n25502 , n1545 );
    not g1830 ( n2756 , n20477 );
    or g1831 ( n779 , n8345 , n24628 );
    not g1832 ( n739 , n25814 );
    and g1833 ( n11349 , n27183 , n2150 );
    or g1834 ( n17435 , n25748 , n3751 );
    or g1835 ( n7404 , n15676 , n21116 );
    or g1836 ( n11939 , n1656 , n11397 );
    or g1837 ( n22709 , n12709 , n8085 );
    and g1838 ( n20147 , n4352 , n11683 );
    xnor g1839 ( n23650 , n20134 , n15237 );
    or g1840 ( n5702 , n24229 , n5801 );
    and g1841 ( n20598 , n7644 , n11235 );
    or g1842 ( n18019 , n19848 , n6979 );
    and g1843 ( n3644 , n14431 , n25739 );
    nor g1844 ( n25407 , n3840 , n11254 );
    or g1845 ( n18401 , n14655 , n9565 );
    and g1846 ( n16330 , n15061 , n14892 );
    not g1847 ( n8415 , n19707 );
    and g1848 ( n24356 , n9417 , n11558 );
    or g1849 ( n17364 , n2520 , n2267 );
    xnor g1850 ( n6838 , n22119 , n9252 );
    xnor g1851 ( n3421 , n1163 , n24620 );
    not g1852 ( n23084 , n6246 );
    xnor g1853 ( n5637 , n19005 , n24618 );
    or g1854 ( n6252 , n524 , n14736 );
    or g1855 ( n10697 , n13590 , n22370 );
    nor g1856 ( n15224 , n19616 , n26673 );
    and g1857 ( n7291 , n5015 , n18246 );
    xnor g1858 ( n23032 , n19156 , n24706 );
    or g1859 ( n7611 , n6111 , n16868 );
    and g1860 ( n22904 , n11331 , n17988 );
    xnor g1861 ( n3728 , n19594 , n25627 );
    nor g1862 ( n13290 , n10184 , n22470 );
    xnor g1863 ( n10766 , n20151 , n19042 );
    xnor g1864 ( n15919 , n8974 , n14289 );
    or g1865 ( n18772 , n16819 , n5017 );
    or g1866 ( n7699 , n9732 , n26441 );
    and g1867 ( n5738 , n569 , n8110 );
    or g1868 ( n1135 , n27068 , n10505 );
    xnor g1869 ( n8215 , n7220 , n17920 );
    not g1870 ( n5212 , n12168 );
    xnor g1871 ( n9487 , n4602 , n12402 );
    nor g1872 ( n24103 , n16544 , n2160 );
    xnor g1873 ( n1239 , n22397 , n12191 );
    or g1874 ( n21027 , n18384 , n12952 );
    xnor g1875 ( n13650 , n1688 , n3544 );
    and g1876 ( n23859 , n27125 , n26595 );
    xnor g1877 ( n14941 , n4973 , n17563 );
    xnor g1878 ( n14300 , n21140 , n24456 );
    not g1879 ( n17812 , n12145 );
    not g1880 ( n20808 , n22748 );
    not g1881 ( n5341 , n14066 );
    xnor g1882 ( n17813 , n26724 , n1777 );
    xnor g1883 ( n24977 , n26875 , n6131 );
    xnor g1884 ( n10196 , n6442 , n6828 );
    xnor g1885 ( n11738 , n8828 , n6443 );
    xnor g1886 ( n3832 , n6797 , n22568 );
    xnor g1887 ( n8762 , n6895 , n4858 );
    nor g1888 ( n13126 , n23317 , n38 );
    nor g1889 ( n20789 , n26982 , n2679 );
    xnor g1890 ( n12125 , n5657 , n5704 );
    nor g1891 ( n12427 , n5914 , n790 );
    or g1892 ( n26357 , n26059 , n7672 );
    and g1893 ( n2354 , n18274 , n24383 );
    nor g1894 ( n22 , n3743 , n3038 );
    nor g1895 ( n4473 , n19680 , n18341 );
    and g1896 ( n10232 , n8064 , n449 );
    xnor g1897 ( n13841 , n8030 , n4050 );
    xnor g1898 ( n18888 , n22690 , n4736 );
    and g1899 ( n19580 , n26547 , n15163 );
    not g1900 ( n22968 , n17277 );
    nor g1901 ( n25548 , n9069 , n22169 );
    xnor g1902 ( n5024 , n23764 , n21533 );
    or g1903 ( n8029 , n122 , n15227 );
    nor g1904 ( n2616 , n23146 , n21585 );
    or g1905 ( n16370 , n14186 , n27170 );
    xnor g1906 ( n24133 , n12370 , n11613 );
    nor g1907 ( n10090 , n25370 , n23819 );
    xnor g1908 ( n13230 , n4502 , n13760 );
    not g1909 ( n401 , n19905 );
    xor g1910 ( n25647 , n11707 , n14829 );
    and g1911 ( n17702 , n2735 , n5628 );
    not g1912 ( n13553 , n18632 );
    or g1913 ( n8469 , n9361 , n2947 );
    xnor g1914 ( n2470 , n21333 , n232 );
    not g1915 ( n13982 , n13006 );
    or g1916 ( n17233 , n9257 , n5798 );
    and g1917 ( n17802 , n26797 , n14654 );
    or g1918 ( n8142 , n27038 , n19374 );
    xnor g1919 ( n9726 , n10196 , n20741 );
    xnor g1920 ( n14687 , n1802 , n6038 );
    or g1921 ( n116 , n20023 , n12734 );
    or g1922 ( n1776 , n17954 , n23767 );
    or g1923 ( n13233 , n21188 , n10011 );
    or g1924 ( n14173 , n19277 , n6327 );
    xnor g1925 ( n8349 , n18664 , n9077 );
    nor g1926 ( n22155 , n20966 , n17938 );
    or g1927 ( n8357 , n8212 , n1782 );
    or g1928 ( n24332 , n3594 , n1504 );
    xnor g1929 ( n115 , n16723 , n24618 );
    xnor g1930 ( n4284 , n1380 , n11220 );
    nor g1931 ( n2975 , n2750 , n7543 );
    and g1932 ( n15119 , n6348 , n6116 );
    not g1933 ( n24813 , n11817 );
    not g1934 ( n18787 , n7775 );
    xnor g1935 ( n7406 , n16821 , n21545 );
    xnor g1936 ( n14996 , n22956 , n11952 );
    not g1937 ( n3632 , n26311 );
    nor g1938 ( n20768 , n1690 , n1000 );
    or g1939 ( n14485 , n12940 , n6157 );
    xnor g1940 ( n10409 , n11214 , n2078 );
    xnor g1941 ( n8296 , n22892 , n24298 );
    xnor g1942 ( n1733 , n24091 , n2272 );
    and g1943 ( n9383 , n18151 , n6414 );
    or g1944 ( n5327 , n10494 , n26304 );
    xnor g1945 ( n11287 , n14826 , n17458 );
    or g1946 ( n23327 , n17780 , n12430 );
    and g1947 ( n20202 , n22626 , n18765 );
    xnor g1948 ( n18302 , n8571 , n10872 );
    or g1949 ( n20969 , n25680 , n14348 );
    xnor g1950 ( n19378 , n10837 , n1576 );
    not g1951 ( n13062 , n23432 );
    or g1952 ( n13537 , n20777 , n2461 );
    not g1953 ( n14255 , n17064 );
    nor g1954 ( n9991 , n19588 , n13329 );
    nor g1955 ( n10147 , n4479 , n23724 );
    and g1956 ( n14001 , n19361 , n15918 );
    nor g1957 ( n6930 , n16932 , n6913 );
    or g1958 ( n21947 , n17999 , n17982 );
    or g1959 ( n25154 , n25506 , n14237 );
    xnor g1960 ( n15190 , n25880 , n18609 );
    and g1961 ( n542 , n1144 , n9299 );
    and g1962 ( n22876 , n15550 , n2347 );
    xnor g1963 ( n185 , n24862 , n3906 );
    or g1964 ( n4352 , n4085 , n16547 );
    or g1965 ( n15966 , n8845 , n22773 );
    or g1966 ( n237 , n24004 , n12900 );
    and g1967 ( n2386 , n160 , n25275 );
    xnor g1968 ( n16759 , n17881 , n25068 );
    or g1969 ( n5761 , n2409 , n25057 );
    or g1970 ( n11610 , n18737 , n2328 );
    and g1971 ( n3944 , n12997 , n13532 );
    or g1972 ( n1219 , n16319 , n19170 );
    and g1973 ( n23527 , n94 , n9476 );
    not g1974 ( n339 , n9926 );
    and g1975 ( n26977 , n2527 , n23507 );
    xnor g1976 ( n16746 , n10650 , n22253 );
    or g1977 ( n5900 , n9883 , n13885 );
    xnor g1978 ( n3794 , n18390 , n13587 );
    nor g1979 ( n3750 , n16880 , n21734 );
    xnor g1980 ( n6418 , n12911 , n1222 );
    and g1981 ( n8034 , n3466 , n19917 );
    xnor g1982 ( n7052 , n2085 , n5169 );
    not g1983 ( n20089 , n12384 );
    or g1984 ( n23815 , n10043 , n25252 );
    not g1985 ( n5569 , n26216 );
    or g1986 ( n12052 , n25445 , n244 );
    and g1987 ( n26889 , n21588 , n15449 );
    xnor g1988 ( n8722 , n6931 , n17612 );
    not g1989 ( n9290 , n9460 );
    and g1990 ( n11341 , n12923 , n204 );
    xnor g1991 ( n2695 , n2155 , n16938 );
    and g1992 ( n12577 , n689 , n19627 );
    not g1993 ( n17610 , n26752 );
    or g1994 ( n10690 , n25841 , n3053 );
    xnor g1995 ( n8672 , n26886 , n1099 );
    not g1996 ( n19229 , n2146 );
    or g1997 ( n19293 , n19797 , n3903 );
    not g1998 ( n2071 , n14480 );
    or g1999 ( n2182 , n10696 , n72 );
    or g2000 ( n25162 , n11804 , n17755 );
    or g2001 ( n14807 , n17248 , n21020 );
    xnor g2002 ( n16319 , n25030 , n1549 );
    or g2003 ( n25534 , n26036 , n7832 );
    xnor g2004 ( n10210 , n2432 , n15017 );
    not g2005 ( n23175 , n8850 );
    nor g2006 ( n24050 , n22550 , n7465 );
    xnor g2007 ( n4410 , n25081 , n17560 );
    and g2008 ( n18432 , n3493 , n24087 );
    or g2009 ( n2603 , n10313 , n26932 );
    nor g2010 ( n17234 , n3405 , n9665 );
    not g2011 ( n3939 , n17204 );
    or g2012 ( n14141 , n3915 , n17411 );
    or g2013 ( n18369 , n1879 , n670 );
    not g2014 ( n14700 , n6734 );
    and g2015 ( n5197 , n5061 , n6016 );
    or g2016 ( n23496 , n5567 , n19152 );
    xnor g2017 ( n23754 , n12310 , n6575 );
    or g2018 ( n13882 , n6805 , n8679 );
    or g2019 ( n8829 , n19890 , n12810 );
    xnor g2020 ( n18970 , n26663 , n20087 );
    not g2021 ( n15 , n21143 );
    xnor g2022 ( n20287 , n11802 , n9112 );
    xnor g2023 ( n23100 , n9765 , n20213 );
    nor g2024 ( n21756 , n6032 , n13623 );
    xnor g2025 ( n11408 , n27016 , n14947 );
    xnor g2026 ( n11787 , n8363 , n2816 );
    not g2027 ( n22071 , n1752 );
    or g2028 ( n4157 , n18207 , n25511 );
    and g2029 ( n18573 , n15636 , n25139 );
    or g2030 ( n9522 , n25628 , n27129 );
    or g2031 ( n9348 , n2176 , n19561 );
    nor g2032 ( n8203 , n25470 , n12898 );
    xnor g2033 ( n21919 , n19222 , n6691 );
    not g2034 ( n9404 , n25441 );
    and g2035 ( n20435 , n23011 , n23971 );
    xnor g2036 ( n23145 , n27109 , n3884 );
    nor g2037 ( n10397 , n24247 , n558 );
    or g2038 ( n19918 , n20497 , n16482 );
    not g2039 ( n1091 , n14323 );
    or g2040 ( n8104 , n18734 , n14870 );
    xnor g2041 ( n6445 , n15457 , n15997 );
    not g2042 ( n21910 , n1278 );
    not g2043 ( n19047 , n14648 );
    nor g2044 ( n11187 , n20151 , n22428 );
    and g2045 ( n26171 , n995 , n229 );
    xnor g2046 ( n17081 , n12950 , n8083 );
    nor g2047 ( n12841 , n801 , n10760 );
    or g2048 ( n12817 , n22725 , n11480 );
    and g2049 ( n12336 , n13777 , n15370 );
    or g2050 ( n26831 , n23430 , n20628 );
    xnor g2051 ( n2546 , n19702 , n19270 );
    xnor g2052 ( n3960 , n4236 , n22846 );
    or g2053 ( n2791 , n5993 , n13104 );
    or g2054 ( n13931 , n10209 , n19442 );
    and g2055 ( n4805 , n20831 , n26690 );
    not g2056 ( n26300 , n21210 );
    or g2057 ( n2685 , n22820 , n19137 );
    nor g2058 ( n13515 , n11302 , n20948 );
    nor g2059 ( n14000 , n26255 , n27102 );
    xnor g2060 ( n14843 , n15603 , n15901 );
    or g2061 ( n21372 , n26895 , n13543 );
    not g2062 ( n2085 , n4759 );
    xnor g2063 ( n12725 , n3654 , n20996 );
    and g2064 ( n23499 , n4390 , n2381 );
    not g2065 ( n17360 , n23890 );
    and g2066 ( n8963 , n5397 , n17825 );
    or g2067 ( n14489 , n4144 , n25634 );
    nor g2068 ( n26377 , n10903 , n24584 );
    or g2069 ( n20766 , n3428 , n25216 );
    xnor g2070 ( n1891 , n19008 , n2524 );
    nor g2071 ( n3114 , n12265 , n5728 );
    xnor g2072 ( n6470 , n13055 , n20172 );
    nor g2073 ( n21829 , n5374 , n23002 );
    or g2074 ( n14159 , n3736 , n4790 );
    xnor g2075 ( n10797 , n12717 , n25679 );
    xnor g2076 ( n22355 , n7628 , n23982 );
    xnor g2077 ( n21746 , n4749 , n12385 );
    xnor g2078 ( n19642 , n10590 , n3677 );
    and g2079 ( n1812 , n12107 , n10853 );
    not g2080 ( n5172 , n6379 );
    and g2081 ( n3226 , n15861 , n4887 );
    xnor g2082 ( n15406 , n20937 , n21596 );
    xnor g2083 ( n25418 , n13748 , n24923 );
    and g2084 ( n8517 , n9614 , n6890 );
    xnor g2085 ( n24035 , n26495 , n5789 );
    not g2086 ( n26769 , n26935 );
    nor g2087 ( n4159 , n2713 , n25271 );
    xnor g2088 ( n18693 , n2584 , n10698 );
    xnor g2089 ( n20594 , n10198 , n6119 );
    or g2090 ( n18214 , n20112 , n26102 );
    nor g2091 ( n1785 , n8196 , n3992 );
    xnor g2092 ( n6772 , n15389 , n23913 );
    or g2093 ( n13902 , n8647 , n26226 );
    nor g2094 ( n23957 , n14761 , n26460 );
    and g2095 ( n3065 , n1556 , n13974 );
    xnor g2096 ( n5062 , n4934 , n18279 );
    and g2097 ( n22935 , n19586 , n18147 );
    and g2098 ( n6277 , n13666 , n1131 );
    nor g2099 ( n16155 , n13668 , n835 );
    or g2100 ( n7565 , n21979 , n23135 );
    or g2101 ( n25909 , n24311 , n17430 );
    xnor g2102 ( n17853 , n22378 , n22619 );
    and g2103 ( n138 , n26648 , n8817 );
    and g2104 ( n3607 , n7066 , n9413 );
    and g2105 ( n4699 , n3506 , n26414 );
    or g2106 ( n14921 , n7396 , n27178 );
    nor g2107 ( n10209 , n12650 , n11220 );
    xnor g2108 ( n8660 , n20638 , n10512 );
    xnor g2109 ( n8320 , n16100 , n23139 );
    xnor g2110 ( n11313 , n4663 , n8409 );
    and g2111 ( n18063 , n8129 , n8972 );
    or g2112 ( n25335 , n647 , n1773 );
    or g2113 ( n18842 , n6209 , n2597 );
    not g2114 ( n8227 , n2111 );
    and g2115 ( n15509 , n15920 , n13545 );
    xnor g2116 ( n19982 , n19411 , n5978 );
    or g2117 ( n15480 , n10319 , n23812 );
    xnor g2118 ( n7086 , n26008 , n17201 );
    or g2119 ( n24205 , n2102 , n19560 );
    nor g2120 ( n5907 , n19406 , n21905 );
    and g2121 ( n20152 , n26870 , n7902 );
    xnor g2122 ( n2586 , n26011 , n4154 );
    xnor g2123 ( n25106 , n20999 , n3353 );
    nor g2124 ( n18221 , n20137 , n17077 );
    nor g2125 ( n13991 , n11525 , n11258 );
    and g2126 ( n23485 , n17896 , n1475 );
    and g2127 ( n18144 , n20375 , n16075 );
    xnor g2128 ( n25104 , n18047 , n22933 );
    or g2129 ( n6479 , n16910 , n502 );
    or g2130 ( n23906 , n10190 , n5478 );
    xnor g2131 ( n23667 , n7604 , n11580 );
    or g2132 ( n23112 , n5406 , n11145 );
    xnor g2133 ( n25852 , n20011 , n17953 );
    xnor g2134 ( n7271 , n23352 , n22953 );
    not g2135 ( n14249 , n10765 );
    or g2136 ( n14426 , n2979 , n23258 );
    or g2137 ( n3434 , n22867 , n12334 );
    nor g2138 ( n15369 , n26654 , n3554 );
    xnor g2139 ( n4451 , n1675 , n20220 );
    and g2140 ( n25881 , n1571 , n23833 );
    nor g2141 ( n3423 , n19888 , n13308 );
    xnor g2142 ( n13648 , n10152 , n10581 );
    and g2143 ( n21274 , n13173 , n10006 );
    or g2144 ( n16749 , n11328 , n21255 );
    xnor g2145 ( n24579 , n19219 , n27197 );
    nor g2146 ( n9725 , n7674 , n16468 );
    nor g2147 ( n26123 , n2057 , n19603 );
    and g2148 ( n10524 , n23021 , n4690 );
    not g2149 ( n7953 , n13775 );
    not g2150 ( n15897 , n3012 );
    xnor g2151 ( n8487 , n1542 , n12916 );
    or g2152 ( n20281 , n13822 , n767 );
    or g2153 ( n11466 , n23114 , n6362 );
    or g2154 ( n5422 , n11188 , n21316 );
    and g2155 ( n17541 , n6185 , n11646 );
    and g2156 ( n20979 , n26284 , n12403 );
    not g2157 ( n12040 , n2732 );
    or g2158 ( n23614 , n4085 , n3211 );
    or g2159 ( n12431 , n10274 , n17636 );
    xnor g2160 ( n17978 , n24717 , n2979 );
    or g2161 ( n20884 , n26899 , n4743 );
    xnor g2162 ( n11095 , n24985 , n185 );
    or g2163 ( n15103 , n3984 , n22153 );
    nor g2164 ( n18012 , n2341 , n2967 );
    not g2165 ( n22261 , n3306 );
    or g2166 ( n3558 , n20224 , n23881 );
    not g2167 ( n5523 , n24474 );
    buf g2168 ( n8492 , n15931 );
    xnor g2169 ( n7779 , n13745 , n26460 );
    xnor g2170 ( n19363 , n10710 , n23529 );
    or g2171 ( n11626 , n25129 , n9446 );
    xnor g2172 ( n4762 , n14507 , n17488 );
    xnor g2173 ( n4890 , n10081 , n890 );
    xnor g2174 ( n5178 , n12633 , n9900 );
    or g2175 ( n19499 , n1203 , n24556 );
    and g2176 ( n22556 , n9045 , n4437 );
    xnor g2177 ( n24721 , n21644 , n18555 );
    or g2178 ( n12074 , n12458 , n26373 );
    and g2179 ( n547 , n9258 , n19250 );
    and g2180 ( n1345 , n1615 , n20856 );
    xnor g2181 ( n3663 , n24291 , n17196 );
    not g2182 ( n839 , n12342 );
    xnor g2183 ( n15758 , n10468 , n20770 );
    xnor g2184 ( n27177 , n12513 , n25568 );
    nor g2185 ( n19168 , n23313 , n16345 );
    not g2186 ( n1626 , n8391 );
    xnor g2187 ( n23453 , n7785 , n7817 );
    xnor g2188 ( n6394 , n24665 , n5704 );
    and g2189 ( n20895 , n26258 , n10154 );
    xnor g2190 ( n27055 , n1365 , n23333 );
    or g2191 ( n2435 , n8016 , n21911 );
    nor g2192 ( n5939 , n14230 , n10185 );
    or g2193 ( n22451 , n3599 , n5366 );
    or g2194 ( n20212 , n25726 , n5200 );
    xnor g2195 ( n5804 , n23084 , n3253 );
    or g2196 ( n13849 , n2970 , n3793 );
    xnor g2197 ( n9653 , n20295 , n23659 );
    xnor g2198 ( n22294 , n1686 , n1292 );
    not g2199 ( n17755 , n3031 );
    or g2200 ( n2763 , n21324 , n1446 );
    or g2201 ( n14020 , n10794 , n10400 );
    and g2202 ( n18855 , n1003 , n8931 );
    not g2203 ( n14033 , n1414 );
    not g2204 ( n20289 , n387 );
    or g2205 ( n1955 , n17768 , n8517 );
    and g2206 ( n16565 , n18749 , n4156 );
    or g2207 ( n20090 , n5572 , n7684 );
    or g2208 ( n18127 , n14560 , n4267 );
    xnor g2209 ( n19355 , n20828 , n6751 );
    xnor g2210 ( n7684 , n2398 , n107 );
    xnor g2211 ( n22933 , n8938 , n4255 );
    and g2212 ( n11051 , n405 , n4561 );
    xnor g2213 ( n16858 , n23878 , n2035 );
    xnor g2214 ( n9415 , n19863 , n2210 );
    not g2215 ( n16856 , n24488 );
    or g2216 ( n21992 , n25914 , n20359 );
    xnor g2217 ( n17902 , n15957 , n23697 );
    or g2218 ( n8543 , n821 , n17584 );
    xnor g2219 ( n18582 , n11215 , n19533 );
    not g2220 ( n26085 , n23235 );
    and g2221 ( n11983 , n21831 , n25448 );
    and g2222 ( n23102 , n13480 , n22769 );
    not g2223 ( n8719 , n8406 );
    xnor g2224 ( n17735 , n16132 , n22857 );
    and g2225 ( n26792 , n3629 , n10474 );
    or g2226 ( n18403 , n16903 , n17061 );
    or g2227 ( n25159 , n5068 , n14715 );
    xnor g2228 ( n15105 , n2980 , n12514 );
    and g2229 ( n26261 , n24321 , n18885 );
    xnor g2230 ( n24501 , n18229 , n25509 );
    xnor g2231 ( n21532 , n1437 , n17784 );
    and g2232 ( n20764 , n6608 , n19654 );
    and g2233 ( n23389 , n17603 , n22608 );
    xnor g2234 ( n25195 , n8713 , n24736 );
    nor g2235 ( n21715 , n3937 , n21295 );
    xnor g2236 ( n5769 , n2355 , n16223 );
    buf g2237 ( n11381 , n10777 );
    or g2238 ( n11686 , n24848 , n23972 );
    and g2239 ( n11327 , n2562 , n5823 );
    nor g2240 ( n11870 , n13136 , n26065 );
    not g2241 ( n24701 , n1162 );
    or g2242 ( n4653 , n17376 , n8842 );
    nor g2243 ( n15006 , n7769 , n26625 );
    xnor g2244 ( n11746 , n15512 , n22607 );
    or g2245 ( n7603 , n19068 , n9925 );
    and g2246 ( n15174 , n18027 , n4866 );
    and g2247 ( n19547 , n13982 , n15092 );
    xnor g2248 ( n17023 , n6381 , n13914 );
    and g2249 ( n26721 , n22896 , n26345 );
    xnor g2250 ( n12417 , n22449 , n7157 );
    not g2251 ( n17047 , n4537 );
    and g2252 ( n20960 , n16919 , n7628 );
    and g2253 ( n22541 , n19822 , n17760 );
    xnor g2254 ( n10466 , n10882 , n8406 );
    or g2255 ( n21916 , n3366 , n15670 );
    and g2256 ( n13120 , n9001 , n20995 );
    and g2257 ( n3535 , n2315 , n17375 );
    xnor g2258 ( n543 , n7888 , n5500 );
    xnor g2259 ( n18810 , n13884 , n7917 );
    xnor g2260 ( n20267 , n20796 , n5140 );
    or g2261 ( n22052 , n12811 , n11822 );
    nor g2262 ( n10067 , n19106 , n2680 );
    xnor g2263 ( n22635 , n22093 , n26743 );
    not g2264 ( n15796 , n13490 );
    not g2265 ( n18554 , n14230 );
    xnor g2266 ( n9750 , n15241 , n15146 );
    or g2267 ( n26502 , n7338 , n10899 );
    and g2268 ( n23780 , n3797 , n2203 );
    or g2269 ( n7922 , n26577 , n3052 );
    or g2270 ( n1167 , n16743 , n16875 );
    not g2271 ( n6137 , n3477 );
    not g2272 ( n26648 , n12440 );
    or g2273 ( n8049 , n20409 , n19117 );
    and g2274 ( n21514 , n16743 , n24485 );
    xnor g2275 ( n17382 , n25089 , n10253 );
    or g2276 ( n2624 , n13459 , n593 );
    not g2277 ( n22724 , n21222 );
    or g2278 ( n7078 , n8547 , n22045 );
    xnor g2279 ( n6463 , n16162 , n10251 );
    xnor g2280 ( n23086 , n18551 , n8632 );
    xnor g2281 ( n20772 , n20131 , n17418 );
    xnor g2282 ( n12329 , n13431 , n13943 );
    xnor g2283 ( n4182 , n26830 , n8415 );
    not g2284 ( n19615 , n26803 );
    not g2285 ( n4109 , n7706 );
    or g2286 ( n741 , n18485 , n2731 );
    or g2287 ( n8977 , n6204 , n5065 );
    xnor g2288 ( n25373 , n16482 , n13333 );
    xnor g2289 ( n22082 , n1271 , n26647 );
    nor g2290 ( n1103 , n8847 , n3993 );
    xnor g2291 ( n6003 , n9212 , n3456 );
    not g2292 ( n16618 , n24901 );
    xnor g2293 ( n4443 , n6259 , n24152 );
    or g2294 ( n2594 , n20326 , n5694 );
    or g2295 ( n22190 , n22882 , n21572 );
    nor g2296 ( n19195 , n10557 , n12381 );
    xnor g2297 ( n23864 , n23501 , n10563 );
    and g2298 ( n1257 , n1709 , n24961 );
    and g2299 ( n4550 , n22031 , n20824 );
    xnor g2300 ( n20574 , n20542 , n9575 );
    xnor g2301 ( n18002 , n26277 , n23778 );
    and g2302 ( n157 , n26510 , n11246 );
    xnor g2303 ( n14593 , n23017 , n23853 );
    xnor g2304 ( n22761 , n4244 , n7345 );
    not g2305 ( n9711 , n1845 );
    not g2306 ( n1329 , n5438 );
    xnor g2307 ( n16516 , n8838 , n4828 );
    and g2308 ( n11125 , n21867 , n8557 );
    and g2309 ( n38 , n13886 , n17242 );
    or g2310 ( n9029 , n22250 , n1071 );
    xnor g2311 ( n7640 , n3885 , n19208 );
    nor g2312 ( n16854 , n12398 , n23586 );
    and g2313 ( n2091 , n12622 , n26289 );
    or g2314 ( n13795 , n9053 , n22015 );
    nor g2315 ( n3879 , n23895 , n13976 );
    xnor g2316 ( n7950 , n19528 , n24782 );
    nor g2317 ( n23884 , n17004 , n24496 );
    nor g2318 ( n11316 , n23099 , n17517 );
    or g2319 ( n1964 , n6168 , n4537 );
    nor g2320 ( n23500 , n22849 , n16824 );
    and g2321 ( n19318 , n21528 , n7488 );
    xnor g2322 ( n23196 , n19905 , n3030 );
    not g2323 ( n7910 , n24203 );
    or g2324 ( n8684 , n20379 , n10677 );
    and g2325 ( n6452 , n932 , n2666 );
    and g2326 ( n21798 , n15103 , n25325 );
    and g2327 ( n8592 , n13052 , n4635 );
    xnor g2328 ( n14189 , n5441 , n2426 );
    xnor g2329 ( n2371 , n19213 , n25730 );
    xnor g2330 ( n13943 , n25049 , n23451 );
    or g2331 ( n23093 , n24582 , n14116 );
    xnor g2332 ( n18599 , n9272 , n16764 );
    or g2333 ( n2227 , n8451 , n7555 );
    or g2334 ( n8968 , n18514 , n15182 );
    not g2335 ( n5629 , n8297 );
    or g2336 ( n6258 , n26725 , n24292 );
    xnor g2337 ( n10908 , n26622 , n11471 );
    or g2338 ( n24952 , n18014 , n20619 );
    or g2339 ( n3702 , n23030 , n8381 );
    xnor g2340 ( n8282 , n4665 , n24278 );
    nor g2341 ( n6268 , n25913 , n15568 );
    or g2342 ( n16945 , n19339 , n21770 );
    xnor g2343 ( n19456 , n5739 , n4293 );
    xnor g2344 ( n6359 , n16313 , n25736 );
    not g2345 ( n6071 , n20417 );
    or g2346 ( n5861 , n787 , n9973 );
    xnor g2347 ( n3916 , n18145 , n19196 );
    nor g2348 ( n6027 , n14153 , n16466 );
    xnor g2349 ( n5936 , n10914 , n11892 );
    xnor g2350 ( n24993 , n14765 , n12650 );
    nor g2351 ( n21428 , n2651 , n4400 );
    nor g2352 ( n11826 , n481 , n11220 );
    xnor g2353 ( n12144 , n1444 , n15239 );
    xnor g2354 ( n11403 , n6297 , n17016 );
    nor g2355 ( n17676 , n17277 , n12869 );
    nor g2356 ( n3127 , n9445 , n5812 );
    or g2357 ( n13335 , n10277 , n1082 );
    or g2358 ( n19053 , n16806 , n16005 );
    or g2359 ( n19959 , n15244 , n23952 );
    and g2360 ( n11405 , n17581 , n4330 );
    and g2361 ( n22559 , n8101 , n9468 );
    not g2362 ( n15137 , n3071 );
    or g2363 ( n23332 , n19083 , n7450 );
    nor g2364 ( n8644 , n20059 , n15603 );
    nor g2365 ( n708 , n15580 , n4913 );
    xnor g2366 ( n3211 , n11549 , n14223 );
    or g2367 ( n18501 , n9863 , n19480 );
    and g2368 ( n17191 , n8069 , n4044 );
    and g2369 ( n18064 , n9607 , n14935 );
    xnor g2370 ( n20427 , n1197 , n25061 );
    xnor g2371 ( n5522 , n9206 , n23792 );
    xnor g2372 ( n5365 , n13359 , n4665 );
    or g2373 ( n2516 , n18814 , n802 );
    or g2374 ( n22235 , n726 , n26849 );
    and g2375 ( n24443 , n10382 , n24001 );
    not g2376 ( n19556 , n26248 );
    and g2377 ( n1770 , n23574 , n18923 );
    or g2378 ( n24515 , n23182 , n5542 );
    or g2379 ( n15646 , n11884 , n13313 );
    or g2380 ( n14925 , n23687 , n12025 );
    not g2381 ( n18786 , n2565 );
    not g2382 ( n5934 , n2900 );
    xnor g2383 ( n4368 , n14549 , n25861 );
    not g2384 ( n18581 , n11048 );
    not g2385 ( n21721 , n22395 );
    xnor g2386 ( n16264 , n6792 , n410 );
    nor g2387 ( n1281 , n7682 , n3952 );
    not g2388 ( n26124 , n3040 );
    not g2389 ( n11268 , n11383 );
    or g2390 ( n9545 , n23937 , n282 );
    xnor g2391 ( n12063 , n2570 , n7569 );
    or g2392 ( n17021 , n16594 , n23250 );
    or g2393 ( n27000 , n19372 , n25902 );
    xnor g2394 ( n985 , n13574 , n9341 );
    xnor g2395 ( n102 , n14079 , n19670 );
    xnor g2396 ( n15339 , n23827 , n27070 );
    not g2397 ( n2576 , n18157 );
    nor g2398 ( n1680 , n4877 , n11135 );
    not g2399 ( n4468 , n23974 );
    or g2400 ( n23992 , n8066 , n23340 );
    xnor g2401 ( n14393 , n20110 , n1147 );
    xnor g2402 ( n14391 , n9188 , n10612 );
    nor g2403 ( n1591 , n21740 , n12547 );
    and g2404 ( n21932 , n3941 , n2701 );
    or g2405 ( n27123 , n14882 , n21072 );
    or g2406 ( n5450 , n23390 , n1411 );
    not g2407 ( n6535 , n7073 );
    and g2408 ( n14994 , n9698 , n1818 );
    xnor g2409 ( n7256 , n13706 , n2033 );
    or g2410 ( n19092 , n19161 , n22405 );
    xnor g2411 ( n5832 , n13820 , n5541 );
    and g2412 ( n1287 , n2458 , n1732 );
    and g2413 ( n23373 , n11229 , n9741 );
    not g2414 ( n22219 , n3721 );
    or g2415 ( n3157 , n23920 , n25920 );
    or g2416 ( n6784 , n7521 , n9871 );
    or g2417 ( n17346 , n3349 , n10501 );
    and g2418 ( n9960 , n5538 , n24111 );
    not g2419 ( n19520 , n27170 );
    xnor g2420 ( n19968 , n16089 , n9316 );
    and g2421 ( n22690 , n4839 , n17133 );
    or g2422 ( n4131 , n14228 , n14770 );
    xnor g2423 ( n6383 , n22936 , n10596 );
    or g2424 ( n22827 , n8010 , n19086 );
    xnor g2425 ( n15969 , n7307 , n9728 );
    or g2426 ( n2609 , n24103 , n2025 );
    xnor g2427 ( n3229 , n2545 , n3740 );
    xnor g2428 ( n17436 , n872 , n10214 );
    not g2429 ( n2967 , n23068 );
    and g2430 ( n12388 , n25741 , n19942 );
    nor g2431 ( n2234 , n10098 , n263 );
    and g2432 ( n3798 , n3313 , n4367 );
    and g2433 ( n24381 , n22290 , n13018 );
    nor g2434 ( n18385 , n17351 , n21850 );
    and g2435 ( n6584 , n24417 , n4719 );
    not g2436 ( n13391 , n9850 );
    and g2437 ( n5560 , n19618 , n18707 );
    or g2438 ( n8560 , n18088 , n11173 );
    and g2439 ( n1578 , n1802 , n7331 );
    not g2440 ( n20129 , n25384 );
    or g2441 ( n24075 , n8199 , n22638 );
    nor g2442 ( n21036 , n18880 , n15456 );
    xnor g2443 ( n11025 , n5490 , n7599 );
    xnor g2444 ( n8744 , n4135 , n13610 );
    or g2445 ( n17053 , n25187 , n23728 );
    xnor g2446 ( n9093 , n23368 , n19793 );
    or g2447 ( n16023 , n19024 , n5893 );
    nor g2448 ( n4070 , n25603 , n14389 );
    xnor g2449 ( n2555 , n17332 , n9759 );
    xnor g2450 ( n16074 , n24170 , n24085 );
    or g2451 ( n26558 , n12196 , n18289 );
    or g2452 ( n2024 , n11915 , n21864 );
    xnor g2453 ( n4738 , n7827 , n9505 );
    xnor g2454 ( n4897 , n19010 , n10212 );
    and g2455 ( n11117 , n21171 , n10121 );
    xnor g2456 ( n25218 , n13505 , n10895 );
    xnor g2457 ( n7163 , n19608 , n15378 );
    xnor g2458 ( n20602 , n26351 , n26225 );
    and g2459 ( n13938 , n8820 , n13197 );
    xnor g2460 ( n12734 , n14918 , n16694 );
    or g2461 ( n14452 , n8266 , n7538 );
    xnor g2462 ( n27042 , n10852 , n9898 );
    xnor g2463 ( n608 , n20076 , n21082 );
    xnor g2464 ( n8090 , n20437 , n20151 );
    xnor g2465 ( n18609 , n21287 , n9967 );
    or g2466 ( n17327 , n23069 , n18153 );
    and g2467 ( n93 , n13006 , n20266 );
    or g2468 ( n21601 , n11392 , n6654 );
    or g2469 ( n4220 , n2576 , n13853 );
    not g2470 ( n6242 , n17132 );
    nor g2471 ( n2309 , n1895 , n20972 );
    not g2472 ( n12928 , n18486 );
    xnor g2473 ( n1027 , n16972 , n2895 );
    nor g2474 ( n17800 , n12655 , n11214 );
    xnor g2475 ( n20578 , n10522 , n23024 );
    nor g2476 ( n13757 , n1333 , n19051 );
    or g2477 ( n10769 , n5302 , n19116 );
    xnor g2478 ( n24908 , n6153 , n19775 );
    and g2479 ( n21722 , n14011 , n17309 );
    and g2480 ( n20828 , n10697 , n7075 );
    or g2481 ( n6016 , n15302 , n12912 );
    and g2482 ( n18718 , n18086 , n24777 );
    and g2483 ( n16298 , n5134 , n2830 );
    or g2484 ( n9640 , n10392 , n20897 );
    or g2485 ( n24976 , n20894 , n18022 );
    and g2486 ( n20295 , n1460 , n20783 );
    xnor g2487 ( n23429 , n23889 , n20616 );
    and g2488 ( n17937 , n6750 , n19058 );
    not g2489 ( n14514 , n16092 );
    xnor g2490 ( n1636 , n2820 , n13973 );
    not g2491 ( n18981 , n26334 );
    and g2492 ( n482 , n25976 , n4292 );
    xnor g2493 ( n11251 , n19033 , n17037 );
    not g2494 ( n9035 , n20192 );
    or g2495 ( n11558 , n4667 , n21654 );
    and g2496 ( n26329 , n2279 , n21232 );
    nor g2497 ( n11891 , n20604 , n23331 );
    not g2498 ( n26144 , n1822 );
    not g2499 ( n17607 , n22537 );
    and g2500 ( n12936 , n8703 , n25290 );
    not g2501 ( n2057 , n27185 );
    or g2502 ( n17522 , n4858 , n6895 );
    or g2503 ( n8899 , n9135 , n24194 );
    and g2504 ( n12753 , n6572 , n20710 );
    and g2505 ( n20617 , n10207 , n20084 );
    not g2506 ( n7297 , n860 );
    or g2507 ( n18964 , n10976 , n9757 );
    xnor g2508 ( n476 , n1689 , n20036 );
    xnor g2509 ( n21894 , n13512 , n10934 );
    or g2510 ( n24526 , n2047 , n1048 );
    xnor g2511 ( n11351 , n27087 , n24274 );
    or g2512 ( n1628 , n1750 , n21321 );
    not g2513 ( n16458 , n15564 );
    not g2514 ( n11248 , n12119 );
    xnor g2515 ( n1976 , n2242 , n6449 );
    xnor g2516 ( n4856 , n21843 , n14998 );
    not g2517 ( n7808 , n16025 );
    xnor g2518 ( n13683 , n9115 , n18586 );
    and g2519 ( n3980 , n11917 , n22193 );
    nor g2520 ( n13933 , n11919 , n26510 );
    or g2521 ( n10004 , n10992 , n25438 );
    xnor g2522 ( n26706 , n13688 , n25462 );
    or g2523 ( n9136 , n2268 , n19153 );
    not g2524 ( n7823 , n17180 );
    xnor g2525 ( n13001 , n22363 , n11848 );
    and g2526 ( n21170 , n3278 , n12710 );
    not g2527 ( n552 , n15090 );
    not g2528 ( n13401 , n22771 );
    or g2529 ( n2446 , n25620 , n17407 );
    xnor g2530 ( n14257 , n10567 , n14421 );
    xnor g2531 ( n19908 , n21774 , n20980 );
    not g2532 ( n22807 , n15654 );
    or g2533 ( n23507 , n25599 , n7232 );
    xnor g2534 ( n11974 , n3397 , n2889 );
    or g2535 ( n24995 , n9945 , n22227 );
    xnor g2536 ( n369 , n8244 , n21226 );
    or g2537 ( n26802 , n17296 , n21181 );
    not g2538 ( n16283 , n21385 );
    or g2539 ( n5373 , n18290 , n12875 );
    xnor g2540 ( n16321 , n16276 , n1348 );
    or g2541 ( n16020 , n8079 , n21736 );
    or g2542 ( n14948 , n19119 , n21833 );
    or g2543 ( n6197 , n4703 , n10926 );
    and g2544 ( n9278 , n18561 , n1488 );
    and g2545 ( n18085 , n22688 , n3474 );
    and g2546 ( n17996 , n26618 , n12658 );
    not g2547 ( n11243 , n12379 );
    or g2548 ( n25361 , n20780 , n7819 );
    not g2549 ( n27160 , n4196 );
    xnor g2550 ( n25927 , n6724 , n22405 );
    xnor g2551 ( n25948 , n11429 , n12315 );
    or g2552 ( n5912 , n26186 , n1028 );
    and g2553 ( n22621 , n24057 , n2910 );
    xnor g2554 ( n563 , n15896 , n12295 );
    xnor g2555 ( n9567 , n13925 , n21538 );
    not g2556 ( n21605 , n10614 );
    xnor g2557 ( n25802 , n16825 , n7020 );
    and g2558 ( n12026 , n11777 , n16644 );
    or g2559 ( n20396 , n26264 , n19454 );
    not g2560 ( n20734 , n22414 );
    or g2561 ( n10535 , n11455 , n14870 );
    or g2562 ( n24781 , n8922 , n10553 );
    xnor g2563 ( n8530 , n8520 , n20506 );
    not g2564 ( n11079 , n23303 );
    or g2565 ( n15434 , n26273 , n7186 );
    nor g2566 ( n21697 , n5318 , n7439 );
    and g2567 ( n620 , n19897 , n26987 );
    xnor g2568 ( n8163 , n25992 , n17298 );
    or g2569 ( n13665 , n4913 , n17525 );
    not g2570 ( n21422 , n3246 );
    xnor g2571 ( n14187 , n26426 , n12205 );
    nor g2572 ( n15168 , n19952 , n17444 );
    nor g2573 ( n8761 , n12863 , n13046 );
    xnor g2574 ( n8846 , n24488 , n24996 );
    and g2575 ( n11606 , n6758 , n24361 );
    and g2576 ( n15478 , n17884 , n24010 );
    xnor g2577 ( n14195 , n1822 , n1813 );
    not g2578 ( n21846 , n4426 );
    xnor g2579 ( n2813 , n20387 , n7077 );
    or g2580 ( n20685 , n12327 , n14447 );
    xnor g2581 ( n23694 , n8389 , n17454 );
    or g2582 ( n24159 , n7671 , n8354 );
    or g2583 ( n25703 , n17737 , n7744 );
    and g2584 ( n16588 , n4963 , n2818 );
    nor g2585 ( n9893 , n23272 , n14826 );
    and g2586 ( n12276 , n23250 , n11209 );
    or g2587 ( n8023 , n11652 , n12639 );
    not g2588 ( n2490 , n24884 );
    xnor g2589 ( n2228 , n5946 , n2445 );
    and g2590 ( n26087 , n19652 , n22610 );
    xnor g2591 ( n19933 , n14195 , n13533 );
    and g2592 ( n1940 , n21010 , n22678 );
    or g2593 ( n20510 , n25775 , n1397 );
    xnor g2594 ( n10349 , n24450 , n14533 );
    not g2595 ( n15787 , n8380 );
    nor g2596 ( n12245 , n10964 , n3314 );
    xnor g2597 ( n9406 , n15268 , n18737 );
    not g2598 ( n21564 , n4908 );
    and g2599 ( n21250 , n1858 , n24921 );
    nor g2600 ( n7453 , n2210 , n19863 );
    xnor g2601 ( n24039 , n1812 , n3233 );
    or g2602 ( n8764 , n19682 , n7041 );
    xnor g2603 ( n23852 , n939 , n2283 );
    xnor g2604 ( n27022 , n17345 , n11935 );
    not g2605 ( n6468 , n22772 );
    xnor g2606 ( n15691 , n2723 , n5806 );
    or g2607 ( n2912 , n22007 , n67 );
    not g2608 ( n4559 , n21497 );
    xnor g2609 ( n21254 , n9128 , n16816 );
    xnor g2610 ( n3842 , n13521 , n9420 );
    nor g2611 ( n9887 , n17447 , n12968 );
    or g2612 ( n25718 , n17977 , n11875 );
    xnor g2613 ( n4873 , n17986 , n3947 );
    or g2614 ( n7185 , n328 , n15490 );
    xnor g2615 ( n7298 , n19326 , n4855 );
    xnor g2616 ( n10217 , n4125 , n19477 );
    xnor g2617 ( n23000 , n12489 , n15753 );
    or g2618 ( n4567 , n8146 , n5285 );
    xnor g2619 ( n25267 , n663 , n24327 );
    and g2620 ( n18146 , n416 , n10981 );
    and g2621 ( n17773 , n16259 , n4394 );
    nor g2622 ( n7392 , n17606 , n24936 );
    or g2623 ( n17839 , n5948 , n15415 );
    not g2624 ( n10997 , n17371 );
    not g2625 ( n13967 , n23849 );
    nor g2626 ( n3514 , n17120 , n26510 );
    xnor g2627 ( n27028 , n3161 , n11630 );
    nor g2628 ( n13212 , n22637 , n12837 );
    or g2629 ( n1251 , n19898 , n8319 );
    or g2630 ( n7631 , n20342 , n4570 );
    xnor g2631 ( n20832 , n2415 , n19514 );
    or g2632 ( n2762 , n13975 , n14163 );
    xnor g2633 ( n8179 , n22776 , n15305 );
    nor g2634 ( n19018 , n11936 , n9531 );
    xnor g2635 ( n6746 , n9194 , n16913 );
    or g2636 ( n8879 , n13814 , n5815 );
    and g2637 ( n21534 , n17136 , n12662 );
    or g2638 ( n1260 , n6551 , n5527 );
    not g2639 ( n2653 , n4016 );
    and g2640 ( n25590 , n11764 , n10349 );
    xnor g2641 ( n22892 , n22549 , n16722 );
    and g2642 ( n21278 , n7961 , n20561 );
    not g2643 ( n11745 , n5026 );
    not g2644 ( n26793 , n9251 );
    xnor g2645 ( n14011 , n9964 , n5438 );
    and g2646 ( n10664 , n22051 , n22649 );
    not g2647 ( n10920 , n11592 );
    xnor g2648 ( n9728 , n3271 , n2757 );
    or g2649 ( n13416 , n26019 , n21407 );
    and g2650 ( n2839 , n19961 , n13077 );
    not g2651 ( n590 , n7304 );
    nor g2652 ( n6607 , n6243 , n4751 );
    xnor g2653 ( n15216 , n8614 , n23895 );
    and g2654 ( n1188 , n14495 , n25251 );
    and g2655 ( n19773 , n27026 , n351 );
    xnor g2656 ( n20709 , n4079 , n2758 );
    nor g2657 ( n2007 , n3057 , n7054 );
    and g2658 ( n1755 , n24513 , n845 );
    xnor g2659 ( n24042 , n12785 , n21762 );
    not g2660 ( n18925 , n7725 );
    nor g2661 ( n9628 , n23126 , n17369 );
    or g2662 ( n20912 , n23454 , n8647 );
    not g2663 ( n13530 , n14489 );
    xnor g2664 ( n2217 , n1739 , n4913 );
    xnor g2665 ( n12351 , n18621 , n4957 );
    xnor g2666 ( n10407 , n16362 , n6296 );
    nor g2667 ( n13646 , n2314 , n5407 );
    xnor g2668 ( n8653 , n21143 , n1842 );
    or g2669 ( n19966 , n16386 , n5739 );
    nor g2670 ( n2104 , n9693 , n12457 );
    nor g2671 ( n16787 , n23974 , n8309 );
    nor g2672 ( n14778 , n17906 , n4372 );
    xnor g2673 ( n4396 , n12869 , n822 );
    xnor g2674 ( n19338 , n8952 , n25240 );
    and g2675 ( n7029 , n26151 , n3221 );
    not g2676 ( n312 , n16906 );
    xnor g2677 ( n23851 , n17744 , n19033 );
    not g2678 ( n10995 , n18006 );
    not g2679 ( n25067 , n22309 );
    nor g2680 ( n19471 , n19618 , n18707 );
    xnor g2681 ( n13602 , n562 , n8219 );
    or g2682 ( n14144 , n22040 , n24707 );
    xnor g2683 ( n13759 , n9108 , n8873 );
    xnor g2684 ( n24742 , n20102 , n23751 );
    xnor g2685 ( n21299 , n12733 , n25972 );
    xnor g2686 ( n4146 , n4046 , n20668 );
    or g2687 ( n8976 , n21644 , n4426 );
    or g2688 ( n18605 , n1273 , n1070 );
    or g2689 ( n7150 , n24851 , n10711 );
    xnor g2690 ( n25426 , n13097 , n17225 );
    not g2691 ( n24058 , n19981 );
    xnor g2692 ( n17859 , n3914 , n23962 );
    or g2693 ( n8373 , n710 , n8398 );
    not g2694 ( n21930 , n15240 );
    not g2695 ( n14327 , n3920 );
    not g2696 ( n19085 , n6712 );
    xnor g2697 ( n20220 , n20777 , n2461 );
    xnor g2698 ( n13293 , n26464 , n20057 );
    xnor g2699 ( n24506 , n24323 , n8581 );
    or g2700 ( n13616 , n3439 , n1995 );
    not g2701 ( n17658 , n11329 );
    xnor g2702 ( n14446 , n11989 , n3526 );
    or g2703 ( n26533 , n21847 , n4980 );
    xnor g2704 ( n6551 , n19160 , n14835 );
    xnor g2705 ( n2966 , n13627 , n4847 );
    or g2706 ( n10827 , n26404 , n9751 );
    not g2707 ( n3601 , n16496 );
    not g2708 ( n15313 , n14314 );
    and g2709 ( n3575 , n8448 , n15892 );
    xnor g2710 ( n26098 , n2029 , n13776 );
    not g2711 ( n11652 , n9934 );
    xnor g2712 ( n5430 , n13878 , n2942 );
    not g2713 ( n20030 , n5340 );
    or g2714 ( n2068 , n14953 , n1581 );
    nor g2715 ( n5007 , n8232 , n20749 );
    and g2716 ( n10273 , n24653 , n10746 );
    or g2717 ( n24621 , n17959 , n25221 );
    not g2718 ( n12550 , n20499 );
    and g2719 ( n26173 , n15878 , n21011 );
    nor g2720 ( n7849 , n1009 , n18145 );
    xnor g2721 ( n20906 , n7855 , n20161 );
    and g2722 ( n17401 , n5796 , n25856 );
    xnor g2723 ( n11034 , n2994 , n25872 );
    or g2724 ( n5533 , n2432 , n20633 );
    and g2725 ( n1926 , n23916 , n6827 );
    xnor g2726 ( n7781 , n4887 , n6298 );
    not g2727 ( n12869 , n17186 );
    xnor g2728 ( n21298 , n12934 , n6349 );
    nor g2729 ( n3025 , n5624 , n13490 );
    and g2730 ( n4268 , n18368 , n12428 );
    nor g2731 ( n23502 , n11302 , n17213 );
    or g2732 ( n25010 , n21527 , n20509 );
    not g2733 ( n18767 , n2499 );
    or g2734 ( n8040 , n20345 , n9320 );
    not g2735 ( n25764 , n19741 );
    xnor g2736 ( n14849 , n632 , n23955 );
    or g2737 ( n1641 , n14000 , n7816 );
    or g2738 ( n16631 , n9365 , n13543 );
    xnor g2739 ( n2545 , n27041 , n3582 );
    not g2740 ( n19634 , n4812 );
    nor g2741 ( n20476 , n26876 , n3730 );
    not g2742 ( n2322 , n10728 );
    not g2743 ( n12720 , n24919 );
    nor g2744 ( n10893 , n17995 , n4222 );
    or g2745 ( n13554 , n294 , n23020 );
    or g2746 ( n884 , n26510 , n11246 );
    or g2747 ( n1902 , n24375 , n9942 );
    not g2748 ( n22454 , n9372 );
    and g2749 ( n23343 , n5790 , n14398 );
    nor g2750 ( n7189 , n2151 , n26425 );
    and g2751 ( n4433 , n574 , n24689 );
    or g2752 ( n21333 , n2979 , n24764 );
    nor g2753 ( n11725 , n3173 , n25393 );
    and g2754 ( n18633 , n4625 , n9523 );
    or g2755 ( n1962 , n27012 , n1737 );
    nor g2756 ( n19619 , n839 , n15709 );
    or g2757 ( n3404 , n13292 , n21911 );
    or g2758 ( n26855 , n19076 , n3903 );
    and g2759 ( n21758 , n4351 , n25153 );
    and g2760 ( n23037 , n23227 , n16315 );
    nor g2761 ( n18077 , n11314 , n7689 );
    or g2762 ( n19503 , n9157 , n23931 );
    xnor g2763 ( n10979 , n6353 , n12391 );
    and g2764 ( n25396 , n26628 , n26960 );
    or g2765 ( n5080 , n23658 , n17121 );
    not g2766 ( n12405 , n2841 );
    or g2767 ( n2074 , n23416 , n18597 );
    not g2768 ( n14725 , n2394 );
    not g2769 ( n11146 , n26713 );
    or g2770 ( n23516 , n14066 , n23432 );
    nor g2771 ( n20088 , n9490 , n23693 );
    xnor g2772 ( n26935 , n26837 , n13251 );
    not g2773 ( n1994 , n7652 );
    nor g2774 ( n16030 , n5960 , n13490 );
    and g2775 ( n5209 , n17965 , n1744 );
    nor g2776 ( n2257 , n6841 , n8439 );
    and g2777 ( n25981 , n21606 , n26422 );
    or g2778 ( n13690 , n23573 , n6637 );
    not g2779 ( n246 , n626 );
    nor g2780 ( n27092 , n9940 , n8013 );
    nor g2781 ( n11438 , n15432 , n18883 );
    and g2782 ( n6391 , n15905 , n27118 );
    nor g2783 ( n9384 , n9497 , n23751 );
    not g2784 ( n16942 , n23220 );
    nor g2785 ( n14302 , n12042 , n11308 );
    not g2786 ( n13389 , n7692 );
    and g2787 ( n21576 , n11460 , n27056 );
    xnor g2788 ( n10246 , n655 , n6397 );
    xnor g2789 ( n6626 , n22198 , n5337 );
    xnor g2790 ( n6876 , n3373 , n2892 );
    and g2791 ( n13839 , n24355 , n21935 );
    xnor g2792 ( n15435 , n9058 , n20286 );
    nor g2793 ( n7055 , n15220 , n3846 );
    not g2794 ( n302 , n23277 );
    and g2795 ( n6874 , n3170 , n23699 );
    and g2796 ( n2070 , n18658 , n15035 );
    and g2797 ( n19561 , n17861 , n24190 );
    and g2798 ( n26082 , n25855 , n26461 );
    and g2799 ( n26949 , n13783 , n13590 );
    and g2800 ( n20392 , n2621 , n2364 );
    xnor g2801 ( n14353 , n25020 , n14607 );
    or g2802 ( n21048 , n1815 , n26735 );
    buf g2803 ( n26460 , n5703 );
    not g2804 ( n11501 , n18229 );
    or g2805 ( n3182 , n2384 , n18873 );
    xnor g2806 ( n13776 , n18765 , n21975 );
    or g2807 ( n9589 , n24462 , n6748 );
    and g2808 ( n7932 , n1497 , n4184 );
    not g2809 ( n20216 , n8540 );
    or g2810 ( n20793 , n19531 , n26872 );
    or g2811 ( n25728 , n10761 , n3985 );
    or g2812 ( n22228 , n12955 , n5220 );
    or g2813 ( n25339 , n7923 , n5998 );
    xnor g2814 ( n23299 , n16687 , n6449 );
    or g2815 ( n3787 , n18192 , n9473 );
    or g2816 ( n12462 , n6650 , n11260 );
    not g2817 ( n6195 , n18630 );
    or g2818 ( n3683 , n26738 , n6666 );
    xnor g2819 ( n470 , n11136 , n6435 );
    and g2820 ( n16086 , n7092 , n24486 );
    or g2821 ( n8852 , n11425 , n9967 );
    xnor g2822 ( n809 , n23077 , n12266 );
    and g2823 ( n6979 , n8275 , n7220 );
    or g2824 ( n7114 , n21450 , n24821 );
    or g2825 ( n11874 , n682 , n14811 );
    or g2826 ( n11645 , n3853 , n23372 );
    xnor g2827 ( n242 , n5477 , n6433 );
    not g2828 ( n19493 , n16261 );
    and g2829 ( n4140 , n26564 , n7471 );
    xnor g2830 ( n12916 , n20065 , n2184 );
    xnor g2831 ( n22557 , n9354 , n3722 );
    xnor g2832 ( n4449 , n21537 , n18274 );
    or g2833 ( n15063 , n22261 , n10117 );
    or g2834 ( n14524 , n19494 , n2387 );
    nor g2835 ( n4703 , n26536 , n19607 );
    or g2836 ( n19651 , n4887 , n5045 );
    xnor g2837 ( n25887 , n6122 , n23200 );
    not g2838 ( n21083 , n8399 );
    not g2839 ( n13035 , n17982 );
    not g2840 ( n18994 , n5582 );
    xnor g2841 ( n23735 , n2320 , n26053 );
    nor g2842 ( n4771 , n3472 , n15790 );
    or g2843 ( n9870 , n11542 , n7057 );
    not g2844 ( n2462 , n25617 );
    or g2845 ( n22941 , n11171 , n26026 );
    xnor g2846 ( n10540 , n4430 , n3218 );
    xnor g2847 ( n3630 , n25074 , n12956 );
    xnor g2848 ( n18399 , n10666 , n19856 );
    and g2849 ( n25552 , n16105 , n6118 );
    and g2850 ( n11789 , n8094 , n11051 );
    xnor g2851 ( n1394 , n10611 , n24879 );
    or g2852 ( n20010 , n18203 , n15910 );
    and g2853 ( n12937 , n6110 , n16990 );
    or g2854 ( n26221 , n1783 , n2587 );
    xnor g2855 ( n12733 , n3028 , n13965 );
    and g2856 ( n5811 , n8614 , n21162 );
    xnor g2857 ( n18522 , n22554 , n25381 );
    and g2858 ( n21610 , n2743 , n1584 );
    xor g2859 ( n1386 , n13032 , n12188 );
    nor g2860 ( n7027 , n1777 , n4812 );
    or g2861 ( n19014 , n4039 , n8742 );
    xnor g2862 ( n1470 , n15041 , n26553 );
    or g2863 ( n11825 , n21936 , n46 );
    or g2864 ( n17698 , n10191 , n26463 );
    or g2865 ( n8478 , n13370 , n25644 );
    xnor g2866 ( n3012 , n3071 , n1305 );
    and g2867 ( n805 , n23090 , n3353 );
    or g2868 ( n2848 , n13909 , n520 );
    or g2869 ( n15863 , n23441 , n9926 );
    xnor g2870 ( n4775 , n25187 , n11619 );
    xnor g2871 ( n17149 , n15073 , n19814 );
    nor g2872 ( n16593 , n14114 , n14111 );
    and g2873 ( n4880 , n16033 , n7121 );
    and g2874 ( n3341 , n1969 , n20729 );
    or g2875 ( n2730 , n1689 , n9450 );
    xnor g2876 ( n27049 , n20077 , n19494 );
    xnor g2877 ( n2401 , n4706 , n905 );
    or g2878 ( n12394 , n24461 , n26095 );
    and g2879 ( n10308 , n6845 , n4211 );
    or g2880 ( n16650 , n1138 , n17000 );
    or g2881 ( n9690 , n9110 , n25442 );
    or g2882 ( n26500 , n18521 , n3802 );
    and g2883 ( n12807 , n11445 , n25587 );
    or g2884 ( n24946 , n3013 , n19436 );
    xnor g2885 ( n4958 , n2718 , n9291 );
    and g2886 ( n1645 , n19675 , n24173 );
    or g2887 ( n66 , n6677 , n25026 );
    or g2888 ( n25722 , n24650 , n13033 );
    or g2889 ( n3362 , n25524 , n16234 );
    not g2890 ( n2268 , n12593 );
    or g2891 ( n16157 , n15827 , n15073 );
    nor g2892 ( n9824 , n15251 , n4422 );
    or g2893 ( n9921 , n19321 , n19737 );
    xnor g2894 ( n803 , n19311 , n992 );
    xnor g2895 ( n6492 , n24789 , n19252 );
    and g2896 ( n20456 , n18155 , n16027 );
    xnor g2897 ( n9827 , n8142 , n22835 );
    xnor g2898 ( n8330 , n6631 , n7339 );
    nor g2899 ( n16534 , n13577 , n12341 );
    xnor g2900 ( n18965 , n19905 , n2547 );
    not g2901 ( n22507 , n19425 );
    not g2902 ( n8077 , n9240 );
    xnor g2903 ( n5674 , n6041 , n14550 );
    xnor g2904 ( n11235 , n3401 , n1249 );
    or g2905 ( n7485 , n16635 , n24450 );
    or g2906 ( n22790 , n25916 , n18570 );
    and g2907 ( n4789 , n5029 , n23263 );
    xnor g2908 ( n9190 , n13912 , n11980 );
    or g2909 ( n18106 , n8 , n19678 );
    xnor g2910 ( n16839 , n21713 , n26835 );
    not g2911 ( n13803 , n8479 );
    xnor g2912 ( n13727 , n9974 , n24138 );
    xnor g2913 ( n16054 , n5542 , n22372 );
    xnor g2914 ( n4148 , n23039 , n4590 );
    xnor g2915 ( n2253 , n21508 , n10183 );
    or g2916 ( n17527 , n17018 , n26968 );
    or g2917 ( n25559 , n8678 , n3882 );
    not g2918 ( n14757 , n22864 );
    xnor g2919 ( n4482 , n8456 , n5605 );
    nor g2920 ( n14383 , n22247 , n21126 );
    xnor g2921 ( n1350 , n16970 , n11287 );
    and g2922 ( n27024 , n9729 , n4985 );
    xnor g2923 ( n20755 , n1149 , n8349 );
    or g2924 ( n22522 , n25119 , n3719 );
    or g2925 ( n9773 , n20245 , n8006 );
    or g2926 ( n753 , n20479 , n9222 );
    not g2927 ( n2911 , n19285 );
    and g2928 ( n22307 , n22565 , n5656 );
    and g2929 ( n23316 , n20040 , n16555 );
    and g2930 ( n26519 , n5400 , n9512 );
    nor g2931 ( n7378 , n2659 , n1941 );
    or g2932 ( n12326 , n725 , n24804 );
    or g2933 ( n24921 , n4279 , n13566 );
    and g2934 ( n14461 , n1515 , n19207 );
    nor g2935 ( n9081 , n1689 , n17095 );
    or g2936 ( n20234 , n5075 , n25768 );
    nor g2937 ( n18028 , n23359 , n15454 );
    and g2938 ( n6699 , n26998 , n3592 );
    or g2939 ( n17072 , n2104 , n10609 );
    xnor g2940 ( n14767 , n18015 , n3027 );
    xnor g2941 ( n10280 , n23996 , n5685 );
    not g2942 ( n733 , n5704 );
    xnor g2943 ( n17071 , n19048 , n25007 );
    not g2944 ( n26421 , n2383 );
    buf g2945 ( n21263 , n12211 );
    or g2946 ( n7789 , n9583 , n15566 );
    xnor g2947 ( n13837 , n22342 , n16993 );
    and g2948 ( n1879 , n23304 , n1465 );
    or g2949 ( n9167 , n21481 , n14867 );
    or g2950 ( n4209 , n5230 , n9682 );
    or g2951 ( n21831 , n9924 , n26216 );
    not g2952 ( n586 , n3614 );
    or g2953 ( n15609 , n12636 , n4633 );
    or g2954 ( n991 , n778 , n23769 );
    or g2955 ( n5515 , n19630 , n3361 );
    not g2956 ( n14710 , n22764 );
    xnor g2957 ( n1119 , n18605 , n24144 );
    and g2958 ( n10194 , n11100 , n22513 );
    nor g2959 ( n6650 , n25781 , n2155 );
    xnor g2960 ( n15894 , n12019 , n17585 );
    not g2961 ( n6764 , n15780 );
    not g2962 ( n18173 , n6659 );
    and g2963 ( n18056 , n17160 , n5927 );
    and g2964 ( n3196 , n13882 , n8058 );
    xnor g2965 ( n4930 , n11309 , n26452 );
    xnor g2966 ( n1907 , n13951 , n12507 );
    or g2967 ( n26567 , n13497 , n22631 );
    xnor g2968 ( n21253 , n17124 , n15979 );
    or g2969 ( n15305 , n27 , n25973 );
    xnor g2970 ( n9864 , n4256 , n20946 );
    or g2971 ( n9667 , n4383 , n3808 );
    xnor g2972 ( n26330 , n21544 , n18924 );
    xnor g2973 ( n4269 , n23819 , n25370 );
    xnor g2974 ( n27036 , n5156 , n13460 );
    or g2975 ( n797 , n1103 , n18389 );
    and g2976 ( n18524 , n19105 , n9010 );
    not g2977 ( n333 , n2568 );
    or g2978 ( n7495 , n4893 , n21451 );
    or g2979 ( n14088 , n405 , n13842 );
    and g2980 ( n25885 , n23327 , n25945 );
    or g2981 ( n12206 , n1680 , n479 );
    and g2982 ( n14167 , n11536 , n8684 );
    and g2983 ( n23380 , n21599 , n26324 );
    not g2984 ( n3116 , n8638 );
    not g2985 ( n16751 , n16426 );
    and g2986 ( n21064 , n600 , n12497 );
    or g2987 ( n14490 , n19551 , n2705 );
    xnor g2988 ( n9686 , n23580 , n26350 );
    or g2989 ( n18879 , n7338 , n22355 );
    or g2990 ( n21518 , n24649 , n14719 );
    or g2991 ( n6960 , n13061 , n23552 );
    and g2992 ( n14041 , n17394 , n9727 );
    not g2993 ( n16531 , n4514 );
    not g2994 ( n20100 , n8687 );
    and g2995 ( n5196 , n16485 , n14745 );
    or g2996 ( n14553 , n3139 , n23037 );
    or g2997 ( n18109 , n18775 , n20825 );
    xnor g2998 ( n13447 , n20950 , n15376 );
    or g2999 ( n4985 , n57 , n7539 );
    nor g3000 ( n14479 , n5521 , n1803 );
    or g3001 ( n15027 , n15602 , n3690 );
    and g3002 ( n24388 , n23832 , n19238 );
    not g3003 ( n4185 , n23939 );
    nor g3004 ( n1373 , n27175 , n5474 );
    or g3005 ( n12062 , n19006 , n22180 );
    or g3006 ( n23223 , n12612 , n14048 );
    and g3007 ( n2647 , n22148 , n10566 );
    and g3008 ( n9276 , n11368 , n8939 );
    xnor g3009 ( n24167 , n24817 , n8896 );
    and g3010 ( n15526 , n12114 , n25796 );
    or g3011 ( n9232 , n23895 , n8491 );
    or g3012 ( n25078 , n17558 , n26403 );
    and g3013 ( n14930 , n16654 , n7824 );
    xnor g3014 ( n12610 , n15023 , n13113 );
    or g3015 ( n11868 , n1373 , n1080 );
    xnor g3016 ( n23488 , n21817 , n9057 );
    xnor g3017 ( n15282 , n3798 , n23140 );
    nor g3018 ( n26907 , n18079 , n21460 );
    or g3019 ( n2225 , n6499 , n5002 );
    nor g3020 ( n10078 , n18792 , n15417 );
    or g3021 ( n25672 , n24310 , n16116 );
    or g3022 ( n12376 , n19899 , n18608 );
    xnor g3023 ( n15496 , n26737 , n12975 );
    nor g3024 ( n15249 , n7457 , n32 );
    xnor g3025 ( n12761 , n1685 , n3785 );
    nor g3026 ( n21229 , n9888 , n3827 );
    and g3027 ( n18896 , n18274 , n24202 );
    and g3028 ( n6325 , n10422 , n19383 );
    not g3029 ( n15507 , n12236 );
    xnor g3030 ( n16092 , n14197 , n12808 );
    or g3031 ( n4666 , n5612 , n3144 );
    xnor g3032 ( n3132 , n2941 , n655 );
    not g3033 ( n12769 , n19219 );
    not g3034 ( n6199 , n16423 );
    and g3035 ( n5665 , n19992 , n3427 );
    or g3036 ( n4447 , n19640 , n13916 );
    or g3037 ( n7790 , n17234 , n7993 );
    and g3038 ( n51 , n25943 , n12118 );
    or g3039 ( n7283 , n19616 , n13359 );
    xnor g3040 ( n23628 , n24357 , n16346 );
    and g3041 ( n19498 , n15348 , n9722 );
    xnor g3042 ( n6974 , n4753 , n3366 );
    xnor g3043 ( n19376 , n23061 , n7305 );
    or g3044 ( n19693 , n3685 , n19821 );
    xnor g3045 ( n16662 , n7019 , n10665 );
    xnor g3046 ( n17064 , n20987 , n7635 );
    not g3047 ( n21772 , n8763 );
    xnor g3048 ( n25449 , n8230 , n21024 );
    not g3049 ( n13737 , n23170 );
    xnor g3050 ( n13303 , n17374 , n9006 );
    or g3051 ( n6487 , n24168 , n1617 );
    not g3052 ( n20275 , n16832 );
    and g3053 ( n4600 , n8384 , n11067 );
    nor g3054 ( n18894 , n16830 , n20032 );
    and g3055 ( n4296 , n13402 , n20322 );
    nor g3056 ( n5054 , n23290 , n20185 );
    xnor g3057 ( n21859 , n20575 , n23725 );
    or g3058 ( n22184 , n8098 , n22344 );
    nor g3059 ( n13874 , n22183 , n25595 );
    xnor g3060 ( n9442 , n8952 , n7841 );
    not g3061 ( n1230 , n13123 );
    not g3062 ( n24947 , n3909 );
    xnor g3063 ( n11116 , n7304 , n10095 );
    or g3064 ( n17429 , n27052 , n4944 );
    xnor g3065 ( n23655 , n16831 , n10582 );
    xnor g3066 ( n885 , n7593 , n5101 );
    xnor g3067 ( n3973 , n12592 , n10267 );
    xnor g3068 ( n5701 , n16150 , n14010 );
    xnor g3069 ( n16073 , n22012 , n8688 );
    not g3070 ( n11694 , n7008 );
    or g3071 ( n15047 , n18613 , n5526 );
    xnor g3072 ( n26317 , n24858 , n18763 );
    xnor g3073 ( n27139 , n18795 , n18854 );
    not g3074 ( n17559 , n26098 );
    xnor g3075 ( n22153 , n21836 , n18020 );
    or g3076 ( n21464 , n12132 , n239 );
    and g3077 ( n18816 , n21895 , n4303 );
    or g3078 ( n15112 , n14995 , n11430 );
    or g3079 ( n7720 , n6601 , n3600 );
    and g3080 ( n5957 , n24136 , n18806 );
    xnor g3081 ( n10111 , n10566 , n16108 );
    xnor g3082 ( n25958 , n16609 , n7949 );
    not g3083 ( n13422 , n25586 );
    not g3084 ( n7627 , n15975 );
    not g3085 ( n13357 , n5386 );
    xnor g3086 ( n16176 , n130 , n5247 );
    or g3087 ( n16069 , n25037 , n9183 );
    nor g3088 ( n20471 , n2145 , n5521 );
    not g3089 ( n9909 , n20361 );
    xnor g3090 ( n957 , n7957 , n12412 );
    and g3091 ( n12335 , n26158 , n8262 );
    and g3092 ( n282 , n1235 , n23700 );
    and g3093 ( n7582 , n709 , n3337 );
    and g3094 ( n7098 , n3522 , n25338 );
    and g3095 ( n26944 , n7434 , n23025 );
    not g3096 ( n18587 , n13885 );
    xnor g3097 ( n19039 , n16094 , n26660 );
    and g3098 ( n26247 , n21777 , n4685 );
    and g3099 ( n3384 , n2420 , n23807 );
    xnor g3100 ( n13197 , n1606 , n13607 );
    or g3101 ( n8544 , n17252 , n22338 );
    and g3102 ( n14681 , n1283 , n2427 );
    or g3103 ( n14929 , n8180 , n5734 );
    xnor g3104 ( n4670 , n21285 , n12907 );
    or g3105 ( n6017 , n15361 , n3044 );
    xnor g3106 ( n2532 , n5244 , n255 );
    and g3107 ( n516 , n10796 , n15653 );
    or g3108 ( n6955 , n17617 , n16426 );
    and g3109 ( n8797 , n16427 , n17888 );
    xnor g3110 ( n14544 , n10664 , n14606 );
    or g3111 ( n7334 , n8835 , n19544 );
    or g3112 ( n6854 , n26892 , n17200 );
    nor g3113 ( n1178 , n7072 , n9851 );
    xnor g3114 ( n11710 , n6322 , n16422 );
    xnor g3115 ( n25133 , n4637 , n17074 );
    and g3116 ( n14209 , n8459 , n404 );
    nor g3117 ( n24819 , n21469 , n16017 );
    or g3118 ( n20813 , n9716 , n1495 );
    or g3119 ( n22693 , n21373 , n13182 );
    xnor g3120 ( n10222 , n148 , n2113 );
    and g3121 ( n20050 , n13256 , n25780 );
    xnor g3122 ( n18148 , n15091 , n26693 );
    not g3123 ( n728 , n21155 );
    xnor g3124 ( n11104 , n12470 , n11455 );
    and g3125 ( n6520 , n24377 , n20514 );
    xnor g3126 ( n9759 , n23835 , n2950 );
    xnor g3127 ( n15291 , n11609 , n26386 );
    nor g3128 ( n1289 , n10357 , n20284 );
    not g3129 ( n19738 , n10228 );
    and g3130 ( n14029 , n24490 , n3930 );
    not g3131 ( n9227 , n21723 );
    or g3132 ( n13272 , n23156 , n26813 );
    nor g3133 ( n4503 , n23290 , n15742 );
    not g3134 ( n8739 , n23755 );
    xnor g3135 ( n6847 , n18824 , n2596 );
    or g3136 ( n19206 , n1958 , n1187 );
    not g3137 ( n11144 , n18105 );
    not g3138 ( n396 , n9396 );
    or g3139 ( n7577 , n6659 , n20384 );
    and g3140 ( n18872 , n21984 , n6255 );
    xnor g3141 ( n11765 , n21850 , n17351 );
    and g3142 ( n9183 , n9573 , n17480 );
    not g3143 ( n1956 , n337 );
    xnor g3144 ( n25006 , n26148 , n26323 );
    xnor g3145 ( n19780 , n7165 , n16099 );
    xnor g3146 ( n9807 , n6925 , n10505 );
    not g3147 ( n12644 , n18672 );
    not g3148 ( n7923 , n9380 );
    and g3149 ( n9465 , n7237 , n15087 );
    and g3150 ( n26256 , n25333 , n3847 );
    nor g3151 ( n22606 , n7566 , n586 );
    nor g3152 ( n29 , n16738 , n12860 );
    and g3153 ( n12847 , n3460 , n11452 );
    or g3154 ( n21165 , n13719 , n6710 );
    xnor g3155 ( n20366 , n23381 , n21417 );
    and g3156 ( n10069 , n9697 , n19251 );
    nor g3157 ( n14339 , n14710 , n2416 );
    or g3158 ( n22374 , n709 , n3337 );
    xnor g3159 ( n13096 , n9334 , n13045 );
    not g3160 ( n16750 , n20072 );
    xnor g3161 ( n14198 , n4080 , n16394 );
    or g3162 ( n11602 , n3977 , n4136 );
    xnor g3163 ( n14036 , n15526 , n4382 );
    xnor g3164 ( n15126 , n20254 , n14687 );
    xnor g3165 ( n16051 , n23837 , n22092 );
    or g3166 ( n4469 , n19838 , n11083 );
    nor g3167 ( n14113 , n14923 , n12050 );
    nor g3168 ( n20775 , n5976 , n2694 );
    and g3169 ( n13295 , n206 , n13020 );
    xnor g3170 ( n18312 , n18068 , n20826 );
    xnor g3171 ( n14968 , n18496 , n25331 );
    xnor g3172 ( n637 , n11108 , n18988 );
    buf g3173 ( n21969 , n12417 );
    or g3174 ( n1031 , n1186 , n12317 );
    or g3175 ( n6619 , n31 , n16065 );
    not g3176 ( n5716 , n20958 );
    or g3177 ( n3039 , n22179 , n1944 );
    not g3178 ( n4862 , n20336 );
    and g3179 ( n22109 , n8984 , n62 );
    nor g3180 ( n26814 , n7974 , n8399 );
    and g3181 ( n15994 , n12925 , n8919 );
    or g3182 ( n25341 , n26580 , n5428 );
    xnor g3183 ( n24636 , n12796 , n21809 );
    and g3184 ( n257 , n1270 , n4428 );
    nor g3185 ( n4486 , n19277 , n23430 );
    and g3186 ( n7612 , n16495 , n12401 );
    and g3187 ( n14165 , n8433 , n2292 );
    nor g3188 ( n25928 , n22215 , n26350 );
    or g3189 ( n13519 , n16709 , n22771 );
    or g3190 ( n27152 , n3155 , n14697 );
    nor g3191 ( n25621 , n16910 , n15975 );
    nor g3192 ( n10381 , n27199 , n4003 );
    xnor g3193 ( n16379 , n8460 , n10064 );
    or g3194 ( n22555 , n23298 , n19131 );
    or g3195 ( n9209 , n12341 , n5727 );
    nor g3196 ( n19613 , n187 , n10549 );
    xnor g3197 ( n4121 , n14680 , n20359 );
    xnor g3198 ( n24961 , n7480 , n13347 );
    nor g3199 ( n19813 , n21876 , n18121 );
    xnor g3200 ( n11751 , n19049 , n14097 );
    xnor g3201 ( n20199 , n8052 , n24618 );
    or g3202 ( n8429 , n10499 , n2248 );
    not g3203 ( n2842 , n6678 );
    xnor g3204 ( n14723 , n6954 , n17730 );
    xnor g3205 ( n20076 , n16891 , n21602 );
    or g3206 ( n11699 , n20334 , n13493 );
    and g3207 ( n7498 , n8213 , n26657 );
    xnor g3208 ( n10733 , n2291 , n25629 );
    xnor g3209 ( n27079 , n9153 , n11053 );
    or g3210 ( n7451 , n18516 , n26714 );
    xnor g3211 ( n6281 , n26691 , n7563 );
    xnor g3212 ( n4943 , n11088 , n22843 );
    not g3213 ( n13498 , n14299 );
    xnor g3214 ( n11336 , n14346 , n26797 );
    nor g3215 ( n26442 , n21929 , n9575 );
    xnor g3216 ( n2041 , n648 , n7271 );
    xor g3217 ( n13511 , n8163 , n13752 );
    not g3218 ( n3397 , n1455 );
    not g3219 ( n22077 , n15894 );
    not g3220 ( n23720 , n822 );
    and g3221 ( n3612 , n20009 , n23980 );
    or g3222 ( n999 , n4602 , n8250 );
    or g3223 ( n25508 , n24949 , n789 );
    nor g3224 ( n18190 , n6372 , n11784 );
    xnor g3225 ( n273 , n12652 , n21309 );
    or g3226 ( n3217 , n6993 , n15706 );
    or g3227 ( n25233 , n21350 , n18049 );
    and g3228 ( n13594 , n5934 , n25517 );
    not g3229 ( n1728 , n21956 );
    or g3230 ( n21727 , n4502 , n16618 );
    or g3231 ( n13758 , n16678 , n25384 );
    not g3232 ( n14455 , n13521 );
    nor g3233 ( n25190 , n18585 , n12993 );
    and g3234 ( n7744 , n24505 , n12460 );
    and g3235 ( n5829 , n16609 , n22666 );
    xnor g3236 ( n11134 , n13147 , n12730 );
    xnor g3237 ( n10633 , n3562 , n19694 );
    xnor g3238 ( n23284 , n3846 , n15220 );
    not g3239 ( n9770 , n9222 );
    nor g3240 ( n20399 , n25846 , n4800 );
    and g3241 ( n2337 , n6557 , n17673 );
    not g3242 ( n10469 , n4245 );
    xnor g3243 ( n18570 , n22378 , n24630 );
    not g3244 ( n11337 , n11070 );
    and g3245 ( n3898 , n18476 , n27042 );
    xnor g3246 ( n12216 , n23083 , n8724 );
    xnor g3247 ( n21513 , n25036 , n9983 );
    not g3248 ( n16234 , n3959 );
    not g3249 ( n25461 , n2191 );
    xnor g3250 ( n12838 , n17333 , n19247 );
    or g3251 ( n1341 , n21674 , n5090 );
    or g3252 ( n8435 , n13459 , n17183 );
    nor g3253 ( n10770 , n14408 , n3486 );
    or g3254 ( n9235 , n21538 , n11335 );
    xor g3255 ( n6315 , n11378 , n3515 );
    xnor g3256 ( n20069 , n8124 , n24100 );
    or g3257 ( n12738 , n329 , n21735 );
    or g3258 ( n21379 , n25854 , n9379 );
    nor g3259 ( n8228 , n13490 , n7751 );
    or g3260 ( n21761 , n4752 , n7674 );
    or g3261 ( n20156 , n6273 , n21206 );
    or g3262 ( n6101 , n10687 , n5910 );
    not g3263 ( n21055 , n13031 );
    and g3264 ( n4385 , n8928 , n9231 );
    not g3265 ( n3365 , n17003 );
    and g3266 ( n14789 , n658 , n25339 );
    nor g3267 ( n18952 , n20205 , n2218 );
    xnor g3268 ( n19925 , n8774 , n22198 );
    and g3269 ( n16491 , n6537 , n21311 );
    and g3270 ( n20928 , n7770 , n13413 );
    or g3271 ( n4888 , n13681 , n17307 );
    xnor g3272 ( n24514 , n15127 , n3846 );
    or g3273 ( n19892 , n976 , n17050 );
    and g3274 ( n17752 , n25299 , n17907 );
    xnor g3275 ( n8111 , n2858 , n5521 );
    or g3276 ( n9774 , n15939 , n18927 );
    or g3277 ( n24459 , n3275 , n2800 );
    and g3278 ( n17004 , n11113 , n5917 );
    xnor g3279 ( n3176 , n16291 , n13044 );
    and g3280 ( n6032 , n12035 , n2609 );
    nor g3281 ( n11147 , n17826 , n10554 );
    nor g3282 ( n421 , n4469 , n5987 );
    xnor g3283 ( n16638 , n9912 , n7547 );
    xnor g3284 ( n20008 , n11615 , n8052 );
    not g3285 ( n23645 , n7460 );
    and g3286 ( n3119 , n891 , n17364 );
    not g3287 ( n11583 , n20151 );
    not g3288 ( n17444 , n9219 );
    or g3289 ( n22686 , n18625 , n17249 );
    and g3290 ( n12142 , n6100 , n19965 );
    and g3291 ( n17247 , n19743 , n2683 );
    nor g3292 ( n6124 , n3577 , n25171 );
    xnor g3293 ( n12438 , n851 , n5255 );
    nor g3294 ( n11075 , n21749 , n26744 );
    not g3295 ( n23008 , n20296 );
    not g3296 ( n1406 , n20235 );
    xnor g3297 ( n12540 , n10726 , n23481 );
    or g3298 ( n10172 , n9424 , n15413 );
    or g3299 ( n21112 , n19144 , n9170 );
    and g3300 ( n7553 , n26722 , n15074 );
    or g3301 ( n20194 , n2792 , n21113 );
    or g3302 ( n26534 , n20134 , n9192 );
    xnor g3303 ( n16060 , n25219 , n21425 );
    xnor g3304 ( n19627 , n7184 , n23107 );
    not g3305 ( n18203 , n19245 );
    and g3306 ( n16533 , n8231 , n13565 );
    not g3307 ( n22766 , n8774 );
    xnor g3308 ( n7408 , n7029 , n18372 );
    or g3309 ( n4527 , n10837 , n23890 );
    xnor g3310 ( n24712 , n26235 , n22439 );
    or g3311 ( n21419 , n8334 , n19946 );
    xnor g3312 ( n1527 , n20683 , n17882 );
    xnor g3313 ( n10454 , n23590 , n510 );
    not g3314 ( n20134 , n5337 );
    xnor g3315 ( n20285 , n4626 , n604 );
    or g3316 ( n6836 , n17256 , n14693 );
    or g3317 ( n13496 , n7586 , n2467 );
    not g3318 ( n16602 , n6422 );
    nor g3319 ( n18728 , n17052 , n439 );
    and g3320 ( n12298 , n22309 , n10711 );
    and g3321 ( n6157 , n24060 , n11345 );
    xnor g3322 ( n1008 , n9468 , n15241 );
    or g3323 ( n1149 , n20865 , n517 );
    or g3324 ( n14798 , n22987 , n13357 );
    xnor g3325 ( n8849 , n26468 , n12838 );
    and g3326 ( n3435 , n26825 , n1271 );
    or g3327 ( n26975 , n6023 , n20649 );
    or g3328 ( n149 , n19462 , n8131 );
    xnor g3329 ( n7260 , n25367 , n20163 );
    not g3330 ( n19149 , n3366 );
    and g3331 ( n11863 , n3268 , n14062 );
    xnor g3332 ( n8240 , n1720 , n6543 );
    xnor g3333 ( n6062 , n8827 , n1881 );
    nor g3334 ( n27033 , n4199 , n11118 );
    not g3335 ( n8210 , n619 );
    xor g3336 ( n22120 , n15891 , n9493 );
    not g3337 ( n7223 , n20291 );
    and g3338 ( n20683 , n24174 , n22145 );
    and g3339 ( n17621 , n22094 , n21920 );
    xnor g3340 ( n15625 , n6222 , n9744 );
    not g3341 ( n15423 , n5416 );
    xnor g3342 ( n8751 , n10228 , n11473 );
    and g3343 ( n13193 , n25151 , n214 );
    not g3344 ( n24645 , n4834 );
    xnor g3345 ( n10565 , n19975 , n3121 );
    xnor g3346 ( n25033 , n13360 , n13124 );
    or g3347 ( n4842 , n15604 , n18001 );
    xnor g3348 ( n16423 , n20499 , n18689 );
    or g3349 ( n19492 , n10894 , n11484 );
    and g3350 ( n16365 , n878 , n2123 );
    not g3351 ( n1850 , n10970 );
    or g3352 ( n4635 , n18789 , n1535 );
    xnor g3353 ( n4225 , n14974 , n11246 );
    or g3354 ( n11511 , n975 , n25618 );
    not g3355 ( n776 , n18880 );
    and g3356 ( n13467 , n26493 , n4842 );
    xnor g3357 ( n7802 , n20544 , n12071 );
    xnor g3358 ( n24315 , n17760 , n25373 );
    and g3359 ( n23445 , n21232 , n7471 );
    or g3360 ( n7883 , n13286 , n26080 );
    and g3361 ( n16255 , n19449 , n22757 );
    xnor g3362 ( n15839 , n26399 , n3710 );
    xnor g3363 ( n11136 , n9545 , n2232 );
    and g3364 ( n3729 , n2644 , n289 );
    and g3365 ( n3734 , n1278 , n22695 );
    or g3366 ( n11202 , n15293 , n24644 );
    xnor g3367 ( n22413 , n12646 , n19725 );
    and g3368 ( n26402 , n13734 , n6019 );
    or g3369 ( n3375 , n18013 , n12926 );
    or g3370 ( n11762 , n4227 , n11050 );
    not g3371 ( n10807 , n3827 );
    or g3372 ( n19510 , n5822 , n7963 );
    xnor g3373 ( n11842 , n16857 , n26131 );
    and g3374 ( n25216 , n19506 , n1897 );
    not g3375 ( n6750 , n16439 );
    or g3376 ( n6890 , n2380 , n25253 );
    or g3377 ( n15674 , n23406 , n20962 );
    xnor g3378 ( n23559 , n19601 , n10800 );
    nor g3379 ( n7967 , n8526 , n12232 );
    xnor g3380 ( n6121 , n17183 , n20036 );
    and g3381 ( n12338 , n12085 , n9277 );
    nor g3382 ( n9661 , n11924 , n10986 );
    and g3383 ( n13705 , n24769 , n25401 );
    or g3384 ( n25388 , n24008 , n5 );
    xnor g3385 ( n331 , n1045 , n1603 );
    nor g3386 ( n26678 , n658 , n21095 );
    or g3387 ( n4587 , n22631 , n1167 );
    and g3388 ( n18706 , n3567 , n8137 );
    and g3389 ( n3464 , n5355 , n5000 );
    or g3390 ( n15571 , n5140 , n20796 );
    xnor g3391 ( n26934 , n7102 , n12249 );
    or g3392 ( n20866 , n18485 , n19228 );
    xnor g3393 ( n565 , n22379 , n767 );
    xnor g3394 ( n2488 , n19989 , n18639 );
    and g3395 ( n5481 , n18808 , n1874 );
    xnor g3396 ( n19120 , n15696 , n23545 );
    nor g3397 ( n17710 , n21539 , n6200 );
    or g3398 ( n9895 , n13855 , n1246 );
    or g3399 ( n15554 , n25041 , n16205 );
    or g3400 ( n5188 , n18573 , n15830 );
    or g3401 ( n18368 , n21386 , n21287 );
    or g3402 ( n3227 , n9039 , n12286 );
    nor g3403 ( n3092 , n17940 , n111 );
    xnor g3404 ( n14190 , n9224 , n21449 );
    xnor g3405 ( n1629 , n7413 , n15285 );
    or g3406 ( n1456 , n11302 , n19876 );
    and g3407 ( n11862 , n23709 , n14268 );
    or g3408 ( n3442 , n11370 , n3837 );
    or g3409 ( n6906 , n13584 , n1830 );
    xnor g3410 ( n3588 , n15892 , n3739 );
    and g3411 ( n20549 , n27086 , n5504 );
    xnor g3412 ( n17526 , n4435 , n8533 );
    nor g3413 ( n16236 , n19540 , n25637 );
    xnor g3414 ( n4613 , n13214 , n19144 );
    nor g3415 ( n16017 , n9713 , n1471 );
    xnor g3416 ( n398 , n10117 , n23250 );
    and g3417 ( n16410 , n4884 , n8091 );
    xnor g3418 ( n3603 , n12061 , n1887 );
    or g3419 ( n7618 , n14293 , n20409 );
    and g3420 ( n18936 , n15294 , n15270 );
    or g3421 ( n12786 , n25527 , n16171 );
    or g3422 ( n23137 , n14569 , n20658 );
    not g3423 ( n23634 , n25504 );
    xnor g3424 ( n18531 , n2409 , n14071 );
    and g3425 ( n16006 , n5965 , n9200 );
    not g3426 ( n472 , n4858 );
    nor g3427 ( n22675 , n9655 , n20946 );
    nor g3428 ( n16717 , n24048 , n19683 );
    xnor g3429 ( n19569 , n1199 , n11698 );
    nor g3430 ( n9818 , n20359 , n23704 );
    not g3431 ( n1584 , n10949 );
    and g3432 ( n367 , n25914 , n198 );
    xnor g3433 ( n11261 , n18796 , n2667 );
    not g3434 ( n7343 , n16794 );
    xnor g3435 ( n24274 , n18880 , n2978 );
    xnor g3436 ( n3355 , n22247 , n21126 );
    or g3437 ( n21091 , n2252 , n22020 );
    or g3438 ( n14690 , n6218 , n7669 );
    or g3439 ( n1678 , n24367 , n15991 );
    or g3440 ( n3493 , n16267 , n4299 );
    nor g3441 ( n12363 , n3967 , n8338 );
    not g3442 ( n24131 , n21848 );
    and g3443 ( n18868 , n5672 , n21086 );
    xnor g3444 ( n5587 , n17587 , n25958 );
    or g3445 ( n25535 , n12272 , n16709 );
    not g3446 ( n14856 , n22274 );
    xnor g3447 ( n7703 , n6727 , n5182 );
    not g3448 ( n14094 , n25781 );
    xnor g3449 ( n18583 , n6409 , n4477 );
    and g3450 ( n25352 , n19634 , n27184 );
    and g3451 ( n26482 , n13944 , n23871 );
    not g3452 ( n6724 , n19161 );
    or g3453 ( n11065 , n13689 , n19004 );
    xnor g3454 ( n16117 , n2089 , n25094 );
    xor g3455 ( n21914 , n13976 , n10250 );
    not g3456 ( n19157 , n15077 );
    or g3457 ( n26948 , n25269 , n23641 );
    not g3458 ( n22659 , n13150 );
    not g3459 ( n9615 , n25924 );
    not g3460 ( n18008 , n26167 );
    xnor g3461 ( n26334 , n9061 , n314 );
    or g3462 ( n8611 , n7893 , n19701 );
    and g3463 ( n15862 , n21023 , n19537 );
    and g3464 ( n8808 , n6347 , n10589 );
    and g3465 ( n754 , n13662 , n7589 );
    nor g3466 ( n10119 , n12673 , n25220 );
    or g3467 ( n21535 , n15411 , n1079 );
    or g3468 ( n9472 , n6912 , n18488 );
    or g3469 ( n20635 , n19662 , n5930 );
    xnor g3470 ( n5409 , n5329 , n1 );
    or g3471 ( n13816 , n22631 , n21078 );
    and g3472 ( n23113 , n4137 , n7789 );
    xnor g3473 ( n9593 , n726 , n25749 );
    nor g3474 ( n1108 , n3770 , n24801 );
    xnor g3475 ( n19372 , n12289 , n12892 );
    xnor g3476 ( n22569 , n25228 , n5337 );
    or g3477 ( n19029 , n27043 , n27170 );
    nor g3478 ( n18121 , n6919 , n1755 );
    or g3479 ( n15782 , n22290 , n12878 );
    and g3480 ( n9122 , n8698 , n22788 );
    xnor g3481 ( n8510 , n12190 , n21368 );
    xnor g3482 ( n21679 , n2191 , n26053 );
    or g3483 ( n22096 , n25707 , n10510 );
    xnor g3484 ( n15739 , n24495 , n22764 );
    xnor g3485 ( n5243 , n6399 , n14738 );
    not g3486 ( n23814 , n22625 );
    or g3487 ( n16545 , n6313 , n25529 );
    xnor g3488 ( n11285 , n4512 , n24201 );
    xnor g3489 ( n10785 , n11729 , n10718 );
    xnor g3490 ( n11936 , n9250 , n885 );
    xnor g3491 ( n1993 , n5213 , n4812 );
    nor g3492 ( n8235 , n9627 , n8712 );
    nor g3493 ( n14995 , n25021 , n11841 );
    xnor g3494 ( n12461 , n14820 , n6257 );
    or g3495 ( n17719 , n19511 , n8857 );
    and g3496 ( n25991 , n8316 , n18284 );
    and g3497 ( n16939 , n7640 , n3509 );
    nor g3498 ( n5989 , n2565 , n25490 );
    and g3499 ( n10471 , n2226 , n17146 );
    xnor g3500 ( n23691 , n8661 , n24786 );
    xnor g3501 ( n7134 , n22296 , n4936 );
    xnor g3502 ( n13573 , n10017 , n20349 );
    and g3503 ( n25253 , n5534 , n19693 );
    xnor g3504 ( n2619 , n10149 , n12047 );
    nor g3505 ( n122 , n8964 , n11764 );
    and g3506 ( n3572 , n4565 , n2600 );
    xnor g3507 ( n21858 , n14808 , n25358 );
    and g3508 ( n5586 , n710 , n8398 );
    not g3509 ( n17141 , n9440 );
    xnor g3510 ( n4826 , n25475 , n23697 );
    not g3511 ( n7254 , n5752 );
    not g3512 ( n20939 , n18358 );
    or g3513 ( n20189 , n5302 , n19484 );
    or g3514 ( n20370 , n4957 , n22688 );
    nor g3515 ( n12024 , n6814 , n10763 );
    or g3516 ( n10293 , n24572 , n95 );
    and g3517 ( n19415 , n15916 , n392 );
    and g3518 ( n11990 , n15466 , n3969 );
    or g3519 ( n15187 , n24134 , n8164 );
    xnor g3520 ( n21586 , n12018 , n19453 );
    and g3521 ( n10435 , n8513 , n10709 );
    not g3522 ( n21442 , n21458 );
    or g3523 ( n21808 , n13924 , n22449 );
    or g3524 ( n7241 , n11100 , n22513 );
    or g3525 ( n2558 , n7208 , n23968 );
    not g3526 ( n26768 , n13667 );
    not g3527 ( n16594 , n16507 );
    and g3528 ( n25593 , n3251 , n3530 );
    not g3529 ( n3764 , n4294 );
    or g3530 ( n19275 , n1075 , n137 );
    xnor g3531 ( n11207 , n7657 , n25926 );
    or g3532 ( n1633 , n11855 , n25366 );
    xnor g3533 ( n22596 , n4562 , n3136 );
    xnor g3534 ( n12487 , n8451 , n4537 );
    or g3535 ( n2400 , n2722 , n9390 );
    and g3536 ( n18280 , n20056 , n17692 );
    xnor g3537 ( n6714 , n18319 , n6267 );
    or g3538 ( n14221 , n15553 , n16883 );
    or g3539 ( n11492 , n11177 , n13137 );
    and g3540 ( n11722 , n9386 , n17691 );
    or g3541 ( n1165 , n7082 , n23466 );
    not g3542 ( n4003 , n25221 );
    xnor g3543 ( n17338 , n20862 , n6876 );
    xnor g3544 ( n23714 , n20900 , n9350 );
    or g3545 ( n10600 , n11081 , n12023 );
    or g3546 ( n20380 , n12387 , n6057 );
    or g3547 ( n11912 , n19584 , n6279 );
    not g3548 ( n7970 , n26705 );
    and g3549 ( n12466 , n11530 , n11545 );
    or g3550 ( n10149 , n21635 , n13295 );
    not g3551 ( n17864 , n3187 );
    and g3552 ( n6505 , n11780 , n12254 );
    xnor g3553 ( n26104 , n23907 , n25731 );
    or g3554 ( n17473 , n18814 , n9037 );
    not g3555 ( n5240 , n19665 );
    nor g3556 ( n8987 , n21984 , n4440 );
    or g3557 ( n12005 , n6426 , n2362 );
    or g3558 ( n1295 , n26543 , n26244 );
    not g3559 ( n3354 , n21175 );
    nor g3560 ( n5836 , n21066 , n23789 );
    not g3561 ( n22958 , n26797 );
    and g3562 ( n23626 , n18096 , n14377 );
    and g3563 ( n9651 , n18855 , n20925 );
    nor g3564 ( n6564 , n4338 , n24430 );
    or g3565 ( n6827 , n437 , n26945 );
    nor g3566 ( n7571 , n6038 , n12171 );
    or g3567 ( n16292 , n18952 , n16966 );
    and g3568 ( n11004 , n604 , n4626 );
    xnor g3569 ( n26810 , n2503 , n20929 );
    xnor g3570 ( n2214 , n16076 , n13660 );
    nor g3571 ( n3033 , n5260 , n16130 );
    xnor g3572 ( n19379 , n16274 , n23849 );
    not g3573 ( n19254 , n485 );
    and g3574 ( n8791 , n2955 , n6191 );
    or g3575 ( n23889 , n7842 , n23989 );
    or g3576 ( n8500 , n22442 , n3131 );
    or g3577 ( n25745 , n14695 , n847 );
    nor g3578 ( n12096 , n1497 , n4184 );
    xnor g3579 ( n1420 , n7143 , n3625 );
    and g3580 ( n10460 , n24248 , n10640 );
    nor g3581 ( n3731 , n27068 , n8508 );
    or g3582 ( n18493 , n26564 , n7471 );
    and g3583 ( n518 , n6860 , n10539 );
    and g3584 ( n18001 , n2011 , n18845 );
    not g3585 ( n26170 , n5750 );
    xnor g3586 ( n27096 , n17309 , n1909 );
    or g3587 ( n20561 , n3831 , n21366 );
    and g3588 ( n4751 , n19999 , n26561 );
    nor g3589 ( n11753 , n2815 , n10455 );
    or g3590 ( n3309 , n401 , n17410 );
    or g3591 ( n13762 , n6039 , n9394 );
    xnor g3592 ( n6944 , n8876 , n4975 );
    not g3593 ( n4033 , n19108 );
    and g3594 ( n21681 , n12947 , n24449 );
    xnor g3595 ( n22884 , n4775 , n20235 );
    nor g3596 ( n24083 , n13357 , n506 );
    or g3597 ( n22579 , n9600 , n19701 );
    and g3598 ( n15044 , n20555 , n17246 );
    xnor g3599 ( n5085 , n5696 , n23463 );
    or g3600 ( n12365 , n24486 , n7092 );
    and g3601 ( n21542 , n4169 , n25300 );
    xnor g3602 ( n16887 , n22862 , n16543 );
    or g3603 ( n22417 , n13731 , n21038 );
    not g3604 ( n3853 , n12265 );
    or g3605 ( n9630 , n18018 , n1337 );
    not g3606 ( n11649 , n26726 );
    and g3607 ( n84 , n22486 , n14266 );
    or g3608 ( n17148 , n17951 , n14084 );
    or g3609 ( n19671 , n5779 , n2103 );
    xnor g3610 ( n23337 , n19610 , n9159 );
    or g3611 ( n24440 , n10066 , n18565 );
    nor g3612 ( n4285 , n25797 , n10611 );
    or g3613 ( n18650 , n6092 , n26261 );
    or g3614 ( n10824 , n6247 , n11867 );
    or g3615 ( n12867 , n11826 , n7205 );
    or g3616 ( n6722 , n16389 , n13700 );
    xnor g3617 ( n6178 , n2430 , n16550 );
    or g3618 ( n17619 , n21486 , n12338 );
    and g3619 ( n4981 , n18637 , n9916 );
    or g3620 ( n7413 , n4728 , n969 );
    xnor g3621 ( n11592 , n10806 , n21160 );
    and g3622 ( n16501 , n17904 , n683 );
    not g3623 ( n14293 , n1099 );
    xnor g3624 ( n4934 , n7876 , n25435 );
    not g3625 ( n26505 , n3700 );
    nor g3626 ( n8775 , n9469 , n3237 );
    and g3627 ( n2066 , n24850 , n22706 );
    and g3628 ( n17985 , n3626 , n21099 );
    nor g3629 ( n23330 , n11121 , n19494 );
    or g3630 ( n19586 , n21867 , n19155 );
    or g3631 ( n4135 , n3948 , n4551 );
    not g3632 ( n22428 , n18416 );
    nor g3633 ( n21708 , n21556 , n23068 );
    or g3634 ( n25108 , n12576 , n17287 );
    and g3635 ( n24385 , n1522 , n14138 );
    or g3636 ( n7736 , n25778 , n7223 );
    or g3637 ( n3024 , n16654 , n7824 );
    not g3638 ( n19856 , n6458 );
    nor g3639 ( n970 , n3069 , n18485 );
    xnor g3640 ( n15489 , n578 , n24622 );
    nor g3641 ( n12795 , n24327 , n25967 );
    and g3642 ( n14727 , n24362 , n10007 );
    not g3643 ( n23620 , n26853 );
    xnor g3644 ( n4382 , n5360 , n10493 );
    xnor g3645 ( n21733 , n24763 , n18089 );
    or g3646 ( n3467 , n27182 , n9033 );
    and g3647 ( n100 , n9107 , n18008 );
    or g3648 ( n3295 , n6488 , n10521 );
    xnor g3649 ( n22818 , n18318 , n3946 );
    xnor g3650 ( n9409 , n19368 , n24828 );
    or g3651 ( n7067 , n24432 , n14327 );
    and g3652 ( n5785 , n6299 , n7096 );
    not g3653 ( n15487 , n11036 );
    xnor g3654 ( n25871 , n13839 , n2575 );
    or g3655 ( n22947 , n24614 , n5830 );
    nor g3656 ( n15682 , n5580 , n3359 );
    nor g3657 ( n18761 , n24990 , n19502 );
    not g3658 ( n2818 , n24796 );
    xnor g3659 ( n7351 , n26865 , n15839 );
    or g3660 ( n474 , n7000 , n19535 );
    or g3661 ( n21872 , n14496 , n14552 );
    not g3662 ( n6366 , n14184 );
    and g3663 ( n25307 , n17641 , n8336 );
    not g3664 ( n22260 , n5387 );
    or g3665 ( n7696 , n24062 , n4911 );
    and g3666 ( n26955 , n6231 , n13107 );
    not g3667 ( n311 , n13465 );
    xnor g3668 ( n3281 , n5743 , n17967 );
    nor g3669 ( n1096 , n9873 , n20558 );
    xnor g3670 ( n674 , n6698 , n21295 );
    and g3671 ( n3706 , n7974 , n2759 );
    and g3672 ( n20627 , n14483 , n18747 );
    nor g3673 ( n14683 , n19460 , n12586 );
    nor g3674 ( n21141 , n8322 , n3468 );
    or g3675 ( n13150 , n26744 , n16240 );
    not g3676 ( n22123 , n18578 );
    not g3677 ( n16486 , n26619 );
    and g3678 ( n19259 , n13701 , n14270 );
    xnor g3679 ( n8022 , n11657 , n12426 );
    or g3680 ( n7126 , n21016 , n19254 );
    not g3681 ( n22550 , n11605 );
    or g3682 ( n14742 , n8396 , n12539 );
    nor g3683 ( n73 , n18451 , n27034 );
    or g3684 ( n25420 , n22261 , n20094 );
    or g3685 ( n24224 , n22418 , n23443 );
    and g3686 ( n87 , n4757 , n3598 );
    or g3687 ( n3188 , n9701 , n6076 );
    and g3688 ( n22087 , n26093 , n10529 );
    not g3689 ( n13842 , n23775 );
    xnor g3690 ( n18806 , n8197 , n1927 );
    and g3691 ( n17307 , n12899 , n3534 );
    or g3692 ( n19753 , n3620 , n14753 );
    xnor g3693 ( n24788 , n19942 , n11387 );
    xnor g3694 ( n23597 , n654 , n13932 );
    and g3695 ( n23599 , n13180 , n10103 );
    not g3696 ( n4338 , n20980 );
    or g3697 ( n12722 , n21066 , n11497 );
    xnor g3698 ( n6956 , n6899 , n1883 );
    not g3699 ( n17605 , n25355 );
    or g3700 ( n4809 , n874 , n9043 );
    xnor g3701 ( n20822 , n25110 , n2570 );
    or g3702 ( n13545 , n1559 , n4348 );
    not g3703 ( n10112 , n5954 );
    xnor g3704 ( n933 , n17943 , n4306 );
    xnor g3705 ( n5228 , n9312 , n3336 );
    nor g3706 ( n8218 , n26344 , n1433 );
    not g3707 ( n1672 , n5206 );
    or g3708 ( n10393 , n6221 , n14287 );
    or g3709 ( n8618 , n5223 , n23136 );
    xnor g3710 ( n12353 , n15146 , n10125 );
    nor g3711 ( n13540 , n3256 , n16300 );
    nor g3712 ( n21631 , n23591 , n24690 );
    not g3713 ( n24690 , n20624 );
    xnor g3714 ( n13336 , n1143 , n12817 );
    xnor g3715 ( n15908 , n18452 , n6397 );
    xnor g3716 ( n26630 , n24202 , n9595 );
    not g3717 ( n7326 , n22355 );
    nor g3718 ( n9039 , n3319 , n10255 );
    or g3719 ( n582 , n15865 , n3415 );
    xnor g3720 ( n23165 , n14391 , n6293 );
    xnor g3721 ( n3445 , n6077 , n24767 );
    xnor g3722 ( n5597 , n5722 , n402 );
    not g3723 ( n3724 , n12319 );
    not g3724 ( n18070 , n8302 );
    and g3725 ( n21744 , n1654 , n24245 );
    xnor g3726 ( n24265 , n12208 , n12522 );
    xnor g3727 ( n22727 , n3680 , n2697 );
    or g3728 ( n871 , n24116 , n19797 );
    or g3729 ( n8211 , n24545 , n26364 );
    or g3730 ( n4875 , n649 , n16374 );
    xnor g3731 ( n3955 , n14349 , n19142 );
    or g3732 ( n5173 , n10307 , n23633 );
    not g3733 ( n12474 , n3984 );
    and g3734 ( n8788 , n23444 , n15561 );
    nor g3735 ( n25759 , n21634 , n7930 );
    xnor g3736 ( n25178 , n3031 , n8017 );
    not g3737 ( n678 , n25413 );
    xnor g3738 ( n9752 , n22043 , n12121 );
    or g3739 ( n20892 , n24471 , n5209 );
    xnor g3740 ( n21765 , n5937 , n18719 );
    or g3741 ( n9804 , n12714 , n18584 );
    xnor g3742 ( n3871 , n6040 , n26280 );
    or g3743 ( n16231 , n14569 , n26661 );
    and g3744 ( n20164 , n8829 , n4452 );
    xnor g3745 ( n26131 , n5974 , n19313 );
    or g3746 ( n20778 , n25314 , n19335 );
    xnor g3747 ( n18142 , n7083 , n18037 );
    not g3748 ( n15860 , n10351 );
    xnor g3749 ( n6367 , n4288 , n24646 );
    and g3750 ( n1601 , n4759 , n4818 );
    nor g3751 ( n18240 , n3311 , n1139 );
    and g3752 ( n7269 , n20134 , n15237 );
    or g3753 ( n10572 , n21826 , n17670 );
    or g3754 ( n12820 , n20383 , n3341 );
    and g3755 ( n4672 , n12312 , n16107 );
    nor g3756 ( n6117 , n1956 , n16594 );
    xnor g3757 ( n12034 , n16672 , n2252 );
    and g3758 ( n15542 , n5767 , n23435 );
    not g3759 ( n21984 , n16906 );
    not g3760 ( n7644 , n10352 );
    not g3761 ( n9525 , n4639 );
    not g3762 ( n18710 , n26007 );
    buf g3763 ( n11321 , n19499 );
    and g3764 ( n12255 , n12069 , n16115 );
    and g3765 ( n23941 , n3273 , n20414 );
    and g3766 ( n26209 , n4371 , n11849 );
    and g3767 ( n6313 , n24072 , n14312 );
    and g3768 ( n13872 , n13081 , n18451 );
    and g3769 ( n22840 , n5326 , n15669 );
    nor g3770 ( n6855 , n8851 , n9944 );
    xnor g3771 ( n2249 , n22693 , n19722 );
    and g3772 ( n24692 , n21933 , n668 );
    not g3773 ( n16560 , n10377 );
    or g3774 ( n6493 , n4807 , n5059 );
    or g3775 ( n4630 , n12650 , n18486 );
    nor g3776 ( n26019 , n23589 , n12891 );
    nor g3777 ( n20975 , n21613 , n6242 );
    nor g3778 ( n13469 , n45 , n15657 );
    xnor g3779 ( n11002 , n42 , n5348 );
    and g3780 ( n4494 , n21242 , n6167 );
    xnor g3781 ( n11297 , n23161 , n3383 );
    xnor g3782 ( n6961 , n16158 , n24085 );
    xnor g3783 ( n4963 , n24293 , n12765 );
    xnor g3784 ( n18201 , n5571 , n9672 );
    nor g3785 ( n4544 , n20213 , n9765 );
    and g3786 ( n5692 , n22281 , n8537 );
    or g3787 ( n19837 , n22420 , n15862 );
    not g3788 ( n22021 , n18812 );
    or g3789 ( n12653 , n27039 , n18656 );
    xnor g3790 ( n23303 , n22176 , n12384 );
    xnor g3791 ( n197 , n24635 , n11800 );
    or g3792 ( n3364 , n23895 , n4446 );
    not g3793 ( n21420 , n18934 );
    xnor g3794 ( n15586 , n12828 , n3602 );
    xnor g3795 ( n7432 , n18984 , n5856 );
    xnor g3796 ( n10204 , n19113 , n2731 );
    xnor g3797 ( n21365 , n16005 , n17081 );
    and g3798 ( n3654 , n3255 , n18169 );
    not g3799 ( n23506 , n4978 );
    or g3800 ( n13312 , n4868 , n10993 );
    or g3801 ( n19138 , n22924 , n15745 );
    and g3802 ( n3441 , n11652 , n5047 );
    xnor g3803 ( n9860 , n22049 , n24196 );
    xnor g3804 ( n19938 , n14932 , n17623 );
    xnor g3805 ( n12302 , n18670 , n135 );
    and g3806 ( n25581 , n2906 , n14187 );
    xnor g3807 ( n26573 , n7128 , n24030 );
    nor g3808 ( n25172 , n25007 , n24286 );
    nor g3809 ( n377 , n11172 , n7325 );
    or g3810 ( n10497 , n10650 , n17978 );
    nor g3811 ( n9681 , n8186 , n20040 );
    or g3812 ( n16756 , n13637 , n2622 );
    and g3813 ( n20957 , n4155 , n13031 );
    or g3814 ( n21552 , n21621 , n813 );
    xnor g3815 ( n27170 , n15084 , n16615 );
    nor g3816 ( n18521 , n17641 , n12198 );
    or g3817 ( n23595 , n7306 , n8374 );
    or g3818 ( n8213 , n11583 , n20544 );
    xnor g3819 ( n20748 , n4950 , n97 );
    not g3820 ( n2121 , n19454 );
    or g3821 ( n22348 , n21599 , n26324 );
    and g3822 ( n22833 , n10886 , n9542 );
    and g3823 ( n8298 , n6857 , n14400 );
    xnor g3824 ( n12783 , n2911 , n9072 );
    xnor g3825 ( n14975 , n25120 , n3582 );
    or g3826 ( n4233 , n7224 , n26663 );
    xnor g3827 ( n19920 , n20455 , n3828 );
    nor g3828 ( n5578 , n1558 , n3918 );
    xnor g3829 ( n25079 , n6218 , n25464 );
    xnor g3830 ( n27060 , n866 , n17155 );
    xnor g3831 ( n22080 , n3839 , n21774 );
    nor g3832 ( n26088 , n17381 , n13649 );
    not g3833 ( n10266 , n14524 );
    or g3834 ( n2294 , n3290 , n5873 );
    and g3835 ( n14261 , n8543 , n12028 );
    and g3836 ( n6234 , n10761 , n3985 );
    and g3837 ( n15392 , n8147 , n9650 );
    and g3838 ( n3761 , n11141 , n9189 );
    or g3839 ( n21494 , n22760 , n7576 );
    xnor g3840 ( n23673 , n10767 , n15062 );
    nor g3841 ( n2236 , n13443 , n23923 );
    or g3842 ( n15804 , n6136 , n10708 );
    not g3843 ( n11409 , n15670 );
    xnor g3844 ( n8889 , n13468 , n3705 );
    xnor g3845 ( n8731 , n15693 , n3391 );
    and g3846 ( n3358 , n18029 , n16779 );
    xnor g3847 ( n26674 , n26038 , n5522 );
    and g3848 ( n24294 , n8284 , n25361 );
    or g3849 ( n24687 , n4295 , n11151 );
    or g3850 ( n20585 , n153 , n26301 );
    and g3851 ( n6538 , n21592 , n14709 );
    xnor g3852 ( n16290 , n18885 , n2116 );
    and g3853 ( n7737 , n21578 , n1295 );
    and g3854 ( n7208 , n16722 , n21101 );
    and g3855 ( n25755 , n15117 , n13716 );
    or g3856 ( n10880 , n11402 , n7854 );
    or g3857 ( n27045 , n10443 , n25537 );
    xnor g3858 ( n21032 , n13098 , n3056 );
    nor g3859 ( n6215 , n16449 , n4185 );
    not g3860 ( n6753 , n18290 );
    xnor g3861 ( n15642 , n21508 , n19393 );
    nor g3862 ( n15928 , n11938 , n25126 );
    nor g3863 ( n16101 , n6138 , n3317 );
    and g3864 ( n5358 , n11046 , n18890 );
    and g3865 ( n12533 , n19234 , n1365 );
    xnor g3866 ( n16251 , n2044 , n7130 );
    xnor g3867 ( n25210 , n22913 , n441 );
    or g3868 ( n22128 , n13731 , n8920 );
    xnor g3869 ( n1147 , n10405 , n7731 );
    xnor g3870 ( n19114 , n23862 , n14538 );
    nor g3871 ( n8423 , n20075 , n18158 );
    xnor g3872 ( n11882 , n2979 , n9554 );
    or g3873 ( n17080 , n10740 , n17564 );
    or g3874 ( n25822 , n12576 , n25475 );
    xnor g3875 ( n1580 , n5294 , n17279 );
    and g3876 ( n16390 , n5808 , n7696 );
    or g3877 ( n17875 , n25101 , n15174 );
    and g3878 ( n18153 , n15673 , n21003 );
    xnor g3879 ( n9503 , n643 , n17804 );
    xnor g3880 ( n20162 , n24705 , n26444 );
    or g3881 ( n19961 , n932 , n10739 );
    and g3882 ( n6545 , n23092 , n22228 );
    xnor g3883 ( n19337 , n7925 , n15926 );
    xnor g3884 ( n8178 , n26495 , n19701 );
    or g3885 ( n20858 , n23957 , n3825 );
    and g3886 ( n7687 , n21921 , n14214 );
    xnor g3887 ( n21308 , n12351 , n6503 );
    xnor g3888 ( n16794 , n21662 , n6773 );
    or g3889 ( n8634 , n18333 , n12509 );
    xnor g3890 ( n26584 , n4377 , n18961 );
    xnor g3891 ( n4010 , n19755 , n6367 );
    and g3892 ( n26092 , n16524 , n17539 );
    xnor g3893 ( n3017 , n4600 , n9981 );
    xnor g3894 ( n21824 , n17127 , n17731 );
    xnor g3895 ( n12288 , n5951 , n17383 );
    xnor g3896 ( n21620 , n24448 , n9534 );
    not g3897 ( n23932 , n8656 );
    or g3898 ( n1130 , n23296 , n5413 );
    and g3899 ( n25851 , n13358 , n25453 );
    nor g3900 ( n27052 , n4692 , n21469 );
    xnor g3901 ( n4273 , n14620 , n17077 );
    or g3902 ( n20085 , n12821 , n6596 );
    not g3903 ( n24970 , n6699 );
    xnor g3904 ( n23663 , n1033 , n8619 );
    nor g3905 ( n22983 , n21138 , n3187 );
    not g3906 ( n10581 , n1700 );
    or g3907 ( n17111 , n20165 , n5721 );
    not g3908 ( n20829 , n1738 );
    xnor g3909 ( n4954 , n26553 , n23775 );
    and g3910 ( n6377 , n10181 , n2066 );
    not g3911 ( n12906 , n4108 );
    xnor g3912 ( n7935 , n1874 , n1313 );
    not g3913 ( n14564 , n21492 );
    xnor g3914 ( n22831 , n5354 , n14972 );
    and g3915 ( n19408 , n7564 , n10952 );
    or g3916 ( n6417 , n23063 , n15265 );
    or g3917 ( n16197 , n1816 , n19013 );
    xnor g3918 ( n9917 , n1758 , n10878 );
    or g3919 ( n3579 , n14002 , n16396 );
    not g3920 ( n26486 , n12531 );
    and g3921 ( n17460 , n18663 , n11820 );
    xnor g3922 ( n10022 , n19729 , n10745 );
    xnor g3923 ( n16640 , n6955 , n22457 );
    xnor g3924 ( n10772 , n15086 , n17971 );
    nor g3925 ( n8362 , n23884 , n17289 );
    and g3926 ( n5499 , n22727 , n17411 );
    or g3927 ( n774 , n16582 , n17808 );
    or g3928 ( n16335 , n16983 , n14411 );
    xnor g3929 ( n21545 , n18203 , n16366 );
    or g3930 ( n7878 , n2916 , n24559 );
    and g3931 ( n17824 , n808 , n12102 );
    and g3932 ( n23291 , n22231 , n24640 );
    or g3933 ( n23344 , n13502 , n11224 );
    not g3934 ( n8462 , n26763 );
    xnor g3935 ( n25406 , n20478 , n1204 );
    xnor g3936 ( n6700 , n17640 , n13217 );
    not g3937 ( n11098 , n9653 );
    or g3938 ( n6730 , n11405 , n18305 );
    not g3939 ( n1739 , n17525 );
    or g3940 ( n7135 , n24836 , n10329 );
    and g3941 ( n6005 , n23278 , n7493 );
    buf g3942 ( n21247 , n5178 );
    xnor g3943 ( n23259 , n2421 , n5337 );
    and g3944 ( n7576 , n2138 , n5035 );
    xnor g3945 ( n25999 , n15229 , n8050 );
    or g3946 ( n16385 , n19701 , n13074 );
    nor g3947 ( n9049 , n21608 , n7721 );
    or g3948 ( n13744 , n13102 , n14199 );
    not g3949 ( n27027 , n16285 );
    xnor g3950 ( n14830 , n10688 , n1169 );
    xnor g3951 ( n8480 , n4684 , n2471 );
    or g3952 ( n27119 , n22585 , n23226 );
    or g3953 ( n26879 , n19911 , n10472 );
    xnor g3954 ( n24373 , n26357 , n7976 );
    or g3955 ( n25911 , n10102 , n12661 );
    or g3956 ( n21677 , n11166 , n5358 );
    xnor g3957 ( n7616 , n1508 , n13928 );
    xnor g3958 ( n10949 , n18220 , n20634 );
    xnor g3959 ( n15355 , n16260 , n26804 );
    or g3960 ( n7380 , n19371 , n15960 );
    xnor g3961 ( n13215 , n13953 , n18950 );
    xnor g3962 ( n19590 , n16477 , n11697 );
    and g3963 ( n23524 , n9836 , n16676 );
    and g3964 ( n9588 , n20489 , n26913 );
    not g3965 ( n19594 , n8422 );
    not g3966 ( n24212 , n21112 );
    not g3967 ( n6401 , n18703 );
    xnor g3968 ( n27015 , n8141 , n18094 );
    and g3969 ( n17076 , n14246 , n13272 );
    xnor g3970 ( n8119 , n22560 , n23575 );
    xnor g3971 ( n27102 , n3182 , n21854 );
    or g3972 ( n27053 , n24358 , n24665 );
    and g3973 ( n20055 , n11651 , n12906 );
    or g3974 ( n17509 , n7330 , n2479 );
    nor g3975 ( n6086 , n88 , n14453 );
    or g3976 ( n18086 , n17479 , n12821 );
    nor g3977 ( n22925 , n15189 , n1364 );
    or g3978 ( n1217 , n2350 , n19487 );
    and g3979 ( n9718 , n2915 , n10224 );
    xnor g3980 ( n22634 , n6045 , n16690 );
    or g3981 ( n2905 , n24478 , n1623 );
    nor g3982 ( n14601 , n17664 , n5115 );
    xnor g3983 ( n12813 , n22332 , n21934 );
    xnor g3984 ( n24795 , n15258 , n11775 );
    or g3985 ( n4219 , n6932 , n5973 );
    xnor g3986 ( n8027 , n16000 , n16692 );
    and g3987 ( n7874 , n3105 , n27097 );
    or g3988 ( n24676 , n27046 , n14282 );
    or g3989 ( n11212 , n7935 , n18608 );
    not g3990 ( n9565 , n13258 );
    and g3991 ( n21187 , n9380 , n24686 );
    xnor g3992 ( n4478 , n3462 , n7703 );
    xnor g3993 ( n7395 , n7466 , n21721 );
    or g3994 ( n18980 , n8672 , n5296 );
    or g3995 ( n11852 , n26654 , n9538 );
    not g3996 ( n16586 , n9250 );
    xnor g3997 ( n18982 , n1094 , n10644 );
    not g3998 ( n15580 , n17251 );
    nor g3999 ( n12410 , n8721 , n1040 );
    nor g4000 ( n17226 , n15910 , n8609 );
    and g4001 ( n13916 , n10544 , n6163 );
    nor g4002 ( n14104 , n1163 , n18901 );
    or g4003 ( n2123 , n8208 , n18718 );
    and g4004 ( n13341 , n14798 , n10162 );
    not g4005 ( n10398 , n23212 );
    or g4006 ( n4054 , n23514 , n15132 );
    xnor g4007 ( n21673 , n12734 , n20023 );
    or g4008 ( n13512 , n14284 , n4276 );
    or g4009 ( n10809 , n8542 , n7029 );
    not g4010 ( n8991 , n10633 );
    not g4011 ( n5475 , n22404 );
    and g4012 ( n1258 , n2688 , n8163 );
    or g4013 ( n16997 , n10416 , n5107 );
    nor g4014 ( n6898 , n18472 , n20745 );
    xnor g4015 ( n25765 , n21606 , n26786 );
    and g4016 ( n231 , n10083 , n7762 );
    xnor g4017 ( n10041 , n14513 , n12063 );
    or g4018 ( n18281 , n24978 , n17278 );
    or g4019 ( n21933 , n2903 , n25120 );
    and g4020 ( n18833 , n26310 , n14799 );
    or g4021 ( n26490 , n26470 , n21654 );
    nor g4022 ( n7714 , n17101 , n552 );
    nor g4023 ( n25298 , n24074 , n23464 );
    xnor g4024 ( n17692 , n12017 , n8169 );
    and g4025 ( n578 , n19405 , n15115 );
    xnor g4026 ( n10306 , n9028 , n25240 );
    xnor g4027 ( n5265 , n4034 , n3291 );
    xnor g4028 ( n8302 , n24831 , n4349 );
    not g4029 ( n20948 , n3786 );
    xnor g4030 ( n24372 , n17408 , n20235 );
    or g4031 ( n9927 , n14692 , n9387 );
    and g4032 ( n23886 , n15992 , n6093 );
    xnor g4033 ( n7457 , n19207 , n12424 );
    and g4034 ( n18111 , n16633 , n9923 );
    and g4035 ( n5662 , n4778 , n1787 );
    and g4036 ( n16855 , n3449 , n22195 );
    xnor g4037 ( n9358 , n21692 , n24812 );
    or g4038 ( n25750 , n7712 , n13972 );
    xnor g4039 ( n10427 , n13976 , n16903 );
    xnor g4040 ( n4134 , n9116 , n10466 );
    or g4041 ( n8811 , n22244 , n12834 );
    nor g4042 ( n14149 , n8001 , n20516 );
    and g4043 ( n22292 , n2835 , n26262 );
    xnor g4044 ( n10447 , n3280 , n8117 );
    nor g4045 ( n16222 , n19816 , n9421 );
    buf g4046 ( n13359 , n17180 );
    or g4047 ( n23569 , n15513 , n6690 );
    or g4048 ( n6696 , n24718 , n22677 );
    and g4049 ( n25978 , n26198 , n2982 );
    nor g4050 ( n20924 , n18496 , n25331 );
    or g4051 ( n1315 , n759 , n22848 );
    nor g4052 ( n1870 , n11363 , n6590 );
    or g4053 ( n20246 , n17305 , n7817 );
    or g4054 ( n3070 , n22814 , n26355 );
    nor g4055 ( n1161 , n3837 , n12184 );
    not g4056 ( n2633 , n23432 );
    xnor g4057 ( n1519 , n19235 , n6799 );
    or g4058 ( n16408 , n20581 , n24109 );
    xnor g4059 ( n2583 , n12946 , n21067 );
    xnor g4060 ( n1735 , n20507 , n25086 );
    xnor g4061 ( n22376 , n644 , n12868 );
    and g4062 ( n25866 , n20921 , n25106 );
    nor g4063 ( n20991 , n14539 , n12878 );
    or g4064 ( n22976 , n4555 , n11736 );
    and g4065 ( n16991 , n18856 , n7413 );
    xnor g4066 ( n17343 , n22021 , n1441 );
    xnor g4067 ( n23495 , n22655 , n13189 );
    not g4068 ( n11350 , n19863 );
    nor g4069 ( n18966 , n302 , n16672 );
    nor g4070 ( n10102 , n23170 , n20655 );
    and g4071 ( n3926 , n21414 , n24577 );
    not g4072 ( n19757 , n25977 );
    nor g4073 ( n20229 , n15688 , n26912 );
    and g4074 ( n19436 , n12519 , n21571 );
    or g4075 ( n18733 , n7106 , n12750 );
    and g4076 ( n25980 , n21937 , n17431 );
    nor g4077 ( n20140 , n12098 , n21522 );
    xnor g4078 ( n18500 , n13724 , n17398 );
    or g4079 ( n9918 , n2281 , n17343 );
    not g4080 ( n5410 , n26189 );
    or g4081 ( n16976 , n26319 , n9610 );
    xnor g4082 ( n8274 , n18947 , n10331 );
    nor g4083 ( n1272 , n24031 , n19033 );
    and g4084 ( n27064 , n17341 , n2672 );
    or g4085 ( n23149 , n5019 , n25851 );
    and g4086 ( n17764 , n13118 , n4694 );
    xnor g4087 ( n13439 , n21066 , n12509 );
    not g4088 ( n3526 , n2981 );
    xnor g4089 ( n26965 , n23089 , n9830 );
    nor g4090 ( n26407 , n20011 , n5697 );
    and g4091 ( n14178 , n780 , n15811 );
    or g4092 ( n705 , n11455 , n9940 );
    nor g4093 ( n24530 , n19509 , n4924 );
    or g4094 ( n16819 , n11378 , n9754 );
    and g4095 ( n21950 , n18684 , n3688 );
    not g4096 ( n19218 , n15764 );
    xnor g4097 ( n24578 , n4251 , n23361 );
    not g4098 ( n6693 , n19647 );
    xnor g4099 ( n6483 , n5983 , n2265 );
    xnor g4100 ( n9685 , n18371 , n7933 );
    xnor g4101 ( n5176 , n16638 , n12380 );
    not g4102 ( n19057 , n8629 );
    xnor g4103 ( n9476 , n9319 , n1810 );
    not g4104 ( n12251 , n24137 );
    not g4105 ( n7167 , n25430 );
    and g4106 ( n5116 , n25010 , n7087 );
    xnor g4107 ( n10430 , n12338 , n26856 );
    not g4108 ( n11695 , n13479 );
    and g4109 ( n12334 , n9209 , n25992 );
    and g4110 ( n12527 , n6609 , n21220 );
    or g4111 ( n8474 , n18593 , n1544 );
    nor g4112 ( n19950 , n7818 , n7320 );
    not g4113 ( n23740 , n18727 );
    not g4114 ( n23589 , n23203 );
    and g4115 ( n8902 , n23795 , n22883 );
    and g4116 ( n15900 , n25043 , n17901 );
    nor g4117 ( n17543 , n24417 , n15271 );
    nor g4118 ( n22703 , n26999 , n3990 );
    xor g4119 ( n5599 , n7074 , n3559 );
    not g4120 ( n8714 , n10797 );
    xnor g4121 ( n20997 , n644 , n154 );
    or g4122 ( n3035 , n20700 , n26240 );
    or g4123 ( n15386 , n5368 , n3360 );
    or g4124 ( n4183 , n23845 , n20548 );
    and g4125 ( n10337 , n20613 , n14138 );
    or g4126 ( n10850 , n561 , n16278 );
    or g4127 ( n2752 , n19673 , n22743 );
    or g4128 ( n12748 , n4365 , n16303 );
    nor g4129 ( n3908 , n25164 , n10689 );
    nor g4130 ( n6499 , n11893 , n11337 );
    xnor g4131 ( n2456 , n14251 , n1742 );
    or g4132 ( n10787 , n3959 , n11810 );
    xnor g4133 ( n1267 , n17265 , n17458 );
    not g4134 ( n26289 , n15883 );
    or g4135 ( n15061 , n19163 , n10513 );
    or g4136 ( n15444 , n7237 , n16351 );
    or g4137 ( n23773 , n22447 , n7047 );
    and g4138 ( n13824 , n18410 , n11762 );
    not g4139 ( n8068 , n21095 );
    or g4140 ( n3863 , n9752 , n4467 );
    not g4141 ( n816 , n5794 );
    nor g4142 ( n20132 , n26529 , n3939 );
    and g4143 ( n8059 , n2121 , n4213 );
    or g4144 ( n14245 , n24866 , n3826 );
    or g4145 ( n19011 , n10346 , n2163 );
    nor g4146 ( n17099 , n16022 , n18575 );
    xnor g4147 ( n10183 , n9207 , n19577 );
    and g4148 ( n20812 , n4483 , n3566 );
    not g4149 ( n23209 , n3769 );
    or g4150 ( n965 , n8144 , n17792 );
    xnor g4151 ( n2878 , n5996 , n2528 );
    or g4152 ( n18618 , n3666 , n3926 );
    or g4153 ( n26933 , n20924 , n7869 );
    not g4154 ( n25038 , n3324 );
    xnor g4155 ( n22625 , n7609 , n21496 );
    and g4156 ( n4727 , n18814 , n9037 );
    or g4157 ( n11635 , n21867 , n22248 );
    not g4158 ( n11152 , n20604 );
    xnor g4159 ( n13988 , n6566 , n9509 );
    not g4160 ( n17883 , n197 );
    xnor g4161 ( n5548 , n6025 , n13941 );
    xnor g4162 ( n11330 , n6771 , n5074 );
    or g4163 ( n9250 , n6117 , n25901 );
    xnor g4164 ( n17421 , n2364 , n803 );
    and g4165 ( n21329 , n6742 , n7510 );
    or g4166 ( n10952 , n13268 , n11729 );
    and g4167 ( n5269 , n192 , n12706 );
    or g4168 ( n2712 , n20575 , n11933 );
    or g4169 ( n15005 , n19973 , n14794 );
    and g4170 ( n17223 , n2566 , n4894 );
    and g4171 ( n24884 , n11763 , n2888 );
    nor g4172 ( n10894 , n14016 , n22282 );
    xnor g4173 ( n24475 , n13289 , n14927 );
    or g4174 ( n19659 , n15826 , n20438 );
    and g4175 ( n11123 , n4589 , n6370 );
    not g4176 ( n24098 , n10117 );
    and g4177 ( n210 , n22708 , n3757 );
    or g4178 ( n7908 , n7537 , n21724 );
    xnor g4179 ( n5367 , n2878 , n13775 );
    and g4180 ( n25402 , n15447 , n24951 );
    xnor g4181 ( n5224 , n8745 , n26913 );
    xnor g4182 ( n6462 , n22219 , n12514 );
    xnor g4183 ( n14947 , n16396 , n18295 );
    not g4184 ( n16474 , n11926 );
    or g4185 ( n18561 , n8101 , n9468 );
    or g4186 ( n2859 , n16568 , n183 );
    not g4187 ( n2864 , n12679 );
    or g4188 ( n937 , n10554 , n330 );
    and g4189 ( n7846 , n1355 , n20363 );
    xnor g4190 ( n325 , n23235 , n8253 );
    and g4191 ( n7499 , n2006 , n22453 );
    and g4192 ( n22101 , n13569 , n7374 );
    xnor g4193 ( n20693 , n8695 , n19932 );
    not g4194 ( n17616 , n81 );
    xnor g4195 ( n19873 , n14611 , n742 );
    xnor g4196 ( n15477 , n20561 , n3735 );
    nor g4197 ( n23043 , n11615 , n23018 );
    or g4198 ( n262 , n15717 , n15611 );
    or g4199 ( n23676 , n19 , n24875 );
    or g4200 ( n12393 , n2309 , n15845 );
    not g4201 ( n4558 , n25656 );
    xnor g4202 ( n1572 , n24481 , n21905 );
    xnor g4203 ( n7775 , n13068 , n826 );
    and g4204 ( n1206 , n16761 , n19169 );
    not g4205 ( n14937 , n23475 );
    or g4206 ( n16367 , n8513 , n415 );
    and g4207 ( n20971 , n19430 , n20337 );
    xnor g4208 ( n9775 , n2071 , n8285 );
    not g4209 ( n21433 , n26185 );
    xnor g4210 ( n16080 , n171 , n10260 );
    xnor g4211 ( n15643 , n13363 , n2828 );
    xnor g4212 ( n19063 , n1631 , n21247 );
    or g4213 ( n16958 , n7088 , n20393 );
    not g4214 ( n23970 , n20564 );
    and g4215 ( n20938 , n11692 , n16710 );
    and g4216 ( n6666 , n1871 , n18083 );
    nor g4217 ( n20345 , n13967 , n9655 );
    or g4218 ( n15945 , n13309 , n24278 );
    nor g4219 ( n13244 , n10441 , n6727 );
    or g4220 ( n10450 , n6275 , n2075 );
    and g4221 ( n4526 , n140 , n22354 );
    xnor g4222 ( n1238 , n1145 , n11794 );
    xnor g4223 ( n1292 , n14761 , n26460 );
    and g4224 ( n3841 , n16387 , n507 );
    or g4225 ( n3457 , n643 , n17804 );
    or g4226 ( n3866 , n19398 , n20050 );
    nor g4227 ( n12857 , n17458 , n23064 );
    xnor g4228 ( n14059 , n2714 , n24837 );
    not g4229 ( n8000 , n17999 );
    or g4230 ( n351 , n269 , n24719 );
    not g4231 ( n8496 , n6281 );
    not g4232 ( n2801 , n650 );
    or g4233 ( n25545 , n7292 , n546 );
    not g4234 ( n12422 , n14444 );
    or g4235 ( n8924 , n10863 , n16581 );
    or g4236 ( n25410 , n9661 , n14850 );
    or g4237 ( n11777 , n4045 , n23688 );
    xnor g4238 ( n12211 , n27083 , n3508 );
    xnor g4239 ( n26461 , n21681 , n256 );
    xnor g4240 ( n8041 , n23626 , n16149 );
    xnor g4241 ( n18707 , n1343 , n26748 );
    not g4242 ( n8713 , n26583 );
    not g4243 ( n23244 , n1639 );
    xnor g4244 ( n18694 , n16427 , n17888 );
    not g4245 ( n4031 , n14723 );
    and g4246 ( n4430 , n25136 , n15005 );
    and g4247 ( n18565 , n8953 , n6594 );
    and g4248 ( n5600 , n1294 , n1585 );
    or g4249 ( n795 , n2483 , n6079 );
    and g4250 ( n11726 , n1064 , n11436 );
    or g4251 ( n17611 , n12682 , n817 );
    or g4252 ( n18082 , n10655 , n18064 );
    xnor g4253 ( n16684 , n22967 , n24542 );
    xnor g4254 ( n23103 , n13197 , n17674 );
    nor g4255 ( n4286 , n18514 , n11597 );
    not g4256 ( n14643 , n19158 );
    or g4257 ( n23378 , n19830 , n21457 );
    or g4258 ( n5076 , n21764 , n16026 );
    or g4259 ( n14227 , n12920 , n18557 );
    xnor g4260 ( n10829 , n12744 , n816 );
    xnor g4261 ( n15226 , n26215 , n22083 );
    nor g4262 ( n10029 , n10918 , n5633 );
    or g4263 ( n766 , n25168 , n17094 );
    or g4264 ( n11218 , n1327 , n13201 );
    or g4265 ( n9428 , n11554 , n2964 );
    or g4266 ( n25090 , n17013 , n23974 );
    or g4267 ( n20420 , n22841 , n9935 );
    or g4268 ( n24730 , n22963 , n7110 );
    or g4269 ( n17879 , n23084 , n3870 );
    nor g4270 ( n8425 , n25074 , n10053 );
    xnor g4271 ( n17142 , n17483 , n24573 );
    and g4272 ( n7845 , n24906 , n8397 );
    and g4273 ( n13855 , n8100 , n2481 );
    nor g4274 ( n15395 , n23359 , n19444 );
    not g4275 ( n14465 , n12956 );
    or g4276 ( n8459 , n11186 , n26054 );
    or g4277 ( n3937 , n571 , n23499 );
    or g4278 ( n26297 , n19282 , n23709 );
    or g4279 ( n11142 , n22462 , n10994 );
    xnor g4280 ( n4154 , n7149 , n22871 );
    nor g4281 ( n16567 , n14230 , n19922 );
    and g4282 ( n23824 , n13871 , n20746 );
    not g4283 ( n17725 , n11751 );
    not g4284 ( n19814 , n11539 );
    or g4285 ( n4965 , n15055 , n5270 );
    nor g4286 ( n2556 , n9247 , n18715 );
    xnor g4287 ( n8140 , n8569 , n13119 );
    xnor g4288 ( n3827 , n24777 , n5940 );
    and g4289 ( n16782 , n13346 , n15592 );
    and g4290 ( n2018 , n5775 , n15934 );
    and g4291 ( n14959 , n18069 , n1130 );
    and g4292 ( n12133 , n25661 , n25182 );
    not g4293 ( n7605 , n6175 );
    not g4294 ( n22182 , n25251 );
    nor g4295 ( n24785 , n26209 , n10462 );
    or g4296 ( n8262 , n5204 , n1761 );
    and g4297 ( n3948 , n17333 , n14783 );
    nor g4298 ( n15577 , n23095 , n22332 );
    not g4299 ( n10184 , n11736 );
    not g4300 ( n22651 , n16722 );
    xnor g4301 ( n17687 , n764 , n8798 );
    xnor g4302 ( n22121 , n16119 , n4739 );
    or g4303 ( n26457 , n21691 , n16158 );
    or g4304 ( n26284 , n3968 , n6070 );
    xnor g4305 ( n14267 , n22109 , n18168 );
    nor g4306 ( n15529 , n12446 , n1112 );
    and g4307 ( n19010 , n5761 , n7955 );
    not g4308 ( n9880 , n18151 );
    xnor g4309 ( n4232 , n15743 , n2809 );
    and g4310 ( n7186 , n4414 , n17019 );
    not g4311 ( n13378 , n8285 );
    xnor g4312 ( n3158 , n20250 , n1682 );
    xnor g4313 ( n12322 , n16412 , n25214 );
    or g4314 ( n10256 , n25259 , n14757 );
    and g4315 ( n2902 , n2155 , n7097 );
    and g4316 ( n13584 , n12126 , n7023 );
    not g4317 ( n427 , n14424 );
    and g4318 ( n9207 , n22931 , n3701 );
    xnor g4319 ( n19686 , n24802 , n9359 );
    not g4320 ( n4569 , n3247 );
    not g4321 ( n7364 , n19560 );
    xnor g4322 ( n19924 , n4866 , n1809 );
    or g4323 ( n14128 , n10146 , n21753 );
    xnor g4324 ( n22407 , n24202 , n18274 );
    and g4325 ( n25340 , n12197 , n10068 );
    or g4326 ( n20961 , n16783 , n21891 );
    nor g4327 ( n930 , n22527 , n19820 );
    xnor g4328 ( n18511 , n24066 , n12555 );
    nor g4329 ( n23719 , n23547 , n25569 );
    xnor g4330 ( n21426 , n2360 , n22764 );
    or g4331 ( n22094 , n8261 , n18905 );
    not g4332 ( n21066 , n18333 );
    not g4333 ( n8937 , n5696 );
    or g4334 ( n11813 , n12918 , n1758 );
    or g4335 ( n5828 , n15684 , n1852 );
    nor g4336 ( n14578 , n115 , n22859 );
    or g4337 ( n25013 , n18485 , n12811 );
    not g4338 ( n20011 , n7825 );
    xnor g4339 ( n17589 , n2093 , n18520 );
    nor g4340 ( n14800 , n5714 , n1222 );
    and g4341 ( n2484 , n3537 , n7542 );
    not g4342 ( n21209 , n2953 );
    xnor g4343 ( n48 , n17034 , n23951 );
    and g4344 ( n25031 , n7929 , n24581 );
    and g4345 ( n18007 , n4707 , n19622 );
    xnor g4346 ( n10725 , n25120 , n23272 );
    nor g4347 ( n20836 , n25514 , n13696 );
    xnor g4348 ( n16582 , n14489 , n18317 );
    and g4349 ( n13219 , n3259 , n21720 );
    or g4350 ( n24994 , n9466 , n21798 );
    xnor g4351 ( n17729 , n4542 , n18295 );
    xnor g4352 ( n16261 , n1990 , n14548 );
    or g4353 ( n8696 , n29 , n14372 );
    or g4354 ( n10264 , n18746 , n26452 );
    or g4355 ( n15043 , n10061 , n5027 );
    nor g4356 ( n6768 , n21333 , n20098 );
    and g4357 ( n517 , n18564 , n9562 );
    or g4358 ( n20390 , n9755 , n18048 );
    and g4359 ( n24733 , n16839 , n19030 );
    not g4360 ( n20075 , n24051 );
    or g4361 ( n1228 , n7768 , n1345 );
    xnor g4362 ( n14364 , n3839 , n10363 );
    xnor g4363 ( n4869 , n12298 , n22400 );
    and g4364 ( n817 , n6258 , n18801 );
    or g4365 ( n12974 , n9310 , n24115 );
    or g4366 ( n3059 , n10622 , n501 );
    xnor g4367 ( n14217 , n11662 , n11775 );
    or g4368 ( n2167 , n20991 , n20699 );
    xnor g4369 ( n11254 , n1241 , n11803 );
    xnor g4370 ( n4937 , n8656 , n9380 );
    nor g4371 ( n17848 , n6051 , n15053 );
    and g4372 ( n134 , n16393 , n16627 );
    xnor g4373 ( n709 , n14959 , n3183 );
    or g4374 ( n10083 , n26901 , n22807 );
    and g4375 ( n1900 , n7812 , n495 );
    xnor g4376 ( n6344 , n12673 , n25220 );
    or g4377 ( n16431 , n11513 , n4111 );
    nor g4378 ( n14866 , n22173 , n12593 );
    and g4379 ( n7480 , n25143 , n25988 );
    or g4380 ( n1471 , n2079 , n12095 );
    xnor g4381 ( n14048 , n22128 , n3151 );
    or g4382 ( n8867 , n25628 , n23432 );
    xnor g4383 ( n16816 , n3608 , n24263 );
    xnor g4384 ( n9699 , n26440 , n7990 );
    and g4385 ( n18915 , n23081 , n6205 );
    or g4386 ( n14497 , n16680 , n15692 );
    and g4387 ( n1875 , n26071 , n1425 );
    not g4388 ( n15337 , n10915 );
    or g4389 ( n8424 , n15217 , n15241 );
    or g4390 ( n23090 , n2080 , n1319 );
    or g4391 ( n18351 , n8910 , n19321 );
    xnor g4392 ( n11866 , n6127 , n4642 );
    not g4393 ( n18130 , n18479 );
    not g4394 ( n14042 , n22031 );
    and g4395 ( n21754 , n1390 , n7495 );
    or g4396 ( n16863 , n1161 , n377 );
    not g4397 ( n18715 , n3663 );
    or g4398 ( n5797 , n6788 , n18590 );
    xnor g4399 ( n19323 , n16603 , n11300 );
    or g4400 ( n13267 , n26777 , n17 );
    xnor g4401 ( n18418 , n1390 , n10240 );
    xnor g4402 ( n12386 , n5823 , n6513 );
    xnor g4403 ( n15382 , n3820 , n3684 );
    or g4404 ( n18957 , n22017 , n22671 );
    and g4405 ( n19416 , n26916 , n24288 );
    not g4406 ( n11135 , n13356 );
    and g4407 ( n23504 , n5740 , n14653 );
    or g4408 ( n16867 , n6872 , n16559 );
    and g4409 ( n27082 , n12418 , n21959 );
    not g4410 ( n16205 , n18907 );
    xnor g4411 ( n9088 , n8614 , n25972 );
    and g4412 ( n18188 , n11099 , n26751 );
    nor g4413 ( n4056 , n11457 , n15636 );
    not g4414 ( n25451 , n9889 );
    nor g4415 ( n6574 , n11938 , n19472 );
    or g4416 ( n23702 , n21915 , n2509 );
    nor g4417 ( n3334 , n17125 , n10532 );
    xnor g4418 ( n24861 , n4957 , n7421 );
    or g4419 ( n25182 , n3408 , n2484 );
    or g4420 ( n9933 , n6039 , n10199 );
    and g4421 ( n10936 , n17732 , n20823 );
    xnor g4422 ( n829 , n13063 , n6278 );
    or g4423 ( n27013 , n11750 , n9270 );
    xnor g4424 ( n16596 , n26293 , n26128 );
    not g4425 ( n18335 , n7773 );
    nor g4426 ( n19596 , n4230 , n8378 );
    not g4427 ( n1719 , n3705 );
    xnor g4428 ( n9707 , n20169 , n1949 );
    nor g4429 ( n16947 , n23487 , n6556 );
    and g4430 ( n9263 , n21124 , n3295 );
    xnor g4431 ( n18488 , n16204 , n26117 );
    not g4432 ( n19702 , n18972 );
    and g4433 ( n4053 , n22743 , n2346 );
    xnor g4434 ( n23619 , n9785 , n16199 );
    nor g4435 ( n6547 , n10602 , n21721 );
    not g4436 ( n22812 , n4491 );
    or g4437 ( n11357 , n16211 , n4256 );
    or g4438 ( n16664 , n21937 , n14007 );
    and g4439 ( n18396 , n8903 , n3950 );
    or g4440 ( n20188 , n862 , n20386 );
    or g4441 ( n10121 , n25161 , n8287 );
    xnor g4442 ( n18116 , n12446 , n1112 );
    xnor g4443 ( n8206 , n16478 , n3461 );
    and g4444 ( n15788 , n15148 , n452 );
    or g4445 ( n7299 , n18499 , n19009 );
    nor g4446 ( n23695 , n21276 , n23061 );
    not g4447 ( n24221 , n5718 );
    nor g4448 ( n3197 , n3908 , n16490 );
    or g4449 ( n3517 , n3016 , n7827 );
    or g4450 ( n7700 , n26495 , n5789 );
    and g4451 ( n5199 , n22060 , n594 );
    and g4452 ( n6667 , n2708 , n12528 );
    and g4453 ( n25269 , n6781 , n25477 );
    and g4454 ( n14069 , n5373 , n14558 );
    xnor g4455 ( n19118 , n19245 , n9584 );
    not g4456 ( n12441 , n21184 );
    or g4457 ( n5014 , n21649 , n20192 );
    xnor g4458 ( n5427 , n6180 , n25487 );
    xnor g4459 ( n1309 , n23583 , n22531 );
    xnor g4460 ( n11970 , n22938 , n13732 );
    or g4461 ( n10168 , n8910 , n19201 );
    xnor g4462 ( n17235 , n16042 , n11955 );
    xnor g4463 ( n9833 , n25350 , n3889 );
    xnor g4464 ( n2229 , n10372 , n12152 );
    nor g4465 ( n13547 , n13569 , n7374 );
    xnor g4466 ( n19486 , n25804 , n13350 );
    not g4467 ( n23091 , n14393 );
    nor g4468 ( n1299 , n7566 , n22640 );
    not g4469 ( n3359 , n1528 );
    or g4470 ( n14388 , n21610 , n6151 );
    and g4471 ( n4226 , n14884 , n18533 );
    xnor g4472 ( n19271 , n4495 , n15666 );
    xnor g4473 ( n5195 , n2152 , n25156 );
    xnor g4474 ( n17452 , n7913 , n23541 );
    nor g4475 ( n20695 , n8411 , n945 );
    and g4476 ( n5460 , n16034 , n10451 );
    nor g4477 ( n2264 , n23864 , n12693 );
    or g4478 ( n17523 , n12474 , n23109 );
    or g4479 ( n24909 , n20416 , n12563 );
    nor g4480 ( n8636 , n3515 , n93 );
    or g4481 ( n22650 , n6264 , n3804 );
    and g4482 ( n17680 , n22672 , n16404 );
    and g4483 ( n3417 , n6981 , n11825 );
    nor g4484 ( n15463 , n23529 , n9124 );
    nor g4485 ( n2692 , n24615 , n1742 );
    xnor g4486 ( n8017 , n6729 , n10792 );
    xnor g4487 ( n1724 , n18715 , n6178 );
    xnor g4488 ( n3508 , n1019 , n11011 );
    xnor g4489 ( n20613 , n13019 , n10108 );
    xnor g4490 ( n9426 , n19312 , n17928 );
    and g4491 ( n13032 , n24674 , n19846 );
    and g4492 ( n6 , n24004 , n12900 );
    or g4493 ( n8045 , n18220 , n8420 );
    or g4494 ( n20584 , n8372 , n20378 );
    not g4495 ( n1864 , n19515 );
    and g4496 ( n14080 , n7704 , n21318 );
    or g4497 ( n3974 , n771 , n23383 );
    and g4498 ( n2513 , n15110 , n19292 );
    and g4499 ( n18654 , n26926 , n22245 );
    or g4500 ( n25274 , n18473 , n4812 );
    not g4501 ( n4395 , n18895 );
    or g4502 ( n26926 , n25250 , n18793 );
    xnor g4503 ( n7608 , n22895 , n27200 );
    or g4504 ( n14413 , n19359 , n9781 );
    xnor g4505 ( n3063 , n23559 , n11481 );
    or g4506 ( n27162 , n1030 , n19240 );
    and g4507 ( n21431 , n19770 , n12022 );
    or g4508 ( n13203 , n16205 , n26823 );
    or g4509 ( n19056 , n2915 , n10224 );
    nor g4510 ( n18908 , n11792 , n22571 );
    or g4511 ( n26395 , n2986 , n25422 );
    xnor g4512 ( n3189 , n3568 , n22934 );
    xnor g4513 ( n925 , n16064 , n19460 );
    and g4514 ( n5124 , n14436 , n8992 );
    or g4515 ( n22587 , n22919 , n24506 );
    buf g4516 ( n18639 , n3223 );
    or g4517 ( n12866 , n25208 , n26299 );
    xnor g4518 ( n26303 , n24037 , n13812 );
    or g4519 ( n17661 , n7043 , n10616 );
    or g4520 ( n25371 , n23555 , n18269 );
    not g4521 ( n16572 , n16302 );
    not g4522 ( n3133 , n2408 );
    xnor g4523 ( n22548 , n7972 , n12659 );
    nor g4524 ( n17217 , n12019 , n2512 );
    or g4525 ( n6717 , n17160 , n5927 );
    and g4526 ( n2987 , n8023 , n19447 );
    xnor g4527 ( n19756 , n17594 , n4738 );
    xnor g4528 ( n16221 , n23012 , n1851 );
    xnor g4529 ( n17159 , n6226 , n4564 );
    and g4530 ( n11869 , n21807 , n1417 );
    or g4531 ( n15543 , n5145 , n9886 );
    and g4532 ( n2213 , n10570 , n13374 );
    xnor g4533 ( n12658 , n4981 , n15152 );
    and g4534 ( n21393 , n13781 , n26793 );
    nor g4535 ( n8605 , n13480 , n16544 );
    and g4536 ( n15237 , n246 , n17401 );
    or g4537 ( n23828 , n13503 , n25575 );
    and g4538 ( n13259 , n15107 , n15954 );
    xnor g4539 ( n8629 , n17645 , n10945 );
    xnor g4540 ( n14342 , n26679 , n26419 );
    nor g4541 ( n13092 , n25514 , n4361 );
    and g4542 ( n24382 , n6834 , n5165 );
    xnor g4543 ( n20233 , n19127 , n21727 );
    xnor g4544 ( n6263 , n27183 , n4185 );
    or g4545 ( n12691 , n22149 , n23134 );
    not g4546 ( n16975 , n22686 );
    not g4547 ( n2000 , n13158 );
    nor g4548 ( n14162 , n14907 , n25238 );
    or g4549 ( n18533 , n2446 , n15969 );
    and g4550 ( n26244 , n18702 , n22668 );
    xnor g4551 ( n3743 , n10918 , n9731 );
    xnor g4552 ( n4835 , n20489 , n26913 );
    or g4553 ( n11562 , n25054 , n10138 );
    and g4554 ( n6938 , n4722 , n6403 );
    xnor g4555 ( n24458 , n7903 , n6450 );
    and g4556 ( n4918 , n7335 , n11578 );
    xnor g4557 ( n24056 , n19444 , n2979 );
    nor g4558 ( n2480 , n24924 , n20876 );
    and g4559 ( n26026 , n2153 , n5018 );
    or g4560 ( n4274 , n6492 , n17718 );
    xnor g4561 ( n26689 , n25431 , n16824 );
    and g4562 ( n7875 , n12619 , n20115 );
    and g4563 ( n6668 , n18320 , n12653 );
    xnor g4564 ( n7308 , n20130 , n10599 );
    and g4565 ( n24235 , n20481 , n2620 );
    xnor g4566 ( n17671 , n6295 , n9709 );
    and g4567 ( n669 , n13647 , n18109 );
    xnor g4568 ( n19248 , n15739 , n12507 );
    xnor g4569 ( n17472 , n5685 , n189 );
    and g4570 ( n6767 , n4604 , n8116 );
    xnor g4571 ( n649 , n13645 , n12001 );
    xnor g4572 ( n4753 , n22066 , n25130 );
    and g4573 ( n7165 , n25391 , n19855 );
    or g4574 ( n22373 , n2821 , n13594 );
    or g4575 ( n20882 , n14910 , n21250 );
    xnor g4576 ( n19331 , n3920 , n1993 );
    xnor g4577 ( n23875 , n13360 , n26544 );
    or g4578 ( n18178 , n4309 , n14727 );
    xnor g4579 ( n20247 , n26186 , n19556 );
    not g4580 ( n505 , n3037 );
    xnor g4581 ( n1622 , n26180 , n10650 );
    or g4582 ( n16737 , n7662 , n16616 );
    xnor g4583 ( n25949 , n15064 , n12861 );
    or g4584 ( n25517 , n14564 , n9809 );
    not g4585 ( n218 , n12125 );
    nor g4586 ( n4717 , n22724 , n19614 );
    or g4587 ( n7219 , n1257 , n1369 );
    or g4588 ( n1828 , n7584 , n13221 );
    xnor g4589 ( n23480 , n10600 , n18683 );
    or g4590 ( n8127 , n23347 , n23452 );
    not g4591 ( n19061 , n25693 );
    buf g4592 ( n16244 , n15972 );
    xnor g4593 ( n18771 , n13018 , n22290 );
    or g4594 ( n12963 , n22631 , n8819 );
    and g4595 ( n72 , n25301 , n26679 );
    xnor g4596 ( n9133 , n23948 , n3193 );
    and g4597 ( n14788 , n17284 , n7896 );
    xnor g4598 ( n24955 , n24600 , n3641 );
    or g4599 ( n26125 , n26722 , n15074 );
    or g4600 ( n13380 , n7948 , n1583 );
    or g4601 ( n18844 , n2077 , n11749 );
    and g4602 ( n5649 , n23038 , n23286 );
    and g4603 ( n3200 , n4190 , n10328 );
    xnor g4604 ( n23588 , n15674 , n25503 );
    nor g4605 ( n12136 , n3276 , n268 );
    or g4606 ( n17271 , n25436 , n8162 );
    xnor g4607 ( n12616 , n20934 , n2306 );
    xnor g4608 ( n14782 , n8369 , n15120 );
    nor g4609 ( n12572 , n17900 , n16459 );
    not g4610 ( n17397 , n18139 );
    or g4611 ( n4716 , n10381 , n1772 );
    or g4612 ( n5820 , n25650 , n7177 );
    xnor g4613 ( n15705 , n14165 , n17729 );
    not g4614 ( n2125 , n2886 );
    nor g4615 ( n7187 , n15309 , n3846 );
    or g4616 ( n17174 , n24752 , n4082 );
    xnor g4617 ( n4887 , n5698 , n27173 );
    nor g4618 ( n21161 , n22433 , n10158 );
    and g4619 ( n25862 , n3571 , n4607 );
    not g4620 ( n23806 , n8317 );
    nor g4621 ( n10990 , n10201 , n11336 );
    and g4622 ( n19879 , n12240 , n14833 );
    or g4623 ( n15372 , n22485 , n1100 );
    xnor g4624 ( n9881 , n17545 , n8750 );
    or g4625 ( n11435 , n12533 , n7942 );
    or g4626 ( n4023 , n1298 , n8203 );
    nor g4627 ( n13576 , n14251 , n26946 );
    not g4628 ( n23760 , n3552 );
    not g4629 ( n8220 , n12094 );
    and g4630 ( n21510 , n24131 , n25260 );
    nor g4631 ( n24691 , n26417 , n6789 );
    or g4632 ( n18397 , n24031 , n17993 );
    not g4633 ( n13715 , n2987 );
    or g4634 ( n1651 , n94 , n9476 );
    and g4635 ( n24175 , n8747 , n3212 );
    xnor g4636 ( n16555 , n11341 , n25365 );
    xnor g4637 ( n9558 , n6743 , n23152 );
    and g4638 ( n10401 , n15125 , n11929 );
    xnor g4639 ( n10718 , n11314 , n25738 );
    or g4640 ( n23553 , n24018 , n1654 );
    xnor g4641 ( n25786 , n23497 , n21004 );
    not g4642 ( n13117 , n17606 );
    and g4643 ( n1033 , n19612 , n24459 );
    xnor g4644 ( n4277 , n22292 , n14589 );
    and g4645 ( n21413 , n9618 , n14629 );
    xnor g4646 ( n13987 , n9151 , n7569 );
    or g4647 ( n21347 , n20128 , n7862 );
    xnor g4648 ( n24451 , n21973 , n24916 );
    xnor g4649 ( n585 , n12702 , n12507 );
    xnor g4650 ( n1683 , n24638 , n442 );
    or g4651 ( n9307 , n5908 , n792 );
    or g4652 ( n4779 , n7431 , n26178 );
    nor g4653 ( n3801 , n14528 , n16019 );
    or g4654 ( n16151 , n15622 , n633 );
    xnor g4655 ( n18513 , n4864 , n13266 );
    and g4656 ( n9489 , n5760 , n13954 );
    or g4657 ( n19599 , n12554 , n21083 );
    nor g4658 ( n12768 , n8773 , n10610 );
    or g4659 ( n24321 , n7892 , n15734 );
    or g4660 ( n27109 , n23868 , n2154 );
    or g4661 ( n26246 , n18220 , n21577 );
    and g4662 ( n23104 , n21812 , n14568 );
    not g4663 ( n12845 , n14996 );
    not g4664 ( n7471 , n22744 );
    or g4665 ( n8080 , n7551 , n20535 );
    not g4666 ( n13535 , n22824 );
    xnor g4667 ( n16536 , n25824 , n2349 );
    xnor g4668 ( n5411 , n25313 , n24859 );
    nor g4669 ( n12666 , n24788 , n6025 );
    not g4670 ( n4883 , n9431 );
    and g4671 ( n59 , n19395 , n5497 );
    nor g4672 ( n21702 , n10514 , n6105 );
    and g4673 ( n11230 , n21775 , n2793 );
    xnor g4674 ( n2698 , n20738 , n3158 );
    and g4675 ( n13287 , n27120 , n25504 );
    xnor g4676 ( n23789 , n6594 , n6559 );
    or g4677 ( n13805 , n7453 , n20847 );
    xnor g4678 ( n17028 , n125 , n2659 );
    nor g4679 ( n16670 , n26629 , n19904 );
    or g4680 ( n13892 , n24947 , n19277 );
    xnor g4681 ( n25520 , n3258 , n12108 );
    and g4682 ( n6426 , n12513 , n25568 );
    or g4683 ( n1311 , n20053 , n6887 );
    or g4684 ( n16936 , n24193 , n10977 );
    not g4685 ( n16548 , n11336 );
    and g4686 ( n4052 , n20028 , n18087 );
    and g4687 ( n3144 , n3372 , n2451 );
    xnor g4688 ( n2092 , n5973 , n26838 );
    or g4689 ( n3251 , n4858 , n602 );
    or g4690 ( n17361 , n24181 , n21938 );
    buf g4691 ( n9469 , n3051 );
    or g4692 ( n20980 , n12831 , n8554 );
    not g4693 ( n5516 , n16158 );
    or g4694 ( n10428 , n18297 , n22378 );
    nor g4695 ( n24216 , n23791 , n7083 );
    xnor g4696 ( n25550 , n7076 , n14005 );
    nor g4697 ( n24565 , n13839 , n14218 );
    nor g4698 ( n13751 , n15761 , n12445 );
    and g4699 ( n813 , n25492 , n8029 );
    or g4700 ( n15330 , n12768 , n18508 );
    and g4701 ( n11397 , n26434 , n18543 );
    or g4702 ( n5735 , n3945 , n21998 );
    xnor g4703 ( n21751 , n17499 , n11474 );
    nor g4704 ( n24230 , n24164 , n23475 );
    not g4705 ( n20556 , n21295 );
    not g4706 ( n10425 , n5706 );
    xnor g4707 ( n14466 , n26362 , n17827 );
    xnor g4708 ( n6718 , n6112 , n16797 );
    not g4709 ( n13492 , n20005 );
    xnor g4710 ( n12808 , n4409 , n10125 );
    nor g4711 ( n9198 , n20045 , n14510 );
    and g4712 ( n16542 , n22662 , n16762 );
    and g4713 ( n20469 , n13816 , n14997 );
    nor g4714 ( n20981 , n19404 , n14700 );
    or g4715 ( n628 , n13641 , n16000 );
    xnor g4716 ( n14527 , n6446 , n20060 );
    xnor g4717 ( n4255 , n3136 , n2409 );
    not g4718 ( n12612 , n20959 );
    not g4719 ( n24358 , n12495 );
    and g4720 ( n24227 , n27104 , n13317 );
    xnor g4721 ( n25805 , n25297 , n23857 );
    or g4722 ( n15078 , n11498 , n6316 );
    and g4723 ( n1014 , n23112 , n2 );
    nor g4724 ( n12269 , n13990 , n3744 );
    and g4725 ( n6429 , n1098 , n20448 );
    or g4726 ( n7888 , n26548 , n14658 );
    not g4727 ( n23230 , n1118 );
    not g4728 ( n6916 , n14902 );
    nor g4729 ( n8138 , n12341 , n13945 );
    and g4730 ( n16377 , n460 , n26666 );
    or g4731 ( n77 , n15292 , n15752 );
    not g4732 ( n12068 , n6912 );
    xnor g4733 ( n12488 , n114 , n16093 );
    nor g4734 ( n4270 , n25021 , n10593 );
    nor g4735 ( n27062 , n16705 , n14244 );
    nor g4736 ( n4710 , n14963 , n11579 );
    not g4737 ( n26819 , n8772 );
    xnor g4738 ( n21193 , n20542 , n13697 );
    and g4739 ( n5575 , n21749 , n2298 );
    or g4740 ( n26959 , n8782 , n18643 );
    and g4741 ( n10532 , n15402 , n7309 );
    and g4742 ( n7738 , n3818 , n9795 );
    or g4743 ( n26540 , n6521 , n6659 );
    and g4744 ( n5610 , n23402 , n9283 );
    xnor g4745 ( n5903 , n17849 , n22136 );
    not g4746 ( n1794 , n23779 );
    and g4747 ( n13207 , n9301 , n7718 );
    and g4748 ( n9163 , n11385 , n5422 );
    and g4749 ( n43 , n2592 , n20882 );
    or g4750 ( n3172 , n12454 , n11481 );
    xnor g4751 ( n25474 , n6369 , n3164 );
    nor g4752 ( n4797 , n13319 , n15490 );
    and g4753 ( n25993 , n21388 , n1228 );
    xnor g4754 ( n24330 , n26233 , n21561 );
    not g4755 ( n21698 , n513 );
    xnor g4756 ( n26492 , n14495 , n4271 );
    xnor g4757 ( n2402 , n15405 , n3940 );
    and g4758 ( n11703 , n15564 , n11499 );
    and g4759 ( n23117 , n24673 , n20451 );
    or g4760 ( n12840 , n3150 , n25439 );
    xnor g4761 ( n16905 , n479 , n8701 );
    or g4762 ( n7804 , n23200 , n16077 );
    and g4763 ( n1358 , n2113 , n148 );
    xnor g4764 ( n15365 , n287 , n26160 );
    xnor g4765 ( n414 , n11220 , n12507 );
    not g4766 ( n16345 , n8805 );
    not g4767 ( n255 , n16373 );
    xnor g4768 ( n9268 , n24237 , n19592 );
    nor g4769 ( n9637 , n63 , n13671 );
    xnor g4770 ( n12408 , n12429 , n23424 );
    and g4771 ( n14770 , n1135 , n11839 );
    xnor g4772 ( n14194 , n6232 , n13472 );
    xnor g4773 ( n11271 , n4626 , n21509 );
    xnor g4774 ( n7376 , n26101 , n14046 );
    or g4775 ( n22970 , n21436 , n22983 );
    or g4776 ( n3966 , n23776 , n7417 );
    not g4777 ( n23353 , n348 );
    or g4778 ( n26873 , n621 , n18688 );
    nor g4779 ( n22658 , n20011 , n17953 );
    and g4780 ( n6601 , n24031 , n17993 );
    or g4781 ( n5308 , n18837 , n1321 );
    or g4782 ( n16941 , n20022 , n15141 );
    xnor g4783 ( n13008 , n23160 , n7678 );
    nor g4784 ( n11668 , n23209 , n11755 );
    not g4785 ( n6309 , n2324 );
    or g4786 ( n22118 , n13766 , n6297 );
    or g4787 ( n3430 , n12657 , n10092 );
    or g4788 ( n9185 , n3480 , n7850 );
    and g4789 ( n20752 , n18218 , n7430 );
    or g4790 ( n17594 , n1479 , n16032 );
    xnor g4791 ( n26274 , n14175 , n13658 );
    and g4792 ( n22210 , n2424 , n84 );
    xnor g4793 ( n13884 , n6737 , n17544 );
    xnor g4794 ( n441 , n22662 , n5048 );
    or g4795 ( n16652 , n11226 , n15893 );
    and g4796 ( n5889 , n6687 , n9837 );
    nor g4797 ( n18562 , n23141 , n2035 );
    xnor g4798 ( n21788 , n16197 , n24936 );
    xnor g4799 ( n18791 , n3138 , n24245 );
    not g4800 ( n24575 , n11099 );
    nor g4801 ( n17951 , n24868 , n23268 );
    or g4802 ( n21524 , n15628 , n21722 );
    not g4803 ( n22200 , n11289 );
    nor g4804 ( n3620 , n9671 , n4858 );
    xnor g4805 ( n23411 , n7350 , n1480 );
    or g4806 ( n13084 , n7237 , n4873 );
    and g4807 ( n23075 , n5159 , n11377 );
    nor g4808 ( n5363 , n13953 , n17323 );
    or g4809 ( n5323 , n24949 , n16423 );
    xnor g4810 ( n10141 , n8557 , n24739 );
    nor g4811 ( n8015 , n18598 , n17077 );
    and g4812 ( n7786 , n8885 , n4023 );
    xnor g4813 ( n22006 , n848 , n7864 );
    not g4814 ( n5601 , n5713 );
    not g4815 ( n7422 , n16413 );
    xnor g4816 ( n11234 , n22874 , n25765 );
    nor g4817 ( n21373 , n19258 , n10919 );
    or g4818 ( n4830 , n26798 , n6951 );
    and g4819 ( n23122 , n13591 , n22114 );
    xnor g4820 ( n21728 , n4570 , n17591 );
    and g4821 ( n25794 , n6169 , n26302 );
    not g4822 ( n1046 , n3804 );
    buf g4823 ( n10013 , n14125 );
    and g4824 ( n26260 , n10951 , n13372 );
    xnor g4825 ( n2849 , n3530 , n15857 );
    and g4826 ( n22737 , n11922 , n13639 );
    xnor g4827 ( n7229 , n19622 , n19322 );
    and g4828 ( n25977 , n13707 , n14854 );
    and g4829 ( n14916 , n21429 , n9083 );
    xnor g4830 ( n5850 , n15732 , n9075 );
    and g4831 ( n12930 , n23261 , n24460 );
    and g4832 ( n10341 , n18880 , n26594 );
    or g4833 ( n11024 , n6393 , n7948 );
    and g4834 ( n4831 , n14556 , n1442 );
    and g4835 ( n7899 , n24537 , n11210 );
    or g4836 ( n19169 , n22733 , n16403 );
    xnor g4837 ( n14786 , n23709 , n14268 );
    xnor g4838 ( n7669 , n6749 , n1589 );
    nor g4839 ( n15707 , n8386 , n3217 );
    or g4840 ( n2138 , n2409 , n14071 );
    and g4841 ( n15566 , n16805 , n6906 );
    xnor g4842 ( n24910 , n17485 , n17555 );
    xnor g4843 ( n15057 , n11210 , n24537 );
    xnor g4844 ( n11708 , n726 , n26849 );
    and g4845 ( n24833 , n12594 , n21452 );
    or g4846 ( n1137 , n24116 , n21556 );
    not g4847 ( n8794 , n13372 );
    or g4848 ( n18069 , n9671 , n5205 );
    xnor g4849 ( n15067 , n8436 , n14677 );
    xnor g4850 ( n21045 , n20896 , n6435 );
    or g4851 ( n24199 , n8979 , n9856 );
    or g4852 ( n11012 , n14708 , n19257 );
    not g4853 ( n18814 , n20986 );
    or g4854 ( n14869 , n21127 , n4588 );
    xnor g4855 ( n12964 , n14142 , n10766 );
    or g4856 ( n18380 , n7342 , n5372 );
    nor g4857 ( n22208 , n13775 , n11830 );
    and g4858 ( n26652 , n13427 , n16646 );
    and g4859 ( n9840 , n23218 , n22266 );
    xnor g4860 ( n23816 , n647 , n26408 );
    or g4861 ( n293 , n22732 , n3887 );
    xnor g4862 ( n17398 , n1685 , n15633 );
    nor g4863 ( n15620 , n2432 , n11137 );
    xnor g4864 ( n12319 , n3119 , n7534 );
    or g4865 ( n916 , n2217 , n15038 );
    xnor g4866 ( n5591 , n7689 , n11314 );
    xnor g4867 ( n24711 , n2847 , n16 );
    xnor g4868 ( n4688 , n9485 , n16839 );
    or g4869 ( n17682 , n14736 , n15274 );
    xnor g4870 ( n17856 , n21457 , n20790 );
    or g4871 ( n6594 , n23425 , n12560 );
    and g4872 ( n11373 , n19306 , n14235 );
    xnor g4873 ( n16278 , n23157 , n1863 );
    xnor g4874 ( n21158 , n25929 , n10013 );
    or g4875 ( n13413 , n26172 , n8938 );
    nor g4876 ( n17977 , n22651 , n24552 );
    or g4877 ( n23370 , n5297 , n6697 );
    and g4878 ( n13146 , n5131 , n19674 );
    or g4879 ( n9629 , n20405 , n23113 );
    or g4880 ( n5753 , n22197 , n5927 );
    xnor g4881 ( n17146 , n2894 , n82 );
    and g4882 ( n22308 , n22442 , n22253 );
    not g4883 ( n5987 , n960 );
    xnor g4884 ( n15812 , n8342 , n10906 );
    or g4885 ( n7249 , n20596 , n8771 );
    and g4886 ( n15024 , n14076 , n8901 );
    or g4887 ( n25796 , n16193 , n16001 );
    and g4888 ( n3995 , n17664 , n5115 );
    or g4889 ( n13978 , n26717 , n20020 );
    or g4890 ( n2344 , n5079 , n5008 );
    and g4891 ( n19046 , n4490 , n13167 );
    xnor g4892 ( n6055 , n20597 , n21623 );
    xnor g4893 ( n26269 , n2312 , n25891 );
    xnor g4894 ( n15469 , n11089 , n4955 );
    and g4895 ( n3793 , n15013 , n17961 );
    nor g4896 ( n11133 , n23161 , n22237 );
    or g4897 ( n22816 , n6750 , n19058 );
    and g4898 ( n2873 , n23676 , n5287 );
    or g4899 ( n3418 , n5688 , n6680 );
    or g4900 ( n1473 , n21674 , n22597 );
    or g4901 ( n24349 , n1841 , n25127 );
    xnor g4902 ( n18332 , n25496 , n26566 );
    and g4903 ( n1938 , n22743 , n4708 );
    xnor g4904 ( n8217 , n11028 , n7817 );
    not g4905 ( n7680 , n12766 );
    xnor g4906 ( n14412 , n25497 , n470 );
    and g4907 ( n13738 , n11927 , n14876 );
    xnor g4908 ( n17639 , n20052 , n4182 );
    not g4909 ( n21118 , n22879 );
    or g4910 ( n16892 , n840 , n24620 );
    or g4911 ( n12719 , n24375 , n25119 );
    and g4912 ( n5008 , n2936 , n20430 );
    nor g4913 ( n14472 , n20053 , n18395 );
    and g4914 ( n854 , n9082 , n24346 );
    xnor g4915 ( n24245 , n18461 , n11841 );
    or g4916 ( n20977 , n25142 , n3828 );
    and g4917 ( n269 , n11390 , n7970 );
    or g4918 ( n14213 , n21133 , n25387 );
    xnor g4919 ( n27195 , n9509 , n9554 );
    nor g4920 ( n25506 , n4901 , n20051 );
    and g4921 ( n24 , n24143 , n12420 );
    and g4922 ( n23186 , n445 , n10142 );
    not g4923 ( n4230 , n3878 );
    xnor g4924 ( n12219 , n14684 , n1667 );
    xnor g4925 ( n16626 , n26936 , n20718 );
    xnor g4926 ( n857 , n21081 , n24004 );
    nor g4927 ( n8836 , n6658 , n20141 );
    not g4928 ( n21325 , n4937 );
    xnor g4929 ( n10790 , n12751 , n20982 );
    xnor g4930 ( n19385 , n6994 , n19542 );
    and g4931 ( n6709 , n8958 , n21014 );
    or g4932 ( n5291 , n19516 , n16412 );
    xnor g4933 ( n13667 , n17259 , n7211 );
    or g4934 ( n10580 , n14336 , n7952 );
    or g4935 ( n2067 , n11656 , n1970 );
    or g4936 ( n7093 , n25024 , n25681 );
    and g4937 ( n13041 , n26756 , n26862 );
    and g4938 ( n3389 , n5379 , n3703 );
    or g4939 ( n432 , n14747 , n21445 );
    not g4940 ( n16693 , n23509 );
    or g4941 ( n8326 , n19446 , n3931 );
    xnor g4942 ( n8803 , n8995 , n25925 );
    or g4943 ( n6269 , n17378 , n16603 );
    nor g4944 ( n8270 , n9180 , n15884 );
    or g4945 ( n9484 , n7130 , n12851 );
    not g4946 ( n6935 , n20413 );
    xnor g4947 ( n15672 , n24821 , n5706 );
    or g4948 ( n26474 , n14936 , n20423 );
    xnor g4949 ( n24148 , n2482 , n26149 );
    and g4950 ( n3102 , n11912 , n11421 );
    not g4951 ( n3540 , n26725 );
    or g4952 ( n24703 , n20173 , n7829 );
    and g4953 ( n16700 , n18922 , n4455 );
    nor g4954 ( n26325 , n14140 , n20822 );
    or g4955 ( n16691 , n4657 , n26617 );
    not g4956 ( n19433 , n19388 );
    and g4957 ( n673 , n11126 , n23906 );
    or g4958 ( n21301 , n12342 , n4811 );
    xnor g4959 ( n12390 , n16521 , n7139 );
    or g4960 ( n14329 , n1406 , n6502 );
    xnor g4961 ( n9208 , n19058 , n16439 );
    xnor g4962 ( n9835 , n4434 , n13453 );
    or g4963 ( n6984 , n2790 , n5517 );
    or g4964 ( n901 , n3490 , n666 );
    and g4965 ( n25152 , n13253 , n22276 );
    xnor g4966 ( n20557 , n16018 , n1435 );
    or g4967 ( n16796 , n5036 , n23882 );
    xnor g4968 ( n23289 , n21461 , n26169 );
    xnor g4969 ( n10854 , n22436 , n100 );
    xnor g4970 ( n25277 , n14719 , n24215 );
    xnor g4971 ( n3711 , n12626 , n4272 );
    or g4972 ( n1189 , n16712 , n17664 );
    xnor g4973 ( n4595 , n9338 , n4585 );
    or g4974 ( n24084 , n11312 , n2568 );
    not g4975 ( n25524 , n9832 );
    not g4976 ( n15433 , n17664 );
    or g4977 ( n23742 , n18710 , n15355 );
    nor g4978 ( n23818 , n8266 , n13495 );
    xnor g4979 ( n12179 , n10892 , n721 );
    not g4980 ( n22774 , n21763 );
    xnor g4981 ( n1620 , n22640 , n2013 );
    or g4982 ( n10784 , n12354 , n22392 );
    nor g4983 ( n15852 , n4964 , n8259 );
    or g4984 ( n12084 , n15084 , n21161 );
    nor g4985 ( n3013 , n26805 , n18404 );
    or g4986 ( n17357 , n10131 , n3690 );
    xnor g4987 ( n17299 , n3500 , n12905 );
    or g4988 ( n16063 , n20471 , n15308 );
    nor g4989 ( n19422 , n9605 , n11806 );
    nor g4990 ( n24844 , n15901 , n10220 );
    and g4991 ( n3553 , n21580 , n16229 );
    xnor g4992 ( n6630 , n16990 , n20480 );
    or g4993 ( n882 , n25094 , n3049 );
    xnor g4994 ( n5279 , n15153 , n9340 );
    xnor g4995 ( n18504 , n918 , n11356 );
    nor g4996 ( n9492 , n21606 , n26422 );
    not g4997 ( n16960 , n2316 );
    not g4998 ( n13577 , n11302 );
    or g4999 ( n19232 , n16101 , n8034 );
    or g5000 ( n13346 , n13561 , n12593 );
    not g5001 ( n22609 , n25196 );
    xnor g5002 ( n18653 , n16021 , n6550 );
    xnor g5003 ( n2112 , n3606 , n24643 );
    or g5004 ( n10536 , n12576 , n18563 );
    xnor g5005 ( n22498 , n26050 , n10372 );
    xnor g5006 ( n8906 , n23470 , n2021 );
    nor g5007 ( n2500 , n20923 , n11871 );
    xnor g5008 ( n1589 , n655 , n5386 );
    xnor g5009 ( n9990 , n23427 , n3795 );
    and g5010 ( n8599 , n535 , n2705 );
    xnor g5011 ( n11967 , n20972 , n1895 );
    not g5012 ( n24183 , n27100 );
    xnor g5013 ( n7079 , n24209 , n18339 );
    nor g5014 ( n22443 , n27099 , n24367 );
    not g5015 ( n24519 , n24886 );
    or g5016 ( n8978 , n4479 , n11986 );
    xnor g5017 ( n14691 , n7373 , n3480 );
    xnor g5018 ( n19208 , n7693 , n7566 );
    or g5019 ( n23376 , n15209 , n5952 );
    or g5020 ( n14328 , n8569 , n10791 );
    not g5021 ( n9114 , n26741 );
    xnor g5022 ( n25659 , n26446 , n12433 );
    or g5023 ( n1296 , n12238 , n11518 );
    nor g5024 ( n26918 , n12944 , n6864 );
    xnor g5025 ( n4129 , n1654 , n4256 );
    xnor g5026 ( n9467 , n1532 , n15058 );
    xnor g5027 ( n11267 , n9494 , n9227 );
    xnor g5028 ( n7514 , n13526 , n17713 );
    not g5029 ( n13152 , n3828 );
    not g5030 ( n1779 , n9151 );
    and g5031 ( n17474 , n11098 , n15175 );
    or g5032 ( n7120 , n26344 , n27146 );
    and g5033 ( n18484 , n3863 , n21204 );
    or g5034 ( n7965 , n10028 , n20682 );
    nor g5035 ( n8711 , n15114 , n25389 );
    xnor g5036 ( n25249 , n12241 , n3986 );
    and g5037 ( n25364 , n13127 , n1828 );
    nor g5038 ( n18954 , n23200 , n6122 );
    and g5039 ( n23802 , n4212 , n549 );
    and g5040 ( n22329 , n24638 , n12057 );
    nor g5041 ( n12603 , n3037 , n14385 );
    and g5042 ( n23426 , n3097 , n3764 );
    and g5043 ( n10231 , n14248 , n24108 );
    not g5044 ( n23724 , n1991 );
    and g5045 ( n12778 , n2914 , n13449 );
    xnor g5046 ( n17700 , n2894 , n12675 );
    or g5047 ( n23432 , n18028 , n1785 );
    or g5048 ( n7971 , n8099 , n17426 );
    xnor g5049 ( n16110 , n16363 , n19396 );
    xnor g5050 ( n21924 , n3102 , n16574 );
    or g5051 ( n4607 , n14369 , n4549 );
    not g5052 ( n13129 , n15142 );
    xnor g5053 ( n24992 , n14736 , n3529 );
    nor g5054 ( n8501 , n4715 , n16507 );
    not g5055 ( n15202 , n15979 );
    xnor g5056 ( n18193 , n19764 , n722 );
    not g5057 ( n24671 , n14637 );
    or g5058 ( n2959 , n22105 , n23277 );
    nor g5059 ( n14362 , n24351 , n12113 );
    or g5060 ( n7085 , n11413 , n15509 );
    or g5061 ( n24720 , n16881 , n4167 );
    or g5062 ( n17983 , n8948 , n14680 );
    not g5063 ( n23583 , n25609 );
    or g5064 ( n18732 , n12093 , n3535 );
    or g5065 ( n9850 , n11112 , n26817 );
    or g5066 ( n344 , n19754 , n11308 );
    not g5067 ( n9226 , n3623 );
    xnor g5068 ( n15558 , n9265 , n14355 );
    or g5069 ( n22839 , n10659 , n23126 );
    or g5070 ( n18946 , n19161 , n19254 );
    xnor g5071 ( n17689 , n14148 , n11503 );
    and g5072 ( n23868 , n17605 , n4263 );
    or g5073 ( n9292 , n23720 , n17186 );
    xnor g5074 ( n3901 , n25533 , n23854 );
    xnor g5075 ( n12479 , n18290 , n12875 );
    not g5076 ( n14268 , n10843 );
    nor g5077 ( n23953 , n19330 , n19703 );
    and g5078 ( n22519 , n16465 , n5449 );
    and g5079 ( n15973 , n23339 , n16950 );
    xnor g5080 ( n20084 , n22747 , n26438 );
    or g5081 ( n22229 , n11690 , n1914 );
    xnor g5082 ( n3872 , n23512 , n6341 );
    nor g5083 ( n21647 , n11441 , n7688 );
    or g5084 ( n21802 , n24791 , n2291 );
    nor g5085 ( n294 , n26334 , n8792 );
    nor g5086 ( n16995 , n6218 , n25464 );
    xnor g5087 ( n22909 , n24104 , n3344 );
    xnor g5088 ( n5607 , n4609 , n170 );
    xnor g5089 ( n22435 , n13471 , n15879 );
    and g5090 ( n23701 , n7259 , n2019 );
    xnor g5091 ( n3642 , n10396 , n7526 );
    nor g5092 ( n193 , n10274 , n8052 );
    xnor g5093 ( n22795 , n24663 , n26224 );
    or g5094 ( n15729 , n8713 , n54 );
    and g5095 ( n16282 , n13083 , n4131 );
    or g5096 ( n9301 , n12002 , n27102 );
    or g5097 ( n10185 , n15977 , n5638 );
    and g5098 ( n10695 , n8621 , n7760 );
    or g5099 ( n11345 , n16030 , n14916 );
    xnor g5100 ( n8065 , n5728 , n12265 );
    or g5101 ( n24713 , n15738 , n17490 );
    xnor g5102 ( n19842 , n11427 , n17972 );
    xnor g5103 ( n19358 , n15813 , n15671 );
    not g5104 ( n22110 , n800 );
    xnor g5105 ( n400 , n23701 , n23100 );
    xnor g5106 ( n7671 , n24163 , n7138 );
    nor g5107 ( n320 , n16937 , n16971 );
    not g5108 ( n1003 , n19372 );
    not g5109 ( n25838 , n8643 );
    xnor g5110 ( n7358 , n4436 , n13297 );
    or g5111 ( n14205 , n8367 , n5203 );
    xnor g5112 ( n2784 , n17301 , n27132 );
    xnor g5113 ( n17333 , n313 , n11463 );
    or g5114 ( n13804 , n446 , n21839 );
    xnor g5115 ( n3665 , n2634 , n4163 );
    xnor g5116 ( n15879 , n1662 , n20946 );
    and g5117 ( n24000 , n11455 , n14870 );
    and g5118 ( n16462 , n8568 , n1600 );
    xnor g5119 ( n16503 , n19646 , n19770 );
    xnor g5120 ( n1243 , n11119 , n26863 );
    not g5121 ( n2862 , n2355 );
    not g5122 ( n56 , n6478 );
    not g5123 ( n3138 , n5789 );
    or g5124 ( n2708 , n22724 , n24939 );
    not g5125 ( n5163 , n3445 );
    xnor g5126 ( n15635 , n17982 , n20986 );
    and g5127 ( n14703 , n21 , n23513 );
    xnor g5128 ( n6787 , n11006 , n23457 );
    not g5129 ( n24302 , n8371 );
    and g5130 ( n5712 , n25144 , n5972 );
    and g5131 ( n15657 , n1769 , n11076 );
    xnor g5132 ( n2173 , n18440 , n21914 );
    xnor g5133 ( n20761 , n22257 , n17859 );
    xnor g5134 ( n21013 , n7341 , n11254 );
    or g5135 ( n19831 , n9294 , n11351 );
    or g5136 ( n24922 , n26452 , n21025 );
    xnor g5137 ( n5493 , n16642 , n19630 );
    nor g5138 ( n8886 , n17854 , n23724 );
    not g5139 ( n5318 , n2184 );
    nor g5140 ( n15740 , n987 , n626 );
    or g5141 ( n2863 , n21021 , n18355 );
    xnor g5142 ( n1354 , n11121 , n19494 );
    and g5143 ( n7095 , n644 , n12868 );
    not g5144 ( n13435 , n21596 );
    xnor g5145 ( n6145 , n16476 , n15539 );
    xnor g5146 ( n26050 , n864 , n17684 );
    or g5147 ( n24547 , n20112 , n847 );
    xnor g5148 ( n23140 , n18341 , n19680 );
    and g5149 ( n6816 , n16784 , n15500 );
    and g5150 ( n21020 , n8872 , n17443 );
    xnor g5151 ( n15501 , n4636 , n6263 );
    xnor g5152 ( n10129 , n26946 , n978 );
    and g5153 ( n21177 , n8244 , n8431 );
    nor g5154 ( n17688 , n17536 , n19060 );
    or g5155 ( n24336 , n17949 , n22033 );
    or g5156 ( n14358 , n3836 , n4459 );
    xnor g5157 ( n12623 , n20429 , n12587 );
    nor g5158 ( n6448 , n17088 , n5241 );
    and g5159 ( n584 , n221 , n10523 );
    not g5160 ( n7281 , n690 );
    and g5161 ( n10203 , n24222 , n15091 );
    or g5162 ( n1745 , n4230 , n16290 );
    xnor g5163 ( n12203 , n1243 , n6698 );
    and g5164 ( n3721 , n13804 , n26759 );
    or g5165 ( n17691 , n16241 , n3885 );
    nor g5166 ( n12579 , n16924 , n8624 );
    and g5167 ( n1388 , n21351 , n20587 );
    xnor g5168 ( n7918 , n19392 , n18901 );
    xnor g5169 ( n25243 , n23286 , n13004 );
    not g5170 ( n17479 , n5579 );
    or g5171 ( n10575 , n13967 , n9788 );
    or g5172 ( n19447 , n20518 , n10922 );
    and g5173 ( n2487 , n14336 , n9349 );
    xnor g5174 ( n16445 , n21601 , n26776 );
    and g5175 ( n25563 , n4066 , n23439 );
    or g5176 ( n16564 , n1037 , n233 );
    and g5177 ( n8281 , n3734 , n14257 );
    or g5178 ( n15619 , n1508 , n23314 );
    and g5179 ( n19729 , n6075 , n23733 );
    or g5180 ( n11681 , n13016 , n13226 );
    nor g5181 ( n22730 , n19862 , n10155 );
    xnor g5182 ( n20824 , n12286 , n6525 );
    not g5183 ( n3403 , n2757 );
    or g5184 ( n23579 , n26904 , n10250 );
    xnor g5185 ( n15555 , n27030 , n15057 );
    xnor g5186 ( n12395 , n7098 , n7820 );
    buf g5187 ( n23002 , n11416 );
    and g5188 ( n9368 , n1278 , n19956 );
    or g5189 ( n23570 , n14816 , n12744 );
    or g5190 ( n15222 , n11454 , n19364 );
    xnor g5191 ( n22304 , n4108 , n18148 );
    or g5192 ( n24639 , n1181 , n14458 );
    or g5193 ( n1743 , n5165 , n12889 );
    xnor g5194 ( n170 , n23529 , n20700 );
    or g5195 ( n9013 , n20201 , n20231 );
    not g5196 ( n12763 , n23683 );
    not g5197 ( n12296 , n15047 );
    and g5198 ( n14552 , n12703 , n5959 );
    not g5199 ( n14545 , n5549 );
    xnor g5200 ( n13373 , n13853 , n18157 );
    and g5201 ( n6941 , n738 , n1920 );
    not g5202 ( n7983 , n18904 );
    xnor g5203 ( n14265 , n13977 , n20148 );
    or g5204 ( n4772 , n25886 , n2862 );
    or g5205 ( n19380 , n2038 , n2574 );
    not g5206 ( n9830 , n25918 );
    or g5207 ( n24287 , n15248 , n1014 );
    and g5208 ( n18550 , n18946 , n6322 );
    not g5209 ( n9679 , n8856 );
    and g5210 ( n19325 , n8269 , n21757 );
    xnor g5211 ( n14040 , n21872 , n3041 );
    not g5212 ( n25604 , n15867 );
    xnor g5213 ( n17746 , n1046 , n9213 );
    xnor g5214 ( n16249 , n25860 , n4961 );
    nor g5215 ( n14086 , n22247 , n19502 );
    or g5216 ( n5102 , n17226 , n2984 );
    and g5217 ( n11783 , n27159 , n19929 );
    or g5218 ( n9170 , n12593 , n13714 );
    and g5219 ( n24978 , n5025 , n23162 );
    not g5220 ( n8668 , n2664 );
    or g5221 ( n9517 , n13474 , n20462 );
    not g5222 ( n360 , n1842 );
    or g5223 ( n22199 , n12443 , n10664 );
    xnor g5224 ( n8773 , n8304 , n18771 );
    or g5225 ( n2822 , n18891 , n16364 );
    or g5226 ( n24780 , n2597 , n10682 );
    nor g5227 ( n12708 , n16092 , n2279 );
    xnor g5228 ( n8511 , n6570 , n25684 );
    and g5229 ( n7531 , n8311 , n8062 );
    and g5230 ( n7444 , n17598 , n17926 );
    xnor g5231 ( n15594 , n10092 , n12657 );
    nor g5232 ( n15895 , n15826 , n21585 );
    and g5233 ( n4987 , n8916 , n25473 );
    or g5234 ( n26020 , n17118 , n23730 );
    xnor g5235 ( n1121 , n17311 , n14172 );
    xnor g5236 ( n19087 , n25378 , n26630 );
    xnor g5237 ( n16360 , n26091 , n12667 );
    xnor g5238 ( n18337 , n4246 , n14511 );
    and g5239 ( n24254 , n4889 , n8263 );
    not g5240 ( n2645 , n21728 );
    xnor g5241 ( n13755 , n7587 , n18745 );
    and g5242 ( n13051 , n14915 , n22997 );
    and g5243 ( n23712 , n2549 , n3998 );
    xnor g5244 ( n8409 , n9200 , n2540 );
    and g5245 ( n26459 , n7146 , n3549 );
    nor g5246 ( n26551 , n4715 , n10117 );
    xnor g5247 ( n15176 , n18205 , n80 );
    or g5248 ( n15907 , n7742 , n11853 );
    or g5249 ( n2315 , n13858 , n5445 );
    nor g5250 ( n17373 , n19350 , n24331 );
    and g5251 ( n8336 , n537 , n21221 );
    not g5252 ( n10008 , n22335 );
    xnor g5253 ( n12436 , n23699 , n11844 );
    or g5254 ( n9131 , n12351 , n6503 );
    or g5255 ( n6613 , n14627 , n21259 );
    not g5256 ( n9095 , n23541 );
    not g5257 ( n7689 , n9888 );
    and g5258 ( n24572 , n15905 , n2510 );
    or g5259 ( n26277 , n19351 , n11863 );
    not g5260 ( n13071 , n2109 );
    or g5261 ( n6763 , n2500 , n11718 );
    nor g5262 ( n7681 , n13027 , n24929 );
    and g5263 ( n6440 , n23739 , n24498 );
    not g5264 ( n22783 , n82 );
    xnor g5265 ( n1113 , n26914 , n14620 );
    xnor g5266 ( n18152 , n7315 , n12705 );
    not g5267 ( n528 , n23842 );
    xnor g5268 ( n11467 , n10823 , n11194 );
    not g5269 ( n9683 , n10919 );
    and g5270 ( n12202 , n19361 , n20060 );
    or g5271 ( n15183 , n8525 , n4754 );
    xnor g5272 ( n21797 , n14365 , n25516 );
    xnor g5273 ( n20996 , n27200 , n2583 );
    nor g5274 ( n1959 , n10500 , n12493 );
    not g5275 ( n295 , n25252 );
    and g5276 ( n1824 , n5757 , n20818 );
    or g5277 ( n3520 , n6204 , n23254 );
    not g5278 ( n17867 , n5779 );
    nor g5279 ( n2563 , n2242 , n12810 );
    xnor g5280 ( n11658 , n23936 , n17620 );
    xnor g5281 ( n7231 , n2418 , n6303 );
    xnor g5282 ( n10362 , n21929 , n9575 );
    not g5283 ( n21460 , n21736 );
    xnor g5284 ( n12003 , n3427 , n24793 );
    xnor g5285 ( n4624 , n22245 , n9268 );
    xnor g5286 ( n6872 , n17604 , n25102 );
    or g5287 ( n10140 , n2272 , n26927 );
    xnor g5288 ( n21825 , n18978 , n25576 );
    xnor g5289 ( n2899 , n372 , n5085 );
    xnor g5290 ( n13176 , n18113 , n10557 );
    or g5291 ( n23449 , n12845 , n3623 );
    or g5292 ( n8463 , n2421 , n11243 );
    or g5293 ( n2464 , n26130 , n3661 );
    nor g5294 ( n10704 , n21693 , n15875 );
    xnor g5295 ( n18372 , n8455 , n13727 );
    not g5296 ( n9130 , n16240 );
    xnor g5297 ( n16675 , n7731 , n2328 );
    or g5298 ( n26773 , n12480 , n7318 );
    xnor g5299 ( n13199 , n18536 , n8577 );
    or g5300 ( n17290 , n21764 , n23900 );
    not g5301 ( n2812 , n2145 );
    not g5302 ( n9534 , n7340 );
    not g5303 ( n23807 , n8906 );
    xnor g5304 ( n3461 , n16547 , n19872 );
    xnor g5305 ( n7477 , n24137 , n18943 );
    xnor g5306 ( n1570 , n9246 , n7139 );
    or g5307 ( n19235 , n4545 , n1297 );
    not g5308 ( n10989 , n34 );
    not g5309 ( n22642 , n20374 );
    and g5310 ( n22065 , n21336 , n5536 );
    xnor g5311 ( n5117 , n24318 , n2013 );
    not g5312 ( n16002 , n6104 );
    or g5313 ( n20710 , n10971 , n17241 );
    and g5314 ( n3670 , n24245 , n3138 );
    xnor g5315 ( n2438 , n17035 , n2680 );
    or g5316 ( n19910 , n1565 , n1893 );
    nor g5317 ( n4359 , n22634 , n26942 );
    or g5318 ( n5281 , n17507 , n6277 );
    xnor g5319 ( n8834 , n16707 , n21749 );
    xnor g5320 ( n19932 , n10168 , n7267 );
    or g5321 ( n11531 , n11404 , n12804 );
    not g5322 ( n17061 , n14584 );
    xnor g5323 ( n26608 , n5538 , n20234 );
    or g5324 ( n2544 , n13618 , n2213 );
    or g5325 ( n2745 , n13734 , n6019 );
    and g5326 ( n1018 , n12301 , n26467 );
    xnor g5327 ( n22738 , n8499 , n17314 );
    or g5328 ( n11977 , n23133 , n23252 );
    nor g5329 ( n5968 , n22210 , n24496 );
    not g5330 ( n23616 , n25059 );
    nor g5331 ( n5553 , n14163 , n15512 );
    or g5332 ( n12378 , n10181 , n11056 );
    not g5333 ( n19159 , n12912 );
    xnor g5334 ( n8297 , n6538 , n9847 );
    xnor g5335 ( n7295 , n6079 , n26168 );
    xnor g5336 ( n6873 , n10903 , n4767 );
    nor g5337 ( n3865 , n12631 , n2867 );
    or g5338 ( n5322 , n7642 , n25907 );
    and g5339 ( n3420 , n14612 , n1400 );
    nor g5340 ( n22917 , n23187 , n20031 );
    nor g5341 ( n12407 , n6955 , n19390 );
    or g5342 ( n13876 , n25271 , n21649 );
    and g5343 ( n19438 , n23974 , n17013 );
    or g5344 ( n23547 , n4505 , n24757 );
    xnor g5345 ( n17147 , n4775 , n49 );
    nor g5346 ( n3813 , n12639 , n24091 );
    and g5347 ( n6473 , n892 , n10888 );
    xnor g5348 ( n4867 , n8446 , n21940 );
    xnor g5349 ( n1503 , n25063 , n11898 );
    and g5350 ( n15468 , n6146 , n4456 );
    or g5351 ( n8663 , n2640 , n3476 );
    and g5352 ( n20989 , n15891 , n9319 );
    or g5353 ( n21135 , n23896 , n11595 );
    and g5354 ( n17347 , n10117 , n19825 );
    nor g5355 ( n24755 , n12797 , n22327 );
    or g5356 ( n25686 , n951 , n7498 );
    xnor g5357 ( n7794 , n18436 , n13759 );
    xnor g5358 ( n461 , n14425 , n10638 );
    xnor g5359 ( n8988 , n11371 , n3370 );
    xnor g5360 ( n16218 , n16636 , n1114 );
    xnor g5361 ( n501 , n23482 , n3616 );
    not g5362 ( n19239 , n12281 );
    not g5363 ( n21974 , n1269 );
    nor g5364 ( n4852 , n2856 , n15798 );
    and g5365 ( n15752 , n6821 , n17527 );
    xnor g5366 ( n13141 , n14447 , n1604 );
    nor g5367 ( n5446 , n7837 , n1973 );
    and g5368 ( n5824 , n14853 , n5423 );
    and g5369 ( n1160 , n22937 , n1676 );
    nor g5370 ( n343 , n21747 , n26422 );
    not g5371 ( n209 , n10254 );
    or g5372 ( n3578 , n3936 , n16328 );
    not g5373 ( n26695 , n14684 );
    xnor g5374 ( n13501 , n23518 , n6902 );
    or g5375 ( n13149 , n26341 , n11204 );
    xnor g5376 ( n23565 , n6935 , n25194 );
    xnor g5377 ( n1837 , n5149 , n26024 );
    or g5378 ( n2016 , n356 , n1606 );
    xnor g5379 ( n2290 , n14680 , n5031 );
    xnor g5380 ( n26072 , n17379 , n12421 );
    and g5381 ( n10632 , n23160 , n13863 );
    or g5382 ( n18316 , n12880 , n16229 );
    or g5383 ( n24748 , n11011 , n10217 );
    xnor g5384 ( n4870 , n18948 , n5096 );
    xnor g5385 ( n25792 , n10879 , n12413 );
    or g5386 ( n1659 , n15748 , n21882 );
    or g5387 ( n21596 , n18893 , n2913 );
    and g5388 ( n23633 , n15069 , n20157 );
    xnor g5389 ( n17739 , n5565 , n20500 );
    and g5390 ( n9325 , n13263 , n22596 );
    or g5391 ( n6695 , n24590 , n20835 );
    xnor g5392 ( n23787 , n6711 , n2117 );
    nor g5393 ( n5638 , n25926 , n9646 );
    or g5394 ( n7522 , n14654 , n10577 );
    or g5395 ( n872 , n25088 , n5837 );
    xnor g5396 ( n15617 , n21580 , n18446 );
    or g5397 ( n22102 , n11733 , n14215 );
    or g5398 ( n3357 , n6416 , n9229 );
    xnor g5399 ( n19851 , n23076 , n17511 );
    not g5400 ( n25485 , n25547 );
    or g5401 ( n2118 , n21083 , n25974 );
    xnor g5402 ( n6819 , n12807 , n12966 );
    or g5403 ( n23841 , n16848 , n11356 );
    nor g5404 ( n16820 , n5905 , n8167 );
    or g5405 ( n16805 , n12553 , n14872 );
    not g5406 ( n15114 , n22290 );
    xnor g5407 ( n24745 , n24800 , n22463 );
    not g5408 ( n7183 , n2471 );
    and g5409 ( n26535 , n24583 , n9063 );
    and g5410 ( n3106 , n10526 , n14512 );
    or g5411 ( n14834 , n20836 , n13961 );
    and g5412 ( n23484 , n5400 , n3149 );
    or g5413 ( n9721 , n23237 , n9551 );
    not g5414 ( n14405 , n22885 );
    and g5415 ( n4924 , n16865 , n8470 );
    or g5416 ( n15838 , n26433 , n690 );
    and g5417 ( n3613 , n25286 , n9769 );
    or g5418 ( n12521 , n16573 , n1714 );
    and g5419 ( n16413 , n24006 , n25363 );
    and g5420 ( n3003 , n322 , n23934 );
    or g5421 ( n4681 , n17584 , n3425 );
    xnor g5422 ( n18024 , n18184 , n19572 );
    not g5423 ( n18770 , n6725 );
    nor g5424 ( n11880 , n12161 , n3072 );
    not g5425 ( n12212 , n8645 );
    and g5426 ( n11172 , n3837 , n12184 );
    and g5427 ( n26549 , n2170 , n9811 );
    or g5428 ( n4997 , n15577 , n13552 );
    nor g5429 ( n12307 , n12363 , n18468 );
    xnor g5430 ( n4404 , n7821 , n25128 );
    xnor g5431 ( n567 , n10016 , n2401 );
    or g5432 ( n5216 , n20371 , n8445 );
    xnor g5433 ( n2140 , n20937 , n424 );
    or g5434 ( n11106 , n25523 , n25455 );
    or g5435 ( n14338 , n619 , n14880 );
    and g5436 ( n13879 , n8867 , n18411 );
    or g5437 ( n15262 , n12961 , n2551 );
    and g5438 ( n7142 , n24311 , n17430 );
    xnor g5439 ( n15645 , n10710 , n9372 );
    xnor g5440 ( n5236 , n5438 , n13714 );
    or g5441 ( n2549 , n4941 , n9749 );
    not g5442 ( n3791 , n1662 );
    xnor g5443 ( n14819 , n9543 , n6480 );
    xnor g5444 ( n1927 , n8431 , n21547 );
    not g5445 ( n12453 , n7030 );
    or g5446 ( n14049 , n23489 , n20134 );
    or g5447 ( n24350 , n11523 , n6380 );
    and g5448 ( n9382 , n12565 , n9280 );
    and g5449 ( n16171 , n6978 , n6740 );
    xnor g5450 ( n24166 , n10320 , n3924 );
    xnor g5451 ( n3207 , n18797 , n24280 );
    xnor g5452 ( n1069 , n17821 , n2295 );
    and g5453 ( n2408 , n15331 , n18638 );
    xnor g5454 ( n19985 , n818 , n9942 );
    not g5455 ( n21891 , n4981 );
    not g5456 ( n24375 , n23923 );
    xnor g5457 ( n21144 , n20060 , n19361 );
    or g5458 ( n25411 , n15146 , n5532 );
    xnor g5459 ( n7172 , n5598 , n19728 );
    nor g5460 ( n6569 , n5266 , n3724 );
    or g5461 ( n2277 , n2056 , n14615 );
    xnor g5462 ( n26206 , n1803 , n5521 );
    xnor g5463 ( n20163 , n25972 , n10250 );
    nor g5464 ( n12443 , n10125 , n18326 );
    and g5465 ( n26723 , n12090 , n8487 );
    xnor g5466 ( n12304 , n21938 , n8072 );
    or g5467 ( n13996 , n25669 , n1453 );
    and g5468 ( n19847 , n16547 , n15 );
    or g5469 ( n6266 , n21994 , n20465 );
    or g5470 ( n16050 , n26230 , n19101 );
    or g5471 ( n1166 , n11246 , n14974 );
    and g5472 ( n21836 , n26034 , n13726 );
    not g5473 ( n25998 , n21522 );
    xnor g5474 ( n16354 , n6204 , n7674 );
    and g5475 ( n16899 , n895 , n5565 );
    xor g5476 ( n14655 , n6743 , n20385 );
    and g5477 ( n5999 , n26064 , n10930 );
    xnor g5478 ( n16327 , n26033 , n5126 );
    xnor g5479 ( n6098 , n12673 , n2300 );
    or g5480 ( n4437 , n3085 , n24747 );
    or g5481 ( n5757 , n17539 , n16524 );
    or g5482 ( n6952 , n12525 , n20928 );
    or g5483 ( n22672 , n1099 , n3379 );
    xnor g5484 ( n17371 , n7913 , n14090 );
    xnor g5485 ( n8455 , n7875 , n3063 );
    not g5486 ( n6267 , n12964 );
    or g5487 ( n18556 , n6206 , n9708 );
    or g5488 ( n20439 , n10438 , n23947 );
    xnor g5489 ( n12721 , n9615 , n19737 );
    and g5490 ( n18194 , n16754 , n9374 );
    xnor g5491 ( n23325 , n19218 , n14957 );
    or g5492 ( n13712 , n19588 , n19549 );
    or g5493 ( n13676 , n8743 , n11468 );
    or g5494 ( n18160 , n26891 , n8613 );
    xnor g5495 ( n13375 , n20271 , n10229 );
    or g5496 ( n27169 , n18992 , n7454 );
    or g5497 ( n4420 , n11938 , n3614 );
    and g5498 ( n6253 , n19429 , n14610 );
    xnor g5499 ( n5976 , n26218 , n3480 );
    xnor g5500 ( n25380 , n16117 , n8891 );
    and g5501 ( n20330 , n13918 , n20810 );
    and g5502 ( n10046 , n7631 , n2673 );
    and g5503 ( n5421 , n1713 , n14445 );
    or g5504 ( n25912 , n3601 , n22456 );
    and g5505 ( n18172 , n20700 , n26240 );
    xnor g5506 ( n7430 , n8211 , n16811 );
    not g5507 ( n1951 , n11893 );
    or g5508 ( n7443 , n26649 , n3980 );
    and g5509 ( n12183 , n14580 , n14195 );
    xnor g5510 ( n14045 , n15106 , n10508 );
    and g5511 ( n8786 , n22365 , n23122 );
    or g5512 ( n22837 , n2342 , n5213 );
    nor g5513 ( n5223 , n11736 , n10995 );
    not g5514 ( n13739 , n10875 );
    and g5515 ( n14447 , n21334 , n18399 );
    xnor g5516 ( n9391 , n24074 , n21969 );
    or g5517 ( n23195 , n18632 , n2608 );
    xnor g5518 ( n23779 , n2530 , n26572 );
    and g5519 ( n15522 , n16856 , n21081 );
    or g5520 ( n14673 , n14703 , n9221 );
    or g5521 ( n10621 , n9014 , n16208 );
    xnor g5522 ( n15834 , n11667 , n21398 );
    or g5523 ( n21574 , n8466 , n10082 );
    and g5524 ( n9815 , n11074 , n21872 );
    xnor g5525 ( n7996 , n8153 , n19355 );
    not g5526 ( n16848 , n2999 );
    nor g5527 ( n13283 , n12811 , n3260 );
    xnor g5528 ( n7534 , n1799 , n11580 );
    and g5529 ( n4372 , n5043 , n24726 );
    or g5530 ( n26257 , n25914 , n4941 );
    xnor g5531 ( n7233 , n26049 , n15642 );
    not g5532 ( n4780 , n11775 );
    xnor g5533 ( n22782 , n9037 , n23188 );
    nor g5534 ( n15223 , n12278 , n73 );
    or g5535 ( n549 , n7524 , n10314 );
    xnor g5536 ( n3641 , n10410 , n5493 );
    nor g5537 ( n17205 , n5006 , n9372 );
    nor g5538 ( n3231 , n20595 , n2322 );
    or g5539 ( n21655 , n23979 , n2690 );
    or g5540 ( n7690 , n6923 , n21647 );
    and g5541 ( n16831 , n21902 , n7154 );
    xnor g5542 ( n71 , n14486 , n16744 );
    xnor g5543 ( n1701 , n4805 , n25416 );
    xnor g5544 ( n23965 , n24617 , n6988 );
    not g5545 ( n24818 , n20092 );
    and g5546 ( n14292 , n14958 , n23822 );
    xnor g5547 ( n24875 , n13829 , n6145 );
    not g5548 ( n428 , n22122 );
    xnor g5549 ( n3247 , n22520 , n6974 );
    and g5550 ( n520 , n4678 , n17377 );
    xor g5551 ( n21354 , n17728 , n23586 );
    and g5552 ( n22936 , n8628 , n1035 );
    not g5553 ( n12076 , n19768 );
    or g5554 ( n19778 , n10839 , n22293 );
    or g5555 ( n24411 , n11745 , n6825 );
    xnor g5556 ( n2537 , n11620 , n17796 );
    or g5557 ( n3953 , n13389 , n20536 );
    and g5558 ( n3550 , n2247 , n19715 );
    xnor g5559 ( n12751 , n23376 , n19882 );
    xnor g5560 ( n17106 , n16300 , n5392 );
    or g5561 ( n10137 , n22743 , n4708 );
    xnor g5562 ( n24708 , n7693 , n19472 );
    or g5563 ( n25158 , n13417 , n23026 );
    not g5564 ( n10312 , n9314 );
    and g5565 ( n26143 , n2871 , n18376 );
    xnor g5566 ( n3669 , n25629 , n3795 );
    or g5567 ( n22081 , n23650 , n25115 );
    or g5568 ( n17181 , n14683 , n26010 );
    and g5569 ( n14024 , n23065 , n27055 );
    xnor g5570 ( n15867 , n16570 , n8214 );
    or g5571 ( n24053 , n19941 , n9345 );
    or g5572 ( n19574 , n24638 , n12057 );
    not g5573 ( n6126 , n17426 );
    not g5574 ( n20937 , n25772 );
    nor g5575 ( n19516 , n4409 , n25967 );
    xnor g5576 ( n5768 , n14116 , n12012 );
    or g5577 ( n2254 , n26452 , n2999 );
    not g5578 ( n21126 , n14782 );
    and g5579 ( n648 , n26063 , n14115 );
    or g5580 ( n26621 , n1293 , n15921 );
    and g5581 ( n11522 , n26725 , n17212 );
    xnor g5582 ( n11416 , n3093 , n25264 );
    and g5583 ( n4808 , n714 , n25357 );
    xnor g5584 ( n15783 , n24929 , n13027 );
    and g5585 ( n480 , n12979 , n986 );
    or g5586 ( n20807 , n5650 , n16360 );
    or g5587 ( n19771 , n15850 , n22206 );
    and g5588 ( n22975 , n11600 , n16843 );
    or g5589 ( n26000 , n2743 , n16312 );
    xnor g5590 ( n20278 , n2659 , n11926 );
    or g5591 ( n4604 , n13671 , n10275 );
    nor g5592 ( n27136 , n11152 , n21735 );
    not g5593 ( n15921 , n27193 );
    or g5594 ( n6331 , n22475 , n22794 );
    and g5595 ( n2739 , n8450 , n23042 );
    nor g5596 ( n23153 , n9096 , n25937 );
    or g5597 ( n7068 , n3878 , n20755 );
    xnor g5598 ( n23892 , n10153 , n15737 );
    not g5599 ( n9296 , n14761 );
    xnor g5600 ( n1227 , n5208 , n2387 );
    nor g5601 ( n22988 , n25581 , n1210 );
    xnor g5602 ( n26583 , n12669 , n10233 );
    xnor g5603 ( n15345 , n17668 , n6392 );
    xnor g5604 ( n20720 , n19061 , n9935 );
    nor g5605 ( n26411 , n19393 , n21508 );
    and g5606 ( n20408 , n11519 , n2681 );
    and g5607 ( n439 , n23621 , n23260 );
    and g5608 ( n13603 , n9136 , n7136 );
    or g5609 ( n15688 , n834 , n4106 );
    or g5610 ( n2681 , n27106 , n8264 );
    and g5611 ( n9768 , n7353 , n3830 );
    not g5612 ( n11756 , n12078 );
    or g5613 ( n26636 , n14495 , n25251 );
    and g5614 ( n4118 , n18681 , n12135 );
    not g5615 ( n23464 , n12417 );
    not g5616 ( n22436 , n17095 );
    and g5617 ( n14056 , n10522 , n19110 );
    not g5618 ( n7169 , n10980 );
    or g5619 ( n25804 , n19847 , n11878 );
    xnor g5620 ( n22016 , n5301 , n23319 );
    and g5621 ( n4663 , n16426 , n16774 );
    or g5622 ( n23286 , n13938 , n17489 );
    xnor g5623 ( n4552 , n19600 , n14278 );
    or g5624 ( n13009 , n1793 , n10702 );
    xnor g5625 ( n4898 , n27143 , n4371 );
    xnor g5626 ( n20044 , n8715 , n10611 );
    and g5627 ( n9424 , n3945 , n3393 );
    not g5628 ( n11186 , n2035 );
    and g5629 ( n11404 , n20323 , n11118 );
    or g5630 ( n8766 , n20425 , n12332 );
    xnor g5631 ( n17383 , n17408 , n4326 );
    xnor g5632 ( n21584 , n17397 , n5077 );
    xnor g5633 ( n26901 , n9251 , n22309 );
    xnor g5634 ( n20336 , n20244 , n27134 );
    xnor g5635 ( n6921 , n18451 , n13081 );
    or g5636 ( n7559 , n11725 , n14075 );
    xnor g5637 ( n7117 , n11597 , n17351 );
    and g5638 ( n14496 , n13453 , n4434 );
    not g5639 ( n13976 , n14584 );
    xnor g5640 ( n11197 , n26363 , n1553 );
    xnor g5641 ( n9851 , n10742 , n25245 );
    xnor g5642 ( n25739 , n1566 , n18711 );
    xnor g5643 ( n13113 , n10383 , n2690 );
    or g5644 ( n21284 , n13765 , n11540 );
    xnor g5645 ( n19955 , n24730 , n16277 );
    nor g5646 ( n4543 , n7817 , n11028 );
    not g5647 ( n13953 , n23076 );
    not g5648 ( n10485 , n2043 );
    xnor g5649 ( n24744 , n18651 , n25307 );
    xnor g5650 ( n24263 , n17567 , n18628 );
    and g5651 ( n23981 , n10117 , n22261 );
    and g5652 ( n24957 , n26164 , n24770 );
    nor g5653 ( n23687 , n13280 , n3136 );
    and g5654 ( n21056 , n318 , n23770 );
    xnor g5655 ( n12973 , n24759 , n17930 );
    and g5656 ( n10445 , n24185 , n12499 );
    xnor g5657 ( n27032 , n19446 , n17069 );
    or g5658 ( n1460 , n10683 , n10109 );
    xnor g5659 ( n15885 , n4680 , n7478 );
    xnor g5660 ( n16844 , n7071 , n428 );
    or g5661 ( n25695 , n18401 , n8289 );
    or g5662 ( n22590 , n12950 , n19210 );
    xnor g5663 ( n22934 , n22001 , n4519 );
    or g5664 ( n26199 , n21458 , n8891 );
    or g5665 ( n10290 , n22395 , n12991 );
    xnor g5666 ( n5414 , n26947 , n5231 );
    xnor g5667 ( n4060 , n26706 , n21143 );
    xnor g5668 ( n5471 , n26256 , n3261 );
    xnor g5669 ( n9129 , n15253 , n9984 );
    or g5670 ( n15687 , n21964 , n15961 );
    xnor g5671 ( n1104 , n26295 , n16896 );
    xnor g5672 ( n22317 , n13498 , n23240 );
    xnor g5673 ( n18877 , n18159 , n14716 );
    xnor g5674 ( n22771 , n20882 , n23685 );
    xnor g5675 ( n5780 , n10451 , n16034 );
    and g5676 ( n6165 , n9615 , n12774 );
    not g5677 ( n23791 , n18037 );
    or g5678 ( n10223 , n19371 , n18 );
    and g5679 ( n5461 , n7226 , n23727 );
    or g5680 ( n26910 , n20775 , n20808 );
    or g5681 ( n69 , n11133 , n430 );
    xnor g5682 ( n2370 , n14345 , n25381 );
    or g5683 ( n7549 , n8521 , n4652 );
    xnor g5684 ( n9498 , n23446 , n2623 );
    xnor g5685 ( n23517 , n23226 , n26150 );
    and g5686 ( n26985 , n15296 , n9478 );
    and g5687 ( n6057 , n16987 , n11807 );
    and g5688 ( n11776 , n17975 , n4202 );
    or g5689 ( n22132 , n6814 , n23463 );
    or g5690 ( n5713 , n22332 , n4104 );
    and g5691 ( n22092 , n8464 , n5248 );
    not g5692 ( n26413 , n7554 );
    and g5693 ( n4786 , n19844 , n12299 );
    xnor g5694 ( n1754 , n13846 , n15652 );
    or g5695 ( n13514 , n1997 , n11981 );
    xnor g5696 ( n16350 , n18082 , n23915 );
    or g5697 ( n3259 , n13237 , n14394 );
    and g5698 ( n22989 , n26074 , n19753 );
    or g5699 ( n929 , n2485 , n1625 );
    xnor g5700 ( n12470 , n634 , n4334 );
    or g5701 ( n12374 , n1077 , n18731 );
    and g5702 ( n19412 , n9907 , n18243 );
    nor g5703 ( n419 , n22557 , n1952 );
    or g5704 ( n10376 , n4368 , n17660 );
    or g5705 ( n7929 , n19258 , n9683 );
    xnor g5706 ( n5333 , n4108 , n11013 );
    or g5707 ( n25455 , n5579 , n26831 );
    and g5708 ( n1389 , n8358 , n24344 );
    and g5709 ( n2663 , n16261 , n23013 );
    xnor g5710 ( n4675 , n11320 , n11252 );
    and g5711 ( n11006 , n8442 , n249 );
    xnor g5712 ( n21628 , n12832 , n8238 );
    not g5713 ( n10464 , n2072 );
    or g5714 ( n14175 , n6382 , n25577 );
    xnor g5715 ( n15142 , n23961 , n7310 );
    nor g5716 ( n10227 , n25931 , n13053 );
    not g5717 ( n8230 , n3180 );
    or g5718 ( n13606 , n531 , n18769 );
    not g5719 ( n7316 , n23535 );
    or g5720 ( n18871 , n10452 , n25558 );
    not g5721 ( n17967 , n13518 );
    or g5722 ( n18951 , n2731 , n26879 );
    xnor g5723 ( n22789 , n11477 , n13915 );
    or g5724 ( n5630 , n18334 , n4433 );
    or g5725 ( n6472 , n13454 , n20789 );
    or g5726 ( n6045 , n17328 , n6947 );
    xnor g5727 ( n12705 , n10509 , n26417 );
    not g5728 ( n4195 , n4499 );
    and g5729 ( n15949 , n6474 , n16750 );
    nor g5730 ( n20383 , n2035 , n2675 );
    xnor g5731 ( n2602 , n22901 , n861 );
    xnor g5732 ( n12157 , n20063 , n15036 );
    xnor g5733 ( n17930 , n14733 , n19905 );
    xnor g5734 ( n23107 , n20127 , n23970 );
    or g5735 ( n16587 , n22943 , n24380 );
    and g5736 ( n19335 , n4496 , n5369 );
    xnor g5737 ( n17311 , n18249 , n26219 );
    not g5738 ( n9696 , n814 );
    or g5739 ( n21192 , n23940 , n18541 );
    not g5740 ( n26197 , n3228 );
    not g5741 ( n17960 , n9768 );
    xnor g5742 ( n16465 , n4578 , n10411 );
    xnor g5743 ( n21294 , n5105 , n14790 );
    not g5744 ( n23927 , n17914 );
    and g5745 ( n27202 , n20072 , n3639 );
    nor g5746 ( n8466 , n15077 , n6486 );
    nor g5747 ( n8323 , n5596 , n2340 );
    nor g5748 ( n11328 , n9244 , n10509 );
    and g5749 ( n14408 , n4469 , n23545 );
    xnor g5750 ( n14649 , n6057 , n10679 );
    nor g5751 ( n4654 , n14155 , n7339 );
    and g5752 ( n9846 , n14574 , n9092 );
    xnor g5753 ( n4978 , n6520 , n6837 );
    not g5754 ( n9018 , n22933 );
    not g5755 ( n13848 , n4712 );
    not g5756 ( n15713 , n18251 );
    nor g5757 ( n12178 , n5337 , n25228 );
    and g5758 ( n3000 , n2355 , n16223 );
    or g5759 ( n11097 , n24388 , n23927 );
    or g5760 ( n214 , n11191 , n4261 );
    xnor g5761 ( n941 , n11578 , n2261 );
    or g5762 ( n8012 , n4940 , n18409 );
    xnor g5763 ( n15111 , n20084 , n13117 );
    xnor g5764 ( n7568 , n5998 , n16078 );
    xnor g5765 ( n9509 , n8278 , n23166 );
    and g5766 ( n17501 , n20470 , n18634 );
    not g5767 ( n19529 , n3147 );
    xnor g5768 ( n20859 , n16458 , n8685 );
    xnor g5769 ( n723 , n19666 , n6148 );
    not g5770 ( n9789 , n21050 );
    xnor g5771 ( n8986 , n20358 , n3960 );
    not g5772 ( n7785 , n17305 );
    or g5773 ( n26633 , n16750 , n19828 );
    xnor g5774 ( n23659 , n25749 , n7377 );
    xnor g5775 ( n13463 , n4744 , n1999 );
    and g5776 ( n4416 , n15863 , n5239 );
    or g5777 ( n4303 , n743 , n20861 );
    nor g5778 ( n11339 , n690 , n25700 );
    or g5779 ( n4563 , n11294 , n24732 );
    xnor g5780 ( n10127 , n21749 , n26744 );
    nor g5781 ( n8498 , n22083 , n26499 );
    xnor g5782 ( n4695 , n5167 , n6773 );
    nor g5783 ( n18857 , n15767 , n19658 );
    nor g5784 ( n13857 , n14148 , n14275 );
    not g5785 ( n11143 , n632 );
    not g5786 ( n25101 , n16239 );
    nor g5787 ( n14404 , n5669 , n21575 );
    or g5788 ( n20041 , n14631 , n19769 );
    xnor g5789 ( n15793 , n13836 , n15065 );
    not g5790 ( n10622 , n22191 );
    xnor g5791 ( n7209 , n22197 , n16459 );
    not g5792 ( n23352 , n12445 );
    or g5793 ( n11931 , n9023 , n12307 );
    or g5794 ( n18938 , n25068 , n8324 );
    not g5795 ( n8522 , n19840 );
    xnor g5796 ( n16849 , n9789 , n19762 );
    xnor g5797 ( n1316 , n20151 , n17959 );
    or g5798 ( n3232 , n3018 , n9185 );
    and g5799 ( n19466 , n11694 , n18040 );
    or g5800 ( n11941 , n22776 , n18767 );
    nor g5801 ( n371 , n11736 , n2320 );
    nor g5802 ( n10944 , n7060 , n13821 );
    and g5803 ( n10887 , n12376 , n22967 );
    not g5804 ( n10181 , n20478 );
    xnor g5805 ( n8540 , n3881 , n3964 );
    not g5806 ( n189 , n24654 );
    and g5807 ( n18492 , n25169 , n15078 );
    not g5808 ( n4715 , n23250 );
    not g5809 ( n26447 , n25249 );
    or g5810 ( n25338 , n22745 , n10198 );
    xnor g5811 ( n21216 , n26895 , n12315 );
    xnor g5812 ( n1791 , n17793 , n24881 );
    xnor g5813 ( n12314 , n23913 , n16376 );
    xnor g5814 ( n5387 , n950 , n22789 );
    xnor g5815 ( n9314 , n473 , n6430 );
    or g5816 ( n4187 , n3542 , n2014 );
    xnor g5817 ( n23637 , n4668 , n18373 );
    xnor g5818 ( n5424 , n18739 , n3911 );
    xnor g5819 ( n20441 , n2953 , n10996 );
    and g5820 ( n4289 , n3294 , n14177 );
    not g5821 ( n10446 , n10383 );
    xnor g5822 ( n26232 , n4719 , n23582 );
    and g5823 ( n4754 , n14034 , n24546 );
    nor g5824 ( n10192 , n401 , n3030 );
    and g5825 ( n5250 , n9352 , n6269 );
    or g5826 ( n2241 , n8851 , n15212 );
    and g5827 ( n15473 , n22254 , n22699 );
    xnor g5828 ( n10508 , n14130 , n12861 );
    xnor g5829 ( n23505 , n16738 , n12860 );
    or g5830 ( n6557 , n16351 , n2721 );
    or g5831 ( n136 , n3199 , n3373 );
    xnor g5832 ( n18664 , n13185 , n1450 );
    nor g5833 ( n25876 , n13154 , n15891 );
    xnor g5834 ( n27145 , n6197 , n2149 );
    and g5835 ( n13961 , n17890 , n6009 );
    or g5836 ( n20650 , n26417 , n11482 );
    and g5837 ( n9223 , n19161 , n22405 );
    and g5838 ( n3542 , n13171 , n13633 );
    and g5839 ( n11940 , n15021 , n11663 );
    nor g5840 ( n2495 , n16443 , n13166 );
    not g5841 ( n3752 , n12274 );
    and g5842 ( n23418 , n20367 , n13630 );
    and g5843 ( n8652 , n20878 , n13024 );
    not g5844 ( n7242 , n21860 );
    or g5845 ( n1412 , n9854 , n14955 );
    xnor g5846 ( n732 , n15534 , n25572 );
    nor g5847 ( n10190 , n14750 , n12470 );
    and g5848 ( n12174 , n15416 , n13554 );
    or g5849 ( n16598 , n13353 , n12317 );
    xnor g5850 ( n10224 , n13811 , n18454 );
    xnor g5851 ( n1586 , n12456 , n5404 );
    xnor g5852 ( n1169 , n15546 , n24937 );
    and g5853 ( n26731 , n4119 , n9310 );
    xnor g5854 ( n5093 , n13303 , n12546 );
    and g5855 ( n25842 , n21711 , n9630 );
    or g5856 ( n24395 , n11111 , n286 );
    xnor g5857 ( n8884 , n23112 , n20443 );
    not g5858 ( n26201 , n12502 );
    xnor g5859 ( n26641 , n19415 , n15874 );
    or g5860 ( n14242 , n21649 , n17846 );
    nor g5861 ( n20581 , n2481 , n23201 );
    and g5862 ( n18199 , n23376 , n26108 );
    not g5863 ( n8935 , n18002 );
    xnor g5864 ( n14125 , n3501 , n6152 );
    or g5865 ( n21389 , n5329 , n2694 );
    xnor g5866 ( n20268 , n19911 , n14570 );
    nor g5867 ( n5849 , n15182 , n21915 );
    or g5868 ( n1333 , n10997 , n16486 );
    and g5869 ( n8035 , n9517 , n18015 );
    xnor g5870 ( n15353 , n6598 , n14063 );
    xnor g5871 ( n23319 , n5238 , n9456 );
    and g5872 ( n9929 , n8852 , n7888 );
    xnor g5873 ( n27130 , n8478 , n7905 );
    nor g5874 ( n24282 , n8292 , n5916 );
    not g5875 ( n17414 , n13089 );
    or g5876 ( n13692 , n3423 , n21065 );
    nor g5877 ( n10719 , n25505 , n23843 );
    xnor g5878 ( n19058 , n26182 , n12314 );
    xnor g5879 ( n3459 , n20769 , n4756 );
    or g5880 ( n16888 , n9003 , n11876 );
    and g5881 ( n19819 , n22141 , n6886 );
    not g5882 ( n22614 , n2958 );
    xnor g5883 ( n25574 , n14557 , n16249 );
    or g5884 ( n9063 , n23848 , n26792 );
    not g5885 ( n24750 , n7186 );
    or g5886 ( n26702 , n12572 , n8063 );
    xnor g5887 ( n11206 , n9096 , n6127 );
    or g5888 ( n14744 , n940 , n25787 );
    not g5889 ( n744 , n4588 );
    or g5890 ( n14540 , n21937 , n7953 );
    or g5891 ( n8384 , n15894 , n7329 );
    not g5892 ( n23271 , n2111 );
    or g5893 ( n20305 , n8680 , n11192 );
    and g5894 ( n16908 , n4287 , n1670 );
    or g5895 ( n8086 , n16896 , n781 );
    nor g5896 ( n898 , n8875 , n18655 );
    not g5897 ( n13693 , n16886 );
    not g5898 ( n7709 , n25808 );
    not g5899 ( n12110 , n26135 );
    not g5900 ( n18158 , n15996 );
    or g5901 ( n6008 , n4676 , n8980 );
    and g5902 ( n2137 , n11455 , n9940 );
    or g5903 ( n22777 , n6843 , n14871 );
    not g5904 ( n23018 , n16696 );
    or g5905 ( n18423 , n14818 , n16631 );
    not g5906 ( n18404 , n21948 );
    or g5907 ( n19654 , n3807 , n12536 );
    xnor g5908 ( n15280 , n5196 , n1878 );
    and g5909 ( n6766 , n21557 , n14485 );
    xnor g5910 ( n12913 , n19170 , n3608 );
    xnor g5911 ( n10679 , n9142 , n26565 );
    not g5912 ( n14774 , n16077 );
    or g5913 ( n5141 , n13590 , n13783 );
    and g5914 ( n11440 , n2377 , n12246 );
    xnor g5915 ( n23247 , n1538 , n8523 );
    xnor g5916 ( n6527 , n20151 , n20429 );
    not g5917 ( n5244 , n20415 );
    xnor g5918 ( n2705 , n841 , n13718 );
    and g5919 ( n2335 , n13330 , n7182 );
    and g5920 ( n2267 , n4568 , n14023 );
    not g5921 ( n8430 , n25043 );
    and g5922 ( n26920 , n8569 , n10791 );
    nor g5923 ( n10958 , n14718 , n468 );
    or g5924 ( n16010 , n24684 , n12880 );
    and g5925 ( n3205 , n21507 , n14037 );
    or g5926 ( n26108 , n5330 , n1386 );
    not g5927 ( n19719 , n19230 );
    or g5928 ( n4698 , n1009 , n152 );
    not g5929 ( n16778 , n8374 );
    not g5930 ( n5709 , n13069 );
    or g5931 ( n14030 , n4081 , n21810 );
    not g5932 ( n26782 , n25926 );
    xnor g5933 ( n447 , n14033 , n22797 );
    nor g5934 ( n13637 , n5211 , n12811 );
    or g5935 ( n12602 , n15796 , n23095 );
    and g5936 ( n23024 , n23837 , n7137 );
    not g5937 ( n22289 , n7716 );
    xnor g5938 ( n6349 , n6043 , n4764 );
    nor g5939 ( n12760 , n25749 , n7377 );
    or g5940 ( n7510 , n21942 , n16908 );
    xnor g5941 ( n4760 , n25993 , n3421 );
    and g5942 ( n12532 , n13382 , n13068 );
    nor g5943 ( n16209 , n25038 , n23745 );
    nor g5944 ( n8334 , n10712 , n26512 );
    not g5945 ( n2738 , n12029 );
    or g5946 ( n10325 , n3190 , n23141 );
    or g5947 ( n16416 , n13753 , n16792 );
    nor g5948 ( n20894 , n10650 , n22253 );
    or g5949 ( n11890 , n1360 , n24257 );
    or g5950 ( n4945 , n24000 , n21215 );
    not g5951 ( n16513 , n23661 );
    xnor g5952 ( n9145 , n25917 , n3959 );
    or g5953 ( n7826 , n21744 , n1900 );
    xnor g5954 ( n18059 , n25579 , n21032 );
    or g5955 ( n15853 , n15629 , n18614 );
    nor g5956 ( n17055 , n24358 , n20951 );
    and g5957 ( n18963 , n16494 , n5486 );
    and g5958 ( n6382 , n23486 , n11734 );
    xnor g5959 ( n27046 , n26575 , n11284 );
    and g5960 ( n5567 , n528 , n13627 );
    not g5961 ( n8153 , n24151 );
    not g5962 ( n2399 , n3524 );
    xnor g5963 ( n8600 , n10562 , n4632 );
    xnor g5964 ( n18876 , n12968 , n16244 );
    not g5965 ( n19667 , n12626 );
    and g5966 ( n10553 , n444 , n8142 );
    and g5967 ( n24423 , n8007 , n4244 );
    xnor g5968 ( n16793 , n12441 , n19379 );
    or g5969 ( n10955 , n21375 , n16109 );
    xnor g5970 ( n7708 , n7011 , n11395 );
    xnor g5971 ( n4847 , n19152 , n23842 );
    or g5972 ( n9101 , n9260 , n10093 );
    or g5973 ( n14813 , n16609 , n22666 );
    xnor g5974 ( n7221 , n11406 , n15929 );
    or g5975 ( n23665 , n20206 , n6105 );
    or g5976 ( n3427 , n4073 , n17566 );
    and g5977 ( n22951 , n12862 , n14503 );
    xnor g5978 ( n6141 , n7446 , n9691 );
    xnor g5979 ( n21125 , n11114 , n14345 );
    or g5980 ( n7853 , n22323 , n24405 );
    xnor g5981 ( n4614 , n9167 , n14656 );
    and g5982 ( n7273 , n26112 , n19207 );
    or g5983 ( n22617 , n19200 , n26803 );
    or g5984 ( n20873 , n16179 , n11164 );
    xnor g5985 ( n19674 , n5010 , n22481 );
    and g5986 ( n4167 , n2441 , n806 );
    nor g5987 ( n10840 , n20754 , n593 );
    xnor g5988 ( n13626 , n14834 , n24265 );
    not g5989 ( n17599 , n21206 );
    and g5990 ( n10043 , n18742 , n14319 );
    xnor g5991 ( n5485 , n4433 , n22508 );
    and g5992 ( n1944 , n21217 , n697 );
    or g5993 ( n10747 , n13166 , n22340 );
    and g5994 ( n13632 , n10900 , n10087 );
    xnor g5995 ( n10342 , n23582 , n16738 );
    xnor g5996 ( n1773 , n19812 , n23652 );
    not g5997 ( n4603 , n22476 );
    and g5998 ( n22995 , n7266 , n17533 );
    and g5999 ( n25500 , n14654 , n12664 );
    xnor g6000 ( n4626 , n25699 , n22290 );
    or g6001 ( n15320 , n2022 , n1903 );
    nor g6002 ( n24285 , n13405 , n22253 );
    nor g6003 ( n18704 , n9741 , n11229 );
    not g6004 ( n20338 , n11936 );
    not g6005 ( n14288 , n8694 );
    xnor g6006 ( n18416 , n5525 , n25694 );
    or g6007 ( n26070 , n20321 , n3861 );
    xnor g6008 ( n11295 , n26368 , n19118 );
    not g6009 ( n4342 , n4957 );
    xnor g6010 ( n1049 , n12967 , n5028 );
    not g6011 ( n7882 , n13685 );
    xnor g6012 ( n1505 , n16845 , n3228 );
    or g6013 ( n9277 , n706 , n7771 );
    or g6014 ( n11460 , n5611 , n25694 );
    and g6015 ( n15413 , n23598 , n23604 );
    and g6016 ( n886 , n21526 , n18732 );
    xnor g6017 ( n2688 , n14524 , n16223 );
    and g6018 ( n24863 , n12004 , n12289 );
    not g6019 ( n9244 , n2418 );
    or g6020 ( n1462 , n6356 , n4665 );
    or g6021 ( n18890 , n7606 , n25092 );
    nor g6022 ( n23641 , n2049 , n9303 );
    xnor g6023 ( n5453 , n7788 , n20013 );
    and g6024 ( n7613 , n13773 , n10778 );
    xnor g6025 ( n10330 , n20195 , n15336 );
    not g6026 ( n12198 , n13578 );
    nor g6027 ( n13223 , n4714 , n5030 );
    not g6028 ( n2815 , n11416 );
    not g6029 ( n8720 , n1592 );
    xnor g6030 ( n23232 , n15842 , n9665 );
    and g6031 ( n21713 , n4620 , n26591 );
    not g6032 ( n3124 , n9557 );
    xnor g6033 ( n15746 , n4792 , n10593 );
    xnor g6034 ( n14720 , n19086 , n18307 );
    not g6035 ( n18665 , n3488 );
    or g6036 ( n8880 , n14654 , n26797 );
    and g6037 ( n18873 , n26612 , n21139 );
    not g6038 ( n15519 , n5832 );
    or g6039 ( n1286 , n9800 , n8905 );
    xnor g6040 ( n12325 , n24970 , n24913 );
    or g6041 ( n785 , n10100 , n22898 );
    not g6042 ( n25929 , n13695 );
    or g6043 ( n3717 , n4520 , n10699 );
    nor g6044 ( n21350 , n13459 , n24786 );
    or g6045 ( n18917 , n1619 , n11684 );
    nor g6046 ( n18471 , n1204 , n25701 );
    xnor g6047 ( n17359 , n3417 , n8934 );
    xnor g6048 ( n22471 , n11302 , n24786 );
    or g6049 ( n24490 , n1458 , n1642 );
    or g6050 ( n2632 , n12929 , n10691 );
    and g6051 ( n21495 , n19282 , n23709 );
    nor g6052 ( n19476 , n12507 , n15739 );
    not g6053 ( n5355 , n25565 );
    nor g6054 ( n5204 , n2453 , n20700 );
    or g6055 ( n3283 , n20213 , n26725 );
    and g6056 ( n23070 , n17416 , n1529 );
    or g6057 ( n15156 , n24355 , n13951 );
    and g6058 ( n15231 , n14759 , n24668 );
    xnor g6059 ( n6148 , n10527 , n3314 );
    or g6060 ( n23116 , n12945 , n19160 );
    not g6061 ( n11393 , n7057 );
    or g6062 ( n17876 , n11147 , n12981 );
    or g6063 ( n22242 , n10123 , n15557 );
    xnor g6064 ( n12001 , n3186 , n5834 );
    not g6065 ( n21935 , n10107 );
    nor g6066 ( n3216 , n8186 , n19282 );
    and g6067 ( n14658 , n24071 , n22900 );
    and g6068 ( n24410 , n4780 , n21922 );
    not g6069 ( n25888 , n20470 );
    xnor g6070 ( n1278 , n8596 , n24732 );
    or g6071 ( n16857 , n24691 , n10336 );
    and g6072 ( n20001 , n23403 , n13880 );
    and g6073 ( n13585 , n22694 , n15183 );
    xnor g6074 ( n17810 , n7072 , n6857 );
    not g6075 ( n7111 , n24937 );
    or g6076 ( n11157 , n6259 , n24152 );
    not g6077 ( n3635 , n643 );
    not g6078 ( n7532 , n24875 );
    and g6079 ( n11448 , n9066 , n22894 );
    and g6080 ( n14343 , n9953 , n4946 );
    xnor g6081 ( n10625 , n5975 , n21675 );
    xnor g6082 ( n2363 , n12016 , n11162 );
    not g6083 ( n9564 , n11974 );
    nor g6084 ( n15251 , n9259 , n12423 );
    and g6085 ( n5988 , n20599 , n16450 );
    or g6086 ( n6792 , n19593 , n7227 );
    xor g6087 ( n17408 , n9014 , n11567 );
    or g6088 ( n4823 , n15284 , n26819 );
    or g6089 ( n775 , n3022 , n7188 );
    and g6090 ( n4025 , n4054 , n14820 );
    xnor g6091 ( n11877 , n26881 , n26651 );
    xnor g6092 ( n5049 , n18477 , n10629 );
    or g6093 ( n17240 , n8315 , n26460 );
    xnor g6094 ( n26298 , n234 , n2755 );
    xnor g6095 ( n2306 , n2331 , n12546 );
    xnor g6096 ( n15765 , n3480 , n7057 );
    xnor g6097 ( n1513 , n758 , n14731 );
    xnor g6098 ( n12607 , n7772 , n2827 );
    and g6099 ( n5389 , n6485 , n26265 );
    and g6100 ( n25613 , n12989 , n23470 );
    or g6101 ( n7084 , n15884 , n26001 );
    xnor g6102 ( n18953 , n18622 , n25893 );
    xnor g6103 ( n26425 , n1184 , n16657 );
    or g6104 ( n13619 , n5796 , n1869 );
    not g6105 ( n20444 , n22225 );
    or g6106 ( n5538 , n2633 , n14058 );
    or g6107 ( n22299 , n23769 , n13747 );
    or g6108 ( n5654 , n14415 , n5822 );
    or g6109 ( n3342 , n18550 , n22259 );
    or g6110 ( n11886 , n18471 , n17706 );
    nor g6111 ( n16286 , n24948 , n11322 );
    or g6112 ( n23157 , n18078 , n10711 );
    xnor g6113 ( n19904 , n12200 , n13215 );
    not g6114 ( n570 , n11841 );
    xnor g6115 ( n5902 , n17536 , n23799 );
    and g6116 ( n12009 , n1314 , n20967 );
    xnor g6117 ( n256 , n20020 , n20145 );
    and g6118 ( n19958 , n1988 , n2687 );
    and g6119 ( n27138 , n9715 , n24527 );
    or g6120 ( n16815 , n22515 , n10467 );
    nor g6121 ( n11808 , n5620 , n23814 );
    xnor g6122 ( n11611 , n17161 , n8282 );
    or g6123 ( n13369 , n2175 , n15384 );
    not g6124 ( n9802 , n20349 );
    nor g6125 ( n1352 , n20169 , n4426 );
    not g6126 ( n1838 , n8732 );
    or g6127 ( n13187 , n1348 , n9784 );
    or g6128 ( n7247 , n13156 , n21321 );
    or g6129 ( n22979 , n6569 , n6989 );
    xnor g6130 ( n25430 , n10275 , n22359 );
    or g6131 ( n222 , n22 , n9674 );
    not g6132 ( n1715 , n7339 );
    not g6133 ( n25715 , n10650 );
    nor g6134 ( n22601 , n11056 , n21276 );
    xnor g6135 ( n19071 , n26629 , n19904 );
    xnor g6136 ( n4231 , n5658 , n21682 );
    xnor g6137 ( n13170 , n19271 , n14045 );
    xnor g6138 ( n7885 , n8964 , n22554 );
    and g6139 ( n17686 , n25997 , n24349 );
    and g6140 ( n2655 , n4291 , n10823 );
    and g6141 ( n13589 , n26199 , n14594 );
    and g6142 ( n19305 , n17759 , n16391 );
    or g6143 ( n27080 , n21317 , n8251 );
    or g6144 ( n17892 , n19962 , n1570 );
    or g6145 ( n18637 , n18786 , n25953 );
    xnor g6146 ( n12088 , n8683 , n15379 );
    not g6147 ( n23013 , n15158 );
    xnor g6148 ( n13045 , n15482 , n5123 );
    nor g6149 ( n19461 , n12535 , n15167 );
    not g6150 ( n9496 , n20754 );
    xnor g6151 ( n16422 , n485 , n4642 );
    and g6152 ( n5458 , n11727 , n25292 );
    and g6153 ( n15744 , n25258 , n6838 );
    not g6154 ( n6255 , n13623 );
    or g6155 ( n25350 , n15116 , n15821 );
    nor g6156 ( n24876 , n3740 , n12232 );
    xnor g6157 ( n12585 , n1558 , n3918 );
    nor g6158 ( n22637 , n11976 , n11437 );
    not g6159 ( n10151 , n1895 );
    not g6160 ( n25099 , n5376 );
    xnor g6161 ( n10843 , n20368 , n6741 );
    and g6162 ( n6947 , n7782 , n10688 );
    or g6163 ( n3224 , n5531 , n22952 );
    or g6164 ( n7770 , n11542 , n3136 );
    not g6165 ( n6025 , n16752 );
    and g6166 ( n23627 , n23068 , n13171 );
    xnor g6167 ( n1712 , n2633 , n5341 );
    or g6168 ( n1688 , n7311 , n5657 );
    xnor g6169 ( n2382 , n15227 , n2794 );
    xnor g6170 ( n19334 , n9399 , n6502 );
    xnor g6171 ( n21658 , n23097 , n6082 );
    xnor g6172 ( n15728 , n16387 , n3673 );
    xnor g6173 ( n22841 , n7771 , n6885 );
    xnor g6174 ( n21645 , n6976 , n10035 );
    nor g6175 ( n13049 , n23631 , n3365 );
    not g6176 ( n17002 , n2328 );
    or g6177 ( n6482 , n14979 , n19106 );
    xnor g6178 ( n25321 , n8819 , n16961 );
    xnor g6179 ( n16013 , n10569 , n5275 );
    not g6180 ( n10086 , n13518 );
    and g6181 ( n9362 , n10933 , n326 );
    or g6182 ( n4536 , n10205 , n2538 );
    and g6183 ( n4304 , n10285 , n471 );
    and g6184 ( n19316 , n21042 , n13512 );
    or g6185 ( n17910 , n6051 , n11302 );
    xnor g6186 ( n23253 , n4705 , n919 );
    xnor g6187 ( n7958 , n19377 , n23784 );
    and g6188 ( n1184 , n5945 , n7067 );
    and g6189 ( n8172 , n16238 , n22334 );
    xnor g6190 ( n2232 , n7092 , n20213 );
    and g6191 ( n184 , n25055 , n4079 );
    xnor g6192 ( n2472 , n17035 , n19515 );
    and g6193 ( n1122 , n21310 , n18620 );
    not g6194 ( n3780 , n7636 );
    not g6195 ( n25376 , n18452 );
    and g6196 ( n24169 , n26388 , n702 );
    not g6197 ( n22549 , n16165 );
    not g6198 ( n9788 , n16274 );
    not g6199 ( n9242 , n4259 );
    and g6200 ( n1486 , n14711 , n20204 );
    and g6201 ( n1564 , n4932 , n19969 );
    and g6202 ( n11757 , n26540 , n8102 );
    and g6203 ( n13177 , n19106 , n8715 );
    xnor g6204 ( n19284 , n20885 , n10537 );
    not g6205 ( n17832 , n3671 );
    not g6206 ( n24806 , n24948 );
    or g6207 ( n6091 , n8679 , n8379 );
    nor g6208 ( n14369 , n7670 , n10485 );
    xnor g6209 ( n3581 , n13981 , n6611 );
    and g6210 ( n23497 , n21813 , n10133 );
    or g6211 ( n25123 , n2415 , n172 );
    or g6212 ( n1650 , n11014 , n23900 );
    or g6213 ( n22195 , n23380 , n17008 );
    xnor g6214 ( n7132 , n7059 , n6202 );
    not g6215 ( n15085 , n23636 );
    xnor g6216 ( n4684 , n9993 , n22201 );
    xnor g6217 ( n17218 , n15773 , n21997 );
    nor g6218 ( n23328 , n16376 , n17467 );
    xnor g6219 ( n2792 , n21381 , n11507 );
    xnor g6220 ( n4855 , n7640 , n17511 );
    xnor g6221 ( n9243 , n21822 , n25617 );
    and g6222 ( n3169 , n7982 , n8907 );
    or g6223 ( n5620 , n6297 , n21587 );
    xnor g6224 ( n433 , n6200 , n12288 );
    and g6225 ( n3308 , n18601 , n19874 );
    nor g6226 ( n12544 , n20235 , n8259 );
    or g6227 ( n10678 , n25444 , n6461 );
    or g6228 ( n18824 , n12130 , n14894 );
    xnor g6229 ( n7083 , n21922 , n14217 );
    xnor g6230 ( n20356 , n14754 , n17366 );
    or g6231 ( n4910 , n9821 , n11838 );
    or g6232 ( n21106 , n15492 , n14478 );
    xnor g6233 ( n19467 , n16967 , n3080 );
    and g6234 ( n5839 , n19901 , n8486 );
    not g6235 ( n14719 , n15378 );
    xnor g6236 ( n25635 , n12650 , n16544 );
    and g6237 ( n1453 , n23682 , n8404 );
    xnor g6238 ( n781 , n4763 , n22304 );
    xnor g6239 ( n2004 , n12549 , n23790 );
    xnor g6240 ( n11969 , n16642 , n964 );
    and g6241 ( n8018 , n15905 , n14996 );
    or g6242 ( n12542 , n10463 , n2647 );
    and g6243 ( n24409 , n21819 , n26737 );
    xnor g6244 ( n26177 , n12662 , n11720 );
    and g6245 ( n13680 , n16436 , n25849 );
    or g6246 ( n24449 , n26231 , n11174 );
    not g6247 ( n21127 , n27134 );
    xnor g6248 ( n6716 , n22613 , n18157 );
    or g6249 ( n22966 , n10036 , n14360 );
    xnor g6250 ( n23388 , n27193 , n1293 );
    and g6251 ( n1367 , n19299 , n4779 );
    and g6252 ( n1782 , n15123 , n23017 );
    xor g6253 ( n2350 , n5462 , n14679 );
    xnor g6254 ( n16758 , n14923 , n7238 );
    or g6255 ( n1613 , n23486 , n11734 );
    not g6256 ( n3714 , n12567 );
    not g6257 ( n13828 , n21501 );
    not g6258 ( n14566 , n5451 );
    xor g6259 ( n20692 , n20425 , n3053 );
    or g6260 ( n19262 , n20259 , n3925 );
    nor g6261 ( n25334 , n12789 , n23180 );
    xnor g6262 ( n5336 , n5905 , n8167 );
    or g6263 ( n404 , n18562 , n18195 );
    or g6264 ( n16708 , n24744 , n14557 );
    not g6265 ( n834 , n4943 );
    xnor g6266 ( n466 , n15062 , n12457 );
    and g6267 ( n14462 , n3446 , n3267 );
    xnor g6268 ( n16837 , n20779 , n24910 );
    not g6269 ( n5611 , n12398 );
    not g6270 ( n8818 , n24312 );
    xnor g6271 ( n7435 , n22181 , n4284 );
    nor g6272 ( n613 , n13152 , n167 );
    or g6273 ( n8093 , n16286 , n13041 );
    not g6274 ( n1236 , n25296 );
    xnor g6275 ( n17544 , n16731 , n26191 );
    xnor g6276 ( n16550 , n18907 , n26823 );
    xnor g6277 ( n9269 , n4979 , n9702 );
    and g6278 ( n21881 , n10030 , n4557 );
    or g6279 ( n17045 , n23974 , n281 );
    nor g6280 ( n1246 , n9920 , n13650 );
    or g6281 ( n13415 , n18394 , n26453 );
    or g6282 ( n9205 , n7666 , n4914 );
    nor g6283 ( n14966 , n21721 , n7466 );
    xnor g6284 ( n12538 , n11924 , n10986 );
    or g6285 ( n21592 , n6904 , n26241 );
    not g6286 ( n112 , n21905 );
    or g6287 ( n19035 , n25674 , n19634 );
    or g6288 ( n8799 , n15743 , n20658 );
    xnor g6289 ( n5609 , n2772 , n21131 );
    nor g6290 ( n13635 , n9700 , n15482 );
    xor g6291 ( n19979 , n9961 , n8589 );
    or g6292 ( n14077 , n13461 , n5746 );
    xnor g6293 ( n6612 , n23468 , n7231 );
    and g6294 ( n3371 , n1509 , n16913 );
    xnor g6295 ( n879 , n25343 , n19261 );
    xnor g6296 ( n5961 , n22031 , n4923 );
    nor g6297 ( n14 , n12522 , n12208 );
    not g6298 ( n13278 , n24704 );
    or g6299 ( n21196 , n5895 , n21817 );
    not g6300 ( n8232 , n3179 );
    and g6301 ( n17809 , n5014 , n18579 );
    and g6302 ( n24783 , n21857 , n10861 );
    not g6303 ( n1199 , n10231 );
    or g6304 ( n1647 , n6478 , n4375 );
    xnor g6305 ( n18271 , n1186 , n26408 );
    and g6306 ( n11318 , n9535 , n11846 );
    or g6307 ( n12215 , n11184 , n6842 );
    or g6308 ( n8026 , n25617 , n13448 );
    or g6309 ( n8169 , n20502 , n19977 );
    or g6310 ( n22171 , n4542 , n8805 );
    xnor g6311 ( n10478 , n5213 , n3468 );
    or g6312 ( n21285 , n27186 , n15194 );
    xnor g6313 ( n25337 , n5774 , n5040 );
    or g6314 ( n18851 , n25370 , n11603 );
    not g6315 ( n6143 , n9450 );
    nor g6316 ( n9007 , n2420 , n23807 );
    xnor g6317 ( n18794 , n18021 , n9486 );
    or g6318 ( n5854 , n23250 , n11209 );
    or g6319 ( n15157 , n13677 , n10451 );
    xnor g6320 ( n629 , n24727 , n7882 );
    not g6321 ( n20053 , n19138 );
    and g6322 ( n1567 , n26305 , n3657 );
    and g6323 ( n18382 , n4862 , n25902 );
    or g6324 ( n13627 , n8344 , n21804 );
    not g6325 ( n3591 , n1773 );
    and g6326 ( n3123 , n18602 , n20992 );
    xnor g6327 ( n14375 , n14188 , n4331 );
    nor g6328 ( n14406 , n26797 , n15077 );
    or g6329 ( n23324 , n26088 , n939 );
    or g6330 ( n14672 , n23234 , n1688 );
    or g6331 ( n25281 , n18321 , n20238 );
    xnor g6332 ( n6586 , n5862 , n18841 );
    and g6333 ( n22445 , n22332 , n22370 );
    or g6334 ( n5623 , n800 , n25547 );
    xnor g6335 ( n1521 , n1672 , n14244 );
    or g6336 ( n24223 , n264 , n20344 );
    xnor g6337 ( n23593 , n4665 , n18558 );
    xnor g6338 ( n15614 , n19870 , n6495 );
    xnor g6339 ( n7607 , n7513 , n20431 );
    and g6340 ( n15215 , n9520 , n26376 );
    xnor g6341 ( n20377 , n8227 , n11947 );
    nor g6342 ( n3113 , n8161 , n6870 );
    xnor g6343 ( n693 , n23569 , n13139 );
    nor g6344 ( n18321 , n16642 , n704 );
    xnor g6345 ( n19523 , n21103 , n629 );
    xnor g6346 ( n15892 , n22553 , n7891 );
    and g6347 ( n14517 , n932 , n10739 );
    xnor g6348 ( n16733 , n1298 , n2148 );
    xnor g6349 ( n4513 , n26005 , n2742 );
    xnor g6350 ( n9635 , n11866 , n21356 );
    xnor g6351 ( n16162 , n7934 , n5608 );
    or g6352 ( n14403 , n8340 , n4580 );
    and g6353 ( n16739 , n411 , n22650 );
    or g6354 ( n9071 , n6782 , n10498 );
    and g6355 ( n8959 , n1268 , n23953 );
    xnor g6356 ( n21849 , n25159 , n24056 );
    or g6357 ( n24553 , n19171 , n24293 );
    and g6358 ( n545 , n3349 , n2919 );
    not g6359 ( n17276 , n14811 );
    not g6360 ( n21261 , n15135 );
    or g6361 ( n13087 , n11685 , n21226 );
    xnor g6362 ( n21927 , n7115 , n3987 );
    or g6363 ( n9224 , n12500 , n20930 );
    and g6364 ( n15854 , n26660 , n26810 );
    or g6365 ( n13974 , n19543 , n4618 );
    nor g6366 ( n9119 , n17287 , n23697 );
    xnor g6367 ( n11017 , n7023 , n5942 );
    xnor g6368 ( n9135 , n18766 , n12186 );
    nor g6369 ( n13080 , n26516 , n16052 );
    xnor g6370 ( n10698 , n12017 , n15807 );
    not g6371 ( n12762 , n25355 );
    or g6372 ( n8458 , n15395 , n15203 );
    nor g6373 ( n1058 , n24301 , n4256 );
    nor g6374 ( n19732 , n27175 , n7056 );
    or g6375 ( n25299 , n23436 , n3276 );
    nor g6376 ( n6330 , n6768 , n20412 );
    xnor g6377 ( n17392 , n1732 , n16887 );
    and g6378 ( n2375 , n9329 , n11528 );
    or g6379 ( n11361 , n2629 , n25124 );
    nor g6380 ( n16046 , n25838 , n26935 );
    and g6381 ( n23896 , n9393 , n24233 );
    xnor g6382 ( n23270 , n2397 , n4554 );
    and g6383 ( n24474 , n27196 , n10393 );
    xnor g6384 ( n11548 , n17191 , n16104 );
    not g6385 ( n818 , n13946 );
    xnor g6386 ( n26838 , n6154 , n23829 );
    or g6387 ( n15613 , n2557 , n8441 );
    or g6388 ( n23611 , n12493 , n16520 );
    not g6389 ( n7258 , n1351 );
    nor g6390 ( n26309 , n24937 , n12436 );
    and g6391 ( n25579 , n660 , n22368 );
    xnor g6392 ( n6791 , n10457 , n11746 );
    xnor g6393 ( n11470 , n9189 , n14857 );
    and g6394 ( n14321 , n19124 , n26381 );
    or g6395 ( n13065 , n4579 , n511 );
    and g6396 ( n23812 , n20640 , n13149 );
    not g6397 ( n5947 , n3504 );
    not g6398 ( n8378 , n20755 );
    or g6399 ( n12589 , n12319 , n24745 );
    nor g6400 ( n10243 , n20770 , n10468 );
    xnor g6401 ( n9901 , n11583 , n13538 );
    xnor g6402 ( n7928 , n2246 , n3668 );
    nor g6403 ( n23413 , n14957 , n19218 );
    not g6404 ( n15065 , n27117 );
    not g6405 ( n8037 , n27202 );
    xnor g6406 ( n7695 , n26892 , n11623 );
    not g6407 ( n2941 , n26253 );
    not g6408 ( n5264 , n12142 );
    or g6409 ( n5821 , n18221 , n16090 );
    or g6410 ( n19553 , n17026 , n3078 );
    xnor g6411 ( n20767 , n93 , n3515 );
    xnor g6412 ( n15749 , n10434 , n3728 );
    or g6413 ( n18029 , n14576 , n25069 );
    xnor g6414 ( n13718 , n4322 , n16029 );
    or g6415 ( n22641 , n18758 , n12407 );
    xnor g6416 ( n7968 , n9299 , n17518 );
    or g6417 ( n2870 , n10533 , n24117 );
    or g6418 ( n15821 , n24549 , n26477 );
    not g6419 ( n26122 , n9215 );
    and g6420 ( n3600 , n13815 , n7449 );
    nor g6421 ( n27048 , n25277 , n21860 );
    and g6422 ( n11529 , n11175 , n18968 );
    and g6423 ( n12560 , n11093 , n26400 );
    not g6424 ( n9665 , n12606 );
    and g6425 ( n2564 , n6104 , n2056 );
    nor g6426 ( n16049 , n420 , n7365 );
    and g6427 ( n11964 , n6206 , n17409 );
    xnor g6428 ( n22472 , n26843 , n18935 );
    xnor g6429 ( n11433 , n16524 , n3785 );
    or g6430 ( n6231 , n16111 , n9219 );
    xnor g6431 ( n3027 , n5445 , n21759 );
    not g6432 ( n21795 , n21599 );
    and g6433 ( n15611 , n8014 , n26446 );
    xnor g6434 ( n1810 , n20075 , n15891 );
    or g6435 ( n10507 , n6554 , n25060 );
    or g6436 ( n14938 , n8370 , n6909 );
    xnor g6437 ( n18674 , n25035 , n16317 );
    or g6438 ( n18009 , n16922 , n1486 );
    xnor g6439 ( n23323 , n9768 , n16321 );
    or g6440 ( n17604 , n25395 , n17648 );
    nor g6441 ( n10038 , n7621 , n2510 );
    and g6442 ( n2634 , n17079 , n16556 );
    xnor g6443 ( n22282 , n90 , n22044 );
    and g6444 ( n743 , n13190 , n15769 );
    xnor g6445 ( n2162 , n4469 , n23545 );
    xnor g6446 ( n26822 , n20825 , n17842 );
    or g6447 ( n19635 , n26325 , n8892 );
    and g6448 ( n6737 , n22446 , n24467 );
    or g6449 ( n140 , n23168 , n8067 );
    or g6450 ( n11907 , n23638 , n16271 );
    xnor g6451 ( n12874 , n24774 , n22660 );
    nor g6452 ( n9650 , n18331 , n1415 );
    and g6453 ( n2587 , n15549 , n22813 );
    and g6454 ( n211 , n2682 , n5577 );
    and g6455 ( n479 , n22168 , n5334 );
    nor g6456 ( n15331 , n5640 , n3674 );
    xnor g6457 ( n10345 , n319 , n8226 );
    nor g6458 ( n8749 , n17911 , n22207 );
    or g6459 ( n12559 , n22029 , n10173 );
    xnor g6460 ( n22714 , n16245 , n21275 );
    xnor g6461 ( n15630 , n20883 , n5859 );
    and g6462 ( n13299 , n17491 , n11977 );
    or g6463 ( n16569 , n17423 , n14584 );
    or g6464 ( n10703 , n22791 , n27064 );
    nor g6465 ( n9958 , n15767 , n18973 );
    or g6466 ( n23028 , n23555 , n11745 );
    not g6467 ( n9456 , n26193 );
    or g6468 ( n26839 , n12788 , n15808 );
    xnor g6469 ( n25556 , n12354 , n24323 );
    nor g6470 ( n16320 , n10312 , n10013 );
    or g6471 ( n15735 , n5849 , n2956 );
    or g6472 ( n9304 , n12348 , n22603 );
    and g6473 ( n5983 , n9475 , n22827 );
    or g6474 ( n1892 , n12702 , n348 );
    nor g6475 ( n4657 , n658 , n22274 );
    not g6476 ( n5284 , n3307 );
    not g6477 ( n10406 , n8881 );
    or g6478 ( n2527 , n10207 , n20084 );
    nor g6479 ( n5484 , n1844 , n54 );
    xnor g6480 ( n6341 , n7156 , n10710 );
    or g6481 ( n20047 , n8658 , n6158 );
    not g6482 ( n3050 , n23207 );
    and g6483 ( n17109 , n20844 , n9059 );
    xnor g6484 ( n3147 , n1614 , n2771 );
    or g6485 ( n10164 , n22176 , n7676 );
    not g6486 ( n10431 , n11210 );
    xnor g6487 ( n17705 , n9083 , n21132 );
    nor g6488 ( n20659 , n16994 , n4964 );
    not g6489 ( n13945 , n26585 );
    and g6490 ( n21793 , n5686 , n11773 );
    and g6491 ( n23243 , n4453 , n12542 );
    nor g6492 ( n17981 , n19652 , n17444 );
    and g6493 ( n20763 , n16610 , n4793 );
    xnor g6494 ( n2560 , n27000 , n7181 );
    or g6495 ( n9982 , n15984 , n26521 );
    nor g6496 ( n20071 , n302 , n11975 );
    xnor g6497 ( n4253 , n11056 , n21276 );
    not g6498 ( n14730 , n20153 );
    and g6499 ( n12503 , n14965 , n25465 );
    or g6500 ( n3210 , n2087 , n17986 );
    or g6501 ( n23949 , n15760 , n23285 );
    xnor g6502 ( n6037 , n1886 , n10096 );
    xnor g6503 ( n135 , n4400 , n2651 );
    xnor g6504 ( n577 , n2509 , n22289 );
    not g6505 ( n16878 , n9632 );
    xnor g6506 ( n20754 , n16691 , n476 );
    not g6507 ( n19442 , n19745 );
    or g6508 ( n2687 , n10816 , n23130 );
    nor g6509 ( n21607 , n15389 , n24468 );
    buf g6510 ( n6510 , n4259 );
    xnor g6511 ( n20073 , n19215 , n395 );
    not g6512 ( n7676 , n23065 );
    and g6513 ( n11693 , n17677 , n17242 );
    or g6514 ( n9450 , n22274 , n24129 );
    and g6515 ( n2949 , n6122 , n1894 );
    or g6516 ( n15829 , n11273 , n7949 );
    xnor g6517 ( n20835 , n14221 , n345 );
    or g6518 ( n17905 , n13386 , n22305 );
    not g6519 ( n13561 , n11503 );
    and g6520 ( n1886 , n15427 , n19201 );
    xnor g6521 ( n13740 , n12837 , n6068 );
    or g6522 ( n14663 , n11189 , n25666 );
    and g6523 ( n19997 , n7889 , n17941 );
    not g6524 ( n24273 , n7270 );
    not g6525 ( n2579 , n23430 );
    nor g6526 ( n9438 , n1834 , n3354 );
    xnor g6527 ( n13186 , n23241 , n24563 );
    and g6528 ( n19109 , n23030 , n4333 );
    and g6529 ( n368 , n21863 , n756 );
    or g6530 ( n20931 , n10452 , n3785 );
    xnor g6531 ( n16346 , n9854 , n3056 );
    or g6532 ( n11532 , n17957 , n30 );
    or g6533 ( n3919 , n11747 , n5648 );
    and g6534 ( n9673 , n4338 , n25106 );
    nor g6535 ( n24752 , n12014 , n7215 );
    not g6536 ( n5917 , n8160 );
    and g6537 ( n12100 , n17399 , n16124 );
    nor g6538 ( n26155 , n9254 , n25657 );
    and g6539 ( n156 , n14452 , n21490 );
    or g6540 ( n12729 , n24810 , n15898 );
    and g6541 ( n13700 , n1788 , n16112 );
    and g6542 ( n19532 , n14837 , n18093 );
    xnor g6543 ( n17256 , n17230 , n21687 );
    xnor g6544 ( n14902 , n6163 , n17829 );
    or g6545 ( n17595 , n25004 , n18409 );
    xnor g6546 ( n11040 , n13569 , n4964 );
    not g6547 ( n15101 , n6178 );
    xnor g6548 ( n1371 , n2844 , n20073 );
    xnor g6549 ( n7881 , n18869 , n13073 );
    xnor g6550 ( n23181 , n993 , n26479 );
    or g6551 ( n11807 , n16634 , n12308 );
    xnor g6552 ( n20970 , n9669 , n20946 );
    or g6553 ( n9698 , n19709 , n9806 );
    xnor g6554 ( n15970 , n25026 , n8669 );
    and g6555 ( n11930 , n26559 , n24354 );
    xnor g6556 ( n10422 , n219 , n13450 );
    and g6557 ( n10663 , n1678 , n6409 );
    and g6558 ( n11222 , n20123 , n5909 );
    and g6559 ( n13061 , n3480 , n7373 );
    nor g6560 ( n5650 , n4869 , n15024 );
    xnor g6561 ( n9474 , n839 , n15709 );
    and g6562 ( n8715 , n9570 , n3637 );
    not g6563 ( n18174 , n19595 );
    or g6564 ( n18795 , n6238 , n14664 );
    nor g6565 ( n1957 , n11118 , n15442 );
    nor g6566 ( n20454 , n14056 , n8915 );
    or g6567 ( n17895 , n5304 , n15437 );
    nor g6568 ( n1140 , n16336 , n16306 );
    or g6569 ( n418 , n16924 , n22395 );
    nor g6570 ( n3162 , n10758 , n14845 );
    nor g6571 ( n11624 , n7284 , n7750 );
    or g6572 ( n23038 , n23745 , n23053 );
    nor g6573 ( n2970 , n8497 , n26914 );
    and g6574 ( n23926 , n20010 , n26368 );
    and g6575 ( n26091 , n26807 , n17677 );
    xnor g6576 ( n15051 , n19556 , n3483 );
    and g6577 ( n18829 , n1757 , n11970 );
    not g6578 ( n260 , n17345 );
    not g6579 ( n7798 , n24847 );
    or g6580 ( n12114 , n12967 , n11030 );
    xnor g6581 ( n21477 , n10053 , n19911 );
    xnor g6582 ( n7596 , n3468 , n23430 );
    xnor g6583 ( n3429 , n5442 , n19752 );
    xnor g6584 ( n26953 , n16396 , n22871 );
    or g6585 ( n13664 , n26095 , n12939 );
    and g6586 ( n23241 , n4772 , n25833 );
    not g6587 ( n4217 , n17553 );
    nor g6588 ( n9044 , n4917 , n23905 );
    not g6589 ( n17987 , n14788 );
    or g6590 ( n10104 , n15795 , n18606 );
    nor g6591 ( n20264 , n5999 , n17762 );
    nor g6592 ( n3503 , n7254 , n14071 );
    or g6593 ( n21351 , n10096 , n26553 );
    xnor g6594 ( n8934 , n24949 , n23681 );
    or g6595 ( n14877 , n4776 , n17420 );
    or g6596 ( n9393 , n3958 , n10746 );
    xnor g6597 ( n5682 , n10445 , n1253 );
    xnor g6598 ( n2904 , n3570 , n8067 );
    nor g6599 ( n15832 , n822 , n12869 );
    and g6600 ( n5477 , n15855 , n11511 );
    or g6601 ( n21990 , n12189 , n542 );
    xnor g6602 ( n23307 , n21147 , n25869 );
    and g6603 ( n15374 , n11857 , n149 );
    or g6604 ( n15441 , n2236 , n754 );
    not g6605 ( n23144 , n3710 );
    xnor g6606 ( n1961 , n22274 , n11192 );
    nor g6607 ( n13184 , n20314 , n10253 );
    not g6608 ( n26974 , n23985 );
    and g6609 ( n20335 , n11561 , n3732 );
    and g6610 ( n6824 , n15454 , n26039 );
    and g6611 ( n15194 , n1134 , n3876 );
    or g6612 ( n6052 , n3479 , n11937 );
    xor g6613 ( n17863 , n16468 , n7674 );
    or g6614 ( n25265 , n21495 , n23255 );
    xnor g6615 ( n21642 , n2782 , n5793 );
    or g6616 ( n25720 , n5602 , n19179 );
    and g6617 ( n14359 , n2108 , n1641 );
    nor g6618 ( n6704 , n2355 , n115 );
    nor g6619 ( n22244 , n14387 , n15007 );
    nor g6620 ( n8332 , n3351 , n9842 );
    or g6621 ( n25421 , n15041 , n13224 );
    nor g6622 ( n23320 , n13033 , n19392 );
    or g6623 ( n10379 , n21636 , n22154 );
    and g6624 ( n12784 , n17250 , n26997 );
    xnor g6625 ( n2920 , n19368 , n5802 );
    xnor g6626 ( n8861 , n3852 , n2431 );
    and g6627 ( n18723 , n19428 , n21553 );
    and g6628 ( n9831 , n25516 , n16242 );
    nor g6629 ( n14515 , n15693 , n24701 );
    not g6630 ( n26892 , n15801 );
    not g6631 ( n10131 , n15602 );
    and g6632 ( n16723 , n1642 , n5512 );
    or g6633 ( n4832 , n5957 , n19997 );
    xnor g6634 ( n8807 , n12143 , n20215 );
    or g6635 ( n18779 , n1864 , n11835 );
    or g6636 ( n4593 , n18444 , n26224 );
    nor g6637 ( n16922 , n20641 , n3443 );
    xnor g6638 ( n11281 , n1533 , n5451 );
    not g6639 ( n23751 , n2352 );
    xnor g6640 ( n14456 , n16213 , n14878 );
    nor g6641 ( n20416 , n146 , n2979 );
    or g6642 ( n20357 , n19949 , n16474 );
    xnor g6643 ( n22584 , n19034 , n26282 );
    and g6644 ( n17695 , n6833 , n2040 );
    xnor g6645 ( n3829 , n5628 , n2054 );
    nor g6646 ( n8208 , n21634 , n5579 );
    and g6647 ( n3942 , n12002 , n11382 );
    not g6648 ( n13745 , n8315 );
    or g6649 ( n27159 , n2117 , n6711 );
    xnor g6650 ( n13297 , n16409 , n23861 );
    xnor g6651 ( n26035 , n27089 , n6814 );
    or g6652 ( n17907 , n19205 , n11068 );
    or g6653 ( n16706 , n17763 , n12908 );
    xnor g6654 ( n12094 , n17266 , n25239 );
    or g6655 ( n26183 , n14193 , n16172 );
    or g6656 ( n9354 , n10982 , n21560 );
    and g6657 ( n18081 , n24107 , n14291 );
    xnor g6658 ( n5091 , n22426 , n20658 );
    or g6659 ( n25046 , n11283 , n23128 );
    or g6660 ( n22165 , n13770 , n12491 );
    or g6661 ( n11917 , n2514 , n5213 );
    not g6662 ( n13919 , n21047 );
    xnor g6663 ( n9423 , n22046 , n24268 );
    and g6664 ( n18688 , n15990 , n2977 );
    not g6665 ( n25799 , n11489 );
    and g6666 ( n7865 , n9947 , n22726 );
    and g6667 ( n20863 , n23838 , n24204 );
    and g6668 ( n24072 , n20314 , n147 );
    and g6669 ( n6765 , n3931 , n11596 );
    or g6670 ( n127 , n10413 , n21881 );
    xnor g6671 ( n1939 , n19473 , n24372 );
    xnor g6672 ( n3516 , n12010 , n10624 );
    or g6673 ( n24445 , n12478 , n3917 );
    xor g6674 ( n14610 , n11022 , n6890 );
    and g6675 ( n9649 , n8983 , n21737 );
    xnor g6676 ( n14444 , n9965 , n26665 );
    not g6677 ( n1753 , n21911 );
    nor g6678 ( n1783 , n12 , n23725 );
    and g6679 ( n19417 , n5932 , n5359 );
    xnor g6680 ( n10732 , n16107 , n6068 );
    not g6681 ( n9479 , n2743 );
    or g6682 ( n20034 , n25313 , n1212 );
    nor g6683 ( n15452 , n17302 , n13784 );
    or g6684 ( n1197 , n22426 , n20620 );
    or g6685 ( n3156 , n26925 , n10199 );
    not g6686 ( n20139 , n10072 );
    xnor g6687 ( n12983 , n17090 , n27120 );
    and g6688 ( n24023 , n9472 , n7611 );
    or g6689 ( n11272 , n20113 , n23930 );
    or g6690 ( n17443 , n12651 , n24779 );
    and g6691 ( n2302 , n26706 , n19872 );
    and g6692 ( n18660 , n6604 , n24871 );
    nor g6693 ( n22954 , n14507 , n18058 );
    xnor g6694 ( n23009 , n19713 , n10820 );
    not g6695 ( n11151 , n20231 );
    and g6696 ( n15104 , n17711 , n8398 );
    and g6697 ( n11982 , n17879 , n15771 );
    and g6698 ( n25743 , n6561 , n19386 );
    xnor g6699 ( n15926 , n8358 , n26189 );
    xnor g6700 ( n21662 , n25926 , n12384 );
    or g6701 ( n408 , n7797 , n8925 );
    not g6702 ( n14226 , n12861 );
    xnor g6703 ( n26113 , n9786 , n22217 );
    or g6704 ( n19665 , n10436 , n16148 );
    or g6705 ( n3382 , n3216 , n20591 );
    not g6706 ( n20112 , n24327 );
    xnor g6707 ( n10214 , n3337 , n26552 );
    and g6708 ( n26283 , n8424 , n26432 );
    or g6709 ( n17341 , n14566 , n20378 );
    and g6710 ( n14449 , n1494 , n7120 );
    or g6711 ( n18348 , n19563 , n15045 );
    not g6712 ( n16459 , n21164 );
    or g6713 ( n9624 , n20152 , n13192 );
    nor g6714 ( n2142 , n25156 , n2152 );
    and g6715 ( n24982 , n19676 , n8812 );
    xnor g6716 ( n500 , n5675 , n1876 );
    and g6717 ( n5915 , n13205 , n120 );
    or g6718 ( n20258 , n19094 , n19156 );
    or g6719 ( n22193 , n15527 , n3894 );
    and g6720 ( n19921 , n19938 , n11623 );
    nor g6721 ( n9853 , n5436 , n9972 );
    and g6722 ( n3852 , n15540 , n23031 );
    or g6723 ( n13797 , n13280 , n13309 );
    or g6724 ( n21059 , n14040 , n24711 );
    nor g6725 ( n1979 , n21622 , n15158 );
    or g6726 ( n10429 , n4338 , n25106 );
    xnor g6727 ( n19238 , n15166 , n20377 );
    or g6728 ( n4932 , n18797 , n11489 );
    and g6729 ( n20225 , n4994 , n6447 );
    xnor g6730 ( n3947 , n25120 , n17458 );
    xnor g6731 ( n14488 , n21064 , n16397 );
    or g6732 ( n13516 , n26997 , n17250 );
    xnor g6733 ( n21900 , n5889 , n6914 );
    or g6734 ( n23049 , n19469 , n6209 );
    and g6735 ( n16119 , n16649 , n6493 );
    or g6736 ( n12159 , n15454 , n23892 );
    and g6737 ( n11255 , n1814 , n5080 );
    not g6738 ( n24705 , n8079 );
    xnor g6739 ( n19935 , n25048 , n22815 );
    xnor g6740 ( n7716 , n13088 , n18987 );
    and g6741 ( n8011 , n7042 , n14159 );
    xnor g6742 ( n16451 , n19297 , n21248 );
    or g6743 ( n13787 , n26093 , n20235 );
    or g6744 ( n8844 , n20138 , n9251 );
    xnor g6745 ( n833 , n16911 , n7773 );
    and g6746 ( n2601 , n23756 , n23194 );
    nor g6747 ( n10120 , n26053 , n2320 );
    xnor g6748 ( n13350 , n17978 , n3134 );
    xnor g6749 ( n1658 , n24567 , n4366 );
    nor g6750 ( n3293 , n4194 , n14643 );
    nor g6751 ( n3499 , n10155 , n1738 );
    xnor g6752 ( n24898 , n6176 , n20849 );
    not g6753 ( n22671 , n4202 );
    xor g6754 ( n23392 , n13343 , n1159 );
    and g6755 ( n2501 , n1747 , n1078 );
    and g6756 ( n5092 , n20100 , n17634 );
    nor g6757 ( n17562 , n10333 , n9717 );
    and g6758 ( n20797 , n11425 , n15957 );
    not g6759 ( n13935 , n2479 );
    or g6760 ( n10717 , n2833 , n7098 );
    or g6761 ( n21371 , n25751 , n23190 );
    or g6762 ( n6945 , n22024 , n23977 );
    xnor g6763 ( n15464 , n14845 , n23572 );
    not g6764 ( n14038 , n16970 );
    not g6765 ( n12741 , n17872 );
    xnor g6766 ( n22533 , n21003 , n16182 );
    not g6767 ( n19150 , n6556 );
    xnor g6768 ( n13403 , n8600 , n19627 );
    or g6769 ( n24852 , n9700 , n9969 );
    or g6770 ( n10491 , n25974 , n6963 );
    or g6771 ( n5237 , n21556 , n2035 );
    and g6772 ( n22955 , n10206 , n22938 );
    xnor g6773 ( n11713 , n10191 , n20006 );
    or g6774 ( n7659 , n24366 , n5438 );
    nor g6775 ( n13770 , n23592 , n468 );
    and g6776 ( n16266 , n26827 , n21303 );
    xnor g6777 ( n10404 , n17700 , n19089 );
    xnor g6778 ( n24965 , n24367 , n27099 );
    xnor g6779 ( n19317 , n7226 , n20693 );
    xnor g6780 ( n1484 , n3070 , n13568 );
    not g6781 ( n7761 , n25555 );
    or g6782 ( n10332 , n21697 , n1542 );
    or g6783 ( n4669 , n8732 , n4651 );
    or g6784 ( n27157 , n11694 , n14521 );
    nor g6785 ( n20422 , n3791 , n7437 );
    nor g6786 ( n3297 , n24590 , n22480 );
    nor g6787 ( n22412 , n7049 , n21219 );
    not g6788 ( n5234 , n13672 );
    nor g6789 ( n5044 , n17415 , n16822 );
    xnor g6790 ( n12047 , n101 , n21643 );
    nor g6791 ( n26120 , n3550 , n5171 );
    nor g6792 ( n23848 , n5077 , n17397 );
    nor g6793 ( n25916 , n4245 , n5599 );
    and g6794 ( n5310 , n21178 , n8357 );
    nor g6795 ( n9216 , n14536 , n1320 );
    xnor g6796 ( n25250 , n24235 , n2345 );
    not g6797 ( n300 , n18068 );
    nor g6798 ( n20814 , n26557 , n10048 );
    or g6799 ( n26503 , n3721 , n1855 );
    and g6800 ( n19975 , n22052 , n19231 );
    nor g6801 ( n26129 , n8827 , n8176 );
    xnor g6802 ( n8550 , n6552 , n21045 );
    or g6803 ( n5000 , n19962 , n19527 );
    not g6804 ( n25886 , n25974 );
    nor g6805 ( n22763 , n3710 , n26399 );
    nor g6806 ( n8118 , n18300 , n13303 );
    not g6807 ( n11014 , n26046 );
    or g6808 ( n3482 , n21117 , n20700 );
    and g6809 ( n15228 , n23483 , n26938 );
    or g6810 ( n9794 , n16210 , n2731 );
    xnor g6811 ( n10021 , n24502 , n13617 );
    and g6812 ( n13388 , n18926 , n2705 );
    nor g6813 ( n21307 , n20271 , n11693 );
    or g6814 ( n1485 , n19818 , n12388 );
    xnor g6815 ( n23669 , n23607 , n11812 );
    or g6816 ( n12404 , n6255 , n8704 );
    or g6817 ( n17644 , n8792 , n3764 );
    xnor g6818 ( n16387 , n10300 , n24829 );
    nor g6819 ( n12478 , n13851 , n7010 );
    xnor g6820 ( n18346 , n2718 , n14981 );
    and g6821 ( n23542 , n3892 , n6942 );
    and g6822 ( n12625 , n24153 , n1445 );
    not g6823 ( n8253 , n1245 );
    or g6824 ( n20784 , n19340 , n7241 );
    and g6825 ( n24573 , n23098 , n20550 );
    or g6826 ( n25970 , n6571 , n12549 );
    not g6827 ( n17647 , n23894 );
    or g6828 ( n4444 , n10227 , n3102 );
    xnor g6829 ( n20592 , n26556 , n5438 );
    and g6830 ( n22990 , n752 , n11504 );
    xnor g6831 ( n10897 , n24379 , n18810 );
    nor g6832 ( n14939 , n11383 , n23558 );
    or g6833 ( n4619 , n4436 , n21406 );
    and g6834 ( n16088 , n8977 , n18821 );
    not g6835 ( n20266 , n6933 );
    not g6836 ( n19607 , n3751 );
    or g6837 ( n18805 , n15182 , n2996 );
    nor g6838 ( n13411 , n481 , n13951 );
    xnor g6839 ( n9845 , n14106 , n16880 );
    not g6840 ( n10249 , n10454 );
    and g6841 ( n21150 , n24804 , n17015 );
    and g6842 ( n9587 , n18345 , n22700 );
    xnor g6843 ( n11576 , n15440 , n3147 );
    xnor g6844 ( n15275 , n15412 , n10731 );
    xnor g6845 ( n6678 , n21848 , n11230 );
    xnor g6846 ( n24538 , n21693 , n15875 );
    not g6847 ( n12921 , n19618 );
    xnor g6848 ( n11344 , n25622 , n19186 );
    xnor g6849 ( n20727 , n25360 , n2102 );
    not g6850 ( n3415 , n22782 );
    nor g6851 ( n13483 , n5538 , n5772 );
    nor g6852 ( n17649 , n22274 , n22591 );
    xnor g6853 ( n15499 , n14870 , n8888 );
    nor g6854 ( n25783 , n18351 , n5690 );
    and g6855 ( n6951 , n1628 , n24971 );
    xnor g6856 ( n6392 , n2168 , n9502 );
    and g6857 ( n24914 , n22805 , n10297 );
    xnor g6858 ( n22322 , n21020 , n13703 );
    or g6859 ( n18234 , n23913 , n7274 );
    and g6860 ( n25060 , n8738 , n17700 );
    or g6861 ( n2475 , n2130 , n16921 );
    and g6862 ( n9654 , n15323 , n25177 );
    nor g6863 ( n8532 , n20638 , n3540 );
    or g6864 ( n17769 , n5321 , n22628 );
    or g6865 ( n18695 , n23744 , n5380 );
    and g6866 ( n531 , n1742 , n1798 );
    xnor g6867 ( n22341 , n8894 , n24441 );
    xnor g6868 ( n23213 , n5783 , n11432 );
    or g6869 ( n23726 , n5440 , n4326 );
    and g6870 ( n17352 , n1573 , n4652 );
    or g6871 ( n24204 , n23228 , n10460 );
    or g6872 ( n10302 , n4963 , n2818 );
    xnor g6873 ( n5055 , n23801 , n16646 );
    and g6874 ( n15306 , n20860 , n15020 );
    and g6875 ( n4036 , n4149 , n24799 );
    xnor g6876 ( n11743 , n22636 , n16971 );
    and g6877 ( n5509 , n7334 , n5925 );
    not g6878 ( n16351 , n14826 );
    xnor g6879 ( n6375 , n1171 , n5456 );
    and g6880 ( n2622 , n16817 , n24401 );
    nor g6881 ( n20079 , n20478 , n26030 );
    or g6882 ( n25039 , n19422 , n14082 );
    xnor g6883 ( n15701 , n23272 , n14826 );
    and g6884 ( n26642 , n23580 , n8925 );
    not g6885 ( n3783 , n4007 );
    or g6886 ( n5878 , n6261 , n292 );
    or g6887 ( n23811 , n4530 , n14165 );
    xnor g6888 ( n2981 , n1244 , n11779 );
    nor g6889 ( n17083 , n16483 , n18846 );
    or g6890 ( n23439 , n12503 , n13362 );
    and g6891 ( n15677 , n7247 , n6002 );
    and g6892 ( n7124 , n9187 , n4870 );
    not g6893 ( n24593 , n21894 );
    or g6894 ( n6992 , n6847 , n2051 );
    xnor g6895 ( n897 , n7162 , n21226 );
    or g6896 ( n17672 , n5933 , n625 );
    and g6897 ( n14416 , n19481 , n12052 );
    not g6898 ( n24823 , n15332 );
    and g6899 ( n6832 , n25663 , n16721 );
    and g6900 ( n27029 , n1702 , n2733 );
    or g6901 ( n4297 , n4859 , n14584 );
    not g6902 ( n12457 , n15985 );
    and g6903 ( n2539 , n7621 , n7217 );
    and g6904 ( n1327 , n20138 , n26093 );
    or g6905 ( n15410 , n1340 , n16561 );
    and g6906 ( n18796 , n18937 , n11942 );
    or g6907 ( n16268 , n1472 , n14057 );
    and g6908 ( n14751 , n6039 , n9394 );
    xnor g6909 ( n19424 , n5944 , n21231 );
    nor g6910 ( n7106 , n3791 , n7330 );
    not g6911 ( n2246 , n10114 );
    nor g6912 ( n16881 , n10049 , n6790 );
    xnor g6913 ( n1344 , n18956 , n10427 );
    or g6914 ( n1670 , n22053 , n1388 );
    or g6915 ( n4907 , n26204 , n24360 );
    not g6916 ( n8434 , n23630 );
    or g6917 ( n21090 , n19493 , n25521 );
    xnor g6918 ( n15610 , n18203 , n18909 );
    not g6919 ( n3236 , n7406 );
    xnor g6920 ( n16729 , n17468 , n20021 );
    and g6921 ( n11305 , n23027 , n9734 );
    or g6922 ( n205 , n21340 , n24266 );
    or g6923 ( n21023 , n21306 , n9440 );
    xnor g6924 ( n20149 , n6419 , n20607 );
    not g6925 ( n21965 , n27081 );
    or g6926 ( n11759 , n19898 , n12531 );
    and g6927 ( n26840 , n7148 , n23 );
    and g6928 ( n13972 , n2763 , n15330 );
    and g6929 ( n27201 , n13823 , n14166 );
    or g6930 ( n26084 , n26603 , n6280 );
    or g6931 ( n26911 , n10184 , n27037 );
    nor g6932 ( n3139 , n1558 , n11566 );
    not g6933 ( n21988 , n7486 );
    or g6934 ( n10426 , n8006 , n19514 );
    xnor g6935 ( n24807 , n26516 , n10278 );
    or g6936 ( n165 , n20750 , n24843 );
    or g6937 ( n17554 , n12720 , n19192 );
    not g6938 ( n21113 , n12367 );
    xnor g6939 ( n4160 , n18195 , n18177 );
    or g6940 ( n8269 , n16712 , n24278 );
    xnor g6941 ( n23853 , n12902 , n14198 );
    or g6942 ( n23345 , n19082 , n19321 );
    and g6943 ( n17384 , n22631 , n22613 );
    not g6944 ( n22315 , n9990 );
    and g6945 ( n20567 , n23250 , n16856 );
    or g6946 ( n26110 , n21304 , n15468 );
    not g6947 ( n23161 , n16232 );
    xnor g6948 ( n8945 , n12466 , n5022 );
    xnor g6949 ( n23405 , n13171 , n23068 );
    not g6950 ( n19875 , n16729 );
    xnor g6951 ( n14998 , n16994 , n4964 );
    xnor g6952 ( n4487 , n22021 , n2145 );
    xnor g6953 ( n61 , n5212 , n18145 );
    and g6954 ( n12095 , n25205 , n6839 );
    xnor g6955 ( n2868 , n6667 , n22509 );
    xnor g6956 ( n18999 , n6370 , n13070 );
    xnor g6957 ( n16809 , n24711 , n4760 );
    xnor g6958 ( n11920 , n12660 , n27188 );
    not g6959 ( n25114 , n8527 );
    xnor g6960 ( n860 , n3403 , n4193 );
    xnor g6961 ( n22646 , n15992 , n6093 );
    not g6962 ( n16203 , n8280 );
    xnor g6963 ( n26406 , n24961 , n1709 );
    or g6964 ( n18206 , n20674 , n5010 );
    nor g6965 ( n1935 , n17959 , n17728 );
    xnor g6966 ( n4905 , n25318 , n16544 );
    xnor g6967 ( n5680 , n23904 , n9521 );
    xnor g6968 ( n10504 , n15628 , n18532 );
    and g6969 ( n22536 , n20365 , n14127 );
    not g6970 ( n2776 , n15902 );
    nor g6971 ( n6092 , n9291 , n9077 );
    and g6972 ( n17787 , n18182 , n9336 );
    and g6973 ( n10054 , n18884 , n3224 );
    and g6974 ( n6015 , n5003 , n22941 );
    and g6975 ( n15774 , n26542 , n21403 );
    xnor g6976 ( n25630 , n11849 , n7191 );
    or g6977 ( n22328 , n26864 , n18796 );
    not g6978 ( n23477 , n14090 );
    and g6979 ( n5892 , n9443 , n20188 );
    xnor g6980 ( n477 , n11441 , n22106 );
    xnor g6981 ( n24460 , n2325 , n19248 );
    and g6982 ( n18330 , n6496 , n7307 );
    or g6983 ( n7383 , n11899 , n27201 );
    xnor g6984 ( n19578 , n12022 , n8277 );
    nor g6985 ( n3142 , n16244 , n18759 );
    xnor g6986 ( n1378 , n7871 , n8261 );
    and g6987 ( n4517 , n24797 , n13063 );
    and g6988 ( n10480 , n24135 , n3134 );
    xnor g6989 ( n3149 , n24779 , n21344 );
    or g6990 ( n23074 , n23750 , n22254 );
    xnor g6991 ( n24897 , n2460 , n8439 );
    and g6992 ( n25618 , n18449 , n12588 );
    or g6993 ( n9279 , n11728 , n12641 );
    and g6994 ( n23511 , n4701 , n25675 );
    xnor g6995 ( n1717 , n17751 , n23879 );
    or g6996 ( n4696 , n4555 , n11455 );
    not g6997 ( n5445 , n7387 );
    or g6998 ( n17546 , n15059 , n13207 );
    xnor g6999 ( n13981 , n583 , n13714 );
    or g7000 ( n1818 , n26407 , n3532 );
    xnor g7001 ( n18421 , n6358 , n8962 );
    and g7002 ( n14513 , n9281 , n15621 );
    or g7003 ( n6035 , n7018 , n6737 );
    and g7004 ( n23490 , n7026 , n17835 );
    and g7005 ( n11985 , n16141 , n7533 );
    or g7006 ( n19864 , n11303 , n13133 );
    nor g7007 ( n20371 , n21113 , n23760 );
    or g7008 ( n11715 , n17192 , n26944 );
    xnor g7009 ( n7066 , n17611 , n2030 );
    xnor g7010 ( n11650 , n2188 , n2802 );
    and g7011 ( n8304 , n25968 , n18242 );
    not g7012 ( n1079 , n17555 );
    xnor g7013 ( n18304 , n295 , n27135 );
    nor g7014 ( n15129 , n21912 , n9291 );
    not g7015 ( n15868 , n19305 );
    and g7016 ( n20228 , n914 , n139 );
    xnor g7017 ( n24715 , n6722 , n925 );
    xnor g7018 ( n581 , n22596 , n13263 );
    or g7019 ( n16105 , n1672 , n14244 );
    or g7020 ( n15018 , n17645 , n26405 );
    not g7021 ( n9285 , n4651 );
    xnor g7022 ( n5259 , n20613 , n1599 );
    or g7023 ( n6793 , n22269 , n20217 );
    nor g7024 ( n18378 , n10152 , n7981 );
    and g7025 ( n17656 , n12755 , n24438 );
    xnor g7026 ( n16430 , n7291 , n11128 );
    nor g7027 ( n17757 , n22219 , n4781 );
    and g7028 ( n10839 , n18737 , n2328 );
    and g7029 ( n2247 , n17918 , n24669 );
    and g7030 ( n10810 , n726 , n26849 );
    not g7031 ( n2341 , n20929 );
    xnor g7032 ( n21678 , n26031 , n17154 );
    or g7033 ( n20204 , n5514 , n24175 );
    or g7034 ( n16027 , n13327 , n21401 );
    or g7035 ( n22678 , n20776 , n18660 );
    nor g7036 ( n15133 , n19701 , n2829 );
    and g7037 ( n18652 , n26252 , n16765 );
    or g7038 ( n14134 , n19944 , n5704 );
    xnor g7039 ( n21001 , n22338 , n1992 );
    xnor g7040 ( n25964 , n17388 , n13293 );
    or g7041 ( n1097 , n16482 , n11293 );
    xnor g7042 ( n7830 , n16777 , n16788 );
    xnor g7043 ( n18200 , n6524 , n16851 );
    not g7044 ( n26065 , n15534 );
    xnor g7045 ( n434 , n24630 , n8581 );
    or g7046 ( n4735 , n22634 , n17816 );
    or g7047 ( n20367 , n6262 , n8165 );
    or g7048 ( n2910 , n9849 , n17039 );
    xnor g7049 ( n17102 , n10651 , n19515 );
    or g7050 ( n24699 , n4147 , n20862 );
    xnor g7051 ( n4566 , n23352 , n15761 );
    not g7052 ( n1906 , n1456 );
    and g7053 ( n9179 , n25982 , n18262 );
    and g7054 ( n8100 , n17871 , n6894 );
    and g7055 ( n20304 , n8163 , n7173 );
    nor g7056 ( n17929 , n19005 , n24618 );
    and g7057 ( n12400 , n25905 , n17146 );
    nor g7058 ( n19550 , n20721 , n2615 );
    and g7059 ( n2890 , n25411 , n6977 );
    or g7060 ( n12486 , n17474 , n16553 );
    not g7061 ( n4461 , n23767 );
    not g7062 ( n13224 , n23086 );
    xnor g7063 ( n14398 , n2834 , n8545 );
    and g7064 ( n22013 , n15130 , n25567 );
    nor g7065 ( n16383 , n2568 , n22091 );
    and g7066 ( n18389 , n8586 , n23577 );
    xnor g7067 ( n6402 , n7837 , n26545 );
    xnor g7068 ( n23293 , n19127 , n18200 );
    xnor g7069 ( n22439 , n754 , n10547 );
    or g7070 ( n4838 , n1068 , n22594 );
    xnor g7071 ( n6852 , n12291 , n24933 );
    not g7072 ( n19843 , n13784 );
    xnor g7073 ( n3126 , n22570 , n22249 );
    or g7074 ( n25986 , n4550 , n14379 );
    or g7075 ( n11598 , n18341 , n18262 );
    or g7076 ( n6880 , n6129 , n14749 );
    not g7077 ( n8677 , n5532 );
    and g7078 ( n20315 , n4040 , n16009 );
    buf g7079 ( n16573 , n3471 );
    and g7080 ( n26364 , n5021 , n22553 );
    xnor g7081 ( n6583 , n15182 , n26797 );
    xnor g7082 ( n10996 , n5779 , n25001 );
    and g7083 ( n10980 , n5160 , n8901 );
    xnor g7084 ( n24456 , n24855 , n21328 );
    and g7085 ( n9983 , n5523 , n2653 );
    xnor g7086 ( n16871 , n20084 , n10207 );
    or g7087 ( n1873 , n2576 , n8819 );
    and g7088 ( n22119 , n5647 , n20320 );
    xnor g7089 ( n5751 , n8929 , n10012 );
    or g7090 ( n4787 , n23477 , n6794 );
    xnor g7091 ( n6862 , n12372 , n15881 );
    or g7092 ( n2082 , n19579 , n19729 );
    xnor g7093 ( n12148 , n17143 , n7566 );
    and g7094 ( n19871 , n11904 , n11422 );
    not g7095 ( n7740 , n14922 );
    xnor g7096 ( n924 , n10713 , n25494 );
    or g7097 ( n254 , n24428 , n12450 );
    not g7098 ( n4868 , n25475 );
    and g7099 ( n25707 , n25624 , n9653 );
    or g7100 ( n24822 , n4049 , n19529 );
    or g7101 ( n10545 , n9264 , n19990 );
    not g7102 ( n13371 , n13183 );
    not g7103 ( n19406 , n26264 );
    and g7104 ( n5801 , n16530 , n16735 );
    and g7105 ( n1986 , n24566 , n17477 );
    xnor g7106 ( n11514 , n11308 , n3697 );
    and g7107 ( n17751 , n24894 , n25433 );
    or g7108 ( n21690 , n13527 , n16118 );
    xnor g7109 ( n13271 , n24624 , n13565 );
    xnor g7110 ( n20182 , n10481 , n3407 );
    nor g7111 ( n11659 , n21071 , n7906 );
    not g7112 ( n21633 , n1852 );
    xnor g7113 ( n664 , n23993 , n5640 );
    or g7114 ( n17374 , n19438 , n798 );
    xnor g7115 ( n2095 , n12015 , n7840 );
    not g7116 ( n23750 , n23160 );
    nor g7117 ( n16666 , n16430 , n10915 );
    not g7118 ( n4562 , n4423 );
    not g7119 ( n3204 , n4272 );
    or g7120 ( n16766 , n18676 , n6135 );
    or g7121 ( n5941 , n15142 , n20120 );
    nor g7122 ( n19604 , n20049 , n13806 );
    xnor g7123 ( n3751 , n11547 , n3713 );
    or g7124 ( n7591 , n1054 , n6941 );
    or g7125 ( n9052 , n6504 , n3618 );
    xnor g7126 ( n1634 , n25005 , n5195 );
    nor g7127 ( n12091 , n7924 , n11333 );
    or g7128 ( n1375 , n15430 , n25226 );
    not g7129 ( n5740 , n8890 );
    not g7130 ( n9058 , n4235 );
    or g7131 ( n5535 , n18100 , n15743 );
    and g7132 ( n13579 , n3822 , n26357 );
    xnor g7133 ( n1549 , n13460 , n22335 );
    and g7134 ( n13370 , n22375 , n5722 );
    nor g7135 ( n24432 , n5213 , n4812 );
    xnor g7136 ( n10315 , n12422 , n5616 );
    xnor g7137 ( n1844 , n17197 , n19618 );
    or g7138 ( n13433 , n4254 , n21413 );
    xnor g7139 ( n10108 , n2298 , n21749 );
    or g7140 ( n24013 , n12769 , n25405 );
    and g7141 ( n10490 , n13104 , n5993 );
    xnor g7142 ( n11952 , n20929 , n6596 );
    and g7143 ( n16118 , n4337 , n10600 );
    or g7144 ( n2982 , n23491 , n14659 );
    xnor g7145 ( n13031 , n24366 , n18151 );
    not g7146 ( n6209 , n1630 );
    xnor g7147 ( n25147 , n24496 , n22210 );
    nor g7148 ( n2319 , n16938 , n8775 );
    not g7149 ( n14411 , n26703 );
    nor g7150 ( n9764 , n18173 , n25494 );
    xnor g7151 ( n14746 , n22864 , n23165 );
    and g7152 ( n26924 , n25351 , n1331 );
    xnor g7153 ( n17000 , n547 , n8090 );
    nor g7154 ( n21313 , n21222 , n26565 );
    or g7155 ( n21156 , n7305 , n1204 );
    and g7156 ( n7199 , n14137 , n4726 );
    and g7157 ( n3195 , n20524 , n9571 );
    nor g7158 ( n18430 , n10183 , n24824 );
    xnor g7159 ( n23901 , n6331 , n15822 );
    xnor g7160 ( n8732 , n14639 , n15663 );
    xnor g7161 ( n23715 , n17840 , n8834 );
    not g7162 ( n12640 , n13263 );
    or g7163 ( n10544 , n6904 , n3161 );
    or g7164 ( n25234 , n4859 , n9793 );
    or g7165 ( n20950 , n18530 , n12526 );
    xnor g7166 ( n9808 , n12811 , n19514 );
    and g7167 ( n21536 , n19886 , n2391 );
    and g7168 ( n3500 , n24547 , n15151 );
    xnor g7169 ( n14278 , n18655 , n8875 );
    xnor g7170 ( n9486 , n21693 , n20489 );
    or g7171 ( n14608 , n7987 , n10911 );
    nor g7172 ( n9756 , n20964 , n17077 );
    or g7173 ( n26258 , n26717 , n16083 );
    or g7174 ( n25504 , n14024 , n23568 );
    or g7175 ( n17577 , n13760 , n8682 );
    xnor g7176 ( n10967 , n8815 , n946 );
    and g7177 ( n22028 , n9117 , n20943 );
    not g7178 ( n4606 , n24573 );
    or g7179 ( n2 , n5243 , n24961 );
    not g7180 ( n25810 , n14521 );
    xnor g7181 ( n10239 , n11568 , n13194 );
    and g7182 ( n10371 , n6618 , n25911 );
    and g7183 ( n7706 , n1692 , n13791 );
    xnor g7184 ( n26118 , n10138 , n12419 );
    xnor g7185 ( n7667 , n20920 , n22379 );
    not g7186 ( n5012 , n4085 );
    or g7187 ( n15003 , n22225 , n2842 );
    and g7188 ( n23600 , n18900 , n23839 );
    or g7189 ( n18616 , n24899 , n10160 );
    and g7190 ( n23448 , n12390 , n9747 );
    xnor g7191 ( n22819 , n20451 , n19435 );
    nor g7192 ( n19718 , n10964 , n22260 );
    and g7193 ( n21609 , n2163 , n10346 );
    or g7194 ( n9511 , n9079 , n26042 );
    not g7195 ( n7418 , n16276 );
    or g7196 ( n14445 , n22000 , n11572 );
    or g7197 ( n11631 , n8819 , n10869 );
    xnor g7198 ( n26179 , n7863 , n25606 );
    not g7199 ( n5103 , n15705 );
    xnor g7200 ( n1011 , n10357 , n6444 );
    not g7201 ( n17542 , n10125 );
    nor g7202 ( n4227 , n8571 , n25240 );
    not g7203 ( n23536 , n23308 );
    or g7204 ( n8231 , n24118 , n2525 );
    or g7205 ( n13294 , n22642 , n17515 );
    not g7206 ( n17213 , n23587 );
    nor g7207 ( n11728 , n2597 , n13989 );
    and g7208 ( n23462 , n8463 , n24730 );
    buf g7209 ( n1181 , n15339 );
    or g7210 ( n16779 , n20222 , n4096 );
    not g7211 ( n13731 , n8581 );
    and g7212 ( n12122 , n26036 , n7832 );
    xnor g7213 ( n10731 , n18925 , n25150 );
    or g7214 ( n3036 , n20981 , n20646 );
    xnor g7215 ( n2582 , n22064 , n21491 );
    xnor g7216 ( n25001 , n21880 , n11420 );
    xnor g7217 ( n7502 , n20249 , n21352 );
    not g7218 ( n9200 , n26546 );
    xnor g7219 ( n858 , n138 , n10284 );
    not g7220 ( n25987 , n11824 );
    xnor g7221 ( n2887 , n11319 , n13793 );
    not g7222 ( n3515 , n9754 );
    and g7223 ( n9316 , n15525 , n8145 );
    or g7224 ( n22800 , n11268 , n13831 );
    or g7225 ( n2893 , n26597 , n16296 );
    not g7226 ( n12494 , n26942 );
    not g7227 ( n22345 , n1886 );
    nor g7228 ( n18517 , n15426 , n8745 );
    or g7229 ( n20434 , n15858 , n14474 );
    xnor g7230 ( n20706 , n18846 , n16483 );
    xnor g7231 ( n6147 , n16470 , n755 );
    or g7232 ( n18808 , n18227 , n21828 );
    xnor g7233 ( n14989 , n10058 , n10645 );
    and g7234 ( n9647 , n25987 , n14122 );
    not g7235 ( n15932 , n16541 );
    and g7236 ( n22243 , n17978 , n7223 );
    xnor g7237 ( n21511 , n19218 , n985 );
    nor g7238 ( n4594 , n19453 , n12018 );
    xnor g7239 ( n26849 , n16553 , n17112 );
    and g7240 ( n143 , n15271 , n24850 );
    and g7241 ( n15023 , n4878 , n12102 );
    or g7242 ( n2364 , n14430 , n10887 );
    and g7243 ( n17587 , n20258 , n3442 );
    xnor g7244 ( n19266 , n19742 , n19868 );
    not g7245 ( n11428 , n18714 );
    or g7246 ( n24886 , n5026 , n8581 );
    xnor g7247 ( n4362 , n808 , n23333 );
    and g7248 ( n19597 , n19443 , n22799 );
    xnor g7249 ( n101 , n17480 , n22691 );
    nor g7250 ( n4445 , n13152 , n20455 );
    and g7251 ( n13410 , n2857 , n24821 );
    not g7252 ( n835 , n7006 );
    xnor g7253 ( n9796 , n15113 , n24080 );
    and g7254 ( n24017 , n26671 , n7790 );
    nor g7255 ( n17593 , n1319 , n6864 );
    xnor g7256 ( n17104 , n15024 , n25631 );
    nor g7257 ( n19062 , n4625 , n9523 );
    and g7258 ( n11306 , n17128 , n26912 );
    nor g7259 ( n15527 , n8322 , n12811 );
    and g7260 ( n8922 , n26264 , n20326 );
    xnor g7261 ( n20869 , n25717 , n18700 );
    or g7262 ( n20890 , n18726 , n11910 );
    not g7263 ( n5474 , n20594 );
    nor g7264 ( n4012 , n3878 , n22421 );
    xnor g7265 ( n10451 , n16170 , n6149 );
    and g7266 ( n9551 , n4110 , n17283 );
    or g7267 ( n24068 , n23484 , n19286 );
    xnor g7268 ( n5348 , n19816 , n7709 );
    xnor g7269 ( n9763 , n15953 , n3800 );
    nor g7270 ( n1234 , n3776 , n12709 );
    xnor g7271 ( n8106 , n14494 , n13837 );
    or g7272 ( n19362 , n10873 , n4572 );
    and g7273 ( n23556 , n570 , n18461 );
    nor g7274 ( n22167 , n15113 , n24080 );
    and g7275 ( n17634 , n17286 , n20968 );
    or g7276 ( n3392 , n14131 , n26680 );
    xnor g7277 ( n24609 , n22137 , n7887 );
    and g7278 ( n6846 , n8516 , n7565 );
    xnor g7279 ( n6094 , n25092 , n10263 );
    and g7280 ( n23147 , n23040 , n25782 );
    xnor g7281 ( n18254 , n17941 , n3082 );
    xnor g7282 ( n18589 , n17657 , n20546 );
    and g7283 ( n848 , n15494 , n20046 );
    not g7284 ( n12064 , n24166 );
    xnor g7285 ( n14229 , n24554 , n24032 );
    or g7286 ( n3285 , n1406 , n11486 );
    not g7287 ( n5006 , n10710 );
    xnor g7288 ( n13932 , n7832 , n7697 );
    not g7289 ( n7981 , n10437 );
    xnor g7290 ( n11639 , n8338 , n15521 );
    xnor g7291 ( n6184 , n2052 , n13631 );
    nor g7292 ( n9539 , n12802 , n3707 );
    xnor g7293 ( n11772 , n23710 , n5793 );
    and g7294 ( n27084 , n10951 , n1577 );
    or g7295 ( n10823 , n20759 , n6766 );
    xnor g7296 ( n8888 , n24110 , n27036 );
    xnor g7297 ( n5810 , n4801 , n20557 );
    xnor g7298 ( n23300 , n26170 , n23664 );
    or g7299 ( n17128 , n21967 , n4106 );
    xnor g7300 ( n24392 , n9202 , n14790 );
    xnor g7301 ( n6084 , n19629 , n10520 );
    or g7302 ( n9727 , n15585 , n13505 );
    and g7303 ( n23198 , n14440 , n14718 );
    not g7304 ( n4622 , n8806 );
    xnor g7305 ( n20687 , n10004 , n15701 );
    xnor g7306 ( n1138 , n26143 , n7388 );
    or g7307 ( n22748 , n13921 , n16877 );
    xnor g7308 ( n9166 , n5620 , n1640 );
    and g7309 ( n5084 , n8784 , n17350 );
    or g7310 ( n14639 , n2115 , n4357 );
    xnor g7311 ( n18898 , n24217 , n15897 );
    and g7312 ( n10317 , n3635 , n22635 );
    nor g7313 ( n6571 , n9187 , n13368 );
    xnor g7314 ( n15725 , n21469 , n4692 );
    not g7315 ( n14733 , n17410 );
    or g7316 ( n19287 , n14633 , n20897 );
    and g7317 ( n5863 , n13007 , n26401 );
    not g7318 ( n4572 , n21502 );
    nor g7319 ( n21861 , n21374 , n10891 );
    nor g7320 ( n11664 , n21774 , n6564 );
    or g7321 ( n9010 , n3326 , n334 );
    or g7322 ( n21516 , n6841 , n1662 );
    xnor g7323 ( n23924 , n165 , n26874 );
    not g7324 ( n18450 , n6015 );
    xnor g7325 ( n14400 , n3381 , n4816 );
    xnor g7326 ( n4725 , n10565 , n8317 );
    nor g7327 ( n12054 , n14781 , n15703 );
    and g7328 ( n7384 , n1558 , n5050 );
    xnor g7329 ( n23258 , n23520 , n21355 );
    or g7330 ( n8705 , n10890 , n17510 );
    and g7331 ( n17498 , n11359 , n26114 );
    and g7332 ( n16623 , n23757 , n8195 );
    or g7333 ( n5967 , n17255 , n24213 );
    xnor g7334 ( n8734 , n11302 , n12341 );
    or g7335 ( n26356 , n6251 , n18972 );
    xnor g7336 ( n24563 , n1118 , n20489 );
    and g7337 ( n7454 , n22132 , n1306 );
    not g7338 ( n11816 , n26408 );
    not g7339 ( n2385 , n12851 );
    not g7340 ( n6034 , n18277 );
    and g7341 ( n16810 , n7427 , n24113 );
    or g7342 ( n3546 , n16015 , n21713 );
    xnor g7343 ( n21206 , n14590 , n12890 );
    xnor g7344 ( n8036 , n13263 , n18274 );
    or g7345 ( n5166 , n7683 , n15774 );
    xnor g7346 ( n15678 , n14080 , n19319 );
    and g7347 ( n19566 , n22442 , n3131 );
    or g7348 ( n14297 , n2923 , n757 );
    or g7349 ( n2626 , n21386 , n10763 );
    or g7350 ( n7433 , n869 , n7601 );
    xor g7351 ( n15564 , n2263 , n2507 );
    or g7352 ( n17934 , n143 , n8616 );
    not g7353 ( n13028 , n3962 );
    and g7354 ( n23515 , n9178 , n11549 );
    or g7355 ( n1374 , n7341 , n8925 );
    or g7356 ( n22048 , n6982 , n87 );
    and g7357 ( n26271 , n14620 , n26914 );
    not g7358 ( n3190 , n20429 );
    and g7359 ( n24299 , n20973 , n13539 );
    or g7360 ( n26038 , n22776 , n10353 );
    xnor g7361 ( n15681 , n5601 , n4256 );
    xnor g7362 ( n5865 , n12113 , n12917 );
    and g7363 ( n20325 , n5140 , n14158 );
    and g7364 ( n14696 , n8822 , n6459 );
    xnor g7365 ( n20126 , n5232 , n10289 );
    xnor g7366 ( n3964 , n5496 , n19144 );
    or g7367 ( n13630 , n13991 , n5138 );
    xnor g7368 ( n1942 , n5289 , n26826 );
    and g7369 ( n6390 , n2452 , n11007 );
    or g7370 ( n19507 , n19347 , n13228 );
    and g7371 ( n13818 , n23459 , n10603 );
    and g7372 ( n18331 , n10918 , n5633 );
    xnor g7373 ( n16959 , n8358 , n24344 );
    nor g7374 ( n14017 , n10369 , n599 );
    xnor g7375 ( n27173 , n15490 , n24032 );
    nor g7376 ( n3174 , n10633 , n8378 );
    or g7377 ( n11704 , n15623 , n13904 );
    or g7378 ( n10364 , n3127 , n6060 );
    xnor g7379 ( n3911 , n25778 , n7223 );
    nor g7380 ( n13406 , n12929 , n19005 );
    or g7381 ( n15184 , n3253 , n6246 );
    xnor g7382 ( n20048 , n5934 , n12908 );
    or g7383 ( n3057 , n9843 , n2024 );
    nor g7384 ( n4418 , n15426 , n3136 );
    nor g7385 ( n356 , n22558 , n17803 );
    xnor g7386 ( n2779 , n5588 , n9620 );
    xnor g7387 ( n21989 , n21021 , n15918 );
    or g7388 ( n26263 , n21795 , n4762 );
    xnor g7389 ( n14993 , n12811 , n5213 );
    and g7390 ( n17091 , n19459 , n5160 );
    xnor g7391 ( n5905 , n6363 , n16469 );
    xnor g7392 ( n14163 , n22246 , n14975 );
    and g7393 ( n23046 , n22316 , n931 );
    nor g7394 ( n21259 , n4577 , n9799 );
    and g7395 ( n26448 , n7670 , n8227 );
    or g7396 ( n10627 , n6691 , n21753 );
    xnor g7397 ( n3694 , n19423 , n1112 );
    and g7398 ( n21666 , n14233 , n24082 );
    xnor g7399 ( n14089 , n1920 , n17023 );
    or g7400 ( n24153 , n8827 , n4306 );
    and g7401 ( n6410 , n10398 , n12629 );
    and g7402 ( n8857 , n17046 , n18226 );
    not g7403 ( n24503 , n14885 );
    xnor g7404 ( n10077 , n14351 , n18644 );
    not g7405 ( n27144 , n14437 );
    and g7406 ( n16332 , n8780 , n17622 );
    and g7407 ( n52 , n20455 , n2884 );
    xnor g7408 ( n23076 , n5150 , n11433 );
    not g7409 ( n8680 , n27120 );
    or g7410 ( n3676 , n18125 , n10970 );
    not g7411 ( n22093 , n21470 );
    or g7412 ( n7934 , n25658 , n7379 );
    or g7413 ( n24528 , n8777 , n10122 );
    or g7414 ( n26683 , n11559 , n10405 );
    not g7415 ( n6972 , n16888 );
    not g7416 ( n20597 , n592 );
    and g7417 ( n20110 , n17910 , n5546 );
    xnor g7418 ( n8149 , n12257 , n26718 );
    or g7419 ( n3621 , n18797 , n11221 );
    xnor g7420 ( n1716 , n7099 , n2035 );
    and g7421 ( n19644 , n26999 , n14244 );
    and g7422 ( n65 , n8521 , n4652 );
    or g7423 ( n19893 , n1677 , n20264 );
    not g7424 ( n14486 , n20517 );
    not g7425 ( n4240 , n21111 );
    nor g7426 ( n2087 , n25120 , n17458 );
    or g7427 ( n20632 , n2564 , n10695 );
    not g7428 ( n10188 , n11265 );
    xnor g7429 ( n1245 , n10412 , n2992 );
    xnor g7430 ( n15401 , n2187 , n9572 );
    and g7431 ( n26720 , n15436 , n7485 );
    and g7432 ( n13281 , n22118 , n7058 );
    and g7433 ( n5448 , n208 , n2496 );
    and g7434 ( n26339 , n9999 , n9629 );
    and g7435 ( n18815 , n15538 , n7971 );
    not g7436 ( n15512 , n25243 );
    not g7437 ( n14860 , n4719 );
    and g7438 ( n6748 , n3933 , n21079 );
    xnor g7439 ( n22999 , n24245 , n1654 );
    not g7440 ( n21696 , n3643 );
    and g7441 ( n3066 , n21002 , n21906 );
    not g7442 ( n21853 , n13453 );
    xnor g7443 ( n15150 , n24536 , n20150 );
    xnor g7444 ( n10244 , n20461 , n25952 );
    xnor g7445 ( n22217 , n7172 , n11738 );
    xnor g7446 ( n10385 , n26873 , n10680 );
    or g7447 ( n10762 , n26093 , n10529 );
    and g7448 ( n9662 , n26686 , n5571 );
    nor g7449 ( n23601 , n2583 , n17845 );
    or g7450 ( n17265 , n1222 , n15818 );
    xnor g7451 ( n5324 , n15215 , n10910 );
    xnor g7452 ( n25756 , n14742 , n13222 );
    and g7453 ( n3699 , n9854 , n14955 );
    not g7454 ( n22926 , n864 );
    or g7455 ( n12758 , n3670 , n17199 );
    xnor g7456 ( n8776 , n19869 , n23805 );
    not g7457 ( n10918 , n13580 );
    or g7458 ( n5777 , n25096 , n6420 );
    xnor g7459 ( n22502 , n21095 , n25316 );
    or g7460 ( n15708 , n7733 , n16549 );
    and g7461 ( n6647 , n4713 , n14067 );
    nor g7462 ( n12671 , n11211 , n3547 );
    not g7463 ( n658 , n11192 );
    and g7464 ( n21047 , n10339 , n3505 );
    nor g7465 ( n11131 , n27143 , n15572 );
    xnor g7466 ( n14701 , n3168 , n3484 );
    or g7467 ( n22856 , n18438 , n12081 );
    xnor g7468 ( n11210 , n3469 , n10354 );
    and g7469 ( n5937 , n16926 , n18942 );
    nor g7470 ( n913 , n15282 , n23268 );
    or g7471 ( n11233 , n16890 , n18157 );
    xnor g7472 ( n15628 , n14160 , n17170 );
    or g7473 ( n11599 , n20598 , n1491 );
    not g7474 ( n5495 , n10534 );
    not g7475 ( n9523 , n20835 );
    xnor g7476 ( n8577 , n25049 , n2872 );
    nor g7477 ( n4718 , n26483 , n12088 );
    and g7478 ( n8465 , n25421 , n6570 );
    and g7479 ( n13526 , n5726 , n22578 );
    nor g7480 ( n435 , n22342 , n16993 );
    and g7481 ( n25511 , n26959 , n19687 );
    xnor g7482 ( n5817 , n4132 , n4282 );
    xnor g7483 ( n16885 , n3958 , n11002 );
    nor g7484 ( n20952 , n19469 , n9399 );
    nor g7485 ( n11655 , n2518 , n8272 );
    or g7486 ( n10285 , n8343 , n8305 );
    or g7487 ( n24589 , n730 , n7352 );
    or g7488 ( n12528 , n21313 , n20230 );
    and g7489 ( n19626 , n26516 , n16052 );
    xor g7490 ( n940 , n17211 , n4939 );
    not g7491 ( n16022 , n5263 );
    not g7492 ( n7439 , n23109 );
    or g7493 ( n24546 , n9777 , n8502 );
    not g7494 ( n2152 , n16808 );
    or g7495 ( n18226 , n17944 , n24291 );
    xnor g7496 ( n12829 , n15998 , n12386 );
    and g7497 ( n6280 , n5814 , n51 );
    not g7498 ( n26161 , n15698 );
    not g7499 ( n17287 , n9967 );
    not g7500 ( n8509 , n5302 );
    xnor g7501 ( n19354 , n11793 , n9317 );
    xnor g7502 ( n20049 , n13169 , n17696 );
    nor g7503 ( n13058 , n14680 , n25240 );
    and g7504 ( n17851 , n20429 , n22365 );
    or g7505 ( n21902 , n17095 , n26713 );
    xnor g7506 ( n23331 , n26488 , n18907 );
    or g7507 ( n13174 , n19229 , n12929 );
    or g7508 ( n26898 , n15734 , n18664 );
    and g7509 ( n963 , n22015 , n16334 );
    xnor g7510 ( n26829 , n468 , n17911 );
    not g7511 ( n704 , n3746 );
    and g7512 ( n4290 , n22147 , n25720 );
    nor g7513 ( n1937 , n11186 , n12464 );
    not g7514 ( n1215 , n19584 );
    and g7515 ( n2677 , n14537 , n25986 );
    nor g7516 ( n26568 , n5752 , n22780 );
    and g7517 ( n26638 , n3512 , n25970 );
    and g7518 ( n24394 , n10140 , n26525 );
    nor g7519 ( n997 , n9600 , n17613 );
    xnor g7520 ( n10618 , n16793 , n7089 );
    and g7521 ( n5734 , n19808 , n562 );
    or g7522 ( n26730 , n4434 , n23098 );
    and g7523 ( n26383 , n12793 , n16352 );
    and g7524 ( n26635 , n12495 , n24851 );
    not g7525 ( n1190 , n14024 );
    nor g7526 ( n21979 , n20907 , n18107 );
    not g7527 ( n24164 , n13419 );
    xnor g7528 ( n4156 , n21082 , n8026 );
    xnor g7529 ( n26902 , n8221 , n3880 );
    not g7530 ( n63 , n10275 );
    nor g7531 ( n4094 , n4895 , n8393 );
    not g7532 ( n19624 , n17069 );
    or g7533 ( n15934 , n9852 , n10368 );
    not g7534 ( n19888 , n8626 );
    and g7535 ( n4178 , n12111 , n11217 );
    xnor g7536 ( n23872 , n12151 , n7496 );
    xnor g7537 ( n5469 , n2768 , n24327 );
    not g7538 ( n23582 , n7030 );
    not g7539 ( n8571 , n20359 );
    or g7540 ( n19622 , n20695 , n5592 );
    or g7541 ( n21096 , n180 , n6442 );
    or g7542 ( n27023 , n16254 , n22988 );
    or g7543 ( n15954 , n5007 , n22233 );
    and g7544 ( n16603 , n2639 , n8257 );
    xnor g7545 ( n11509 , n11764 , n10349 );
    xnor g7546 ( n27010 , n10505 , n12153 );
    xnor g7547 ( n26958 , n2633 , n4181 );
    xnor g7548 ( n10423 , n14388 , n21575 );
    or g7549 ( n10886 , n7285 , n14600 );
    xnor g7550 ( n11605 , n2219 , n8059 );
    and g7551 ( n5646 , n9174 , n23991 );
    xnor g7552 ( n25957 , n24619 , n19115 );
    not g7553 ( n14301 , n2715 );
    not g7554 ( n12911 , n8292 );
    xnor g7555 ( n12870 , n1131 , n13412 );
    or g7556 ( n24985 , n3410 , n388 );
    nor g7557 ( n14942 , n9827 , n24280 );
    and g7558 ( n22809 , n12871 , n20411 );
    nor g7559 ( n1300 , n5012 , n17578 );
    xnor g7560 ( n4037 , n25126 , n19575 );
    xnor g7561 ( n16448 , n12509 , n7761 );
    xnor g7562 ( n25452 , n4343 , n14976 );
    or g7563 ( n8048 , n2113 , n148 );
    or g7564 ( n4238 , n19903 , n2020 );
    or g7565 ( n22674 , n3356 , n26860 );
    xnor g7566 ( n23749 , n19444 , n20689 );
    and g7567 ( n24257 , n6546 , n6694 );
    or g7568 ( n26631 , n16155 , n5442 );
    nor g7569 ( n13366 , n2540 , n24688 );
    and g7570 ( n14315 , n3475 , n22949 );
    not g7571 ( n22049 , n18519 );
    and g7572 ( n654 , n6573 , n17719 );
    and g7573 ( n14078 , n23094 , n18897 );
    nor g7574 ( n7688 , n25565 , n24374 );
    or g7575 ( n17841 , n24839 , n10219 );
    or g7576 ( n12710 , n14645 , n14429 );
    not g7577 ( n20562 , n23819 );
    xnor g7578 ( n1685 , n26163 , n6850 );
    xnor g7579 ( n14521 , n10635 , n6250 );
    or g7580 ( n12785 , n1679 , n21913 );
    xnor g7581 ( n15277 , n854 , n15206 );
    nor g7582 ( n22664 , n2926 , n17010 );
    or g7583 ( n21519 , n19663 , n8025 );
    and g7584 ( n14360 , n5717 , n4046 );
    not g7585 ( n3931 , n21082 );
    or g7586 ( n11180 , n19888 , n22414 );
    or g7587 ( n26382 , n16044 , n10772 );
    or g7588 ( n12321 , n20181 , n18037 );
    or g7589 ( n17009 , n2142 , n15544 );
    or g7590 ( n7062 , n2944 , n22270 );
    or g7591 ( n26517 , n22817 , n22066 );
    or g7592 ( n19440 , n11089 , n4955 );
    xnor g7593 ( n2943 , n5990 , n7326 );
    xnor g7594 ( n7416 , n9871 , n8240 );
    and g7595 ( n27041 , n2812 , n5736 );
    and g7596 ( n525 , n19271 , n22232 );
    xnor g7597 ( n19948 , n18883 , n21095 );
    not g7598 ( n22410 , n26944 );
    xnor g7599 ( n11730 , n3882 , n22387 );
    xnor g7600 ( n23917 , n6946 , n20124 );
    xnor g7601 ( n24622 , n5261 , n20169 );
    nor g7602 ( n6111 , n11840 , n15423 );
    not g7603 ( n26834 , n7373 );
    or g7604 ( n8883 , n26870 , n7902 );
    not g7605 ( n6085 , n20635 );
    xnor g7606 ( n11801 , n2750 , n7543 );
    nor g7607 ( n10985 , n682 , n3632 );
    or g7608 ( n12922 , n26377 , n25076 );
    or g7609 ( n10182 , n24523 , n22296 );
    xnor g7610 ( n19245 , n10778 , n22574 );
    or g7611 ( n24001 , n21297 , n25993 );
    and g7612 ( n3894 , n18364 , n13655 );
    not g7613 ( n120 , n19922 );
    xnor g7614 ( n13285 , n46 , n26055 );
    nor g7615 ( n616 , n2482 , n7448 );
    or g7616 ( n23308 , n18444 , n25059 );
    or g7617 ( n12858 , n17539 , n246 );
    and g7618 ( n5442 , n21939 , n20298 );
    or g7619 ( n13608 , n553 , n27200 );
    nor g7620 ( n3061 , n15332 , n14792 );
    and g7621 ( n23607 , n1412 , n9848 );
    xnor g7622 ( n271 , n11173 , n12874 );
    xnor g7623 ( n2524 , n12143 , n7258 );
    xnor g7624 ( n22298 , n5821 , n19698 );
    or g7625 ( n15092 , n24230 , n7900 );
    not g7626 ( n18882 , n22442 );
    nor g7627 ( n10661 , n10527 , n4307 );
    xnor g7628 ( n20353 , n23568 , n1660 );
    or g7629 ( n13081 , n19048 , n16955 );
    and g7630 ( n10014 , n514 , n105 );
    nor g7631 ( n11176 , n4076 , n13541 );
    xnor g7632 ( n19681 , n2423 , n24208 );
    xnor g7633 ( n8820 , n1306 , n6364 );
    nor g7634 ( n25744 , n17959 , n13784 );
    and g7635 ( n4580 , n15324 , n4795 );
    xnor g7636 ( n9760 , n25795 , n11587 );
    nor g7637 ( n3160 , n24928 , n24510 );
    and g7638 ( n26865 , n4463 , n11288 );
    xnor g7639 ( n19148 , n24972 , n5429 );
    xnor g7640 ( n11008 , n9921 , n9293 );
    or g7641 ( n11991 , n17463 , n11115 );
    xnor g7642 ( n6119 , n20192 , n12481 );
    nor g7643 ( n1415 , n10029 , n26004 );
    nor g7644 ( n16795 , n4086 , n17858 );
    or g7645 ( n8030 , n13888 , n19316 );
    and g7646 ( n22878 , n23144 , n24371 );
    and g7647 ( n10586 , n4469 , n5987 );
    or g7648 ( n15785 , n22724 , n17610 );
    not g7649 ( n18113 , n7119 );
    and g7650 ( n25889 , n4427 , n4161 );
    not g7651 ( n21015 , n11011 );
    nor g7652 ( n24338 , n17173 , n7731 );
    and g7653 ( n13090 , n168 , n20940 );
    xnor g7654 ( n26399 , n18174 , n7841 );
    and g7655 ( n20662 , n24118 , n2525 );
    xnor g7656 ( n13642 , n354 , n19858 );
    or g7657 ( n24642 , n15887 , n10153 );
    or g7658 ( n7047 , n16467 , n26061 );
    and g7659 ( n19593 , n1215 , n23715 );
    not g7660 ( n4191 , n16638 );
    or g7661 ( n6322 , n17355 , n19036 );
    and g7662 ( n8942 , n16272 , n17024 );
    or g7663 ( n18822 , n2486 , n20015 );
    or g7664 ( n283 , n4243 , n15306 );
    not g7665 ( n7393 , n1999 );
    and g7666 ( n22475 , n7949 , n16609 );
    xnor g7667 ( n2285 , n7457 , n2615 );
    nor g7668 ( n18287 , n2886 , n16609 );
    or g7669 ( n16836 , n1904 , n26667 );
    and g7670 ( n24820 , n13790 , n20679 );
    and g7671 ( n10841 , n26408 , n1186 );
    xnor g7672 ( n15996 , n10126 , n11888 );
    not g7673 ( n13079 , n19730 );
    xnor g7674 ( n3078 , n4716 , n15314 );
    not g7675 ( n4853 , n23605 );
    xnor g7676 ( n914 , n13543 , n19234 );
    and g7677 ( n9638 , n13190 , n23999 );
    and g7678 ( n24718 , n4434 , n23098 );
    xnor g7679 ( n801 , n7542 , n2478 );
    or g7680 ( n1381 , n25590 , n20800 );
    nor g7681 ( n1656 , n17911 , n25331 );
    xnor g7682 ( n1168 , n22906 , n23369 );
    or g7683 ( n18278 , n7226 , n23727 );
    or g7684 ( n13878 , n20553 , n3165 );
    xnor g7685 ( n2517 , n20902 , n5991 );
    not g7686 ( n13979 , n8844 );
    or g7687 ( n26806 , n18327 , n24694 );
    xnor g7688 ( n21232 , n7505 , n25473 );
    not g7689 ( n6206 , n21333 );
    or g7690 ( n8804 , n18189 , n16590 );
    or g7691 ( n23472 , n20470 , n18634 );
    xnor g7692 ( n3617 , n21539 , n13050 );
    and g7693 ( n16949 , n20358 , n16560 );
    nor g7694 ( n5071 , n9888 , n25115 );
    or g7695 ( n1988 , n905 , n7435 );
    or g7696 ( n26372 , n17302 , n18054 );
    or g7697 ( n12498 , n26442 , n11524 );
    nor g7698 ( n26391 , n9124 , n5483 );
    or g7699 ( n2716 , n896 , n22915 );
    and g7700 ( n6528 , n9509 , n6566 );
    nor g7701 ( n22259 , n6724 , n485 );
    or g7702 ( n24426 , n22987 , n6397 );
    xnor g7703 ( n11284 , n3783 , n26452 );
    not g7704 ( n304 , n14330 );
    not g7705 ( n12535 , n919 );
    buf g7706 ( n12891 , n19263 );
    xnor g7707 ( n23514 , n20047 , n9002 );
    xnor g7708 ( n4387 , n22700 , n18345 );
    or g7709 ( n8443 , n23625 , n14101 );
    or g7710 ( n864 , n19201 , n27189 );
    or g7711 ( n15391 , n23913 , n8144 );
    or g7712 ( n9657 , n7168 , n6068 );
    nor g7713 ( n8646 , n12271 , n16233 );
    xnor g7714 ( n23248 , n20435 , n3281 );
    xnor g7715 ( n25656 , n27150 , n253 );
    not g7716 ( n21691 , n24085 );
    not g7717 ( n1192 , n8331 );
    not g7718 ( n19267 , n16233 );
    not g7719 ( n11096 , n11510 );
    or g7720 ( n7626 , n10928 , n1616 );
    xnor g7721 ( n19817 , n24319 , n6971 );
    and g7722 ( n3637 , n14155 , n12004 );
    and g7723 ( n26669 , n21925 , n24763 );
    or g7724 ( n11423 , n4837 , n22995 );
    xnor g7725 ( n23834 , n2100 , n22795 );
    and g7726 ( n12237 , n9003 , n1735 );
    and g7727 ( n7456 , n9097 , n16344 );
    nor g7728 ( n3956 , n11745 , n10017 );
    or g7729 ( n4414 , n14543 , n6988 );
    xnor g7730 ( n18760 , n24312 , n10847 );
    nor g7731 ( n10574 , n24786 , n20754 );
    nor g7732 ( n12362 , n19626 , n151 );
    not g7733 ( n15809 , n15766 );
    not g7734 ( n14543 , n17679 );
    and g7735 ( n15517 , n26186 , n1028 );
    not g7736 ( n17339 , n5599 );
    or g7737 ( n21863 , n15560 , n300 );
    xnor g7738 ( n4000 , n26677 , n26330 );
    or g7739 ( n22866 , n5394 , n19739 );
    xnor g7740 ( n21335 , n12902 , n26634 );
    and g7741 ( n15340 , n18705 , n8083 );
    xnor g7742 ( n24722 , n3354 , n1834 );
    or g7743 ( n14224 , n23832 , n19238 );
    not g7744 ( n20274 , n14941 );
    not g7745 ( n11394 , n19162 );
    nor g7746 ( n8408 , n4786 , n4608 );
    or g7747 ( n23741 , n25221 , n19425 );
    not g7748 ( n22170 , n26452 );
    and g7749 ( n7672 , n12958 , n14413 );
    xnor g7750 ( n25303 , n25877 , n5026 );
    xnor g7751 ( n24340 , n3295 , n12463 );
    nor g7752 ( n2833 , n25289 , n4195 );
    xnor g7753 ( n4124 , n25877 , n10057 );
    and g7754 ( n24759 , n24022 , n1043 );
    xnor g7755 ( n5253 , n21576 , n21559 );
    or g7756 ( n7127 , n9469 , n14094 );
    and g7757 ( n23881 , n8294 , n10476 );
    xnor g7758 ( n3830 , n12543 , n9090 );
    xnor g7759 ( n4893 , n5699 , n20025 );
    or g7760 ( n25845 , n26871 , n15791 );
    and g7761 ( n666 , n2855 , n19287 );
    and g7762 ( n7101 , n10885 , n19276 );
    nor g7763 ( n2207 , n26224 , n18483 );
    xnor g7764 ( n12349 , n27180 , n21511 );
    or g7765 ( n19093 , n16718 , n22218 );
    and g7766 ( n4065 , n5272 , n22526 );
    xnor g7767 ( n9182 , n6324 , n14531 );
    xnor g7768 ( n21874 , n7696 , n11017 );
    nor g7769 ( n1089 , n26318 , n11248 );
    and g7770 ( n8452 , n10310 , n14093 );
    or g7771 ( n3658 , n10071 , n6490 );
    or g7772 ( n8290 , n6508 , n13336 );
    xnor g7773 ( n4756 , n15437 , n8001 );
    xnor g7774 ( n16694 , n6553 , n12446 );
    or g7775 ( n12882 , n18745 , n5510 );
    not g7776 ( n17453 , n25972 );
    not g7777 ( n4605 , n7828 );
    or g7778 ( n3874 , n20733 , n3710 );
    and g7779 ( n12065 , n6165 , n23183 );
    xnor g7780 ( n1671 , n3919 , n26105 );
    or g7781 ( n2437 , n10418 , n19211 );
    nor g7782 ( n384 , n23921 , n130 );
    xnor g7783 ( n15775 , n1122 , n5365 );
    or g7784 ( n764 , n3243 , n17073 );
    xnor g7785 ( n17170 , n1630 , n4326 );
    or g7786 ( n4742 , n16511 , n25825 );
    nor g7787 ( n1224 , n5604 , n7026 );
    nor g7788 ( n19359 , n20131 , n17418 );
    xnor g7789 ( n25815 , n1753 , n19457 );
    or g7790 ( n14286 , n1359 , n7252 );
    xnor g7791 ( n9458 , n18910 , n4168 );
    xnor g7792 ( n7992 , n18401 , n12772 );
    or g7793 ( n26820 , n958 , n9658 );
    not g7794 ( n20059 , n5956 );
    or g7795 ( n4919 , n12562 , n23978 );
    nor g7796 ( n20740 , n15295 , n3195 );
    and g7797 ( n7450 , n18475 , n15197 );
    xnor g7798 ( n11617 , n15743 , n13319 );
    xnor g7799 ( n14919 , n2646 , n22072 );
    xnor g7800 ( n19734 , n19806 , n24024 );
    and g7801 ( n19160 , n20576 , n15349 );
    or g7802 ( n26569 , n20137 , n17601 );
    not g7803 ( n15686 , n10069 );
    or g7804 ( n26659 , n21556 , n21207 );
    or g7805 ( n24672 , n11816 , n8649 );
    nor g7806 ( n25649 , n342 , n14570 );
    and g7807 ( n8940 , n1379 , n9105 );
    or g7808 ( n4197 , n20491 , n20769 );
    not g7809 ( n21288 , n24440 );
    xnor g7810 ( n19236 , n11117 , n21980 );
    not g7811 ( n3094 , n26053 );
    nor g7812 ( n18580 , n24306 , n9116 );
    not g7813 ( n1155 , n20966 );
    and g7814 ( n16193 , n12967 , n11030 );
    or g7815 ( n23839 , n1935 , n17552 );
    xnor g7816 ( n3584 , n16184 , n13247 );
    xnor g7817 ( n10705 , n25036 , n11016 );
    not g7818 ( n2360 , n20687 );
    and g7819 ( n24247 , n27111 , n3391 );
    xnor g7820 ( n16692 , n18861 , n10251 );
    and g7821 ( n4057 , n26503 , n25702 );
    and g7822 ( n25906 , n17770 , n12629 );
    or g7823 ( n5959 , n1107 , n17257 );
    xnor g7824 ( n5110 , n24846 , n16714 );
    and g7825 ( n9716 , n6508 , n21710 );
    not g7826 ( n9957 , n11136 );
    nor g7827 ( n5602 , n21502 , n4017 );
    or g7828 ( n5056 , n823 , n19010 );
    nor g7829 ( n382 , n2764 , n9789 );
    xnor g7830 ( n16689 , n19228 , n4812 );
    or g7831 ( n7112 , n13933 , n24275 );
    nor g7832 ( n9549 , n20117 , n9460 );
    and g7833 ( n23236 , n3110 , n9902 );
    or g7834 ( n3615 , n20688 , n3424 );
    xnor g7835 ( n671 , n21253 , n17664 );
    xnor g7836 ( n25441 , n4016 , n24474 );
    xnor g7837 ( n16076 , n17871 , n12675 );
    and g7838 ( n16526 , n10870 , n8187 );
    and g7839 ( n17724 , n205 , n22842 );
    xnor g7840 ( n10751 , n26410 , n23918 );
    or g7841 ( n4971 , n9076 , n3727 );
    xnor g7842 ( n18574 , n7334 , n6728 );
    and g7843 ( n8740 , n3827 , n5055 );
    xnor g7844 ( n3054 , n25120 , n8526 );
    xnor g7845 ( n13261 , n26625 , n14230 );
    or g7846 ( n16338 , n5729 , n10308 );
    or g7847 ( n3704 , n20874 , n13819 );
    or g7848 ( n24539 , n21672 , n18314 );
    nor g7849 ( n4243 , n5768 , n2300 );
    and g7850 ( n18107 , n7311 , n20273 );
    and g7851 ( n10855 , n12431 , n22189 );
    xnor g7852 ( n5794 , n7499 , n1223 );
    or g7853 ( n10189 , n11544 , n2978 );
    nor g7854 ( n21942 , n16349 , n8094 );
    and g7855 ( n9102 , n16468 , n15511 );
    and g7856 ( n24628 , n5043 , n18133 );
    not g7857 ( n7893 , n21997 );
    or g7858 ( n1596 , n1777 , n837 );
    xnor g7859 ( n22392 , n6775 , n12121 );
    or g7860 ( n3969 , n19631 , n14449 );
    xnor g7861 ( n25222 , n6169 , n6944 );
    nor g7862 ( n24157 , n3582 , n23064 );
    xnor g7863 ( n17713 , n18798 , n25486 );
    or g7864 ( n5174 , n20358 , n3960 );
    and g7865 ( n15012 , n20040 , n8186 );
    and g7866 ( n16577 , n15262 , n15310 );
    and g7867 ( n13505 , n22816 , n23576 );
    nor g7868 ( n8198 , n22651 , n6385 );
    and g7869 ( n11355 , n5774 , n960 );
    xnor g7870 ( n1304 , n7717 , n26313 );
    or g7871 ( n3560 , n6776 , n17917 );
    and g7872 ( n22005 , n4048 , n14433 );
    nor g7873 ( n26988 , n7871 , n8261 );
    or g7874 ( n20381 , n6592 , n19349 );
    not g7875 ( n12377 , n6730 );
    or g7876 ( n7370 , n16854 , n26143 );
    xnor g7877 ( n11391 , n2679 , n25592 );
    xnor g7878 ( n19455 , n6381 , n16376 );
    and g7879 ( n8368 , n25622 , n11945 );
    xnor g7880 ( n25476 , n16948 , n6379 );
    xnor g7881 ( n8950 , n9832 , n3959 );
    xnor g7882 ( n17410 , n11068 , n25474 );
    xnor g7883 ( n7146 , n10107 , n12507 );
    or g7884 ( n26869 , n12451 , n26880 );
    or g7885 ( n6475 , n20409 , n429 );
    or g7886 ( n9739 , n18032 , n9440 );
    xnor g7887 ( n5767 , n25965 , n9808 );
    not g7888 ( n17846 , n5555 );
    and g7889 ( n22067 , n5618 , n12786 );
    and g7890 ( n21184 , n9844 , n16579 );
    or g7891 ( n24640 , n13515 , n23961 );
    buf g7892 ( n7817 , n21858 );
    not g7893 ( n3241 , n7759 );
    or g7894 ( n24520 , n2717 , n10337 );
    nor g7895 ( n8053 , n9412 , n17567 );
    and g7896 ( n17150 , n328 , n15695 );
    nor g7897 ( n26513 , n15427 , n16521 );
    xnor g7898 ( n17931 , n15754 , n3810 );
    or g7899 ( n14546 , n8908 , n10047 );
    xnor g7900 ( n20116 , n21596 , n6352 );
    or g7901 ( n23177 , n7870 , n24759 );
    or g7902 ( n18458 , n24290 , n6526 );
    xnor g7903 ( n2303 , n9476 , n94 );
    xnor g7904 ( n12271 , n8910 , n22392 );
    or g7905 ( n12089 , n3801 , n20440 );
    xor g7906 ( n19483 , n22349 , n15743 );
    xnor g7907 ( n18661 , n3659 , n17635 );
    nor g7908 ( n2079 , n17366 , n14754 );
    xnor g7909 ( n11089 , n18964 , n20397 );
    xnor g7910 ( n25302 , n4644 , n4933 );
    or g7911 ( n21332 , n11880 , n24218 );
    not g7912 ( n26187 , n24536 );
    not g7913 ( n19112 , n12501 );
    nor g7914 ( n25512 , n56 , n4095 );
    or g7915 ( n22214 , n11827 , n16471 );
    or g7916 ( n22277 , n8156 , n24178 );
    and g7917 ( n26304 , n10461 , n10132 );
    and g7918 ( n25543 , n12181 , n14676 );
    xnor g7919 ( n23381 , n4878 , n12692 );
    xnor g7920 ( n16382 , n3823 , n21599 );
    not g7921 ( n14007 , n23913 );
    or g7922 ( n14035 , n11707 , n20926 );
    not g7923 ( n2235 , n5196 );
    not g7924 ( n22477 , n9806 );
    and g7925 ( n6909 , n9660 , n10515 );
    xnor g7926 ( n22872 , n5582 , n9717 );
    and g7927 ( n13418 , n4960 , n11427 );
    xnor g7928 ( n15762 , n17574 , n8335 );
    xnor g7929 ( n26939 , n23345 , n5381 );
    not g7930 ( n13429 , n23731 );
    not g7931 ( n4729 , n16824 );
    not g7932 ( n20124 , n9245 );
    or g7933 ( n206 , n14538 , n23862 );
    and g7934 ( n1947 , n7034 , n20573 );
    xnor g7935 ( n6745 , n21014 , n9004 );
    not g7936 ( n15498 , n15170 );
    xnor g7937 ( n3924 , n3019 , n1279 );
    xnor g7938 ( n9427 , n26443 , n10017 );
    or g7939 ( n18349 , n19575 , n16126 );
    not g7940 ( n26470 , n16968 );
    nor g7941 ( n17355 , n27144 , n6774 );
    not g7942 ( n20 , n19951 );
    xnor g7943 ( n23420 , n15167 , n919 );
    xnor g7944 ( n12463 , n20811 , n3909 );
    xnor g7945 ( n15297 , n16609 , n2886 );
    and g7946 ( n5870 , n10237 , n23846 );
    and g7947 ( n10011 , n16643 , n24110 );
    and g7948 ( n17101 , n10135 , n24863 );
    or g7949 ( n25492 , n11303 , n2429 );
    or g7950 ( n24295 , n26138 , n17340 );
    nor g7951 ( n20572 , n22977 , n23513 );
    xnor g7952 ( n18497 , n3346 , n19311 );
    xnor g7953 ( n22394 , n23353 , n14881 );
    or g7954 ( n4701 , n26658 , n19911 );
    or g7955 ( n20081 , n16755 , n18812 );
    xnor g7956 ( n11818 , n18248 , n16844 );
    xnor g7957 ( n11299 , n9990 , n18097 );
    xnor g7958 ( n22662 , n21494 , n16074 );
    or g7959 ( n12594 , n18838 , n1484 );
    xnor g7960 ( n12476 , n20954 , n21263 );
    or g7961 ( n5029 , n25258 , n6838 );
    nor g7962 ( n22131 , n22191 , n12064 );
    not g7963 ( n2894 , n22272 );
    not g7964 ( n16712 , n15539 );
    xnor g7965 ( n11648 , n7924 , n4767 );
    not g7966 ( n1987 , n14257 );
    not g7967 ( n17578 , n3211 );
    xnor g7968 ( n1703 , n25618 , n16829 );
    not g7969 ( n23670 , n4601 );
    or g7970 ( n3989 , n12603 , n11983 );
    and g7971 ( n26378 , n4843 , n872 );
    or g7972 ( n7998 , n21108 , n8073 );
    and g7973 ( n14075 , n11263 , n1538 );
    nor g7974 ( n2689 , n26180 , n10650 );
    xnor g7975 ( n22835 , n12911 , n26264 );
    not g7976 ( n16889 , n23166 );
    or g7977 ( n22956 , n6421 , n23674 );
    nor g7978 ( n25387 , n13244 , n3462 );
    nor g7979 ( n2404 , n20053 , n23876 );
    and g7980 ( n11061 , n559 , n11705 );
    nor g7981 ( n24478 , n15291 , n13401 );
    or g7982 ( n4411 , n17542 , n4409 );
    or g7983 ( n6409 , n24469 , n9447 );
    xnor g7984 ( n13093 , n27005 , n27188 );
    xnor g7985 ( n18538 , n26882 , n19618 );
    xnor g7986 ( n22829 , n2320 , n11736 );
    nor g7987 ( n12093 , n1798 , n8930 );
    not g7988 ( n8167 , n14488 );
    xnor g7989 ( n22154 , n22932 , n10316 );
    or g7990 ( n7986 , n22238 , n9036 );
    not g7991 ( n14139 , n23773 );
    or g7992 ( n13414 , n26691 , n20036 );
    xnor g7993 ( n13949 , n16994 , n9246 );
    and g7994 ( n1612 , n6337 , n3686 );
    or g7995 ( n11786 , n10207 , n18833 );
    xnor g7996 ( n3264 , n1662 , n7330 );
    and g7997 ( n26778 , n3366 , n4753 );
    xnor g7998 ( n23899 , n14296 , n23374 );
    or g7999 ( n11219 , n18257 , n23098 );
    or g8000 ( n6530 , n20407 , n25093 );
    xnor g8001 ( n4049 , n10822 , n18462 );
    or g8002 ( n16198 , n12414 , n16390 );
    or g8003 ( n484 , n25548 , n3323 );
    or g8004 ( n14676 , n8757 , n25383 );
    and g8005 ( n18730 , n11786 , n6384 );
    nor g8006 ( n4996 , n5960 , n9942 );
    xnor g8007 ( n24569 , n8491 , n23895 );
    and g8008 ( n10434 , n11466 , n2393 );
    xnor g8009 ( n23235 , n16414 , n3902 );
    and g8010 ( n5679 , n26106 , n23324 );
    nor g8011 ( n6042 , n3740 , n3498 );
    or g8012 ( n20332 , n16743 , n24485 );
    xnor g8013 ( n24634 , n1594 , n16602 );
    or g8014 ( n3111 , n2953 , n10681 );
    xnor g8015 ( n16951 , n20164 , n23299 );
    and g8016 ( n1369 , n8755 , n22923 );
    xnor g8017 ( n17220 , n7081 , n17597 );
    and g8018 ( n20871 , n26529 , n3939 );
    xnor g8019 ( n11103 , n12400 , n14534 );
    or g8020 ( n3310 , n16162 , n693 );
    or g8021 ( n10356 , n18936 , n13483 );
    xnor g8022 ( n12057 , n4995 , n24327 );
    and g8023 ( n18233 , n5913 , n4737 );
    xnor g8024 ( n7999 , n14877 , n26359 );
    nor g8025 ( n21664 , n4397 , n26178 );
    or g8026 ( n9410 , n21177 , n21534 );
    and g8027 ( n25093 , n4192 , n15619 );
    not g8028 ( n6713 , n21945 );
    xnor g8029 ( n7554 , n8171 , n4060 );
    nor g8030 ( n24428 , n2036 , n8434 );
    xnor g8031 ( n27110 , n21546 , n17922 );
    or g8032 ( n18122 , n17339 , n15564 );
    not g8033 ( n1467 , n14544 );
    xnor g8034 ( n1429 , n22495 , n3789 );
    buf g8035 ( n1319 , n24692 );
    or g8036 ( n15567 , n15631 , n4 );
    xnor g8037 ( n1807 , n14990 , n18526 );
    xnor g8038 ( n2678 , n9040 , n7769 );
    nor g8039 ( n5763 , n16889 , n4306 );
    xnor g8040 ( n2461 , n810 , n23694 );
    buf g8041 ( n21272 , n1674 );
    or g8042 ( n21880 , n9363 , n23044 );
    not g8043 ( n21117 , n26510 );
    and g8044 ( n4058 , n18100 , n16231 );
    xnor g8045 ( n3834 , n26152 , n21262 );
    or g8046 ( n16436 , n10275 , n22359 );
    or g8047 ( n9916 , n5989 , n15471 );
    and g8048 ( n21179 , n19140 , n17148 );
    not g8049 ( n15042 , n10625 );
    nor g8050 ( n7528 , n7270 , n16902 );
    not g8051 ( n599 , n14693 );
    or g8052 ( n13780 , n12445 , n19255 );
    xnor g8053 ( n24261 , n11246 , n26510 );
    xnor g8054 ( n1053 , n15998 , n9723 );
    nor g8055 ( n13016 , n5750 , n19884 );
    xnor g8056 ( n8756 , n20011 , n5697 );
    xnor g8057 ( n15570 , n12944 , n12614 );
    or g8058 ( n21068 , n13529 , n14720 );
    or g8059 ( n16242 , n22158 , n8717 );
    or g8060 ( n2814 , n13263 , n22596 );
    or g8061 ( n4147 , n11108 , n7327 );
    and g8062 ( n26148 , n23398 , n8183 );
    not g8063 ( n16711 , n22660 );
    xnor g8064 ( n11965 , n26238 , n24259 );
    xnor g8065 ( n11463 , n10485 , n7670 );
    xnor g8066 ( n22124 , n11211 , n17627 );
    not g8067 ( n18485 , n19514 );
    xnor g8068 ( n26414 , n12763 , n3740 );
    and g8069 ( n5699 , n7251 , n26057 );
    or g8070 ( n23646 , n9290 , n196 );
    or g8071 ( n22499 , n5465 , n11537 );
    xnor g8072 ( n16764 , n16637 , n2776 );
    xnor g8073 ( n1602 , n24527 , n12226 );
    nor g8074 ( n19172 , n26689 , n22666 );
    or g8075 ( n4568 , n20667 , n21927 );
    or g8076 ( n9171 , n3402 , n18440 );
    not g8077 ( n25627 , n12749 );
    not g8078 ( n17888 , n5800 );
    xnor g8079 ( n8913 , n6218 , n19652 );
    or g8080 ( n19645 , n18453 , n21657 );
    xnor g8081 ( n22998 , n11864 , n10279 );
    and g8082 ( n25027 , n14822 , n2074 );
    or g8083 ( n7427 , n3363 , n18506 );
    not g8084 ( n7957 , n18941 );
    or g8085 ( n21904 , n8344 , n6794 );
    not g8086 ( n12932 , n19327 );
    not g8087 ( n11938 , n21226 );
    and g8088 ( n4538 , n22696 , n18167 );
    not g8089 ( n6503 , n592 );
    not g8090 ( n19119 , n18792 );
    xnor g8091 ( n20696 , n26496 , n1621 );
    or g8092 ( n19504 , n22133 , n14598 );
    xnor g8093 ( n22450 , n7249 , n5182 );
    xnor g8094 ( n8089 , n26584 , n12204 );
    not g8095 ( n16252 , n4306 );
    or g8096 ( n19822 , n16482 , n13333 );
    not g8097 ( n5440 , n14148 );
    not g8098 ( n22194 , n3945 );
    or g8099 ( n16554 , n7151 , n21427 );
    not g8100 ( n14500 , n18827 );
    and g8101 ( n13997 , n25425 , n20368 );
    or g8102 ( n3910 , n21995 , n25789 );
    or g8103 ( n18627 , n2259 , n10991 );
    or g8104 ( n15283 , n19095 , n4783 );
    or g8105 ( n11687 , n6394 , n9273 );
    xnor g8106 ( n18959 , n11056 , n18157 );
    xnor g8107 ( n7797 , n14732 , n10965 );
    or g8108 ( n2972 , n104 , n20927 );
    or g8109 ( n21588 , n15079 , n5752 );
    nor g8110 ( n18296 , n24704 , n5728 );
    and g8111 ( n23914 , n25972 , n3707 );
    xnor g8112 ( n14252 , n21502 , n4017 );
    or g8113 ( n19808 , n6523 , n14298 );
    xnor g8114 ( n2667 , n25515 , n27066 );
    nor g8115 ( n13332 , n26565 , n20437 );
    or g8116 ( n23963 , n4658 , n11442 );
    or g8117 ( n19288 , n3349 , n12762 );
    or g8118 ( n9862 , n22059 , n25723 );
    nor g8119 ( n18381 , n13231 , n27115 );
    not g8120 ( n8529 , n15264 );
    or g8121 ( n14911 , n22291 , n6874 );
    nor g8122 ( n22024 , n15884 , n25602 );
    and g8123 ( n938 , n9688 , n22466 );
    xnor g8124 ( n20849 , n8508 , n12153 );
    or g8125 ( n9408 , n22523 , n24698 );
    and g8126 ( n3650 , n89 , n10396 );
    and g8127 ( n24207 , n4084 , n26051 );
    or g8128 ( n7800 , n13657 , n15941 );
    not g8129 ( n15734 , n9077 );
    xnor g8130 ( n25855 , n1032 , n19877 );
    and g8131 ( n27113 , n24355 , n1267 );
    xnor g8132 ( n8763 , n22723 , n5692 );
    xnor g8133 ( n4152 , n10857 , n8133 );
    xnor g8134 ( n6078 , n329 , n21735 );
    or g8135 ( n14368 , n382 , n10812 );
    not g8136 ( n19755 , n1853 );
    or g8137 ( n11450 , n12040 , n21459 );
    xnor g8138 ( n17956 , n9579 , n956 );
    not g8139 ( n4549 , n313 );
    xnor g8140 ( n10869 , n11835 , n9179 );
    or g8141 ( n17750 , n1537 , n13246 );
    nor g8142 ( n7017 , n26046 , n23512 );
    nor g8143 ( n22252 , n9631 , n18300 );
    and g8144 ( n200 , n2422 , n1562 );
    nor g8145 ( n4248 , n22346 , n23033 );
    and g8146 ( n9156 , n6050 , n14898 );
    or g8147 ( n16145 , n23752 , n26078 );
    not g8148 ( n19030 , n9485 );
    not g8149 ( n1941 , n15210 );
    or g8150 ( n22231 , n13577 , n11944 );
    or g8151 ( n24236 , n2915 , n23559 );
    xnor g8152 ( n13038 , n7380 , n24191 );
    xnor g8153 ( n9375 , n13359 , n7057 );
    or g8154 ( n429 , n25749 , n18507 );
    or g8155 ( n5576 , n23489 , n6733 );
    nor g8156 ( n23629 , n17423 , n19914 );
    nor g8157 ( n18192 , n17505 , n5465 );
    xnor g8158 ( n19478 , n23052 , n17038 );
    or g8159 ( n9275 , n10008 , n13460 );
    xnor g8160 ( n25209 , n3237 , n2695 );
    not g8161 ( n25967 , n847 );
    xnor g8162 ( n5428 , n2490 , n20447 );
    xnor g8163 ( n22537 , n18044 , n5383 );
    xnor g8164 ( n21159 , n19702 , n23849 );
    xnor g8165 ( n21358 , n10204 , n16158 );
    and g8166 ( n24386 , n1382 , n4252 );
    xnor g8167 ( n22640 , n16450 , n18926 );
    xnor g8168 ( n15170 , n9008 , n23505 );
    and g8169 ( n14372 , n9008 , n16145 );
    xnor g8170 ( n23410 , n4333 , n8869 );
    xnor g8171 ( n4972 , n26938 , n732 );
    and g8172 ( n3965 , n17915 , n26049 );
    xnor g8173 ( n1047 , n7493 , n11860 );
    and g8174 ( n15032 , n24250 , n22263 );
    not g8175 ( n4194 , n15408 );
    or g8176 ( n16827 , n524 , n24947 );
    nor g8177 ( n7942 , n1365 , n19234 );
    or g8178 ( n7920 , n9637 , n13680 );
    nor g8179 ( n12109 , n18003 , n26013 );
    nor g8180 ( n16747 , n13459 , n1689 );
    not g8181 ( n1916 , n10344 );
    or g8182 ( n9045 , n21957 , n14410 );
    or g8183 ( n21318 , n4833 , n24221 );
    nor g8184 ( n26451 , n9883 , n11016 );
    not g8185 ( n13245 , n5307 );
    and g8186 ( n9932 , n23762 , n2053 );
    not g8187 ( n2086 , n3849 );
    and g8188 ( n4641 , n8125 , n2550 );
    xor g8189 ( n6430 , n6122 , n19196 );
    and g8190 ( n24497 , n25028 , n10871 );
    xnor g8191 ( n20403 , n18470 , n10793 );
    or g8192 ( n12757 , n692 , n1991 );
    xnor g8193 ( n20389 , n7803 , n21630 );
    or g8194 ( n15279 , n10751 , n14466 );
    or g8195 ( n17736 , n7517 , n1026 );
    and g8196 ( n17989 , n6715 , n3159 );
    or g8197 ( n4627 , n25043 , n17901 );
    or g8198 ( n8124 , n23758 , n10361 );
    not g8199 ( n2935 , n16051 );
    and g8200 ( n2876 , n25306 , n8038 );
    nor g8201 ( n11643 , n11597 , n12888 );
    not g8202 ( n3677 , n921 );
    xnor g8203 ( n9608 , n10608 , n12587 );
    xnor g8204 ( n11712 , n16463 , n16258 );
    xnor g8205 ( n16460 , n16710 , n11801 );
    and g8206 ( n21289 , n15820 , n21824 );
    and g8207 ( n19564 , n13076 , n17492 );
    or g8208 ( n17283 , n15928 , n8444 );
    and g8209 ( n11885 , n4801 , n11970 );
    nor g8210 ( n399 , n5128 , n22926 );
    xnor g8211 ( n314 , n22764 , n2416 );
    xnor g8212 ( n15794 , n23166 , n18105 );
    or g8213 ( n15449 , n3503 , n1875 );
    xnor g8214 ( n8997 , n17294 , n335 );
    nor g8215 ( n20303 , n2909 , n19312 );
    and g8216 ( n5339 , n18938 , n19957 );
    or g8217 ( n6823 , n3586 , n1285 );
    and g8218 ( n4279 , n16514 , n21825 );
    xnor g8219 ( n26375 , n19434 , n26965 );
    xnor g8220 ( n21309 , n25960 , n1102 );
    xnor g8221 ( n22249 , n11229 , n17195 );
    or g8222 ( n7847 , n4304 , n23876 );
    and g8223 ( n15736 , n2268 , n19153 );
    xnor g8224 ( n21458 , n15478 , n7369 );
    not g8225 ( n18506 , n19228 );
    not g8226 ( n12366 , n18183 );
    or g8227 ( n21395 , n14936 , n15233 );
    xnor g8228 ( n175 , n18772 , n17654 );
    or g8229 ( n4244 , n26465 , n9758 );
    or g8230 ( n9385 , n6438 , n6473 );
    and g8231 ( n3315 , n12400 , n2966 );
    and g8232 ( n2797 , n25778 , n3134 );
    xnor g8233 ( n7580 , n12351 , n14323 );
    or g8234 ( n6512 , n8746 , n620 );
    xnor g8235 ( n10746 , n1978 , n22884 );
    xnor g8236 ( n7053 , n26299 , n25208 );
    or g8237 ( n4234 , n690 , n13036 );
    or g8238 ( n13838 , n26557 , n4670 );
    xnor g8239 ( n6185 , n25595 , n909 );
    or g8240 ( n10118 , n25891 , n2312 );
    or g8241 ( n23519 , n6253 , n20664 );
    xnor g8242 ( n26135 , n4465 , n10271 );
    or g8243 ( n338 , n5211 , n21832 );
    not g8244 ( n12990 , n11589 );
    xnor g8245 ( n13123 , n12436 , n19475 );
    xnor g8246 ( n23986 , n16044 , n8113 );
    not g8247 ( n1262 , n21832 );
    or g8248 ( n13471 , n9027 , n22112 );
    or g8249 ( n1032 , n22151 , n10960 );
    or g8250 ( n9729 , n8713 , n6071 );
    not g8251 ( n2261 , n23285 );
    or g8252 ( n20606 , n3937 , n1243 );
    nor g8253 ( n3248 , n1946 , n6648 );
    not g8254 ( n17806 , n13452 );
    and g8255 ( n5570 , n20453 , n1361 );
    or g8256 ( n8839 , n1829 , n15371 );
    nor g8257 ( n10494 , n2145 , n22021 );
    or g8258 ( n179 , n24050 , n25737 );
    xnor g8259 ( n7131 , n3374 , n27101 );
    and g8260 ( n25127 , n9623 , n3262 );
    not g8261 ( n25726 , n5072 );
    xnor g8262 ( n3686 , n6261 , n19685 );
    and g8263 ( n25121 , n19358 , n25302 );
    and g8264 ( n18266 , n15827 , n15073 );
    and g8265 ( n16510 , n5730 , n4825 );
    and g8266 ( n6931 , n2577 , n4421 );
    nor g8267 ( n22291 , n12396 , n20064 );
    or g8268 ( n20805 , n2187 , n2161 );
    or g8269 ( n12253 , n21886 , n2983 );
    not g8270 ( n14244 , n7833 );
    xnor g8271 ( n20757 , n25345 , n9967 );
    nor g8272 ( n18788 , n15636 , n18255 );
    or g8273 ( n3816 , n16497 , n6848 );
    nor g8274 ( n2957 , n7755 , n21097 );
    not g8275 ( n10802 , n13468 );
    and g8276 ( n784 , n14218 , n7737 );
    and g8277 ( n5747 , n17041 , n25626 );
    or g8278 ( n6937 , n23623 , n5412 );
    and g8279 ( n1368 , n20983 , n18082 );
    and g8280 ( n13800 , n20527 , n2525 );
    xnor g8281 ( n21446 , n25205 , n20356 );
    xnor g8282 ( n9152 , n10314 , n10242 );
    xor g8283 ( n21441 , n26912 , n13038 );
    or g8284 ( n12290 , n16355 , n11371 );
    xnor g8285 ( n19602 , n24168 , n8271 );
    or g8286 ( n1134 , n20826 , n14532 );
    or g8287 ( n9785 , n7914 , n17767 );
    not g8288 ( n19944 , n26979 );
    not g8289 ( n6833 , n23039 );
    xnor g8290 ( n25831 , n13492 , n16536 );
    nor g8291 ( n20853 , n23990 , n16960 );
    and g8292 ( n21122 , n3145 , n10453 );
    nor g8293 ( n275 , n23408 , n22660 );
    or g8294 ( n17107 , n1540 , n13424 );
    xnor g8295 ( n1523 , n4576 , n17302 );
    nor g8296 ( n18591 , n570 , n16211 );
    or g8297 ( n16187 , n7065 , n18480 );
    or g8298 ( n22825 , n26890 , n24117 );
    nor g8299 ( n19865 , n3823 , n12262 );
    or g8300 ( n12915 , n25204 , n19309 );
    xnor g8301 ( n692 , n4422 , n10442 );
    nor g8302 ( n5295 , n20228 , n8717 );
    or g8303 ( n11563 , n14736 , n21226 );
    xnor g8304 ( n8674 , n5122 , n19976 );
    and g8305 ( n1071 , n18957 , n21660 );
    not g8306 ( n4673 , n11810 );
    and g8307 ( n12347 , n9295 , n15786 );
    not g8308 ( n10986 , n3651 );
    or g8309 ( n13181 , n22216 , n539 );
    nor g8310 ( n24397 , n7756 , n20683 );
    or g8311 ( n3782 , n5169 , n2085 );
    and g8312 ( n2098 , n21649 , n17846 );
    nor g8313 ( n13131 , n19701 , n7437 );
    xnor g8314 ( n6544 , n23529 , n10739 );
    or g8315 ( n11520 , n12609 , n6954 );
    or g8316 ( n23440 , n6834 , n5165 );
    and g8317 ( n19859 , n22419 , n20390 );
    xnor g8318 ( n14944 , n3133 , n4379 );
    and g8319 ( n7815 , n15541 , n16043 );
    or g8320 ( n17441 , n13588 , n16318 );
    or g8321 ( n8243 , n18355 , n21822 );
    xnor g8322 ( n1895 , n26716 , n16301 );
    xnor g8323 ( n16366 , n11654 , n8006 );
    not g8324 ( n18318 , n3471 );
    and g8325 ( n14109 , n16968 , n27189 );
    xnor g8326 ( n22716 , n13896 , n4661 );
    or g8327 ( n19786 , n23015 , n24754 );
    or g8328 ( n7336 , n25369 , n21329 );
    not g8329 ( n20056 , n4877 );
    or g8330 ( n15824 , n1558 , n5050 );
    or g8331 ( n20154 , n21792 , n1478 );
    and g8332 ( n10826 , n5226 , n11223 );
    nor g8333 ( n3351 , n9076 , n24805 );
    or g8334 ( n5994 , n3568 , n18202 );
    xnor g8335 ( n18812 , n18918 , n11787 );
    not g8336 ( n16313 , n23833 );
    or g8337 ( n3313 , n8568 , n1600 );
    or g8338 ( n15933 , n11554 , n25521 );
    and g8339 ( n9871 , n7728 , n1699 );
    or g8340 ( n10862 , n21868 , n7892 );
    or g8341 ( n7512 , n1762 , n711 );
    not g8342 ( n19632 , n18314 );
    or g8343 ( n15600 , n11503 , n18151 );
    not g8344 ( n26508 , n15761 );
    nor g8345 ( n12718 , n13650 , n14025 );
    or g8346 ( n19156 , n22426 , n12543 );
    xnor g8347 ( n8130 , n3328 , n14970 );
    or g8348 ( n8627 , n21777 , n4685 );
    xnor g8349 ( n7523 , n23556 , n27089 );
    or g8350 ( n16780 , n13953 , n17511 );
    nor g8351 ( n4241 , n2453 , n22492 );
    and g8352 ( n16850 , n1492 , n6077 );
    or g8353 ( n19124 , n25273 , n25777 );
    xnor g8354 ( n3725 , n9902 , n10913 );
    buf g8355 ( n19731 , n23104 );
    xnor g8356 ( n21472 , n19810 , n12273 );
    or g8357 ( n26361 , n14518 , n18806 );
    or g8358 ( n8007 , n16364 , n15495 );
    or g8359 ( n7322 , n8094 , n5580 );
    xnor g8360 ( n6476 , n69 , n11593 );
    not g8361 ( n8003 , n15643 );
    and g8362 ( n22114 , n17013 , n7799 );
    nor g8363 ( n19209 , n12009 , n10259 );
    or g8364 ( n13771 , n5077 , n13914 );
    and g8365 ( n7342 , n12513 , n8162 );
    or g8366 ( n20007 , n18894 , n5186 );
    xnor g8367 ( n27108 , n161 , n12780 );
    xnor g8368 ( n19834 , n19236 , n21930 );
    or g8369 ( n14588 , n744 , n9363 );
    xnor g8370 ( n18238 , n4394 , n672 );
    nor g8371 ( n15334 , n4201 , n3045 );
    xnor g8372 ( n3555 , n22966 , n24722 );
    xnor g8373 ( n17600 , n16069 , n21673 );
    and g8374 ( n10313 , n407 , n9717 );
    and g8375 ( n14901 , n4034 , n15208 );
    not g8376 ( n10424 , n665 );
    and g8377 ( n26575 , n3309 , n23177 );
    xnor g8378 ( n8335 , n6731 , n7347 );
    and g8379 ( n23459 , n4177 , n19482 );
    and g8380 ( n17795 , n15318 , n7758 );
    not g8381 ( n26747 , n21687 );
    or g8382 ( n1098 , n4132 , n24301 );
    not g8383 ( n25015 , n18125 );
    or g8384 ( n12482 , n16743 , n5194 );
    or g8385 ( n1638 , n9165 , n11319 );
    nor g8386 ( n9925 , n22472 , n9125 );
    and g8387 ( n1115 , n8333 , n7908 );
    nor g8388 ( n15799 , n3681 , n18383 );
    and g8389 ( n9188 , n17512 , n9606 );
    xnor g8390 ( n7518 , n5374 , n23002 );
    nor g8391 ( n26423 , n17663 , n22862 );
    or g8392 ( n25638 , n26845 , n3790 );
    and g8393 ( n22152 , n1462 , n20007 );
    and g8394 ( n13162 , n9378 , n10833 );
    and g8395 ( n13462 , n13531 , n9745 );
    xnor g8396 ( n17563 , n10467 , n593 );
    not g8397 ( n12022 , n19646 );
    or g8398 ( n2648 , n6305 , n9197 );
    not g8399 ( n18754 , n15910 );
    xnor g8400 ( n10873 , n11726 , n8401 );
    nor g8401 ( n14117 , n2915 , n8363 );
    xnor g8402 ( n20302 , n19327 , n21934 );
    and g8403 ( n18219 , n10156 , n26782 );
    and g8404 ( n18084 , n838 , n10676 );
    or g8405 ( n877 , n13103 , n14321 );
    xnor g8406 ( n13455 , n11988 , n17880 );
    or g8407 ( n19790 , n26875 , n18487 );
    xnor g8408 ( n10355 , n13693 , n12650 );
    and g8409 ( n13013 , n4278 , n15074 );
    or g8410 ( n13600 , n22365 , n15359 );
    nor g8411 ( n11513 , n21317 , n19196 );
    not g8412 ( n18867 , n16078 );
    not g8413 ( n25704 , n23653 );
    not g8414 ( n20513 , n19540 );
    or g8415 ( n15621 , n1356 , n13341 );
    xnor g8416 ( n551 , n13231 , n27115 );
    or g8417 ( n9186 , n5113 , n5283 );
    or g8418 ( n4323 , n19304 , n15497 );
    or g8419 ( n3331 , n12534 , n3004 );
    not g8420 ( n20260 , n80 );
    xnor g8421 ( n20458 , n11958 , n11483 );
    not g8422 ( n10571 , n23213 );
    or g8423 ( n10883 , n21471 , n19357 );
    xnor g8424 ( n8135 , n9092 , n13877 );
    and g8425 ( n7600 , n25946 , n12512 );
    or g8426 ( n22803 , n24200 , n14648 );
    and g8427 ( n18541 , n7600 , n16757 );
    xnor g8428 ( n24951 , n26995 , n11658 );
    nor g8429 ( n11166 , n16294 , n2160 );
    xnor g8430 ( n3932 , n11660 , n11512 );
    not g8431 ( n17803 , n19691 );
    or g8432 ( n4541 , n846 , n8407 );
    or g8433 ( n23522 , n22083 , n1304 );
    or g8434 ( n26389 , n3510 , n21523 );
    xnor g8435 ( n24616 , n4635 , n857 );
    or g8436 ( n14644 , n22763 , n26865 );
    or g8437 ( n9882 , n23063 , n11486 );
    xnor g8438 ( n22241 , n26919 , n11322 );
    and g8439 ( n20238 , n17644 , n8924 );
    xnor g8440 ( n7032 , n12629 , n23212 );
    or g8441 ( n5972 , n5512 , n27071 );
    nor g8442 ( n522 , n20937 , n424 );
    xnor g8443 ( n9192 , n22254 , n22699 );
    not g8444 ( n12090 , n6819 );
    not g8445 ( n23905 , n23318 );
    xnor g8446 ( n12620 , n16151 , n18898 );
    xnor g8447 ( n18886 , n7723 , n25892 );
    or g8448 ( n9656 , n20077 , n6794 );
    nor g8449 ( n1918 , n9680 , n7364 );
    or g8450 ( n13083 , n12789 , n23218 );
    and g8451 ( n20876 , n6018 , n10099 );
    xnor g8452 ( n18692 , n330 , n5668 );
    xnor g8453 ( n24298 , n6224 , n11696 );
    nor g8454 ( n12728 , n2308 , n2489 );
    xnor g8455 ( n24537 , n2381 , n22377 );
    xnor g8456 ( n26923 , n20834 , n16273 );
    or g8457 ( n4581 , n26053 , n25461 );
    xnor g8458 ( n12873 , n18233 , n15535 );
    not g8459 ( n24364 , n27146 );
    nor g8460 ( n2106 , n25877 , n10057 );
    or g8461 ( n21387 , n5363 , n9328 );
    nor g8462 ( n86 , n3094 , n2191 );
    or g8463 ( n23367 , n24273 , n14630 );
    or g8464 ( n3395 , n14718 , n23705 );
    xnor g8465 ( n15230 , n13286 , n8514 );
    xnor g8466 ( n20973 , n5179 , n129 );
    or g8467 ( n26736 , n16135 , n9168 );
    nor g8468 ( n7666 , n25240 , n20707 );
    and g8469 ( n9706 , n328 , n19387 );
    and g8470 ( n12927 , n17522 , n9410 );
    or g8471 ( n3449 , n1432 , n12040 );
    or g8472 ( n27016 , n20952 , n20262 );
    or g8473 ( n8916 , n8677 , n15146 );
    nor g8474 ( n26358 , n910 , n12891 );
    or g8475 ( n25776 , n18861 , n693 );
    not g8476 ( n11834 , n22437 );
    or g8477 ( n18764 , n21016 , n23956 );
    or g8478 ( n3864 , n16565 , n11982 );
    or g8479 ( n19812 , n16452 , n26840 );
    xnor g8480 ( n21529 , n21798 , n23969 );
    xnor g8481 ( n5779 , n4062 , n16499 );
    buf g8482 ( n13037 , n10908 );
    and g8483 ( n15810 , n12602 , n24775 );
    nor g8484 ( n18088 , n22660 , n24774 );
    and g8485 ( n8264 , n18309 , n7433 );
    and g8486 ( n3689 , n26530 , n25465 );
    or g8487 ( n22564 , n20702 , n17774 );
    and g8488 ( n15798 , n17402 , n5691 );
    xnor g8489 ( n18940 , n22532 , n15548 );
    nor g8490 ( n26738 , n12650 , n13693 );
    xnor g8491 ( n8728 , n22410 , n15610 );
    and g8492 ( n12163 , n4730 , n14030 );
    xnor g8493 ( n9021 , n11578 , n7335 );
    and g8494 ( n17514 , n20728 , n1036 );
    or g8495 ( n19697 , n22652 , n6267 );
    not g8496 ( n10159 , n604 );
    nor g8497 ( n21257 , n21784 , n18163 );
    and g8498 ( n16804 , n5219 , n24454 );
    nor g8499 ( n487 , n18869 , n10741 );
    and g8500 ( n7813 , n22023 , n1017 );
    and g8501 ( n3700 , n8189 , n24994 );
    or g8502 ( n24906 , n7496 , n12151 );
    not g8503 ( n9067 , n16965 );
    not g8504 ( n18746 , n5098 );
    xnor g8505 ( n8837 , n18947 , n26797 );
    or g8506 ( n7201 , n17578 , n8653 );
    xnor g8507 ( n5167 , n26747 , n9380 );
    not g8508 ( n21392 , n11640 );
    not g8509 ( n2407 , n16803 );
    xnor g8510 ( n27067 , n19110 , n10522 );
    xnor g8511 ( n17074 , n13734 , n6019 );
    nor g8512 ( n17774 , n5919 , n3653 );
    and g8513 ( n2909 , n27117 , n13836 );
    not g8514 ( n25650 , n13851 );
    and g8515 ( n10377 , n9286 , n7629 );
    xnor g8516 ( n20198 , n16009 , n6397 );
    xnor g8517 ( n20029 , n19249 , n12884 );
    and g8518 ( n22284 , n18651 , n25307 );
    and g8519 ( n6529 , n26227 , n23101 );
    or g8520 ( n9634 , n20329 , n25464 );
    nor g8521 ( n16208 , n6502 , n1630 );
    and g8522 ( n19678 , n4581 , n3928 );
    xnor g8523 ( n12864 , n2716 , n18657 );
    not g8524 ( n10969 , n755 );
    and g8525 ( n19522 , n8373 , n18819 );
    and g8526 ( n1495 , n9528 , n13055 );
    xnor g8527 ( n8184 , n14872 , n11903 );
    xnor g8528 ( n25919 , n977 , n2858 );
    xnor g8529 ( n6031 , n9524 , n2788 );
    or g8530 ( n12833 , n23099 , n7402 );
    or g8531 ( n5670 , n22912 , n7484 );
    and g8532 ( n9519 , n13152 , n2688 );
    xnor g8533 ( n23897 , n5555 , n17323 );
    and g8534 ( n14907 , n4515 , n19136 );
    xnor g8535 ( n21234 , n25701 , n1204 );
    xnor g8536 ( n8416 , n14696 , n19552 );
    xnor g8537 ( n24791 , n12664 , n24196 );
    or g8538 ( n14093 , n17103 , n17795 );
    not g8539 ( n23592 , n14130 );
    and g8540 ( n10122 , n9735 , n2595 );
    not g8541 ( n25612 , n11701 );
    nor g8542 ( n2846 , n12929 , n16971 );
    and g8543 ( n12079 , n21273 , n4302 );
    not g8544 ( n2044 , n8728 );
    or g8545 ( n16699 , n8414 , n24617 );
    nor g8546 ( n1259 , n24620 , n22327 );
    xnor g8547 ( n13628 , n21322 , n19531 );
    xnor g8548 ( n8774 , n5133 , n2421 );
    or g8549 ( n9676 , n18591 , n15726 );
    or g8550 ( n24938 , n21247 , n24458 );
    xnor g8551 ( n11578 , n3171 , n3425 );
    nor g8552 ( n9282 , n19360 , n12964 );
    xnor g8553 ( n1971 , n26295 , n16824 );
    and g8554 ( n11574 , n25600 , n24123 );
    xnor g8555 ( n8046 , n7460 , n22068 );
    and g8556 ( n9149 , n7377 , n21125 );
    not g8557 ( n2045 , n5226 );
    not g8558 ( n27002 , n2951 );
    xnor g8559 ( n22692 , n25419 , n17061 );
    and g8560 ( n15777 , n14672 , n2258 );
    nor g8561 ( n113 , n2980 , n12514 );
    nor g8562 ( n20842 , n21597 , n22722 );
    xnor g8563 ( n26431 , n14509 , n825 );
    not g8564 ( n21114 , n18395 );
    xnor g8565 ( n7829 , n5026 , n8581 );
    not g8566 ( n13767 , n24429 );
    xnor g8567 ( n7174 , n6063 , n17862 );
    xnor g8568 ( n3089 , n27198 , n15469 );
    and g8569 ( n14808 , n5724 , n2572 );
    or g8570 ( n651 , n26043 , n6665 );
    and g8571 ( n11618 , n24003 , n15472 );
    or g8572 ( n3954 , n7757 , n16962 );
    not g8573 ( n9273 , n231 );
    not g8574 ( n23898 , n6819 );
    or g8575 ( n26276 , n26329 , n4908 );
    or g8576 ( n13694 , n17066 , n22325 );
    xnor g8577 ( n1012 , n23417 , n9513 );
    xnor g8578 ( n3456 , n10138 , n25054 );
    not g8579 ( n23190 , n14256 );
    xnor g8580 ( n15359 , n14673 , n126 );
    xnor g8581 ( n26740 , n6501 , n20274 );
    or g8582 ( n11038 , n1195 , n21412 );
    xnor g8583 ( n7647 , n2983 , n17519 );
    xnor g8584 ( n4384 , n19048 , n9536 );
    not g8585 ( n2174 , n13460 );
    xnor g8586 ( n20582 , n19563 , n3189 );
    not g8587 ( n11924 , n8847 );
    or g8588 ( n26101 , n2376 , n6644 );
    not g8589 ( n8436 , n13660 );
    not g8590 ( n8682 , n1998 );
    not g8591 ( n7092 , n5296 );
    and g8592 ( n2526 , n12166 , n8346 );
    xnor g8593 ( n17166 , n17107 , n9228 );
    not g8594 ( n14395 , n10917 );
    or g8595 ( n13730 , n14965 , n25465 );
    or g8596 ( n7375 , n19944 , n24366 );
    xnor g8597 ( n17762 , n13481 , n454 );
    xnor g8598 ( n8293 , n1777 , n16029 );
    or g8599 ( n19891 , n9846 , n18099 );
    or g8600 ( n1144 , n25113 , n24839 );
    or g8601 ( n9367 , n4710 , n4526 );
    and g8602 ( n22701 , n9464 , n5294 );
    or g8603 ( n569 , n24786 , n1574 );
    and g8604 ( n855 , n10715 , n12517 );
    and g8605 ( n25089 , n16585 , n2751 );
    nor g8606 ( n18098 , n8745 , n7532 );
    and g8607 ( n7105 , n3923 , n12486 );
    and g8608 ( n26928 , n13264 , n17982 );
    and g8609 ( n301 , n23611 , n6512 );
    xnor g8610 ( n7962 , n13137 , n1288 );
    xnor g8611 ( n4165 , n5642 , n8731 );
    or g8612 ( n16629 , n20975 , n18817 );
    or g8613 ( n3566 , n10716 , n19132 );
    not g8614 ( n23118 , n14921 );
    nor g8615 ( n4462 , n17909 , n9172 );
    or g8616 ( n23335 , n13591 , n3164 );
    and g8617 ( n26355 , n4027 , n19065 );
    or g8618 ( n24384 , n24850 , n12921 );
    and g8619 ( n11323 , n26824 , n25761 );
    and g8620 ( n18118 , n23084 , n3870 );
    nor g8621 ( n1427 , n9957 , n6435 );
    not g8622 ( n15842 , n3405 );
    or g8623 ( n17319 , n8331 , n20176 );
    not g8624 ( n20535 , n22057 );
    xnor g8625 ( n18854 , n11451 , n19770 );
    xnor g8626 ( n10564 , n105 , n2920 );
    or g8627 ( n21039 , n10192 , n20335 );
    xnor g8628 ( n2366 , n22276 , n1113 );
    xnor g8629 ( n23292 , n6442 , n8959 );
    or g8630 ( n1474 , n2377 , n12246 );
    and g8631 ( n23442 , n465 , n24985 );
    or g8632 ( n14924 , n23880 , n15166 );
    nor g8633 ( n17908 , n5990 , n7326 );
    and g8634 ( n1761 , n5237 , n7443 );
    not g8635 ( n3383 , n22294 );
    or g8636 ( n26063 , n26307 , n23799 );
    xnor g8637 ( n9359 , n2664 , n11301 );
    or g8638 ( n18476 , n12016 , n23118 );
    xnor g8639 ( n7 , n11943 , n3369 );
    xnor g8640 ( n10482 , n11203 , n16978 );
    xnor g8641 ( n26885 , n6025 , n24788 );
    nor g8642 ( n10084 , n5043 , n24726 );
    or g8643 ( n7042 , n8784 , n17350 );
    and g8644 ( n17781 , n11495 , n17275 );
    xnor g8645 ( n23067 , n13957 , n23392 );
    xnor g8646 ( n22126 , n3209 , n26685 );
    not g8647 ( n16257 , n5255 );
    xnor g8648 ( n20061 , n20843 , n9879 );
    and g8649 ( n20018 , n16766 , n25174 );
    not g8650 ( n1325 , n15532 );
    or g8651 ( n15584 , n4318 , n5562 );
    nor g8652 ( n17252 , n20429 , n26054 );
    nor g8653 ( n2726 , n6222 , n990 );
    not g8654 ( n25954 , n5260 );
    xnor g8655 ( n8850 , n6681 , n10538 );
    not g8656 ( n5708 , n25813 );
    xor g8657 ( n6896 , n20127 , n23842 );
    or g8658 ( n5791 , n17251 , n7473 );
    not g8659 ( n23512 , n23900 );
    xnor g8660 ( n2760 , n25602 , n15884 );
    or g8661 ( n17503 , n24302 , n5238 );
    or g8662 ( n4104 , n18907 , n18951 );
    or g8663 ( n9144 , n5203 , n8297 );
    and g8664 ( n10976 , n19680 , n18341 );
    xnor g8665 ( n9672 , n16473 , n22597 );
    and g8666 ( n5809 , n641 , n14460 );
    xnor g8667 ( n21355 , n20290 , n9934 );
    xnor g8668 ( n10686 , n10075 , n15959 );
    xnor g8669 ( n24009 , n20823 , n5764 );
    and g8670 ( n2031 , n13508 , n7400 );
    xnor g8671 ( n19685 , n23807 , n26443 );
    xnor g8672 ( n12773 , n15633 , n8097 );
    nor g8673 ( n2287 , n11926 , n2090 );
    and g8674 ( n633 , n1248 , n18222 );
    and g8675 ( n24206 , n2216 , n22873 );
    nor g8676 ( n17726 , n18724 , n138 );
    xnor g8677 ( n16541 , n16715 , n13255 );
    or g8678 ( n25353 , n16521 , n7139 );
    xnor g8679 ( n5788 , n21104 , n6315 );
    not g8680 ( n10760 , n1446 );
    not g8681 ( n4878 , n26901 );
    xnor g8682 ( n2665 , n1618 , n17926 );
    and g8683 ( n5510 , n16167 , n173 );
    or g8684 ( n10339 , n7237 , n15087 );
    or g8685 ( n8188 , n12337 , n18388 );
    xnor g8686 ( n21603 , n16687 , n20906 );
    or g8687 ( n6675 , n10301 , n7001 );
    or g8688 ( n5720 , n26920 , n3913 );
    and g8689 ( n16047 , n12147 , n9485 );
    nor g8690 ( n16254 , n2906 , n14187 );
    not g8691 ( n2274 , n20570 );
    xnor g8692 ( n2596 , n10577 , n24196 );
    and g8693 ( n4629 , n21783 , n26863 );
    xnor g8694 ( n22138 , n537 , n21221 );
    not g8695 ( n4599 , n830 );
    and g8696 ( n8054 , n17268 , n20636 );
    nor g8697 ( n12822 , n8182 , n4659 );
    or g8698 ( n26666 , n10574 , n16266 );
    not g8699 ( n8520 , n7856 );
    or g8700 ( n20374 , n8676 , n4672 );
    xnor g8701 ( n21378 , n26223 , n10950 );
    and g8702 ( n18566 , n14638 , n11071 );
    and g8703 ( n7290 , n21867 , n19155 );
    nor g8704 ( n22518 , n9827 , n25799 );
    nor g8705 ( n9412 , n22071 , n18452 );
    and g8706 ( n5689 , n27142 , n2410 );
    or g8707 ( n23266 , n26217 , n3698 );
    or g8708 ( n25843 , n26972 , n9668 );
    xnor g8709 ( n13922 , n10951 , n15254 );
    and g8710 ( n19765 , n2780 , n24212 );
    nor g8711 ( n28 , n12754 , n2167 );
    xnor g8712 ( n644 , n2053 , n1503 );
    xnor g8713 ( n6628 , n14312 , n14451 );
    and g8714 ( n20800 , n22301 , n14183 );
    xnor g8715 ( n21021 , n6972 , n3161 );
    or g8716 ( n17659 , n19962 , n23793 );
    xnor g8717 ( n1593 , n2776 , n4853 );
    or g8718 ( n12425 , n26704 , n3358 );
    nor g8719 ( n2519 , n13378 , n2071 );
    xnor g8720 ( n15723 , n19154 , n13095 );
    or g8721 ( n5920 , n9818 , n7530 );
    or g8722 ( n13791 , n17099 , n15124 );
    xnor g8723 ( n3915 , n1897 , n7464 );
    nor g8724 ( n4309 , n3554 , n167 );
    not g8725 ( n12774 , n19737 );
    not g8726 ( n14273 , n14381 );
    or g8727 ( n11167 , n21565 , n6911 );
    and g8728 ( n11170 , n17862 , n6063 );
    and g8729 ( n8960 , n20820 , n16058 );
    nor g8730 ( n15149 , n20896 , n6435 );
    xnor g8731 ( n24202 , n22521 , n26913 );
    and g8732 ( n5893 , n469 , n25686 );
    and g8733 ( n3929 , n19945 , n26190 );
    xnor g8734 ( n21256 , n23084 , n3870 );
    xnor g8735 ( n20450 , n20038 , n20947 );
    or g8736 ( n5401 , n14899 , n10408 );
    and g8737 ( n25012 , n22801 , n21033 );
    and g8738 ( n23689 , n20078 , n6676 );
    not g8739 ( n21739 , n3217 );
    not g8740 ( n2336 , n11184 );
    and g8741 ( n7164 , n5393 , n7986 );
    xnor g8742 ( n1376 , n12513 , n8162 );
    and g8743 ( n20135 , n11906 , n14611 );
    xnor g8744 ( n20425 , n1221 , n16597 );
    or g8745 ( n4264 , n22606 , n21381 );
    or g8746 ( n17177 , n18200 , n19127 );
    xnor g8747 ( n10012 , n4326 , n12593 );
    or g8748 ( n19987 , n5267 , n14038 );
    not g8749 ( n6321 , n10017 );
    not g8750 ( n23966 , n21538 );
    or g8751 ( n11360 , n6638 , n6301 );
    xnor g8752 ( n8484 , n17090 , n20986 );
    or g8753 ( n22694 , n10152 , n1700 );
    xnor g8754 ( n11589 , n3195 , n12998 );
    xnor g8755 ( n24576 , n13528 , n17274 );
    not g8756 ( n23572 , n25540 );
    or g8757 ( n16270 , n11586 , n3214 );
    or g8758 ( n1366 , n5882 , n17064 );
    or g8759 ( n1921 , n14204 , n14783 );
    and g8760 ( n13618 , n2312 , n25891 );
    and g8761 ( n15022 , n10158 , n25004 );
    xnor g8762 ( n10779 , n3840 , n8925 );
    xnor g8763 ( n5552 , n26486 , n2858 );
    xnor g8764 ( n4975 , n11499 , n16458 );
    xnor g8765 ( n12126 , n17570 , n11239 );
    or g8766 ( n2307 , n12269 , n10069 );
    or g8767 ( n24070 , n23211 , n17758 );
    and g8768 ( n3784 , n18477 , n2060 );
    or g8769 ( n3592 , n12427 , n23523 );
    or g8770 ( n10842 , n1888 , n6817 );
    and g8771 ( n26496 , n25950 , n16706 );
    xnor g8772 ( n22381 , n24226 , n17412 );
    or g8773 ( n18091 , n3882 , n4112 );
    and g8774 ( n17566 , n15980 , n5083 );
    xnor g8775 ( n6684 , n20337 , n16925 );
    or g8776 ( n10030 , n13633 , n2675 );
    or g8777 ( n11692 , n15675 , n6956 );
    xnor g8778 ( n3978 , n15539 , n17664 );
    xnor g8779 ( n19533 , n23724 , n17854 );
    xnor g8780 ( n11242 , n8713 , n20417 );
    or g8781 ( n6100 , n25632 , n24399 );
    or g8782 ( n12181 , n9872 , n2801 );
    nor g8783 ( n5758 , n1630 , n11121 );
    and g8784 ( n11994 , n2831 , n16409 );
    or g8785 ( n25496 , n14640 , n15904 );
    and g8786 ( n24685 , n12506 , n9819 );
    xnor g8787 ( n15946 , n4964 , n8259 );
    xnor g8788 ( n579 , n14158 , n11381 );
    xnor g8789 ( n6095 , n25757 , n26201 );
    xnor g8790 ( n17411 , n13692 , n12617 );
    not g8791 ( n24280 , n11221 );
    and g8792 ( n24680 , n6259 , n24152 );
    or g8793 ( n19744 , n10542 , n10014 );
    or g8794 ( n6002 , n1108 , n22075 );
    or g8795 ( n2237 , n12153 , n10148 );
    not g8796 ( n16845 , n20189 );
    nor g8797 ( n9177 , n15932 , n2385 );
    and g8798 ( n16109 , n12394 , n25034 );
    or g8799 ( n18436 , n14551 , n16677 );
    xnor g8800 ( n10961 , n16001 , n1049 );
    xnor g8801 ( n21140 , n26328 , n4746 );
    and g8802 ( n18784 , n25664 , n3008 );
    or g8803 ( n16388 , n997 , n21480 );
    xnor g8804 ( n7765 , n25165 , n20308 );
    xnor g8805 ( n26240 , n14340 , n20302 );
    and g8806 ( n95 , n24738 , n17546 );
    not g8807 ( n18617 , n3118 );
    xnor g8808 ( n2436 , n17764 , n25858 );
    and g8809 ( n4001 , n12791 , n16018 );
    or g8810 ( n24120 , n20170 , n1827 );
    and g8811 ( n4138 , n16777 , n13694 );
    not g8812 ( n17979 , n11566 );
    or g8813 ( n25292 , n3575 , n12936 );
    xnor g8814 ( n24309 , n3568 , n6071 );
    xnor g8815 ( n18903 , n13319 , n15490 );
    not g8816 ( n13108 , n27078 );
    and g8817 ( n18568 , n20606 , n5807 );
    xnor g8818 ( n20590 , n6266 , n447 );
    or g8819 ( n2395 , n8770 , n2286 );
    or g8820 ( n16115 , n12473 , n12681 );
    or g8821 ( n5306 , n12354 , n8581 );
    or g8822 ( n15843 , n23445 , n13733 );
    xnor g8823 ( n8329 , n22793 , n15077 );
    and g8824 ( n26774 , n13391 , n21626 );
    xnor g8825 ( n3722 , n337 , n16507 );
    xnor g8826 ( n23174 , n109 , n592 );
    xnor g8827 ( n15438 , n7234 , n21146 );
    xnor g8828 ( n10913 , n26894 , n16573 );
    not g8829 ( n24305 , n21489 );
    xnor g8830 ( n12191 , n56 , n20506 );
    not g8831 ( n25184 , n9817 );
    xnor g8832 ( n15869 , n17289 , n9858 );
    or g8833 ( n19421 , n14621 , n26581 );
    nor g8834 ( n20158 , n3981 , n23805 );
    or g8835 ( n17245 , n16324 , n10075 );
    xnor g8836 ( n14587 , n9789 , n2764 );
    nor g8837 ( n16057 , n1171 , n3407 );
    or g8838 ( n20758 , n1618 , n9218 );
    or g8839 ( n4329 , n20743 , n25019 );
    and g8840 ( n7328 , n12991 , n24700 );
    and g8841 ( n27206 , n23449 , n5382 );
    or g8842 ( n19573 , n3464 , n4217 );
    or g8843 ( n26812 , n6602 , n24465 );
    and g8844 ( n26791 , n14049 , n11360 );
    and g8845 ( n23135 , n25072 , n16458 );
    nor g8846 ( n13659 , n6580 , n16608 );
    and g8847 ( n26664 , n18493 , n15356 );
    xnor g8848 ( n2483 , n8303 , n1733 );
    and g8849 ( n14103 , n4556 , n254 );
    not g8850 ( n25258 , n15447 );
    xnor g8851 ( n12013 , n2163 , n10346 );
    or g8852 ( n16619 , n24327 , n23185 );
    xnor g8853 ( n2133 , n2281 , n6814 );
    and g8854 ( n10696 , n16009 , n12910 );
    xnor g8855 ( n3544 , n4748 , n11486 );
    and g8856 ( n23729 , n9050 , n11789 );
    xnor g8857 ( n16392 , n636 , n24256 );
    and g8858 ( n17167 , n2190 , n17786 );
    and g8859 ( n25434 , n11011 , n10217 );
    or g8860 ( n5190 , n17254 , n14313 );
    xnor g8861 ( n4564 , n14256 , n25751 );
    xnor g8862 ( n12289 , n26661 , n26808 );
    xnor g8863 ( n25017 , n24143 , n13183 );
    not g8864 ( n25713 , n24281 );
    and g8865 ( n6220 , n6598 , n749 );
    xnor g8866 ( n12352 , n402 , n24815 );
    nor g8867 ( n15034 , n5302 , n3694 );
    or g8868 ( n19824 , n26678 , n12532 );
    xnor g8869 ( n16506 , n717 , n10927 );
    or g8870 ( n15455 , n1735 , n20618 );
    or g8871 ( n13601 , n22031 , n20824 );
    xnor g8872 ( n13658 , n9096 , n25937 );
    not g8873 ( n20074 , n429 );
    xnor g8874 ( n8113 , n6030 , n2350 );
    xnor g8875 ( n24988 , n10955 , n12630 );
    or g8876 ( n19302 , n4099 , n13717 );
    or g8877 ( n12401 , n2689 , n21965 );
    not g8878 ( n20043 , n11377 );
    and g8879 ( n9497 , n20102 , n14269 );
    xnor g8880 ( n16359 , n7694 , n7650 );
    xnor g8881 ( n25115 , n10845 , n21705 );
    or g8882 ( n10706 , n8964 , n18126 );
    xnor g8883 ( n3173 , n22180 , n8855 );
    xnor g8884 ( n13743 , n10074 , n1410 );
    and g8885 ( n7332 , n22893 , n8481 );
    buf g8886 ( n5145 , n618 );
    or g8887 ( n13785 , n24635 , n24162 );
    xnor g8888 ( n3077 , n2666 , n932 );
    xnor g8889 ( n10311 , n24443 , n9422 );
    and g8890 ( n21852 , n1422 , n24246 );
    or g8891 ( n25136 , n24209 , n7671 );
    and g8892 ( n20930 , n1229 , n25410 );
    not g8893 ( n18921 , n1618 );
    not g8894 ( n26450 , n15182 );
    nor g8895 ( n26404 , n5172 , n26124 );
    nor g8896 ( n6221 , n12702 , n12507 );
    xnor g8897 ( n9024 , n20259 , n22043 );
    not g8898 ( n9300 , n25192 );
    nor g8899 ( n10487 , n22695 , n1278 );
    and g8900 ( n25278 , n17422 , n9330 );
    xnor g8901 ( n25518 , n10609 , n466 );
    xnor g8902 ( n26989 , n20077 , n3952 );
    not g8903 ( n14750 , n18734 );
    and g8904 ( n20958 , n14297 , n18911 );
    or g8905 ( n13457 , n9649 , n19613 );
    xnor g8906 ( n14350 , n15921 , n7691 );
    xnor g8907 ( n20891 , n18812 , n1222 );
    xnor g8908 ( n5183 , n16605 , n5804 );
    or g8909 ( n23 , n8222 , n3435 );
    xnor g8910 ( n14511 , n2918 , n8305 );
    not g8911 ( n12735 , n11467 );
    nor g8912 ( n13575 , n8930 , n22772 );
    and g8913 ( n4128 , n17740 , n25951 );
    or g8914 ( n17915 , n3411 , n24824 );
    and g8915 ( n7076 , n22441 , n21776 );
    and g8916 ( n13201 , n9251 , n24851 );
    or g8917 ( n22314 , n24227 , n22561 );
    and g8918 ( n1491 , n13279 , n695 );
    xnor g8919 ( n5874 , n3341 , n16858 );
    and g8920 ( n20867 , n15246 , n26338 );
    not g8921 ( n8064 , n1002 );
    not g8922 ( n25900 , n23688 );
    or g8923 ( n15448 , n6357 , n16752 );
    xnor g8924 ( n22695 , n18630 , n8581 );
    and g8925 ( n24197 , n24084 , n23458 );
    or g8926 ( n21146 , n11897 , n4480 );
    xnor g8927 ( n11276 , n11018 , n1525 );
    nor g8928 ( n10026 , n1380 , n10843 );
    nor g8929 ( n9356 , n25038 , n22626 );
    and g8930 ( n5639 , n20281 , n12193 );
    or g8931 ( n21336 , n7775 , n24734 );
    xnor g8932 ( n19551 , n9411 , n12546 );
    or g8933 ( n532 , n3518 , n935 );
    and g8934 ( n23455 , n16029 , n25674 );
    not g8935 ( n8308 , n26964 );
    nor g8936 ( n6653 , n15127 , n13562 );
    and g8937 ( n7200 , n3702 , n15634 );
    nor g8938 ( n8105 , n27114 , n17727 );
    or g8939 ( n16008 , n10448 , n6471 );
    or g8940 ( n20736 , n17501 , n25991 );
    nor g8941 ( n26864 , n9595 , n27066 );
    and g8942 ( n25854 , n5140 , n6705 );
    and g8943 ( n7115 , n13174 , n14263 );
    and g8944 ( n16059 , n26036 , n1505 );
    or g8945 ( n15381 , n9991 , n24061 );
    nor g8946 ( n20605 , n13489 , n20575 );
    not g8947 ( n821 , n22626 );
    and g8948 ( n14407 , n22844 , n1836 );
    xnor g8949 ( n8615 , n20169 , n4426 );
    and g8950 ( n22293 , n11610 , n9965 );
    or g8951 ( n3627 , n15109 , n10125 );
    or g8952 ( n1899 , n10548 , n9333 );
    xnor g8953 ( n21762 , n19084 , n9598 );
    and g8954 ( n6159 , n26682 , n17964 );
    xnor g8955 ( n17461 , n19926 , n2193 );
    not g8956 ( n18869 , n2657 );
    not g8957 ( n24081 , n5882 );
    or g8958 ( n13358 , n10568 , n8309 );
    or g8959 ( n3762 , n24991 , n4321 );
    xnor g8960 ( n5765 , n9079 , n24632 );
    xnor g8961 ( n2832 , n13231 , n9003 );
    and g8962 ( n18388 , n12954 , n21087 );
    xnor g8963 ( n11401 , n11924 , n3993 );
    or g8964 ( n8631 , n20327 , n9538 );
    not g8965 ( n16084 , n24170 );
    or g8966 ( n12716 , n19109 , n5114 );
    and g8967 ( n11432 , n5547 , n6625 );
    or g8968 ( n12619 , n6750 , n11670 );
    nor g8969 ( n10637 , n12944 , n3448 );
    and g8970 ( n19041 , n20446 , n24606 );
    or g8971 ( n12669 , n12872 , n8318 );
    or g8972 ( n18670 , n18600 , n13723 );
    nor g8973 ( n2725 , n7691 , n15921 );
    not g8974 ( n13843 , n5357 );
    or g8975 ( n11076 , n1706 , n13032 );
    nor g8976 ( n25896 , n23849 , n16274 );
    not g8977 ( n4479 , n692 );
    xnor g8978 ( n10322 , n10920 , n18537 );
    or g8979 ( n21899 , n14641 , n11031 );
    xnor g8980 ( n26929 , n4372 , n5350 );
    or g8981 ( n19689 , n26961 , n1639 );
    xnor g8982 ( n16473 , n17419 , n21134 );
    xnor g8983 ( n21577 , n3992 , n11882 );
    or g8984 ( n21452 , n11232 , n15518 );
    not g8985 ( n2939 , n23990 );
    or g8986 ( n15549 , n21509 , n25608 );
    nor g8987 ( n21410 , n15732 , n16058 );
    xnor g8988 ( n9749 , n7177 , n13393 );
    xnor g8989 ( n554 , n24332 , n13504 );
    xnor g8990 ( n18780 , n1384 , n17715 );
    not g8991 ( n3086 , n3581 );
    or g8992 ( n9606 , n22445 , n18492 );
    xnor g8993 ( n16973 , n19941 , n10577 );
    not g8994 ( n13136 , n23885 );
    xnor g8995 ( n18647 , n18907 , n18901 );
    not g8996 ( n2156 , n7305 );
    xnor g8997 ( n6183 , n23812 , n22099 );
    or g8998 ( n5932 , n3050 , n7684 );
    xnor g8999 ( n26220 , n24809 , n434 );
    nor g9000 ( n12167 , n19888 , n24188 );
    nor g9001 ( n22905 , n20478 , n1204 );
    or g9002 ( n8822 , n19789 , n4978 );
    xnor g9003 ( n26069 , n21493 , n15746 );
    and g9004 ( n19418 , n15687 , n22048 );
    or g9005 ( n25675 , n20191 , n20799 );
    xnor g9006 ( n7575 , n3194 , n7147 );
    and g9007 ( n17124 , n3116 , n24980 );
    xnor g9008 ( n10643 , n1079 , n15411 );
    nor g9009 ( n16760 , n15182 , n20065 );
    xnor g9010 ( n13555 , n527 , n6369 );
    not g9011 ( n20628 , n22226 );
    or g9012 ( n683 , n3225 , n9619 );
    not g9013 ( n8389 , n2878 );
    xnor g9014 ( n4739 , n25797 , n10611 );
    xnor g9015 ( n26896 , n5633 , n13580 );
    xnor g9016 ( n25983 , n16261 , n15158 );
    or g9017 ( n2674 , n4028 , n25870 );
    or g9018 ( n7589 , n3100 , n5551 );
    or g9019 ( n7991 , n22069 , n6943 );
    nor g9020 ( n13337 , n11393 , n2409 );
    nor g9021 ( n17439 , n13023 , n9548 );
    or g9022 ( n4460 , n10949 , n22095 );
    nor g9023 ( n20208 , n2252 , n18495 );
    or g9024 ( n7405 , n17368 , n3019 );
    nor g9025 ( n8467 , n1222 , n22021 );
    or g9026 ( n24637 , n26949 , n4641 );
    not g9027 ( n11550 , n7917 );
    not g9028 ( n11646 , n16446 );
    xnor g9029 ( n3387 , n13463 , n25475 );
    not g9030 ( n3496 , n6847 );
    and g9031 ( n20098 , n6206 , n232 );
    and g9032 ( n558 , n3896 , n5502 );
    not g9033 ( n2155 , n3051 );
    or g9034 ( n12896 , n11776 , n19629 );
    xnor g9035 ( n14499 , n4361 , n25514 );
    nor g9036 ( n1880 , n13863 , n23160 );
    nor g9037 ( n14631 , n1340 , n18742 );
    xnor g9038 ( n11474 , n11944 , n15167 );
    or g9039 ( n14285 , n456 , n8437 );
    xnor g9040 ( n3431 , n3019 , n15241 );
    xnor g9041 ( n8491 , n181 , n15766 );
    or g9042 ( n15523 , n22360 , n24776 );
    not g9043 ( n11582 , n19147 );
    or g9044 ( n3447 , n26747 , n24666 );
    xnor g9045 ( n15515 , n16524 , n987 );
    and g9046 ( n1623 , n13519 , n10226 );
    not g9047 ( n812 , n16562 );
    and g9048 ( n12972 , n6795 , n21439 );
    or g9049 ( n25447 , n8948 , n16474 );
    xnor g9050 ( n14280 , n8933 , n11321 );
    nor g9051 ( n18060 , n11711 , n17308 );
    or g9052 ( n14752 , n14104 , n10079 );
    not g9053 ( n21362 , n11815 );
    not g9054 ( n2618 , n4435 );
    and g9055 ( n13955 , n2870 , n14667 );
    or g9056 ( n8043 , n8840 , n25853 );
    not g9057 ( n216 , n21751 );
    xnor g9058 ( n8488 , n23760 , n14528 );
    or g9059 ( n6886 , n24183 , n12605 );
    nor g9060 ( n14665 , n6494 , n8832 );
    not g9061 ( n2768 , n2161 );
    and g9062 ( n21065 , n9428 , n7851 );
    xnor g9063 ( n3671 , n1232 , n19913 );
    and g9064 ( n26571 , n18409 , n4940 );
    xnor g9065 ( n17204 , n20547 , n26511 );
    and g9066 ( n10736 , n26077 , n16751 );
    or g9067 ( n23916 , n21623 , n20597 );
    or g9068 ( n5717 , n4531 , n21833 );
    or g9069 ( n16585 , n9910 , n7319 );
    xnor g9070 ( n7783 , n19888 , n20734 );
    xnor g9071 ( n6963 , n7614 , n4954 );
    xnor g9072 ( n26332 , n26587 , n25406 );
    or g9073 ( n13682 , n19149 , n13133 );
    nor g9074 ( n22942 , n11559 , n6351 );
    xnor g9075 ( n538 , n9373 , n24510 );
    or g9076 ( n596 , n10469 , n11499 );
    and g9077 ( n4668 , n2671 , n26183 );
    xnor g9078 ( n25608 , n13432 , n23174 );
    or g9079 ( n14759 , n8736 , n5914 );
    and g9080 ( n6954 , n26534 , n21199 );
    or g9081 ( n15091 , n9540 , n12825 );
    or g9082 ( n20568 , n7319 , n23488 );
    or g9083 ( n8470 , n4328 , n25298 );
    not g9084 ( n3239 , n1946 );
    or g9085 ( n20559 , n16893 , n19779 );
    nor g9086 ( n17044 , n17929 , n21923 );
    not g9087 ( n21219 , n15333 );
    or g9088 ( n6434 , n20567 , n6849 );
    xnor g9089 ( n10859 , n16458 , n20907 );
    xnor g9090 ( n26775 , n25750 , n6875 );
    xnor g9091 ( n10350 , n11467 , n26015 );
    xnor g9092 ( n26192 , n11929 , n26744 );
    xnor g9093 ( n1416 , n2705 , n535 );
    nor g9094 ( n7581 , n5706 , n24821 );
    or g9095 ( n17622 , n4217 , n18055 );
    and g9096 ( n12248 , n7410 , n8458 );
    or g9097 ( n14214 , n26971 , n10613 );
    not g9098 ( n279 , n15872 );
    xnor g9099 ( n22380 , n2893 , n7039 );
    or g9100 ( n10759 , n14964 , n12803 );
    nor g9101 ( n8354 , n9632 , n197 );
    and g9102 ( n20280 , n5583 , n26631 );
    xnor g9103 ( n24020 , n6877 , n874 );
    xnor g9104 ( n22416 , n16106 , n15000 );
    or g9105 ( n7556 , n15837 , n14844 );
    or g9106 ( n25295 , n25113 , n9881 );
    or g9107 ( n12862 , n12258 , n8964 );
    or g9108 ( n14934 , n5388 , n19341 );
    nor g9109 ( n17448 , n26295 , n16896 );
    nor g9110 ( n15866 , n7059 , n6202 );
    or g9111 ( n8291 , n5071 , n3200 );
    xnor g9112 ( n16072 , n21232 , n22744 );
    xnor g9113 ( n10775 , n24591 , n20767 );
    xnor g9114 ( n26225 , n15894 , n18899 );
    and g9115 ( n20307 , n20396 , n11332 );
    or g9116 ( n7303 , n1437 , n12488 );
    not g9117 ( n13760 , n16626 );
    nor g9118 ( n20965 , n20153 , n2964 );
    or g9119 ( n19820 , n19298 , n1173 );
    not g9120 ( n18115 , n7524 );
    and g9121 ( n19928 , n14143 , n18605 );
    not g9122 ( n7394 , n26831 );
    and g9123 ( n18197 , n18245 , n22965 );
    or g9124 ( n15551 , n11963 , n6203 );
    or g9125 ( n18885 , n1289 , n7813 );
    and g9126 ( n26453 , n15668 , n13482 );
    not g9127 ( n3719 , n1792 );
    and g9128 ( n4609 , n1137 , n12290 );
    and g9129 ( n14453 , n21334 , n15273 );
    xnor g9130 ( n3179 , n1878 , n9335 );
    or g9131 ( n5667 , n5004 , n27171 );
    xnor g9132 ( n6707 , n383 , n16940 );
    or g9133 ( n25557 , n6929 , n22008 );
    not g9134 ( n11317 , n16360 );
    not g9135 ( n11627 , n25317 );
    not g9136 ( n11442 , n15024 );
    nor g9137 ( n5109 , n22404 , n7324 );
    nor g9138 ( n18600 , n25426 , n1532 );
    or g9139 ( n12717 , n5268 , n16095 );
    or g9140 ( n22927 , n6617 , n18941 );
    nor g9141 ( n11364 , n24237 , n19592 );
    and g9142 ( n14043 , n6987 , n18501 );
    xnor g9143 ( n6798 , n14661 , n25322 );
    not g9144 ( n2903 , n3582 );
    or g9145 ( n21211 , n971 , n1926 );
    and g9146 ( n23772 , n12567 , n12279 );
    or g9147 ( n2991 , n22905 , n26587 );
    nor g9148 ( n489 , n5958 , n22349 );
    not g9149 ( n22003 , n18496 );
    and g9150 ( n24843 , n14802 , n5281 );
    not g9151 ( n14677 , n4886 );
    not g9152 ( n19328 , n21860 );
    or g9153 ( n24055 , n1039 , n11110 );
    xnor g9154 ( n7102 , n25167 , n1104 );
    xnor g9155 ( n24706 , n3837 , n24374 );
    or g9156 ( n2258 , n18594 , n20907 );
    xnor g9157 ( n12016 , n22783 , n18578 );
    not g9158 ( n22736 , n9881 );
    xnor g9159 ( n17704 , n3203 , n2935 );
    xnor g9160 ( n3730 , n22229 , n7583 );
    xnor g9161 ( n14845 , n9163 , n11508 );
    xnor g9162 ( n26359 , n10509 , n9244 );
    or g9163 ( n6378 , n26496 , n25800 );
    or g9164 ( n14137 , n3239 , n14649 );
    not g9165 ( n4874 , n17575 );
    or g9166 ( n15388 , n9549 , n7489 );
    nor g9167 ( n25161 , n25381 , n14573 );
    nor g9168 ( n9048 , n22170 , n16848 );
    and g9169 ( n15491 , n23746 , n7269 );
    and g9170 ( n20676 , n5255 , n6446 );
    or g9171 ( n12135 , n22595 , n15421 );
    xnor g9172 ( n20080 , n6823 , n2491 );
    or g9173 ( n17807 , n22887 , n4700 );
    and g9174 ( n26230 , n5055 , n1318 );
    or g9175 ( n18038 , n12400 , n2966 );
    not g9176 ( n7399 , n19568 );
    not g9177 ( n16106 , n18137 );
    or g9178 ( n13397 , n6042 , n5051 );
    nor g9179 ( n19640 , n10683 , n21134 );
    and g9180 ( n14335 , n17260 , n5457 );
    nor g9181 ( n862 , n852 , n11848 );
    nor g9182 ( n23609 , n22379 , n9967 );
    not g9183 ( n18557 , n18263 );
    xnor g9184 ( n3193 , n16793 , n7692 );
    or g9185 ( n24513 , n22558 , n16548 );
    or g9186 ( n22369 , n2498 , n947 );
    or g9187 ( n8752 , n1669 , n16639 );
    and g9188 ( n9360 , n4234 , n18650 );
    and g9189 ( n20665 , n5005 , n2654 );
    nor g9190 ( n26990 , n2230 , n13842 );
    nor g9191 ( n19967 , n6352 , n13435 );
    xnor g9192 ( n5827 , n16822 , n14580 );
    xnor g9193 ( n17163 , n4874 , n11708 );
    or g9194 ( n5647 , n15861 , n4887 );
    not g9195 ( n2460 , n11106 );
    xnor g9196 ( n26698 , n8956 , n8089 );
    and g9197 ( n19990 , n17714 , n453 );
    and g9198 ( n25382 , n6750 , n11670 );
    xnor g9199 ( n10242 , n14688 , n9084 );
    nor g9200 ( n22054 , n11989 , n14087 );
    nor g9201 ( n2928 , n22363 , n27065 );
    and g9202 ( n20240 , n4527 , n5797 );
    not g9203 ( n10911 , n7727 );
    xnor g9204 ( n26656 , n15385 , n24568 );
    or g9205 ( n26106 , n5842 , n3590 );
    and g9206 ( n1737 , n16958 , n18270 );
    and g9207 ( n23446 , n9884 , n20093 );
    xnor g9208 ( n4340 , n20440 , n21731 );
    nor g9209 ( n9416 , n7949 , n16609 );
    xnor g9210 ( n1261 , n27042 , n25415 );
    nor g9211 ( n25199 , n18434 , n20051 );
    and g9212 ( n3225 , n21915 , n2509 );
    or g9213 ( n14259 , n782 , n27042 );
    or g9214 ( n26862 , n21829 , n22465 );
    xnor g9215 ( n16701 , n17824 , n5860 );
    xnor g9216 ( n17466 , n17797 , n27021 );
    not g9217 ( n15891 , n12297 );
    xnor g9218 ( n25908 , n5852 , n16963 );
    and g9219 ( n24312 , n1749 , n15514 );
    not g9220 ( n16470 , n23366 );
    not g9221 ( n13590 , n25119 );
    and g9222 ( n21659 , n1682 , n3318 );
    and g9223 ( n8387 , n12634 , n16920 );
    xnor g9224 ( n22481 , n8456 , n26744 );
    xnor g9225 ( n3016 , n13114 , n16641 );
    xnor g9226 ( n26566 , n24560 , n27139 );
    xnor g9227 ( n20002 , n9747 , n17089 );
    or g9228 ( n8923 , n17630 , n18557 );
    or g9229 ( n22788 , n2799 , n2271 );
    xnor g9230 ( n6703 , n19120 , n5129 );
    xnor g9231 ( n19714 , n2281 , n18755 );
    xnor g9232 ( n2895 , n1345 , n9106 );
    nor g9233 ( n12250 , n17380 , n10962 );
    and g9234 ( n14487 , n26032 , n23171 );
    nor g9235 ( n9920 , n8100 , n2481 );
    or g9236 ( n22362 , n18971 , n1446 );
    xnor g9237 ( n17693 , n15456 , n25365 );
    xnor g9238 ( n14506 , n23285 , n25704 );
    nor g9239 ( n23940 , n20043 , n23264 );
    xnor g9240 ( n19785 , n3802 , n8778 );
    and g9241 ( n9885 , n20625 , n21453 );
    or g9242 ( n24581 , n19668 , n21223 );
    xnor g9243 ( n15992 , n2139 , n3710 );
    xnor g9244 ( n672 , n17411 , n22727 );
    and g9245 ( n21080 , n16154 , n6101 );
    or g9246 ( n8621 , n9310 , n4119 );
    and g9247 ( n9333 , n19991 , n16651 );
    nor g9248 ( n1888 , n11186 , n12821 );
    xnor g9249 ( n14009 , n10053 , n15539 );
    xnor g9250 ( n4176 , n19498 , n8246 );
    not g9251 ( n10296 , n5091 );
    and g9252 ( n26462 , n11113 , n24272 );
    or g9253 ( n9055 , n18714 , n729 );
    not g9254 ( n25291 , n9873 );
    or g9255 ( n11768 , n4986 , n21840 );
    xnor g9256 ( n26888 , n15796 , n8528 );
    xnor g9257 ( n10592 , n2897 , n22358 );
    and g9258 ( n1298 , n21551 , n27013 );
    nor g9259 ( n12596 , n20042 , n24466 );
    xnor g9260 ( n7959 , n22702 , n14074 );
    not g9261 ( n9099 , n1040 );
    not g9262 ( n20488 , n20489 );
    xnor g9263 ( n18977 , n5923 , n17481 );
    or g9264 ( n25836 , n27172 , n20075 );
    not g9265 ( n16843 , n161 );
    and g9266 ( n1607 , n26125 , n26321 );
    nor g9267 ( n16901 , n3740 , n21784 );
    not g9268 ( n12373 , n17274 );
    and g9269 ( n6769 , n5183 , n4448 );
    nor g9270 ( n6597 , n20630 , n25312 );
    xnor g9271 ( n24816 , n16609 , n12906 );
    not g9272 ( n2790 , n21981 );
    and g9273 ( n24182 , n12757 , n3507 );
    and g9274 ( n907 , n573 , n19345 );
    or g9275 ( n10270 , n11399 , n15483 );
    or g9276 ( n9436 , n18506 , n5226 );
    xnor g9277 ( n9218 , n9876 , n3330 );
    or g9278 ( n1746 , n26133 , n16570 );
    xnor g9279 ( n12569 , n5600 , n8022 );
    or g9280 ( n7463 , n16366 , n18203 );
    xnor g9281 ( n15814 , n24392 , n21779 );
    nor g9282 ( n1310 , n15722 , n1184 );
    not g9283 ( n17323 , n18950 );
    xnor g9284 ( n23862 , n2803 , n9645 );
    or g9285 ( n24588 , n18754 , n24499 );
    xnor g9286 ( n26795 , n10418 , n3593 );
    or g9287 ( n9906 , n4934 , n14061 );
    or g9288 ( n17950 , n24267 , n5897 );
    and g9289 ( n2181 , n17665 , n1496 );
    not g9290 ( n20327 , n20770 );
    or g9291 ( n26320 , n631 , n12734 );
    xnor g9292 ( n24112 , n9100 , n26264 );
    nor g9293 ( n13377 , n16707 , n20120 );
    not g9294 ( n11806 , n5408 );
    and g9295 ( n25109 , n15396 , n25578 );
    xnor g9296 ( n11301 , n21839 , n16544 );
    nor g9297 ( n621 , n23235 , n8253 );
    or g9298 ( n1436 , n15740 , n2243 );
    not g9299 ( n10156 , n7657 );
    or g9300 ( n22097 , n19608 , n2730 );
    xnor g9301 ( n2860 , n1393 , n8936 );
    and g9302 ( n18542 , n12554 , n20711 );
    xnor g9303 ( n25748 , n22609 , n22829 );
    or g9304 ( n4949 , n26762 , n21555 );
    and g9305 ( n26140 , n8117 , n3280 );
    xnor g9306 ( n3076 , n13502 , n27069 );
    and g9307 ( n17520 , n4386 , n10583 );
    xnor g9308 ( n13825 , n12658 , n8232 );
    or g9309 ( n26922 , n4915 , n5052 );
    and g9310 ( n11864 , n4627 , n13334 );
    xnor g9311 ( n1648 , n1970 , n22043 );
    and g9312 ( n8444 , n13087 , n13433 );
    nor g9313 ( n14781 , n26363 , n21596 );
    xnor g9314 ( n8724 , n15657 , n14124 );
    not g9315 ( n26688 , n25751 );
    not g9316 ( n5304 , n8001 );
    xnor g9317 ( n3117 , n8745 , n24278 );
    not g9318 ( n4132 , n9655 );
    nor g9319 ( n17354 , n11751 , n3245 );
    and g9320 ( n23809 , n16476 , n15008 );
    not g9321 ( n17706 , n19508 );
    and g9322 ( n24487 , n8704 , n18665 );
    or g9323 ( n26416 , n22703 , n10299 );
    or g9324 ( n8654 , n1819 , n15521 );
    not g9325 ( n13696 , n19804 );
    not g9326 ( n18735 , n26239 );
    or g9327 ( n18968 , n18823 , n20147 );
    xnor g9328 ( n20786 , n17141 , n3299 );
    xnor g9329 ( n24784 , n26664 , n17538 );
    or g9330 ( n12283 , n12316 , n19168 );
    nor g9331 ( n4218 , n21632 , n26510 );
    nor g9332 ( n2722 , n461 , n22387 );
    or g9333 ( n8061 , n8643 , n26769 );
    or g9334 ( n22950 , n6215 , n4636 );
    and g9335 ( n15848 , n22676 , n11588 );
    xnor g9336 ( n11252 , n25221 , n22507 );
    xnor g9337 ( n18265 , n11454 , n8458 );
    nor g9338 ( n14374 , n19941 , n10577 );
    and g9339 ( n21223 , n25388 , n16288 );
    xnor g9340 ( n22583 , n6034 , n21934 );
    and g9341 ( n24740 , n21653 , n21617 );
    or g9342 ( n12035 , n446 , n11045 );
    or g9343 ( n17797 , n9738 , n6048 );
    or g9344 ( n9034 , n15433 , n24875 );
    xnor g9345 ( n6444 , n8783 , n7979 );
    xnor g9346 ( n18071 , n20910 , n6155 );
    and g9347 ( n21962 , n5960 , n17830 );
    xnor g9348 ( n2804 , n25339 , n12700 );
    or g9349 ( n26491 , n9365 , n9095 );
    not g9350 ( n1594 , n13503 );
    not g9351 ( n19076 , n1690 );
    xnor g9352 ( n9847 , n2113 , n14345 );
    nor g9353 ( n8098 , n19219 , n25251 );
    not g9354 ( n23126 , n26512 );
    or g9355 ( n21571 , n20812 , n3135 );
    and g9356 ( n18267 , n9400 , n11154 );
    nor g9357 ( n19970 , n5103 , n21565 );
    xnor g9358 ( n16543 , n15561 , n19708 );
    or g9359 ( n5369 , n13713 , n20001 );
    nor g9360 ( n12132 , n10146 , n11152 );
    or g9361 ( n25824 , n1725 , n39 );
    xnor g9362 ( n15120 , n2111 , n16473 );
    and g9363 ( n8502 , n20531 , n7645 );
    or g9364 ( n11570 , n4277 , n13685 );
    or g9365 ( n3504 , n1654 , n2425 );
    and g9366 ( n8709 , n4722 , n14323 );
    or g9367 ( n15493 , n13912 , n11980 );
    xnor g9368 ( n3803 , n685 , n25586 );
    nor g9369 ( n11191 , n11209 , n5495 );
    or g9370 ( n13111 , n13751 , n3128 );
    or g9371 ( n22949 , n17293 , n12298 );
    or g9372 ( n18671 , n18003 , n26058 );
    and g9373 ( n3165 , n26361 , n18470 );
    or g9374 ( n6994 , n727 , n15637 );
    nor g9375 ( n10044 , n13494 , n23983 );
    and g9376 ( n19351 , n26797 , n16221 );
    xnor g9377 ( n25446 , n9817 , n13189 );
    not g9378 ( n3547 , n26522 );
    nor g9379 ( n5950 , n2336 , n19366 );
    xnor g9380 ( n8249 , n23657 , n23035 );
    xnor g9381 ( n17367 , n19971 , n6685 );
    or g9382 ( n8927 , n8858 , n23602 );
    and g9383 ( n14057 , n6868 , n5087 );
    and g9384 ( n16235 , n884 , n4617 );
    or g9385 ( n18551 , n240 , n3113 );
    not g9386 ( n15696 , n17056 );
    or g9387 ( n15993 , n26828 , n16070 );
    or g9388 ( n10566 , n20362 , n3548 );
    xnor g9389 ( n9364 , n13121 , n5049 );
    xnor g9390 ( n14271 , n16945 , n15758 );
    or g9391 ( n25580 , n25025 , n8356 );
    or g9392 ( n14724 , n4040 , n18006 );
    or g9393 ( n5583 , n22723 , n7006 );
    xnor g9394 ( n3379 , n23249 , n5077 );
    or g9395 ( n18870 , n16294 , n2944 );
    xnor g9396 ( n23594 , n23983 , n13494 );
    or g9397 ( n15402 , n25452 , n507 );
    xnor g9398 ( n20521 , n22517 , n9226 );
    nor g9399 ( n23239 , n6595 , n6199 );
    xnor g9400 ( n19360 , n17283 , n9429 );
    not g9401 ( n14378 , n1596 );
    xnor g9402 ( n2499 , n19856 , n21687 );
    or g9403 ( n21468 , n9670 , n2873 );
    and g9404 ( n25560 , n20064 , n215 );
    xnor g9405 ( n19589 , n24781 , n21426 );
    and g9406 ( n20467 , n25095 , n7078 );
    xnor g9407 ( n16071 , n19361 , n15918 );
    not g9408 ( n26650 , n20863 );
    and g9409 ( n16300 , n1748 , n11353 );
    xnor g9410 ( n25653 , n5159 , n16734 );
    xnor g9411 ( n10599 , n10500 , n12493 );
    and g9412 ( n23322 , n7237 , n4873 );
    or g9413 ( n2108 , n12546 , n14614 );
    not g9414 ( n16037 , n21080 );
    xnor g9415 ( n15286 , n17184 , n24487 );
    or g9416 ( n25943 , n25441 , n21620 );
    nor g9417 ( n23478 , n18227 , n17397 );
    or g9418 ( n14250 , n5818 , n7365 );
    xnor g9419 ( n9069 , n4093 , n752 );
    and g9420 ( n3992 , n4962 , n23214 );
    xnor g9421 ( n19682 , n23706 , n5984 );
    not g9422 ( n23705 , n25331 );
    xnor g9423 ( n21967 , n23708 , n26808 );
    nor g9424 ( n3831 , n25194 , n6935 );
    or g9425 ( n13986 , n14140 , n20009 );
    xnor g9426 ( n20966 , n19016 , n12039 );
    and g9427 ( n9169 , n16780 , n8188 );
    or g9428 ( n17041 , n15415 , n12119 );
    xnor g9429 ( n17842 , n22716 , n23912 );
    and g9430 ( n20644 , n16508 , n6976 );
    or g9431 ( n16289 , n20681 , n15754 );
    xnor g9432 ( n23371 , n13733 , n16072 );
    nor g9433 ( n2916 , n6356 , n8418 );
    and g9434 ( n25065 , n8766 , n10690 );
    and g9435 ( n25255 , n23281 , n20557 );
    not g9436 ( n15185 , n2382 );
    and g9437 ( n3913 , n5543 , n22409 );
    and g9438 ( n15840 , n5123 , n15482 );
    or g9439 ( n1022 , n19477 , n2114 );
    xnor g9440 ( n2093 , n22417 , n3595 );
    and g9441 ( n8616 , n23001 , n5293 );
    or g9442 ( n26653 , n17092 , n10543 );
    and g9443 ( n6968 , n17509 , n9307 );
    or g9444 ( n574 , n12508 , n25942 );
    nor g9445 ( n19704 , n20296 , n20862 );
    nor g9446 ( n6565 , n5211 , n15910 );
    not g9447 ( n18055 , n22683 );
    xnor g9448 ( n9888 , n8263 , n2904 );
    xnor g9449 ( n10245 , n3149 , n5400 );
    not g9450 ( n24945 , n25186 );
    and g9451 ( n4002 , n3024 , n4949 );
    nor g9452 ( n17185 , n24890 , n10411 );
    not g9453 ( n15417 , n21833 );
    or g9454 ( n13427 , n13028 , n11579 );
    or g9455 ( n3177 , n15685 , n5477 );
    xnor g9456 ( n21438 , n4213 , n19454 );
    xnor g9457 ( n19191 , n27144 , n23980 );
    and g9458 ( n7321 , n23841 , n556 );
    xor g9459 ( n27192 , n18758 , n20259 );
    and g9460 ( n15457 , n2825 , n15948 );
    and g9461 ( n13226 , n5533 , n12080 );
    not g9462 ( n15138 , n25523 );
    nor g9463 ( n21563 , n7991 , n3133 );
    xnor g9464 ( n24900 , n4492 , n23002 );
    and g9465 ( n3381 , n14595 , n18367 );
    or g9466 ( n26049 , n8932 , n7795 );
    xnor g9467 ( n8422 , n1737 , n15607 );
    buf g9468 ( n12522 , n18137 );
    not g9469 ( n3380 , n13884 );
    xor g9470 ( n2489 , n26491 , n7894 );
    xnor g9471 ( n12236 , n10844 , n8615 );
    not g9472 ( n2036 , n3014 );
    nor g9473 ( n17944 , n19303 , n15313 );
    or g9474 ( n9710 , n16033 , n15852 );
    and g9475 ( n22505 , n11153 , n14639 );
    not g9476 ( n7517 , n2013 );
    or g9477 ( n6922 , n3904 , n1653 );
    xnor g9478 ( n6541 , n23197 , n11276 );
    xnor g9479 ( n22832 , n11459 , n1837 );
    or g9480 ( n13721 , n450 , n16028 );
    xnor g9481 ( n18405 , n5545 , n4953 );
    or g9482 ( n18167 , n12245 , n19666 );
    not g9483 ( n24617 , n3002 );
    or g9484 ( n14258 , n3320 , n7879 );
    or g9485 ( n5681 , n1751 , n12008 );
    not g9486 ( n25327 , n21216 );
    or g9487 ( n15980 , n8858 , n5886 );
    and g9488 ( n14264 , n1745 , n4135 );
    and g9489 ( n13361 , n1587 , n1685 );
    xnor g9490 ( n6012 , n26242 , n24147 );
    and g9491 ( n7599 , n18062 , n8478 );
    xnor g9492 ( n25427 , n22972 , n8003 );
    xnor g9493 ( n4201 , n14582 , n8946 );
    xnor g9494 ( n11496 , n26967 , n12203 );
    xnor g9495 ( n23803 , n23999 , n13190 );
    or g9496 ( n4391 , n8996 , n9955 );
    xnor g9497 ( n4682 , n5555 , n21649 );
    and g9498 ( n26249 , n5778 , n4965 );
    nor g9499 ( n8787 , n8931 , n1003 );
    xnor g9500 ( n5660 , n7536 , n19200 );
    and g9501 ( n19936 , n8727 , n21075 );
    and g9502 ( n24980 , n26064 , n9095 );
    xnor g9503 ( n9204 , n26490 , n11168 );
    not g9504 ( n23631 , n12375 );
    xnor g9505 ( n24654 , n1347 , n7962 );
    nor g9506 ( n16625 , n12971 , n17953 );
    xnor g9507 ( n10055 , n13330 , n12256 );
    or g9508 ( n17231 , n26514 , n23176 );
    and g9509 ( n20688 , n6770 , n1175 );
    or g9510 ( n14833 , n3416 , n3167 );
    or g9511 ( n9028 , n10125 , n8522 );
    xnor g9512 ( n2660 , n331 , n24616 );
    and g9513 ( n4608 , n4296 , n11019 );
    or g9514 ( n10640 , n842 , n1543 );
    xnor g9515 ( n2690 , n12541 , n26901 );
    nor g9516 ( n3249 , n7455 , n17255 );
    xnor g9517 ( n21800 , n3580 , n24724 );
    or g9518 ( n18828 , n642 , n4127 );
    and g9519 ( n20491 , n5304 , n15437 );
    nor g9520 ( n1207 , n21627 , n5415 );
    nor g9521 ( n12945 , n3009 , n6011 );
    or g9522 ( n14594 , n5518 , n3194 );
    nor g9523 ( n6622 , n11953 , n13896 );
    and g9524 ( n14579 , n23813 , n3912 );
    not g9525 ( n18054 , n4576 );
    and g9526 ( n7197 , n5657 , n14395 );
    xnor g9527 ( n16984 , n24774 , n3460 );
    xnor g9528 ( n128 , n13329 , n15884 );
    nor g9529 ( n1597 , n4957 , n7421 );
    nor g9530 ( n22177 , n12686 , n5642 );
    and g9531 ( n19726 , n17184 , n24487 );
    xnor g9532 ( n4989 , n27142 , n9312 );
    and g9533 ( n20052 , n2594 , n21991 );
    or g9534 ( n1561 , n8597 , n8194 );
    or g9535 ( n13002 , n14942 , n3497 );
    xnor g9536 ( n21101 , n20711 , n16396 );
    xnor g9537 ( n4366 , n17213 , n11302 );
    and g9538 ( n14186 , n1458 , n21372 );
    xnor g9539 ( n299 , n19357 , n21649 );
    not g9540 ( n14204 , n6232 );
    xnor g9541 ( n16339 , n8471 , n21402 );
    not g9542 ( n3006 , n7044 );
    or g9543 ( n17766 , n15453 , n26012 );
    nor g9544 ( n23797 , n9222 , n25054 );
    or g9545 ( n25578 , n1797 , n1837 );
    and g9546 ( n26291 , n24825 , n8009 );
    and g9547 ( n4090 , n12056 , n9892 );
    not g9548 ( n16349 , n14790 );
    or g9549 ( n12523 , n2202 , n19072 );
    not g9550 ( n20206 , n5140 );
    not g9551 ( n10741 , n10482 );
    xnor g9552 ( n22895 , n10440 , n385 );
    xnor g9553 ( n9238 , n16507 , n23250 );
    or g9554 ( n20337 , n22054 , n5473 );
    not g9555 ( n18624 , n25278 );
    xnor g9556 ( n24956 , n13104 , n26420 );
    and g9557 ( n16686 , n18835 , n26416 );
    xnor g9558 ( n12469 , n12781 , n9989 );
    xnor g9559 ( n25462 , n24004 , n12900 );
    nor g9560 ( n12067 , n10470 , n4062 );
    or g9561 ( n9381 , n18730 , n17753 );
    nor g9562 ( n16528 , n11143 , n10709 );
    or g9563 ( n14571 , n25624 , n9653 );
    or g9564 ( n22268 , n10024 , n26141 );
    and g9565 ( n13311 , n23835 , n10947 );
    xnor g9566 ( n25360 , n23881 , n5615 );
    or g9567 ( n20236 , n11785 , n19713 );
    and g9568 ( n19147 , n9927 , n19635 );
    xnor g9569 ( n18993 , n2498 , n26013 );
    nor g9570 ( n22741 , n11578 , n2261 );
    xnor g9571 ( n21239 , n15539 , n24278 );
    xnor g9572 ( n9504 , n20039 , n8694 );
    or g9573 ( n9528 , n6508 , n21710 );
    xnor g9574 ( n26150 , n13846 , n17090 );
    not g9575 ( n4995 , n23185 );
    not g9576 ( n22207 , n18953 );
    not g9577 ( n7470 , n13567 );
    nor g9578 ( n3099 , n13899 , n15242 );
    nor g9579 ( n16800 , n11273 , n23086 );
    or g9580 ( n20545 , n1264 , n26635 );
    or g9581 ( n3267 , n4803 , n20408 );
    or g9582 ( n20097 , n19894 , n22517 );
    nor g9583 ( n12500 , n9373 , n7677 );
    xnor g9584 ( n22654 , n16518 , n23649 );
    not g9585 ( n20150 , n5929 );
    nor g9586 ( n27001 , n9274 , n9814 );
    not g9587 ( n15795 , n7656 );
    not g9588 ( n251 , n26915 );
    not g9589 ( n402 , n22375 );
    and g9590 ( n4857 , n15427 , n10168 );
    or g9591 ( n20024 , n12976 , n18007 );
    and g9592 ( n2362 , n9343 , n15656 );
    not g9593 ( n20365 , n12950 );
    not g9594 ( n10791 , n13119 );
    nor g9595 ( n13365 , n20089 , n21216 );
    or g9596 ( n7796 , n23757 , n8195 );
    or g9597 ( n155 , n3791 , n26876 );
    or g9598 ( n7275 , n4380 , n2998 );
    nor g9599 ( n26788 , n22619 , n22043 );
    not g9600 ( n5745 , n12152 );
    or g9601 ( n26614 , n17996 , n4597 );
    or g9602 ( n12510 , n15756 , n6484 );
    or g9603 ( n2256 , n131 , n23542 );
    or g9604 ( n11342 , n2780 , n2000 );
    nor g9605 ( n15050 , n4603 , n26536 );
    or g9606 ( n4488 , n3185 , n21996 );
    xnor g9607 ( n454 , n1136 , n11667 );
    or g9608 ( n15882 , n14739 , n15458 );
    nor g9609 ( n18057 , n20376 , n6202 );
    nor g9610 ( n24014 , n12699 , n8688 );
    not g9611 ( n10500 , n25685 );
    xnor g9612 ( n18831 , n1216 , n18680 );
    or g9613 ( n21660 , n6140 , n22352 );
    or g9614 ( n15431 , n22336 , n15724 );
    xnor g9615 ( n2149 , n24517 , n26327 );
    and g9616 ( n19628 , n14519 , n14208 );
    or g9617 ( n20657 , n18912 , n18198 );
    xnor g9618 ( n24284 , n26580 , n18768 );
    or g9619 ( n2751 , n20178 , n20508 );
    xnor g9620 ( n24161 , n5897 , n12886 );
    xnor g9621 ( n2280 , n25471 , n23842 );
    or g9622 ( n23618 , n14502 , n18230 );
    or g9623 ( n23909 , n21580 , n16229 );
    xnor g9624 ( n17180 , n210 , n15873 );
    or g9625 ( n20157 , n17793 , n20114 );
    xnor g9626 ( n16833 , n22392 , n8920 );
    xnor g9627 ( n12910 , n1381 , n19070 );
    or g9628 ( n22805 , n3318 , n1682 );
    or g9629 ( n27126 , n14017 , n19750 );
    and g9630 ( n26821 , n9155 , n19490 );
    xnor g9631 ( n9247 , n17275 , n13014 );
    and g9632 ( n493 , n18046 , n1025 );
    or g9633 ( n19049 , n21141 , n26165 );
    nor g9634 ( n920 , n4360 , n17368 );
    and g9635 ( n971 , n21623 , n6503 );
    not g9636 ( n11229 , n14078 );
    or g9637 ( n5628 , n15398 , n21752 );
    xnor g9638 ( n9508 , n15868 , n7988 );
    or g9639 ( n3896 , n24623 , n26638 );
    not g9640 ( n24883 , n15254 );
    not g9641 ( n20196 , n14394 );
    and g9642 ( n11555 , n6588 , n2988 );
    and g9643 ( n17840 , n16992 , n451 );
    or g9644 ( n9516 , n8700 , n24884 );
    not g9645 ( n11988 , n3323 );
    nor g9646 ( n10623 , n2342 , n20245 );
    not g9647 ( n6760 , n14510 );
    nor g9648 ( n759 , n11901 , n10201 );
    or g9649 ( n19931 , n15200 , n8783 );
    and g9650 ( n16480 , n15284 , n26819 );
    nor g9651 ( n13888 , n14288 , n20039 );
    or g9652 ( n23762 , n11898 , n25063 );
    nor g9653 ( n17615 , n1281 , n13169 );
    or g9654 ( n12581 , n22540 , n21041 );
    and g9655 ( n12491 , n19918 , n7404 );
    or g9656 ( n15031 , n359 , n22710 );
    or g9657 ( n24912 , n16540 , n9288 );
    not g9658 ( n26691 , n24786 );
    not g9659 ( n8024 , n19649 );
    or g9660 ( n9127 , n25144 , n5972 );
    and g9661 ( n8360 , n21678 , n684 );
    xnor g9662 ( n20731 , n12308 , n9145 );
    xnor g9663 ( n20523 , n13567 , n1730 );
    and g9664 ( n2610 , n19657 , n17772 );
    and g9665 ( n13167 , n13378 , n10444 );
    or g9666 ( n4161 , n8078 , n15143 );
    or g9667 ( n22567 , n8344 , n13913 );
    or g9668 ( n1213 , n6721 , n7857 );
    xnor g9669 ( n16219 , n10914 , n1481 );
    not g9670 ( n24660 , n18585 );
    or g9671 ( n26002 , n15168 , n26720 );
    xnor g9672 ( n7979 , n26660 , n25643 );
    and g9673 ( n24846 , n19864 , n12581 );
    nor g9674 ( n2520 , n15884 , n2412 );
    or g9675 ( n2449 , n8382 , n7644 );
    nor g9676 ( n13188 , n26691 , n8661 );
    and g9677 ( n207 , n13460 , n10008 );
    or g9678 ( n2504 , n21118 , n2331 );
    xnor g9679 ( n11078 , n7219 , n21834 );
    not g9680 ( n17744 , n20724 );
    not g9681 ( n10568 , n10411 );
    or g9682 ( n22014 , n18737 , n6109 );
    or g9683 ( n10472 , n13708 , n23085 );
    or g9684 ( n16170 , n5922 , n6624 );
    or g9685 ( n9299 , n14 , n16897 );
    or g9686 ( n25747 , n6164 , n25942 );
    xnor g9687 ( n15001 , n11220 , n2944 );
    or g9688 ( n7246 , n25896 , n21184 );
    nor g9689 ( n15272 , n10586 , n15253 );
    and g9690 ( n18731 , n5753 , n5632 );
    not g9691 ( n24351 , n12917 );
    xnor g9692 ( n9313 , n7565 , n22390 );
    xnor g9693 ( n9222 , n24046 , n10929 );
    nor g9694 ( n10987 , n5785 , n16353 );
    nor g9695 ( n5230 , n2057 , n21930 );
    xnor g9696 ( n26903 , n25872 , n19618 );
    not g9697 ( n8695 , n23727 );
    and g9698 ( n2503 , n3069 , n11654 );
    or g9699 ( n26984 , n11384 , n16812 );
    xnor g9700 ( n5046 , n14591 , n14986 );
    or g9701 ( n27196 , n13873 , n24355 );
    xnor g9702 ( n12039 , n17351 , n16507 );
    xnor g9703 ( n26159 , n10921 , n21357 );
    xnor g9704 ( n24283 , n16709 , n12272 );
    or g9705 ( n17486 , n7935 , n11552 );
    and g9706 ( n23973 , n10430 , n18575 );
    and g9707 ( n10940 , n25157 , n26281 );
    xnor g9708 ( n14518 , n1944 , n897 );
    and g9709 ( n11633 , n10311 , n14713 );
    and g9710 ( n7397 , n24588 , n5102 );
    or g9711 ( n7300 , n1757 , n11970 );
    not g9712 ( n23920 , n677 );
    not g9713 ( n24495 , n14448 );
    not g9714 ( n18983 , n26304 );
    and g9715 ( n26728 , n26956 , n7021 );
    not g9716 ( n13109 , n21900 );
    or g9717 ( n4841 , n11756 , n21175 );
    not g9718 ( n19392 , n638 );
    xnor g9719 ( n24724 , n13539 , n20532 );
    xnor g9720 ( n1621 , n1704 , n3356 );
    xnor g9721 ( n12941 , n17327 , n10360 );
    or g9722 ( n16044 , n14655 , n79 );
    xnor g9723 ( n22514 , n8869 , n8381 );
    not g9724 ( n21632 , n1112 );
    and g9725 ( n10578 , n27139 , n24560 );
    not g9726 ( n20299 , n8864 );
    and g9727 ( n16791 , n3937 , n1243 );
    and g9728 ( n24189 , n4147 , n20862 );
    and g9729 ( n19281 , n4431 , n11925 );
    xnor g9730 ( n5731 , n166 , n4376 );
    not g9731 ( n15650 , n5125 );
    and g9732 ( n21432 , n2731 , n16210 );
    not g9733 ( n10689 , n14453 );
    or g9734 ( n21775 , n9053 , n23488 );
    xnor g9735 ( n25606 , n8106 , n13262 );
    and g9736 ( n6600 , n22298 , n19751 );
    xnor g9737 ( n13793 , n21412 , n9821 );
    and g9738 ( n3470 , n26997 , n19059 );
    and g9739 ( n8303 , n12597 , n19099 );
    and g9740 ( n11684 , n26275 , n16434 );
    or g9741 ( n22580 , n7741 , n3123 );
    xnor g9742 ( n25192 , n12032 , n2083 );
    xnor g9743 ( n1428 , n11273 , n7949 );
    or g9744 ( n9031 , n5225 , n21652 );
    xnor g9745 ( n19222 , n25352 , n26823 );
    not g9746 ( n79 , n22970 );
    nor g9747 ( n12575 , n26673 , n15539 );
    or g9748 ( n5490 , n18391 , n16421 );
    or g9749 ( n26811 , n572 , n21076 );
    or g9750 ( n16732 , n15608 , n24423 );
    xnor g9751 ( n13926 , n11954 , n9593 );
    or g9752 ( n26936 , n26990 , n25012 );
    or g9753 ( n15116 , n11707 , n15214 );
    and g9754 ( n23606 , n4696 , n8515 );
    not g9755 ( n6705 , n8079 );
    not g9756 ( n16443 , n6154 );
    xnor g9757 ( n21986 , n11932 , n20720 );
    or g9758 ( n22279 , n18914 , n4629 );
    xnor g9759 ( n19356 , n15500 , n16784 );
    xnor g9760 ( n22497 , n15007 , n14387 );
    not g9761 ( n7685 , n23180 );
    xnor g9762 ( n5350 , n14265 , n2938 );
    and g9763 ( n9955 , n3821 , n24781 );
    and g9764 ( n21040 , n237 , n13688 );
    nor g9765 ( n19513 , n4868 , n25345 );
    and g9766 ( n2384 , n2146 , n212 );
    or g9767 ( n8793 , n10357 , n20621 );
    xnor g9768 ( n3596 , n14130 , n23463 );
    or g9769 ( n1338 , n2522 , n15764 );
    or g9770 ( n25625 , n6764 , n5328 );
    or g9771 ( n14427 , n25400 , n25975 );
    not g9772 ( n24580 , n25739 );
    xnor g9773 ( n597 , n16513 , n6999 );
    nor g9774 ( n26603 , n9983 , n16173 );
    not g9775 ( n5030 , n9559 );
    and g9776 ( n24126 , n5075 , n682 );
    or g9777 ( n25753 , n23818 , n9360 );
    or g9778 ( n25488 , n16943 , n22264 );
    xnor g9779 ( n17843 , n13944 , n7759 );
    xnor g9780 ( n11792 , n11789 , n26107 );
    or g9781 ( n8081 , n2341 , n24620 );
    nor g9782 ( n3972 , n9402 , n2439 );
    xnor g9783 ( n14880 , n3578 , n18181 );
    nor g9784 ( n21092 , n19639 , n11207 );
    not g9785 ( n713 , n17235 );
    xnor g9786 ( n2072 , n24921 , n6714 );
    or g9787 ( n5134 , n348 , n6679 );
    and g9788 ( n7188 , n15545 , n16461 );
    nor g9789 ( n21621 , n27037 , n17605 );
    xnor g9790 ( n24399 , n15046 , n1156 );
    xnor g9791 ( n9963 , n10306 , n3710 );
    or g9792 ( n13823 , n3136 , n5752 );
    nor g9793 ( n23979 , n15023 , n10446 );
    xnor g9794 ( n1691 , n12453 , n14762 );
    or g9795 ( n5137 , n1426 , n10105 );
    xnor g9796 ( n21451 , n24544 , n657 );
    xnor g9797 ( n24881 , n12751 , n7798 );
    nor g9798 ( n3664 , n19025 , n16482 );
    xnor g9799 ( n7924 , n21791 , n22262 );
    or g9800 ( n15962 , n8740 , n19638 );
    xnor g9801 ( n18686 , n15405 , n2223 );
    not g9802 ( n3776 , n22399 );
    or g9803 ( n13175 , n12642 , n5508 );
    nor g9804 ( n19760 , n6492 , n9523 );
    or g9805 ( n20760 , n16091 , n3012 );
    xnor g9806 ( n19791 , n1584 , n2743 );
    or g9807 ( n24333 , n1658 , n384 );
    and g9808 ( n22992 , n5854 , n24066 );
    nor g9809 ( n9659 , n27149 , n15414 );
    xnor g9810 ( n16469 , n15182 , n17351 );
    xnor g9811 ( n13189 , n4563 , n23295 );
    nor g9812 ( n20518 , n9934 , n2272 );
    xnor g9813 ( n13722 , n4827 , n15316 );
    or g9814 ( n15505 , n23457 , n11006 );
    nor g9815 ( n6623 , n24919 , n25261 );
    or g9816 ( n23282 , n3942 , n26328 );
    or g9817 ( n23785 , n13635 , n13067 );
    or g9818 ( n25801 , n1326 , n2854 );
    and g9819 ( n587 , n7801 , n8548 );
    or g9820 ( n6878 , n2628 , n22554 );
    or g9821 ( n17057 , n26895 , n2387 );
    or g9822 ( n1363 , n20365 , n22571 );
    or g9823 ( n7707 , n12289 , n552 );
    or g9824 ( n22117 , n21609 , n20763 );
    xnor g9825 ( n20947 , n22363 , n27065 );
    and g9826 ( n16785 , n19659 , n6646 );
    xnor g9827 ( n1419 , n2842 , n23678 );
    or g9828 ( n14667 , n26314 , n14443 );
    or g9829 ( n14433 , n22413 , n23302 );
    or g9830 ( n23349 , n23129 , n9577 );
    and g9831 ( n6316 , n9794 , n8503 );
    or g9832 ( n17165 , n23164 , n16771 );
    or g9833 ( n10056 , n3324 , n8612 );
    not g9834 ( n16774 , n26077 );
    xnor g9835 ( n7944 , n12040 , n21085 );
    nor g9836 ( n3817 , n17423 , n8614 );
    or g9837 ( n12828 , n2805 , n1524 );
    and g9838 ( n20874 , n5696 , n7871 );
    and g9839 ( n23952 , n21054 , n21808 );
    not g9840 ( n7168 , n18745 );
    or g9841 ( n5497 , n8347 , n9019 );
    xnor g9842 ( n847 , n5421 , n13021 );
    or g9843 ( n9495 , n12973 , n15867 );
    and g9844 ( n24448 , n13084 , n14212 );
    and g9845 ( n3754 , n25305 , n16749 );
    xnor g9846 ( n17662 , n24818 , n3981 );
    xnor g9847 ( n26016 , n16778 , n18691 );
    xnor g9848 ( n25008 , n13577 , n11374 );
    xnor g9849 ( n11119 , n15696 , n2109 );
    xnor g9850 ( n13853 , n25727 , n4253 );
    or g9851 ( n19537 , n3114 , n20347 );
    xnor g9852 ( n14548 , n1682 , n18157 );
    nor g9853 ( n361 , n13490 , n15769 );
    or g9854 ( n24328 , n1163 , n5668 );
    not g9855 ( n5806 , n5787 );
    and g9856 ( n15414 , n952 , n3647 );
    nor g9857 ( n1110 , n2858 , n977 );
    xnor g9858 ( n4158 , n3861 , n2809 );
    or g9859 ( n15825 , n25021 , n20137 );
    or g9860 ( n653 , n20964 , n18345 );
    xnor g9861 ( n26743 , n4435 , n274 );
    xnor g9862 ( n9952 , n11830 , n13775 );
    or g9863 ( n24931 , n14260 , n4268 );
    and g9864 ( n12286 , n19100 , n12074 );
    not g9865 ( n12317 , n3186 );
    not g9866 ( n24008 , n8255 );
    or g9867 ( n17096 , n27183 , n23939 );
    nor g9868 ( n18992 , n11901 , n4938 );
    or g9869 ( n25542 , n21117 , n1112 );
    and g9870 ( n14871 , n5654 , n17482 );
    nor g9871 ( n4645 , n16949 , n3919 );
    nor g9872 ( n22216 , n23285 , n25704 );
    not g9873 ( n18838 , n15058 );
    xnor g9874 ( n14324 , n19128 , n7440 );
    nor g9875 ( n26897 , n12962 , n1960 );
    or g9876 ( n6860 , n8101 , n21912 );
    xnor g9877 ( n12632 , n196 , n9460 );
    not g9878 ( n25282 , n3279 );
    or g9879 ( n24548 , n24603 , n13022 );
    or g9880 ( n7843 , n24059 , n2741 );
    or g9881 ( n26734 , n1635 , n1592 );
    or g9882 ( n22689 , n11847 , n1247 );
    and g9883 ( n25112 , n21593 , n7787 );
    nor g9884 ( n19717 , n24072 , n14312 );
    not g9885 ( n12889 , n4956 );
    or g9886 ( n22140 , n2251 , n20549 );
    not g9887 ( n1364 , n17815 );
    not g9888 ( n944 , n17940 );
    nor g9889 ( n5221 , n16590 , n26090 );
    xnor g9890 ( n1196 , n8725 , n4077 );
    not g9891 ( n5165 , n24298 );
    nor g9892 ( n17838 , n16840 , n8302 );
    xnor g9893 ( n21943 , n2157 , n26136 );
    or g9894 ( n6274 , n19531 , n21322 );
    xnor g9895 ( n13407 , n15330 , n16595 );
    and g9896 ( n4144 , n15636 , n18255 );
    not g9897 ( n12887 , n24677 );
    and g9898 ( n8748 , n15100 , n11793 );
    xnor g9899 ( n2105 , n5632 , n16895 );
    xnor g9900 ( n16258 , n10749 , n7066 );
    xnor g9901 ( n3041 , n18504 , n11630 );
    xnor g9902 ( n22160 , n24700 , n26180 );
    or g9903 ( n23991 , n13571 , n26028 );
    or g9904 ( n10282 , n24150 , n7919 );
    xnor g9905 ( n3484 , n21424 , n14767 );
    not g9906 ( n20316 , n11497 );
    nor g9907 ( n1806 , n16166 , n10407 );
    or g9908 ( n2977 , n18673 , n20953 );
    xnor g9909 ( n7061 , n12681 , n577 );
    or g9910 ( n14503 , n15504 , n5441 );
    xor g9911 ( n4310 , n286 , n6294 );
    and g9912 ( n11908 , n10935 , n1711 );
    or g9913 ( n19782 , n1198 , n8593 );
    xnor g9914 ( n5633 , n21600 , n14261 );
    or g9915 ( n19178 , n18444 , n17028 );
    or g9916 ( n6674 , n2031 , n21369 );
    not g9917 ( n24021 , n27082 );
    or g9918 ( n4948 , n24605 , n10524 );
    not g9919 ( n17067 , n20528 );
    xnor g9920 ( n9761 , n25093 , n10315 );
    not g9921 ( n23843 , n15723 );
    nor g9922 ( n1866 , n24327 , n663 );
    or g9923 ( n4101 , n23281 , n20557 );
    not g9924 ( n7455 , n22895 );
    xnor g9925 ( n10780 , n6305 , n1691 );
    not g9926 ( n23012 , n10082 );
    xnor g9927 ( n7072 , n6181 , n4590 );
    xnor g9928 ( n6038 , n25623 , n145 );
    xnor g9929 ( n2901 , n8087 , n2041 );
    and g9930 ( n24663 , n12932 , n22930 );
    and g9931 ( n24062 , n3915 , n17411 );
    xnor g9932 ( n23790 , n1350 , n13368 );
    nor g9933 ( n21486 , n14226 , n1255 );
    xnor g9934 ( n23660 , n4642 , n17658 );
    xnor g9935 ( n14381 , n10722 , n3893 );
    xnor g9936 ( n16353 , n9911 , n4120 );
    xnor g9937 ( n8594 , n16016 , n21797 );
    or g9938 ( n4612 , n2180 , n20848 );
    or g9939 ( n22430 , n27089 , n12657 );
    not g9940 ( n21038 , n13714 );
    not g9941 ( n1652 , n12646 );
    xnor g9942 ( n14294 , n3021 , n973 );
    not g9943 ( n16483 , n7802 );
    or g9944 ( n23922 , n25663 , n647 );
    or g9945 ( n12268 , n21632 , n7751 );
    nor g9946 ( n19462 , n24044 , n12657 );
    not g9947 ( n27057 , n7991 );
    xnor g9948 ( n5329 , n18303 , n18558 );
    or g9949 ( n18984 , n17717 , n21953 );
    or g9950 ( n4122 , n3984 , n18251 );
    not g9951 ( n13591 , n268 );
    not g9952 ( n10025 , n21140 );
    not g9953 ( n8895 , n8455 );
    xnor g9954 ( n11960 , n3349 , n6397 );
    or g9955 ( n14854 , n10365 , n2951 );
    and g9956 ( n21018 , n11434 , n5322 );
    xnor g9957 ( n15922 , n22852 , n5236 );
    nor g9958 ( n22000 , n2421 , n5337 );
    or g9959 ( n18491 , n23426 , n25885 );
    not g9960 ( n6943 , n16212 );
    and g9961 ( n24406 , n6708 , n16416 );
    or g9962 ( n15751 , n24804 , n7809 );
    not g9963 ( n11499 , n5599 );
    xnor g9964 ( n18691 , n13907 , n2858 );
    not g9965 ( n16755 , n1222 );
    or g9966 ( n13772 , n1490 , n9253 );
    not g9967 ( n6270 , n19836 );
    and g9968 ( n21901 , n12392 , n20648 );
    or g9969 ( n22937 , n20389 , n2864 );
    and g9970 ( n7795 , n7103 , n17849 );
    xnor g9971 ( n5634 , n467 , n27108 );
    or g9972 ( n12073 , n306 , n26307 );
    not g9973 ( n17447 , n15972 );
    or g9974 ( n10870 , n12306 , n26545 );
    or g9975 ( n503 , n6753 , n23529 );
    xnor g9976 ( n652 , n5 , n8255 );
    nor g9977 ( n2339 , n17098 , n14273 );
    and g9978 ( n19581 , n14088 , n23826 );
    xnor g9979 ( n12890 , n26528 , n12888 );
    xnor g9980 ( n7039 , n16465 , n5449 );
    not g9981 ( n22491 , n23650 );
    nor g9982 ( n24607 , n18537 , n24617 );
    and g9983 ( n272 , n17822 , n10607 );
    and g9984 ( n20502 , n12702 , n348 );
    or g9985 ( n18104 , n10606 , n24743 );
    or g9986 ( n18955 , n9233 , n15108 );
    and g9987 ( n18207 , n8782 , n18643 );
    nor g9988 ( n3490 , n25270 , n1339 );
    or g9989 ( n7459 , n15422 , n2908 );
    and g9990 ( n24331 , n21129 , n15159 );
    nor g9991 ( n8700 , n4518 , n12990 );
    xnor g9992 ( n9559 , n9437 , n17720 );
    nor g9993 ( n26333 , n14601 , n25297 );
    or g9994 ( n443 , n14569 , n12004 );
    nor g9995 ( n15358 , n4181 , n2633 );
    not g9996 ( n17379 , n8402 );
    xnor g9997 ( n6345 , n16038 , n23901 );
    and g9998 ( n7617 , n2175 , n4484 );
    not g9999 ( n20133 , n4119 );
    or g10000 ( n16260 , n10401 , n17437 );
    not g10001 ( n14647 , n24679 );
    or g10002 ( n21769 , n16813 , n11894 );
    nor g10003 ( n12451 , n18649 , n3984 );
    not g10004 ( n6515 , n26017 );
    or g10005 ( n4788 , n22612 , n12360 );
    or g10006 ( n486 , n22315 , n23877 );
    xnor g10007 ( n8994 , n14791 , n9557 );
    not g10008 ( n7374 , n3213 );
    xnor g10009 ( n6437 , n2905 , n6807 );
    or g10010 ( n25782 , n16884 , n5250 );
    and g10011 ( n4422 , n20398 , n1517 );
    and g10012 ( n24614 , n21824 , n11877 );
    or g10013 ( n12977 , n4977 , n11320 );
    not g10014 ( n17316 , n10124 );
    and g10015 ( n8591 , n13302 , n11202 );
    or g10016 ( n26121 , n15269 , n19377 );
    and g10017 ( n7282 , n17020 , n17034 );
    or g10018 ( n26998 , n16203 , n17816 );
    and g10019 ( n22628 , n12233 , n25392 );
    or g10020 ( n3797 , n10622 , n24166 );
    xnor g10021 ( n13850 , n23761 , n19040 );
    not g10022 ( n1973 , n26545 );
    nor g10023 ( n19838 , n16351 , n13549 );
    xnor g10024 ( n25688 , n22836 , n15636 );
    not g10025 ( n25737 , n10667 );
    xnor g10026 ( n9787 , n17978 , n10650 );
    nor g10027 ( n4697 , n12386 , n2696 );
    xnor g10028 ( n20397 , n20044 , n7421 );
    not g10029 ( n4149 , n22492 );
    or g10030 ( n10519 , n8492 , n20528 );
    not g10031 ( n26299 , n15970 );
    or g10032 ( n10935 , n10832 , n8352 );
    and g10033 ( n24779 , n2277 , n26037 );
    xnor g10034 ( n9046 , n11820 , n11277 );
    xnor g10035 ( n26529 , n23689 , n24198 );
    not g10036 ( n10037 , n1293 );
    not g10037 ( n15639 , n4467 );
    xnor g10038 ( n11246 , n24799 , n22492 );
    or g10039 ( n23301 , n24962 , n5644 );
    nor g10040 ( n6304 , n13677 , n26752 );
    or g10041 ( n21003 , n1781 , n26045 );
    or g10042 ( n20503 , n26000 , n12137 );
    xnor g10043 ( n16034 , n23122 , n12587 );
    xnor g10044 ( n15462 , n7086 , n20462 );
    or g10045 ( n9866 , n8198 , n11150 );
    or g10046 ( n6712 , n218 , n4605 );
    or g10047 ( n19723 , n16799 , n25148 );
    and g10048 ( n10081 , n4993 , n9994 );
    or g10049 ( n17965 , n7254 , n9599 );
    xnor g10050 ( n12606 , n9105 , n4449 );
    or g10051 ( n7398 , n3029 , n16348 );
    xnor g10052 ( n6477 , n19581 , n12848 );
    not g10053 ( n14145 , n1689 );
    nor g10054 ( n25716 , n26162 , n21386 );
    nor g10055 ( n11244 , n7168 , n17547 );
    and g10056 ( n18656 , n3137 , n2838 );
    or g10057 ( n6166 , n5460 , n7668 );
    not g10058 ( n12924 , n3843 );
    xnor g10059 ( n21893 , n23862 , n4854 );
    xnor g10060 ( n22513 , n18008 , n14230 );
    or g10061 ( n3822 , n16359 , n13257 );
    or g10062 ( n24234 , n405 , n26109 );
    or g10063 ( n18932 , n6910 , n25563 );
    xnor g10064 ( n20384 , n24422 , n4319 );
    nor g10065 ( n24019 , n21272 , n3203 );
    and g10066 ( n22405 , n21227 , n19813 );
    or g10067 ( n25573 , n23288 , n3055 );
    xnor g10068 ( n18437 , n23780 , n25033 );
    xnor g10069 ( n16957 , n7652 , n16559 );
    not g10070 ( n14625 , n16608 );
    and g10071 ( n5558 , n22310 , n19209 );
    xnor g10072 ( n17637 , n3015 , n21272 );
    not g10073 ( n5338 , n13941 );
    not g10074 ( n21004 , n22413 );
    and g10075 ( n7869 , n21282 , n19246 );
    xnor g10076 ( n14092 , n9942 , n2210 );
    nor g10077 ( n13488 , n7693 , n3909 );
    xnor g10078 ( n17229 , n5886 , n1839 );
    xnor g10079 ( n11101 , n13211 , n16809 );
    or g10080 ( n17267 , n20527 , n2525 );
    nor g10081 ( n15790 , n19429 , n23519 );
    xnor g10082 ( n27021 , n18283 , n6924 );
    not g10083 ( n11958 , n12081 );
    and g10084 ( n20560 , n26660 , n17826 );
    or g10085 ( n16372 , n2967 , n18907 );
    xnor g10086 ( n18708 , n13213 , n16011 );
    xnor g10087 ( n18905 , n12502 , n4320 );
    not g10088 ( n20271 , n17166 );
    xnor g10089 ( n9900 , n835 , n20826 );
    or g10090 ( n20398 , n24305 , n8823 );
    or g10091 ( n26164 , n17911 , n17674 );
    xnor g10092 ( n15649 , n20470 , n4590 );
    nor g10093 ( n20864 , n16928 , n19940 );
    not g10094 ( n9733 , n22795 );
    xnor g10095 ( n8084 , n26950 , n1945 );
    not g10096 ( n10620 , n3319 );
    or g10097 ( n7633 , n13298 , n25231 );
    xnor g10098 ( n3895 , n966 , n12446 );
    nor g10099 ( n27167 , n25139 , n15636 );
    nor g10100 ( n10416 , n25724 , n24503 );
    and g10101 ( n11027 , n26107 , n21636 );
    xnor g10102 ( n12081 , n9109 , n21354 );
    or g10103 ( n8157 , n24005 , n15528 );
    or g10104 ( n8737 , n26660 , n26810 );
    xnor g10105 ( n26930 , n14890 , n16375 );
    xnor g10106 ( n10737 , n22290 , n12562 );
    and g10107 ( n26409 , n8571 , n10872 );
    or g10108 ( n16835 , n4917 , n13841 );
    and g10109 ( n25554 , n13750 , n20024 );
    xnor g10110 ( n2279 , n2123 , n1996 );
    or g10111 ( n14027 , n12815 , n8441 );
    xnor g10112 ( n9341 , n19514 , n19228 );
    and g10113 ( n13711 , n3460 , n16667 );
    not g10114 ( n3257 , n14163 );
    xnor g10115 ( n23503 , n7010 , n13851 );
    and g10116 ( n22751 , n9514 , n17204 );
    xnor g10117 ( n8587 , n26992 , n7437 );
    xnor g10118 ( n22457 , n9200 , n18758 );
    or g10119 ( n6376 , n18850 , n15153 );
    not g10120 ( n17195 , n4583 );
    and g10121 ( n297 , n4592 , n24502 );
    xnor g10122 ( n5744 , n11579 , n8067 );
    or g10123 ( n9443 , n22363 , n17291 );
    xnor g10124 ( n11955 , n24135 , n20291 );
    or g10125 ( n15130 , n11997 , n18798 );
    nor g10126 ( n20732 , n16573 , n26894 );
    not g10127 ( n20508 , n14417 );
    or g10128 ( n12678 , n6306 , n25396 );
    nor g10129 ( n27190 , n23559 , n12048 );
    nor g10130 ( n7501 , n18451 , n13081 );
    and g10131 ( n20386 , n20226 , n21136 );
    nor g10132 ( n3396 , n3668 , n2246 );
    xnor g10133 ( n10950 , n2570 , n10250 );
    nor g10134 ( n22576 , n15332 , n8753 );
    and g10135 ( n26880 , n1514 , n6922 );
    xnor g10136 ( n12680 , n4400 , n17739 );
    xnor g10137 ( n22162 , n2884 , n20455 );
    and g10138 ( n26045 , n3991 , n13431 );
    xnor g10139 ( n23467 , n20645 , n21180 );
    or g10140 ( n22239 , n21073 , n502 );
    xnor g10141 ( n22772 , n21564 , n11412 );
    xnor g10142 ( n12177 , n4970 , n2454 );
    nor g10143 ( n23989 , n22602 , n12257 );
    xnor g10144 ( n11900 , n15204 , n12956 );
    or g10145 ( n20940 , n2930 , n12885 );
    xnor g10146 ( n23857 , n17664 , n5115 );
    or g10147 ( n4389 , n26833 , n22875 );
    nor g10148 ( n22288 , n12068 , n18535 );
    and g10149 ( n14299 , n26347 , n12393 );
    and g10150 ( n7646 , n17245 , n8506 );
    xnor g10151 ( n15447 , n4474 , n23215 );
    not g10152 ( n20509 , n26174 );
    xnor g10153 ( n8437 , n373 , n737 );
    not g10154 ( n23211 , n7876 );
    not g10155 ( n23273 , n18924 );
    xnor g10156 ( n4408 , n2432 , n11137 );
    and g10157 ( n4821 , n8737 , n7699 );
    nor g10158 ( n796 , n24612 , n9770 );
    and g10159 ( n24741 , n16008 , n24287 );
    xnor g10160 ( n15234 , n26629 , n18690 );
    xnor g10161 ( n25575 , n23357 , n26958 );
    or g10162 ( n14853 , n7198 , n16439 );
    not g10163 ( n14979 , n25797 );
    or g10164 ( n21699 , n25926 , n20385 );
    or g10165 ( n18456 , n17458 , n17265 );
    xnor g10166 ( n10694 , n17309 , n2096 );
    or g10167 ( n26014 , n7670 , n8227 );
    xnor g10168 ( n14201 , n13960 , n10405 );
    not g10169 ( n21780 , n12744 );
    nor g10170 ( n19214 , n22194 , n6104 );
    not g10171 ( n18126 , n14504 );
    or g10172 ( n6507 , n23365 , n12770 );
    or g10173 ( n8392 , n13092 , n19237 );
    or g10174 ( n18699 , n10810 , n17575 );
    and g10175 ( n26615 , n23514 , n15132 );
    nor g10176 ( n20652 , n15109 , n8677 );
    and g10177 ( n14838 , n19788 , n1468 );
    or g10178 ( n21251 , n3914 , n1717 );
    xnor g10179 ( n4822 , n4914 , n19338 );
    and g10180 ( n8365 , n14213 , n14847 );
    not g10181 ( n11552 , n24080 );
    nor g10182 ( n17121 , n17973 , n26009 );
    or g10183 ( n6066 , n15905 , n27118 );
    or g10184 ( n18358 , n1790 , n20660 );
    and g10185 ( n12375 , n22573 , n8400 );
    nor g10186 ( n8112 , n20955 , n24322 );
    not g10187 ( n17261 , n3786 );
    xnor g10188 ( n13965 , n17415 , n7593 );
    or g10189 ( n24894 , n3180 , n10249 );
    or g10190 ( n18748 , n7825 , n8511 );
    or g10191 ( n23764 , n11659 , n4928 );
    or g10192 ( n16992 , n7769 , n15245 );
    and g10193 ( n24118 , n5167 , n4170 );
    xnor g10194 ( n21293 , n23136 , n15779 );
    or g10195 ( n23944 , n8642 , n12172 );
    nor g10196 ( n22007 , n16830 , n25688 );
    not g10197 ( n5855 , n25069 );
    and g10198 ( n17313 , n9434 , n5563 );
    or g10199 ( n26842 , n21988 , n8380 );
    xnor g10200 ( n10095 , n18262 , n22588 );
    or g10201 ( n16935 , n14145 , n20036 );
    not g10202 ( n5970 , n17085 );
    not g10203 ( n14955 , n3056 );
    or g10204 ( n23338 , n2212 , n21393 );
    xnor g10205 ( n10905 , n4999 , n27017 );
    not g10206 ( n12961 , n16846 );
    and g10207 ( n1617 , n17789 , n1731 );
    xnor g10208 ( n12228 , n24986 , n9 );
    not g10209 ( n9303 , n781 );
    not g10210 ( n2110 , n7476 );
    or g10211 ( n4211 , n9081 , n19597 );
    and g10212 ( n24011 , n13771 , n14911 );
    xnor g10213 ( n7257 , n3591 , n647 );
    xnor g10214 ( n26251 , n16033 , n15946 );
    xnor g10215 ( n9737 , n24787 , n906 );
    xnor g10216 ( n9420 , n4856 , n23323 );
    xnor g10217 ( n9636 , n3049 , n25094 );
    xnor g10218 ( n2233 , n22195 , n1865 );
    or g10219 ( n8651 , n10092 , n11477 );
    and g10220 ( n2521 , n1740 , n4997 );
    or g10221 ( n10068 , n13038 , n11306 );
    not g10222 ( n19 , n8745 );
    or g10223 ( n12241 , n9964 , n4880 );
    and g10224 ( n7184 , n2894 , n22783 );
    or g10225 ( n14308 , n6664 , n4114 );
    not g10226 ( n18298 , n16263 );
    xnor g10227 ( n24928 , n3389 , n4148 );
    nor g10228 ( n17632 , n26107 , n4376 );
    and g10229 ( n22534 , n10471 , n8600 );
    xnor g10230 ( n14355 , n788 , n21780 );
    or g10231 ( n1861 , n18704 , n5317 );
    xnor g10232 ( n4375 , n23734 , n25927 );
    xnor g10233 ( n23685 , n1894 , n3921 );
    and g10234 ( n26466 , n19776 , n18932 );
    not g10235 ( n5685 , n22340 );
    and g10236 ( n26286 , n11601 , n4546 );
    and g10237 ( n13019 , n13325 , n7176 );
    or g10238 ( n26859 , n6206 , n17409 );
    or g10239 ( n26537 , n17230 , n10792 );
    nor g10240 ( n1116 , n10023 , n22715 );
    xnor g10241 ( n2099 , n21757 , n21239 );
    or g10242 ( n7054 , n22750 , n13728 );
    or g10243 ( n3999 , n6212 , n23375 );
    or g10244 ( n20984 , n15259 , n7833 );
    and g10245 ( n12439 , n8631 , n607 );
    or g10246 ( n15246 , n21117 , n22332 );
    and g10247 ( n8707 , n18737 , n15268 );
    and g10248 ( n21848 , n17400 , n21196 );
    or g10249 ( n25531 , n6812 , n14866 );
    and g10250 ( n1727 , n319 , n23032 );
    xnor g10251 ( n17112 , n11098 , n15175 );
    not g10252 ( n144 , n23529 );
    nor g10253 ( n16853 , n27015 , n22993 );
    or g10254 ( n9334 , n18633 , n24647 );
    or g10255 ( n16132 , n6950 , n23275 );
    xnor g10256 ( n15153 , n4157 , n16503 );
    or g10257 ( n1015 , n25524 , n2562 );
    nor g10258 ( n20566 , n7060 , n19976 );
    or g10259 ( n24209 , n4508 , n13843 );
    and g10260 ( n17008 , n22348 , n7482 );
    not g10261 ( n20998 , n11056 );
    or g10262 ( n17282 , n14642 , n23417 );
    xnor g10263 ( n2802 , n23493 , n1222 );
    and g10264 ( n17793 , n12083 , n7989 );
    and g10265 ( n2052 , n19553 , n24195 );
    and g10266 ( n8742 , n6635 , n121 );
    or g10267 ( n24737 , n1404 , n18262 );
    or g10268 ( n11763 , n12767 , n1658 );
    and g10269 ( n17545 , n4621 , n10748 );
    and g10270 ( n4920 , n21527 , n20509 );
    xnor g10271 ( n21024 , n10454 , n102 );
    xnor g10272 ( n13830 , n24170 , n18537 );
    or g10273 ( n2414 , n17069 , n19446 );
    xnor g10274 ( n15495 , n21434 , n2715 );
    or g10275 ( n13020 , n4510 , n24741 );
    nor g10276 ( n22482 , n23609 , n14335 );
    or g10277 ( n26114 , n7480 , n8122 );
    or g10278 ( n2394 , n14100 , n2284 );
    or g10279 ( n14325 , n10051 , n11047 );
    not g10280 ( n19989 , n16097 );
    or g10281 ( n7294 , n15 , n26706 );
    xnor g10282 ( n18526 , n1028 , n1994 );
    nor g10283 ( n7560 , n12930 , n22084 );
    or g10284 ( n16036 , n8886 , n2898 );
    not g10285 ( n12123 , n19893 );
    and g10286 ( n19491 , n13042 , n12721 );
    buf g10287 ( n9502 , n75 );
    xnor g10288 ( n14905 , n7561 , n3443 );
    and g10289 ( n5933 , n4957 , n22688 );
    or g10290 ( n25386 , n3419 , n25554 );
    not g10291 ( n22095 , n17690 );
    and g10292 ( n17194 , n24522 , n4450 );
    not g10293 ( n17728 , n12964 );
    xnor g10294 ( n14005 , n4307 , n10964 );
    or g10295 ( n3453 , n17789 , n1731 );
    or g10296 ( n1174 , n15799 , n12496 );
    not g10297 ( n23707 , n8497 );
    and g10298 ( n21955 , n17535 , n6552 );
    not g10299 ( n17502 , n19477 );
    not g10300 ( n14980 , n24169 );
    xnor g10301 ( n12060 , n11118 , n4199 );
    xnor g10302 ( n11779 , n13960 , n12990 );
    or g10303 ( n9016 , n17708 , n2769 );
    nor g10304 ( n17440 , n24584 , n13802 );
    xnor g10305 ( n10924 , n18703 , n22530 );
    xnor g10306 ( n5789 , n9307 , n21963 );
    xnor g10307 ( n24219 , n22729 , n18744 );
    or g10308 ( n10040 , n4856 , n14455 );
    or g10309 ( n6425 , n2613 , n20851 );
    xnor g10310 ( n8901 , n8518 , n17677 );
    or g10311 ( n4423 , n6385 , n8844 );
    or g10312 ( n2292 , n9298 , n17339 );
    and g10313 ( n20646 , n6801 , n16395 );
    xnor g10314 ( n1760 , n20980 , n4516 );
    and g10315 ( n25118 , n8899 , n20873 );
    or g10316 ( n4556 , n3014 , n23630 );
    or g10317 ( n5622 , n23592 , n23463 );
    or g10318 ( n13394 , n22658 , n4006 );
    xnor g10319 ( n12826 , n14365 , n11993 );
    xnor g10320 ( n20012 , n26822 , n22404 );
    and g10321 ( n12672 , n24434 , n20585 );
    or g10322 ( n12164 , n333 , n4798 );
    or g10323 ( n9623 , n22206 , n9559 );
    or g10324 ( n24110 , n17348 , n15335 );
    nor g10325 ( n730 , n12385 , n4749 );
    and g10326 ( n19973 , n24209 , n7671 );
    or g10327 ( n18329 , n3409 , n2310 );
    and g10328 ( n15568 , n26390 , n1489 );
    not g10329 ( n10146 , n25643 );
    not g10330 ( n17088 , n23660 );
    or g10331 ( n25910 , n24850 , n16083 );
    not g10332 ( n10533 , n18434 );
    or g10333 ( n22368 , n6905 , n11587 );
    or g10334 ( n23278 , n767 , n8806 );
    or g10335 ( n9265 , n18966 , n19796 );
    nor g10336 ( n736 , n23030 , n20829 );
    and g10337 ( n24063 , n26393 , n13267 );
    and g10338 ( n23029 , n21749 , n11676 );
    nor g10339 ( n1356 , n19033 , n17037 );
    nor g10340 ( n2805 , n1406 , n1978 );
    and g10341 ( n388 , n16014 , n262 );
    xnor g10342 ( n24138 , n6847 , n12070 );
    not g10343 ( n6508 , n14388 );
    and g10344 ( n3736 , n8553 , n15502 );
    or g10345 ( n4991 , n3169 , n8729 );
    and g10346 ( n20401 , n18883 , n25146 );
    or g10347 ( n4216 , n15189 , n24320 );
    or g10348 ( n23774 , n9598 , n21570 );
    not g10349 ( n7619 , n6185 );
    and g10350 ( n18424 , n9099 , n19067 );
    and g10351 ( n15797 , n22374 , n5118 );
    nor g10352 ( n10307 , n21540 , n18768 );
    not g10353 ( n7818 , n5077 );
    not g10354 ( n24090 , n8009 );
    xnor g10355 ( n2383 , n25453 , n18743 );
    and g10356 ( n8547 , n6847 , n2051 );
    or g10357 ( n21026 , n13711 , n26586 );
    or g10358 ( n9061 , n5907 , n24407 );
    xnor g10359 ( n8489 , n25410 , n21000 );
    xnor g10360 ( n4923 , n19628 , n2999 );
    and g10361 ( n18648 , n17616 , n21391 );
    and g10362 ( n8595 , n11961 , n22863 );
    xnor g10363 ( n17362 , n21287 , n25331 );
    or g10364 ( n17748 , n10430 , n18575 );
    nor g10365 ( n18902 , n4695 , n17371 );
    and g10366 ( n16647 , n25274 , n3888 );
    xnor g10367 ( n2150 , n17989 , n20706 );
    or g10368 ( n10348 , n14311 , n6335 );
    or g10369 ( n19554 , n12390 , n9747 );
    xnor g10370 ( n8993 , n1598 , n12041 );
    and g10371 ( n1233 , n25443 , n26761 );
    xnor g10372 ( n5403 , n22005 , n19854 );
    not g10373 ( n23249 , n12739 );
    or g10374 ( n26032 , n9479 , n3506 );
    xnor g10375 ( n23364 , n8472 , n23905 );
    or g10376 ( n1392 , n16952 , n14756 );
    xnor g10377 ( n21164 , n9410 , n8762 );
    xnor g10378 ( n7363 , n5138 , n14669 );
    and g10379 ( n26554 , n4363 , n13097 );
    xnor g10380 ( n4295 , n17935 , n8111 );
    nor g10381 ( n2130 , n1876 , n5675 );
    not g10382 ( n19241 , n5868 );
    or g10383 ( n7821 , n20265 , n23297 );
    nor g10384 ( n9488 , n12288 , n7932 );
    or g10385 ( n313 , n11754 , n19885 );
    or g10386 ( n17024 , n23500 , n4831 );
    not g10387 ( n19373 , n21417 );
    or g10388 ( n10253 , n23064 , n25818 );
    not g10389 ( n3622 , n14957 );
    not g10390 ( n1960 , n11980 );
    or g10391 ( n18588 , n11753 , n19928 );
    and g10392 ( n12536 , n1649 , n165 );
    xnor g10393 ( n696 , n1080 , n16356 );
    not g10394 ( n617 , n12751 );
    xnor g10395 ( n960 , n8386 , n7641 );
    or g10396 ( n6866 , n22767 , n7022 );
    or g10397 ( n4628 , n22626 , n18765 );
    or g10398 ( n9734 , n22935 , n12881 );
    or g10399 ( n16169 , n16029 , n12088 );
    or g10400 ( n309 , n11569 , n4921 );
    xnor g10401 ( n6881 , n26939 , n10057 );
    xnor g10402 ( n11352 , n1124 , n25999 );
    or g10403 ( n6516 , n12097 , n9000 );
    not g10404 ( n1232 , n23019 );
    xnor g10405 ( n11508 , n24529 , n18171 );
    not g10406 ( n10743 , n12204 );
    xnor g10407 ( n494 , n15112 , n26035 );
    nor g10408 ( n1423 , n11901 , n17911 );
    not g10409 ( n14718 , n17911 );
    and g10410 ( n11085 , n705 , n20047 );
    or g10411 ( n8039 , n5335 , n5143 );
    or g10412 ( n22529 , n11605 , n24399 );
    not g10413 ( n24630 , n25556 );
    not g10414 ( n22755 , n3169 );
    and g10415 ( n4245 , n25556 , n12169 );
    or g10416 ( n19937 , n26723 , n2205 );
    nor g10417 ( n9309 , n11580 , n1799 );
    or g10418 ( n16488 , n8553 , n15502 );
    nor g10419 ( n5262 , n990 , n19097 );
    xnor g10420 ( n11063 , n19773 , n2885 );
    or g10421 ( n5879 , n14830 , n6468 );
    not g10422 ( n15074 , n18687 );
    and g10423 ( n12261 , n6094 , n12877 );
    xnor g10424 ( n18344 , n17233 , n8160 );
    xnor g10425 ( n24228 , n15656 , n27177 );
    and g10426 ( n1042 , n16927 , n16652 );
    not g10427 ( n3407 , n10199 );
    nor g10428 ( n21119 , n6883 , n14681 );
    xnor g10429 ( n25918 , n24123 , n9377 );
    or g10430 ( n17336 , n18496 , n20201 );
    nor g10431 ( n727 , n17295 , n14289 );
    and g10432 ( n23197 , n25545 , n9585 );
    xnor g10433 ( n3319 , n11142 , n20703 );
    not g10434 ( n2141 , n4100 );
    or g10435 ( n25623 , n17331 , n11291 );
    xnor g10436 ( n11507 , n586 , n7566 );
    xnor g10437 ( n23915 , n22715 , n25900 );
    not g10438 ( n10357 , n3623 );
    not g10439 ( n698 , n20840 );
    not g10440 ( n8013 , n9135 );
    and g10441 ( n22759 , n2262 , n11735 );
    or g10442 ( n171 , n15974 , n2593 );
    or g10443 ( n2170 , n15652 , n8151 );
    xnor g10444 ( n13317 , n4896 , n2146 );
    xnor g10445 ( n4278 , n903 , n996 );
    xnor g10446 ( n3120 , n12504 , n24975 );
    xnor g10447 ( n5357 , n1349 , n23065 );
    and g10448 ( n12995 , n3695 , n10953 );
    nor g10449 ( n381 , n528 , n25471 );
    not g10450 ( n2914 , n6381 );
    or g10451 ( n25880 , n1058 , n2521 );
    xnor g10452 ( n7097 , n5245 , n26893 );
    or g10453 ( n2843 , n17887 , n18417 );
    and g10454 ( n22218 , n3450 , n10293 );
    xnor g10455 ( n6532 , n20700 , n26510 );
    or g10456 ( n562 , n5931 , n25711 );
    nor g10457 ( n3140 , n2036 , n12391 );
    and g10458 ( n2474 , n6717 , n24912 );
    xnor g10459 ( n17432 , n38 , n19098 );
    xnor g10460 ( n20927 , n18624 , n21505 );
    and g10461 ( n11754 , n9598 , n21570 );
    xnor g10462 ( n6903 , n23160 , n8067 );
    or g10463 ( n24751 , n24381 , n40 );
    xnor g10464 ( n7438 , n4108 , n26689 );
    xnor g10465 ( n13998 , n19797 , n3903 );
    and g10466 ( n24854 , n22617 , n19091 );
    or g10467 ( n6656 , n3538 , n23515 );
    xnor g10468 ( n25293 , n4226 , n4548 );
    nor g10469 ( n24610 , n4490 , n21846 );
    nor g10470 ( n14442 , n6309 , n17572 );
    not g10471 ( n12267 , n16949 );
    xnor g10472 ( n19389 , n19809 , n25223 );
    or g10473 ( n22164 , n5719 , n17911 );
    xnor g10474 ( n18967 , n13460 , n11455 );
    or g10475 ( n26464 , n6452 , n8475 );
    or g10476 ( n5613 , n26450 , n23109 );
    nor g10477 ( n6882 , n22736 , n12741 );
    xnor g10478 ( n10124 , n26283 , n16847 );
    nor g10479 ( n20913 , n1587 , n16524 );
    xnor g10480 ( n8570 , n16024 , n8355 );
    or g10481 ( n8970 , n1611 , n6718 );
    not g10482 ( n26925 , n10481 );
    xnor g10483 ( n14839 , n4538 , n8776 );
    xnor g10484 ( n21154 , n1610 , n18685 );
    and g10485 ( n20702 , n22422 , n18648 );
    and g10486 ( n8783 , n12601 , n591 );
    and g10487 ( n12137 , n8045 , n13779 );
    and g10488 ( n17551 , n25974 , n6963 );
    xnor g10489 ( n6918 , n10169 , n19132 );
    and g10490 ( n13475 , n15871 , n10572 );
    nor g10491 ( n19761 , n8614 , n25972 );
    and g10492 ( n2134 , n5089 , n6059 );
    or g10493 ( n13363 , n15854 , n4821 );
    and g10494 ( n20265 , n17251 , n23967 );
    not g10495 ( n27150 , n13041 );
    xnor g10496 ( n4141 , n15087 , n15147 );
    nor g10497 ( n6883 , n21288 , n26522 );
    xnor g10498 ( n14172 , n7374 , n13613 );
    xnor g10499 ( n12772 , n23467 , n6030 );
    and g10500 ( n11979 , n26356 , n3838 );
    and g10501 ( n12726 , n965 , n7483 );
    or g10502 ( n5215 , n19239 , n4513 );
    xnor g10503 ( n5385 , n18710 , n5621 );
    xnor g10504 ( n23630 , n22785 , n3638 );
    not g10505 ( n15633 , n7285 );
    not g10506 ( n26015 , n11986 );
    or g10507 ( n20729 , n17116 , n7717 );
    not g10508 ( n15287 , n16581 );
    xnor g10509 ( n1019 , n4639 , n7506 );
    xnor g10510 ( n27044 , n19352 , n12593 );
    nor g10511 ( n5831 , n13789 , n6971 );
    or g10512 ( n12823 , n658 , n2723 );
    and g10513 ( n9311 , n17126 , n18112 );
    and g10514 ( n10912 , n12853 , n4535 );
    xnor g10515 ( n9898 , n20564 , n8721 );
    xnor g10516 ( n21907 , n7316 , n25068 );
    xnor g10517 ( n15816 , n18476 , n12144 );
    xnor g10518 ( n11720 , n8431 , n8244 );
    and g10519 ( n4510 , n10448 , n6471 );
    not g10520 ( n4749 , n13022 );
    or g10521 ( n3928 , n86 , n11543 );
    or g10522 ( n18182 , n4722 , n14323 );
    or g10523 ( n25177 , n18924 , n12701 );
    and g10524 ( n9447 , n17668 , n11167 );
    xnor g10525 ( n2931 , n27144 , n6774 );
    xnor g10526 ( n5615 , n9069 , n20470 );
    or g10527 ( n25767 , n24659 , n590 );
    nor g10528 ( n22149 , n4360 , n25923 );
    xnor g10529 ( n2226 , n19962 , n7139 );
    and g10530 ( n6989 , n7263 , n24968 );
    and g10531 ( n7947 , n20332 , n20987 );
    and g10532 ( n10730 , n1877 , n7265 );
    or g10533 ( n14349 , n7831 , n6005 );
    or g10534 ( n26481 , n17002 , n18274 );
    not g10535 ( n12652 , n5607 );
    xnor g10536 ( n10235 , n22700 , n9655 );
    and g10537 ( n21923 , n21346 , n19548 );
    not g10538 ( n18920 , n15161 );
    and g10539 ( n9257 , n12702 , n11144 );
    or g10540 ( n8147 , n21652 , n21600 );
    or g10541 ( n13024 , n954 , n6208 );
    and g10542 ( n2837 , n17554 , n11203 );
    not g10543 ( n25004 , n9507 );
    and g10544 ( n9978 , n1611 , n6718 );
    xnor g10545 ( n23605 , n7858 , n21294 );
    xnor g10546 ( n14957 , n6942 , n24953 );
    xor g10547 ( n17089 , n12390 , n6948 );
    or g10548 ( n6621 , n7437 , n26992 );
    nor g10549 ( n21467 , n23678 , n2842 );
    or g10550 ( n14688 , n9950 , n16332 );
    not g10551 ( n26914 , n3730 );
    xnor g10552 ( n15964 , n2978 , n20040 );
    nor g10553 ( n6026 , n16210 , n166 );
    and g10554 ( n13905 , n9639 , n22580 );
    xnor g10555 ( n14886 , n27152 , n15794 );
    and g10556 ( n24500 , n14680 , n8948 );
    and g10557 ( n18891 , n17266 , n25239 );
    or g10558 ( n952 , n26688 , n16727 );
    not g10559 ( n5160 , n14919 );
    and g10560 ( n9732 , n3018 , n16366 );
    and g10561 ( n14238 , n8559 , n9579 );
    xnor g10562 ( n10761 , n16826 , n6636 );
    xnor g10563 ( n721 , n12149 , n1952 );
    xnor g10564 ( n11911 , n12246 , n25204 );
    not g10565 ( n24805 , n964 );
    xnor g10566 ( n21537 , n24390 , n13426 );
    xnor g10567 ( n6006 , n17379 , n16353 );
    or g10568 ( n5129 , n8759 , n20456 );
    nor g10569 ( n12473 , n22289 , n2509 );
    xnor g10570 ( n16683 , n3224 , n7873 );
    buf g10571 ( n7130 , n16541 );
    xnor g10572 ( n19223 , n23204 , n7474 );
    or g10573 ( n700 , n24905 , n6033 );
    nor g10574 ( n25344 , n23936 , n1386 );
    or g10575 ( n17356 , n8324 , n5574 );
    nor g10576 ( n18673 , n8540 , n2399 );
    or g10577 ( n1566 , n24695 , n2088 );
    or g10578 ( n16912 , n17115 , n5675 );
    xnor g10579 ( n19857 , n11302 , n2146 );
    xnor g10580 ( n22191 , n19206 , n11556 );
    xnor g10581 ( n8507 , n8515 , n14599 );
    not g10582 ( n17994 , n16295 );
    xnor g10583 ( n15118 , n18087 , n10350 );
    xnor g10584 ( n23109 , n209 , n1288 );
    xnor g10585 ( n2433 , n11580 , n24620 );
    and g10586 ( n18682 , n10399 , n13322 );
    and g10587 ( n21704 , n12464 , n25352 );
    nor g10588 ( n23182 , n4022 , n9569 );
    or g10589 ( n15377 , n26358 , n1986 );
    or g10590 ( n26576 , n13646 , n16137 );
    xnor g10591 ( n24782 , n5112 , n5417 );
    xnor g10592 ( n25956 , n7466 , n6659 );
    not g10593 ( n990 , n7949 );
    or g10594 ( n22316 , n7841 , n9445 );
    and g10595 ( n17438 , n17470 , n25998 );
    not g10596 ( n24929 , n24990 );
    or g10597 ( n4011 , n3541 , n9219 );
    not g10598 ( n13348 , n10046 );
    xnor g10599 ( n23318 , n10172 , n11104 );
    nor g10600 ( n25227 , n10632 , n1824 );
    not g10601 ( n18850 , n2666 );
    not g10602 ( n5320 , n8025 );
    and g10603 ( n2898 , n3406 , n19126 );
    xnor g10604 ( n8692 , n643 , n22635 );
    or g10605 ( n19250 , n5887 , n10541 );
    xnor g10606 ( n7840 , n26422 , n21747 );
    not g10607 ( n16311 , n26520 );
    xnor g10608 ( n5191 , n16496 , n22456 );
    or g10609 ( n11851 , n24083 , n7409 );
    xnor g10610 ( n8159 , n1491 , n794 );
    not g10611 ( n6262 , n11525 );
    or g10612 ( n18464 , n23737 , n6361 );
    xnor g10613 ( n6174 , n12811 , n3260 );
    or g10614 ( n2159 , n24170 , n23460 );
    or g10615 ( n18249 , n13731 , n24630 );
    xnor g10616 ( n9809 , n7197 , n14609 );
    and g10617 ( n9611 , n13414 , n25233 );
    xnor g10618 ( n8750 , n14008 , n3785 );
    nor g10619 ( n16378 , n14740 , n14698 );
    or g10620 ( n26426 , n4265 , n12995 );
    or g10621 ( n8394 , n16561 , n18139 );
    or g10622 ( n13536 , n9978 , n5598 );
    or g10623 ( n3292 , n4594 , n21348 );
    xnor g10624 ( n18636 , n6917 , n2323 );
    or g10625 ( n22913 , n11959 , n15312 );
    xnor g10626 ( n17623 , n2210 , n16608 );
    xnor g10627 ( n8620 , n4106 , n4943 );
    not g10628 ( n1141 , n17488 );
    xnor g10629 ( n10651 , n2838 , n2438 );
    xnor g10630 ( n3623 , n1824 , n1457 );
    xnor g10631 ( n2734 , n12236 , n19785 );
    and g10632 ( n24743 , n22504 , n2907 );
    xnor g10633 ( n9 , n20517 , n18735 );
    xnor g10634 ( n15929 , n26030 , n20478 );
    xnor g10635 ( n390 , n5678 , n2678 );
    and g10636 ( n12799 , n22911 , n11396 );
    or g10637 ( n11719 , n11473 , n15506 );
    or g10638 ( n14537 , n8358 , n24344 );
    or g10639 ( n5710 , n22492 , n9372 );
    and g10640 ( n4043 , n19677 , n2554 );
    not g10641 ( n19297 , n18024 );
    xnor g10642 ( n9620 , n14361 , n3120 );
    xnor g10643 ( n10639 , n13603 , n6756 );
    not g10644 ( n12356 , n1055 );
    or g10645 ( n15201 , n24164 , n14937 );
    not g10646 ( n8101 , n15241 );
    or g10647 ( n16154 , n6809 , n6847 );
    and g10648 ( n11718 , n4220 , n22869 );
    xnor g10649 ( n8490 , n5927 , n17160 );
    not g10650 ( n24403 , n19177 );
    xnor g10651 ( n20388 , n15351 , n10216 );
    nor g10652 ( n15742 , n632 , n25827 );
    xnor g10653 ( n25538 , n2066 , n20478 );
    not g10654 ( n24603 , n24015 );
    nor g10655 ( n566 , n17784 , n24085 );
    xnor g10656 ( n24446 , n9096 , n485 );
    xnor g10657 ( n923 , n15808 , n4160 );
    xnor g10658 ( n5991 , n16994 , n16521 );
    not g10659 ( n11425 , n23697 );
    and g10660 ( n3769 , n18140 , n7085 );
    and g10661 ( n22166 , n8382 , n7644 );
    nor g10662 ( n15925 , n15271 , n12161 );
    xnor g10663 ( n14384 , n6712 , n5332 );
    xnor g10664 ( n8205 , n6259 , n14838 );
    buf g10665 ( n2694 , n3584 );
    not g10666 ( n27069 , n11224 );
    nor g10667 ( n2927 , n3086 , n18213 );
    or g10668 ( n16864 , n2323 , n6917 );
    not g10669 ( n23746 , n4325 );
    or g10670 ( n3107 , n2612 , n27193 );
    or g10671 ( n3008 , n4102 , n20744 );
    and g10672 ( n22685 , n3283 , n25746 );
    or g10673 ( n4621 , n12002 , n11918 );
    and g10674 ( n11139 , n2542 , n17057 );
    or g10675 ( n23178 , n8155 , n20920 );
    not g10676 ( n16364 , n24599 );
    nor g10677 ( n20016 , n1040 , n12152 );
    nor g10678 ( n8642 , n11533 , n11095 );
    and g10679 ( n6358 , n26787 , n13792 );
    not g10680 ( n23162 , n21235 );
    not g10681 ( n912 , n11719 );
    xnor g10682 ( n22885 , n8910 , n9246 );
    xnor g10683 ( n6249 , n9514 , n3939 );
    or g10684 ( n7951 , n14133 , n7524 );
    or g10685 ( n23756 , n15581 , n5407 );
    xnor g10686 ( n10216 , n17901 , n8430 );
    or g10687 ( n18766 , n26478 , n19721 );
    not g10688 ( n10868 , n21890 );
    or g10689 ( n11636 , n5181 , n11282 );
    nor g10690 ( n16884 , n8328 , n24601 );
    nor g10691 ( n9869 , n13062 , n5341 );
    not g10692 ( n11544 , n19282 );
    and g10693 ( n12901 , n17983 , n10458 );
    xnor g10694 ( n11140 , n16029 , n19228 );
    not g10695 ( n9398 , n15495 );
    xnor g10696 ( n8020 , n2415 , n172 );
    and g10697 ( n22915 , n18828 , n23904 );
    and g10698 ( n3804 , n18675 , n22423 );
    not g10699 ( n14131 , n15220 );
    or g10700 ( n26037 , n16717 , n1817 );
    xnor g10701 ( n22907 , n15306 , n6098 );
    not g10702 ( n22765 , n24935 );
    xnor g10703 ( n10045 , n2964 , n11554 );
    not g10704 ( n2562 , n6513 );
    and g10705 ( n19198 , n7362 , n16143 );
    xnor g10706 ( n16374 , n4128 , n20891 );
    or g10707 ( n18672 , n22212 , n12510 );
    nor g10708 ( n12455 , n19081 , n6283 );
    xnor g10709 ( n6308 , n21616 , n12852 );
    nor g10710 ( n19518 , n17108 , n4008 );
    and g10711 ( n26716 , n12156 , n22242 );
    nor g10712 ( n2434 , n7657 , n25316 );
    not g10713 ( n26875 , n12960 );
    or g10714 ( n9405 , n15315 , n10419 );
    or g10715 ( n6459 , n18216 , n19259 );
    not g10716 ( n349 , n9897 );
    xnor g10717 ( n1674 , n21848 , n7207 );
    not g10718 ( n12929 , n19144 );
    xnor g10719 ( n12108 , n26914 , n8497 );
    nor g10720 ( n12058 , n7486 , n15787 );
    or g10721 ( n10898 , n17333 , n14783 );
    and g10722 ( n23491 , n1672 , n16765 );
    not g10723 ( n141 , n6064 );
    not g10724 ( n22804 , n12663 );
    or g10725 ( n26825 , n19327 , n25624 );
    or g10726 ( n13183 , n8153 , n16333 );
    nor g10727 ( n5494 , n1896 , n8381 );
    or g10728 ( n19776 , n23089 , n12877 );
    xnor g10729 ( n23652 , n20201 , n18496 );
    xnor g10730 ( n4271 , n22182 , n22427 );
    and g10731 ( n26204 , n2323 , n6917 );
    xnor g10732 ( n6965 , n5777 , n18010 );
    or g10733 ( n5926 , n27199 , n20151 );
    or g10734 ( n4072 , n9893 , n22104 );
    or g10735 ( n15318 , n13451 , n949 );
    or g10736 ( n26824 , n25004 , n7375 );
    and g10737 ( n25384 , n17290 , n2034 );
    or g10738 ( n12739 , n15546 , n24922 );
    and g10739 ( n7090 , n1432 , n12040 );
    xnor g10740 ( n7193 , n20259 , n3925 );
    or g10741 ( n18149 , n23477 , n7913 );
    or g10742 ( n7763 , n4277 , n23843 );
    or g10743 ( n8831 , n4486 , n19980 );
    xnor g10744 ( n17288 , n21824 , n11877 );
    or g10745 ( n7475 , n11102 , n20454 );
    and g10746 ( n9197 , n12453 , n2908 );
    or g10747 ( n15823 , n1091 , n15079 );
    xnor g10748 ( n9767 , n6337 , n6128 );
    nor g10749 ( n1443 , n778 , n16291 );
    xnor g10750 ( n4405 , n18421 , n19163 );
    xnor g10751 ( n3122 , n14345 , n14702 );
    or g10752 ( n6725 , n5131 , n11719 );
    or g10753 ( n15648 , n6912 , n25656 );
    not g10754 ( n27156 , n17045 );
    or g10755 ( n20180 , n14431 , n25739 );
    xnor g10756 ( n3037 , n11517 , n20484 );
    or g10757 ( n15844 , n836 , n14696 );
    not g10758 ( n10947 , n2950 );
    or g10759 ( n25591 , n13117 , n18833 );
    not g10760 ( n25050 , n12386 );
    xnor g10761 ( n9713 , n2293 , n6716 );
    xnor g10762 ( n22311 , n15934 , n10864 );
    not g10763 ( n8948 , n5031 );
    and g10764 ( n13517 , n9934 , n20290 );
    nor g10765 ( n22133 , n251 , n8438 );
    xnor g10766 ( n22383 , n4870 , n1350 );
    xnor g10767 ( n23612 , n5824 , n17984 );
    xnor g10768 ( n12072 , n3008 , n22902 );
    xnor g10769 ( n15963 , n22047 , n6352 );
    and g10770 ( n25247 , n98 , n4830 );
    xnor g10771 ( n19775 , n25521 , n11554 );
    xnor g10772 ( n2039 , n2146 , n6785 );
    nor g10773 ( n16669 , n12049 , n10464 );
    nor g10774 ( n14766 , n20639 , n24125 );
    nor g10775 ( n3074 , n24081 , n14255 );
    or g10776 ( n21109 , n4056 , n11555 );
    nor g10777 ( n21476 , n9546 , n14758 );
    nor g10778 ( n13865 , n24358 , n13781 );
    xnor g10779 ( n24736 , n2759 , n8052 );
    and g10780 ( n769 , n8970 , n13536 );
    xnor g10781 ( n26280 , n24465 , n6602 );
    not g10782 ( n24664 , n4183 );
    xnor g10783 ( n4532 , n14032 , n19152 );
    xnor g10784 ( n26703 , n12533 , n24927 );
    or g10785 ( n4456 , n23997 , n15215 );
    and g10786 ( n19993 , n24199 , n14020 );
    and g10787 ( n1024 , n15157 , n8828 );
    not g10788 ( n25041 , n26660 );
    not g10789 ( n18651 , n14576 );
    or g10790 ( n23379 , n11643 , n14590 );
    and g10791 ( n4545 , n3349 , n10501 );
    and g10792 ( n4980 , n13847 , n18206 );
    and g10793 ( n14753 , n20105 , n9589 );
    not g10794 ( n15576 , n8386 );
    or g10795 ( n18112 , n8955 , n5741 );
    and g10796 ( n16265 , n20569 , n3597 );
    and g10797 ( n7622 , n20784 , n2897 );
    not g10798 ( n9068 , n6971 );
    not g10799 ( n12509 , n23789 );
    or g10800 ( n21242 , n8430 , n11701 );
    or g10801 ( n9965 , n22954 , n190 );
    and g10802 ( n934 , n11418 , n14582 );
    and g10803 ( n22593 , n22980 , n13363 );
    not g10804 ( n2997 , n17171 );
    not g10805 ( n481 , n2944 );
    or g10806 ( n4968 , n26146 , n23891 );
    buf g10807 ( n1380 , n1917 );
    and g10808 ( n20619 , n21291 , n14828 );
    and g10809 ( n22151 , n15490 , n328 );
    and g10810 ( n190 , n17011 , n23501 );
    xor g10811 ( n23045 , n14829 , n1165 );
    buf g10812 ( n19390 , n26546 );
    and g10813 ( n10015 , n4507 , n9389 );
    or g10814 ( n14248 , n13535 , n1047 );
    xnor g10815 ( n9040 , n11473 , n15506 );
    xnor g10816 ( n19825 , n21137 , n14130 );
    nor g10817 ( n22673 , n1403 , n5284 );
    xnor g10818 ( n14773 , n24727 , n905 );
    and g10819 ( n19182 , n9634 , n5190 );
    and g10820 ( n22874 , n2972 , n8639 );
    xnor g10821 ( n15881 , n14965 , n10389 );
    xnor g10822 ( n23568 , n15212 , n8174 );
    nor g10823 ( n20407 , n14444 , n5616 );
    xnor g10824 ( n11032 , n9242 , n25240 );
    xnor g10825 ( n12966 , n13137 , n7674 );
    xnor g10826 ( n12567 , n14179 , n19455 );
    nor g10827 ( n12704 , n16683 , n16882 );
    and g10828 ( n16245 , n3392 , n19582 );
    nor g10829 ( n4915 , n9832 , n6513 );
    or g10830 ( n1422 , n16856 , n21081 );
    xnor g10831 ( n4850 , n21597 , n440 );
    not g10832 ( n11278 , n5374 );
    nor g10833 ( n1127 , n5440 , n2724 );
    xnor g10834 ( n10563 , n14603 , n15053 );
    or g10835 ( n12264 , n18994 , n7787 );
    and g10836 ( n15813 , n2740 , n20949 );
    xnor g10837 ( n8824 , n192 , n26884 );
    xnor g10838 ( n17872 , n2267 , n6099 );
    and g10839 ( n20533 , n10218 , n3523 );
    or g10840 ( n4598 , n12126 , n7023 );
    nor g10841 ( n26790 , n4663 , n19390 );
    not g10842 ( n14114 , n4275 );
    or g10843 ( n26074 , n12511 , n19196 );
    nor g10844 ( n11122 , n7524 , n19680 );
    not g10845 ( n22302 , n12015 );
    or g10846 ( n12519 , n5549 , n8302 );
    not g10847 ( n15792 , n23279 );
    and g10848 ( n12664 , n24325 , n10937 );
    xnor g10849 ( n2415 , n12984 , n3468 );
    and g10850 ( n1497 , n16833 , n20592 );
    nor g10851 ( n22732 , n15182 , n12090 );
    xnor g10852 ( n7091 , n10501 , n3349 );
    not g10853 ( n21671 , n16136 );
    not g10854 ( n5479 , n14461 );
    or g10855 ( n7362 , n1118 , n6477 );
    or g10856 ( n17335 , n22770 , n14029 );
    and g10857 ( n3304 , n2351 , n8377 );
    not g10858 ( n11195 , n6501 );
    and g10859 ( n25677 , n8927 , n17574 );
    xnor g10860 ( n870 , n21825 , n16514 );
    not g10861 ( n21634 , n12821 );
    and g10862 ( n975 , n23806 , n17629 );
    and g10863 ( n25042 , n10837 , n1576 );
    xnor g10864 ( n5784 , n26660 , n1163 );
    xnor g10865 ( n4625 , n24982 , n20268 );
    xnor g10866 ( n790 , n4591 , n26562 );
    xnor g10867 ( n6902 , n15447 , n24951 );
    not g10868 ( n8952 , n20707 );
    xnor g10869 ( n8772 , n22946 , n25053 );
    and g10870 ( n6365 , n18030 , n4612 );
    or g10871 ( n25811 , n15178 , n16263 );
    xnor g10872 ( n21789 , n1396 , n15967 );
    and g10873 ( n22033 , n16120 , n19937 );
    or g10874 ( n24401 , n4819 , n210 );
    nor g10875 ( n9094 , n17995 , n462 );
    buf g10876 ( n25156 , n20413 );
    or g10877 ( n10144 , n17083 , n17989 );
    xnor g10878 ( n14202 , n5739 , n16386 );
    not g10879 ( n395 , n4822 );
    and g10880 ( n12677 , n11563 , n24232 );
    and g10881 ( n22084 , n5088 , n26110 );
    not g10882 ( n25171 , n12322 );
    or g10883 ( n10474 , n8580 , n587 );
    or g10884 ( n3774 , n9617 , n10268 );
    nor g10885 ( n22948 , n10470 , n11775 );
    not g10886 ( n19898 , n2858 );
    and g10887 ( n5545 , n25341 , n5173 );
    and g10888 ( n7537 , n643 , n17804 );
    or g10889 ( n10087 , n19950 , n24011 );
    or g10890 ( n21326 , n19794 , n23810 );
    or g10891 ( n23438 , n13117 , n20084 );
    or g10892 ( n2684 , n7759 , n725 );
    and g10893 ( n23156 , n10077 , n9285 );
    xnor g10894 ( n3223 , n17167 , n2546 );
    or g10895 ( n15920 , n23592 , n14440 );
    and g10896 ( n21996 , n11874 , n6994 );
    and g10897 ( n7333 , n16067 , n6937 );
    xnor g10898 ( n1894 , n17139 , n25198 );
    not g10899 ( n18027 , n26119 );
    and g10900 ( n12926 , n24943 , n21027 );
    and g10901 ( n1050 , n16102 , n3922 );
    or g10902 ( n21917 , n616 , n13579 );
    xnor g10903 ( n13270 , n10515 , n16849 );
    not g10904 ( n8792 , n10777 );
    or g10905 ( n25710 , n1953 , n13585 );
    and g10906 ( n22898 , n7901 , n13864 );
    or g10907 ( n26368 , n10619 , n23675 );
    and g10908 ( n1936 , n6675 , n12895 );
    xnor g10909 ( n17948 , n2909 , n9426 );
    not g10910 ( n11657 , n11476 );
    and g10911 ( n11819 , n16664 , n2848 );
    or g10912 ( n2727 , n22275 , n17680 );
    not g10913 ( n12004 , n18 );
    and g10914 ( n21876 , n12650 , n14765 );
    and g10915 ( n720 , n21068 , n11190 );
    not g10916 ( n15389 , n8144 );
    or g10917 ( n11705 , n6803 , n1509 );
    not g10918 ( n26351 , n10560 );
    and g10919 ( n20645 , n7676 , n12512 );
    xnor g10920 ( n21964 , n4022 , n14565 );
    or g10921 ( n18988 , n8572 , n5939 );
    xnor g10922 ( n324 , n14684 , n22588 );
    or g10923 ( n26473 , n16547 , n15 );
    xnor g10924 ( n16744 , n2558 , n14691 );
    and g10925 ( n10584 , n4863 , n23622 );
    not g10926 ( n26293 , n25885 );
    xnor g10927 ( n11426 , n10220 , n15901 );
    and g10928 ( n2883 , n12002 , n27102 );
    or g10929 ( n17182 , n8685 , n21283 );
    xnor g10930 ( n17306 , n9655 , n20946 );
    and g10931 ( n21877 , n26588 , n4573 );
    nor g10932 ( n961 , n24410 , n11662 );
    or g10933 ( n19153 , n744 , n21038 );
    and g10934 ( n23004 , n20049 , n13806 );
    or g10935 ( n17942 , n11676 , n13037 );
    or g10936 ( n23545 , n13411 , n4090 );
    xnor g10937 ( n19894 , n16171 , n5786 );
    xnor g10938 ( n9817 , n17330 , n5414 );
    or g10939 ( n25163 , n337 , n16507 );
    or g10940 ( n17264 , n24263 , n3608 );
    xnor g10941 ( n18721 , n22013 , n17681 );
    or g10942 ( n12759 , n1938 , n25790 );
    or g10943 ( n10673 , n4533 , n6340 );
    xnor g10944 ( n21417 , n5704 , n12315 );
    or g10945 ( n19743 , n1183 , n8582 );
    xnor g10946 ( n3370 , n24620 , n7099 );
    xnor g10947 ( n2961 , n25290 , n10783 );
    or g10948 ( n11927 , n1864 , n17035 );
    xnor g10949 ( n18313 , n2389 , n3007 );
    and g10950 ( n7116 , n2589 , n3087 );
    xnor g10951 ( n12467 , n25186 , n1516 );
    not g10952 ( n11833 , n24182 );
    and g10953 ( n10875 , n12317 , n10394 );
    nor g10954 ( n1734 , n11830 , n18006 );
    not g10955 ( n23487 , n25074 );
    xnor g10956 ( n3968 , n8742 , n21789 );
    nor g10957 ( n26059 , n1405 , n9067 );
    or g10958 ( n20698 , n7915 , n5231 );
    xnor g10959 ( n11415 , n17734 , n10639 );
    not g10960 ( n24778 , n4193 );
    not g10961 ( n24367 , n7221 );
    xnor g10962 ( n8598 , n9332 , n5145 );
    nor g10963 ( n5004 , n13898 , n14275 );
    and g10964 ( n21606 , n7005 , n26820 );
    xor g10965 ( n13518 , n13833 , n1168 );
    or g10966 ( n6577 , n7899 , n22388 );
    not g10967 ( n7973 , n20382 );
    nor g10968 ( n22760 , n11542 , n15079 );
    xnor g10969 ( n13500 , n9819 , n14960 );
    and g10970 ( n4457 , n3520 , n19235 );
    xnor g10971 ( n14765 , n5234 , n12702 );
    xnor g10972 ( n21182 , n25428 , n16522 );
    and g10973 ( n9705 , n20478 , n26030 );
    xnor g10974 ( n16983 , n25316 , n20385 );
    xnor g10975 ( n18792 , n7591 , n23680 );
    or g10976 ( n4252 , n8958 , n21014 );
    not g10977 ( n5852 , n1138 );
    or g10978 ( n13883 , n23526 , n25081 );
    or g10979 ( n26003 , n4446 , n4734 );
    or g10980 ( n19345 , n15317 , n21568 );
    xnor g10981 ( n25619 , n5281 , n13176 );
    and g10982 ( n16411 , n25287 , n23538 );
    not g10983 ( n15426 , n26913 );
    nor g10984 ( n26465 , n5402 , n7361 );
    not g10985 ( n19869 , n1913 );
    not g10986 ( n1182 , n3506 );
    and g10987 ( n8702 , n16153 , n25116 );
    xnor g10988 ( n21549 , n8506 , n11584 );
    xnor g10989 ( n17263 , n3569 , n21013 );
    not g10990 ( n22108 , n8583 );
    not g10991 ( n21871 , n25494 );
    not g10992 ( n9631 , n2331 );
    not g10993 ( n4970 , n21082 );
    or g10994 ( n16435 , n25255 , n17321 );
    and g10995 ( n374 , n15823 , n15606 );
    or g10996 ( n27204 , n21716 , n4457 );
    xnor g10997 ( n16948 , n15484 , n24964 );
    and g10998 ( n17145 , n18740 , n20283 );
    or g10999 ( n11368 , n22510 , n14306 );
    or g11000 ( n4535 , n19718 , n16956 );
    xnor g11001 ( n16232 , n1653 , n8913 );
    or g11002 ( n27050 , n6029 , n758 );
    xnor g11003 ( n4548 , n12944 , n2439 );
    and g11004 ( n22882 , n7809 , n15038 );
    or g11005 ( n8727 , n2416 , n16455 );
    xnor g11006 ( n14414 , n14213 , n18252 );
    or g11007 ( n5632 , n7040 , n12799 );
    xnor g11008 ( n24177 , n20851 , n5385 );
    not g11009 ( n20117 , n196 );
    not g11010 ( n19113 , n26879 );
    not g11011 ( n24152 , n9358 );
    or g11012 ( n7889 , n24136 , n18806 );
    xnor g11013 ( n24847 , n27126 , n26068 );
    not g11014 ( n25228 , n9192 );
    or g11015 ( n24811 , n8077 , n10843 );
    nor g11016 ( n24810 , n4626 , n21509 );
    or g11017 ( n11601 , n27122 , n17251 );
    not g11018 ( n6895 , n13858 );
    and g11019 ( n6158 , n5735 , n9132 );
    or g11020 ( n26166 , n9196 , n12354 );
    or g11021 ( n20911 , n14823 , n12753 );
    not g11022 ( n26367 , n14878 );
    and g11023 ( n5897 , n12951 , n9704 );
    not g11024 ( n13420 , n5673 );
    nor g11025 ( n12534 , n10023 , n6670 );
    and g11026 ( n23985 , n19293 , n659 );
    and g11027 ( n9843 , n4236 , n8239 );
    or g11028 ( n10142 , n4711 , n715 );
    xnor g11029 ( n20092 , n4032 , n17898 );
    xnor g11030 ( n12531 , n15308 , n3202 );
    or g11031 ( n18811 , n16420 , n2233 );
    and g11032 ( n6389 , n17655 , n10144 );
    nor g11033 ( n8813 , n4469 , n23545 );
    or g11034 ( n11795 , n5578 , n1493 );
    or g11035 ( n10237 , n9291 , n1413 );
    xnor g11036 ( n13947 , n26942 , n9498 );
    not g11037 ( n24237 , n25250 );
    and g11038 ( n7914 , n3739 , n15892 );
    not g11039 ( n24468 , n17792 );
    and g11040 ( n12382 , n13105 , n1551 );
    not g11041 ( n3549 , n10422 );
    xnor g11042 ( n235 , n5845 , n9566 );
    and g11043 ( n1965 , n24330 , n5320 );
    not g11044 ( n2218 , n16314 );
    not g11045 ( n17431 , n10706 );
    xnor g11046 ( n10267 , n5322 , n21488 );
    xnor g11047 ( n16314 , n6455 , n25467 );
    and g11048 ( n1846 , n20385 , n23932 );
    or g11049 ( n2278 , n14557 , n16982 );
    xnor g11050 ( n19399 , n5307 , n22646 );
    buf g11051 ( n14528 , n12367 );
    nor g11052 ( n4547 , n2732 , n21085 );
    or g11053 ( n5888 , n26168 , n19660 );
    or g11054 ( n2466 , n14309 , n9611 );
    or g11055 ( n23125 , n6729 , n1106 );
    or g11056 ( n1355 , n20945 , n22953 );
    and g11057 ( n3881 , n12856 , n24703 );
    nor g11058 ( n22209 , n19313 , n20444 );
    xnor g11059 ( n5549 , n23622 , n20199 );
    xnor g11060 ( n7919 , n1493 , n12585 );
    nor g11061 ( n3266 , n7593 , n17415 );
    xnor g11062 ( n9413 , n12805 , n12350 );
    xnor g11063 ( n23610 , n8491 , n25586 );
    and g11064 ( n13580 , n24442 , n4541 );
    xnor g11065 ( n25061 , n16276 , n24374 );
    nor g11066 ( n8999 , n4665 , n7823 );
    or g11067 ( n26033 , n20277 , n17460 );
    nor g11068 ( n21873 , n22597 , n18901 );
    not g11069 ( n9717 , n24842 );
    xnor g11070 ( n1863 , n1040 , n12152 );
    xnor g11071 ( n21590 , n13291 , n2443 );
    and g11072 ( n13689 , n8838 , n1987 );
    and g11073 ( n15585 , n2915 , n10625 );
    nor g11074 ( n5388 , n12078 , n3354 );
    xnor g11075 ( n24256 , n19058 , n9445 );
    or g11076 ( n11820 , n26574 , n5664 );
    or g11077 ( n13977 , n6400 , n18554 );
    xnor g11078 ( n7722 , n5358 , n20726 );
    xnor g11079 ( n2650 , n20051 , n4901 );
    and g11080 ( n6074 , n19934 , n24224 );
    or g11081 ( n26956 , n23705 , n21287 );
    and g11082 ( n14951 , n2254 , n13458 );
    or g11083 ( n18021 , n24716 , n20875 );
    xnor g11084 ( n14451 , n2566 , n23677 );
    and g11085 ( n5254 , n1459 , n8193 );
    and g11086 ( n26080 , n8230 , n20653 );
    xnor g11087 ( n23207 , n18834 , n14231 );
    nor g11088 ( n1559 , n26957 , n14130 );
    and g11089 ( n26217 , n2886 , n16609 );
    not g11090 ( n13529 , n27175 );
    xnor g11091 ( n13557 , n26951 , n22477 );
    xnor g11092 ( n17636 , n3116 , n24980 );
    or g11093 ( n11673 , n8255 , n5 );
    or g11094 ( n24797 , n8539 , n14610 );
    xnor g11095 ( n21630 , n13968 , n18649 );
    or g11096 ( n14434 , n4780 , n15258 );
    or g11097 ( n17890 , n16528 , n4503 );
    xnor g11098 ( n17320 , n25755 , n7358 );
    or g11099 ( n19306 , n14156 , n11552 );
    xnor g11100 ( n18075 , n24323 , n1681 );
    not g11101 ( n10148 , n8508 );
    nor g11102 ( n601 , n19464 , n5108 );
    xnor g11103 ( n13885 , n26000 , n2394 );
    xnor g11104 ( n10713 , n12076 , n8856 );
    and g11105 ( n4908 , n24564 , n15962 );
    nor g11106 ( n12988 , n21520 , n19615 );
    and g11107 ( n15957 , n20964 , n6762 );
    xnor g11108 ( n4649 , n9402 , n6864 );
    xnor g11109 ( n8973 , n20213 , n26725 );
    nor g11110 ( n20589 , n19914 , n24551 );
    or g11111 ( n23482 , n18546 , n25834 );
    xnor g11112 ( n1501 , n17616 , n959 );
    xnor g11113 ( n21827 , n1339 , n21842 );
    xnor g11114 ( n18400 , n12962 , n26662 );
    or g11115 ( n988 , n146 , n16889 );
    xnor g11116 ( n24606 , n22810 , n22120 );
    and g11117 ( n11723 , n7288 , n19064 );
    not g11118 ( n20137 , n7437 );
    or g11119 ( n7488 , n24574 , n16228 );
    not g11120 ( n22061 , n18425 );
    nor g11121 ( n17292 , n15087 , n3257 );
    xnor g11122 ( n15145 , n25894 , n8205 );
    and g11123 ( n2379 , n20586 , n7299 );
    or g11124 ( n7255 , n1418 , n2878 );
    xnor g11125 ( n5256 , n12270 , n15963 );
    and g11126 ( n15253 , n26710 , n15418 );
    and g11127 ( n12912 , n20463 , n13687 );
    xnor g11128 ( n3552 , n291 , n5117 );
    and g11129 ( n6817 , n12221 , n19049 );
    and g11130 ( n15888 , n25004 , n7375 );
    and g11131 ( n19465 , n26312 , n26993 );
    and g11132 ( n19324 , n15027 , n8030 );
    and g11133 ( n2020 , n22161 , n19931 );
    xnor g11134 ( n23473 , n16313 , n15164 );
    or g11135 ( n9121 , n13737 , n16907 );
    not g11136 ( n26433 , n11670 );
    xnor g11137 ( n12070 , n25729 , n3279 );
    or g11138 ( n11641 , n2317 , n5109 );
    and g11139 ( n20916 , n5535 , n23137 );
    nor g11140 ( n21847 , n11566 , n12198 );
    nor g11141 ( n4522 , n6692 , n15661 );
    nor g11142 ( n4799 , n24736 , n8713 );
    or g11143 ( n12156 , n10037 , n19196 );
    or g11144 ( n23105 , n16232 , n22294 );
    or g11145 ( n21887 , n16830 , n18295 );
    xnor g11146 ( n26028 , n19820 , n1057 );
    and g11147 ( n1107 , n7421 , n20044 );
    and g11148 ( n4602 , n12318 , n25955 );
    and g11149 ( n20664 , n2543 , n19810 );
    not g11150 ( n14118 , n16260 );
    and g11151 ( n16641 , n13357 , n11077 );
    and g11152 ( n4906 , n8854 , n19145 );
    nor g11153 ( n16246 , n1553 , n3547 );
    or g11154 ( n24398 , n4615 , n26233 );
    nor g11155 ( n5229 , n1839 , n5886 );
    not g11156 ( n2857 , n9110 );
    or g11157 ( n9715 , n12356 , n1545 );
    and g11158 ( n4097 , n504 , n26135 );
    not g11159 ( n212 , n6785 );
    xnor g11160 ( n22509 , n20470 , n3366 );
    xnor g11161 ( n17279 , n5260 , n16130 );
    or g11162 ( n20078 , n17002 , n7731 );
    xnor g11163 ( n7276 , n12163 , n10139 );
    not g11164 ( n4236 , n14258 );
    nor g11165 ( n9433 , n11580 , n19230 );
    and g11166 ( n24867 , n9143 , n16697 );
    xnor g11167 ( n2954 , n13288 , n18874 );
    nor g11168 ( n20379 , n8722 , n10791 );
    xnor g11169 ( n6726 , n19824 , n22406 );
    xnor g11170 ( n25346 , n17926 , n17598 );
    xnor g11171 ( n21089 , n22742 , n26903 );
    not g11172 ( n25939 , n5231 );
    or g11173 ( n19676 , n13842 , n13708 );
    and g11174 ( n3360 , n8610 , n4689 );
    and g11175 ( n14894 , n5540 , n14179 );
    xnor g11176 ( n23636 , n802 , n21629 );
    xnor g11177 ( n10506 , n9576 , n21599 );
    nor g11178 ( n17708 , n26222 , n12565 );
    xnor g11179 ( n24242 , n21907 , n26054 );
    not g11180 ( n19134 , n6915 );
    or g11181 ( n22337 , n6996 , n8570 );
    and g11182 ( n10366 , n25054 , n10138 );
    xnor g11183 ( n11298 , n13081 , n18729 );
    and g11184 ( n2157 , n8086 , n26948 );
    xnor g11185 ( n24739 , n22203 , n20259 );
    xnor g11186 ( n18974 , n6118 , n1521 );
    or g11187 ( n4417 , n3061 , n2808 );
    xnor g11188 ( n17912 , n6353 , n12242 );
    or g11189 ( n22512 , n17794 , n22551 );
    or g11190 ( n20899 , n6010 , n22989 );
    and g11191 ( n10418 , n4679 , n19102 );
    or g11192 ( n2497 , n23467 , n10772 );
    xnor g11193 ( n7436 , n13458 , n25793 );
    xnor g11194 ( n5050 , n10308 , n7163 );
    or g11195 ( n22860 , n24170 , n24085 );
    and g11196 ( n22352 , n3005 , n9348 );
    nor g11197 ( n20660 , n20088 , n5086 );
    xnor g11198 ( n25460 , n14744 , n691 );
    xnor g11199 ( n3150 , n316 , n24210 );
    and g11200 ( n11378 , n17568 , n3171 );
    nor g11201 ( n27140 , n11714 , n10861 );
    xnor g11202 ( n19741 , n2215 , n8706 );
    or g11203 ( n5035 , n736 , n9148 );
    not g11204 ( n16532 , n4787 );
    or g11205 ( n4730 , n4132 , n2005 );
    not g11206 ( n7359 , n12610 );
    and g11207 ( n16263 , n5879 , n20806 );
    xnor g11208 ( n1893 , n7846 , n9609 );
    or g11209 ( n15538 , n400 , n19478 );
    xnor g11210 ( n22618 , n7619 , n11044 );
    or g11211 ( n25197 , n26766 , n21664 );
    and g11212 ( n22648 , n15102 , n8237 );
    nor g11213 ( n1793 , n26882 , n106 );
    or g11214 ( n20346 , n24972 , n5429 );
    or g11215 ( n5396 , n11205 , n19975 );
    and g11216 ( n21886 , n379 , n20671 );
    not g11217 ( n22408 , n1441 );
    and g11218 ( n9842 , n1290 , n22657 );
    or g11219 ( n3905 , n22116 , n15605 );
    or g11220 ( n8926 , n21969 , n19284 );
    not g11221 ( n18363 , n15392 );
    xnor g11222 ( n4947 , n19096 , n19063 );
    or g11223 ( n17046 , n18643 , n14314 );
    nor g11224 ( n24827 , n21037 , n13899 );
    or g11225 ( n23206 , n21961 , n16121 );
    and g11226 ( n10890 , n21947 , n16525 );
    not g11227 ( n8266 , n690 );
    xnor g11228 ( n20512 , n27184 , n4812 );
    nor g11229 ( n7642 , n11457 , n6385 );
    or g11230 ( n15641 , n7921 , n1065 );
    or g11231 ( n41 , n2773 , n12927 );
    and g11232 ( n12713 , n19672 , n19987 );
    and g11233 ( n15605 , n1189 , n15195 );
    or g11234 ( n603 , n9598 , n7759 );
    xnor g11235 ( n6501 , n21656 , n20519 );
    not g11236 ( n5774 , n6229 );
    not g11237 ( n23708 , n15960 );
    xnor g11238 ( n1081 , n10224 , n11481 );
    not g11239 ( n2721 , n13549 );
    or g11240 ( n20524 , n13577 , n23587 );
    not g11241 ( n17301 , n8957 );
    or g11242 ( n4377 , n21229 , n7036 );
    xnor g11243 ( n17758 , n5704 , n22309 );
    or g11244 ( n47 , n21359 , n23384 );
    xnor g11245 ( n13506 , n24803 , n227 );
    and g11246 ( n1756 , n8804 , n12729 );
    and g11247 ( n2924 , n5705 , n3227 );
    nor g11248 ( n15409 , n27104 , n19005 );
    or g11249 ( n8481 , n23072 , n26384 );
    not g11250 ( n25941 , n15586 );
    not g11251 ( n10255 , n17142 );
    xnor g11252 ( n4106 , n13372 , n1681 );
    xnor g11253 ( n3340 , n23172 , n20578 );
    or g11254 ( n10594 , n17022 , n150 );
    xnor g11255 ( n5687 , n24550 , n4791 );
    or g11256 ( n21121 , n9102 , n19180 );
    xnor g11257 ( n18943 , n9204 , n7359 );
    or g11258 ( n2581 , n1868 , n26791 );
    not g11259 ( n15221 , n9003 );
    xnor g11260 ( n4554 , n5304 , n20516 );
    xnor g11261 ( n12740 , n4292 , n14454 );
    and g11262 ( n14101 , n20753 , n14581 );
    xnor g11263 ( n8366 , n14255 , n5882 );
    xnor g11264 ( n3477 , n22382 , n23326 );
    or g11265 ( n11001 , n10075 , n8225 );
    xnor g11266 ( n14749 , n10286 , n25044 );
    and g11267 ( n17221 , n1595 , n12820 );
    and g11268 ( n25903 , n15809 , n181 );
    and g11269 ( n26268 , n12044 , n11231 );
    xnor g11270 ( n18428 , n25806 , n9445 );
    or g11271 ( n25348 , n2436 , n11714 );
    or g11272 ( n5588 , n4415 , n23859 );
    not g11273 ( n14992 , n2416 );
    and g11274 ( n12257 , n20501 , n14476 );
    and g11275 ( n5664 , n21059 , n10921 );
    nor g11276 ( n7756 , n12343 , n25568 );
    and g11277 ( n13441 , n4413 , n23116 );
    xnor g11278 ( n16595 , n10760 , n10882 );
    xnor g11279 ( n2699 , n7497 , n22863 );
    not g11280 ( n15000 , n12674 );
    and g11281 ( n16336 , n15404 , n10610 );
    or g11282 ( n20368 , n25716 , n25708 );
    or g11283 ( n22453 , n23617 , n21493 );
    xnor g11284 ( n25097 , n25911 , n1724 );
    xnor g11285 ( n3851 , n2510 , n7678 );
    and g11286 ( n5537 , n17841 , n19096 );
    and g11287 ( n19075 , n503 , n25056 );
    not g11288 ( n22501 , n25855 );
    xnor g11289 ( n20673 , n3734 , n25984 );
    not g11290 ( n1105 , n1834 );
    or g11291 ( n10180 , n15918 , n21021 );
    xnor g11292 ( n5868 , n5993 , n1185 );
    or g11293 ( n1468 , n784 , n21692 );
    not g11294 ( n24101 , n2551 );
    nor g11295 ( n18236 , n6753 , n2453 );
    nor g11296 ( n13513 , n21247 , n1631 );
    nor g11297 ( n1669 , n6831 , n7546 );
    xnor g11298 ( n11567 , n6502 , n1630 );
    xnor g11299 ( n18895 , n14735 , n16812 );
    and g11300 ( n22798 , n11796 , n21464 );
    and g11301 ( n17699 , n16789 , n10962 );
    xnor g11302 ( n3987 , n23974 , n8309 );
    xnor g11303 ( n19670 , n1630 , n11121 );
    and g11304 ( n12694 , n20990 , n13344 );
    or g11305 ( n7262 , n13488 , n6520 );
    nor g11306 ( n18352 , n7170 , n19186 );
    nor g11307 ( n3100 , n10146 , n329 );
    and g11308 ( n12993 , n3643 , n24883 );
    or g11309 ( n14037 , n8801 , n5889 );
    not g11310 ( n8239 , n22846 );
    xnor g11311 ( n20879 , n13509 , n4861 );
    nor g11312 ( n6275 , n3832 , n20006 );
    not g11313 ( n24802 , n8170 );
    and g11314 ( n13315 , n5576 , n1763 );
    and g11315 ( n22388 , n25472 , n1966 );
    or g11316 ( n2840 , n20112 , n2161 );
    nor g11317 ( n15658 , n7297 , n304 );
    and g11318 ( n15446 , n24480 , n14634 );
    or g11319 ( n24794 , n14440 , n7523 );
    xnor g11320 ( n19562 , n13677 , n26752 );
    xnor g11321 ( n2444 , n4336 , n24967 );
    or g11322 ( n20373 , n8117 , n3280 );
    xnor g11323 ( n26313 , n15659 , n5213 );
    xnor g11324 ( n24681 , n4685 , n21213 );
    xnor g11325 ( n20707 , n7562 , n5584 );
    or g11326 ( n14212 , n23322 , n12185 );
    and g11327 ( n9738 , n18511 , n14361 );
    xor g11328 ( n513 , n14192 , n3320 );
    not g11329 ( n25521 , n24188 );
    not g11330 ( n13748 , n5288 );
    or g11331 ( n5655 , n5207 , n21284 );
    xnor g11332 ( n956 , n11623 , n19938 );
    xnor g11333 ( n20111 , n5400 , n9512 );
    xnor g11334 ( n17132 , n6755 , n13988 );
    xnor g11335 ( n8379 , n683 , n21299 );
    and g11336 ( n20428 , n18053 , n2844 );
    or g11337 ( n8590 , n11964 , n12345 );
    and g11338 ( n22275 , n1099 , n3379 );
    or g11339 ( n10213 , n11947 , n23271 );
    or g11340 ( n8536 , n25439 , n14782 );
    or g11341 ( n3303 , n944 , n22738 );
    xnor g11342 ( n17940 , n21878 , n17743 );
    or g11343 ( n2595 , n9638 , n18631 );
    or g11344 ( n2772 , n11170 , n8260 );
    xnor g11345 ( n20355 , n11784 , n70 );
    xnor g11346 ( n5168 , n8392 , n27153 );
    xnor g11347 ( n348 , n16704 , n5981 );
    xnor g11348 ( n18243 , n19153 , n27044 );
    not g11349 ( n5429 , n11611 );
    nor g11350 ( n8759 , n17056 , n23545 );
    xnor g11351 ( n6928 , n23464 , n9877 );
    or g11352 ( n7989 , n9206 , n6597 );
    xnor g11353 ( n17412 , n15471 , n17712 );
    or g11354 ( n26687 , n18950 , n17846 );
    or g11355 ( n23850 , n24054 , n14032 );
    xnor g11356 ( n26954 , n25068 , n8324 );
    or g11357 ( n23263 , n25340 , n15744 );
    not g11358 ( n23863 , n14345 );
    nor g11359 ( n10488 , n8472 , n6150 );
    or g11360 ( n10380 , n19297 , n23754 );
    or g11361 ( n21541 , n9294 , n18880 );
    or g11362 ( n12499 , n19546 , n5130 );
    xnor g11363 ( n20795 , n14016 , n21106 );
    or g11364 ( n15021 , n24325 , n21353 );
    xnor g11365 ( n13558 , n22205 , n26288 );
    xnor g11366 ( n24967 , n23161 , n22237 );
    xnor g11367 ( n16823 , n9928 , n6785 );
    and g11368 ( n16403 , n20931 , n6144 );
    and g11369 ( n16570 , n1873 , n10814 );
    and g11370 ( n24901 , n17164 , n18726 );
    not g11371 ( n14138 , n1599 );
    xnor g11372 ( n24378 , n22567 , n4532 );
    xnor g11373 ( n23911 , n2944 , n13951 );
    xor g11374 ( n21498 , n13108 , n5026 );
    and g11375 ( n6643 , n16335 , n23893 );
    not g11376 ( n11502 , n502 );
    xnor g11377 ( n274 , n14208 , n2547 );
    xnor g11378 ( n11918 , n13313 , n18959 );
    and g11379 ( n17162 , n24025 , n20951 );
    xnor g11380 ( n24210 , n7436 , n5098 );
    or g11381 ( n11007 , n17066 , n22773 );
    not g11382 ( n24960 , n8551 );
    xnor g11383 ( n11431 , n19594 , n6235 );
    or g11384 ( n9677 , n7361 , n14885 );
    xnor g11385 ( n2054 , n16393 , n11653 );
    xnor g11386 ( n1129 , n19227 , n19005 );
    and g11387 ( n11324 , n25957 , n19247 );
    not g11388 ( n1176 , n3136 );
    xnor g11389 ( n26290 , n19797 , n24620 );
    nor g11390 ( n2486 , n10660 , n8897 );
    xnor g11391 ( n9191 , n5725 , n1499 );
    or g11392 ( n6552 , n225 , n26181 );
    and g11393 ( n21470 , n14851 , n3036 );
    xnor g11394 ( n2817 , n20700 , n12875 );
    or g11395 ( n4994 , n7569 , n1779 );
    xnor g11396 ( n9981 , n21841 , n12693 );
    and g11397 ( n406 , n20155 , n24424 );
    or g11398 ( n12247 , n2230 , n18295 );
    nor g11399 ( n4986 , n9133 , n393 );
    and g11400 ( n9997 , n23561 , n10364 );
    and g11401 ( n20848 , n11778 , n21121 );
    xnor g11402 ( n19414 , n13181 , n16447 );
    nor g11403 ( n24595 , n13419 , n23475 );
    and g11404 ( n14567 , n23614 , n17611 );
    xnor g11405 ( n25858 , n4119 , n1525 );
    and g11406 ( n8905 , n21061 , n22956 );
    or g11407 ( n12200 , n7487 , n16571 );
    xnor g11408 ( n25215 , n12368 , n2881 );
    xnor g11409 ( n20176 , n23642 , n24309 );
    xnor g11410 ( n24365 , n15884 , n5213 );
    xnor g11411 ( n5733 , n19643 , n9694 );
    or g11412 ( n21819 , n10013 , n25971 );
    or g11413 ( n2381 , n9119 , n9929 );
    nor g11414 ( n12327 , n21334 , n18399 );
    xnor g11415 ( n2794 , n25394 , n8964 );
    nor g11416 ( n13713 , n21489 , n11151 );
    xnor g11417 ( n2993 , n2731 , n4812 );
    xnor g11418 ( n11174 , n15090 , n20608 );
    and g11419 ( n11638 , n20336 , n23233 );
    and g11420 ( n1466 , n3782 , n8474 );
    or g11421 ( n7649 , n22670 , n21050 );
    and g11422 ( n7548 , n20948 , n5946 );
    and g11423 ( n6849 , n5663 , n4945 );
    not g11424 ( n3862 , n3554 );
    and g11425 ( n6380 , n13275 , n14427 );
    xnor g11426 ( n22683 , n18351 , n9024 );
    nor g11427 ( n20062 , n9600 , n3791 );
    nor g11428 ( n22223 , n22009 , n24839 );
    xnor g11429 ( n1784 , n15284 , n8772 );
    xnor g11430 ( n17927 , n24303 , n1027 );
    not g11431 ( n26086 , n16971 );
    or g11432 ( n24667 , n19763 , n4922 );
    not g11433 ( n21520 , n19955 );
    xnor g11434 ( n17663 , n23149 , n7240 );
    nor g11435 ( n15890 , n20415 , n14852 );
    or g11436 ( n5287 , n18098 , n13530 );
    xnor g11437 ( n19184 , n16671 , n20690 );
    nor g11438 ( n16600 , n23063 , n19494 );
    not g11439 ( n21565 , n75 );
    and g11440 ( n2947 , n26621 , n5136 );
    xnor g11441 ( n22414 , n5468 , n16801 );
    and g11442 ( n14058 , n26246 , n20778 );
    or g11443 ( n12233 , n9675 , n11723 );
    xnor g11444 ( n11497 , n24027 , n24956 );
    and g11445 ( n2259 , n16162 , n693 );
    xnor g11446 ( n15574 , n10625 , n19454 );
    and g11447 ( n20697 , n9232 , n11042 );
    nor g11448 ( n6134 , n11740 , n19941 );
    not g11449 ( n10501 , n9550 );
    and g11450 ( n4397 , n1398 , n20548 );
    xnor g11451 ( n1332 , n26570 , n15105 );
    xnor g11452 ( n10479 , n12139 , n17891 );
    not g11453 ( n15147 , n14163 );
    or g11454 ( n229 , n3525 , n17935 );
    xnor g11455 ( n25826 , n9414 , n538 );
    nor g11456 ( n18420 , n14336 , n20077 );
    or g11457 ( n26685 , n17494 , n15450 );
    not g11458 ( n26957 , n14440 );
    or g11459 ( n6840 , n5846 , n21950 );
    or g11460 ( n4212 , n16003 , n489 );
    or g11461 ( n13396 , n13643 , n6466 );
    xnor g11462 ( n24927 , n10158 , n1136 );
    not g11463 ( n13485 , n3716 );
    xnor g11464 ( n7100 , n25034 , n7975 );
    not g11465 ( n530 , n21267 );
    not g11466 ( n23208 , n24736 );
    nor g11467 ( n22224 , n6355 , n8589 );
    and g11468 ( n3361 , n19621 , n27204 );
    or g11469 ( n20459 , n11655 , n4644 );
    nor g11470 ( n17208 , n8492 , n25739 );
    or g11471 ( n17946 , n20562 , n13109 );
    xnor g11472 ( n20840 , n4406 , n8810 );
    xnor g11473 ( n7598 , n14712 , n10714 );
    or g11474 ( n20888 , n6641 , n17952 );
    or g11475 ( n21303 , n20645 , n21475 );
    or g11476 ( n5492 , n12129 , n26173 );
    xnor g11477 ( n18874 , n13158 , n8309 );
    not g11478 ( n15038 , n25100 );
    xnor g11479 ( n4685 , n26004 , n26896 );
    xnor g11480 ( n10520 , n22671 , n17975 );
    nor g11481 ( n191 , n14637 , n11210 );
    xnor g11482 ( n22002 , n24677 , n10866 );
    and g11483 ( n15772 , n9642 , n6331 );
    xnor g11484 ( n10709 , n13140 , n4158 );
    xnor g11485 ( n16828 , n16455 , n2416 );
    or g11486 ( n1494 , n12096 , n9488 );
    xnor g11487 ( n23964 , n22671 , n22017 );
    xnor g11488 ( n14970 , n6141 , n5028 );
    or g11489 ( n21099 , n12435 , n16281 );
    and g11490 ( n26089 , n15188 , n24725 );
    xnor g11491 ( n14679 , n16662 , n7769 );
    xnor g11492 ( n13578 , n15451 , n1949 );
    nor g11493 ( n14551 , n5342 , n17559 );
    or g11494 ( n16343 , n18266 , n11814 );
    not g11495 ( n25533 , n5110 );
    not g11496 ( n21104 , n5017 );
    xnor g11497 ( n23876 , n11197 , n25878 );
    or g11498 ( n6217 , n14406 , n19643 );
    xnor g11499 ( n12742 , n2830 , n22394 );
    or g11500 ( n9590 , n11286 , n7392 );
    xnor g11501 ( n14577 , n11486 , n20235 );
    or g11502 ( n5962 , n20059 , n17671 );
    xnor g11503 ( n21175 , n17868 , n4141 );
    and g11504 ( n11204 , n17745 , n15843 );
    not g11505 ( n14127 , n15914 );
    xnor g11506 ( n24536 , n26338 , n18166 );
    and g11507 ( n3917 , n25149 , n12948 );
    or g11508 ( n13238 , n25099 , n20455 );
    xnor g11509 ( n12406 , n12691 , n25080 );
    nor g11510 ( n7419 , n19869 , n676 );
    nor g11511 ( n5364 , n905 , n24727 );
    xnor g11512 ( n15663 , n21 , n20923 );
    not g11513 ( n5266 , n24745 );
    or g11514 ( n6676 , n15311 , n7574 );
    and g11515 ( n22490 , n17214 , n15907 );
    or g11516 ( n3821 , n22764 , n2360 );
    xnor g11517 ( n21205 , n10070 , n26483 );
    or g11518 ( n3137 , n17035 , n2680 );
    and g11519 ( n9747 , n12955 , n7353 );
    not g11520 ( n10681 , n25001 );
    xnor g11521 ( n7001 , n14873 , n9452 );
    not g11522 ( n20051 , n24117 );
    and g11523 ( n18412 , n11459 , n18781 );
    xnor g11524 ( n1170 , n20427 , n24860 );
    xnor g11525 ( n17504 , n2360 , n17458 );
    or g11526 ( n16177 , n24765 , n23447 );
    or g11527 ( n15855 , n23806 , n17629 );
    or g11528 ( n10963 , n1978 , n17055 );
    nor g11529 ( n15293 , n18506 , n19514 );
    not g11530 ( n9015 , n16981 );
    nor g11531 ( n2856 , n19514 , n2415 );
    xnor g11532 ( n25359 , n14122 , n22300 );
    or g11533 ( n1520 , n1110 , n9553 );
    xnor g11534 ( n4712 , n6033 , n21658 );
    not g11535 ( n20131 , n26557 );
    nor g11536 ( n605 , n13301 , n23313 );
    or g11537 ( n4287 , n14790 , n342 );
    and g11538 ( n4324 , n20212 , n6472 );
    not g11539 ( n27147 , n24194 );
    or g11540 ( n7075 , n12303 , n2406 );
    and g11541 ( n1903 , n17595 , n14134 );
    and g11542 ( n18494 , n18848 , n20038 );
    and g11543 ( n17216 , n5312 , n7800 );
    and g11544 ( n15483 , n6040 , n26812 );
    not g11545 ( n21321 , n4008 );
    not g11546 ( n12802 , n15009 );
    xnor g11547 ( n23935 , n19436 , n9792 );
    xnor g11548 ( n16574 , n13053 , n24150 );
    xnor g11549 ( n17684 , n13949 , n5128 );
    and g11550 ( n24918 , n13434 , n390 );
    xnor g11551 ( n18166 , n26510 , n22332 );
    not g11552 ( n17532 , n11667 );
    xnor g11553 ( n26713 , n15125 , n9130 );
    or g11554 ( n7895 , n23877 , n25918 );
    or g11555 ( n11541 , n11788 , n5301 );
    not g11556 ( n26227 , n4199 );
    xnor g11557 ( n4601 , n1452 , n14236 );
    not g11558 ( n9053 , n3740 );
    and g11559 ( n4373 , n14948 , n6973 );
    or g11560 ( n5606 , n13188 , n5738 );
    or g11561 ( n24071 , n20964 , n20946 );
    and g11562 ( n2243 , n7228 , n2991 );
    xnor g11563 ( n11304 , n6168 , n7555 );
    or g11564 ( n3824 , n18990 , n673 );
    or g11565 ( n11735 , n21307 , n25103 );
    nor g11566 ( n12636 , n9204 , n12251 );
    not g11567 ( n18606 , n669 );
    not g11568 ( n2656 , n1708 );
    nor g11569 ( n2269 , n8647 , n24343 );
    and g11570 ( n23187 , n16889 , n8278 );
    or g11571 ( n12951 , n20737 , n919 );
    nor g11572 ( n18773 , n15433 , n15539 );
    or g11573 ( n3110 , n18318 , n20171 );
    and g11574 ( n4914 , n3095 , n22199 );
    xnor g11575 ( n23939 , n11782 , n5591 );
    xnor g11576 ( n21857 , n12685 , n11274 );
    xnor g11577 ( n1253 , n15271 , n5822 );
    nor g11578 ( n19332 , n8732 , n15914 );
    or g11579 ( n6534 , n7952 , n3952 );
    xnor g11580 ( n19217 , n16765 , n26999 );
    and g11581 ( n17893 , n12215 , n4979 );
    and g11582 ( n24800 , n5104 , n3997 );
    and g11583 ( n16639 , n24676 , n19407 );
    xnor g11584 ( n25712 , n24026 , n5780 );
    or g11585 ( n23733 , n4876 , n11819 );
    or g11586 ( n4521 , n2428 , n4280 );
    or g11587 ( n21646 , n17862 , n6063 );
    xnor g11588 ( n17518 , n17390 , n21247 );
    or g11589 ( n24670 , n17993 , n23145 );
    or g11590 ( n20540 , n24007 , n22028 );
    xnor g11591 ( n332 , n9953 , n9487 );
    xnor g11592 ( n23257 , n24745 , n3724 );
    nor g11593 ( n11413 , n821 , n8856 );
    xnor g11594 ( n129 , n8856 , n22442 );
    or g11595 ( n13437 , n4236 , n21476 );
    not g11596 ( n12381 , n7946 );
    and g11597 ( n11406 , n25910 , n13009 );
    xnor g11598 ( n9940 , n21962 , n13074 );
    xnor g11599 ( n25944 , n3337 , n709 );
    and g11600 ( n12071 , n14736 , n3529 );
    or g11601 ( n12635 , n9663 , n1526 );
    nor g11602 ( n15717 , n3284 , n8003 );
    nor g11603 ( n16680 , n20032 , n7149 );
    xnor g11604 ( n11262 , n26425 , n2151 );
    nor g11605 ( n10816 , n9909 , n1694 );
    nor g11606 ( n12642 , n5131 , n19674 );
    nor g11607 ( n23718 , n12875 , n12652 );
    xnor g11608 ( n23643 , n16971 , n19144 );
    xnor g11609 ( n21302 , n16751 , n24021 );
    nor g11610 ( n27039 , n13897 , n13159 );
    not g11611 ( n10281 , n26645 );
    or g11612 ( n22838 , n15375 , n22483 );
    not g11613 ( n26883 , n3260 );
    or g11614 ( n25205 , n17588 , n5155 );
    xnor g11615 ( n16597 , n9026 , n11273 );
    or g11616 ( n9524 , n26411 , n3965 );
    nor g11617 ( n7994 , n3976 , n16882 );
    not g11618 ( n5466 , n2909 );
    or g11619 ( n26781 , n20250 , n1682 );
    xnor g11620 ( n1156 , n26594 , n18880 );
    nor g11621 ( n2251 , n1662 , n26962 );
    nor g11622 ( n8347 , n4692 , n26023 );
    or g11623 ( n19021 , n4412 , n22109 );
    or g11624 ( n8588 , n19862 , n16223 );
    xnor g11625 ( n13928 , n21841 , n17994 );
    xnor g11626 ( n16690 , n5077 , n13851 );
    or g11627 ( n16498 , n16374 , n23181 );
    not g11628 ( n2980 , n17558 );
    or g11629 ( n20282 , n18901 , n638 );
    and g11630 ( n7900 , n7264 , n21515 );
    xnor g11631 ( n17882 , n25568 , n16880 );
    and g11632 ( n9973 , n4229 , n26973 );
    xnor g11633 ( n24260 , n20937 , n7810 );
    or g11634 ( n178 , n26271 , n25152 );
    nor g11635 ( n9663 , n23487 , n26658 );
    and g11636 ( n12685 , n21983 , n25557 );
    not g11637 ( n8931 , n434 );
    or g11638 ( n22547 , n6393 , n2028 );
    not g11639 ( n22342 , n8660 );
    not g11640 ( n10821 , n19312 );
    nor g11641 ( n3326 , n13995 , n21981 );
    and g11642 ( n25030 , n7541 , n20632 );
    not g11643 ( n13643 , n3743 );
    or g11644 ( n24142 , n5675 , n5424 );
    not g11645 ( n25368 , n8933 );
    xnor g11646 ( n3884 , n12090 , n8487 );
    xnor g11647 ( n826 , n21095 , n11192 );
    not g11648 ( n19658 , n26226 );
    and g11649 ( n8120 , n5912 , n14990 );
    and g11650 ( n5463 , n21190 , n18458 );
    and g11651 ( n22847 , n17722 , n6792 );
    or g11652 ( n9357 , n26367 , n8930 );
    or g11653 ( n7159 , n21926 , n19468 );
    xnor g11654 ( n13144 , n18306 , n3726 );
    xnor g11655 ( n26239 , n5086 , n20670 );
    xnor g11656 ( n10076 , n21923 , n5637 );
    not g11657 ( n18393 , n18944 );
    and g11658 ( n9327 , n17828 , n11361 );
    or g11659 ( n23079 , n20782 , n4702 );
    or g11660 ( n24253 , n24772 , n24207 );
    not g11661 ( n14311 , n11414 );
    and g11662 ( n5268 , n15189 , n24320 );
    or g11663 ( n4689 , n16636 , n20877 );
    xnor g11664 ( n1435 , n8732 , n14127 );
    xnor g11665 ( n11799 , n6356 , n4665 );
    and g11666 ( n21072 , n2032 , n19782 );
    or g11667 ( n2673 , n12857 , n1931 );
    xnor g11668 ( n19216 , n26298 , n26625 );
    not g11669 ( n20525 , n9342 );
    and g11670 ( n25584 , n619 , n14880 );
    nor g11671 ( n706 , n10499 , n9512 );
    and g11672 ( n22286 , n7437 , n26992 );
    and g11673 ( n1030 , n20417 , n3568 );
    or g11674 ( n14303 , n18738 , n9457 );
    and g11675 ( n6818 , n17336 , n19812 );
    and g11676 ( n7977 , n19012 , n25456 );
    and g11677 ( n13679 , n19446 , n3931 );
    xnor g11678 ( n13216 , n9962 , n24028 );
    xnor g11679 ( n6403 , n7651 , n581 );
    not g11680 ( n12955 , n7139 );
    nor g11681 ( n23288 , n22351 , n24093 );
    or g11682 ( n25091 , n1280 , n24787 );
    or g11683 ( n14392 , n15009 , n12733 );
    and g11684 ( n22070 , n10338 , n425 );
    xnor g11685 ( n26794 , n12231 , n26821 );
    not g11686 ( n5319 , n6449 );
    or g11687 ( n16081 , n25941 , n9269 );
    or g11688 ( n17258 , n9869 , n16066 );
    or g11689 ( n17280 , n16227 , n6513 );
    xnor g11690 ( n9771 , n22852 , n18229 );
    nor g11691 ( n23228 , n26189 , n24180 );
    not g11692 ( n4299 , n1917 );
    xnor g11693 ( n15961 , n21041 , n7838 );
    and g11694 ( n25366 , n8429 , n16039 );
    and g11695 ( n10373 , n15258 , n2420 );
    xnor g11696 ( n21945 , n20525 , n12806 );
    nor g11697 ( n26760 , n5965 , n9200 );
    xnor g11698 ( n7507 , n16131 , n2922 );
    and g11699 ( n21286 , n5539 , n23019 );
    not g11700 ( n22398 , n21967 );
    or g11701 ( n21908 , n13490 , n6333 );
    nor g11702 ( n9239 , n9875 , n25562 );
    xnor g11703 ( n15548 , n11010 , n17183 );
    xnor g11704 ( n20633 , n12595 , n4682 );
    or g11705 ( n22720 , n14809 , n21736 );
    and g11706 ( n14525 , n18496 , n20201 );
    not g11707 ( n13053 , n7919 );
    xnor g11708 ( n24684 , n12193 , n10174 );
    or g11709 ( n1425 , n3499 , n14315 );
    nor g11710 ( n4904 , n16476 , n15539 );
    xnor g11711 ( n8862 , n22277 , n3628 );
    or g11712 ( n6050 , n24417 , n10027 );
    or g11713 ( n22041 , n7130 , n3075 );
    or g11714 ( n23590 , n1329 , n5512 );
    and g11715 ( n22022 , n17736 , n15951 );
    and g11716 ( n10300 , n7355 , n18273 );
    or g11717 ( n20256 , n329 , n6541 );
    or g11718 ( n10801 , n23478 , n12684 );
    nor g11719 ( n14920 , n11452 , n23068 );
    not g11720 ( n13286 , n6299 );
    or g11721 ( n21492 , n16750 , n9015 );
    xnor g11722 ( n4005 , n2009 , n7767 );
    xnor g11723 ( n14154 , n13206 , n17035 );
    and g11724 ( n5930 , n20742 , n26861 );
    not g11725 ( n22585 , n17090 );
    and g11726 ( n7717 , n7283 , n24915 );
    or g11727 ( n25821 , n14366 , n8477 );
    xnor g11728 ( n24439 , n23819 , n22861 );
    or g11729 ( n22900 , n773 , n12798 );
    xnor g11730 ( n24979 , n7657 , n25316 );
    not g11731 ( n7319 , n8526 );
    and g11732 ( n1582 , n13210 , n14890 );
    and g11733 ( n8554 , n18552 , n1315 );
    or g11734 ( n24424 , n18424 , n3837 );
    or g11735 ( n21805 , n9793 , n22361 );
    xor g11736 ( n6132 , n17339 , n6502 );
    xnor g11737 ( n15127 , n14903 , n9302 );
    or g11738 ( n20226 , n2766 , n18248 );
    nor g11739 ( n19310 , n10201 , n24043 );
    not g11740 ( n18741 , n15865 );
    not g11741 ( n19453 , n24171 );
    xnor g11742 ( n6998 , n14906 , n23565 );
    or g11743 ( n20571 , n23722 , n5324 );
    nor g11744 ( n12129 , n14902 , n4288 );
    or g11745 ( n19231 , n26027 , n19198 );
    xnor g11746 ( n14097 , n2035 , n12821 );
    not g11747 ( n11365 , n14749 );
    xnor g11748 ( n13736 , n5629 , n7377 );
    or g11749 ( n4671 , n20429 , n22909 );
    not g11750 ( n24455 , n25653 );
    xnor g11751 ( n6152 , n15769 , n13190 );
    or g11752 ( n23998 , n8820 , n13197 );
    not g11753 ( n5918 , n13951 );
    or g11754 ( n21618 , n18776 , n1770 );
    not g11755 ( n12554 , n16396 );
    xnor g11756 ( n24016 , n6068 , n18745 );
    not g11757 ( n20125 , n10204 );
    and g11758 ( n12155 , n9816 , n11 );
    or g11759 ( n8058 , n25283 , n13193 );
    or g11760 ( n18604 , n19949 , n11285 );
    xnor g11761 ( n25208 , n10079 , n1820 );
    and g11762 ( n14732 , n19133 , n19014 );
    not g11763 ( n6028 , n25302 );
    or g11764 ( n8479 , n15636 , n9656 );
    or g11765 ( n802 , n20089 , n5998 );
    nor g11766 ( n24290 , n26875 , n5530 );
    or g11767 ( n9907 , n5149 , n26703 );
    or g11768 ( n21991 , n24282 , n23712 );
    not g11769 ( n20538 , n1530 );
    and g11770 ( n24991 , n26213 , n24773 );
    or g11771 ( n714 , n14870 , n8888 );
    not g11772 ( n27030 , n22388 );
    or g11773 ( n16087 , n24338 , n20110 );
    not g11774 ( n23936 , n5818 );
    not g11775 ( n5045 , n21427 );
    xnor g11776 ( n6155 , n20338 , n9531 );
    not g11777 ( n22230 , n23763 );
    or g11778 ( n21617 , n18073 , n6767 );
    xnor g11779 ( n8246 , n19940 , n14705 );
    or g11780 ( n26996 , n18921 , n1028 );
    xnor g11781 ( n26780 , n8752 , n23796 );
    not g11782 ( n2204 , n24225 );
    or g11783 ( n26686 , n22597 , n16473 );
    xnor g11784 ( n8685 , n11503 , n18151 );
    and g11785 ( n20583 , n14431 , n22587 );
    and g11786 ( n11809 , n22590 , n19053 );
    not g11787 ( n25818 , n17591 );
    xnor g11788 ( n3897 , n1336 , n6265 );
    xnor g11789 ( n17557 , n12042 , n11514 );
    xnor g11790 ( n548 , n15067 , n11079 );
    and g11791 ( n13930 , n1252 , n23427 );
    and g11792 ( n12339 , n8048 , n13942 );
    or g11793 ( n12490 , n20737 , n20036 );
    or g11794 ( n26679 , n26532 , n526 );
    xnor g11795 ( n21968 , n15787 , n11408 );
    xnor g11796 ( n3708 , n18584 , n19803 );
    or g11797 ( n11388 , n4665 , n24278 );
    or g11798 ( n5725 , n15840 , n8364 );
    xnor g11799 ( n21244 , n8779 , n18290 );
    nor g11800 ( n11957 , n12639 , n26986 );
    xnor g11801 ( n24842 , n19983 , n18433 );
    xnor g11802 ( n22632 , n21517 , n8582 );
    xnor g11803 ( n8267 , n26040 , n17228 );
    xnor g11804 ( n17827 , n26536 , n4603 );
    and g11805 ( n13597 , n22337 , n19290 );
    xnor g11806 ( n3595 , n7829 , n12593 );
    or g11807 ( n17491 , n26007 , n15126 );
    xnor g11808 ( n18050 , n26870 , n25864 );
    or g11809 ( n5249 , n21760 , n11589 );
    xnor g11810 ( n19804 , n18590 , n25225 );
    or g11811 ( n22526 , n16730 , n11066 );
    or g11812 ( n7019 , n173 , n18008 );
    not g11813 ( n10109 , n11630 );
    and g11814 ( n19779 , n26398 , n17886 );
    not g11815 ( n10951 , n1200 );
    and g11816 ( n16695 , n2235 , n3556 );
    xnor g11817 ( n2535 , n6384 , n21788 );
    nor g11818 ( n20717 , n14777 , n3236 );
    not g11819 ( n21194 , n12430 );
    nor g11820 ( n23283 , n12709 , n19989 );
    and g11821 ( n17296 , n17995 , n4222 );
    and g11822 ( n9201 , n21186 , n2215 );
    xnor g11823 ( n8971 , n20656 , n9845 );
    or g11824 ( n23925 , n17414 , n19478 );
    xnor g11825 ( n25731 , n16468 , n17351 );
    nor g11826 ( n20311 , n14139 , n14838 );
    nor g11827 ( n3753 , n8068 , n1128 );
    xnor g11828 ( n10927 , n23383 , n771 );
    not g11829 ( n23664 , n2249 );
    not g11830 ( n5678 , n15245 );
    or g11831 ( n21641 , n9557 , n16158 );
    and g11832 ( n23132 , n16268 , n1647 );
    and g11833 ( n16159 , n11745 , n18249 );
    xnor g11834 ( n4966 , n19101 , n11797 );
    xnor g11835 ( n2788 , n15808 , n16713 );
    or g11836 ( n17868 , n27190 , n2531 );
    or g11837 ( n7955 , n18960 , n14982 );
    and g11838 ( n9254 , n11016 , n9883 );
    or g11839 ( n24255 , n11089 , n972 );
    xnor g11840 ( n21911 , n24509 , n18065 );
    and g11841 ( n1201 , n9652 , n901 );
    and g11842 ( n3536 , n23497 , n22413 );
    not g11843 ( n2219 , n1536 );
    not g11844 ( n10343 , n24992 );
    and g11845 ( n21304 , n18097 , n20354 );
    xnor g11846 ( n22321 , n7800 , n5626 );
    xnor g11847 ( n20647 , n1654 , n21997 );
    or g11848 ( n7021 , n14613 , n6777 );
    or g11849 ( n5379 , n22851 , n17610 );
    and g11850 ( n20887 , n22019 , n13064 );
    and g11851 ( n27103 , n10769 , n1174 );
    xnor g11852 ( n17168 , n9348 , n24712 );
    xnor g11853 ( n20301 , n7806 , n19933 );
    not g11854 ( n1173 , n14044 );
    or g11855 ( n15876 , n23894 , n4851 );
    xnor g11856 ( n10386 , n27114 , n4569 );
    or g11857 ( n3501 , n2459 , n24838 );
    and g11858 ( n15450 , n4971 , n9306 );
    not g11859 ( n167 , n10392 );
    nor g11860 ( n8546 , n17664 , n21253 );
    or g11861 ( n8337 , n7841 , n8952 );
    xnor g11862 ( n20219 , n24746 , n4119 );
    xnor g11863 ( n5904 , n2800 , n8584 );
    or g11864 ( n25003 , n25903 , n20697 );
    and g11865 ( n9234 , n6726 , n18202 );
    and g11866 ( n21692 , n25308 , n17777 );
    and g11867 ( n10813 , n14928 , n1614 );
    xnor g11868 ( n6543 , n16539 , n15362 );
    or g11869 ( n8074 , n5898 , n24182 );
    not g11870 ( n18742 , n19117 );
    xnor g11871 ( n5524 , n9674 , n24585 );
    and g11872 ( n2854 , n15068 , n5630 );
    and g11873 ( n23134 , n26984 , n24720 );
    or g11874 ( n6719 , n5016 , n12839 );
    or g11875 ( n22873 , n13593 , n13845 );
    or g11876 ( n25 , n11919 , n19037 );
    and g11877 ( n8021 , n15768 , n16592 );
    or g11878 ( n11035 , n2713 , n20479 );
    xnor g11879 ( n8944 , n19825 , n10117 );
    and g11880 ( n25727 , n20511 , n11272 );
    or g11881 ( n1305 , n15162 , n19936 );
    or g11882 ( n14898 , n20498 , n15486 );
    xnor g11883 ( n24932 , n20280 , n515 );
    xnor g11884 ( n6289 , n13596 , n7805 );
    xnor g11885 ( n3330 , n23822 , n1637 );
    xnor g11886 ( n19108 , n6053 , n1907 );
    not g11887 ( n23317 , n25178 );
    or g11888 ( n4899 , n5451 , n17858 );
    or g11889 ( n25374 , n21708 , n13604 );
    and g11890 ( n24313 , n26986 , n12639 );
    or g11891 ( n7552 , n25121 , n14161 );
    xnor g11892 ( n22251 , n9135 , n27147 );
    not g11893 ( n10509 , n17115 );
    xnor g11894 ( n20413 , n11979 , n6822 );
    or g11895 ( n15443 , n3996 , n20916 );
    and g11896 ( n22551 , n5941 , n7964 );
    not g11897 ( n9017 , n15821 );
    or g11898 ( n20419 , n1768 , n19069 );
    not g11899 ( n18755 , n17343 );
    xnor g11900 ( n827 , n11151 , n4295 );
    xnor g11901 ( n9513 , n8264 , n15765 );
    and g11902 ( n26597 , n11743 , n13301 );
    or g11903 ( n18783 , n12175 , n12949 );
    or g11904 ( n10099 , n4857 , n7193 );
    and g11905 ( n18365 , n15824 , n18490 );
    or g11906 ( n5723 , n6498 , n20906 );
    and g11907 ( n20449 , n23549 , n764 );
    xnor g11908 ( n26598 , n9743 , n17806 );
    or g11909 ( n25847 , n3589 , n18223 );
    or g11910 ( n3899 , n5466 , n10821 );
    or g11911 ( n10338 , n8991 , n20755 );
    or g11912 ( n11766 , n2579 , n3468 );
    xnor g11913 ( n25131 , n22631 , n2117 );
    and g11914 ( n11399 , n6602 , n24465 );
    or g11915 ( n4889 , n14963 , n3570 );
    xnor g11916 ( n26546 , n2028 , n17853 );
    and g11917 ( n23788 , n22554 , n1414 );
    or g11918 ( n8359 , n3204 , n12626 );
    nor g11919 ( n25025 , n19042 , n19360 );
    xnor g11920 ( n17206 , n8266 , n13495 );
    xnor g11921 ( n23999 , n17634 , n8687 );
    xnor g11922 ( n7719 , n9957 , n2659 );
    xnor g11923 ( n23509 , n11895 , n5451 );
    or g11924 ( n17540 , n13384 , n4459 );
    nor g11925 ( n1360 , n24473 , n3614 );
    or g11926 ( n6899 , n10 , n23407 );
    or g11927 ( n11761 , n528 , n13627 );
    or g11928 ( n13030 , n15369 , n12580 );
    and g11929 ( n21926 , n7722 , n154 );
    xnor g11930 ( n1237 , n3938 , n6481 );
    xnor g11931 ( n20333 , n8377 , n13155 );
    not g11932 ( n6708 , n25807 );
    or g11933 ( n24006 , n18425 , n7970 );
    and g11934 ( n21366 , n2026 , n14906 );
    and g11935 ( n17039 , n25904 , n20657 );
    and g11936 ( n1919 , n5594 , n15708 );
    or g11937 ( n4952 , n10736 , n4663 );
    xnor g11938 ( n15393 , n11151 , n21489 );
    xnor g11939 ( n8072 , n10622 , n265 );
    xnor g11940 ( n14107 , n9979 , n15805 );
    or g11941 ( n1789 , n15660 , n24814 );
    and g11942 ( n2372 , n2454 , n4970 );
    nor g11943 ( n9812 , n2804 , n18129 );
    not g11944 ( n602 , n1138 );
    xnor g11945 ( n3643 , n20089 , n16502 );
    or g11946 ( n9038 , n860 , n14330 );
    and g11947 ( n6102 , n2278 , n7093 );
    not g11948 ( n23995 , n25689 );
    nor g11949 ( n5437 , n7693 , n19472 );
    not g11950 ( n24624 , n2525 );
    xnor g11951 ( n19495 , n20604 , n21735 );
    nor g11952 ( n23744 , n2816 , n26486 );
    not g11953 ( n16064 , n25520 );
    nor g11954 ( n6408 , n2562 , n8244 );
    xnor g11955 ( n20483 , n21400 , n19081 );
    not g11956 ( n7745 , n22495 );
    xnor g11957 ( n3976 , n23975 , n16645 );
    or g11958 ( n18479 , n9655 , n21908 );
    nor g11959 ( n14740 , n6613 , n6703 );
    not g11960 ( n13729 , n9172 );
    and g11961 ( n23972 , n16836 , n10798 );
    xnor g11962 ( n11670 , n26352 , n22679 );
    xnor g11963 ( n20651 , n26962 , n3730 );
    or g11964 ( n1583 , n12354 , n19321 );
    or g11965 ( n23461 , n19139 , n211 );
    and g11966 ( n12082 , n11038 , n10058 );
    not g11967 ( n17923 , n26291 );
    xnor g11968 ( n22691 , n10451 , n17741 );
    or g11969 ( n2425 , n13783 , n26394 );
    nor g11970 ( n1929 , n19476 , n2325 );
    xnor g11971 ( n21527 , n20899 , n11960 );
    or g11972 ( n16139 , n18981 , n11381 );
    xnor g11973 ( n22372 , n9569 , n21317 );
    and g11974 ( n4364 , n13307 , n14784 );
    xnor g11975 ( n24793 , n24990 , n19502 );
    or g11976 ( n4192 , n21841 , n16295 );
    or g11977 ( n16189 , n23436 , n9003 );
    xnor g11978 ( n5541 , n21764 , n23529 );
    not g11979 ( n18383 , n6861 );
    xnor g11980 ( n17317 , n13108 , n11174 );
    xnor g11981 ( n3219 , n23396 , n1121 );
    xnor g11982 ( n14772 , n19879 , n2282 );
    and g11983 ( n11656 , n7948 , n1583 );
    xnor g11984 ( n17982 , n1967 , n26989 );
    nor g11985 ( n23560 , n24116 , n20929 );
    or g11986 ( n2028 , n19082 , n24630 );
    and g11987 ( n20405 , n4242 , n17388 );
    or g11988 ( n24635 , n1365 , n25924 );
    or g11989 ( n3450 , n15905 , n2510 );
    xnor g11990 ( n25660 , n24902 , n8623 );
    or g11991 ( n26388 , n23539 , n14488 );
    or g11992 ( n12957 , n7722 , n154 );
    xnor g11993 ( n2696 , n15605 , n22575 );
    not g11994 ( n12239 , n13734 );
    and g11995 ( n3938 , n4142 , n19504 );
    xnor g11996 ( n19886 , n10615 , n6078 );
    or g11997 ( n22148 , n23216 , n15093 );
    nor g11998 ( n26428 , n1181 , n11428 );
    not g11999 ( n14612 , n1949 );
    not g12000 ( n24180 , n8358 );
    and g12001 ( n15141 , n26372 , n8080 );
    xnor g12002 ( n14796 , n2218 , n18483 );
    xnor g12003 ( n6996 , n11869 , n20198 );
    or g12004 ( n2803 , n4258 , n25922 );
    and g12005 ( n14522 , n26858 , n17327 );
    nor g12006 ( n20474 , n25972 , n21378 );
    nor g12007 ( n23119 , n14744 , n17936 );
    or g12008 ( n1094 , n16625 , n15032 );
    and g12009 ( n23080 , n15595 , n20781 );
    nor g12010 ( n26514 , n4040 , n3349 );
    xnor g12011 ( n21225 , n16122 , n4115 );
    and g12012 ( n8670 , n20622 , n25880 );
    and g12013 ( n15726 , n1588 , n22229 );
    or g12014 ( n12280 , n20613 , n14138 );
    nor g12015 ( n7286 , n1406 , n4940 );
    not g12016 ( n2432 , n10116 );
    nor g12017 ( n8252 , n18290 , n25160 );
    or g12018 ( n3765 , n11187 , n547 );
    xnor g12019 ( n422 , n651 , n11845 );
    or g12020 ( n27203 , n866 , n9449 );
    and g12021 ( n1065 , n14420 , n15664 );
    not g12022 ( n1533 , n8724 );
    nor g12023 ( n15134 , n9679 , n22442 );
    not g12024 ( n88 , n25164 );
    xnor g12025 ( n248 , n20569 , n14120 );
    and g12026 ( n18530 , n7566 , n22640 );
    xnor g12027 ( n18820 , n19946 , n12627 );
    nor g12028 ( n23351 , n15058 , n1532 );
    and g12029 ( n6461 , n603 , n16505 );
    nor g12030 ( n4977 , n4003 , n22507 );
    xnor g12031 ( n14531 , n2242 , n12810 );
    or g12032 ( n2672 , n16575 , n2379 );
    xnor g12033 ( n12667 , n19090 , n20271 );
    not g12034 ( n26580 , n21540 );
    xnor g12035 ( n9085 , n3228 , n22470 );
    or g12036 ( n3432 , n17014 , n17646 );
    and g12037 ( n26637 , n20318 , n13345 );
    not g12038 ( n3587 , n24399 );
    xnor g12039 ( n7913 , n19234 , n21398 );
    and g12040 ( n12359 , n19731 , n23993 );
    xnor g12041 ( n13217 , n4708 , n19216 );
    not g12042 ( n20099 , n9219 );
    nor g12043 ( n24845 , n12481 , n9227 );
    not g12044 ( n11485 , n26708 );
    or g12045 ( n6261 , n22919 , n23044 );
    xnor g12046 ( n742 , n25465 , n26530 );
    not g12047 ( n14269 , n2969 );
    and g12048 ( n20743 , n4854 , n23862 );
    or g12049 ( n16495 , n4574 , n25715 );
    nor g12050 ( n16103 , n18995 , n17143 );
    xnor g12051 ( n13122 , n7483 , n10774 );
    or g12052 ( n20922 , n13154 , n3918 );
    or g12053 ( n24317 , n8352 , n22960 );
    xnor g12054 ( n15598 , n18547 , n26504 );
    or g12055 ( n6103 , n5122 , n6483 );
    xnor g12056 ( n881 , n8814 , n21158 );
    or g12057 ( n20123 , n5924 , n16201 );
    and g12058 ( n7217 , n18300 , n9411 );
    xnor g12059 ( n5851 , n17626 , n2246 );
    xnor g12060 ( n8375 , n10152 , n7981 );
    or g12061 ( n5352 , n5025 , n23162 );
    and g12062 ( n11959 , n6908 , n9098 );
    nor g12063 ( n4208 , n25036 , n11016 );
    or g12064 ( n21169 , n417 , n4499 );
    or g12065 ( n14825 , n13367 , n13074 );
    xnor g12066 ( n6329 , n6492 , n20835 );
    xnor g12067 ( n26964 , n6827 , n6055 );
    xnor g12068 ( n24934 , n25340 , n76 );
    xnor g12069 ( n18512 , n1505 , n26036 );
    xnor g12070 ( n17993 , n19182 , n22563 );
    xnor g12071 ( n4184 , n10784 , n6881 );
    or g12072 ( n14312 , n10985 , n24122 );
    or g12073 ( n13542 , n13224 , n21089 );
    nor g12074 ( n1568 , n24355 , n1267 );
    or g12075 ( n18415 , n11315 , n24918 );
    xnor g12076 ( n21203 , n25060 , n14832 );
    or g12077 ( n2033 , n13184 , n13962 );
    xnor g12078 ( n1552 , n7442 , n8767 );
    nor g12079 ( n20680 , n8987 , n14245 );
    not g12080 ( n4938 , n23463 );
    xnor g12081 ( n12754 , n7073 , n13010 );
    xnor g12082 ( n5742 , n15329 , n13135 );
    or g12083 ( n25469 , n6877 , n9108 );
    or g12084 ( n11190 , n19732 , n14296 );
    xnor g12085 ( n1820 , n1163 , n18901 );
    nor g12086 ( n15711 , n15905 , n23168 );
    xnor g12087 ( n17219 , n25148 , n21521 );
    or g12088 ( n322 , n21083 , n7520 );
    xnor g12089 ( n6783 , n9485 , n12147 );
    or g12090 ( n11620 , n16056 , n13540 );
    xnor g12091 ( n3311 , n413 , n5409 );
    or g12092 ( n8421 , n14306 , n2599 );
    or g12093 ( n24195 , n12582 , n6681 );
    or g12094 ( n14595 , n23141 , n22981 );
    xnor g12095 ( n8946 , n8399 , n8052 );
    not g12096 ( n17660 , n1512 );
    not g12097 ( n868 , n4775 );
    xnor g12098 ( n5286 , n20040 , n9396 );
    xnor g12099 ( n13963 , n25558 , n18904 );
    xnor g12100 ( n1518 , n18127 , n2402 );
    not g12101 ( n13989 , n19494 );
    xnor g12102 ( n76 , n15447 , n6838 );
    xnor g12103 ( n4204 , n3926 , n492 );
    or g12104 ( n25308 , n19383 , n10422 );
    xnor g12105 ( n24704 , n1485 , n24518 );
    not g12106 ( n18189 , n4626 );
    nor g12107 ( n15368 , n18419 , n22005 );
    not g12108 ( n13124 , n16392 );
    xnor g12109 ( n7210 , n17156 , n4872 );
    nor g12110 ( n21421 , n19634 , n2731 );
    xnor g12111 ( n710 , n17894 , n1982 );
    or g12112 ( n17707 , n18649 , n11278 );
    xnor g12113 ( n6924 , n15731 , n12300 );
    or g12114 ( n8095 , n10002 , n21861 );
    xnor g12115 ( n8933 , n19120 , n16027 );
    xnor g12116 ( n25539 , n15755 , n14468 );
    or g12117 ( n16838 , n4709 , n16088 );
    or g12118 ( n21528 , n18926 , n2705 );
    not g12119 ( n24774 , n2059 );
    and g12120 ( n18402 , n6007 , n24641 );
    or g12121 ( n26281 , n25190 , n24281 );
    and g12122 ( n7227 , n18415 , n19369 );
    or g12123 ( n16165 , n11486 , n13781 );
    buf g12124 ( n24286 , n14083 );
    and g12125 ( n21684 , n24670 , n2182 );
    not g12126 ( n21107 , n9274 );
    or g12127 ( n25317 , n337 , n5340 );
    xnor g12128 ( n8331 , n11661 , n324 );
    and g12129 ( n2260 , n23537 , n11010 );
    or g12130 ( n2373 , n22487 , n13645 );
    xnor g12131 ( n11525 , n11608 , n17693 );
    xnor g12132 ( n18544 , n21276 , n18157 );
    xnor g12133 ( n19312 , n17659 , n3833 );
    or g12134 ( n23672 , n24845 , n9641 );
    xnor g12135 ( n3563 , n14235 , n9796 );
    not g12136 ( n20620 , n3830 );
    or g12137 ( n20294 , n23320 , n19564 );
    buf g12138 ( n20920 , n18953 );
    not g12139 ( n13353 , n5834 );
    nor g12140 ( n7921 , n14612 , n20169 );
    and g12141 ( n5225 , n10395 , n15476 );
    or g12142 ( n25951 , n22994 , n9025 );
    not g12143 ( n9780 , n9749 );
    xnor g12144 ( n15090 , n19023 , n8330 );
    xnor g12145 ( n22090 , n188 , n25551 );
    not g12146 ( n7448 , n13257 );
    and g12147 ( n12175 , n22820 , n19137 );
    or g12148 ( n5871 , n4544 , n23701 );
    xnor g12149 ( n21502 , n8287 , n12483 );
    xnor g12150 ( n19432 , n5318 , n3943 );
    or g12151 ( n12537 , n12673 , n21529 );
    or g12152 ( n573 , n21701 , n21547 );
    xnor g12153 ( n9980 , n4570 , n17458 );
    not g12154 ( n11577 , n18729 );
    or g12155 ( n13382 , n8068 , n11192 );
    and g12156 ( n6808 , n10575 , n7246 );
    and g12157 ( n16943 , n6859 , n17600 );
    and g12158 ( n17818 , n17675 , n26412 );
    and g12159 ( n19983 , n26976 , n22947 );
    or g12160 ( n1627 , n5883 , n20764 );
    xnor g12161 ( n15093 , n1787 , n10618 );
    nor g12162 ( n6320 , n12204 , n22478 );
    nor g12163 ( n23425 , n14967 , n20013 );
    or g12164 ( n15035 , n23464 , n25966 );
    xnor g12165 ( n26847 , n5676 , n22381 );
    or g12166 ( n17158 , n22749 , n5468 );
    or g12167 ( n11530 , n6051 , n593 );
    and g12168 ( n18528 , n5349 , n3990 );
    not g12169 ( n19194 , n25383 );
    and g12170 ( n20711 , n13898 , n7311 );
    or g12171 ( n12083 , n11941 , n1890 );
    or g12172 ( n24108 , n888 , n25977 );
    or g12173 ( n15525 , n23631 , n24935 );
    xnor g12174 ( n15205 , n16686 , n14047 );
    or g12175 ( n2871 , n832 , n11938 );
    not g12176 ( n14969 , n6891 );
    xnor g12177 ( n722 , n3045 , n4201 );
    not g12178 ( n6089 , n9168 );
    nor g12179 ( n18014 , n19085 , n24592 );
    or g12180 ( n3023 , n113 , n2604 );
    and g12181 ( n3101 , n7046 , n7853 );
    and g12182 ( n9331 , n10646 , n12106 );
    and g12183 ( n26410 , n20237 , n13111 );
    or g12184 ( n9544 , n1427 , n25497 );
    xnor g12185 ( n18089 , n9942 , n10739 );
    not g12186 ( n6063 , n2443 );
    xnor g12187 ( n224 , n1928 , n21256 );
    or g12188 ( n9560 , n14710 , n2219 );
    or g12189 ( n4337 , n23852 , n17430 );
    not g12190 ( n26895 , n6794 );
    or g12191 ( n24303 , n6813 , n14347 );
    or g12192 ( n20101 , n5727 , n3477 );
    xnor g12193 ( n22340 , n5681 , n9461 );
    xnor g12194 ( n9194 , n11099 , n915 );
    xnor g12195 ( n23888 , n4147 , n6700 );
    nor g12196 ( n18717 , n2155 , n7097 );
    xnor g12197 ( n14106 , n19772 , n2571 );
    or g12198 ( n20739 , n18749 , n4156 );
    or g12199 ( n12830 , n15447 , n24951 );
    xnor g12200 ( n14136 , n16198 , n8184 );
    or g12201 ( n5546 , n16534 , n5070 );
    or g12202 ( n6118 , n26052 , n8054 );
    and g12203 ( n12689 , n26555 , n18795 );
    xnor g12204 ( n25892 , n22260 , n10964 );
    nor g12205 ( n23728 , n6502 , n19494 );
    and g12206 ( n25107 , n9894 , n14793 );
    and g12207 ( n7243 , n10247 , n14253 );
    and g12208 ( n18013 , n6369 , n527 );
    or g12209 ( n22823 , n7377 , n21125 );
    or g12210 ( n20341 , n4502 , n25536 );
    or g12211 ( n13078 , n4022 , n13110 );
    not g12212 ( n20175 , n4122 );
    xnor g12213 ( n21533 , n6713 , n14528 );
    and g12214 ( n7816 , n22996 , n163 );
    or g12215 ( n11400 , n6239 , n25685 );
    or g12216 ( n3262 , n13223 , n5545 );
    and g12217 ( n13609 , n27157 , n16802 );
    or g12218 ( n9810 , n20466 , n23323 );
    or g12219 ( n26542 , n10743 , n26584 );
    or g12220 ( n24463 , n4727 , n11207 );
    xnor g12221 ( n21173 , n12721 , n24095 );
    xnor g12222 ( n24258 , n2317 , n25385 );
    xnor g12223 ( n8417 , n17146 , n12207 );
    and g12224 ( n26714 , n24240 , n4406 );
    and g12225 ( n25975 , n6735 , n6045 );
    or g12226 ( n19929 , n3074 , n2220 );
    and g12227 ( n13911 , n26481 , n16976 );
    nor g12228 ( n20070 , n2187 , n9572 );
    xnor g12229 ( n14102 , n90 , n23994 );
    nor g12230 ( n2807 , n305 , n2610 );
    or g12231 ( n8601 , n18742 , n14319 );
    xnor g12232 ( n24289 , n25039 , n5279 );
    xnor g12233 ( n18395 , n11197 , n17766 );
    and g12234 ( n26154 , n22985 , n3156 );
    and g12235 ( n10463 , n23216 , n15093 );
    xnor g12236 ( n4221 , n3774 , n7754 );
    xnor g12237 ( n6043 , n13322 , n18698 );
    or g12238 ( n27205 , n23091 , n18735 );
    and g12239 ( n4733 , n13452 , n9743 );
    not g12240 ( n10486 , n6279 );
    xnor g12241 ( n947 , n11628 , n17325 );
    xnor g12242 ( n2761 , n21452 , n9467 );
    not g12243 ( n4497 , n10185 );
    xnor g12244 ( n24393 , n1380 , n3324 );
    or g12245 ( n7858 , n7003 , n2480 );
    nor g12246 ( n5612 , n1346 , n442 );
    or g12247 ( n21199 , n12178 , n7116 );
    or g12248 ( n11972 , n6154 , n23996 );
    nor g12249 ( n9948 , n25265 , n23773 );
    or g12250 ( n12597 , n25331 , n2189 );
    not g12251 ( n24343 , n26733 );
    nor g12252 ( n1829 , n18855 , n20925 );
    not g12253 ( n10277 , n18006 );
    or g12254 ( n23226 , n22176 , n120 );
    xnor g12255 ( n2275 , n21520 , n19615 );
    and g12256 ( n19330 , n8305 , n2918 );
    or g12257 ( n19656 , n23306 , n9201 );
    nor g12258 ( n20956 , n27008 , n21194 );
    or g12259 ( n10748 , n20200 , n9156 );
    not g12260 ( n2223 , n881 );
    or g12261 ( n26671 , n15842 , n12606 );
    nor g12262 ( n25882 , n3018 , n2731 );
    not g12263 ( n24815 , n14380 );
    xnor g12264 ( n26620 , n6385 , n18171 );
    xnor g12265 ( n25202 , n14596 , n23635 );
    xnor g12266 ( n3118 , n520 , n6593 );
    not g12267 ( n2919 , n25355 );
    nor g12268 ( n773 , n23095 , n1112 );
    or g12269 ( n2139 , n26318 , n15860 );
    not g12270 ( n7938 , n22378 );
    or g12271 ( n24502 , n4113 , n21278 );
    xnor g12272 ( n8863 , n12878 , n14539 );
    not g12273 ( n10157 , n19335 );
    xnor g12274 ( n2320 , n17695 , n7692 );
    xnor g12275 ( n2491 , n23098 , n4434 );
    or g12276 ( n21501 , n17035 , n1872 );
    or g12277 ( n18164 , n9539 , n12255 );
    and g12278 ( n1579 , n20912 , n2245 );
    xnor g12279 ( n5737 , n9621 , n17367 );
    and g12280 ( n606 , n14242 , n12595 );
    and g12281 ( n21770 , n14529 , n9477 );
    xnor g12282 ( n22400 , n25073 , n12152 );
    xnor g12283 ( n13812 , n12232 , n3740 );
    not g12284 ( n10948 , n16945 );
    xnor g12285 ( n9984 , n4469 , n960 );
    and g12286 ( n25141 , n20890 , n24952 );
    xnor g12287 ( n17415 , n20797 , n2978 );
    and g12288 ( n20529 , n18278 , n19932 );
    xnor g12289 ( n12357 , n1639 , n5128 );
    xnor g12290 ( n16965 , n5450 , n5469 );
    and g12291 ( n3048 , n18026 , n6188 );
    and g12292 ( n21810 , n8440 , n2304 );
    nor g12293 ( n3029 , n2698 , n16961 );
    xnor g12294 ( n8174 , n12612 , n20794 );
    xnor g12295 ( n21324 , n24751 , n8604 );
    xnor g12296 ( n12660 , n6812 , n2614 );
    xnor g12297 ( n26639 , n7331 , n12171 );
    xnor g12298 ( n10139 , n21322 , n25345 );
    or g12299 ( n4525 , n7378 , n634 );
    xnor g12300 ( n6661 , n2926 , n12586 );
    not g12301 ( n6357 , n24788 );
    or g12302 ( n17451 , n9832 , n11831 );
    nor g12303 ( n7941 , n8813 , n10770 );
    or g12304 ( n1676 , n7590 , n16413 );
    or g12305 ( n10830 , n22257 , n22287 );
    or g12306 ( n5245 , n17188 , n24408 );
    or g12307 ( n14711 , n48 , n1309 );
    xnor g12308 ( n1200 , n24323 , n6775 );
    xnor g12309 ( n22508 , n2976 , n13262 );
    nor g12310 ( n8447 , n17718 , n7020 );
    and g12311 ( n4611 , n418 , n16726 );
    nor g12312 ( n15847 , n10116 , n15017 );
    xnor g12313 ( n4151 , n19994 , n6329 );
    or g12314 ( n6224 , n26469 , n3867 );
    or g12315 ( n14592 , n12261 , n22221 );
    or g12316 ( n14530 , n544 , n8170 );
    and g12317 ( n17437 , n12759 , n18156 );
    or g12318 ( n22676 , n8875 , n259 );
    xnor g12319 ( n14121 , n13272 , n25346 );
    nor g12320 ( n10677 , n20369 , n19034 );
    not g12321 ( n9597 , n7241 );
    not g12322 ( n6079 , n19660 );
    not g12323 ( n4361 , n6335 );
    xnor g12324 ( n5139 , n19273 , n18347 );
    nor g12325 ( n540 , n17679 , n8414 );
    or g12326 ( n14291 , n288 , n2144 );
    or g12327 ( n1441 , n6510 , n20482 );
    or g12328 ( n14653 , n26895 , n6611 );
    and g12329 ( n17 , n6274 , n3277 );
    or g12330 ( n1390 , n6892 , n14428 );
    nor g12331 ( n12021 , n3241 , n13944 );
    or g12332 ( n12690 , n5553 , n18716 );
    xnor g12333 ( n26237 , n20762 , n2468 );
    and g12334 ( n11872 , n17698 , n10450 );
    or g12335 ( n9579 , n18056 , n2474 );
    and g12336 ( n4974 , n18794 , n16038 );
    not g12337 ( n16294 , n11220 );
    xnor g12338 ( n18208 , n6385 , n8869 );
    nor g12339 ( n15244 , n17664 , n7532 );
    or g12340 ( n27056 , n6061 , n12685 );
    xnor g12341 ( n14480 , n2538 , n19857 );
    nor g12342 ( n7109 , n25779 , n26161 );
    not g12343 ( n13205 , n10792 );
    or g12344 ( n3655 , n11481 , n23493 );
    and g12345 ( n9134 , n5149 , n26703 );
    or g12346 ( n27077 , n3784 , n13121 );
    or g12347 ( n25286 , n6485 , n18676 );
    or g12348 ( n4305 , n3519 , n7687 );
    or g12349 ( n403 , n6811 , n10860 );
    and g12350 ( n24809 , n3213 , n8143 );
    and g12351 ( n22226 , n10568 , n5848 );
    and g12352 ( n22661 , n27000 , n6292 );
    nor g12353 ( n18408 , n10324 , n9779 );
    not g12354 ( n2377 , n25204 );
    or g12355 ( n19870 , n13629 , n3693 );
    and g12356 ( n4258 , n4086 , n1533 );
    or g12357 ( n22060 , n21857 , n10861 );
    xnor g12358 ( n13022 , n7969 , n21827 );
    xnor g12359 ( n21731 , n21113 , n16019 );
    nor g12360 ( n13390 , n25376 , n1752 );
    not g12361 ( n12048 , n2055 );
    or g12362 ( n15089 , n7360 , n18598 );
    xnor g12363 ( n9709 , n2586 , n11743 );
    not g12364 ( n22227 , n2244 );
    nor g12365 ( n5144 , n26703 , n7615 );
    and g12366 ( n25935 , n15018 , n8426 );
    and g12367 ( n4597 , n11200 , n8723 );
    nor g12368 ( n8567 , n4301 , n16330 );
    or g12369 ( n694 , n22958 , n19157 );
    and g12370 ( n1852 , n24811 , n11500 );
    xnor g12371 ( n15820 , n10351 , n26318 );
    and g12372 ( n201 , n5467 , n19110 );
    xnor g12373 ( n16902 , n24952 , n22371 );
    xnor g12374 ( n22378 , n26166 , n4124 );
    and g12375 ( n9025 , n13254 , n24570 );
    not g12376 ( n1786 , n9605 );
    xnor g12377 ( n8608 , n17340 , n15303 );
    nor g12378 ( n16635 , n19610 , n18539 );
    xnor g12379 ( n8725 , n1577 , n14405 );
    or g12380 ( n20577 , n17789 , n15337 );
    not g12381 ( n19258 , n8943 );
    or g12382 ( n25116 , n8301 , n20449 );
    xnor g12383 ( n5568 , n24850 , n22706 );
    nor g12384 ( n2585 , n3740 , n2545 );
    and g12385 ( n23280 , n16628 , n7028 );
    not g12386 ( n8771 , n10104 );
    xnor g12387 ( n16262 , n20289 , n9300 );
    or g12388 ( n8426 , n14479 , n17060 );
    not g12389 ( n26601 , n13471 );
    xnor g12390 ( n23423 , n17483 , n18504 );
    and g12391 ( n24104 , n26494 , n365 );
    or g12392 ( n1548 , n22443 , n23938 );
    or g12393 ( n22864 , n5084 , n8011 );
    xnor g12394 ( n4734 , n22350 , n2747 );
    or g12395 ( n20974 , n12932 , n22370 );
    or g12396 ( n6372 , n6724 , n11329 );
    xnor g12397 ( n3606 , n4074 , n15593 );
    and g12398 ( n5973 , n3487 , n20889 );
    nor g12399 ( n11256 , n22723 , n20923 );
    or g12400 ( n26157 , n25721 , n24067 );
    nor g12401 ( n17192 , n18909 , n18203 );
    and g12402 ( n13891 , n576 , n13969 );
    and g12403 ( n5305 , n2840 , n19079 );
    xnor g12404 ( n8088 , n13046 , n15216 );
    or g12405 ( n3858 , n13659 , n14932 );
    not g12406 ( n14777 , n22079 );
    xnor g12407 ( n2295 , n24403 , n26768 );
    not g12408 ( n7058 , n24860 );
    xnor g12409 ( n26741 , n290 , n24086 );
    xor g12410 ( n497 , n7242 , n3311 );
    or g12411 ( n18138 , n17120 , n7751 );
    or g12412 ( n5003 , n446 , n25318 );
    xnor g12413 ( n2929 , n929 , n1376 );
    and g12414 ( n21381 , n1407 , n7655 );
    xnor g12415 ( n8898 , n14417 , n3054 );
    or g12416 ( n23396 , n8931 , n24809 );
    xnor g12417 ( n6342 , n12068 , n18535 );
    xnor g12418 ( n8519 , n4508 , n5357 );
    or g12419 ( n3081 , n14080 , n24494 );
    and g12420 ( n10782 , n22081 , n21382 );
    not g12421 ( n8539 , n21073 );
    xnor g12422 ( n4836 , n11985 , n18116 );
    xnor g12423 ( n5296 , n14348 , n22393 );
    or g12424 ( n15321 , n963 , n13071 );
    xnor g12425 ( n23855 , n1844 , n21300 );
    xnor g12426 ( n10692 , n9891 , n14461 );
    or g12427 ( n1967 , n26895 , n5512 );
    not g12428 ( n9859 , n22325 );
    xnor g12429 ( n6022 , n4488 , n15803 );
    nor g12430 ( n2063 , n6685 , n19971 );
    not g12431 ( n12345 , n16150 );
    or g12432 ( n15367 , n25099 , n4442 );
    nor g12433 ( n9782 , n12161 , n106 );
    and g12434 ( n5955 , n11424 , n12692 );
    xnor g12435 ( n6135 , n14045 , n9936 );
    or g12436 ( n8541 , n18008 , n17869 );
    not g12437 ( n7350 , n1910 );
    xnor g12438 ( n17651 , n1837 , n9961 );
    xnor g12439 ( n26102 , n26997 , n19059 );
    and g12440 ( n7863 , n25747 , n17661 );
    nor g12441 ( n20865 , n20284 , n3779 );
    not g12442 ( n16466 , n19845 );
    and g12443 ( n27073 , n10604 , n17424 );
    xnor g12444 ( n21157 , n12711 , n3436 );
    xor g12445 ( n11377 , n10164 , n12983 );
    and g12446 ( n3802 , n8556 , n18259 );
    xnor g12447 ( n20096 , n22614 , n8234 );
    or g12448 ( n21611 , n580 , n3053 );
    or g12449 ( n19992 , n3150 , n24929 );
    xnor g12450 ( n24972 , n21112 , n8309 );
    nor g12451 ( n10323 , n14695 , n10125 );
    xnor g12452 ( n9873 , n508 , n12518 );
    and g12453 ( n1322 , n8101 , n21912 );
    xnor g12454 ( n23401 , n5118 , n25944 );
    not g12455 ( n3625 , n19478 );
    and g12456 ( n16934 , n19440 , n27198 );
    and g12457 ( n13564 , n8851 , n15212 );
    or g12458 ( n16926 , n10097 , n18002 );
    xnor g12459 ( n17417 , n21912 , n15241 );
    and g12460 ( n9211 , n18136 , n24976 );
    and g12461 ( n5412 , n4919 , n17222 );
    or g12462 ( n5021 , n24383 , n6403 );
    xnor g12463 ( n2478 , n1777 , n21832 );
    or g12464 ( n383 , n14930 , n4002 );
    xnor g12465 ( n11395 , n17295 , n14289 );
    not g12466 ( n24239 , n6095 );
    not g12467 ( n22562 , n9986 );
    nor g12468 ( n16216 , n5112 , n5417 );
    xnor g12469 ( n12617 , n20365 , n22571 );
    xor g12470 ( n7886 , n19110 , n2470 );
    or g12471 ( n10852 , n22123 , n82 );
    and g12472 ( n24214 , n1338 , n27180 );
    xnor g12473 ( n8028 , n21291 , n218 );
    or g12474 ( n8189 , n4514 , n5111 );
    or g12475 ( n6294 , n5558 , n23280 );
    xnor g12476 ( n24226 , n19871 , n25996 );
    or g12477 ( n6771 , n5499 , n17773 );
    xnor g12478 ( n13247 , n25074 , n10053 );
    not g12479 ( n7561 , n48 );
    xnor g12480 ( n23874 , n1817 , n159 );
    xnor g12481 ( n26789 , n14317 , n25797 );
    nor g12482 ( n8868 , n4699 , n16946 );
    not g12483 ( n17286 , n24768 );
    and g12484 ( n12316 , n596 , n22790 );
    xnor g12485 ( n22326 , n25855 , n26461 );
    xnor g12486 ( n8649 , n8652 , n16973 );
    xnor g12487 ( n26968 , n20794 , n23333 );
    or g12488 ( n25433 , n102 , n15192 );
    and g12489 ( n7012 , n21134 , n4930 );
    not g12490 ( n6235 , n7100 );
    or g12491 ( n26349 , n4942 , n13147 );
    not g12492 ( n3946 , n1714 );
    and g12493 ( n22074 , n6218 , n9296 );
    or g12494 ( n895 , n14519 , n3164 );
    xnor g12495 ( n10547 , n9942 , n23923 );
    not g12496 ( n19444 , n23258 );
    not g12497 ( n25405 , n25251 );
    and g12498 ( n24122 , n4655 , n16629 );
    xnor g12499 ( n8982 , n21657 , n22241 );
    or g12500 ( n9082 , n8032 , n14394 );
    and g12501 ( n23523 , n8667 , n16977 );
    or g12502 ( n22500 , n2997 , n6445 );
    xnor g12503 ( n24859 , n17090 , n22173 );
    and g12504 ( n15851 , n10641 , n3469 );
    and g12505 ( n15486 , n158 , n21053 );
    xnor g12506 ( n18315 , n9557 , n24170 );
    and g12507 ( n16089 , n16606 , n5896 );
    xnor g12508 ( n10665 , n22274 , n22591 );
    or g12509 ( n11892 , n16147 , n11367 );
    not g12510 ( n18103 , n7249 );
    and g12511 ( n4223 , n6734 , n3 );
    not g12512 ( n19003 , n6082 );
    not g12513 ( n3485 , n450 );
    xnor g12514 ( n4215 , n18930 , n9126 );
    xnor g12515 ( n14946 , n6492 , n17718 );
    xnor g12516 ( n13621 , n13252 , n9463 );
    and g12517 ( n25841 , n20425 , n12332 );
    and g12518 ( n19526 , n14724 , n9555 );
    or g12519 ( n25832 , n12014 , n1222 );
    and g12520 ( n15173 , n21261 , n18204 );
    xnor g12521 ( n19751 , n2876 , n19193 );
    xnor g12522 ( n18619 , n11670 , n16439 );
    xor g12523 ( n15346 , n24624 , n21095 );
    not g12524 ( n22176 , n6773 );
    xnor g12525 ( n6254 , n4065 , n7479 );
    and g12526 ( n20224 , n20470 , n14052 );
    xnor g12527 ( n6894 , n7311 , n13781 );
    xnor g12528 ( n22203 , n22619 , n6775 );
    and g12529 ( n16012 , n528 , n17556 );
    or g12530 ( n927 , n1319 , n3448 );
    or g12531 ( n3705 , n14091 , n6693 );
    not g12532 ( n19527 , n24049 );
    not g12533 ( n21842 , n10392 );
    xnor g12534 ( n6133 , n23486 , n16663 );
    nor g12535 ( n3473 , n15883 , n11096 );
    and g12536 ( n9091 , n12508 , n25942 );
    or g12537 ( n17834 , n22290 , n12562 );
    xnor g12538 ( n14437 , n23447 , n11225 );
    and g12539 ( n2284 , n20503 , n5153 );
    and g12540 ( n17614 , n21954 , n21548 );
    not g12541 ( n5875 , n15119 );
    xnor g12542 ( n11108 , n8436 , n16167 );
    xnor g12543 ( n22928 , n8381 , n18295 );
    not g12544 ( n16129 , n20040 );
    and g12545 ( n21878 , n24780 , n16134 );
    or g12546 ( n26142 , n18035 , n92 );
    xnor g12547 ( n2116 , n7892 , n15734 );
    nor g12548 ( n3811 , n26508 , n61 );
    and g12549 ( n21437 , n12657 , n10092 );
    or g12550 ( n16014 , n10124 , n18734 );
    nor g12551 ( n15066 , n26093 , n5745 );
    and g12552 ( n12285 , n24594 , n15912 );
    and g12553 ( n5641 , n20489 , n21693 );
    and g12554 ( n10512 , n12962 , n26662 );
    or g12555 ( n10526 , n26790 , n13366 );
    nor g12556 ( n12526 , n1299 , n19411 );
    and g12557 ( n3021 , n21102 , n8005 );
    nor g12558 ( n14627 , n16294 , n12507 );
    nor g12559 ( n25369 , n15580 , n9050 );
    and g12560 ( n9437 , n5249 , n9516 );
    xnor g12561 ( n9556 , n15688 , n11169 );
    or g12562 ( n4946 , n25639 , n12648 );
    or g12563 ( n9585 , n4582 , n19993 );
    and g12564 ( n10344 , n18186 , n1664 );
    xnor g12565 ( n6279 , n12382 , n26754 );
    and g12566 ( n19154 , n14726 , n18695 );
    or g12567 ( n1968 , n27188 , n8890 );
    nor g12568 ( n6484 , n2585 , n7179 );
    or g12569 ( n16950 , n1775 , n21170 );
    xnor g12570 ( n1539 , n11159 , n9477 );
    not g12571 ( n13376 , n26191 );
    xnor g12572 ( n1482 , n7935 , n11552 );
    not g12573 ( n4400 , n18500 );
    or g12574 ( n11183 , n23304 , n17069 );
    xnor g12575 ( n3082 , n18806 , n24136 );
    nor g12576 ( n2380 , n3257 , n3677 );
    nor g12577 ( n25507 , n19327 , n21934 );
    not g12578 ( n24658 , n21473 );
    or g12579 ( n7848 , n5277 , n19123 );
    not g12580 ( n11257 , n10631 );
    xnor g12581 ( n17493 , n23147 , n6536 );
    nor g12582 ( n6581 , n16257 , n4119 );
    not g12583 ( n16709 , n15291 );
    xnor g12584 ( n2365 , n24786 , n20036 );
    and g12585 ( n2575 , n16622 , n23946 );
    nor g12586 ( n25596 , n557 , n16006 );
    or g12587 ( n5971 , n586 , n21825 );
    or g12588 ( n6694 , n7661 , n459 );
    xnor g12589 ( n11029 , n14323 , n14071 );
    xnor g12590 ( n7338 , n20230 , n18034 );
    xnor g12591 ( n5969 , n23212 , n2728 );
    and g12592 ( n7156 , n2341 , n2503 );
    not g12593 ( n21734 , n25568 );
    or g12594 ( n17783 , n23055 , n3696 );
    xnor g12595 ( n12291 , n26635 , n12399 );
    and g12596 ( n16152 , n8672 , n5296 );
    xnor g12597 ( n3208 , n23902 , n7132 );
    and g12598 ( n25848 , n17357 , n20419 );
    xnor g12599 ( n14047 , n9110 , n13282 );
    and g12600 ( n10922 , n12520 , n26933 );
    not g12601 ( n9693 , n15062 );
    not g12602 ( n14151 , n8418 );
    nor g12603 ( n2144 , n17370 , n11061 );
    or g12604 ( n19133 , n14133 , n4024 );
    not g12605 ( n5328 , n12169 );
    not g12606 ( n506 , n24326 );
    xnor g12607 ( n23950 , n3887 , n327 );
    xnor g12608 ( n12297 , n8336 , n2985 );
    or g12609 ( n23821 , n20446 , n24606 );
    xnor g12610 ( n17455 , n2812 , n5736 );
    xnor g12611 ( n15437 , n26360 , n110 );
    xnor g12612 ( n12145 , n2256 , n20694 );
    or g12613 ( n24769 , n16002 , n3945 );
    or g12614 ( n25453 , n2846 , n23087 );
    not g12615 ( n22715 , n16324 );
    nor g12616 ( n12189 , n21247 , n17390 );
    and g12617 ( n19226 , n3958 , n10746 );
    and g12618 ( n17318 , n17834 , n22663 );
    xnor g12619 ( n21912 , n1286 , n15645 );
    not g12620 ( n9969 , n19940 );
    or g12621 ( n14370 , n13131 , n5528 );
    nor g12622 ( n23976 , n13037 , n13129 );
    nor g12623 ( n12303 , n25119 , n21934 );
    or g12624 ( n632 , n19267 , n4177 );
    and g12625 ( n1543 , n21241 , n10060 );
    or g12626 ( n10162 , n7051 , n6749 );
    or g12627 ( n19766 , n15517 , n8120 );
    and g12628 ( n10542 , n5802 , n19368 );
    not g12629 ( n19605 , n10884 );
    nor g12630 ( n25342 , n19673 , n5462 );
    or g12631 ( n15559 , n26451 , n26155 );
    or g12632 ( n7852 , n13162 , n23346 );
    xnor g12633 ( n14762 , n15431 , n25310 );
    and g12634 ( n16452 , n26224 , n8672 );
    xnor g12635 ( n15342 , n22654 , n21915 );
    xnor g12636 ( n11132 , n3808 , n923 );
    or g12637 ( n2714 , n10078 , n4373 );
    xnor g12638 ( n11354 , n26324 , n12262 );
    or g12639 ( n7044 , n11324 , n20168 );
    xor g12640 ( n2288 , n4304 , n21114 );
    xnor g12641 ( n22463 , n27118 , n7678 );
    and g12642 ( n13657 , n22879 , n12616 );
    or g12643 ( n26436 , n21489 , n4085 );
    xnor g12644 ( n498 , n20296 , n17338 );
    nor g12645 ( n10259 , n12046 , n6072 );
    or g12646 ( n11612 , n1509 , n16913 );
    xnor g12647 ( n15014 , n5140 , n6105 );
    xnor g12648 ( n14298 , n11305 , n3001 );
    or g12649 ( n11943 , n15983 , n23117 );
    xnor g12650 ( n3781 , n6969 , n22339 );
    and g12651 ( n7415 , n7844 , n9541 );
    xnor g12652 ( n1512 , n15288 , n12361 );
    not g12653 ( n5760 , n8151 );
    and g12654 ( n843 , n20373 , n1375 );
    or g12655 ( n21312 , n8322 , n19081 );
    nor g12656 ( n26878 , n24116 , n11580 );
    xnor g12657 ( n16126 , n16234 , n4673 );
    and g12658 ( n23468 , n2396 , n432 );
    xnor g12659 ( n23955 , n23290 , n10709 );
    xnor g12660 ( n18883 , n15652 , n4939 );
    or g12661 ( n18128 , n19375 , n9278 );
    xnor g12662 ( n24608 , n4750 , n7859 );
    or g12663 ( n17097 , n23359 , n11898 );
    xnor g12664 ( n2305 , n4941 , n9780 );
    and g12665 ( n46 , n8561 , n4470 );
    or g12666 ( n2635 , n10366 , n16814 );
    or g12667 ( n19292 , n11429 , n12969 );
    nor g12668 ( n16767 , n10773 , n22470 );
    or g12669 ( n4048 , n21686 , n17191 );
    xnor g12670 ( n16233 , n8596 , n15508 );
    and g12671 ( n8969 , n12264 , n27137 );
    or g12672 ( n15750 , n10044 , n24999 );
    nor g12673 ( n20809 , n25953 , n24460 );
    xnor g12674 ( n1223 , n24043 , n10201 );
    and g12675 ( n8265 , n2421 , n11243 );
    or g12676 ( n15634 , n24555 , n5985 );
    nor g12677 ( n4582 , n16988 , n20442 );
    xnor g12678 ( n14960 , n13492 , n23763 );
    xnor g12679 ( n7824 , n10667 , n19636 );
    xnor g12680 ( n1821 , n10477 , n6548 );
    xnor g12681 ( n24136 , n13854 , n18503 );
    nor g12682 ( n25024 , n21547 , n6003 );
    and g12683 ( n11068 , n6482 , n8710 );
    or g12684 ( n14191 , n17065 , n11124 );
    nor g12685 ( n12712 , n10053 , n5329 );
    or g12686 ( n23682 , n6833 , n24615 );
    xnor g12687 ( n6088 , n15572 , n2989 );
    and g12688 ( n4102 , n11089 , n972 );
    not g12689 ( n16731 , n13284 );
    nor g12690 ( n25553 , n12900 , n1255 );
    or g12691 ( n2936 , n5244 , n16373 );
    not g12692 ( n12055 , n24714 );
    xnor g12693 ( n2367 , n1308 , n7734 );
    nor g12694 ( n3531 , n4075 , n12120 );
    or g12695 ( n7766 , n1742 , n14251 );
    or g12696 ( n3221 , n12305 , n24817 );
    xnor g12697 ( n5496 , n24519 , n12161 );
    and g12698 ( n3028 , n24792 , n18299 );
    or g12699 ( n26381 , n25940 , n22325 );
    or g12700 ( n15110 , n27071 , n18595 );
    or g12701 ( n8673 , n19949 , n11136 );
    not g12702 ( n17790 , n17311 );
    nor g12703 ( n17814 , n4304 , n19413 );
    xnor g12704 ( n1162 , n12103 , n9448 );
    or g12705 ( n2447 , n12914 , n6846 );
    or g12706 ( n16414 , n24414 , n22434 );
    xnor g12707 ( n11182 , n11977 , n10059 );
    or g12708 ( n994 , n7094 , n21163 );
    xnor g12709 ( n6283 , n15730 , n2331 );
    not g12710 ( n15514 , n19431 );
    nor g12711 ( n7778 , n1279 , n14875 );
    xnor g12712 ( n20288 , n9711 , n19064 );
    xnor g12713 ( n19303 , n18913 , n15352 );
    nor g12714 ( n10492 , n1594 , n16602 );
    nor g12715 ( n23968 , n16781 , n15777 );
    and g12716 ( n25708 , n22430 , n9676 );
    xnor g12717 ( n12188 , n23779 , n11615 );
    not g12718 ( n393 , n1924 );
    nor g12719 ( n6870 , n15743 , n2809 );
    or g12720 ( n4903 , n9296 , n25915 );
    xnor g12721 ( n4885 , n17390 , n22736 );
    or g12722 ( n26908 , n21937 , n25355 );
    or g12723 ( n12069 , n7716 , n22654 );
    xnor g12724 ( n15956 , n3209 , n9306 );
    and g12725 ( n615 , n26222 , n12565 );
    not g12726 ( n11697 , n15108 );
    nor g12727 ( n20750 , n10557 , n18113 );
    xnor g12728 ( n14731 , n22861 , n4426 );
    xnor g12729 ( n7272 , n20620 , n14575 );
    nor g12730 ( n8579 , n14996 , n10357 );
    not g12731 ( n13821 , n6483 );
    xnor g12732 ( n14044 , n13731 , n13714 );
    not g12733 ( n15259 , n16705 );
    nor g12734 ( n4650 , n19842 , n7258 );
    or g12735 ( n5340 , n3228 , n20189 );
    or g12736 ( n23483 , n649 , n26065 );
    xnor g12737 ( n4502 , n25718 , n4634 );
    and g12738 ( n15988 , n21395 , n10856 );
    nor g12739 ( n17129 , n16751 , n25018 );
    buf g12740 ( n5914 , n8280 );
    not g12741 ( n24366 , n1152 );
    xnor g12742 ( n6423 , n21471 , n19357 );
    xnor g12743 ( n8767 , n9399 , n9507 );
    and g12744 ( n10668 , n11976 , n11437 );
    xnor g12745 ( n1618 , n22354 , n5744 );
    and g12746 ( n6811 , n11485 , n11582 );
    xnor g12747 ( n6912 , n18881 , n25016 );
    or g12748 ( n3268 , n26797 , n16221 );
    not g12749 ( n10904 , n13262 );
    xnor g12750 ( n16040 , n17184 , n18587 );
    or g12751 ( n10805 , n6239 , n8319 );
    not g12752 ( n12066 , n20013 );
    xnor g12753 ( n14541 , n15650 , n15691 );
    not g12754 ( n544 , n9359 );
    xnor g12755 ( n345 , n6908 , n26972 );
    and g12756 ( n3287 , n2241 , n16418 );
    or g12757 ( n11362 , n26122 , n26306 );
    and g12758 ( n19249 , n4698 , n14623 );
    not g12759 ( n16642 , n3217 );
    and g12760 ( n4276 , n19746 , n22693 );
    xnor g12761 ( n13798 , n10471 , n13403 );
    not g12762 ( n15049 , n19039 );
    xnor g12763 ( n16142 , n24661 , n15462 );
    nor g12764 ( n7155 , n8708 , n9402 );
    nor g12765 ( n12965 , n19460 , n16064 );
    and g12766 ( n9320 , n13861 , n4021 );
    and g12767 ( n5676 , n25206 , n10502 );
    or g12768 ( n6720 , n7099 , n18888 );
    nor g12769 ( n7880 , n23039 , n4590 );
    or g12770 ( n13662 , n2314 , n25643 );
    nor g12771 ( n11881 , n24557 , n15630 );
    xnor g12772 ( n3713 , n1082 , n10277 );
    or g12773 ( n19185 , n9351 , n16360 );
    and g12774 ( n1500 , n7822 , n24543 );
    not g12775 ( n5886 , n10024 );
    xnor g12776 ( n4811 , n16075 , n9370 );
    nor g12777 ( n24765 , n776 , n13494 );
    or g12778 ( n22996 , n21078 , n13725 );
    or g12779 ( n11954 , n12140 , n8791 );
    xnor g12780 ( n6875 , n17333 , n14783 );
    or g12781 ( n8633 , n9493 , n12297 );
    or g12782 ( n169 , n16853 , n8768 );
    xnor g12783 ( n24015 , n11061 , n1971 );
    xnor g12784 ( n7049 , n21882 , n26694 );
    or g12785 ( n9837 , n844 , n3103 );
    xnor g12786 ( n21487 , n23262 , n12931 );
    or g12787 ( n25522 , n14052 , n18925 );
    nor g12788 ( n2329 , n23582 , n16738 );
    xnor g12789 ( n8170 , n19159 , n23399 );
    or g12790 ( n22461 , n18581 , n12567 );
    or g12791 ( n25272 , n11996 , n7430 );
    or g12792 ( n13970 , n25408 , n15781 );
    and g12793 ( n6073 , n5395 , n11991 );
    not g12794 ( n5512 , n12315 );
    or g12795 ( n315 , n17978 , n3134 );
    and g12796 ( n9791 , n1792 , n19521 );
    and g12797 ( n10173 , n7461 , n26464 );
    xnor g12798 ( n20068 , n10602 , n22395 );
    xnor g12799 ( n26992 , n22142 , n26081 );
    xnor g12800 ( n24461 , n25980 , n15182 );
    and g12801 ( n20769 , n3453 , n6487 );
    and g12802 ( n14316 , n1341 , n7821 );
    xnor g12803 ( n12518 , n2312 , n10378 );
    and g12804 ( n17567 , n13078 , n19183 );
    and g12805 ( n12914 , n21101 , n17779 );
    or g12806 ( n25478 , n2482 , n19104 );
    xnor g12807 ( n10135 , n15490 , n18 );
    xnor g12808 ( n20210 , n6489 , n16743 );
    xnor g12809 ( n20231 , n6049 , n23816 );
    and g12810 ( n16897 , n4392 , n14834 );
    xnor g12811 ( n27135 , n18742 , n14319 );
    xnor g12812 ( n12169 , n5816 , n5438 );
    and g12813 ( n9379 , n15571 , n16838 );
    xnor g12814 ( n3465 , n2843 , n25232 );
    xnor g12815 ( n26234 , n7963 , n6590 );
    nor g12816 ( n8802 , n6523 , n24479 );
    and g12817 ( n26052 , n10333 , n2100 );
    not g12818 ( n27099 , n24444 );
    or g12819 ( n8193 , n11862 , n23070 );
    xnor g12820 ( n2611 , n17607 , n23366 );
    nor g12821 ( n12641 , n26991 , n23330 );
    xnor g12822 ( n17337 , n24895 , n21970 );
    xnor g12823 ( n20293 , n6937 , n17843 );
    or g12824 ( n22258 , n7165 , n23239 );
    xnor g12825 ( n23268 , n9895 , n15537 );
    not g12826 ( n2724 , n14275 );
    and g12827 ( n24787 , n6958 , n2912 );
    or g12828 ( n10134 , n14619 , n26251 );
    and g12829 ( n16450 , n14566 , n11895 );
    not g12830 ( n7410 , n11454 );
    nor g12831 ( n19398 , n8119 , n26135 );
    xnor g12832 ( n24828 , n5679 , n20839 );
    and g12833 ( n15665 , n17630 , n18557 );
    xnor g12834 ( n10866 , n17250 , n11044 );
    not g12835 ( n12112 , n21620 );
    and g12836 ( n17654 , n11834 , n5788 );
    not g12837 ( n24590 , n6492 );
    xnor g12838 ( n19858 , n16271 , n3117 );
    or g12839 ( n495 , n8981 , n22593 );
    not g12840 ( n4029 , n2530 );
    and g12841 ( n4 , n2159 , n5056 );
    and g12842 ( n23256 , n17707 , n27133 );
    xnor g12843 ( n4260 , n17250 , n15241 );
    xnor g12844 ( n4477 , n17517 , n23099 );
    not g12845 ( n18621 , n5034 );
    nor g12846 ( n751 , n5031 , n6510 );
    and g12847 ( n18804 , n11972 , n19507 );
    or g12848 ( n17281 , n25671 , n17040 );
    nor g12849 ( n16952 , n25365 , n15456 );
    and g12850 ( n11050 , n21992 , n13289 );
    or g12851 ( n23838 , n5410 , n8358 );
    and g12852 ( n19123 , n16341 , n11218 );
    xnor g12853 ( n1741 , n8720 , n3803 );
    xnor g12854 ( n9146 , n15310 , n5844 );
    not g12855 ( n11921 , n23216 );
    nor g12856 ( n9297 , n26170 , n23664 );
    or g12857 ( n1585 , n21821 , n25530 );
    and g12858 ( n2040 , n22851 , n5988 );
    not g12859 ( n508 , n14199 );
    xnor g12860 ( n8958 , n3704 , n9021 );
    xnor g12861 ( n12905 , n23704 , n2659 );
    or g12862 ( n19917 , n20814 , n22936 );
    or g12863 ( n13675 , n12567 , n12279 );
    not g12864 ( n5433 , n16411 );
    not g12865 ( n6948 , n477 );
    or g12866 ( n18900 , n27199 , n12964 );
    or g12867 ( n7730 , n26634 , n7314 );
    xnor g12868 ( n14015 , n6895 , n20462 );
    xnor g12869 ( n2038 , n26190 , n12355 );
    xnor g12870 ( n16397 , n11533 , n14398 );
    xnor g12871 ( n25045 , n3136 , n5752 );
    nor g12872 ( n17407 , n24656 , n13583 );
    and g12873 ( n11586 , n19568 , n162 );
    nor g12874 ( n12030 , n27053 , n12544 );
    and g12875 ( n11340 , n18709 , n27016 );
    and g12876 ( n9347 , n212 , n9928 );
    not g12877 ( n12971 , n2608 );
    and g12878 ( n26296 , n14510 , n8994 );
    xnor g12879 ( n19402 , n2036 , n2891 );
    or g12880 ( n6651 , n23537 , n11010 );
    not g12881 ( n13822 , n22793 );
    and g12882 ( n6761 , n17319 , n9511 );
    or g12883 ( n6735 , n25650 , n5077 );
    not g12884 ( n23315 , n6387 );
    and g12885 ( n17571 , n11966 , n6722 );
    or g12886 ( n15416 , n15576 , n21739 );
    and g12887 ( n17561 , n8690 , n9363 );
    and g12888 ( n20499 , n23949 , n17093 );
    not g12889 ( n13343 , n6372 );
    or g12890 ( n12056 , n5918 , n2944 );
    or g12891 ( n16297 , n7632 , n14384 );
    xnor g12892 ( n17117 , n8083 , n18705 );
    not g12893 ( n4116 , n25995 );
    or g12894 ( n2644 , n7146 , n3549 );
    xnor g12895 ( n5786 , n17959 , n6861 );
    or g12896 ( n20473 , n22256 , n16220 );
    not g12897 ( n13280 , n3480 );
    or g12898 ( n22486 , n1831 , n10022 );
    and g12899 ( n1210 , n11700 , n13398 );
    xnor g12900 ( n5096 , n23709 , n19282 );
    nor g12901 ( n11854 , n12464 , n18907 );
    and g12902 ( n20185 , n21597 , n22722 );
    nor g12903 ( n24314 , n1432 , n2852 );
    not g12904 ( n25787 , n17694 );
    and g12905 ( n14945 , n14128 , n2256 );
    and g12906 ( n19885 , n23774 , n24751 );
    or g12907 ( n17179 , n26191 , n13284 );
    and g12908 ( n26622 , n16402 , n24944 );
    and g12909 ( n6140 , n22439 , n26235 );
    xnor g12910 ( n3628 , n13539 , n20973 );
    and g12911 ( n5362 , n7951 , n15443 );
    xnor g12912 ( n18139 , n6208 , n10177 );
    not g12913 ( n21400 , n13963 );
    not g12914 ( n2314 , n329 );
    nor g12915 ( n18305 , n8428 , n25961 );
    or g12916 ( n5015 , n21856 , n24163 );
    xnor g12917 ( n6829 , n1118 , n10053 );
    or g12918 ( n3647 , n4686 , n21836 );
    or g12919 ( n1948 , n34 , n13625 );
    xnor g12920 ( n8482 , n24488 , n23250 );
    xnor g12921 ( n22857 , n3346 , n8044 );
    and g12922 ( n21401 , n19129 , n20855 );
    not g12923 ( n10105 , n12419 );
    nor g12924 ( n23943 , n23798 , n12217 );
    and g12925 ( n25620 , n5101 , n17423 );
    or g12926 ( n26606 , n10156 , n12416 );
    not g12927 ( n14119 , n6590 );
    or g12928 ( n16613 , n11580 , n2035 );
    xnor g12929 ( n5978 , n22640 , n7566 );
    nor g12930 ( n22185 , n1209 , n13599 );
    nor g12931 ( n68 , n6731 , n7347 );
    or g12932 ( n17801 , n23315 , n14463 );
    not g12933 ( n9340 , n15458 );
    xnor g12934 ( n19393 , n3732 , n23196 );
    and g12935 ( n4069 , n2631 , n7559 );
    nor g12936 ( n17065 , n20151 , n5852 );
    xnor g12937 ( n22704 , n7407 , n9625 );
    or g12938 ( n7412 , n1259 , n44 );
    xnor g12939 ( n665 , n12077 , n3596 );
    not g12940 ( n25566 , n18213 );
    or g12941 ( n26563 , n8895 , n13727 );
    or g12942 ( n26755 , n10273 , n24648 );
    xnor g12943 ( n3559 , n27188 , n4326 );
    xnor g12944 ( n2819 , n12771 , n5025 );
    or g12945 ( n17894 , n2877 , n20457 );
    xnor g12946 ( n18108 , n16070 , n20008 );
    not g12947 ( n6841 , n7330 );
    xnor g12948 ( n17598 , n12677 , n10974 );
    not g12949 ( n23114 , n10751 );
    xnor g12950 ( n11005 , n19407 , n25398 );
    not g12951 ( n22397 , n14057 );
    or g12952 ( n16632 , n14401 , n26306 );
    and g12953 ( n14914 , n8200 , n21192 );
    or g12954 ( n15084 , n23477 , n1365 );
    or g12955 ( n21227 , n12702 , n13672 );
    and g12956 ( n10879 , n3775 , n23221 );
    not g12957 ( n23725 , n11933 );
    or g12958 ( n238 , n2445 , n7511 );
    nor g12959 ( n6869 , n13957 , n13343 );
    nor g12960 ( n21475 , n27120 , n23264 );
    and g12961 ( n5550 , n12578 , n16671 );
    and g12962 ( n611 , n23396 , n17790 );
    and g12963 ( n23997 , n6464 , n7351 );
    and g12964 ( n21931 , n5345 , n17363 );
    nor g12965 ( n26478 , n12258 , n14774 );
    not g12966 ( n7331 , n6038 );
    and g12967 ( n23390 , n22198 , n24493 );
    xnor g12968 ( n6237 , n5465 , n17505 );
    xnor g12969 ( n14971 , n1765 , n25119 );
    nor g12970 ( n17032 , n20845 , n26848 );
    nor g12971 ( n12458 , n5288 , n24923 );
    or g12972 ( n8468 , n16034 , n10451 );
    or g12973 ( n15595 , n25021 , n26495 );
    xnor g12974 ( n23958 , n22098 , n7174 );
    or g12975 ( n1010 , n16767 , n23606 );
    not g12976 ( n21814 , n4062 );
    xnor g12977 ( n20025 , n25974 , n19005 );
    or g12978 ( n10328 , n3970 , n4059 );
    xnor g12979 ( n25113 , n3572 , n3148 );
    xnor g12980 ( n3638 , n21652 , n5225 );
    not g12981 ( n2169 , n19531 );
    and g12982 ( n14379 , n13601 , n20540 );
    xnor g12983 ( n6172 , n19875 , n9737 );
    xnor g12984 ( n17585 , n20794 , n25471 );
    nor g12985 ( n21281 , n12343 , n14106 );
    not g12986 ( n11840 , n323 );
    not g12987 ( n17010 , n17530 );
    xnor g12988 ( n2201 , n1112 , n7751 );
    and g12989 ( n23427 , n20536 , n2749 );
    xnor g12990 ( n1057 , n2093 , n22173 );
    xnor g12991 ( n24344 , n2924 , n13669 );
    or g12992 ( n828 , n4967 , n18559 );
    not g12993 ( n24731 , n6135 );
    xnor g12994 ( n4086 , n14210 , n21078 );
    or g12995 ( n2053 , n25791 , n15088 );
    not g12996 ( n17584 , n26986 );
    xnor g12997 ( n16520 , n8443 , n5170 );
    or g12998 ( n13458 , n11179 , n6668 );
    or g12999 ( n8575 , n7827 , n23203 );
    and g13000 ( n20534 , n20798 , n9878 );
    xnor g13001 ( n7089 , n10937 , n16376 );
    or g13002 ( n18150 , n21260 , n24121 );
    or g13003 ( n130 , n13800 , n25766 );
    nor g13004 ( n4686 , n25751 , n21850 );
    xnor g13005 ( n19896 , n3393 , n1465 );
    xnor g13006 ( n4345 , n13502 , n21055 );
    xnor g13007 ( n2507 , n14148 , n14275 );
    not g13008 ( n8395 , n14102 );
    nor g13009 ( n18912 , n9877 , n23464 );
    and g13010 ( n21657 , n23584 , n26020 );
    xnor g13011 ( n10408 , n23740 , n2858 );
    and g13012 ( n25853 , n11859 , n15770 );
    xnor g13013 ( n2440 , n5656 , n21005 );
    not g13014 ( n20982 , n12696 );
    xnor g13015 ( n17138 , n15849 , n7278 );
    or g13016 ( n22752 , n2842 , n20933 );
    or g13017 ( n1463 , n19469 , n13989 );
    or g13018 ( n13180 , n16221 , n21444 );
    or g13019 ( n21139 , n25588 , n25613 );
    xnor g13020 ( n24425 , n18983 , n4487 );
    or g13021 ( n2682 , n21380 , n15659 );
    or g13022 ( n20166 , n20589 , n26021 );
    xnor g13023 ( n26693 , n14633 , n2886 );
    and g13024 ( n24587 , n6996 , n8570 );
    or g13025 ( n3982 , n2230 , n19227 );
    and g13026 ( n1263 , n17077 , n14620 );
    or g13027 ( n5577 , n24607 , n7903 );
    or g13028 ( n20701 , n19541 , n25749 );
    and g13029 ( n3338 , n5141 , n24637 );
    xnor g13030 ( n10974 , n19042 , n23586 );
    nor g13031 ( n20801 , n26450 , n17351 );
    xnor g13032 ( n26285 , n8163 , n2688 );
    not g13033 ( n10155 , n18171 );
    not g13034 ( n22600 , n25115 );
    or g13035 ( n11290 , n15044 , n12377 );
    xnor g13036 ( n26216 , n4985 , n11242 );
    nor g13037 ( n2332 , n8003 , n22972 );
    or g13038 ( n23356 , n6871 , n18328 );
    xnor g13039 ( n26943 , n25732 , n11565 );
    xnor g13040 ( n23960 , n11337 , n11893 );
    or g13041 ( n18722 , n21280 , n7002 );
    or g13042 ( n8060 , n14778 , n13510 );
    or g13043 ( n26578 , n20978 , n25243 );
    and g13044 ( n8207 , n9147 , n24597 );
    and g13045 ( n26360 , n20504 , n14896 );
    or g13046 ( n23662 , n21879 , n8853 );
    and g13047 ( n19754 , n21956 , n17700 );
    and g13048 ( n21375 , n24461 , n26095 );
    nor g13049 ( n16347 , n9107 , n18360 );
    not g13050 ( n5826 , n6265 );
    nor g13051 ( n19083 , n839 , n6139 );
    xnor g13052 ( n18137 , n13219 , n19376 );
    xnor g13053 ( n3799 , n7242 , n880 );
    or g13054 ( n18185 , n26069 , n23277 );
    and g13055 ( n24808 , n8435 , n9580 );
    and g13056 ( n15398 , n20076 , n4970 );
    not g13057 ( n1387 , n10699 );
    not g13058 ( n15229 , n20014 );
    nor g13059 ( n22886 , n20127 , n19927 );
    or g13060 ( n9070 , n4149 , n12875 );
    not g13061 ( n12018 , n11671 );
    xnor g13062 ( n15835 , n3045 , n9376 );
    nor g13063 ( n20184 , n4326 , n3952 );
    or g13064 ( n2571 , n7124 , n16510 );
    xnor g13065 ( n7698 , n14729 , n1976 );
    or g13066 ( n10921 , n438 , n18784 );
    or g13067 ( n9580 , n3422 , n22525 );
    nor g13068 ( n12196 , n24237 , n4017 );
    and g13069 ( n19095 , n5329 , n2694 );
    xnor g13070 ( n10846 , n16882 , n3976 );
    or g13071 ( n21688 , n25068 , n23535 );
    or g13072 ( n7440 , n6869 , n1159 );
    or g13073 ( n20818 , n26092 , n24930 );
    or g13074 ( n16067 , n7759 , n10479 );
    xnor g13075 ( n7988 , n22772 , n8930 );
    or g13076 ( n6839 , n17856 , n18790 );
    not g13077 ( n20433 , n17824 );
    xnor g13078 ( n26942 , n24308 , n13075 );
    and g13079 ( n5781 , n2058 , n10112 );
    or g13080 ( n15037 , n15154 , n19445 );
    and g13081 ( n8643 , n17371 , n4695 );
    not g13082 ( n8647 , n271 );
    xnor g13083 ( n26675 , n5370 , n9685 );
    nor g13084 ( n2084 , n23913 , n3710 );
    not g13085 ( n21485 , n15190 );
    and g13086 ( n3709 , n18994 , n7787 );
    not g13087 ( n18269 , n10057 );
    not g13088 ( n4859 , n10250 );
    xnor g13089 ( n15828 , n19701 , n7437 );
    and g13090 ( n18440 , n7602 , n4475 );
    nor g13091 ( n13163 , n905 , n4706 );
    nor g13092 ( n17378 , n6270 , n27121 );
    or g13093 ( n19344 , n24890 , n4665 );
    xnor g13094 ( n15716 , n720 , n6888 );
    xnor g13095 ( n18509 , n5459 , n6467 );
    not g13096 ( n19926 , n23776 );
    xnor g13097 ( n12361 , n18255 , n15636 );
    or g13098 ( n16055 , n7161 , n16411 );
    and g13099 ( n2286 , n8921 , n26734 );
    not g13100 ( n6200 , n4184 );
    or g13101 ( n9030 , n11980 , n19446 );
    or g13102 ( n25448 , n8021 , n25309 );
    or g13103 ( n6844 , n21613 , n8974 );
    and g13104 ( n16021 , n18244 , n4107 );
    not g13105 ( n9373 , n24928 );
    nor g13106 ( n14492 , n10758 , n13562 );
    not g13107 ( n22862 , n11295 );
    or g13108 ( n2835 , n23428 , n8649 );
    xnor g13109 ( n20519 , n13945 , n12341 );
    or g13110 ( n22384 , n18114 , n1 );
    or g13111 ( n15690 , n18761 , n5665 );
    xnor g13112 ( n19708 , n8006 , n5211 );
    xnor g13113 ( n9992 , n13891 , n11140 );
    or g13114 ( n13316 , n1414 , n4005 );
    and g13115 ( n18703 , n2789 , n13640 );
    or g13116 ( n5502 , n22318 , n1162 );
    and g13117 ( n3486 , n375 , n25771 );
    and g13118 ( n5086 , n22299 , n13294 );
    or g13119 ( n174 , n22737 , n3767 );
    xnor g13120 ( n23585 , n3467 , n19456 );
    xnor g13121 ( n11538 , n156 , n22058 );
    xnor g13122 ( n5818 , n212 , n17150 );
    or g13123 ( n14574 , n21777 , n15392 );
    xnor g13124 ( n18010 , n4230 , n8378 );
    not g13125 ( n14158 , n24219 );
    or g13126 ( n26753 , n12505 , n24497 );
    xnor g13127 ( n2389 , n24436 , n21885 );
    and g13128 ( n20926 , n7577 , n15731 );
    or g13129 ( n14987 , n24540 , n14901 );
    xnor g13130 ( n5142 , n974 , n18668 );
    xnor g13131 ( n15328 , n22972 , n3945 );
    xnor g13132 ( n5556 , n7787 , n23722 );
    xnor g13133 ( n13958 , n7014 , n13611 );
    xnor g13134 ( n21212 , n24902 , n25572 );
    not g13135 ( n9212 , n16814 );
    and g13136 ( n4709 , n6204 , n23898 );
    or g13137 ( n19434 , n25823 , n2018 );
    and g13138 ( n1430 , n24532 , n18021 );
    and g13139 ( n25541 , n19699 , n24526 );
    and g13140 ( n3433 , n12787 , n2016 );
    and g13141 ( n16318 , n25776 , n628 );
    xnor g13142 ( n19404 , n15924 , n2680 );
    or g13143 ( n1795 , n19061 , n13436 );
    or g13144 ( n16676 , n9471 , n6589 );
    or g13145 ( n15627 , n17251 , n23967 );
    xnor g13146 ( n2827 , n23631 , n22765 );
    xnor g13147 ( n7630 , n25995 , n21115 );
    xnor g13148 ( n22581 , n12734 , n631 );
    xnor g13149 ( n26282 , n8722 , n13119 );
    and g13150 ( n1145 , n1932 , n14526 );
    not g13151 ( n12996 , n18145 );
    xnor g13152 ( n8283 , n7805 , n7657 );
    and g13153 ( n15763 , n7089 , n16793 );
    xnor g13154 ( n22953 , n18614 , n19420 );
    or g13155 ( n24683 , n331 , n684 );
    xnor g13156 ( n7045 , n9655 , n13074 );
    xnor g13157 ( n20415 , n11883 , n14064 );
    and g13158 ( n16549 , n3676 , n9224 );
    not g13159 ( n15454 , n9554 );
    and g13160 ( n11160 , n9070 , n10842 );
    and g13161 ( n18593 , n2085 , n5169 );
    xnor g13162 ( n9937 , n6319 , n442 );
    xnor g13163 ( n21252 , n17734 , n23253 );
    xnor g13164 ( n13266 , n9535 , n2615 );
    or g13165 ( n10518 , n23808 , n20887 );
    xnor g13166 ( n22776 , n9993 , n25926 );
    xnor g13167 ( n19446 , n19545 , n25749 );
    nor g13168 ( n11622 , n8371 , n4410 );
    xnor g13169 ( n10489 , n11396 , n14797 );
    xnor g13170 ( n3426 , n11693 , n13375 );
    or g13171 ( n19031 , n9913 , n20428 );
    nor g13172 ( n2637 , n11363 , n14119 );
    or g13173 ( n5271 , n5355 , n17659 );
    xnor g13174 ( n22687 , n9333 , n14666 );
    not g13175 ( n19884 , n8635 );
    nor g13176 ( n12282 , n25974 , n2355 );
    xnor g13177 ( n21399 , n23421 , n10846 );
    or g13178 ( n18839 , n9262 , n16934 );
    or g13179 ( n19981 , n4256 , n5713 );
    and g13180 ( n9262 , n11089 , n4955 );
    nor g13181 ( n16085 , n25324 , n1630 );
    or g13182 ( n9037 , n26782 , n20089 );
    xor g13183 ( n915 , n7325 , n15232 );
    not g13184 ( n20737 , n15167 );
    xnor g13185 ( n9989 , n10218 , n19547 );
    xnor g13186 ( n21970 , n20771 , n18639 );
    or g13187 ( n20501 , n5304 , n13115 );
    xnor g13188 ( n5805 , n3785 , n21 );
    xnor g13189 ( n15039 , n18295 , n16223 );
    xnor g13190 ( n18577 , n11499 , n18570 );
    and g13191 ( n19860 , n21360 , n2311 );
    xnor g13192 ( n6655 , n13067 , n25735 );
    xor g13193 ( n25416 , n7991 , n13323 );
    and g13194 ( n22305 , n24737 , n25767 );
    or g13195 ( n10865 , n176 , n1452 );
    or g13196 ( n25878 , n5836 , n17788 );
    xnor g13197 ( n24141 , n5909 , n15401 );
    and g13198 ( n23066 , n22011 , n17042 );
    or g13199 ( n2921 , n6533 , n24685 );
    not g13200 ( n4658 , n4869 );
    or g13201 ( n1379 , n18274 , n24383 );
    not g13202 ( n23793 , n15508 );
    xnor g13203 ( n13151 , n9717 , n407 );
    and g13204 ( n12045 , n15699 , n25732 );
    and g13205 ( n15335 , n10292 , n20559 );
    or g13206 ( n26097 , n12471 , n23533 );
    xnor g13207 ( n11671 , n7415 , n8242 );
    and g13208 ( n17241 , n21892 , n20779 );
    or g13209 ( n5906 , n23304 , n1465 );
    not g13210 ( n25779 , n3078 );
    xnor g13211 ( n2573 , n13806 , n20351 );
    or g13212 ( n22611 , n23830 , n19342 );
    xnor g13213 ( n25813 , n24075 , n20941 );
    not g13214 ( n147 , n11721 );
    xnor g13215 ( n10660 , n22951 , n14561 );
    or g13216 ( n11037 , n7705 , n19016 );
    xnor g13217 ( n18875 , n16500 , n8678 );
    xnor g13218 ( n804 , n20051 , n18434 );
    not g13219 ( n23302 , n18265 );
    or g13220 ( n15360 , n19632 , n6085 );
    xnor g13221 ( n5325 , n20116 , n12054 );
    or g13222 ( n9642 , n12562 , n12351 );
    and g13223 ( n14803 , n15135 , n25712 );
    nor g13224 ( n2340 , n26443 , n10017 );
    and g13225 ( n10991 , n19954 , n9596 );
    xnor g13226 ( n21082 , n21345 , n9190 );
    or g13227 ( n20653 , n4834 , n23823 );
    or g13228 ( n19876 , n17090 , n6773 );
    and g13229 ( n13169 , n5704 , n5512 );
    not g13230 ( n15007 , n4513 );
    and g13231 ( n7239 , n12434 , n11681 );
    xnor g13232 ( n9616 , n17146 , n4004 );
    xnor g13233 ( n16798 , n12332 , n20692 );
    xnor g13234 ( n26585 , n420 , n18219 );
    not g13235 ( n7503 , n8622 );
    nor g13236 ( n27149 , n25586 , n8491 );
    not g13237 ( n1252 , n3795 );
    and g13238 ( n12120 , n21539 , n6200 );
    or g13239 ( n18523 , n2102 , n598 );
    and g13240 ( n21264 , n18237 , n2847 );
    or g13241 ( n10589 , n25763 , n13145 );
    xnor g13242 ( n10864 , n1705 , n9456 );
    or g13243 ( n21440 , n16453 , n12033 );
    and g13244 ( n5642 , n21383 , n13624 );
    not g13245 ( n4744 , n766 );
    not g13246 ( n2467 , n25718 );
    nor g13247 ( n13326 , n18157 , n2698 );
    nor g13248 ( n21826 , n7335 , n4319 );
    not g13249 ( n7177 , n7010 );
    xnor g13250 ( n25770 , n5847 , n27188 );
    buf g13251 ( n12493 , n24425 );
    or g13252 ( n20412 , n4341 , n5069 );
    not g13253 ( n20020 , n3072 );
    and g13254 ( n347 , n25 , n23382 );
    not g13255 ( n14735 , n21688 );
    not g13256 ( n3093 , n15421 );
    or g13257 ( n13434 , n22644 , n8918 );
    and g13258 ( n10822 , n12846 , n10968 );
    and g13259 ( n9165 , n9821 , n11838 );
    xnor g13260 ( n25214 , n25967 , n4409 );
    or g13261 ( n21944 , n3136 , n4423 );
    xnor g13262 ( n23722 , n16936 , n7515 );
    xnor g13263 ( n3183 , n4999 , n19196 );
    nor g13264 ( n7807 , n21982 , n5760 );
    nor g13265 ( n3011 , n1387 , n2782 );
    not g13266 ( n21070 , n6549 );
    and g13267 ( n16361 , n22362 , n26589 );
    not g13268 ( n21248 , n20080 );
    buf g13269 ( n9883 , n21510 );
    or g13270 ( n7259 , n12962 , n18322 );
    nor g13271 ( n935 , n9347 , n3723 );
    xnor g13272 ( n16083 , n23930 , n14055 );
    nor g13273 ( n8630 , n18371 , n7933 );
    or g13274 ( n3277 , n9587 , n18816 );
    xnor g13275 ( n3741 , n26915 , n14598 );
    xnor g13276 ( n152 , n7498 , n14180 );
    or g13277 ( n891 , n19588 , n8041 );
    and g13278 ( n11828 , n19152 , n22567 );
    and g13279 ( n12259 , n13781 , n10917 );
    or g13280 ( n10900 , n18035 , n3279 );
    or g13281 ( n5618 , n18383 , n17959 );
    and g13282 ( n27106 , n3480 , n11393 );
    nor g13283 ( n6788 , n19680 , n17360 );
    xnor g13284 ( n10973 , n17386 , n5073 );
    not g13285 ( n4181 , n25628 );
    and g13286 ( n2176 , n6851 , n2656 );
    buf g13287 ( n19200 , n19955 );
    xnor g13288 ( n4901 , n20193 , n16768 );
    and g13289 ( n2715 , n4297 , n9171 );
    xnor g13290 ( n27101 , n17198 , n19170 );
    or g13291 ( n21061 , n7930 , n20929 );
    not g13292 ( n17568 , n3425 );
    xnor g13293 ( n21176 , n15181 , n9503 );
    or g13294 ( n25193 , n16760 , n7415 );
    not g13295 ( n9108 , n16874 );
    and g13296 ( n19009 , n26606 , n16914 );
    and g13297 ( n20553 , n14518 , n18806 );
    and g13298 ( n25367 , n1226 , n26610 );
    not g13299 ( n22964 , n2850 );
    xnor g13300 ( n16097 , n6089 , n25476 );
    not g13301 ( n8372 , n1558 );
    nor g13302 ( n22944 , n6397 , n10995 );
    and g13303 ( n18889 , n22268 , n11931 );
    or g13304 ( n26435 , n11363 , n12161 );
    and g13305 ( n3825 , n25522 , n484 );
    xnor g13306 ( n10283 , n15766 , n6105 );
    not g13307 ( n6561 , n10076 );
    xnor g13308 ( n14768 , n13846 , n26625 );
    or g13309 ( n20934 , n8949 , n20469 );
    xnor g13310 ( n14482 , n6694 , n21707 );
    and g13311 ( n5529 , n7954 , n4157 );
    and g13312 ( n10384 , n14719 , n24215 );
    not g13313 ( n1726 , n25843 );
    not g13314 ( n26919 , n791 );
    not g13315 ( n22370 , n21934 );
    or g13316 ( n5979 , n14086 , n25077 );
    xnor g13317 ( n3760 , n509 , n403 );
    or g13318 ( n11082 , n19074 , n15936 );
    xnor g13319 ( n20668 , n15417 , n24578 );
    not g13320 ( n11477 , n26851 );
    not g13321 ( n13206 , n22121 );
    and g13322 ( n10167 , n23141 , n1370 );
    xnor g13323 ( n13284 , n19149 , n11409 );
    and g13324 ( n2127 , n5479 , n9891 );
    not g13325 ( n16514 , n3614 );
    xnor g13326 ( n15343 , n10660 , n8897 );
    and g13327 ( n3693 , n10380 , n1548 );
    not g13328 ( n16210 , n4376 );
    and g13329 ( n21729 , n25376 , n2378 );
    and g13330 ( n10884 , n10747 , n9578 );
    xnor g13331 ( n13444 , n22012 , n18883 );
    or g13332 ( n2591 , n9706 , n24554 );
    or g13333 ( n20806 , n15056 , n13572 );
    xnor g13334 ( n8182 , n19433 , n13951 );
    xnor g13335 ( n9215 , n8831 , n20539 );
    and g13336 ( n19286 , n26029 , n17582 );
    or g13337 ( n17668 , n26760 , n25596 );
    not g13338 ( n8704 , n6032 );
    xnor g13339 ( n23083 , n7799 , n24879 );
    xnor g13340 ( n21834 , n6471 , n15489 );
    or g13341 ( n26 , n13332 , n6112 );
    or g13342 ( n4498 , n16477 , n10767 );
    or g13343 ( n13140 , n23793 , n8596 );
    nor g13344 ( n16776 , n4199 , n6529 );
    xnor g13345 ( n2853 , n7732 , n4898 );
    not g13346 ( n25377 , n11293 );
    or g13347 ( n25645 , n12513 , n8395 );
    xnor g13348 ( n23372 , n20129 , n24035 );
    or g13349 ( n6081 , n15049 , n5139 );
    not g13350 ( n24889 , n2186 );
    or g13351 ( n11175 , n6456 , n17978 );
    nor g13352 ( n11009 , n6729 , n11192 );
    xnor g13353 ( n6988 , n12635 , n17791 );
    not g13354 ( n9569 , n8251 );
    not g13355 ( n9196 , n24323 );
    and g13356 ( n6777 , n20095 , n6980 );
    or g13357 ( n4882 , n1898 , n14395 );
    and g13358 ( n3583 , n19035 , n3539 );
    xnor g13359 ( n16803 , n10730 , n14399 );
    xnor g13360 ( n12433 , n3284 , n15643 );
    nor g13361 ( n9684 , n19609 , n19132 );
    or g13362 ( n14903 , n3956 , n23167 );
    or g13363 ( n22441 , n19460 , n17530 );
    or g13364 ( n8967 , n17979 , n13578 );
    xnor g13365 ( n3806 , n162 , n26174 );
    xnor g13366 ( n3735 , n18975 , n8411 );
    or g13367 ( n3771 , n19384 , n14041 );
    not g13368 ( n18535 , n18488 );
    or g13369 ( n22032 , n17817 , n19900 );
    xnor g13370 ( n1922 , n15769 , n13490 );
    nor g13371 ( n13929 , n8185 , n18402 );
    not g13372 ( n609 , n16840 );
    and g13373 ( n3723 , n17608 , n2591 );
    nor g13374 ( n15015 , n18031 , n21537 );
    xnor g13375 ( n26444 , n953 , n14501 );
    and g13376 ( n25191 , n8181 , n15953 );
    not g13377 ( n146 , n11898 );
    xnor g13378 ( n22452 , n5629 , n15546 );
    and g13379 ( n11130 , n5215 , n14368 );
    and g13380 ( n19977 , n1892 , n26277 );
    not g13381 ( n5143 , n307 );
    or g13382 ( n4740 , n26618 , n12658 );
    or g13383 ( n17413 , n14289 , n17132 );
    or g13384 ( n26827 , n8680 , n16611 );
    nor g13385 ( n8010 , n20512 , n25726 );
    xnor g13386 ( n3307 , n21192 , n13003 );
    or g13387 ( n23040 , n16993 , n3829 );
    or g13388 ( n23761 , n19921 , n14238 );
    xnor g13389 ( n17006 , n18464 , n5548 );
    and g13390 ( n12270 , n12722 , n20236 );
    xnor g13391 ( n4810 , n23350 , n2303 );
    not g13392 ( n26735 , n6053 );
    or g13393 ( n24651 , n20417 , n3568 );
    or g13394 ( n19746 , n12380 , n4191 );
    nor g13395 ( n11449 , n10481 , n3407 );
    or g13396 ( n9286 , n26312 , n8079 );
    or g13397 ( n26960 , n16041 , n5659 );
    xnor g13398 ( n9494 , n13160 , n12148 );
    and g13399 ( n25528 , n10650 , n17978 );
    or g13400 ( n2368 , n9210 , n2729 );
    not g13401 ( n19673 , n7769 );
    or g13402 ( n20105 , n472 , n23586 );
    or g13403 ( n8333 , n15135 , n25712 );
    or g13404 ( n17941 , n19268 , n20452 );
    or g13405 ( n14420 , n13378 , n9323 );
    not g13406 ( n1905 , n4201 );
    and g13407 ( n12737 , n6424 , n15720 );
    not g13408 ( n5122 , n7060 );
    not g13409 ( n13886 , n24926 );
    and g13410 ( n22525 , n12823 , n2674 );
    xnor g13411 ( n24696 , n3018 , n9557 );
    nor g13412 ( n3682 , n10049 , n7621 );
    or g13413 ( n15349 , n14129 , n18286 );
    or g13414 ( n16371 , n23776 , n20556 );
    nor g13415 ( n22396 , n15659 , n6988 );
    nor g13416 ( n23164 , n17593 , n21376 );
    or g13417 ( n2455 , n21934 , n18277 );
    xnor g13418 ( n22863 , n5785 , n6006 );
    nor g13419 ( n640 , n11670 , n8266 );
    nor g13420 ( n1775 , n15073 , n19814 );
    or g13421 ( n14279 , n10492 , n13467 );
    xnor g13422 ( n4777 , n940 , n26763 );
    not g13423 ( n24040 , n5789 );
    nor g13424 ( n26670 , n5891 , n26100 );
    xnor g13425 ( n5856 , n23321 , n6300 );
    xnor g13426 ( n19364 , n16066 , n1712 );
    or g13427 ( n12087 , n17425 , n4068 );
    and g13428 ( n18744 , n5318 , n3943 );
    and g13429 ( n13908 , n13138 , n2068 );
    and g13430 ( n13324 , n2791 , n24027 );
    or g13431 ( n2203 , n22131 , n24064 );
    or g13432 ( n21794 , n2184 , n23109 );
    and g13433 ( n5843 , n26646 , n4329 );
    and g13434 ( n11894 , n24794 , n7826 );
    nor g13435 ( n11236 , n12406 , n16203 );
    and g13436 ( n13525 , n14510 , n7292 );
    and g13437 ( n13125 , n11049 , n15097 );
    xnor g13438 ( n8225 , n15786 , n12177 );
    and g13439 ( n26994 , n10136 , n19519 );
    and g13440 ( n8131 , n2626 , n5821 );
    and g13441 ( n6060 , n7405 , n3350 );
    xnor g13442 ( n12687 , n14335 , n7356 );
    or g13443 ( n23108 , n8782 , n24561 );
    not g13444 ( n26890 , n4901 );
    xnor g13445 ( n7505 , n15146 , n5532 );
    or g13446 ( n20504 , n23208 , n26583 );
    xnor g13447 ( n16440 , n13416 , n20339 );
    xnor g13448 ( n24604 , n18819 , n18011 );
    xnor g13449 ( n7356 , n22379 , n9967 );
    or g13450 ( n21364 , n23157 , n20016 );
    or g13451 ( n1588 , n11841 , n17077 );
    not g13452 ( n20599 , n18926 );
    and g13453 ( n12263 , n7648 , n5289 );
    not g13454 ( n7237 , n23272 );
    or g13455 ( n14281 , n13894 , n10277 );
    or g13456 ( n14847 , n27057 , n2408 );
    xnor g13457 ( n4583 , n312 , n799 );
    or g13458 ( n13134 , n19759 , n23941 );
    and g13459 ( n19027 , n5696 , n23463 );
    or g13460 ( n18442 , n277 , n5112 );
    xnor g13461 ( n1465 , n20559 , n14657 );
    xnor g13462 ( n5559 , n10931 , n12615 );
    or g13463 ( n998 , n22599 , n17897 );
    nor g13464 ( n5729 , n19608 , n15378 );
    and g13465 ( n23552 , n2770 , n2558 );
    and g13466 ( n9326 , n8153 , n19355 );
    or g13467 ( n21813 , n2987 , n13905 );
    or g13468 ( n16344 , n11364 , n18654 );
    and g13469 ( n7194 , n15167 , n25330 );
    and g13470 ( n758 , n2624 , n23336 );
    and g13471 ( n7312 , n2358 , n1208 );
    xnor g13472 ( n17082 , n16697 , n9143 );
    xnor g13473 ( n13614 , n9655 , n23849 );
    or g13474 ( n2778 , n25668 , n18336 );
    nor g13475 ( n1051 , n25524 , n16325 );
    and g13476 ( n19343 , n23062 , n5166 );
    xnor g13477 ( n25984 , n1987 , n11161 );
    xnor g13478 ( n21719 , n17701 , n18092 );
    or g13479 ( n4262 , n18296 , n14207 );
    not g13480 ( n1336 , n23597 );
    or g13481 ( n9537 , n19935 , n8195 );
    xnor g13482 ( n1090 , n19157 , n22878 );
    and g13483 ( n4860 , n12719 , n22187 );
    or g13484 ( n3511 , n4868 , n11425 );
    xnor g13485 ( n992 , n5346 , n19121 );
    not g13486 ( n22158 , n16016 );
    and g13487 ( n16228 , n4899 , n1256 );
    and g13488 ( n24450 , n9444 , n12425 );
    or g13489 ( n11036 , n8265 , n23462 );
    and g13490 ( n14084 , n5658 , n15966 );
    nor g13491 ( n15198 , n7743 , n13263 );
    xnor g13492 ( n13043 , n1173 , n91 );
    and g13493 ( n8073 , n11057 , n10149 );
    and g13494 ( n25652 , n21904 , n17057 );
    not g13495 ( n22859 , n8352 );
    nor g13496 ( n4776 , n21780 , n788 );
    xnor g13497 ( n5042 , n26240 , n20700 );
    or g13498 ( n1409 , n7836 , n19343 );
    nor g13499 ( n21363 , n3868 , n13259 );
    and g13500 ( n5982 , n23726 , n7659 );
    or g13501 ( n22161 , n10146 , n26660 );
    or g13502 ( n13279 , n14955 , n13098 );
    xnor g13503 ( n26068 , n1658 , n19464 );
    or g13504 ( n4044 , n24856 , n17724 );
    and g13505 ( n25924 , n22128 , n5306 );
    and g13506 ( n12023 , n24771 , n22046 );
    and g13507 ( n4059 , n21815 , n11012 );
    or g13508 ( n26626 , n25941 , n13958 );
    xnor g13509 ( n9633 , n5311 , n11717 );
    not g13510 ( n23456 , n13133 );
    xnor g13511 ( n26420 , n5718 , n22643 );
    and g13512 ( n53 , n18220 , n20634 );
    or g13513 ( n3278 , n20505 , n11539 );
    not g13514 ( n16024 , n886 );
    not g13515 ( n24661 , n6102 );
    xnor g13516 ( n13610 , n4230 , n16290 );
    nor g13517 ( n3633 , n3601 , n23894 );
    or g13518 ( n5462 , n6400 , n17864 );
    and g13519 ( n18631 , n17123 , n21026 );
    nor g13520 ( n11750 , n25164 , n6285 );
    not g13521 ( n1909 , n9289 );
    and g13522 ( n20526 , n1015 , n26922 );
    not g13523 ( n2559 , n22631 );
    not g13524 ( n6203 , n9512 );
    or g13525 ( n1492 , n24485 , n14356 );
    xnor g13526 ( n7236 , n14039 , n4396 );
    xnor g13527 ( n17792 , n10329 , n23222 );
    and g13528 ( n17249 , n13721 , n16353 );
    or g13529 ( n7251 , n6209 , n4326 );
    xnor g13530 ( n16688 , n10073 , n6683 );
    not g13531 ( n22139 , n8997 );
    xnor g13532 ( n6196 , n23290 , n1939 );
    or g13533 ( n8557 , n19082 , n8910 );
    xnor g13534 ( n23240 , n7750 , n7284 );
    and g13535 ( n18536 , n23742 , n6425 );
    or g13536 ( n24591 , n11790 , n8279 );
    xnor g13537 ( n6387 , n3060 , n3979 );
    xnor g13538 ( n6169 , n20322 , n19334 );
    xnor g13539 ( n23543 , n3018 , n18537 );
    xnor g13540 ( n5911 , n19537 , n26668 );
    or g13541 ( n9697 , n23497 , n22413 );
    or g13542 ( n23205 , n21681 , n15373 );
    and g13543 ( n11747 , n25457 , n9949 );
    nor g13544 ( n8801 , n10405 , n25370 );
    xnor g13545 ( n25864 , n10782 , n15150 );
    and g13546 ( n5361 , n7877 , n21591 );
    or g13547 ( n4507 , n24403 , n13667 );
    xnor g13548 ( n12364 , n15110 , n22940 );
    not g13549 ( n25663 , n19941 );
    not g13550 ( n17547 , n5510 );
    xnor g13551 ( n3564 , n12470 , n14750 );
    xnor g13552 ( n25198 , n61 , n15761 );
    or g13553 ( n9230 , n11338 , n12633 );
    and g13554 ( n19342 , n74 , n22984 );
    xnor g13555 ( n27163 , n3557 , n14985 );
    nor g13556 ( n4849 , n16364 , n7680 );
    or g13557 ( n14467 , n25126 , n22097 );
    not g13558 ( n11240 , n1218 );
    and g13559 ( n12308 , n11021 , n26507 );
    or g13560 ( n15199 , n386 , n21758 );
    not g13561 ( n23639 , n9179 );
    or g13562 ( n13962 , n11072 , n18728 );
    xnor g13563 ( n22914 , n7054 , n3057 );
    not g13564 ( n13980 , n21451 );
    nor g13565 ( n20955 , n8520 , n17590 );
    xnor g13566 ( n11688 , n17043 , n23103 );
    or g13567 ( n10522 , n4534 , n10654 );
    or g13568 ( n6318 , n12530 , n23657 );
    or g13569 ( n9056 , n5977 , n8894 );
    or g13570 ( n26362 , n8209 , n19479 );
    or g13571 ( n5147 , n17453 , n16903 );
    or g13572 ( n6977 , n3452 , n555 );
    not g13573 ( n26506 , n3483 );
    xnor g13574 ( n18232 , n23519 , n4092 );
    and g13575 ( n25809 , n17021 , n1010 );
    nor g13576 ( n19996 , n11459 , n18781 );
    xnor g13577 ( n18311 , n8513 , n8578 );
    or g13578 ( n22991 , n2423 , n2197 );
    or g13579 ( n22334 , n7571 , n21484 );
    or g13580 ( n1013 , n10424 , n21206 );
    and g13581 ( n1321 , n4669 , n7556 );
    xnor g13582 ( n24269 , n17705 , n22421 );
    or g13583 ( n19555 , n21951 , n10383 );
    nor g13584 ( n22053 , n22849 , n405 );
    not g13585 ( n10978 , n22097 );
    xnor g13586 ( n19691 , n12576 , n18130 );
    xnor g13587 ( n12192 , n1194 , n7881 );
    xnor g13588 ( n20418 , n20444 , n12112 );
    xnor g13589 ( n5205 , n19739 , n25883 );
    xnor g13590 ( n18210 , n10514 , n6105 );
    or g13591 ( n20636 , n13304 , n14416 );
    or g13592 ( n15575 , n13189 , n18258 );
    xnor g13593 ( n12992 , n7159 , n21818 );
    and g13594 ( n12695 , n12879 , n9338 );
    xnor g13595 ( n9054 , n11036 , n22618 );
    nor g13596 ( n23124 , n26344 , n14754 );
    xnor g13597 ( n21049 , n15417 , n18792 );
    xnor g13598 ( n10033 , n23162 , n19241 );
    nor g13599 ( n8746 , n6946 , n20124 );
    or g13600 ( n17059 , n16648 , n13377 );
    xnor g13601 ( n24870 , n7823 , n1 );
    or g13602 ( n20735 , n16415 , n8465 );
    and g13603 ( n16467 , n21784 , n18163 );
    or g13604 ( n12015 , n1582 , n17699 );
    nor g13605 ( n13510 , n26749 , n2938 );
    xnor g13606 ( n13556 , n12758 , n8760 );
    and g13607 ( n26596 , n24417 , n24907 );
    not g13608 ( n7776 , n9809 );
    not g13609 ( n24359 , n14080 );
    or g13610 ( n16651 , n1423 , n5346 );
    xnor g13611 ( n11386 , n18458 , n5470 );
    or g13612 ( n8327 , n20597 , n109 );
    xnor g13613 ( n1996 , n22492 , n25523 );
    or g13614 ( n1969 , n8322 , n15659 );
    xnor g13615 ( n21833 , n380 , n824 );
    xnor g13616 ( n14215 , n24124 , n10838 );
    or g13617 ( n4413 , n13137 , n3274 );
    and g13618 ( n25081 , n23869 , n22127 );
    not g13619 ( n19502 , n3150 );
    xnor g13620 ( n20072 , n13543 , n6794 );
    xnor g13621 ( n6431 , n23459 , n6196 );
    xnor g13622 ( n26604 , n19531 , n1999 );
    or g13623 ( n21757 , n16454 , n10584 );
    or g13624 ( n1702 , n15221 , n21853 );
    and g13625 ( n15421 , n24652 , n26418 );
    and g13626 ( n13985 , n5255 , n25289 );
    not g13627 ( n14344 , n7593 );
    and g13628 ( n23044 , n23470 , n9009 );
    and g13629 ( n19946 , n25754 , n12294 );
    or g13630 ( n14143 , n23002 , n13556 );
    xnor g13631 ( n26387 , n26968 , n25336 );
    xnor g13632 ( n11382 , n15523 , n7711 );
    and g13633 ( n25933 , n17069 , n19446 );
    or g13634 ( n6090 , n12973 , n19742 );
    not g13635 ( n14341 , n2728 );
    not g13636 ( n26946 , n15961 );
    and g13637 ( n11637 , n8713 , n54 );
    nor g13638 ( n23088 , n387 , n12293 );
    or g13639 ( n15412 , n16216 , n18356 );
    xnor g13640 ( n20898 , n25376 , n2378 );
    xnor g13641 ( n16979 , n6670 , n10023 );
    nor g13642 ( n12582 , n21998 , n25779 );
    or g13643 ( n26547 , n20497 , n21997 );
    or g13644 ( n21171 , n2628 , n15383 );
    not g13645 ( n10230 , n5490 );
    or g13646 ( n24054 , n13913 , n13843 );
    or g13647 ( n3014 , n23386 , n15374 );
    or g13648 ( n12019 , n4087 , n4667 );
    xnor g13649 ( n6706 , n558 , n2765 );
    or g13650 ( n7727 , n24065 , n20307 );
    xnor g13651 ( n25487 , n8305 , n22253 );
    or g13652 ( n27088 , n19192 , n15511 );
    not g13653 ( n1088 , n7207 );
    not g13654 ( n15616 , n26306 );
    or g13655 ( n18051 , n22285 , n25998 );
    xnor g13656 ( n1808 , n9979 , n27007 );
    xnor g13657 ( n521 , n25495 , n9152 );
    or g13658 ( n11269 , n1786 , n5408 );
    and g13659 ( n15045 , n3568 , n18202 );
    xnor g13660 ( n23688 , n19995 , n1008 );
    or g13661 ( n1556 , n22135 , n1609 );
    xnor g13662 ( n19909 , n13990 , n2307 );
    or g13663 ( n17094 , n9318 , n1022 );
    or g13664 ( n23171 , n13817 , n272 );
    xnor g13665 ( n15352 , n6691 , n21753 );
    or g13666 ( n22578 , n20158 , n4538 );
    or g13667 ( n17030 , n11592 , n14003 );
    and g13668 ( n13313 , n22572 , n12752 );
    and g13669 ( n26233 , n27166 , n10850 );
    nor g13670 ( n15553 , n15164 , n16313 );
    xnor g13671 ( n20689 , n25231 , n11109 );
    not g13672 ( n14397 , n18326 );
    not g13673 ( n7160 , n4288 );
    or g13674 ( n18124 , n22134 , n11940 );
    xnor g13675 ( n23361 , n10201 , n6814 );
    or g13676 ( n8237 , n12579 , n14043 );
    xnor g13677 ( n25519 , n11066 , n1552 );
    xnor g13678 ( n9120 , n15787 , n7486 );
    xnor g13679 ( n18734 , n495 , n22999 );
    xnor g13680 ( n14156 , n9320 , n13614 );
    or g13681 ( n18832 , n6584 , n4474 );
    xnor g13682 ( n25839 , n24686 , n25451 );
    xnor g13683 ( n4198 , n12477 , n18035 );
    and g13684 ( n3243 , n13039 , n6043 );
    and g13685 ( n5773 , n10302 , n2273 );
    or g13686 ( n27133 , n23781 , n22904 );
    and g13687 ( n21339 , n11914 , n17158 );
    or g13688 ( n19672 , n20342 , n14826 );
    not g13689 ( n18031 , n16744 );
    xnor g13690 ( n15958 , n6964 , n22064 );
    nor g13691 ( n9829 , n11220 , n4299 );
    xnor g13692 ( n7180 , n19078 , n18039 );
    nor g13693 ( n12872 , n18269 , n5026 );
    nor g13694 ( n24905 , n6082 , n23097 );
    or g13695 ( n9754 , n2995 , n17428 );
    and g13696 ( n10999 , n19025 , n21962 );
    xnor g13697 ( n25413 , n9721 , n3916 );
    xnor g13698 ( n5120 , n4684 , n23220 );
    or g13699 ( n20792 , n19081 , n26316 );
    nor g13700 ( n10166 , n23168 , n3962 );
    and g13701 ( n16852 , n24301 , n9669 );
    or g13702 ( n26112 , n14936 , n6502 );
    xnor g13703 ( n12279 , n23394 , n2305 );
    and g13704 ( n19468 , n14592 , n12957 );
    xnor g13705 ( n22371 , n22382 , n26471 );
    xnor g13706 ( n26081 , n26224 , n18483 );
    or g13707 ( n5975 , n15083 , n22431 );
    and g13708 ( n18275 , n1651 , n23350 );
    and g13709 ( n3510 , n16604 , n23348 );
    not g13710 ( n22571 , n949 );
    not g13711 ( n22363 , n852 );
    and g13712 ( n10193 , n16825 , n17703 );
    or g13713 ( n22570 , n4849 , n26245 );
    or g13714 ( n9543 , n24391 , n12704 );
    or g13715 ( n8639 , n12250 , n24525 );
    or g13716 ( n2851 , n3000 , n26385 );
    not g13717 ( n6842 , n19366 );
    or g13718 ( n10828 , n15943 , n19591 );
    xnor g13719 ( n10059 , n18710 , n21796 );
    and g13720 ( n17272 , n19974 , n22440 );
    or g13721 ( n10433 , n20956 , n6699 );
    not g13722 ( n2750 , n15675 );
    or g13723 ( n17747 , n9099 , n5745 );
    xnor g13724 ( n22327 , n17783 , n16337 );
    not g13725 ( n2126 , n23591 );
    or g13726 ( n20551 , n26782 , n11088 );
    or g13727 ( n6845 , n14145 , n22436 );
    or g13728 ( n8031 , n4645 , n7985 );
    or g13729 ( n19077 , n2579 , n19081 );
    or g13730 ( n1438 , n15884 , n5213 );
    and g13731 ( n37 , n24316 , n12745 );
    or g13732 ( n13918 , n23837 , n23242 );
    xnor g13733 ( n18102 , n17251 , n4913 );
    or g13734 ( n19690 , n22155 , n11823 );
    xnor g13735 ( n7634 , n5528 , n15828 );
    or g13736 ( n8972 , n8754 , n10344 );
    buf g13737 ( n8930 , n18429 );
    nor g13738 ( n8078 , n20151 , n20429 );
    xnor g13739 ( n2612 , n10037 , n13148 );
    or g13740 ( n24192 , n12513 , n8162 );
    not g13741 ( n4955 , n6925 );
    and g13742 ( n8929 , n13714 , n1329 );
    xnor g13743 ( n7280 , n18658 , n11928 );
    and g13744 ( n21906 , n4882 , n12637 );
    nor g13745 ( n6702 , n3498 , n14289 );
    not g13746 ( n20344 , n25415 );
    xnor g13747 ( n11928 , n5949 , n21969 );
    xnor g13748 ( n7686 , n19091 , n2275 );
    and g13749 ( n15591 , n3172 , n17238 );
    and g13750 ( n21700 , n13677 , n10451 );
    nor g13751 ( n24521 , n8367 , n726 );
    and g13752 ( n10336 , n24142 , n10569 );
    xnor g13753 ( n887 , n1471 , n3152 );
    xnor g13754 ( n6559 , n25296 , n23717 );
    or g13755 ( n26400 , n9216 , n25107 );
    not g13756 ( n18179 , n8814 );
    or g13757 ( n19213 , n21218 , n9815 );
    and g13758 ( n9641 , n12953 , n22328 );
    nor g13759 ( n13765 , n481 , n15474 );
    or g13760 ( n1718 , n26789 , n11733 );
    and g13761 ( n719 , n14358 , n6986 );
    nor g13762 ( n3153 , n19482 , n4177 );
    xnor g13763 ( n27112 , n21130 , n18154 );
    xnor g13764 ( n25603 , n3954 , n18611 );
    xnor g13765 ( n771 , n26889 , n6961 );
    xnor g13766 ( n4063 , n16722 , n6385 );
    xnor g13767 ( n25812 , n23254 , n27008 );
    not g13768 ( n11052 , n17784 );
    not g13769 ( n5783 , n7670 );
    not g13770 ( n19828 , n20819 );
    xnor g13771 ( n18291 , n14886 , n933 );
    or g13772 ( n11263 , n2023 , n19489 );
    or g13773 ( n17043 , n20985 , n25304 );
    xnor g13774 ( n13761 , n13436 , n25693 );
    not g13775 ( n22386 , n16701 );
    xnor g13776 ( n25155 , n6989 , n23257 );
    or g13777 ( n10888 , n22948 , n18165 );
    or g13778 ( n25995 , n9874 , n6816 );
    or g13779 ( n11307 , n8419 , n23727 );
    and g13780 ( n10198 , n10473 , n25429 );
    not g13781 ( n11831 , n16117 );
    xnor g13782 ( n18045 , n9237 , n24508 );
    or g13783 ( n1274 , n13237 , n5568 );
    not g13784 ( n2492 , n23346 );
    and g13785 ( n10872 , n14695 , n15473 );
    xnor g13786 ( n24798 , n22626 , n3324 );
    xnor g13787 ( n23693 , n22314 , n22473 );
    or g13788 ( n27128 , n707 , n21418 );
    or g13789 ( n7901 , n1646 , n4191 );
    xnor g13790 ( n24156 , n24045 , n21433 );
    not g13791 ( n4298 , n17705 );
    nor g13792 ( n26184 , n5098 , n7436 );
    or g13793 ( n5992 , n12583 , n25593 );
    xnor g13794 ( n10116 , n27014 , n10322 );
    xnor g13795 ( n17462 , n10001 , n21263 );
    and g13796 ( n9159 , n21974 , n22284 );
    nor g13797 ( n15025 , n6814 , n8084 );
    not g13798 ( n223 , n21223 );
    nor g13799 ( n11897 , n7234 , n15360 );
    xnor g13800 ( n18862 , n18247 , n2409 );
    nor g13801 ( n19264 , n9359 , n24802 );
    and g13802 ( n26341 , n162 , n20509 );
    xnor g13803 ( n6115 , n4504 , n14577 );
    xnor g13804 ( n4008 , n11621 , n23965 );
    xnor g13805 ( n19534 , n6631 , n24732 );
    and g13806 ( n8842 , n26168 , n19660 );
    or g13807 ( n4463 , n15415 , n4395 );
    xnor g13808 ( n24841 , n17874 , n20802 );
    and g13809 ( n12935 , n5635 , n17153 );
    not g13810 ( n22278 , n25632 );
    not g13811 ( n5185 , n13719 );
    or g13812 ( n19853 , n25407 , n20979 );
    or g13813 ( n18074 , n15204 , n18478 );
    xnor g13814 ( n3869 , n21722 , n10504 );
    xnor g13815 ( n25540 , n405 , n4561 );
    xnor g13816 ( n25793 , n26452 , n2999 );
    and g13817 ( n5590 , n18428 , n16793 );
    xnor g13818 ( n24171 , n3009 , n21729 );
    or g13819 ( n13670 , n535 , n2705 );
    nor g13820 ( n7472 , n23161 , n3383 );
    and g13821 ( n25219 , n6097 , n11686 );
    nor g13822 ( n13428 , n25900 , n22715 );
    xnor g13823 ( n7284 , n15788 , n12556 );
    not g13824 ( n17110 , n3460 );
    and g13825 ( n13449 , n23863 , n11114 );
    nor g13826 ( n10088 , n9554 , n8176 );
    nor g13827 ( n11283 , n6610 , n7752 );
    or g13828 ( n6635 , n18100 , n16231 );
    or g13829 ( n18120 , n25957 , n19247 );
    xnor g13830 ( n15273 , n5998 , n14352 );
    or g13831 ( n25145 , n21883 , n15615 );
    xnor g13832 ( n10820 , n18333 , n11497 );
    not g13833 ( n26178 , n1552 );
    not g13834 ( n4706 , n19486 );
    not g13835 ( n19872 , n21143 );
    xnor g13836 ( n243 , n25127 , n19734 );
    xnor g13837 ( n19403 , n4652 , n8521 );
    xnor g13838 ( n21353 , n25849 , n7167 );
    or g13839 ( n23975 , n19088 , n17516 );
    xnor g13840 ( n5703 , n10072 , n21159 );
    nor g13841 ( n20730 , n21334 , n15273 );
    and g13842 ( n22135 , n18724 , n138 );
    and g13843 ( n12684 , n9144 , n25236 );
    or g13844 ( n1283 , n20292 , n15119 );
    and g13845 ( n23262 , n20276 , n16292 );
    xnor g13846 ( n9022 , n23044 , n22201 );
    or g13847 ( n12173 , n1597 , n26924 );
    not g13848 ( n5525 , n6413 );
    xnor g13849 ( n23784 , n16471 , n12835 );
    or g13850 ( n16120 , n20796 , n26444 );
    or g13851 ( n2032 , n17626 , n25241 );
    xnor g13852 ( n23305 , n21569 , n13151 );
    nor g13853 ( n415 , n25566 , n16233 );
    or g13854 ( n21129 , n14718 , n14440 );
    or g13855 ( n18866 , n6600 , n18910 );
    xnor g13856 ( n19368 , n7653 , n579 );
    and g13857 ( n7742 , n4049 , n19529 );
    or g13858 ( n17722 , n25931 , n1510 );
    xnor g13859 ( n17936 , n4028 , n17569 );
    xnor g13860 ( n9403 , n14220 , n10362 );
    or g13861 ( n10073 , n17105 , n24819 );
    xnor g13862 ( n9566 , n25452 , n3673 );
    xnor g13863 ( n2185 , n5205 , n23586 );
    nor g13864 ( n15364 , n13349 , n8856 );
    not g13865 ( n9935 , n7131 );
    nor g13866 ( n13817 , n1182 , n2743 );
    or g13867 ( n23770 , n5590 , n18682 );
    xnor g13868 ( n25069 , n17442 , n15424 );
    not g13869 ( n4518 , n21760 );
    xnor g13870 ( n9435 , n7512 , n6133 );
    and g13871 ( n1218 , n16358 , n21331 );
    and g13872 ( n13228 , n1219 , n3374 );
    and g13873 ( n928 , n12369 , n15646 );
    or g13874 ( n23948 , n15747 , n11994 );
    and g13875 ( n22750 , n3188 , n9862 );
    xnor g13876 ( n16645 , n19282 , n2978 );
    or g13877 ( n2430 , n21421 , n16647 );
    not g13878 ( n17098 , n15883 );
    nor g13879 ( n1447 , n8155 , n17287 );
    xnor g13880 ( n25938 , n21447 , n7779 );
    or g13881 ( n13318 , n16824 , n25353 );
    xnor g13882 ( n3733 , n17952 , n22756 );
    nor g13883 ( n1054 , n2914 , n13914 );
    or g13884 ( n26595 , n17352 , n4043 );
    or g13885 ( n7287 , n19157 , n12138 );
    xnor g13886 ( n6453 , n11211 , n26522 );
    xnor g13887 ( n15243 , n2160 , n19282 );
    nor g13888 ( n8955 , n13425 , n22215 );
    or g13889 ( n6646 , n1018 , n2616 );
    xnor g13890 ( n24860 , n24070 , n661 );
    xnor g13891 ( n18310 , n25961 , n15225 );
    and g13892 ( n4551 , n10898 , n25750 );
    xnor g13893 ( n24834 , n25370 , n4426 );
    and g13894 ( n3580 , n18407 , n18866 );
    and g13895 ( n11092 , n8255 , n5 );
    or g13896 ( n6428 , n26268 , n1258 );
    and g13897 ( n25185 , n15876 , n22367 );
    not g13898 ( n26786 , n26422 );
    xor g13899 ( n15565 , n586 , n21226 );
    and g13900 ( n26995 , n13086 , n14303 );
    or g13901 ( n7812 , n1654 , n24245 );
    or g13902 ( n2347 , n17100 , n24390 );
    or g13903 ( n13128 , n23230 , n20488 );
    xnor g13904 ( n13622 , n18371 , n21151 );
    and g13905 ( n23666 , n18344 , n2965 );
    xnor g13906 ( n3554 , n15777 , n5857 );
    and g13907 ( n1148 , n119 , n20459 );
    xnor g13908 ( n11674 , n550 , n7928 );
    nor g13909 ( n1265 , n11382 , n17607 );
    not g13910 ( n19215 , n20530 );
    xnor g13911 ( n19142 , n2944 , n22270 );
    or g13912 ( n18242 , n15640 , n1221 );
    or g13913 ( n19984 , n14856 , n11192 );
    xnor g13914 ( n24347 , n19124 , n6897 );
    or g13915 ( n24858 , n25201 , n4057 );
    and g13916 ( n181 , n11043 , n25117 );
    buf g13917 ( n6692 , n2324 );
    xnor g13918 ( n1778 , n4003 , n17959 );
    and g13919 ( n10954 , n13670 , n17029 );
    xnor g13920 ( n9322 , n14265 , n25667 );
    xnor g13921 ( n10316 , n9003 , n13453 );
    and g13922 ( n11811 , n8326 , n26456 );
    nor g13923 ( n13889 , n8638 , n23018 );
    not g13924 ( n11767 , n3535 );
    xnor g13925 ( n5700 , n6396 , n26740 );
    or g13926 ( n27116 , n1672 , n16765 );
    not g13927 ( n22426 , n14575 );
    or g13928 ( n9178 , n12900 , n16547 );
    xnor g13929 ( n25080 , n7841 , n22918 );
    or g13930 ( n168 , n12094 , n25724 );
    not g13931 ( n3391 , n21626 );
    xnor g13932 ( n5813 , n17250 , n10125 );
    xnor g13933 ( n19117 , n23 , n20626 );
    not g13934 ( n23071 , n18466 );
    not g13935 ( n26008 , n19638 );
    nor g13936 ( n23419 , n21937 , n11736 );
    nor g13937 ( n3327 , n17739 , n4400 );
    xnor g13938 ( n15261 , n19960 , n16140 );
    not g13939 ( n18473 , n2731 );
    xnor g13940 ( n18520 , n4245 , n18577 );
    xnor g13941 ( n17741 , n7217 , n8324 );
    xnor g13942 ( n26707 , n21662 , n14943 );
    and g13943 ( n26472 , n9204 , n12251 );
    xnor g13944 ( n1714 , n12972 , n16719 );
    and g13945 ( n6892 , n15628 , n21722 );
    or g13946 ( n6757 , n26415 , n24088 );
    nor g13947 ( n15599 , n8625 , n7291 );
    not g13948 ( n26717 , n12161 );
    xnor g13949 ( n26484 , n6179 , n18345 );
    xnor g13950 ( n11489 , n14062 , n8837 );
    not g13951 ( n7902 , n25864 );
    xnor g13952 ( n379 , n26009 , n7354 );
    or g13953 ( n1248 , n3173 , n2841 );
    and g13954 ( n26176 , n750 , n11520 );
    nor g13955 ( n3698 , n18287 , n406 );
    xnor g13956 ( n25515 , n3434 , n2301 );
    nor g13957 ( n26809 , n14113 , n8172 );
    not g13958 ( n15583 , n18877 );
    xnor g13959 ( n22563 , n6204 , n3795 );
    nor g13960 ( n17116 , n5213 , n24617 );
    not g13961 ( n26997 , n11044 );
    and g13962 ( n20227 , n15838 , n2398 );
    xnor g13963 ( n24052 , n10932 , n26764 );
    nor g13964 ( n5019 , n2780 , n10411 );
    xnor g13965 ( n25355 , n16535 , n15908 );
    and g13966 ( n21791 , n5704 , n24665 );
    xnor g13967 ( n20057 , n20970 , n13367 );
    not g13968 ( n26255 , n21078 );
    xnor g13969 ( n2199 , n5990 , n21208 );
    xnor g13970 ( n8784 , n18492 , n12813 );
    nor g13971 ( n17254 , n20536 , n3349 );
    and g13972 ( n18836 , n9103 , n3342 );
    nor g13973 ( n11855 , n12861 , n15064 );
    xnor g13974 ( n3573 , n2675 , n5139 );
    and g13975 ( n6286 , n2836 , n18436 );
    not g13976 ( n14923 , n19982 );
    or g13977 ( n3567 , n1541 , n25495 );
    nor g13978 ( n26640 , n20009 , n23980 );
    or g13979 ( n15786 , n20251 , n10942 );
    nor g13980 ( n17831 , n22222 , n7761 );
    xnor g13981 ( n16674 , n26010 , n6661 );
    or g13982 ( n25149 , n7111 , n926 );
    xnor g13983 ( n15319 , n5451 , n3918 );
    and g13984 ( n25040 , n4304 , n19413 );
    xnor g13985 ( n6859 , n22218 , n3431 );
    not g13986 ( n24862 , n23612 );
    xnor g13987 ( n7767 , n21764 , n5483 );
    not g13988 ( n10934 , n9504 );
    or g13989 ( n13773 , n3468 , n15289 );
    nor g13990 ( n5895 , n3582 , n21784 );
    not g13991 ( n10666 , n5167 );
    nor g13992 ( n21423 , n23352 , n25659 );
    nor g13993 ( n18327 , n18338 , n18672 );
    nor g13994 ( n15055 , n13783 , n22332 );
    or g13995 ( n4335 , n25566 , n3581 );
    or g13996 ( n12954 , n14486 , n18735 );
    not g13997 ( n15875 , n2233 );
    not g13998 ( n24902 , n16374 );
    or g13999 ( n23267 , n6935 , n16808 );
    or g14000 ( n6282 , n2812 , n8363 );
    or g14001 ( n18697 , n14402 , n20785 );
    xnor g14002 ( n21449 , n25015 , n1850 );
    or g14003 ( n5282 , n16872 , n25027 );
    and g14004 ( n8904 , n21450 , n4870 );
    not g14005 ( n11384 , n25923 );
    xnor g14006 ( n25568 , n19772 , n6866 );
    xnor g14007 ( n15779 , n10995 , n11736 );
    xnor g14008 ( n14387 , n986 , n3122 );
    or g14009 ( n22896 , n20037 , n1207 );
    and g14010 ( n8951 , n23125 , n15080 );
    xnor g14011 ( n14685 , n8512 , n2819 );
    nor g14012 ( n10909 , n306 , n13936 );
    xnor g14013 ( n8521 , n9132 , n3611 );
    xnor g14014 ( n4015 , n20120 , n13129 );
    not g14015 ( n15267 , n15475 );
    xnor g14016 ( n21397 , n790 , n5914 );
    or g14017 ( n4750 , n18408 , n4283 );
    xnor g14018 ( n22476 , n21937 , n10706 );
    xnor g14019 ( n26185 , n21 , n23513 );
    and g14020 ( n2799 , n19531 , n26872 );
    and g14021 ( n1153 , n14173 , n9772 );
    or g14022 ( n9195 , n15173 , n6415 );
    or g14023 ( n27014 , n9956 , n24294 );
    not g14024 ( n15193 , n24496 );
    or g14025 ( n6326 , n26423 , n21530 );
    and g14026 ( n5921 , n458 , n26101 );
    xnor g14027 ( n13808 , n25330 , n15167 );
    xnor g14028 ( n10051 , n2379 , n15319 );
    and g14029 ( n4318 , n14899 , n10408 );
    or g14030 ( n16740 , n12688 , n26249 );
    nor g14031 ( n13392 , n20707 , n9780 );
    or g14032 ( n9839 , n22273 , n9605 );
    or g14033 ( n6449 , n21756 , n17178 );
    not g14034 ( n2775 , n5236 );
    or g14035 ( n4332 , n6120 , n23197 );
    nor g14036 ( n14560 , n5990 , n21208 );
    and g14037 ( n12415 , n13763 , n118 );
    xnor g14038 ( n7519 , n20376 , n6202 );
    and g14039 ( n7527 , n23219 , n23764 );
    and g14040 ( n25037 , n17741 , n10451 );
    or g14041 ( n15653 , n23029 , n17840 );
    nor g14042 ( n25762 , n8496 , n1574 );
    xnor g14043 ( n5214 , n18994 , n2100 );
    xnor g14044 ( n17529 , n662 , n18736 );
    not g14045 ( n19391 , n3836 );
    or g14046 ( n9154 , n3622 , n15764 );
    xnor g14047 ( n24969 , n2493 , n9442 );
    nor g14048 ( n23276 , n14936 , n5740 );
    xnor g14049 ( n10585 , n21489 , n4085 );
    and g14050 ( n16070 , n10580 , n12084 );
    not g14051 ( n15959 , n7216 );
    or g14052 ( n23027 , n13237 , n1066 );
    xnor g14053 ( n23567 , n26939 , n20259 );
    or g14054 ( n13647 , n23912 , n22716 );
    or g14055 ( n16434 , n22687 , n11734 );
    xnor g14056 ( n20624 , n4612 , n7118 );
    xnor g14057 ( n12350 , n14244 , n16705 );
    xnor g14058 ( n17721 , n24525 , n22267 );
    not g14059 ( n15427 , n16994 );
    or g14060 ( n5808 , n5942 , n7023 );
    or g14061 ( n22023 , n3623 , n6444 );
    or g14062 ( n15532 , n12161 , n24886 );
    nor g14063 ( n3495 , n3460 , n19477 );
    not g14064 ( n12149 , n22557 );
    and g14065 ( n5835 , n11183 , n16891 );
    or g14066 ( n192 , n23119 , n16591 );
    not g14067 ( n6660 , n6371 );
    or g14068 ( n22446 , n26512 , n4909 );
    xnor g14069 ( n10034 , n87 , n10129 );
    nor g14070 ( n13807 , n6239 , n20209 );
    or g14071 ( n14053 , n379 , n20671 );
    or g14072 ( n10523 , n10916 , n5835 );
    not g14073 ( n21029 , n18107 );
    not g14074 ( n24329 , n21884 );
    or g14075 ( n5807 , n16791 , n26967 );
    or g14076 ( n14748 , n22751 , n6505 );
    not g14077 ( n25692 , n14458 );
    or g14078 ( n3933 , n16227 , n21226 );
    and g14079 ( n2359 , n9034 , n19959 );
    or g14080 ( n11642 , n3134 , n24135 );
    xnor g14081 ( n11094 , n23941 , n11196 );
    or g14082 ( n23260 , n25571 , n7978 );
    xnor g14083 ( n4828 , n6200 , n14257 );
    xnor g14084 ( n16993 , n21503 , n20269 );
    xnor g14085 ( n2892 , n3199 , n22782 );
    xnor g14086 ( n14891 , n27203 , n25202 );
    xnor g14087 ( n5472 , n1321 , n2665 );
    or g14088 ( n7196 , n16103 , n4990 );
    nor g14089 ( n7907 , n20411 , n9512 );
    and g14090 ( n24848 , n6613 , n8933 );
    and g14091 ( n14429 , n13664 , n6197 );
    nor g14092 ( n20178 , n25120 , n8526 );
    nor g14093 ( n14799 , n1534 , n6201 );
    not g14094 ( n8607 , n25455 );
    or g14095 ( n1408 , n17782 , n16782 );
    or g14096 ( n21639 , n14966 , n19370 );
    or g14097 ( n23563 , n26782 , n11069 );
    xnor g14098 ( n13754 , n27034 , n11995 );
    not g14099 ( n328 , n24032 );
    not g14100 ( n26629 , n1183 );
    xnor g14101 ( n7833 , n25366 , n25949 );
    and g14102 ( n17224 , n5714 , n26409 );
    and g14103 ( n23566 , n10156 , n20551 );
    or g14104 ( n7225 , n13935 , n11841 );
    or g14105 ( n4763 , n3749 , n21342 );
    xnor g14106 ( n9084 , n21089 , n23086 );
    nor g14107 ( n1563 , n25040 , n9060 );
    not g14108 ( n6446 , n851 );
    and g14109 ( n23540 , n23923 , n23874 );
    buf g14110 ( n19460 , n1092 );
    xnor g14111 ( n15132 , n25357 , n15499 );
    and g14112 ( n17490 , n17177 , n18712 );
    and g14113 ( n11769 , n4740 , n26614 );
    or g14114 ( n16173 , n7340 , n24448 );
    not g14115 ( n1061 , n23201 );
    xnor g14116 ( n26826 , n9814 , n9274 );
    or g14117 ( n119 , n18256 , n14958 );
    xnor g14118 ( n13251 , n24624 , n17090 );
    or g14119 ( n18663 , n2371 , n14713 );
    and g14120 ( n1983 , n25788 , n8697 );
    and g14121 ( n2625 , n21301 , n8912 );
    or g14122 ( n8440 , n15796 , n4836 );
    or g14123 ( n1696 , n15321 , n1652 );
    or g14124 ( n20203 , n22030 , n3754 );
    or g14125 ( n13880 , n1954 , n4575 );
    nor g14126 ( n14882 , n13621 , n16130 );
    or g14127 ( n11992 , n14570 , n1528 );
    and g14128 ( n288 , n16824 , n26295 );
    xnor g14129 ( n13631 , n9940 , n8013 );
    and g14130 ( n12839 , n6004 , n18567 );
    or g14131 ( n6549 , n6195 , n20608 );
    and g14132 ( n8730 , n2775 , n22852 );
    or g14133 ( n4747 , n18902 , n8643 );
    xnor g14134 ( n18644 , n19472 , n21226 );
    not g14135 ( n24880 , n10787 );
    xnor g14136 ( n4370 , n26810 , n26660 );
    not g14137 ( n12306 , n7837 );
    or g14138 ( n25429 , n8998 , n25378 );
    or g14139 ( n3576 , n6701 , n7195 );
    xnor g14140 ( n5787 , n24118 , n13271 );
    or g14141 ( n3406 , n23231 , n10114 );
    or g14142 ( n16998 , n1630 , n16147 );
    and g14143 ( n9116 , n5877 , n11626 );
    or g14144 ( n1073 , n777 , n3433 );
    or g14145 ( n264 , n12016 , n17756 );
    nor g14146 ( n27178 , n7428 , n17169 );
    or g14147 ( n11716 , n8118 , n14359 );
    xnor g14148 ( n10484 , n18160 , n687 );
    not g14149 ( n17906 , n14265 );
    or g14150 ( n11505 , n24646 , n4288 );
    xnor g14151 ( n18859 , n18468 , n11639 );
    not g14152 ( n778 , n13044 );
    not g14153 ( n19340 , n22358 );
    or g14154 ( n612 , n25930 , n15940 );
    and g14155 ( n18775 , n23912 , n22716 );
    not g14156 ( n26218 , n7850 );
    xnor g14157 ( n16978 , n16468 , n12720 );
    xnor g14158 ( n18218 , n7070 , n21661 );
    nor g14159 ( n8150 , n17266 , n9151 );
    or g14160 ( n8386 , n14339 , n25705 );
    or g14161 ( n17580 , n10914 , n25014 );
    xnor g14162 ( n1555 , n7041 , n393 );
    or g14163 ( n16614 , n13443 , n13783 );
    not g14164 ( n5547 , n9598 );
    not g14165 ( n21999 , n15710 );
    xnor g14166 ( n10628 , n13937 , n10836 );
    xnor g14167 ( n18743 , n10411 , n8309 );
    or g14168 ( n3026 , n7119 , n14544 );
    or g14169 ( n21920 , n321 , n16577 );
    not g14170 ( n16267 , n10843 );
    xnor g14171 ( n863 , n2610 , n9406 );
    xnor g14172 ( n24599 , n13240 , n18897 );
    or g14173 ( n18543 , n4796 , n20828 );
    not g14174 ( n234 , n15977 );
    or g14175 ( n16161 , n22173 , n17932 );
    and g14176 ( n1455 , n26909 , n17618 );
    and g14177 ( n25705 , n2392 , n9061 );
    and g14178 ( n18696 , n6723 , n5370 );
    and g14179 ( n6374 , n171 , n15680 );
    and g14180 ( n16137 , n12738 , n10615 );
    xnor g14181 ( n12379 , n25422 , n6388 );
    xnor g14182 ( n17196 , n18643 , n15313 );
    not g14183 ( n12923 , n14704 );
    and g14184 ( n6913 , n11280 , n6479 );
    not g14185 ( n1009 , n19196 );
    xnor g14186 ( n19274 , n24051 , n18158 );
    not g14187 ( n5036 , n14391 );
    xnor g14188 ( n13752 , n8110 , n23691 );
    xnor g14189 ( n18919 , n18567 , n2164 );
    and g14190 ( n3656 , n6090 , n17429 );
    nor g14191 ( n11102 , n19110 , n10522 );
    or g14192 ( n12044 , n19152 , n22567 );
    or g14193 ( n13952 , n11125 , n22203 );
    or g14194 ( n23856 , n10084 , n4372 );
    nor g14195 ( n18914 , n17056 , n2109 );
    and g14196 ( n21840 , n9515 , n19559 );
    not g14197 ( n13893 , n8753 );
    and g14198 ( n1493 , n3064 , n22746 );
    not g14199 ( n22421 , n16290 );
    not g14200 ( n25572 , n649 );
    not g14201 ( n17230 , n6729 );
    xnor g14202 ( n8701 , n20056 , n11135 );
    or g14203 ( n9865 , n18344 , n2965 );
    not g14204 ( n21137 , n1097 );
    or g14205 ( n26393 , n20040 , n23983 );
    not g14206 ( n22912 , n3606 );
    and g14207 ( n745 , n26739 , n24046 );
    xnor g14208 ( n14878 , n24720 , n4175 );
    or g14209 ( n24677 , n1880 , n25227 );
    nor g14210 ( n21792 , n15077 , n24112 );
    nor g14211 ( n17017 , n23854 , n25533 );
    or g14212 ( n13064 , n24051 , n20989 );
    and g14213 ( n21830 , n3738 , n20193 );
    xnor g14214 ( n26905 , n21296 , n23229 );
    not g14215 ( n4922 , n13175 );
    and g14216 ( n25628 , n146 , n6832 );
    xnor g14217 ( n20104 , n21619 , n22974 );
    xnor g14218 ( n4259 , n814 , n4121 );
    nor g14219 ( n14572 , n19170 , n3608 );
    not g14220 ( n18847 , n8119 );
    or g14221 ( n1858 , n6267 , n18319 );
    not g14222 ( n4038 , n16291 );
    xnor g14223 ( n20723 , n14388 , n19892 );
    not g14224 ( n21977 , n19583 );
    or g14225 ( n4584 , n6373 , n13567 );
    or g14226 ( n17400 , n2903 , n22015 );
    xnor g14227 ( n5706 , n5047 , n9934 );
    or g14228 ( n16673 , n26086 , n19144 );
    xnor g14229 ( n5954 , n22539 , n6798 );
    or g14230 ( n17363 , n22403 , n22681 );
    not g14231 ( n18371 , n13844 );
    or g14232 ( n15460 , n3745 , n21074 );
    or g14233 ( n16865 , n10854 , n21969 );
    or g14234 ( n22801 , n8381 , n23775 );
    and g14235 ( n18555 , n26691 , n7563 );
    not g14236 ( n21867 , n20259 );
    and g14237 ( n22449 , n18423 , n19029 );
    or g14238 ( n10658 , n14899 , n23308 );
    nor g14239 ( n5037 , n2242 , n6449 );
    not g14240 ( n10513 , n18421 );
    and g14241 ( n21334 , n23563 , n21699 );
    or g14242 ( n12061 , n25690 , n7273 );
    or g14243 ( n2441 , n26062 , n25068 );
    or g14244 ( n7648 , n21107 , n4675 );
    xnor g14245 ( n15465 , n2204 , n20252 );
    xnor g14246 ( n4007 , n17752 , n8383 );
    xnor g14247 ( n24176 , n8771 , n7897 );
    or g14248 ( n3678 , n13977 , n15006 );
    nor g14249 ( n24310 , n3097 , n26667 );
    xnor g14250 ( n26605 , n14500 , n26784 );
    and g14251 ( n19480 , n26701 , n4233 );
    or g14252 ( n19508 , n5560 , n16944 );
    nor g14253 ( n26133 , n20923 , n5288 );
    not g14254 ( n16400 , n24485 );
    xnor g14255 ( n25631 , n4869 , n11317 );
    not g14256 ( n6831 , n14282 );
    or g14257 ( n10292 , n6104 , n19985 );
    or g14258 ( n10562 , n19962 , n12955 );
    and g14259 ( n9137 , n680 , n4948 );
    or g14260 ( n5314 , n6352 , n21288 );
    nor g14261 ( n15338 , n3570 , n575 );
    xnor g14262 ( n21504 , n3506 , n9934 );
    or g14263 ( n8442 , n9396 , n11817 );
    not g14264 ( n9944 , n25471 );
    nor g14265 ( n11456 , n5495 , n9366 );
    or g14266 ( n19506 , n3260 , n20512 );
    not g14267 ( n25930 , n13190 );
    xnor g14268 ( n10390 , n19290 , n20872 );
    and g14269 ( n27155 , n15489 , n6471 );
    and g14270 ( n24509 , n23741 , n12977 );
    or g14271 ( n14270 , n24276 , n578 );
    buf g14272 ( n4542 , n1238 );
    or g14273 ( n21310 , n20032 , n19227 );
    nor g14274 ( n22978 , n15534 , n25572 );
    xnor g14275 ( n27017 , n14183 , n11509 );
    not g14276 ( n3967 , n15521 );
    and g14277 ( n19848 , n16427 , n1807 );
    nor g14278 ( n11380 , n17230 , n3447 );
    or g14279 ( n9330 , n7581 , n16933 );
    and g14280 ( n10848 , n3368 , n23531 );
    nor g14281 ( n12485 , n9399 , n9507 );
    nor g14282 ( n16575 , n5451 , n3918 );
    and g14283 ( n13252 , n831 , n5871 );
    or g14284 ( n17849 , n23603 , n9720 );
    or g14285 ( n22623 , n3734 , n10487 );
    and g14286 ( n20721 , n7457 , n32 );
    xnor g14287 ( n2697 , n725 , n7759 );
    and g14288 ( n4068 , n20246 , n6017 );
    or g14289 ( n26763 , n15380 , n22576 );
    and g14290 ( n21724 , n3457 , n15181 );
    not g14291 ( n5417 , n7376 );
    xnor g14292 ( n12931 , n1759 , n25331 );
    or g14293 ( n3773 , n286 , n13379 );
    xnor g14294 ( n4929 , n26529 , n17204 );
    or g14295 ( n6604 , n7561 , n2849 );
    or g14296 ( n13052 , n24004 , n21081 );
    and g14297 ( n4246 , n22297 , n1633 );
    not g14298 ( n6239 , n24425 );
    xnor g14299 ( n1869 , n22281 , n8537 );
    xnor g14300 ( n13473 , n21288 , n25238 );
    and g14301 ( n22539 , n15632 , n5278 );
    or g14302 ( n5152 , n698 , n18404 );
    or g14303 ( n2351 , n26056 , n9314 );
    not g14304 ( n11551 , n20001 );
    xnor g14305 ( n8214 , n5506 , n20923 );
    or g14306 ( n25275 , n25837 , n5481 );
    or g14307 ( n5315 , n11144 , n12702 );
    or g14308 ( n25662 , n4691 , n4988 );
    and g14309 ( n12008 , n1795 , n10824 );
    not g14310 ( n27107 , n22465 );
    or g14311 ( n13946 , n25643 , n27141 );
    and g14312 ( n24619 , n20914 , n4528 );
    xnor g14313 ( n11161 , n6825 , n21498 );
    or g14314 ( n7381 , n11903 , n14872 );
    and g14315 ( n9619 , n23702 , n1038 );
    xnor g14316 ( n7216 , n25537 , n14971 );
    or g14317 ( n9959 , n17151 , n3572 );
    or g14318 ( n7964 , n13862 , n23976 );
    or g14319 ( n4078 , n3217 , n3746 );
    and g14320 ( n27171 , n16188 , n1566 );
    or g14321 ( n1766 , n12143 , n1351 );
    and g14322 ( n15166 , n7936 , n2962 );
    and g14323 ( n4790 , n16488 , n5725 );
    or g14324 ( n14582 , n15022 , n13125 );
    not g14325 ( n2090 , n18302 );
    or g14326 ( n3273 , n5183 , n4448 );
    xnor g14327 ( n12529 , n19116 , n3945 );
    and g14328 ( n6950 , n7935 , n11552 );
    xnor g14329 ( n8165 , n19194 , n14805 );
    and g14330 ( n11114 , n26241 , n918 );
    nor g14331 ( n13351 , n22358 , n9597 );
    xnor g14332 ( n15470 , n27123 , n6884 );
    nor g14333 ( n9740 , n15405 , n2223 );
    not g14334 ( n10251 , n693 );
    or g14335 ( n21282 , n9779 , n20205 );
    xnor g14336 ( n7391 , n23193 , n14154 );
    or g14337 ( n26376 , n8298 , n5124 );
    nor g14338 ( n12442 , n9671 , n19042 );
    xnor g14339 ( n81 , n9246 , n7876 );
    or g14340 ( n25583 , n21467 , n23870 );
    xnor g14341 ( n19568 , n24082 , n11447 );
    not g14342 ( n4083 , n10320 );
    xnor g14343 ( n10590 , n15584 , n21030 );
    or g14344 ( n25187 , n6764 , n8344 );
    nor g14345 ( n13546 , n16016 , n14365 );
    not g14346 ( n24371 , n2139 );
    and g14347 ( n1359 , n16476 , n19 );
    or g14348 ( n7961 , n6262 , n18975 );
    xnor g14349 ( n6885 , n13333 , n9512 );
    nor g14350 ( n22116 , n2045 , n19228 );
    xnor g14351 ( n9376 , n23404 , n7753 );
    xnor g14352 ( n1117 , n25643 , n20604 );
    not g14353 ( n8162 , n22282 );
    xnor g14354 ( n24281 , n17162 , n17147 );
    nor g14355 ( n19260 , n18814 , n25471 );
    xnor g14356 ( n17928 , n27084 , n19696 );
    nor g14357 ( n24662 , n5715 , n20554 );
    nor g14358 ( n19000 , n27188 , n4326 );
    and g14359 ( n18048 , n10889 , n6696 );
    xnor g14360 ( n24853 , n15609 , n1560 );
    and g14361 ( n15978 , n16180 , n19463 );
    xnor g14362 ( n26872 , n204 , n14704 );
    or g14363 ( n1517 , n21128 , n13252 );
    xnor g14364 ( n2990 , n22332 , n7751 );
    not g14365 ( n5746 , n11932 );
    nor g14366 ( n5068 , n11740 , n3591 );
    xnor g14367 ( n26754 , n21749 , n919 );
    xnor g14368 ( n21328 , n6734 , n19404 );
    not g14369 ( n13913 , n5208 );
    or g14370 ( n7628 , n22975 , n18144 );
    xnor g14371 ( n8441 , n26021 , n4984 );
    and g14372 ( n14505 , n14604 , n2851 );
    not g14373 ( n20393 , n14156 );
    xnor g14374 ( n25173 , n5708 , n1181 );
    or g14375 ( n9501 , n6229 , n7212 );
    or g14376 ( n15159 , n23198 , n10822 );
    and g14377 ( n17499 , n12618 , n7595 );
    xnor g14378 ( n145 , n23509 , n7731 );
    not g14379 ( n12262 , n6359 );
    or g14380 ( n25134 , n2125 , n20829 );
    or g14381 ( n11748 , n5512 , n18962 );
    xnor g14382 ( n5360 , n21200 , n18549 );
    and g14383 ( n6395 , n17664 , n21253 );
    and g14384 ( n8160 , n2917 , n3771 );
    and g14385 ( n4016 , n2605 , n3683 );
    not g14386 ( n23242 , n4391 );
    or g14387 ( n13047 , n19513 , n22137 );
    not g14388 ( n21469 , n7391 );
    nor g14389 ( n8345 , n5043 , n18133 );
    or g14390 ( n15561 , n902 , n19620 );
    not g14391 ( n24552 , n13708 );
    or g14392 ( n16757 , n11377 , n16611 );
    or g14393 ( n2661 , n25981 , n27003 );
    or g14394 ( n11154 , n14814 , n6419 );
    xnor g14395 ( n1510 , n516 , n10020 );
    xnor g14396 ( n2568 , n226 , n18544 );
    not g14397 ( n8980 , n13250 );
    and g14398 ( n25132 , n18765 , n4659 );
    or g14399 ( n22145 , n16880 , n18357 );
    xnor g14400 ( n6354 , n13218 , n17472 );
    and g14401 ( n488 , n25586 , n8491 );
    or g14402 ( n15802 , n11449 , n26154 );
    xnor g14403 ( n24989 , n4086 , n8724 );
    not g14404 ( n8572 , n4708 );
    xnor g14405 ( n23007 , n20979 , n10779 );
    or g14406 ( n17326 , n7305 , n830 );
    and g14407 ( n8364 , n16563 , n9334 );
    xnor g14408 ( n15411 , n4641 , n7746 );
    and g14409 ( n24251 , n25078 , n3023 );
    xnor g14410 ( n25468 , n21011 , n16299 );
    or g14411 ( n9248 , n8256 , n17815 );
    or g14412 ( n4983 , n21 , n23513 );
    xnor g14413 ( n7558 , n20540 , n26126 );
    buf g14414 ( n593 , n13220 );
    not g14415 ( n10441 , n5182 );
    and g14416 ( n16921 , n20650 , n4968 );
    and g14417 ( n26586 , n21581 , n14741 );
    xnor g14418 ( n9979 , n23333 , n16502 );
    not g14419 ( n19255 , n25659 );
    or g14420 ( n13720 , n25237 , n13336 );
    not g14421 ( n23329 , n14661 );
    and g14422 ( n11371 , n21583 , n16756 );
    xnor g14423 ( n11128 , n4613 , n10076 );
    or g14424 ( n20122 , n26596 , n6399 );
    xnor g14425 ( n13491 , n13494 , n3425 );
    nor g14426 ( n24892 , n21471 , n24612 );
    and g14427 ( n19171 , n13026 , n13906 );
    or g14428 ( n16075 , n27048 , n24530 );
    and g14429 ( n2166 , n19097 , n5333 );
    or g14430 ( n20987 , n10373 , n25082 );
    or g14431 ( n27141 , n9557 , n21944 );
    xnor g14432 ( n2534 , n8195 , n19935 );
    not g14433 ( n4591 , n3214 );
    xnor g14434 ( n7573 , n1705 , n5354 );
    or g14435 ( n2471 , n1106 , n26770 );
    or g14436 ( n20193 , n4996 , n26669 );
    and g14437 ( n16518 , n22111 , n13971 );
    xnor g14438 ( n16841 , n7637 , n3377 );
    or g14439 ( n20677 , n14171 , n16739 );
    and g14440 ( n24613 , n23647 , n24465 );
    or g14441 ( n19878 , n23773 , n9358 );
    xnor g14442 ( n14888 , n3606 , n7484 );
    and g14443 ( n20543 , n8843 , n9071 );
    xnor g14444 ( n8505 , n8157 , n22899 );
    xnor g14445 ( n15846 , n24628 , n9322 );
    xnor g14446 ( n14706 , n16058 , n18532 );
    xnor g14447 ( n2615 , n26260 , n4139 );
    xnor g14448 ( n11682 , n11969 , n7302 );
    and g14449 ( n16748 , n1009 , n4999 );
    or g14450 ( n5671 , n20988 , n26955 );
    nor g14451 ( n3856 , n7008 , n25810 );
    and g14452 ( n10462 , n11311 , n12903 );
    or g14453 ( n26593 , n13591 , n3909 );
    or g14454 ( n14709 , n25326 , n17752 );
    xnor g14455 ( n25166 , n7670 , n3253 );
    or g14456 ( n3401 , n19032 , n23802 );
    or g14457 ( n19407 , n13408 , n2450 );
    or g14458 ( n18529 , n14625 , n2210 );
    xnor g14459 ( n22091 , n13852 , n4009 );
    or g14460 ( n20395 , n3315 , n6214 );
    xnor g14461 ( n9626 , n14021 , n14202 );
    or g14462 ( n7458 , n22666 , n18148 );
    xnor g14463 ( n15815 , n2182 , n12814 );
    or g14464 ( n9481 , n19624 , n14625 );
    xnor g14465 ( n20967 , n15266 , n3506 );
    or g14466 ( n1990 , n7623 , n16736 );
    not g14467 ( n12547 , n18905 );
    not g14468 ( n22515 , n13220 );
    and g14469 ( n15048 , n26757 , n12504 );
    or g14470 ( n11666 , n1896 , n11457 );
    and g14471 ( n10721 , n7496 , n12151 );
    and g14472 ( n9023 , n8338 , n3967 );
    or g14473 ( n10726 , n17836 , n9684 );
    and g14474 ( n18387 , n26560 , n9272 );
    nor g14475 ( n11179 , n401 , n14519 );
    not g14476 ( n10274 , n23369 );
    xnor g14477 ( n9452 , n25739 , n26443 );
    and g14478 ( n20241 , n17062 , n21906 );
    or g14479 ( n16894 , n16261 , n23013 );
    and g14480 ( n25902 , n19387 , n1395 );
    xnor g14481 ( n6219 , n19303 , n8782 );
    or g14482 ( n26646 , n8416 , n101 );
    xnor g14483 ( n11803 , n16261 , n24188 );
    xnor g14484 ( n19247 , n9562 , n19409 );
    xnor g14485 ( n26189 , n215 , n14702 );
    or g14486 ( n5125 , n24686 , n9889 );
    and g14487 ( n5648 , n19197 , n26099 );
    or g14488 ( n21515 , n22411 , n3951 );
    or g14489 ( n1732 , n1242 , n21031 );
    not g14490 ( n17645 , n5521 );
    xor g14491 ( n27197 , n25405 , n20406 );
    or g14492 ( n4881 , n5767 , n23435 );
    not g14493 ( n15073 , n20505 );
    or g14494 ( n4998 , n21905 , n24481 );
    and g14495 ( n7036 , n16655 , n3339 );
    or g14496 ( n9001 , n19427 , n18500 );
    xnor g14497 ( n25592 , n13352 , n2233 );
    and g14498 ( n5059 , n13782 , n9568 );
    not g14499 ( n2048 , n7924 );
    xnor g14500 ( n8817 , n12125 , n25327 );
    xnor g14501 ( n6107 , n24851 , n12495 );
    or g14502 ( n2172 , n12513 , n14106 );
    or g14503 ( n21583 , n9180 , n2514 );
    or g14504 ( n20816 , n23788 , n4249 );
    xnor g14505 ( n17855 , n1818 , n13557 );
    xnor g14506 ( n11439 , n3360 , n26006 );
    xnor g14507 ( n24320 , n11930 , n1277 );
    xnor g14508 ( n2826 , n5241 , n1177 );
    xnor g14509 ( n2422 , n14462 , n5784 );
    xnor g14510 ( n12920 , n25991 , n1840 );
    not g14511 ( n25007 , n23187 );
    or g14512 ( n2945 , n2099 , n21948 );
    not g14513 ( n10749 , n9413 );
    xnor g14514 ( n10750 , n24645 , n13714 );
    not g14515 ( n26498 , n5450 );
    nor g14516 ( n12686 , n15693 , n21626 );
    nor g14517 ( n15974 , n12068 , n4558 );
    xnor g14518 ( n5111 , n15414 , n23610 );
    nor g14519 ( n5331 , n25007 , n19048 );
    not g14520 ( n20796 , n8079 );
    and g14521 ( n1045 , n17631 , n24068 );
    not g14522 ( n5530 , n1344 );
    not g14523 ( n17350 , n22456 );
    or g14524 ( n6097 , n6613 , n8933 );
    or g14525 ( n19219 , n13528 , n12373 );
    and g14526 ( n7289 , n681 , n18491 );
    and g14527 ( n4250 , n23438 , n7603 );
    nor g14528 ( n15864 , n1536 , n21743 );
    not g14529 ( n11453 , n23026 );
    or g14530 ( n5087 , n22740 , n24169 );
    xnor g14531 ( n890 , n17605 , n25533 );
    xnor g14532 ( n10605 , n5934 , n7776 );
    xnor g14533 ( n6822 , n17716 , n14704 );
    xnor g14534 ( n18628 , n18452 , n1752 );
    xnor g14535 ( n13202 , n972 , n11155 );
    xnor g14536 ( n4464 , n13489 , n20575 );
    and g14537 ( n22647 , n15075 , n19800 );
    not g14538 ( n959 , n9966 );
    and g14539 ( n23191 , n21801 , n15597 );
    or g14540 ( n3998 , n13392 , n23394 );
    or g14541 ( n26494 , n19277 , n13963 );
    or g14542 ( n15181 , n18209 , n8047 );
    or g14543 ( n15086 , n11069 , n6743 );
    or g14544 ( n7304 , n17439 , n24966 );
    not g14545 ( n19028 , n19786 );
    not g14546 ( n21896 , n22634 );
    nor g14547 ( n3256 , n3809 , n8406 );
    and g14548 ( n16432 , n1715 , n19371 );
    xnor g14549 ( n5927 , n7153 , n15325 );
    and g14550 ( n17105 , n9713 , n1471 );
    or g14551 ( n13334 , n15900 , n15351 );
    xnor g14552 ( n21726 , n3184 , n7209 );
    not g14553 ( n17483 , n7436 );
    or g14554 ( n2733 , n20642 , n22932 );
    or g14555 ( n6889 , n12453 , n2908 );
    xnor g14556 ( n631 , n8786 , n25381 );
    and g14557 ( n8785 , n16998 , n10134 );
    not g14558 ( n3015 , n5701 );
    xnor g14559 ( n14421 , n3861 , n6631 );
    xnor g14560 ( n21629 , n20043 , n20986 );
    or g14561 ( n23946 , n740 , n14318 );
    xnor g14562 ( n19070 , n17605 , n4263 );
    or g14563 ( n14068 , n16464 , n4844 );
    nor g14564 ( n12655 , n3405 , n24165 );
    not g14565 ( n1882 , n12754 );
    xnor g14566 ( n4175 , n16812 , n25923 );
    not g14567 ( n4307 , n17159 );
    xnor g14568 ( n18065 , n16077 , n26300 );
    xnor g14569 ( n8306 , n12721 , n13465 );
    or g14570 ( n5877 , n8773 , n11657 );
    xnor g14571 ( n14361 , n24246 , n14883 );
    xnor g14572 ( n18036 , n16993 , n24601 );
    nor g14573 ( n22089 , n23849 , n19702 );
    nor g14574 ( n19439 , n2995 , n15678 );
    xnor g14575 ( n27070 , n575 , n22198 );
    nor g14576 ( n18101 , n11378 , n22110 );
    xnor g14577 ( n25614 , n11383 , n16859 );
    xnor g14578 ( n15303 , n21071 , n8945 );
    xnor g14579 ( n11903 , n10808 , n3077 );
    buf g14580 ( n15767 , n271 );
    not g14581 ( n23050 , n4115 );
    and g14582 ( n19609 , n10169 , n7133 );
    or g14583 ( n6539 , n17005 , n12117 );
    xnor g14584 ( n17791 , n8006 , n19514 );
    or g14585 ( n26083 , n10265 , n241 );
    xnor g14586 ( n19396 , n1336 , n3843 );
    or g14587 ( n12982 , n10003 , n8929 );
    not g14588 ( n9574 , n6658 );
    xnor g14589 ( n117 , n11209 , n5495 );
    not g14590 ( n18700 , n26608 );
    and g14591 ( n20910 , n14146 , n2437 );
    and g14592 ( n20255 , n11357 , n10286 );
    nor g14593 ( n12218 , n13190 , n9318 );
    and g14594 ( n18308 , n6338 , n3070 );
    xnor g14595 ( n11138 , n264 , n1261 );
    xnor g14596 ( n17998 , n14159 , n5770 );
    xnor g14597 ( n18909 , n22226 , n23430 );
    and g14598 ( n11540 , n7062 , n14349 );
    xnor g14599 ( n5841 , n24971 , n9687 );
    not g14600 ( n27199 , n17959 );
    or g14601 ( n12392 , n19297 , n24042 );
    xnor g14602 ( n4026 , n20196 , n26748 );
    nor g14603 ( n11033 , n20032 , n25974 );
    or g14604 ( n1515 , n6764 , n6611 );
    or g14605 ( n9769 , n12122 , n19320 );
    or g14606 ( n14332 , n12468 , n22224 );
    and g14607 ( n16581 , n21019 , n10433 );
    xnor g14608 ( n3483 , n23729 , n22597 );
    xnor g14609 ( n735 , n5227 , n2140 );
    or g14610 ( n21012 , n25334 , n18978 );
    or g14611 ( n92 , n5077 , n12739 );
    and g14612 ( n9755 , n18504 , n17483 );
    or g14613 ( n397 , n13757 , n25654 );
    xnor g14614 ( n10199 , n23292 , n11423 );
    xnor g14615 ( n4172 , n7611 , n6342 );
    xnor g14616 ( n23551 , n2057 , n21930 );
    nor g14617 ( n11732 , n7305 , n23061 );
    or g14618 ( n15606 , n25897 , n17573 );
    xnor g14619 ( n13794 , n8285 , n20036 );
    xnor g14620 ( n22391 , n21450 , n24821 );
    or g14621 ( n600 , n20393 , n26832 );
    or g14622 ( n2548 , n26572 , n4029 );
    or g14623 ( n7203 , n505 , n9748 );
    xnor g14624 ( n463 , n11437 , n13740 );
    not g14625 ( n3949 , n1543 );
    xnor g14626 ( n9002 , n9940 , n11455 );
    xnor g14627 ( n17972 , n21824 , n15820 );
    xnor g14628 ( n13732 , n20365 , n14127 );
    xnor g14629 ( n3298 , n17005 , n25303 );
    xnor g14630 ( n8226 , n23032 , n22863 );
    and g14631 ( n19381 , n5723 , n6324 );
    xnor g14632 ( n20102 , n7659 , n7031 );
    xnor g14633 ( n2950 , n2206 , n24412 );
    xnor g14634 ( n23767 , n20526 , n24139 );
    or g14635 ( n17916 , n8943 , n9683 );
    and g14636 ( n3636 , n24972 , n5429 );
    xnor g14637 ( n13698 , n24125 , n20639 );
    xnor g14638 ( n18545 , n14158 , n5140 );
    not g14639 ( n22365 , n12587 );
    xnor g14640 ( n19137 , n4096 , n22778 );
    xnor g14641 ( n7496 , n11722 , n1316 );
    xnor g14642 ( n492 , n21420 , n9820 );
    not g14643 ( n11603 , n863 );
    or g14644 ( n202 , n17701 , n10531 );
    xnor g14645 ( n6495 , n23865 , n19200 );
    or g14646 ( n17988 , n22074 , n15484 );
    and g14647 ( n5132 , n17212 , n14634 );
    xnor g14648 ( n19103 , n17762 , n22433 );
    nor g14649 ( n8538 , n22964 , n21060 );
    or g14650 ( n11709 , n7328 , n20493 );
    buf g14651 ( n26344 , n24873 );
    or g14652 ( n1769 , n25139 , n1794 );
    xnor g14653 ( n4956 , n8201 , n20317 );
    not g14654 ( n2208 , n2221 );
    xnor g14655 ( n25996 , n21378 , n25972 );
    and g14656 ( n21913 , n15782 , n14334 );
    or g14657 ( n5393 , n26957 , n18662 );
    or g14658 ( n24107 , n604 , n4626 );
    xnor g14659 ( n4736 , n22597 , n18901 );
    and g14660 ( n19375 , n6750 , n13328 );
    and g14661 ( n10335 , n6894 , n2894 );
    and g14662 ( n3043 , n8568 , n13140 );
    or g14663 ( n12176 , n3091 , n26031 );
    and g14664 ( n9610 , n13225 , n10115 );
    and g14665 ( n22545 , n2915 , n23559 );
    and g14666 ( n19350 , n22626 , n25038 );
    xnor g14667 ( n677 , n9052 , n4982 );
    or g14668 ( n16826 , n19944 , n1451 );
    xnor g14669 ( n17405 , n20077 , n22433 );
    xnor g14670 ( n6164 , n1093 , n3718 );
    nor g14671 ( n18216 , n832 , n23506 );
    and g14672 ( n4114 , n10005 , n12691 );
    xnor g14673 ( n7636 , n25089 , n11721 );
    or g14674 ( n21305 , n19074 , n8581 );
    xnor g14675 ( n16182 , n3239 , n1464 );
    xnor g14676 ( n9575 , n24920 , n26806 );
    and g14677 ( n20953 , n15674 , n17270 );
    and g14678 ( n2913 , n3081 , n19512 );
    nor g14679 ( n4539 , n22198 , n8774 );
    xnor g14680 ( n14180 , n8964 , n1293 );
    or g14681 ( n2836 , n16874 , n18589 );
    nor g14682 ( n22845 , n7149 , n22871 );
    or g14683 ( n14031 , n25345 , n18479 );
    xnor g14684 ( n15975 , n4485 , n19906 );
    or g14685 ( n4839 , n9050 , n16210 );
    or g14686 ( n17878 , n23493 , n8405 );
    or g14687 ( n10641 , n16822 , n23329 );
    not g14688 ( n20249 , n23034 );
    xnor g14689 ( n24911 , n25171 , n3577 );
    and g14690 ( n7414 , n9779 , n24663 );
    xnor g14691 ( n24154 , n20649 , n15565 );
    xnor g14692 ( n3265 , n22782 , n24455 );
    xnor g14693 ( n22404 , n16676 , n16612 );
    or g14694 ( n26645 , n21674 , n5791 );
    and g14695 ( n18987 , n7953 , n20908 );
    not g14696 ( n17572 , n10897 );
    or g14697 ( n17745 , n21232 , n7471 );
    and g14698 ( n18645 , n18306 , n3303 );
    xnor g14699 ( n19625 , n18107 , n10859 );
    xnor g14700 ( n16900 , n14332 , n3662 );
    xnor g14701 ( n27117 , n19962 , n15508 );
    xnor g14702 ( n3649 , n11532 , n8375 );
    xnor g14703 ( n3726 , n111 , n17940 );
    not g14704 ( n19201 , n9246 );
    or g14705 ( n15069 , n12751 , n24847 );
    xnor g14706 ( n22669 , n9394 , n6039 );
    or g14707 ( n7982 , n24130 , n16531 );
    xnor g14708 ( n17679 , n21007 , n3018 );
    and g14709 ( n8156 , n9210 , n2729 );
    nor g14710 ( n22265 , n14158 , n11381 );
    not g14711 ( n20964 , n2289 );
    and g14712 ( n2951 , n1650 , n3272 );
    and g14713 ( n10268 , n21837 , n25845 );
    or g14714 ( n17776 , n5025 , n12771 );
    not g14715 ( n7906 , n17808 );
    not g14716 ( n22069 , n11006 );
    xnor g14717 ( n2324 , n13867 , n1922 );
    or g14718 ( n12943 , n11924 , n13072 );
    nor g14719 ( n24963 , n11824 , n14152 );
    nor g14720 ( n22868 , n26054 , n21907 );
    xnor g14721 ( n18679 , n18396 , n16923 );
    nor g14722 ( n18067 , n626 , n21772 );
    and g14723 ( n1070 , n16307 , n14742 );
    or g14724 ( n639 , n3346 , n8044 );
    nor g14725 ( n25868 , n755 , n23366 );
    and g14726 ( n26012 , n5314 , n25878 );
    or g14727 ( n18813 , n15489 , n6471 );
    and g14728 ( n25064 , n11279 , n6336 );
    or g14729 ( n16530 , n20998 , n22281 );
    not g14730 ( n676 , n1741 );
    and g14731 ( n10113 , n2219 , n8059 );
    and g14732 ( n1489 , n14392 , n18164 );
    and g14733 ( n14061 , n8780 , n3154 );
    xnor g14734 ( n3436 , n12049 , n10464 );
    and g14735 ( n15475 , n18176 , n25847 );
    xnor g14736 ( n298 , n14912 , n4989 );
    and g14737 ( n21185 , n24672 , n12748 );
    not g14738 ( n13360 , n24969 );
    or g14739 ( n14377 , n16787 , n7115 );
    buf g14740 ( n23878 , n8988 );
    or g14741 ( n23576 , n17937 , n11253 );
    and g14742 ( n17933 , n23895 , n8491 );
    xnor g14743 ( n2343 , n8397 , n23872 );
    and g14744 ( n6112 , n11946 , n24033 );
    nor g14745 ( n23530 , n1568 , n24571 );
    and g14746 ( n16616 , n27084 , n11307 );
    or g14747 ( n16671 , n14800 , n13824 );
    xnor g14748 ( n12059 , n5143 , n9040 );
    xnor g14749 ( n3261 , n24919 , n21915 );
    and g14750 ( n20251 , n19488 , n18355 );
    or g14751 ( n16557 , n4764 , n6043 );
    or g14752 ( n5565 , n10067 , n12818 );
    not g14753 ( n15644 , n5001 );
    nor g14754 ( n25551 , n16246 , n21119 );
    and g14755 ( n18253 , n10406 , n8947 );
    not g14756 ( n18930 , n22070 );
    nor g14757 ( n24089 , n3839 , n21774 );
    and g14758 ( n3691 , n7625 , n17785 );
    xnor g14759 ( n7755 , n6777 , n17362 );
    xnor g14760 ( n9891 , n10951 , n8794 );
    not g14761 ( n11211 , n14907 );
    nor g14762 ( n9157 , n18345 , n25168 );
    or g14763 ( n19026 , n2382 , n22169 );
    xnor g14764 ( n8376 , n5359 , n19912 );
    and g14765 ( n9397 , n23925 , n16964 );
    and g14766 ( n2753 , n17434 , n16737 );
    not g14767 ( n8008 , n8679 );
    nor g14768 ( n6970 , n7150 , n22062 );
    xnor g14769 ( n6514 , n10103 , n8274 );
    not g14770 ( n27200 , n17845 );
    nor g14771 ( n26145 , n5783 , n6682 );
    and g14772 ( n5415 , n24550 , n22182 );
    xnor g14773 ( n22031 , n11625 , n13959 );
    or g14774 ( n9153 , n24587 , n13597 );
    and g14775 ( n16535 , n24710 , n16431 );
    xnor g14776 ( n25696 , n15143 , n6527 );
    nor g14777 ( n12894 , n15153 , n9340 );
    and g14778 ( n26236 , n14322 , n8726 );
    or g14779 ( n16974 , n25863 , n23626 );
    xnor g14780 ( n7536 , n14144 , n17478 );
    or g14781 ( n13100 , n25886 , n19005 );
    and g14782 ( n19784 , n19651 , n6298 );
    or g14783 ( n10477 , n10815 , n2655 );
    xnor g14784 ( n8717 , n16631 , n17395 );
    nor g14785 ( n40 , n24211 , n8304 );
    xnor g14786 ( n23131 , n1654 , n16482 );
    not g14787 ( n4792 , n17870 );
    xnor g14788 ( n24096 , n21484 , n26639 );
    nor g14789 ( n19004 , n6200 , n6672 );
    or g14790 ( n1475 , n1477 , n3957 );
    or g14791 ( n25206 , n5471 , n2864 );
    xnor g14792 ( n3414 , n5801 , n1004 );
    or g14793 ( n19815 , n20112 , n23746 );
    xnor g14794 ( n16527 , n18741 , n3265 );
    or g14795 ( n22115 , n9180 , n18754 );
    xnor g14796 ( n26915 , n17057 , n27049 );
    xnor g14797 ( n11047 , n26697 , n24439 );
    or g14798 ( n26843 , n26551 , n22035 );
    and g14799 ( n9390 , n11450 , n3489 );
    not g14800 ( n1318 , n14767 );
    and g14801 ( n25668 , n14899 , n18496 );
    xnor g14802 ( n10867 , n25413 , n1293 );
    xnor g14803 ( n11584 , n22715 , n10023 );
    not g14804 ( n2477 , n12541 );
    not g14805 ( n1803 , n26405 );
    or g14806 ( n12703 , n13453 , n4434 );
    or g14807 ( n10399 , n18428 , n16793 );
    xnor g14808 ( n22756 , n14139 , n9358 );
    xnor g14809 ( n6585 , n2244 , n543 );
    or g14810 ( n11528 , n11211 , n13774 );
    xnor g14811 ( n25489 , n15894 , n24378 );
    nor g14812 ( n5146 , n17381 , n23731 );
    or g14813 ( n25988 , n6647 , n9457 );
    nor g14814 ( n10036 , n24578 , n15417 );
    and g14815 ( n22040 , n9598 , n19084 );
    not g14816 ( n19051 , n19625 );
    and g14817 ( n25921 , n1262 , n1084 );
    and g14818 ( n12116 , n13190 , n21632 );
    and g14819 ( n8168 , n15533 , n18839 );
    nor g14820 ( n23121 , n9832 , n3959 );
    or g14821 ( n3475 , n5745 , n25073 );
    not g14822 ( n5112 , n12211 );
    not g14823 ( n24650 , n22597 );
    and g14824 ( n10465 , n16225 , n4680 );
    xnor g14825 ( n10629 , n901 , n8258 );
    or g14826 ( n2710 , n6202 , n2366 );
    or g14827 ( n26446 , n475 , n10517 );
    and g14828 ( n8047 , n1276 , n5311 );
    and g14829 ( n12885 , n3517 , n15377 );
    and g14830 ( n11568 , n21803 , n13768 );
    or g14831 ( n14890 , n1006 , n6531 );
    or g14832 ( n17535 , n6946 , n8485 );
    not g14833 ( n1000 , n3903 );
    xnor g14834 ( n13774 , n24270 , n17958 );
    or g14835 ( n22938 , n12167 , n13956 );
    nor g14836 ( n7175 , n24208 , n2423 );
    xnor g14837 ( n10271 , n23097 , n14749 );
    or g14838 ( n3105 , n280 , n16214 );
    or g14839 ( n6314 , n17562 , n16804 );
    xnor g14840 ( n23967 , n8650 , n20826 );
    not g14841 ( n7925 , n10460 );
    nor g14842 ( n18892 , n8087 , n14795 );
    not g14843 ( n26501 , n24592 );
    not g14844 ( n26162 , n27089 );
    or g14845 ( n13331 , n20435 , n10085 );
    nor g14846 ( n1825 , n16257 , n6861 );
    xnor g14847 ( n21168 , n16220 , n4774 );
    xnor g14848 ( n3509 , n18358 , n14206 );
    xnor g14849 ( n6335 , n7371 , n7438 );
    nor g14850 ( n15302 , n4659 , n1835 );
    not g14851 ( n4800 , n15719 );
    nor g14852 ( n10066 , n1236 , n23717 );
    nor g14853 ( n9800 , n2341 , n6596 );
    and g14854 ( n4783 , n21389 , n413 );
    or g14855 ( n22698 , n24941 , n3961 );
    not g14856 ( n22655 , n13387 );
    xnor g14857 ( n12323 , n17599 , n665 );
    xnor g14858 ( n9792 , n21948 , n26805 );
    or g14859 ( n11237 , n644 , n12868 );
    and g14860 ( n18613 , n24791 , n2291 );
    not g14861 ( n24301 , n20946 );
    and g14862 ( n25546 , n12154 , n12103 );
    and g14863 ( n25595 , n23074 , n26395 );
    and g14864 ( n24574 , n5451 , n1533 );
    xnor g14865 ( n9004 , n18968 , n18753 );
    or g14866 ( n13374 , n22202 , n19983 );
    not g14867 ( n11312 , n15268 );
    and g14868 ( n14331 , n5852 , n16963 );
    xnor g14869 ( n2030 , n17578 , n4085 );
    xnor g14870 ( n22175 , n10833 , n9378 );
    and g14871 ( n26004 , n26003 , n20166 );
    xnor g14872 ( n16093 , n8994 , n14510 );
    and g14873 ( n9361 , n1293 , n15921 );
    or g14874 ( n17019 , n540 , n9342 );
    xnor g14875 ( n15383 , n6977 , n23096 );
    xnor g14876 ( n9897 , n7009 , n4300 );
    nor g14877 ( n3545 , n8964 , n22554 );
    not g14878 ( n4022 , n21317 );
    or g14879 ( n7620 , n13311 , n17332 );
    xnor g14880 ( n19040 , n9935 , n22841 );
    nor g14881 ( n15054 , n12380 , n16638 );
    nor g14882 ( n4615 , n13842 , n23670 );
    and g14883 ( n17709 , n9275 , n25597 );
    or g14884 ( n17123 , n13190 , n23999 );
    xnor g14885 ( n12746 , n13528 , n4417 );
    xnor g14886 ( n3758 , n5864 , n14587 );
    xnor g14887 ( n19835 , n7671 , n197 );
    or g14888 ( n5762 , n14933 , n17386 );
    not g14889 ( n21868 , n21912 );
    xnor g14890 ( n18319 , n2541 , n1722 );
    not g14891 ( n20733 , n8439 );
    xnor g14892 ( n25211 , n22660 , n21753 );
    or g14893 ( n10115 , n381 , n24356 );
    not g14894 ( n13309 , n19911 );
    not g14895 ( n26047 , n17200 );
    or g14896 ( n17732 , n22895 , n17203 );
    xnor g14897 ( n13018 , n25042 , n7421 );
    xnor g14898 ( n1052 , n3780 , n5075 );
    or g14899 ( n18552 , n5498 , n16544 );
    xnor g14900 ( n3080 , n16713 , n17497 );
    xnor g14901 ( n20431 , n3203 , n21272 );
    xnor g14902 ( n26564 , n19753 , n16369 );
    or g14903 ( n11663 , n23328 , n11117 );
    and g14904 ( n20242 , n3260 , n21832 );
    not g14905 ( n11755 , n4485 );
    and g14906 ( n21116 , n1902 , n15441 );
    not g14907 ( n24493 , n7536 );
    or g14908 ( n11311 , n3099 , n23418 );
    and g14909 ( n1125 , n24544 , n21167 );
    xnor g14910 ( n385 , n20455 , n5376 );
    not g14911 ( n17613 , n5817 );
    and g14912 ( n10417 , n17004 , n24496 );
    nor g14913 ( n24772 , n10773 , n13460 );
    and g14914 ( n26952 , n8860 , n4313 );
    xnor g14915 ( n23684 , n19538 , n17227 );
    or g14916 ( n13173 , n5790 , n14398 );
    xnor g14917 ( n14737 , n3132 , n21957 );
    or g14918 ( n17924 , n15697 , n7104 );
    and g14919 ( n7806 , n18316 , n15480 );
    and g14920 ( n19036 , n13440 , n23944 );
    not g14921 ( n14791 , n21944 );
    xnor g14922 ( n6491 , n1765 , n12875 );
    buf g14923 ( n23064 , n8898 );
    xnor g14924 ( n14091 , n18441 , n1117 );
    and g14925 ( n20343 , n24761 , n13746 );
    nor g14926 ( n9432 , n2850 , n19907 );
    or g14927 ( n9542 , n25263 , n18387 );
    nor g14928 ( n22867 , n6051 , n25276 );
    xnor g14929 ( n7570 , n18145 , n26191 );
    and g14930 ( n23246 , n9131 , n15704 );
    not g14931 ( n18655 , n5419 );
    and g14932 ( n2001 , n16930 , n662 );
    not g14933 ( n966 , n18720 );
    not g14934 ( n27183 , n16449 );
    xnor g14935 ( n3001 , n7402 , n7305 );
    xnor g14936 ( n20004 , n22219 , n11553 );
    or g14937 ( n1849 , n1116 , n7646 );
    not g14938 ( n20886 , n14792 );
    or g14939 ( n24233 , n5348 , n19226 );
    or g14940 ( n24594 , n3393 , n1465 );
    or g14941 ( n15541 , n18090 , n1252 );
    xnor g14942 ( n22538 , n17212 , n20411 );
    not g14943 ( n4040 , n6397 );
    xnor g14944 ( n13587 , n9431 , n27076 );
    xnor g14945 ( n2937 , n2213 , n26269 );
    or g14946 ( n18156 , n15125 , n11929 );
    or g14947 ( n2620 , n24562 , n14018 );
    xnor g14948 ( n19577 , n5213 , n19081 );
    and g14949 ( n20799 , n9470 , n15320 );
    not g14950 ( n14628 , n20970 );
    not g14951 ( n23428 , n18035 );
    nor g14952 ( n571 , n17568 , n2978 );
    or g14953 ( n5661 , n7841 , n19595 );
    or g14954 ( n18505 , n16473 , n2111 );
    not g14955 ( n24116 , n24620 );
    and g14956 ( n25766 , n17267 , n23517 );
    and g14957 ( n22665 , n11237 , n10091 );
    or g14958 ( n15771 , n18118 , n1928 );
    and g14959 ( n352 , n7123 , n6615 );
    xnor g14960 ( n7346 , n17001 , n1784 );
    not g14961 ( n2027 , n9498 );
    xnor g14962 ( n3718 , n6319 , n19836 );
    nor g14963 ( n1472 , n56 , n20506 );
    not g14964 ( n19277 , n19081 );
    and g14965 ( n23176 , n11208 , n20899 );
    and g14966 ( n15759 , n11465 , n21109 );
    or g14967 ( n7469 , n10593 , n1662 );
    xnor g14968 ( n9419 , n8357 , n17082 );
    or g14969 ( n19151 , n14961 , n5520 );
    nor g14970 ( n22038 , n2013 , n22640 );
    or g14971 ( n14851 , n14760 , n6734 );
    or g14972 ( n13706 , n20108 , n12411 );
    or g14973 ( n20823 , n21781 , n25549 );
    and g14974 ( n12598 , n7550 , n7858 );
    xnor g14975 ( n22262 , n18409 , n8259 );
    xnor g14976 ( n7240 , n23430 , n19081 );
    xnor g14977 ( n23885 , n4888 , n1572 );
    or g14978 ( n25135 , n19805 , n5125 );
    or g14979 ( n11999 , n840 , n19719 );
    not g14980 ( n14389 , n26177 );
    xnor g14981 ( n8087 , n1206 , n4260 );
    xnor g14982 ( n16479 , n4217 , n22683 );
    xnor g14983 ( n24920 , n18338 , n12644 );
    not g14984 ( n12421 , n25449 );
    not g14985 ( n5616 , n12999 );
    or g14986 ( n9374 , n3604 , n11815 );
    nor g14987 ( n14203 , n14465 , n6356 );
    or g14988 ( n4680 , n4312 , n21903 );
    not g14989 ( n26324 , n3823 );
    nor g14990 ( n6177 , n15633 , n8097 );
    not g14991 ( n22688 , n12075 );
    nor g14992 ( n14073 , n1939 , n13818 );
    or g14993 ( n22946 , n6938 , n1201 );
    xnor g14994 ( n10321 , n10764 , n2253 );
    not g14995 ( n25260 , n11230 );
    xnor g14996 ( n8845 , n14804 , n20579 );
    or g14997 ( n27125 , n4614 , n15132 );
    nor g14998 ( n26945 , n19172 , n7371 );
    not g14999 ( n5697 , n8511 );
    nor g15000 ( n20022 , n11550 , n13884 );
    and g15001 ( n22180 , n14098 , n18124 );
    xnor g15002 ( n24486 , n17897 , n20278 );
    and g15003 ( n5242 , n13902 , n3557 );
    xnor g15004 ( n21258 , n5752 , n14071 );
    xnor g15005 ( n16807 , n26026 , n4905 );
    nor g15006 ( n11087 , n19005 , n12889 );
    not g15007 ( n9680 , n2102 );
    xnor g15008 ( n25062 , n16950 , n11632 );
    or g15009 ( n8703 , n8448 , n15892 );
    nor g15010 ( n20759 , n4938 , n25345 );
    xnor g15011 ( n18667 , n9748 , n3037 );
    not g15012 ( n7682 , n18409 );
    or g15013 ( n8697 , n16326 , n7199 );
    and g15014 ( n12180 , n3605 , n2748 );
    and g15015 ( n10361 , n6108 , n20911 );
    not g15016 ( n5891 , n9011 );
    or g15017 ( n16102 , n24219 , n8792 );
    and g15018 ( n22638 , n916 , n21211 );
    xnor g15019 ( n14606 , n14397 , n10125 );
    xnor g15020 ( n23277 , n9278 , n5561 );
    buf g15021 ( n16880 , n9140 );
    and g15022 ( n1729 , n23115 , n1849 );
    xnor g15023 ( n6637 , n22084 , n4765 );
    nor g15024 ( n12525 , n3124 , n24170 );
    or g15025 ( n14585 , n3938 , n9853 );
    or g15026 ( n1507 , n18212 , n15223 );
    xnor g15027 ( n6837 , n7693 , n3909 );
    nor g15028 ( n8 , n26688 , n14256 );
    and g15029 ( n12051 , n6218 , n7669 );
    and g15030 ( n25959 , n992 , n19311 );
    or g15031 ( n14745 , n19761 , n26684 );
    and g15032 ( n12092 , n9970 , n24413 );
    or g15033 ( n4188 , n19090 , n13085 );
    xnor g15034 ( n8154 , n14130 , n468 );
    not g15035 ( n21804 , n21654 );
    or g15036 ( n5294 , n3231 , n3533 );
    xnor g15037 ( n11420 , n8906 , n2420 );
    xnor g15038 ( n5332 , n24592 , n21291 );
    xnor g15039 ( n15784 , n25582 , n17035 );
    xnor g15040 ( n17711 , n11 , n20331 );
    xnor g15041 ( n25362 , n14915 , n9510 );
    and g15042 ( n19774 , n13316 , n6266 );
    or g15043 ( n21595 , n11672 , n6401 );
    or g15044 ( n7355 , n468 , n22322 );
    xnor g15045 ( n1946 , n16282 , n20714 );
    and g15046 ( n14018 , n23391 , n6763 );
    xnor g15047 ( n13056 , n11229 , n9741 );
    xnor g15048 ( n12765 , n13906 , n13026 );
    or g15049 ( n9193 , n24552 , n24618 );
    or g15050 ( n1744 , n26568 , n13767 );
    or g15051 ( n15673 , n1946 , n1629 );
    not g15052 ( n12208 , n13384 );
    or g15053 ( n15030 , n688 , n7674 );
    xnor g15054 ( n17963 , n21747 , n25397 );
    xnor g15055 ( n21098 , n11394 , n17847 );
    xnor g15056 ( n26545 , n18314 , n20635 );
    not g15057 ( n13066 , n23876 );
    and g15058 ( n18165 , n14434 , n14869 );
    nor g15059 ( n8410 , n12663 , n14974 );
    xnor g15060 ( n26582 , n19564 , n7918 );
    xnor g15061 ( n20239 , n26265 , n6485 );
    or g15062 ( n4452 , n23245 , n3778 );
    not g15063 ( n1923 , n6955 );
    not g15064 ( n27009 , n6362 );
    xnor g15065 ( n22824 , n10998 , n22793 );
    and g15066 ( n5070 , n15578 , n17991 );
    or g15067 ( n26394 , n26660 , n3232 );
    xnor g15068 ( n14865 , n16319 , n23882 );
    not g15069 ( n27114 , n18123 );
    xnor g15070 ( n24028 , n15681 , n13333 );
    and g15071 ( n19272 , n7402 , n23099 );
    or g15072 ( n3855 , n4499 , n16136 );
    xnor g15073 ( n20172 , n21710 , n6508 );
    nor g15074 ( n10475 , n25962 , n17468 );
    nor g15075 ( n14619 , n6209 , n12241 );
    or g15076 ( n8171 , n134 , n17702 );
    xnor g15077 ( n49 , n5740 , n25770 );
    or g15078 ( n14978 , n11452 , n3460 );
    not g15079 ( n1637 , n8272 );
    not g15080 ( n4317 , n4104 );
    xnor g15081 ( n18005 , n4479 , n23724 );
    xnor g15082 ( n14550 , n24184 , n25923 );
    or g15083 ( n24738 , n1587 , n13303 );
    xnor g15084 ( n25018 , n19527 , n21993 );
    xnor g15085 ( n4553 , n21406 , n11165 );
    xnor g15086 ( n9605 , n19687 , n6219 );
    xnor g15087 ( n21680 , n16997 , n60 );
    not g15088 ( n1631 , n10219 );
    xnor g15089 ( n26745 , n15907 , n24404 );
    or g15090 ( n23363 , n25868 , n13200 );
    not g15091 ( n9877 , n19284 );
    xnor g15092 ( n5158 , n18019 , n186 );
    and g15093 ( n25577 , n3774 , n1613 );
    not g15094 ( n22906 , n17636 );
    or g15095 ( n24022 , n13897 , n22121 );
    xnor g15096 ( n10596 , n20131 , n10048 );
    or g15097 ( n9825 , n6400 , n11069 );
    and g15098 ( n4388 , n16614 , n4238 );
    xnor g15099 ( n23422 , n12567 , n11048 );
    xnor g15100 ( n20107 , n17108 , n4008 );
    xnor g15101 ( n9431 , n26286 , n16492 );
    or g15102 ( n3557 , n12053 , n7527 );
    xnor g15103 ( n17712 , n2565 , n23261 );
    and g15104 ( n2338 , n12389 , n23143 );
    xnor g15105 ( n148 , n5299 , n15546 );
    and g15106 ( n13178 , n4623 , n373 );
    xnor g15107 ( n17176 , n21235 , n5025 );
    and g15108 ( n18390 , n2712 , n26221 );
    nor g15109 ( n10876 , n10587 , n9163 );
    xnor g15110 ( n23354 , n17672 , n2832 );
    not g15111 ( n9392 , n9901 );
    nor g15112 ( n8254 , n12971 , n13553 );
    or g15113 ( n8346 , n19611 , n22582 );
    nor g15114 ( n10414 , n17035 , n13206 );
    not g15115 ( n20438 , n21585 );
    and g15116 ( n21074 , n18276 , n17086 );
    not g15117 ( n6522 , n9022 );
    or g15118 ( n17029 , n228 , n9239 );
    not g15119 ( n7348 , n274 );
    and g15120 ( n17548 , n17966 , n5762 );
    nor g15121 ( n1848 , n11044 , n4325 );
    xnor g15122 ( n17811 , n5673 , n16146 );
    nor g15123 ( n14624 , n26748 , n20196 );
    not g15124 ( n14356 , n24907 );
    xnor g15125 ( n3 , n16348 , n25321 );
    or g15126 ( n3489 , n4547 , n7540 );
    xnor g15127 ( n4501 , n5194 , n12161 );
    and g15128 ( n20360 , n8223 , n10678 );
    or g15129 ( n4495 , n26519 , n6194 );
    xnor g15130 ( n19570 , n12782 , n17811 );
    xnor g15131 ( n996 , n10571 , n9431 );
    xnor g15132 ( n21710 , n1143 , n11709 );
    not g15133 ( n24111 , n20234 );
    or g15134 ( n23577 , n9432 , n24803 );
    or g15135 ( n4450 , n8018 , n16700 );
    and g15136 ( n5830 , n19011 , n22117 );
    and g15137 ( n1653 , n23858 , n24702 );
    and g15138 ( n18860 , n478 , n19421 );
    not g15139 ( n14087 , n11047 );
    not g15140 ( n575 , n6733 );
    or g15141 ( n23398 , n12751 , n12696 );
    nor g15142 ( n21100 , n15427 , n14337 );
    xnor g15143 ( n26208 , n11747 , n15161 );
    not g15144 ( n8197 , n20887 );
    nor g15145 ( n4969 , n4883 , n27076 );
    or g15146 ( n17056 , n22366 , n5550 );
    xnor g15147 ( n21094 , n8438 , n3741 );
    or g15148 ( n26852 , n17725 , n1562 );
    xnor g15149 ( n21160 , n5211 , n21832 );
    nor g15150 ( n23057 , n7470 , n1730 );
    xnor g15151 ( n19854 , n12248 , n1696 );
    or g15152 ( n22401 , n12891 , n9266 );
    and g15153 ( n24694 , n9719 , n21639 );
    nor g15154 ( n6843 , n12002 , n11056 );
    and g15155 ( n2531 , n25311 , n380 );
    or g15156 ( n15579 , n26450 , n6819 );
    or g15157 ( n2621 , n992 , n19311 );
    xnor g15158 ( n26405 , n5714 , n26409 );
    xnor g15159 ( n19583 , n26979 , n18962 );
    xnor g15160 ( n11644 , n13261 , n22591 );
    or g15161 ( n2019 , n19525 , n25862 );
    nor g15162 ( n20674 , n26744 , n8456 );
    not g15163 ( n18749 , n9971 );
    or g15164 ( n3336 , n12698 , n18443 );
    xnor g15165 ( n16769 , n25494 , n1314 );
    nor g15166 ( n10003 , n2268 , n4326 );
    xnor g15167 ( n25685 , n23080 , n2133 );
    xnor g15168 ( n20610 , n10405 , n23974 );
    xnor g15169 ( n8688 , n14869 , n24795 );
    or g15170 ( n26468 , n16601 , n18580 );
    nor g15171 ( n359 , n23024 , n10522 );
    xnor g15172 ( n24184 , n15472 , n22821 );
    not g15173 ( n12299 , n11019 );
    and g15174 ( n177 , n19437 , n18640 );
    and g15175 ( n27087 , n3511 , n11602 );
    or g15176 ( n5881 , n25015 , n4890 );
    nor g15177 ( n19546 , n14431 , n25877 );
    and g15178 ( n278 , n8654 , n1094 );
    or g15179 ( n6229 , n24370 , n18868 );
    or g15180 ( n25473 , n10166 , n26652 );
    or g15181 ( n17785 , n15301 , n24789 );
    not g15182 ( n6610 , n10083 );
    xnor g15183 ( n1370 , n12501 , n8067 );
    nor g15184 ( n12224 , n23396 , n17790 );
    or g15185 ( n19449 , n2694 , n7823 );
    and g15186 ( n6497 , n26259 , n10016 );
    or g15187 ( n16775 , n8155 , n15077 );
    xnor g15188 ( n23034 , n11762 , n20190 );
    not g15189 ( n22247 , n25439 );
    xnor g15190 ( n19737 , n26979 , n5704 );
    or g15191 ( n26099 , n21036 , n4118 );
    and g15192 ( n1958 , n25068 , n17881 );
    xnor g15193 ( n12848 , n342 , n14570 );
    or g15194 ( n12919 , n7731 , n19858 );
    xnor g15195 ( n8432 , n17429 , n22255 );
    xnor g15196 ( n12119 , n17542 , n19840 );
    and g15197 ( n19715 , n23397 , n5398 );
    and g15198 ( n24962 , n11151 , n4295 );
    xnor g15199 ( n5170 , n12317 , n1186 );
    xnor g15200 ( n15857 , n602 , n4858 );
    or g15201 ( n2008 , n18335 , n16911 );
    xnor g15202 ( n16025 , n3925 , n12121 );
    xnor g15203 ( n14609 , n1552 , n27006 );
    or g15204 ( n9336 , n27063 , n10203 );
    xnor g15205 ( n14635 , n21480 , n14225 );
    or g15206 ( n24777 , n3329 , n23358 );
    xnor g15207 ( n917 , n15038 , n2217 );
    xnor g15208 ( n20495 , n4916 , n18346 );
    and g15209 ( n19544 , n5147 , n20350 );
    xnor g15210 ( n18790 , n24218 , n4501 );
    xnor g15211 ( n18945 , n16660 , n25687 );
    nor g15212 ( n14940 , n3161 , n11630 );
    or g15213 ( n3512 , n1350 , n6637 );
    and g15214 ( n14422 , n16477 , n10767 );
    nor g15215 ( n3975 , n6895 , n20462 );
    or g15216 ( n1072 , n21888 , n18044 );
    nor g15217 ( n4254 , n21846 , n19608 );
    and g15218 ( n7425 , n10391 , n10383 );
    and g15219 ( n13917 , n19510 , n5175 );
    not g15220 ( n4125 , n2114 );
    xnor g15221 ( n820 , n13772 , n14668 );
    or g15222 ( n11527 , n6800 , n22152 );
    or g15223 ( n1932 , n14936 , n25324 );
    or g15224 ( n9083 , n275 , n12133 );
    or g15225 ( n10975 , n10909 , n2541 );
    or g15226 ( n208 , n18269 , n10784 );
    and g15227 ( n27043 , n14818 , n16631 );
    xnor g15228 ( n982 , n2627 , n26489 );
    xnor g15229 ( n5404 , n9897 , n19132 );
    and g15230 ( n24095 , n23137 , n13320 );
    or g15231 ( n10682 , n5512 , n5067 );
    not g15232 ( n21973 , n4118 );
    nor g15233 ( n13856 , n139 , n914 );
    xnor g15234 ( n4509 , n25835 , n7519 );
    or g15235 ( n24316 , n6760 , n21649 );
    or g15236 ( n15578 , n18814 , n17090 );
    xnor g15237 ( n12147 , n18365 , n12850 );
    xnor g15238 ( n20443 , n24961 , n5243 );
    or g15239 ( n14889 , n9813 , n953 );
    or g15240 ( n10006 , n23343 , n21064 );
    xnor g15241 ( n980 , n14655 , n22970 );
    nor g15242 ( n1291 , n3465 , n2244 );
    or g15243 ( n11625 , n12136 , n15531 );
    or g15244 ( n20322 , n7311 , n15780 );
    or g15245 ( n15115 , n2519 , n8951 );
    xnor g15246 ( n852 , n2778 , n21504 );
    not g15247 ( n9050 , n26107 );
    xnor g15248 ( n19488 , n7213 , n9172 );
    or g15249 ( n21787 , n10881 , n17324 );
    or g15250 ( n16866 , n5400 , n9512 );
    or g15251 ( n19530 , n12996 , n13376 );
    or g15252 ( n22969 , n20909 , n7397 );
    or g15253 ( n6040 , n13080 , n12362 );
    not g15254 ( n16227 , n8244 );
    and g15255 ( n3109 , n11199 , n15757 );
    not g15256 ( n8736 , n12406 );
    nor g15257 ( n14874 , n23791 , n20925 );
    or g15258 ( n24079 , n17899 , n9169 );
    buf g15259 ( n2252 , n17299 );
    or g15260 ( n375 , n14580 , n14195 );
    or g15261 ( n13640 , n20056 , n17692 );
    not g15262 ( n6828 , n14838 );
    not g15263 ( n7952 , n10158 );
    and g15264 ( n20200 , n12002 , n11918 );
    not g15265 ( n9457 , n7805 );
    xnor g15266 ( n18168 , n17690 , n713 );
    not g15267 ( n14573 , n15383 );
    xnor g15268 ( n11181 , n8792 , n26334 );
    and g15269 ( n11575 , n2940 , n2464 );
    or g15270 ( n12010 , n1389 , n2677 );
    xnor g15271 ( n23558 , n21667 , n26387 );
    and g15272 ( n22465 , n4903 , n20858 );
    and g15273 ( n21778 , n15444 , n4072 );
    xnor g15274 ( n13503 , n20314 , n10046 );
    or g15275 ( n576 , n25936 , n16712 );
    or g15276 ( n26799 , n23804 , n10997 );
    xnor g15277 ( n2298 , n19597 , n21785 );
    buf g15278 ( n3356 , n1512 );
    and g15279 ( n17974 , n150 , n17022 );
    not g15280 ( n10452 , n16524 );
    or g15281 ( n3325 , n11244 , n7587 );
    or g15282 ( n8603 , n26580 , n3716 );
    or g15283 ( n26346 , n2975 , n20938 );
    or g15284 ( n5278 , n22319 , n17134 );
    xnor g15285 ( n18429 , n21026 , n23803 );
    xnor g15286 ( n18477 , n15898 , n11271 );
    and g15287 ( n7749 , n21279 , n4389 );
    or g15288 ( n9464 , n25954 , n25241 );
    or g15289 ( n9953 , n2928 , n18494 );
    not g15290 ( n5238 , n4410 );
    xnor g15291 ( n26438 , n15678 , n13475 );
    or g15292 ( n5289 , n17939 , n24214 );
    xnor g15293 ( n25213 , n26724 , n5226 );
    or g15294 ( n4737 , n9887 , n10630 );
    and g15295 ( n228 , n23083 , n17858 );
    xnor g15296 ( n22377 , n2978 , n3425 );
    and g15297 ( n12549 , n9078 , n10759 );
    and g15298 ( n13678 , n7895 , n26349 );
    xnor g15299 ( n13484 , n24743 , n5191 );
    or g15300 ( n2567 , n19949 , n15210 );
    nor g15301 ( n19130 , n493 , n14969 );
    and g15302 ( n16511 , n13109 , n24898 );
    or g15303 ( n21695 , n23121 , n23395 );
    xnor g15304 ( n20616 , n27183 , n2150 );
    or g15305 ( n22367 , n699 , n23661 );
    or g15306 ( n10546 , n15110 , n16701 );
    not g15307 ( n10470 , n15258 );
    nor g15308 ( n9849 , n880 , n19328 );
    not g15309 ( n26363 , n10795 );
    nor g15310 ( n7018 , n13376 , n16731 );
    or g15311 ( n17049 , n8781 , n21058 );
    or g15312 ( n7995 , n10403 , n23956 );
    xnor g15313 ( n22780 , n21506 , n19911 );
    and g15314 ( n10994 , n22739 , n13970 );
    and g15315 ( n22356 , n8793 , n15804 );
    xnor g15316 ( n8553 , n6316 , n18647 );
    nor g15317 ( n6677 , n26660 , n18907 );
    or g15318 ( n21851 , n12202 , n12672 );
    xnor g15319 ( n20670 , n23693 , n10505 );
    not g15320 ( n8738 , n19089 );
    nor g15321 ( n23675 , n5449 , n9647 );
    not g15322 ( n1984 , n354 );
    and g15323 ( n1550 , n27060 , n25543 );
    or g15324 ( n20817 , n10841 , n2386 );
    xnor g15325 ( n12256 , n4194 , n8795 );
    xnor g15326 ( n13489 , n6625 , n9598 );
    or g15327 ( n26761 , n25866 , n14836 );
    xnor g15328 ( n16062 , n13259 , n12252 );
    or g15329 ( n17175 , n20470 , n14052 );
    xnor g15330 ( n24427 , n13303 , n3785 );
    xnor g15331 ( n12424 , n27188 , n6502 );
    or g15332 ( n15100 , n26925 , n9394 );
    not g15333 ( n8624 , n10984 );
    or g15334 ( n17655 , n7802 , n10785 );
    xnor g15335 ( n17703 , n17769 , n7638 );
    and g15336 ( n18195 , n21312 , n13673 );
    nor g15337 ( n5539 , n19465 , n2126 );
    or g15338 ( n16821 , n6759 , n10755 );
    not g15339 ( n13766 , n7272 );
    or g15340 ( n2304 , n361 , n13867 );
    not g15341 ( n10457 , n23375 );
    or g15342 ( n25820 , n24638 , n19327 );
    or g15343 ( n3574 , n7849 , n6123 );
    or g15344 ( n22844 , n22442 , n22253 );
    xnor g15345 ( n23987 , n18585 , n25713 );
    or g15346 ( n21311 , n16542 , n24655 );
    nor g15347 ( n6786 , n20415 , n255 );
    not g15348 ( n8456 , n23587 );
    or g15349 ( n10286 , n3514 , n20867 );
    and g15350 ( n5321 , n11737 , n14274 );
    or g15351 ( n22236 , n20289 , n6184 );
    or g15352 ( n11163 , n25584 , n18435 );
    nor g15353 ( n10496 , n19110 , n26753 );
    or g15354 ( n3738 , n24018 , n13074 );
    or g15355 ( n14371 , n1673 , n14579 );
    xnor g15356 ( n15808 , n3339 , n15252 );
    and g15357 ( n9087 , n25379 , n11625 );
    and g15358 ( n2485 , n644 , n154 );
    or g15359 ( n26163 , n16947 , n25899 );
    or g15360 ( n7386 , n15992 , n6093 );
    xnor g15361 ( n12654 , n21492 , n10605 );
    or g15362 ( n6966 , n14600 , n563 );
    not g15363 ( n19017 , n13625 );
    xnor g15364 ( n13613 , n13569 , n17553 );
    or g15365 ( n21499 , n2055 , n619 );
    or g15366 ( n289 , n26459 , n21195 );
    and g15367 ( n13442 , n25820 , n22032 );
    nor g15368 ( n25201 , n22219 , n12514 );
    and g15369 ( n3497 , n15987 , n9139 );
    and g15370 ( n19078 , n13797 , n13496 );
    and g15371 ( n19426 , n14825 , n10931 );
    xnor g15372 ( n11010 , n370 , n2228 );
    not g15373 ( n17847 , n259 );
    or g15374 ( n22985 , n15072 , n8748 );
    nor g15375 ( n3424 , n3356 , n19758 );
    xnor g15376 ( n10228 , n2346 , n14768 );
    xnor g15377 ( n19322 , n11366 , n11669 );
    nor g15378 ( n25309 , n16339 , n5569 );
    and g15379 ( n20106 , n19042 , n18846 );
    and g15380 ( n12450 , n20903 , n624 );
    xnor g15381 ( n19125 , n2452 , n16484 );
    not g15382 ( n20811 , n24200 );
    or g15383 ( n523 , n18383 , n5255 );
    nor g15384 ( n14964 , n26252 , n7750 );
    xnor g15385 ( n22897 , n2977 , n325 );
    xnor g15386 ( n22255 , n26499 , n22083 );
    or g15387 ( n18407 , n22298 , n19751 );
    xnor g15388 ( n7538 , n10811 , n8965 );
    xnor g15389 ( n19045 , n21542 , n1378 );
    xnor g15390 ( n8286 , n3587 , n22278 );
    and g15391 ( n9184 , n18131 , n13724 );
    or g15392 ( n23255 , n16906 , n16138 );
    not g15393 ( n17143 , n2389 );
    xnor g15394 ( n20671 , n24197 , n10094 );
    xnor g15395 ( n23435 , n589 , n23293 );
    not g15396 ( n21652 , n14261 );
    and g15397 ( n16918 , n1282 , n9167 );
    and g15398 ( n3476 , n8359 , n27040 );
    or g15399 ( n2193 , n21865 , n12628 );
    not g15400 ( n11162 , n17756 );
    or g15401 ( n22997 , n6779 , n14463 );
    xnor g15402 ( n25850 , n18926 , n6513 );
    or g15403 ( n425 , n3174 , n3006 );
    and g15404 ( n16721 , n14293 , n26886 );
    and g15405 ( n12222 , n3405 , n24165 );
    and g15406 ( n26981 , n25542 , n26214 );
    or g15407 ( n15106 , n5619 , n22541 );
    or g15408 ( n21812 , n17579 , n4859 );
    and g15409 ( n12849 , n4436 , n21406 );
    xnor g15410 ( n12272 , n14504 , n8964 );
    xnor g15411 ( n9317 , n9394 , n26925 );
    not g15412 ( n11249 , n23717 );
    not g15413 ( n5436 , n580 );
    or g15414 ( n4784 , n5349 , n3990 );
    and g15415 ( n23988 , n25832 , n2188 );
    or g15416 ( n24597 , n16975 , n24470 );
    nor g15417 ( n1581 , n19023 , n18375 );
    or g15418 ( n14367 , n7678 , n11579 );
    xnor g15419 ( n2189 , n2882 , n17190 );
    or g15420 ( n3104 , n12115 , n23256 );
    nor g15421 ( n8185 , n19974 , n22440 );
    and g15422 ( n15096 , n10554 , n330 );
    nor g15423 ( n24114 , n12258 , n19116 );
    or g15424 ( n25597 , n207 , n25030 );
    not g15425 ( n11559 , n7731 );
    or g15426 ( n6348 , n23789 , n25555 );
    and g15427 ( n7003 , n10096 , n24511 );
    xnor g15428 ( n4163 , n17572 , n6692 );
    xnor g15429 ( n10595 , n18382 , n18142 );
    xnor g15430 ( n25994 , n9891 , n15872 );
    not g15431 ( n23581 , n5674 );
    not g15432 ( n18514 , n17351 );
    or g15433 ( n17020 , n24768 , n1019 );
    xnor g15434 ( n1102 , n10710 , n26510 );
    xnor g15435 ( n11758 , n15557 , n18807 );
    xnor g15436 ( n9609 , n15113 , n26832 );
    xnor g15437 ( n9858 , n17004 , n15193 );
    not g15438 ( n7930 , n6596 );
    or g15439 ( n8843 , n19361 , n15918 );
    xnor g15440 ( n22891 , n19421 , n8217 );
    xnor g15441 ( n26804 , n11158 , n11566 );
    nor g15442 ( n21342 , n6948 , n1911 );
    xnor g15443 ( n20021 , n12956 , n26913 );
    xnor g15444 ( n22624 , n5855 , n7693 );
    xnor g15445 ( n25893 , n6814 , n10763 );
    or g15446 ( n20507 , n20563 , n21191 );
    or g15447 ( n158 , n14431 , n22587 );
    nor g15448 ( n20681 , n2768 , n5924 );
    xnor g15449 ( n20436 , n3969 , n18998 );
    not g15450 ( n26904 , n2570 );
    and g15451 ( n9886 , n2395 , n11259 );
    or g15452 ( n15387 , n10941 , n12901 );
    and g15453 ( n13956 , n15933 , n6153 );
    xnor g15454 ( n25971 , n4187 , n4225 );
    or g15455 ( n8628 , n2939 , n2316 );
    or g15456 ( n7136 , n15736 , n19352 );
    and g15457 ( n823 , n24170 , n23460 );
    and g15458 ( n19995 , n6066 , n7701 );
    xnor g15459 ( n13835 , n21990 , n17427 );
    nor g15460 ( n15604 , n2750 , n25393 );
    and g15461 ( n9583 , n12553 , n14872 );
    and g15462 ( n14112 , n18170 , n3444 );
    or g15463 ( n20270 , n26528 , n25017 );
    not g15464 ( n18247 , n25057 );
    not g15465 ( n18474 , n14845 );
    or g15466 ( n15425 , n21520 , n24106 );
    nor g15467 ( n16045 , n26241 , n2999 );
    xnor g15468 ( n8117 , n233 , n22583 );
    xnor g15469 ( n13445 , n17674 , n17911 );
    or g15470 ( n13404 , n22585 , n26837 );
    not g15471 ( n6904 , n21134 );
    or g15472 ( n3005 , n22439 , n26235 );
    or g15473 ( n21391 , n19155 , n25458 );
    or g15474 ( n14436 , n1637 , n23822 );
    or g15475 ( n8312 , n6408 , n14815 );
    xnor g15476 ( n10304 , n17069 , n16608 );
    or g15477 ( n13673 , n24127 , n9207 );
    xnor g15478 ( n3836 , n7312 , n4180 );
    xnor g15479 ( n618 , n13240 , n21473 );
    and g15480 ( n24306 , n10882 , n8719 );
    not g15481 ( n180 , n25265 );
    and g15482 ( n17564 , n25932 , n14771 );
    xnor g15483 ( n14816 , n16303 , n4481 );
    xnor g15484 ( n7337 , n17728 , n17959 );
    nor g15485 ( n7151 , n23708 , n6013 );
    xnor g15486 ( n16277 , n11243 , n2421 );
    xnor g15487 ( n25200 , n5875 , n13473 );
    xnor g15488 ( n2642 , n5728 , n24704 );
    nor g15489 ( n15877 , n15439 , n7248 );
    xnor g15490 ( n26117 , n8220 , n7361 );
    or g15491 ( n4235 , n11695 , n2135 );
    xnor g15492 ( n17796 , n19247 , n25957 );
    and g15493 ( n14373 , n7357 , n24332 );
    xnor g15494 ( n2852 , n13234 , n18737 );
    not g15495 ( n23312 , n11747 );
    xnor g15496 ( n18466 , n1601 , n24151 );
    and g15497 ( n13583 , n8655 , n11037 );
    not g15498 ( n7827 , n19263 );
    xnor g15499 ( n24121 , n20018 , n10033 );
    or g15500 ( n5594 , n2657 , n10482 );
    or g15501 ( n4455 , n13361 , n8300 );
    nor g15502 ( n4380 , n19138 , n24984 );
    xnor g15503 ( n1809 , n18027 , n25101 );
    not g15504 ( n14021 , n17040 );
    xnor g15505 ( n8126 , n22824 , n8385 );
    xor g15506 ( n3152 , n21469 , n9713 );
    xnor g15507 ( n2361 , n25774 , n4885 );
    or g15508 ( n14072 , n9094 , n22655 );
    xnor g15509 ( n14459 , n14514 , n24536 );
    not g15510 ( n14818 , n1136 );
    not g15511 ( n11944 , n17261 );
    xnor g15512 ( n9778 , n22689 , n2650 );
    not g15513 ( n24125 , n24932 );
    xnor g15514 ( n11662 , n14588 , n10288 );
    xor g15515 ( n1862 , n13343 , n11784 );
    or g15516 ( n12409 , n24850 , n15271 );
    xnor g15517 ( n12545 , n4210 , n10790 );
    xnor g15518 ( n21238 , n16629 , n1214 );
    not g15519 ( n7543 , n6956 );
    or g15520 ( n7202 , n898 , n10503 );
    or g15521 ( n10247 , n3366 , n4753 );
    not g15522 ( n11158 , n10973 );
    not g15523 ( n6303 , n26371 );
    or g15524 ( n876 , n26980 , n8387 );
    and g15525 ( n1974 , n12247 , n15971 );
    and g15526 ( n18597 , n17797 , n10789 );
    not g15527 ( n20314 , n25089 );
    buf g15528 ( n22820 , n26119 );
    or g15529 ( n6742 , n17251 , n26107 );
    nor g15530 ( n24158 , n4371 , n11849 );
    xnor g15531 ( n504 , n22900 , n13142 );
    xnor g15532 ( n9968 , n1916 , n23749 );
    xnor g15533 ( n5074 , n7023 , n12126 );
    xnor g15534 ( n11458 , n23932 , n20385 );
    and g15535 ( n26245 , n13634 , n16997 );
    xnor g15536 ( n11623 , n22608 , n2101 );
    and g15537 ( n17463 , n23963 , n20807 );
    not g15538 ( n7020 , n17703 );
    xnor g15539 ( n7468 , n4713 , n7805 );
    nor g15540 ( n9284 , n4721 , n5140 );
    xnor g15541 ( n4224 , n1849 , n12034 );
    xnor g15542 ( n21123 , n18932 , n14243 );
    xnor g15543 ( n8398 , n18132 , n14527 );
    not g15544 ( n9595 , n25515 );
    xnor g15545 ( n11698 , n4659 , n8182 );
    xnor g15546 ( n19315 , n14784 , n20058 );
    and g15547 ( n15800 , n25710 , n18162 );
    nor g15548 ( n26649 , n11186 , n7099 );
    xnor g15549 ( n12670 , n9446 , n17372 );
    or g15550 ( n4428 , n16383 , n21742 );
    xnor g15551 ( n9394 , n23292 , n17533 );
    and g15552 ( n21572 , n15751 , n20434 );
    xnor g15553 ( n26103 , n26510 , n1112 );
    not g15554 ( n14516 , n8379 );
    and g15555 ( n8300 , n25459 , n23282 );
    not g15556 ( n8675 , n4967 );
    and g15557 ( n19867 , n5785 , n16353 );
    xnor g15558 ( n17487 , n26872 , n19531 );
    not g15559 ( n18928 , n7752 );
    xnor g15560 ( n964 , n2162 , n7941 );
    nor g15561 ( n20159 , n12509 , n7761 );
    or g15562 ( n9147 , n25540 , n14845 );
    or g15563 ( n1347 , n13390 , n8053 );
    and g15564 ( n17917 , n13542 , n14688 );
    and g15565 ( n19131 , n16557 , n12934 );
    or g15566 ( n23022 , n23921 , n5946 );
    xnor g15567 ( n14458 , n211 , n195 );
    or g15568 ( n23826 , n16061 , n7614 );
    or g15569 ( n23336 , n6192 , n20885 );
    xnor g15570 ( n14584 , n26684 , n9088 );
    xnor g15571 ( n26815 , n21966 , n24269 );
    nor g15572 ( n24836 , n2829 , n23620 );
    or g15573 ( n750 , n23746 , n13161 );
    xnor g15574 ( n17212 , n20074 , n20409 );
    nor g15575 ( n25829 , n14172 , n611 );
    nor g15576 ( n26599 , n1584 , n17690 );
    or g15577 ( n26539 , n24484 , n23995 );
    xnor g15578 ( n11724 , n4535 , n17662 );
    nor g15579 ( n21245 , n25345 , n21322 );
    or g15580 ( n21966 , n24477 , n13091 );
    not g15581 ( n19806 , n11738 );
    nor g15582 ( n15983 , n12145 , n9814 );
    and g15583 ( n13786 , n1541 , n25495 );
    or g15584 ( n13395 , n9309 , n3119 );
    xnor g15585 ( n11209 , n10999 , n23463 );
    or g15586 ( n22726 , n11316 , n10663 );
    xnor g15587 ( n16386 , n1056 , n16689 );
    nor g15588 ( n6029 , n4426 , n13109 );
    xnor g15589 ( n7390 , n25702 , n6462 );
    or g15590 ( n6973 , n23640 , n1083 );
    xnor g15591 ( n9821 , n18801 , n10130 );
    or g15592 ( n21983 , n832 , n15424 );
    or g15593 ( n21539 , n18963 , n19956 );
    not g15594 ( n1405 , n6138 );
    and g15595 ( n20857 , n14870 , n8888 );
    or g15596 ( n4164 , n23666 , n26134 );
    nor g15597 ( n13000 , n13480 , n11544 );
    and g15598 ( n3634 , n3909 , n24200 );
    or g15599 ( n23532 , n524 , n18027 );
    and g15600 ( n6589 , n1805 , n14674 );
    xnor g15601 ( n26337 , n24839 , n22009 );
    xnor g15602 ( n18467 , n1579 , n22822 );
    or g15603 ( n4066 , n1705 , n5354 );
    not g15604 ( n7860 , n6710 );
    or g15605 ( n13734 , n20787 , n13769 );
    xnor g15606 ( n13476 , n4203 , n20207 );
    or g15607 ( n19387 , n15695 , n13502 );
    and g15608 ( n5468 , n11594 , n1342 );
    nor g15609 ( n8483 , n16012 , n20127 );
    xnor g15610 ( n5627 , n20043 , n16611 );
    not g15611 ( n17497 , n7086 );
    xnor g15612 ( n9429 , n10712 , n23586 );
    xnor g15613 ( n25442 , n27161 , n21448 );
    xnor g15614 ( n6046 , n2410 , n23370 );
    nor g15615 ( n9064 , n23144 , n1662 );
    and g15616 ( n15301 , n13263 , n8979 );
    or g15617 ( n20130 , n15149 , n21955 );
    xnor g15618 ( n10800 , n27089 , n8806 );
    xnor g15619 ( n12223 , n25541 , n1575 );
    or g15620 ( n16790 , n24939 , n18416 );
    xnor g15621 ( n9089 , n5709 , n26834 );
    xnor g15622 ( n23285 , n24339 , n17176 );
    or g15623 ( n681 , n3097 , n3764 );
    or g15624 ( n6227 , n11516 , n4513 );
    and g15625 ( n12583 , n4858 , n8224 );
    xnor g15626 ( n12225 , n12243 , n2642 );
    not g15627 ( n19797 , n22327 );
    xnor g15628 ( n19501 , n20235 , n8259 );
    and g15629 ( n24380 , n5391 , n7784 );
    not g15630 ( n8132 , n20054 );
    or g15631 ( n25034 , n15050 , n26700 );
    and g15632 ( n13464 , n7814 , n1393 );
    not g15633 ( n4360 , n16812 );
    not g15634 ( n11066 , n17408 );
    xnor g15635 ( n2352 , n8351 , n25519 );
    not g15636 ( n25691 , n26394 );
    and g15637 ( n13756 , n7517 , n24318 );
    and g15638 ( n20962 , n15899 , n18520 );
    nor g15639 ( n25058 , n11044 , n7619 );
    or g15640 ( n4694 , n13525 , n3691 );
    or g15641 ( n26315 , n17954 , n23608 );
    or g15642 ( n3645 , n5226 , n21205 );
    not g15643 ( n9180 , n5211 );
    nor g15644 ( n14621 , n13037 , n8295 );
    nor g15645 ( n24555 , n2230 , n8869 );
    xnor g15646 ( n5673 , n17194 , n17417 );
    or g15647 ( n13218 , n10291 , n5192 );
    nor g15648 ( n11788 , n4410 , n9456 );
    xnor g15649 ( n16301 , n13775 , n6397 );
    and g15650 ( n16704 , n9801 , n21574 );
    xnor g15651 ( n21046 , n10532 , n4782 );
    xnor g15652 ( n2946 , n24281 , n8492 );
    and g15653 ( n2604 , n8866 , n26570 );
    xnor g15654 ( n8355 , n10501 , n5914 );
    xnor g15655 ( n17108 , n18033 , n10478 );
    xnor g15656 ( n5694 , n3186 , n23224 );
    and g15657 ( n20191 , n13708 , n21083 );
    xnor g15658 ( n18377 , n21917 , n8585 );
    not g15659 ( n22652 , n19360 );
    xnor g15660 ( n7544 , n10017 , n5026 );
    not g15661 ( n24143 , n8313 );
    nor g15662 ( n8092 , n3441 , n8959 );
    xnor g15663 ( n18632 , n25084 , n8366 );
    and g15664 ( n15288 , n11227 , n16370 );
    and g15665 ( n2378 , n4022 , n14565 );
    xnor g15666 ( n5860 , n10383 , n25336 );
    not g15667 ( n2187 , n9054 );
    nor g15668 ( n15326 , n10405 , n23974 );
    and g15669 ( n10269 , n6688 , n1746 );
    or g15670 ( n2550 , n20560 , n14462 );
    xnor g15671 ( n2533 , n25986 , n16959 );
    xnor g15672 ( n26776 , n182 , n17171 );
    xnor g15673 ( n26288 , n8869 , n1738 );
    not g15674 ( n16065 , n8166 );
    or g15675 ( n23683 , n2858 , n18727 );
    and g15676 ( n4239 , n5935 , n13952 );
    xnor g15677 ( n16825 , n14671 , n9707 );
    xnor g15678 ( n15827 , n18805 , n8614 );
    and g15679 ( n20527 , n5167 , n6458 );
    and g15680 ( n13939 , n26200 , n13233 );
    nor g15681 ( n23163 , n24015 , n4749 );
    xnor g15682 ( n1308 , n5089 , n17947 );
    nor g15683 ( n7768 , n9180 , n18537 );
    or g15684 ( n6109 , n14603 , n1141 );
    or g15685 ( n19382 , n22476 , n25748 );
    xnor g15686 ( n6099 , n2412 , n15884 );
    or g15687 ( n23360 , n9598 , n350 );
    and g15688 ( n12468 , n19839 , n6518 );
    and g15689 ( n4848 , n16189 , n7451 );
    or g15690 ( n2508 , n12875 , n7751 );
    or g15691 ( n13213 , n19518 , n15677 );
    or g15692 ( n9947 , n17635 , n20080 );
    not g15693 ( n13329 , n26001 );
    or g15694 ( n17402 , n26658 , n18991 );
    not g15695 ( n10301 , n15688 );
    and g15696 ( n13544 , n11996 , n7430 );
    and g15697 ( n26021 , n20270 , n23379 );
    nor g15698 ( n8796 , n23369 , n22906 );
    not g15699 ( n23800 , n7734 );
    nor g15700 ( n25798 , n24348 , n8332 );
    not g15701 ( n13863 , n2421 );
    or g15702 ( n7643 , n22085 , n15368 );
    not g15703 ( n5095 , n15775 );
    nor g15704 ( n7344 , n528 , n1639 );
    xnor g15705 ( n4719 , n5667 , n26953 );
    and g15706 ( n8975 , n21867 , n22248 );
    and g15707 ( n2397 , n20577 , n6519 );
    and g15708 ( n16056 , n3809 , n8406 );
    not g15709 ( n21097 , n23829 );
    xnor g15710 ( n26590 , n358 , n19274 );
    nor g15711 ( n4440 , n312 , n799 );
    not g15712 ( n8602 , n6808 );
    nor g15713 ( n2348 , n18649 , n3795 );
    and g15714 ( n4207 , n9941 , n9868 );
    not g15715 ( n20245 , n15289 );
    xnor g15716 ( n26520 , n1367 , n8296 );
    or g15717 ( n11353 , n16293 , n5600 );
    xnor g15718 ( n7990 , n17599 , n9093 );
    or g15719 ( n12085 , n6203 , n13333 );
    nor g15720 ( n5867 , n25524 , n16117 );
    xnor g15721 ( n8665 , n21565 , n5103 );
    xnor g15722 ( n17171 , n24253 , n398 );
    and g15723 ( n21640 , n18349 , n25703 );
    xnor g15724 ( n22107 , n25482 , n2901 );
    or g15725 ( n6657 , n19332 , n4001 );
    and g15726 ( n7557 , n3026 , n8752 );
    nor g15727 ( n15640 , n11273 , n9026 );
    xnor g15728 ( n14282 , n10269 , n14135 );
    not g15729 ( n4982 , n13573 );
    or g15730 ( n10171 , n20842 , n5054 );
    and g15731 ( n9298 , n19469 , n25625 );
    xnor g15732 ( n24602 , n10091 , n22376 );
    or g15733 ( n365 , n24387 , n13507 );
    or g15734 ( n25343 , n2296 , n13582 );
    or g15735 ( n2097 , n17838 , n8954 );
    and g15736 ( n23252 , n11616 , n981 );
    or g15737 ( n19336 , n26658 , n1118 );
    not g15738 ( n11871 , n3414 );
    or g15739 ( n16869 , n23068 , n13171 );
    or g15740 ( n12793 , n16244 , n19741 );
    or g15741 ( n16446 , n11243 , n26497 );
    nor g15742 ( n6010 , n1009 , n1742 );
    or g15743 ( n22455 , n22173 , n583 );
    or g15744 ( n25212 , n14974 , n12652 );
    or g15745 ( n7851 , n3162 , n24878 );
    or g15746 ( n7250 , n11008 , n12743 );
    nor g15747 ( n19166 , n11479 , n679 );
    or g15748 ( n11810 , n11566 , n13150 );
    or g15749 ( n13792 , n16347 , n13261 );
    not g15750 ( n15236 , n25359 );
    xnor g15751 ( n26429 , n8514 , n17189 );
    or g15752 ( n9434 , n6485 , n26265 );
    nor g15753 ( n4076 , n8539 , n7627 );
    or g15754 ( n13132 , n10623 , n7613 );
    or g15755 ( n19256 , n7917 , n3380 );
    xnor g15756 ( n22575 , n19228 , n5226 );
    nor g15757 ( n6533 , n23763 , n13492 );
    and g15758 ( n15329 , n14846 , n16297 );
    or g15759 ( n24073 , n3635 , n22635 );
    or g15760 ( n7645 , n9044 , n21183 );
    and g15761 ( n20908 , n10037 , n13148 );
    and g15762 ( n26384 , n27035 , n11163 );
    nor g15763 ( n12472 , n22318 , n3391 );
    or g15764 ( n1440 , n24252 , n10081 );
    and g15765 ( n23658 , n24187 , n19331 );
    or g15766 ( n16772 , n19 , n16476 );
    xnor g15767 ( n25611 , n4832 , n2534 );
    or g15768 ( n15757 , n5781 , n14112 );
    nor g15769 ( n7777 , n6115 , n7385 );
    or g15770 ( n16802 , n3856 , n20834 );
    or g15771 ( n3159 , n12819 , n23186 );
    not g15772 ( n22722 , n20002 );
    not g15773 ( n6877 , n866 );
    and g15774 ( n233 , n20282 , n20294 );
    not g15775 ( n6285 , n14447 );
    and g15776 ( n1576 , n8568 , n23793 );
    xnor g15777 ( n2122 , n1627 , n14773 );
    and g15778 ( n5741 , n18979 , n23138 );
    xnor g15779 ( n10177 , n1099 , n6381 );
    nor g15780 ( n16962 , n14362 , n14240 );
    and g15781 ( n7904 , n20686 , n20507 );
    and g15782 ( n26270 , n26457 , n7063 );
    not g15783 ( n3993 , n13072 );
    xnor g15784 ( n26077 , n5328 , n15780 );
    xnor g15785 ( n14761 , n22234 , n2175 );
    or g15786 ( n5658 , n10668 , n13212 );
    nor g15787 ( n9828 , n14704 , n17716 );
    not g15788 ( n20497 , n5400 );
    xnor g15789 ( n24488 , n9553 , n25919 );
    and g15790 ( n6014 , n9357 , n23155 );
    or g15791 ( n22854 , n9718 , n5425 );
    xnor g15792 ( n1143 , n18314 , n12644 );
    or g15793 ( n26321 , n7553 , n10879 );
    and g15794 ( n22656 , n11030 , n6141 );
    nor g15795 ( n24211 , n22290 , n13018 );
    and g15796 ( n16000 , n5994 , n18348 );
    xnor g15797 ( n21580 , n17231 , n16354 );
    xnor g15798 ( n1481 , n4934 , n20658 );
    xnor g15799 ( n25937 , n24920 , n21639 );
    xnor g15800 ( n10617 , n24589 , n3588 );
    and g15801 ( n16066 , n8790 , n7633 );
    not g15802 ( n6670 , n8225 );
    not g15803 ( n23365 , n16713 );
    or g15804 ( n2494 , n17017 , n19418 );
    or g15805 ( n1076 , n23804 , n21138 );
    or g15806 ( n3250 , n3689 , n20135 );
    and g15807 ( n15651 , n6485 , n18676 );
    xnor g15808 ( n15909 , n25941 , n17495 );
    xnor g15809 ( n11194 , n13494 , n4319 );
    or g15810 ( n26854 , n16812 , n14397 );
    xnor g15811 ( n20317 , n18295 , n25974 );
    or g15812 ( n16272 , n4729 , n10096 );
    xnor g15813 ( n16356 , n13529 , n5474 );
    and g15814 ( n10186 , n23303 , n15067 );
    xnor g15815 ( n10236 , n22118 , n1170 );
    xnor g15816 ( n4489 , n17316 , n18734 );
    not g15817 ( n22615 , n22303 );
    and g15818 ( n16553 , n10213 , n14924 );
    and g15819 ( n14182 , n6904 , n17419 );
    nor g15820 ( n14840 , n19616 , n1118 );
    and g15821 ( n5711 , n26552 , n3337 );
    or g15822 ( n18364 , n23230 , n4665 );
    xnor g15823 ( n8280 , n2595 , n26484 );
    not g15824 ( n2675 , n8988 );
    and g15825 ( n26881 , n26659 , n16187 );
    not g15826 ( n4130 , n7871 );
    and g15827 ( n4020 , n10025 , n24456 );
    not g15828 ( n14536 , n5443 );
    and g15829 ( n18198 , n9181 , n8926 );
    not g15830 ( n5925 , n20961 );
    and g15831 ( n21555 , n1260 , n22555 );
    xnor g15832 ( n13499 , n20138 , n25073 );
    or g15833 ( n15242 , n22792 , n1550 );
    and g15834 ( n17036 , n21535 , n19787 );
    xnor g15835 ( n23424 , n111 , n5587 );
    or g15836 ( n9491 , n16106 , n26964 );
    xnor g15837 ( n20014 , n4303 , n4387 );
    xnor g15838 ( n23951 , n1019 , n24768 );
    and g15839 ( n1625 , n12260 , n25990 );
    or g15840 ( n8123 , n11201 , n26340 );
    and g15841 ( n25189 , n8060 , n9482 );
    nor g15842 ( n5631 , n18191 , n18188 );
    nor g15843 ( n10606 , n16496 , n17350 );
    not g15844 ( n2522 , n985 );
    or g15845 ( n5391 , n18601 , n19874 );
    not g15846 ( n26724 , n9992 );
    nor g15847 ( n27012 , n4100 , n24609 );
    xnor g15848 ( n17172 , n5329 , n10053 );
    and g15849 ( n9148 , n26868 , n22205 );
    or g15850 ( n16035 , n2746 , n4609 );
    not g15851 ( n4798 , n22091 );
    and g15852 ( n23087 , n16673 , n1408 );
    or g15853 ( n3198 , n11736 , n18183 );
    or g15854 ( n2357 , n19849 , n26585 );
    not g15855 ( n9538 , n10468 );
    xnor g15856 ( n21233 , n24403 , n23175 );
    xnor g15857 ( n14475 , n5282 , n17837 );
    and g15858 ( n6419 , n2866 , n19645 );
    not g15859 ( n10608 , n15359 );
    nor g15860 ( n16041 , n9570 , n6785 );
    not g15861 ( n14829 , n15214 );
    nor g15862 ( n18375 , n6631 , n7339 );
    xnor g15863 ( n8858 , n5135 , n7792 );
    xnor g15864 ( n23199 , n8371 , n6464 );
    or g15865 ( n18681 , n4868 , n23820 );
    not g15866 ( n11802 , n16910 );
    not g15867 ( n14795 , n2041 );
    or g15868 ( n26115 , n1029 , n19281 );
    not g15869 ( n15026 , n4293 );
    or g15870 ( n14334 , n2502 , n366 );
    and g15871 ( n20432 , n18525 , n876 );
    xnor g15872 ( n18225 , n22755 , n310 );
    or g15873 ( n3215 , n6027 , n7239 );
    or g15874 ( n21383 , n14515 , n10735 );
    or g15875 ( n10871 , n13163 , n6497 );
    xnor g15876 ( n18339 , n7671 , n4959 );
    xnor g15877 ( n17322 , n3837 , n7325 );
    and g15878 ( n21016 , n8248 , n22917 );
    or g15879 ( n19246 , n2207 , n22142 );
    xnor g15880 ( n10212 , n23460 , n24170 );
    xnor g15881 ( n16369 , n1742 , n19196 );
    or g15882 ( n26130 , n5657 , n733 );
    or g15883 ( n10819 , n2721 , n14826 );
    or g15884 ( n1399 , n16607 , n1244 );
    not g15885 ( n11542 , n2409 );
    or g15886 ( n19289 , n22545 , n7875 );
    or g15887 ( n16525 , n5426 , n8028 );
    or g15888 ( n21243 , n5750 , n2249 );
    xnor g15889 ( n11515 , n19480 , n14787 );
    not g15890 ( n5227 , n20432 );
    xnor g15891 ( n2598 , n13339 , n12562 );
    and g15892 ( n23738 , n19653 , n18132 );
    and g15893 ( n14313 , n11781 , n24396 );
    nor g15894 ( n26887 , n10788 , n16900 );
    nor g15895 ( n26146 , n3946 , n18318 );
    or g15896 ( n7694 , n14722 , n13442 );
    not g15897 ( n6864 , n15969 );
    xnor g15898 ( n11993 , n22591 , n26167 );
    xnor g15899 ( n1480 , n23064 , n3582 );
    or g15900 ( n5375 , n874 , n12267 );
    not g15901 ( n5574 , n2510 );
    not g15902 ( n258 , n8799 );
    or g15903 ( n10642 , n24823 , n13893 );
    not g15904 ( n7041 , n9133 );
    xnor g15905 ( n921 , n15509 , n14304 );
    nor g15906 ( n6054 , n4195 , n21671 );
    or g15907 ( n25437 , n23162 , n5868 );
    xnor g15908 ( n6297 , n7096 , n7876 );
    not g15909 ( n22535 , n6360 );
    xnor g15910 ( n14423 , n21071 , n7906 );
    xnor g15911 ( n23747 , n10117 , n3306 );
    or g15912 ( n21429 , n15796 , n10739 );
    and g15913 ( n16872 , n25237 , n21710 );
    not g15914 ( n12465 , n16126 );
    or g15915 ( n11547 , n2949 , n43 );
    or g15916 ( n12227 , n15240 , n27185 );
    not g15917 ( n26830 , n20687 );
    or g15918 ( n3373 , n22176 , n21662 );
    not g15919 ( n12991 , n7466 );
    xnor g15920 ( n1915 , n4261 , n117 );
    not g15921 ( n27075 , n303 );
    xnor g15922 ( n12502 , n26541 , n4967 );
    or g15923 ( n14674 , n6815 , n19505 );
    xnor g15924 ( n12246 , n27204 , n18545 );
    not g15925 ( n1036 , n18438 );
    or g15926 ( n3060 , n4654 , n25874 );
    and g15927 ( n13502 , n9052 , n11082 );
    or g15928 ( n15915 , n20513 , n12605 );
    or g15929 ( n21581 , n3460 , n16667 );
    xnor g15930 ( n20500 , n3164 , n2547 );
    xnor g15931 ( n22267 , n17380 , n20927 );
    or g15932 ( n70 , n18190 , n3084 );
    or g15933 ( n19484 , n25738 , n11265 );
    xnor g15934 ( n25009 , n11503 , n12593 );
    or g15935 ( n2600 , n14441 , n20240 );
    or g15936 ( n11293 , n9942 , n13946 );
    xnor g15937 ( n19409 , n20284 , n3779 );
    and g15938 ( n5823 , n20378 , n4677 );
    not g15939 ( n25558 , n20923 );
    and g15940 ( n11077 , n13376 , n4643 );
    xnor g15941 ( n12605 , n21474 , n11354 );
    or g15942 ( n13430 , n18506 , n4812 );
    xnor g15943 ( n8729 , n6240 , n19497 );
    xnor g15944 ( n23982 , n1036 , n20728 );
    or g15945 ( n2572 , n23043 , n26622 );
    or g15946 ( n24494 , n22308 , n14407 );
    or g15947 ( n16307 , n26460 , n19649 );
    or g15948 ( n3064 , n19902 , n12535 );
    not g15949 ( n16660 , n18063 );
    or g15950 ( n11396 , n18352 , n2129 );
    xnor g15951 ( n18039 , n3018 , n2731 );
    nor g15952 ( n11680 , n22077 , n21838 );
    and g15953 ( n18852 , n3120 , n14361 );
    not g15954 ( n26497 , n1434 );
    xnor g15955 ( n22474 , n2291 , n24791 );
    or g15956 ( n19829 , n25643 , n20604 );
    xnor g15957 ( n23980 , n1755 , n24993 );
    and g15958 ( n2523 , n741 , n7594 );
    and g15959 ( n10531 , n20425 , n15498 );
    xnor g15960 ( n17805 , n2281 , n1047 );
    nor g15961 ( n6398 , n840 , n11186 );
    xnor g15962 ( n9535 , n10223 , n17078 );
    xnor g15963 ( n10010 , n18588 , n3845 );
    xnor g15964 ( n13652 , n15696 , n13709 );
    or g15965 ( n2069 , n9678 , n1484 );
    xnor g15966 ( n14787 , n23612 , n14488 );
    or g15967 ( n23561 , n20554 , n19058 );
    xnor g15968 ( n6307 , n21993 , n14575 );
    xnor g15969 ( n18975 , n16838 , n20267 );
    xnor g15970 ( n22986 , n16561 , n23596 );
    or g15971 ( n18066 , n20747 , n18540 );
    or g15972 ( n21079 , n2403 , n25125 );
    buf g15973 ( n11554 , n8626 );
    not g15974 ( n4659 , n3955 );
    xnor g15975 ( n18094 , n19005 , n7149 );
    or g15976 ( n20257 , n11550 , n1626 );
    xnor g15977 ( n14320 , n2980 , n4781 );
    or g15978 ( n19105 , n20880 , n376 );
    not g15979 ( n23231 , n3668 );
    xnor g15980 ( n7729 , n27015 , n22993 );
    xnor g15981 ( n8798 , n5527 , n25218 );
    nor g15982 ( n1307 , n6865 , n3727 );
    xnor g15983 ( n22473 , n8418 , n6356 );
    or g15984 ( n21491 , n25480 , n16904 );
    nor g15985 ( n12134 , n19340 , n234 );
    not g15986 ( n19082 , n6775 );
    xnor g15987 ( n25356 , n25011 , n2943 );
    xnor g15988 ( n22122 , n4580 , n5057 );
    xnor g15989 ( n1172 , n26892 , n26047 );
    xnor g15990 ( n17051 , n2160 , n7335 );
    xnor g15991 ( n9217 , n12694 , n22450 );
    nor g15992 ( n26891 , n11840 , n23059 );
    or g15993 ( n17675 , n23800 , n1308 );
    xnor g15994 ( n13551 , n7552 , n26609 );
    xnor g15995 ( n22808 , n14041 , n10359 );
    or g15996 ( n14424 , n20826 , n17326 );
    or g15997 ( n10175 , n12454 , n16755 );
    nor g15998 ( n15260 , n21540 , n13485 );
    or g15999 ( n9470 , n21083 , n13708 );
    xnor g16000 ( n10756 , n5995 , n22627 );
    not g16001 ( n3333 , n21727 );
    or g16002 ( n8311 , n16937 , n14002 );
    or g16003 ( n10931 , n14517 , n2839 );
    xnor g16004 ( n24002 , n8839 , n25852 );
    nor g16005 ( n1202 , n8305 , n2918 );
    or g16006 ( n15710 , n9196 , n6775 );
    nor g16007 ( n8757 , n2017 , n650 );
    xnor g16008 ( n14032 , n8645 , n15635 );
    or g16009 ( n4565 , n9401 , n22121 );
    not g16010 ( n945 , n19569 );
    not g16011 ( n23281 , n2696 );
    xnor g16012 ( n20190 , n2816 , n1222 );
    not g16013 ( n12511 , n1742 );
    nor g16014 ( n15880 , n8422 , n25627 );
    nor g16015 ( n6061 , n18261 , n12398 );
    and g16016 ( n555 , n12244 , n14673 );
    and g16017 ( n5301 , n8421 , n4305 );
    or g16018 ( n24069 , n989 , n22847 );
    or g16019 ( n15013 , n22804 , n21309 );
    or g16020 ( n18923 , n17446 , n11606 );
    or g16021 ( n2584 , n16298 , n3819 );
    or g16022 ( n4402 , n4704 , n14365 );
    and g16023 ( n10630 , n4976 , n15694 );
    xnor g16024 ( n19664 , n2741 , n5581 );
    xnor g16025 ( n18020 , n21850 , n25751 );
    not g16026 ( n17120 , n22332 );
    and g16027 ( n26369 , n19574 , n13185 );
    xnor g16028 ( n6298 , n21070 , n17317 );
    and g16029 ( n10896 , n8978 , n27123 );
    nor g16030 ( n2512 , n20794 , n25471 );
    xnor g16031 ( n12278 , n4181 , n13879 );
    or g16032 ( n2311 , n2668 , n12807 );
    not g16033 ( n22440 , n23435 );
    nor g16034 ( n24582 , n14692 , n14437 );
    or g16035 ( n20860 , n19594 , n12749 );
    xnor g16036 ( n11653 , n25746 , n8973 );
    or g16037 ( n22786 , n20 , n16907 );
    nor g16038 ( n17456 , n18741 , n22782 );
    xnor g16039 ( n18899 , n5972 , n1823 );
    not g16040 ( n2875 , n27126 );
    and g16041 ( n526 , n16916 , n3624 );
    or g16042 ( n15976 , n24806 , n5342 );
    or g16043 ( n21105 , n7973 , n15179 );
    or g16044 ( n24060 , n4132 , n13074 );
    and g16045 ( n8173 , n4875 , n4209 );
    nor g16046 ( n26374 , n16309 , n23873 );
    not g16047 ( n6887 , n24984 );
    and g16048 ( n26127 , n20945 , n22953 );
    xnor g16049 ( n14538 , n13207 , n24427 );
    xnor g16050 ( n17837 , n5669 , n21575 );
    not g16051 ( n18191 , n1570 );
    not g16052 ( n20404 , n25322 );
    or g16053 ( n13236 , n24631 , n352 );
    nor g16054 ( n23771 , n16249 , n14557 );
    not g16055 ( n8155 , n22379 );
    nor g16056 ( n26445 , n19144 , n5496 );
    or g16057 ( n6087 , n303 , n25101 );
    xnor g16058 ( n17922 , n4749 , n24015 );
    xnor g16059 ( n5964 , n13236 , n3355 );
    or g16060 ( n15689 , n25649 , n19581 );
    and g16061 ( n22681 , n7222 , n19601 );
    and g16062 ( n22699 , n22723 , n5692 );
    or g16063 ( n15896 , n2334 , n12598 );
    or g16064 ( n22811 , n20404 , n14661 );
    or g16065 ( n21612 , n23753 , n3240 );
    or g16066 ( n624 , n18465 , n3580 );
    nor g16067 ( n15292 , n21599 , n9576 );
    nor g16068 ( n16454 , n4844 , n8052 );
    and g16069 ( n21821 , n26539 , n8476 );
    and g16070 ( n17897 , n19815 , n2581 );
    and g16071 ( n19155 , n8910 , n25018 );
    or g16072 ( n23933 , n1291 , n4829 );
    and g16073 ( n18044 , n12409 , n17934 );
    or g16074 ( n3269 , n21871 , n6659 );
    and g16075 ( n14132 , n1654 , n7893 );
    xnor g16076 ( n10914 , n12774 , n12121 );
    not g16077 ( n2994 , n5568 );
    and g16078 ( n12805 , n23082 , n9613 );
    not g16079 ( n20883 , n12137 );
    and g16080 ( n25825 , n17919 , n26773 );
    xnor g16081 ( n18425 , n13813 , n17496 );
    xnor g16082 ( n6553 , n962 , n9318 );
    and g16083 ( n12292 , n10426 , n12635 );
    or g16084 ( n14618 , n5407 , n20604 );
    not g16085 ( n12217 , n1674 );
    and g16086 ( n1337 , n18406 , n9959 );
    xnor g16087 ( n22020 , n20854 , n20352 );
    and g16088 ( n18548 , n16252 , n17943 );
    xnor g16089 ( n15914 , n15798 , n20832 );
    or g16090 ( n13256 , n18847 , n12110 );
    xnor g16091 ( n5182 , n11006 , n16212 );
    or g16092 ( n21051 , n144 , n11919 );
    not g16093 ( n6351 , n19858 );
    and g16094 ( n12798 , n12268 , n5573 );
    xnor g16095 ( n13784 , n5988 , n13677 );
    and g16096 ( n21041 , n6405 , n3765 );
    and g16097 ( n23296 , n9671 , n5205 );
    or g16098 ( n3950 , n26079 , n7863 );
    xnor g16099 ( n24913 , n21194 , n27008 );
    xnor g16100 ( n27179 , n7692 , n25464 );
    not g16101 ( n6226 , n19678 );
    or g16102 ( n24761 , n10514 , n10041 );
    xnor g16103 ( n18414 , n19536 , n1764 );
    nor g16104 ( n23069 , n3239 , n1464 );
    xnor g16105 ( n78 , n18035 , n5834 );
    and g16106 ( n25785 , n4411 , n14197 );
    nor g16107 ( n18518 , n570 , n2479 );
    xnor g16108 ( n12078 , n21612 , n23825 );
    or g16109 ( n2577 , n21749 , n2298 );
    not g16110 ( n18223 , n13218 );
    not g16111 ( n18615 , n19262 );
    xnor g16112 ( n21368 , n9076 , n704 );
    or g16113 ( n13138 , n14684 , n1667 );
    xnor g16114 ( n18519 , n7920 , n20976 );
    and g16115 ( n14171 , n16713 , n17497 );
    and g16116 ( n13890 , n10514 , n10041 );
    xnor g16117 ( n5482 , n10135 , n2809 );
    xnor g16118 ( n362 , n20655 , n19951 );
    and g16119 ( n25092 , n14520 , n21712 );
    or g16120 ( n25098 , n27033 , n4207 );
    not g16121 ( n13899 , n26208 );
    nor g16122 ( n5154 , n15282 , n9859 );
    xnor g16123 ( n25385 , n5475 , n7324 );
    xnor g16124 ( n6171 , n14371 , n17997 );
    not g16125 ( n1720 , n2747 );
    not g16126 ( n20376 , n2719 );
    and g16127 ( n7158 , n20994 , n12669 );
    xnor g16128 ( n20421 , n23993 , n19731 );
    xnor g16129 ( n2976 , n19286 , n10245 );
    xnor g16130 ( n14607 , n1522 , n1599 );
    xnor g16131 ( n22159 , n14974 , n12663 );
    or g16132 ( n6338 , n21456 , n22537 );
    and g16133 ( n17575 , n14224 , n11097 );
    or g16134 ( n15524 , n173 , n16167 );
    not g16135 ( n4846 , n5862 );
    and g16136 ( n27124 , n14367 , n11142 );
    not g16137 ( n15164 , n13558 );
    or g16138 ( n18276 , n14337 , n24865 );
    or g16139 ( n4707 , n13899 , n8233 );
    xnor g16140 ( n16713 , n21039 , n14694 );
    xnor g16141 ( n18229 , n24732 , n12892 );
    xnor g16142 ( n9461 , n1519 , n5263 );
    xnor g16143 ( n8662 , n13524 , n9225 );
    xnor g16144 ( n19649 , n12676 , n18791 );
    nor g16145 ( n23237 , n9671 , n10712 );
    or g16146 ( n14629 , n16747 , n15520 );
    xnor g16147 ( n17312 , n26564 , n22744 );
    or g16148 ( n16508 , n14040 , n8477 );
    and g16149 ( n1535 , n1989 , n18369 );
    and g16150 ( n7539 , n17330 , n24140 );
    and g16151 ( n24556 , n18447 , n24350 );
    and g16152 ( n26932 , n341 , n21569 );
    xnor g16153 ( n13477 , n22737 , n17220 );
    and g16154 ( n11083 , n10819 , n1813 );
    and g16155 ( n6579 , n19448 , n21966 );
    not g16156 ( n10049 , n25068 );
    not g16157 ( n4174 , n7082 );
    or g16158 ( n15476 , n18134 , n16539 );
    or g16159 ( n5088 , n23877 , n20354 );
    xnor g16160 ( n18586 , n23800 , n5163 );
    or g16161 ( n7701 , n6391 , n24800 );
    and g16162 ( n11798 , n6456 , n17978 );
    not g16163 ( n19614 , n18820 );
    not g16164 ( n20951 , n13940 );
    or g16165 ( n10060 , n26767 , n21470 );
    or g16166 ( n4179 , n8509 , n17087 );
    xnor g16167 ( n12346 , n20003 , n15343 );
    or g16168 ( n26555 , n19770 , n11451 );
    xnor g16169 ( n8585 , n7071 , n14848 );
    or g16170 ( n6312 , n11011 , n1019 );
    xnor g16171 ( n23139 , n7143 , n10728 );
    nor g16172 ( n13983 , n22083 , n26215 );
    or g16173 ( n18367 , n22868 , n1153 );
    not g16174 ( n11137 , n20485 );
    nor g16175 ( n1537 , n18295 , n16223 );
    not g16176 ( n11889 , n2337 );
    or g16177 ( n760 , n5682 , n3862 );
    and g16178 ( n11804 , n10792 , n17230 );
    nor g16179 ( n19066 , n17203 , n17597 );
    or g16180 ( n1303 , n3334 , n9998 );
    or g16181 ( n19969 , n22518 , n14824 );
    xnor g16182 ( n23238 , n10459 , n12313 );
    or g16183 ( n26619 , n16144 , n18107 );
    or g16184 ( n17521 , n9829 , n22181 );
    or g16185 ( n14006 , n25855 , n26461 );
    or g16186 ( n11634 , n17037 , n21385 );
    nor g16187 ( n20596 , n7656 , n669 );
    xnor g16188 ( n14885 , n1529 , n14786 );
    or g16189 ( n16891 , n14001 , n20543 );
    nor g16190 ( n11595 , n15586 , n17495 );
    or g16191 ( n22331 , n14699 , n21300 );
    nor g16192 ( n747 , n16687 , n5319 );
    xnor g16193 ( n26046 , n8607 , n25523 );
    not g16194 ( n21841 , n23864 );
    xnor g16195 ( n11023 , n3787 , n22818 );
    xnor g16196 ( n24415 , n8021 , n10591 );
    or g16197 ( n7288 , n17091 , n9711 );
    not g16198 ( n21207 , n6691 );
    xnor g16199 ( n6908 , n5035 , n18531 );
    xnor g16200 ( n25328 , n20395 , n21746 );
    xnor g16201 ( n336 , n13424 , n23831 );
    or g16202 ( n2215 , n15806 , n20300 );
    or g16203 ( n19816 , n12301 , n560 );
    not g16204 ( n3727 , n6703 );
    xnor g16205 ( n3513 , n1028 , n1618 );
    and g16206 ( n3808 , n7192 , n11956 );
    and g16207 ( n2956 , n14540 , n16023 );
    not g16208 ( n10106 , n7883 );
    and g16209 ( n19285 , n16796 , n10256 );
    or g16210 ( n4336 , n9740 , n17850 );
    or g16211 ( n15363 , n13967 , n20964 );
    xnor g16212 ( n13747 , n23508 , n22945 );
    xnor g16213 ( n12266 , n19926 , n1243 );
    and g16214 ( n8981 , n13783 , n6341 );
    nor g16215 ( n12130 , n2914 , n16376 );
    xnor g16216 ( n19064 , n1128 , n19948 );
    and g16217 ( n14022 , n25817 , n23052 );
    and g16218 ( n15178 , n22634 , n17816 );
    xnor g16219 ( n14805 , n650 , n9872 );
    xnor g16220 ( n22815 , n4461 , n17954 );
    xnor g16221 ( n3568 , n26234 , n18697 );
    not g16222 ( n15560 , n20826 );
    nor g16223 ( n19818 , n15415 , n25523 );
    not g16224 ( n25639 , n4602 );
    xnor g16225 ( n4064 , n20751 , n16466 );
    and g16226 ( n24698 , n15279 , n23817 );
    xnor g16227 ( n24812 , n14218 , n7737 );
    nor g16228 ( n10982 , n26197 , n4555 );
    or g16229 ( n7192 , n8689 , n21508 );
    or g16230 ( n14876 , n8562 , n8941 );
    xnor g16231 ( n3844 , n150 , n24315 );
    nor g16232 ( n13408 , n25604 , n26499 );
    nor g16233 ( n22468 , n2017 , n11649 );
    xnor g16234 ( n354 , n4502 , n24901 );
    or g16235 ( n103 , n10593 , n5817 );
    or g16236 ( n7718 , n2883 , n4018 );
    and g16237 ( n25422 , n25640 , n5702 );
    or g16238 ( n21803 , n25049 , n20731 );
    xnor g16239 ( n8533 , n26373 , n25418 );
    xnor g16240 ( n15803 , n2566 , n4894 );
    xnor g16241 ( n12570 , n11006 , n10113 );
    and g16242 ( n18622 , n15825 , n14370 );
    xnor g16243 ( n9822 , n8088 , n8624 );
    or g16244 ( n14526 , n7074 , n19000 );
    nor g16245 ( n13909 , n27037 , n23913 );
    or g16246 ( n2011 , n2023 , n15675 );
    nor g16247 ( n11896 , n20102 , n14269 );
    xnor g16248 ( n12204 , n14209 , n6162 );
    xnor g16249 ( n10009 , n12231 , n724 );
    not g16250 ( n23141 , n26054 );
    or g16251 ( n8815 , n12613 , n22680 );
    not g16252 ( n2996 , n25980 );
    not g16253 ( n14958 , n8272 );
    xnor g16254 ( n557 , n24863 , n5252 );
    nor g16255 ( n1771 , n19227 , n24298 );
    xnor g16256 ( n26530 , n1761 , n2817 );
    or g16257 ( n15632 , n8629 , n21352 );
    or g16258 ( n7449 , n20315 , n11869 );
    and g16259 ( n18359 , n6844 , n15040 );
    xnor g16260 ( n24345 , n11809 , n16957 );
    not g16261 ( n26302 , n4786 );
    and g16262 ( n9337 , n1333 , n19051 );
    or g16263 ( n5104 , n1587 , n14008 );
    xnor g16264 ( n20872 , n8570 , n6996 );
    xnor g16265 ( n2042 , n10092 , n23644 );
    not g16266 ( n21771 , n25031 );
    and g16267 ( n13829 , n7367 , n15993 );
    or g16268 ( n26342 , n12258 , n152 );
    and g16269 ( n2541 , n18041 , n21012 );
    or g16270 ( n22708 , n1896 , n25886 );
    nor g16271 ( n724 , n1833 , n9834 );
    or g16272 ( n18015 , n23771 , n907 );
    or g16273 ( n25955 , n2239 , n23415 );
    or g16274 ( n2442 , n17351 , n26528 );
    xnor g16275 ( n21636 , n21172 , n6369 );
    or g16276 ( n4392 , n13384 , n16106 );
    or g16277 ( n1330 , n25693 , n7131 );
    or g16278 ( n16150 , n22243 , n2143 );
    xnor g16279 ( n5231 , n9724 , n17689 );
    or g16280 ( n413 , n24382 , n24262 );
    and g16281 ( n18752 , n3645 , n3747 );
    nor g16282 ( n24437 , n22962 , n12209 );
    xnor g16283 ( n14561 , n27037 , n11736 );
    xnor g16284 ( n18807 , n1293 , n19196 );
    and g16285 ( n589 , n17577 , n20341 );
    xnor g16286 ( n24542 , n18608 , n19899 );
    nor g16287 ( n20292 , n21288 , n25238 );
    not g16288 ( n11165 , n10034 );
    or g16289 ( n12732 , n17970 , n3700 );
    xnor g16290 ( n15009 , n17453 , n26783 );
    not g16291 ( n15626 , n19484 );
    or g16292 ( n5370 , n4133 , n2335 );
    xnor g16293 ( n16500 , n7317 , n21471 );
    not g16294 ( n26327 , n12939 );
    or g16295 ( n16605 , n12021 , n7333 );
    xnor g16296 ( n9914 , n6255 , n21984 );
    and g16297 ( n21031 , n8136 , n14371 );
    or g16298 ( n18406 , n21853 , n17410 );
    xnor g16299 ( n12727 , n14616 , n10573 );
    xnor g16300 ( n7122 , n6915 , n18158 );
    or g16301 ( n1158 , n26907 , n26152 );
    xnor g16302 ( n6265 , n4997 , n9864 );
    and g16303 ( n25165 , n16650 , n4323 );
    nor g16304 ( n4892 , n18798 , n9332 );
    and g16305 ( n8221 , n276 , n15386 );
    and g16306 ( n19069 , n3286 , n785 );
    or g16307 ( n18448 , n3607 , n16463 );
    xnor g16308 ( n21661 , n13489 , n4913 );
    or g16309 ( n21202 , n9064 , n23446 );
    xnor g16310 ( n17269 , n11210 , n14637 );
    nor g16311 ( n3135 , n14545 , n18070 );
    or g16312 ( n13345 , n3495 , n9525 );
    not g16313 ( n21587 , n17016 );
    and g16314 ( n16328 , n19178 , n21147 );
    or g16315 ( n9555 , n22944 , n19249 );
    xnor g16316 ( n7652 , n7116 , n22569 );
    nor g16317 ( n26132 , n23528 , n10852 );
    xnor g16318 ( n3914 , n15752 , n10506 );
    or g16319 ( n24250 , n11116 , n2608 );
    and g16320 ( n12818 , n2744 , n7626 );
    xnor g16321 ( n5997 , n26951 , n27054 );
    nor g16322 ( n7831 , n16633 , n4622 );
    xnor g16323 ( n6879 , n3694 , n5302 );
    or g16324 ( n12429 , n1727 , n8595 );
    or g16325 ( n2358 , n16830 , n26741 );
    nor g16326 ( n9692 , n19134 , n18158 );
    xnor g16327 ( n7373 , n18542 , n25074 );
    xnor g16328 ( n18563 , n4136 , n4826 );
    and g16329 ( n4824 , n10762 , n26050 );
    and g16330 ( n2629 , n11980 , n19446 );
    and g16331 ( n23010 , n19494 , n1458 );
    not g16332 ( n22797 , n4005 );
    not g16333 ( n11848 , n17291 );
    not g16334 ( n22510 , n7072 );
    or g16335 ( n10806 , n85 , n10475 );
    and g16336 ( n14474 , n8327 , n13432 );
    or g16337 ( n15070 , n9076 , n25368 );
    and g16338 ( n20108 , n12017 , n15807 );
    and g16339 ( n13769 , n7926 , n27152 );
    xnor g16340 ( n7764 , n10622 , n12064 );
    or g16341 ( n12106 , n1021 , n11009 );
    or g16342 ( n4662 , n6356 , n4067 );
    and g16343 ( n13148 , n20544 , n12071 );
    and g16344 ( n4644 , n25175 , n18023 );
    xnor g16345 ( n15997 , n18676 , n24731 );
    or g16346 ( n16004 , n21873 , n22690 );
    and g16347 ( n25711 , n22564 , n18671 );
    xnor g16348 ( n9225 , n17010 , n19460 );
    and g16349 ( n2593 , n15648 , n18160 );
    xnor g16350 ( n2345 , n6185 , n10125 );
    not g16351 ( n4492 , n23950 );
    or g16352 ( n8828 , n13388 , n19318 );
    xnor g16353 ( n24030 , n23321 , n20429 );
    xnor g16354 ( n10288 , n15258 , n2420 );
    xnor g16355 ( n10093 , n1190 , n17852 );
    or g16356 ( n10667 , n6058 , n21056 );
    xnor g16357 ( n21732 , n19872 , n21462 );
    nor g16358 ( n3455 , n12341 , n22515 );
    xnor g16359 ( n8321 , n23654 , n19225 );
    xnor g16360 ( n12960 , n14432 , n10283 );
    xnor g16361 ( n10303 , n16247 , n23541 );
    nor g16362 ( n14025 , n10335 , n10141 );
    and g16363 ( n5958 , n1205 , n7494 );
    not g16364 ( n3608 , n757 );
    nor g16365 ( n1557 , n25639 , n21337 );
    or g16366 ( n24346 , n14624 , n5448 );
    xnor g16367 ( n24109 , n11270 , n10732 );
    and g16368 ( n5179 , n217 , n22165 );
    xnor g16369 ( n22778 , n5855 , n14576 );
    nor g16370 ( n22961 , n14532 , n17635 );
    and g16371 ( n9643 , n19679 , n26379 );
    or g16372 ( n21870 , n26238 , n10753 );
    or g16373 ( n20844 , n17734 , n10639 );
    and g16374 ( n4343 , n6619 , n12176 );
    xnor g16375 ( n14589 , n8176 , n8827 );
    xnor g16376 ( n3833 , n6640 , n25565 );
    xnor g16377 ( n9418 , n18415 , n2536 );
    nor g16378 ( n17510 , n25276 , n6137 );
    and g16379 ( n14430 , n19899 , n18608 );
    or g16380 ( n17961 , n8410 , n22826 );
    xnor g16381 ( n14010 , n6206 , n17409 );
    or g16382 ( n2114 , n11223 , n7710 );
    and g16383 ( n10812 , n7649 , n5864 );
    xnor g16384 ( n19457 , n26214 , n26103 );
    not g16385 ( n12229 , n7445 );
    nor g16386 ( n21676 , n3030 , n7407 );
    nor g16387 ( n10768 , n19177 , n26768 );
    nor g16388 ( n17103 , n3483 , n19556 );
    and g16389 ( n16116 , n9186 , n2716 );
    or g16390 ( n19207 , n5816 , n15780 );
    nor g16391 ( n22402 , n11195 , n20274 );
    or g16392 ( n18897 , n17054 , n24063 );
    and g16393 ( n11444 , n7748 , n26203 );
    and g16394 ( n7218 , n15448 , n24034 );
    or g16395 ( n19273 , n970 , n12292 );
    and g16396 ( n5488 , n5440 , n24366 );
    or g16397 ( n5239 , n5455 , n1530 );
    or g16398 ( n20430 , n6786 , n11872 );
    or g16399 ( n22739 , n3785 , n21 );
    xnor g16400 ( n22339 , n23354 , n2950 );
    or g16401 ( n1064 , n18746 , n17483 );
    or g16402 ( n3154 , n24049 , n16025 );
    or g16403 ( n9189 , n17063 , n5843 );
    and g16404 ( n15162 , n2416 , n16455 );
    and g16405 ( n6432 , n468 , n22322 );
    xnor g16406 ( n1972 , n5520 , n24977 );
    xnor g16407 ( n16125 , n26135 , n504 );
    not g16408 ( n26947 , n14048 );
    xnor g16409 ( n23820 , n11468 , n26604 );
    and g16410 ( n2473 , n11016 , n25036 );
    xnor g16411 ( n17496 , n7669 , n6218 );
    xnor g16412 ( n7464 , n20512 , n3260 );
    xnor g16413 ( n2266 , n12465 , n19575 );
    or g16414 ( n12662 , n25876 , n24541 );
    not g16415 ( n726 , n22082 );
    and g16416 ( n25051 , n20101 , n8705 );
    or g16417 ( n8294 , n21222 , n277 );
    or g16418 ( n18087 , n3033 , n22701 );
    and g16419 ( n26079 , n8106 , n10904 );
    not g16420 ( n26202 , n14467 );
    or g16421 ( n14859 , n11938 , n7162 );
    or g16422 ( n24240 , n14979 , n4957 );
    xnor g16423 ( n18241 , n9654 , n20523 );
    and g16424 ( n5985 , n13787 , n20545 );
    xnor g16425 ( n9700 , n3691 , n10272 );
    or g16426 ( n7182 , n15408 , n19111 );
    not g16427 ( n16019 , n2792 );
    not g16428 ( n19902 , n21749 );
    and g16429 ( n21817 , n3367 , n16063 );
    or g16430 ( n10091 , n19811 , n534 );
    or g16431 ( n22263 , n14874 , n22661 );
    or g16432 ( n19881 , n16576 , n10437 );
    or g16433 ( n10218 , n3403 , n24778 );
    not g16434 ( n6030 , n10772 );
    not g16435 ( n18202 , n22934 );
    xnor g16436 ( n3528 , n10226 , n9547 );
    not g16437 ( n7292 , n16988 );
    nor g16438 ( n22775 , n18157 , n26030 );
    or g16439 ( n12254 , n21270 , n19823 );
    xnor g16440 ( n8391 , n2040 , n23039 );
    not g16441 ( n4127 , n19377 );
    nor g16442 ( n4339 , n9108 , n8873 );
    or g16443 ( n21548 , n3438 , n25848 );
    and g16444 ( n14428 , n21524 , n18532 );
    and g16445 ( n22112 , n2508 , n17127 );
    or g16446 ( n6616 , n11525 , n19569 );
    nor g16447 ( n11899 , n1176 , n7254 );
    or g16448 ( n18237 , n4537 , n6446 );
    and g16449 ( n12580 , n9895 , n760 );
    xnor g16450 ( n25532 , n5250 , n18036 );
    or g16451 ( n6336 , n16995 , n25229 );
    not g16452 ( n22333 , n20512 );
    or g16453 ( n5208 , n8645 , n13365 );
    or g16454 ( n23421 , n14508 , n13778 );
    and g16455 ( n14241 , n19094 , n1197 );
    xnor g16456 ( n10483 , n17784 , n24085 );
    xnor g16457 ( n24926 , n21687 , n19922 );
    nor g16458 ( n5258 , n9990 , n7134 );
    or g16459 ( n17650 , n21245 , n12163 );
    and g16460 ( n26845 , n18814 , n802 );
    and g16461 ( n11346 , n26307 , n23799 );
    and g16462 ( n18052 , n25498 , n8132 );
    xnor g16463 ( n3282 , n14195 , n14580 );
    or g16464 ( n17469 , n2811 , n4239 );
    xnor g16465 ( n7635 , n16743 , n24485 );
    nor g16466 ( n561 , n4940 , n7609 );
    xnor g16467 ( n2829 , n12608 , n25323 );
    not g16468 ( n14982 , n12716 );
    or g16469 ( n13007 , n9944 , n20986 );
    nor g16470 ( n12337 , n23076 , n3509 );
    and g16471 ( n9577 , n4806 , n11883 );
    xnor g16472 ( n16243 , n22141 , n10858 );
    and g16473 ( n8289 , n23467 , n10772 );
    and g16474 ( n16281 , n11570 , n21103 );
    and g16475 ( n25088 , n19935 , n8195 );
    xnor g16476 ( n16496 , n10695 , n4794 );
    xnor g16477 ( n1697 , n16546 , n24283 );
    or g16478 ( n4802 , n22254 , n6733 );
    xnor g16479 ( n21856 , n12593 , n13714 );
    and g16480 ( n17515 , n23769 , n13747 );
    not g16481 ( n9076 , n19499 );
    xnor g16482 ( n4484 , n7125 , n24418 );
    and g16483 ( n13699 , n24279 , n6106 );
    and g16484 ( n26335 , n5253 , n20146 );
    xor g16485 ( n4425 , n286 , n7234 );
    and g16486 ( n5420 , n23837 , n4384 );
    or g16487 ( n3571 , n5783 , n2043 );
    xnor g16488 ( n16705 , n7414 , n18496 );
    not g16489 ( n4664 , n21638 );
    nor g16490 ( n23189 , n18035 , n12477 );
    or g16491 ( n19019 , n8454 , n1061 );
    xnor g16492 ( n7030 , n8616 , n3875 );
    not g16493 ( n106 , n16083 );
    xnor g16494 ( n14985 , n19658 , n15767 );
    xnor g16495 ( n5527 , n23770 , n16082 );
    not g16496 ( n1 , n3584 );
    and g16497 ( n4480 , n24395 , n1303 );
    xor g16498 ( n27078 , n5596 , n9427 );
    xnor g16499 ( n14164 , n25624 , n9653 );
    or g16500 ( n2735 , n16627 , n16393 );
    and g16501 ( n24930 , n12378 , n1072 );
    not g16502 ( n22743 , n26625 );
    or g16503 ( n19679 , n5006 , n23529 );
    or g16504 ( n4047 , n17403 , n13288 );
    or g16505 ( n10163 , n7175 , n22621 );
    xnor g16506 ( n12978 , n656 , n1007 );
    or g16507 ( n4496 , n24305 , n20231 );
    and g16508 ( n6625 , n15114 , n25699 );
    xnor g16509 ( n6232 , n25182 , n25211 );
    and g16510 ( n19887 , n25120 , n2903 );
    or g16511 ( n16832 , n21287 , n19981 );
    xnor g16512 ( n17190 , n12900 , n1255 );
    xnor g16513 ( n20352 , n26876 , n21997 );
    or g16514 ( n2190 , n20100 , n18720 );
    or g16515 ( n806 , n23054 , n22630 );
    xnor g16516 ( n8847 , n14290 , n19562 );
    xnor g16517 ( n23414 , n25689 , n6852 );
    not g16518 ( n636 , n6060 );
    and g16519 ( n7490 , n26854 , n19206 );
    and g16520 ( n20498 , n24417 , n10027 );
    and g16521 ( n23020 , n16139 , n2225 );
    or g16522 ( n22187 , n7296 , n3562 );
    and g16523 ( n9036 , n15089 , n16740 );
    xnor g16524 ( n15537 , n5682 , n3554 );
    or g16525 ( n8953 , n11249 , n25296 );
    xnor g16526 ( n24907 , n21139 , n2039 );
    not g16527 ( n15818 , n367 );
    nor g16528 ( n14478 , n14016 , n14102 );
    or g16529 ( n23494 , n6281 , n8661 );
    nor g16530 ( n13717 , n24314 , n9236 );
    or g16531 ( n7206 , n12422 , n12999 );
    not g16532 ( n9765 , n22986 );
    or g16533 ( n18949 , n23124 , n2136 );
    xnor g16534 ( n20058 , n6734 , n3 );
    or g16535 ( n3191 , n6959 , n19819 );
    and g16536 ( n18461 , n5006 , n7156 );
    or g16537 ( n4879 , n19027 , n12647 );
    xnor g16538 ( n24679 , n16968 , n21654 );
    or g16539 ( n23221 , n16917 , n938 );
    or g16540 ( n7784 , n3308 , n18623 );
    xnor g16541 ( n22399 , n12213 , n132 );
    xnor g16542 ( n17200 , n41 , n21718 );
    xnor g16543 ( n25415 , n17892 , n9915 );
    or g16544 ( n11389 , n6603 , n21263 );
    nor g16545 ( n2129 , n13040 , n23204 );
    nor g16546 ( n22306 , n12301 , n26467 );
    or g16547 ( n12903 , n11669 , n9561 );
    xnor g16548 ( n15366 , n14357 , n9714 );
    and g16549 ( n11216 , n19833 , n18178 );
    not g16550 ( n11814 , n10955 );
    and g16551 ( n22713 , n3606 , n24643 );
    and g16552 ( n13541 , n8074 , n22239 );
    or g16553 ( n21624 , n11092 , n6642 );
    not g16554 ( n24855 , n20646 );
    not g16555 ( n20954 , n6603 );
    xnor g16556 ( n5555 , n22876 , n18312 );
    xnor g16557 ( n7403 , n25315 , n21323 );
    or g16558 ( n14686 , n8270 , n5610 );
    xnor g16559 ( n18657 , n26667 , n3097 );
    not g16560 ( n2636 , n17169 );
    xnor g16561 ( n4748 , n7311 , n9399 );
    or g16562 ( n20115 , n25382 , n518 );
    and g16563 ( n2376 , n16366 , n18203 );
    or g16564 ( n19943 , n4236 , n6622 );
    or g16565 ( n3098 , n22968 , n17186 );
    xnor g16566 ( n4186 , n2127 , n2285 );
    and g16567 ( n17516 , n27059 , n23368 );
    xnor g16568 ( n19097 , n406 , n15297 );
    and g16569 ( n12097 , n10546 , n6052 );
    or g16570 ( n2216 , n8818 , n5171 );
    and g16571 ( n8212 , n14198 , n12902 );
    nor g16572 ( n14193 , n19177 , n23175 );
    xnor g16573 ( n23486 , n20817 , n27195 );
    nor g16574 ( n15655 , n3460 , n24774 );
    and g16575 ( n24059 , n22034 , n2110 );
    and g16576 ( n18248 , n25478 , n22143 );
    and g16577 ( n26617 , n19984 , n26978 );
    xnor g16578 ( n7023 , n14663 , n20247 );
    or g16579 ( n17294 , n8707 , n2807 );
    or g16580 ( n8683 , n3995 , n26333 );
    xnor g16581 ( n17901 , n11448 , n1391 );
    or g16582 ( n7533 , n5276 , n16810 );
    xnor g16583 ( n22076 , n13589 , n12476 );
    or g16584 ( n25457 , n16129 , n396 );
    and g16585 ( n25564 , n6645 , n17379 );
    not g16586 ( n1562 , n3245 );
    xnor g16587 ( n9441 , n8381 , n23775 );
    or g16588 ( n21890 , n20429 , n14922 );
    or g16589 ( n17627 , n12671 , n15196 );
    nor g16590 ( n12505 , n21272 , n3015 );
    not g16591 ( n14721 , n23568 );
    or g16592 ( n20746 , n20821 , n7972 );
    or g16593 ( n13077 , n14438 , n13265 );
    nor g16594 ( n2469 , n24031 , n6204 );
    not g16595 ( n26149 , n19104 );
    not g16596 ( n14337 , n4964 );
    or g16597 ( n22842 , n21088 , n11247 );
    or g16598 ( n13012 , n7025 , n7706 );
    xnor g16599 ( n21785 , n1689 , n17095 );
    or g16600 ( n7166 , n4854 , n23862 );
    and g16601 ( n4438 , n22579 , n18834 );
    or g16602 ( n3886 , n7605 , n13518 );
    xnor g16603 ( n4042 , n4447 , n16786 );
    not g16604 ( n24868 , n8845 );
    not g16605 ( n5402 , n2173 );
    xnor g16606 ( n4759 , n5270 , n610 );
    and g16607 ( n22344 , n20406 , n24013 );
    xnor g16608 ( n21508 , n4428 , n17140 );
    or g16609 ( n12501 , n20923 , n7983 );
    xnor g16610 ( n23819 , n14629 , n17244 );
    xnor g16611 ( n9552 , n1375 , n10447 );
    nor g16612 ( n11791 , n13359 , n1 );
    or g16613 ( n21866 , n8423 , n358 );
    xnor g16614 ( n20719 , n931 , n3792 );
    and g16615 ( n16685 , n2008 , n21478 );
    or g16616 ( n17921 , n11993 , n8541 );
    or g16617 ( n15912 , n21236 , n23738 );
    or g16618 ( n26987 , n20070 , n11222 );
    not g16619 ( n8076 , n4923 );
    not g16620 ( n13725 , n27102 );
    not g16621 ( n20329 , n3349 );
    and g16622 ( n25404 , n3098 , n21296 );
    xnor g16623 ( n19098 , n25178 , n25103 );
    xnor g16624 ( n13844 , n23037 , n21409 );
    or g16625 ( n21197 , n21435 , n9643 );
    xnor g16626 ( n24097 , n14333 , n9532 );
    nor g16627 ( n11785 , n18333 , n20316 );
    xnor g16628 ( n2885 , n5471 , n12679 );
    nor g16629 ( n12591 , n22254 , n8067 );
    or g16630 ( n16180 , n18514 , n25261 );
    or g16631 ( n7774 , n4053 , n13846 );
    or g16632 ( n7113 , n25109 , n7187 );
    xnor g16633 ( n17900 , n9010 , n5707 );
    xnor g16634 ( n18933 , n27111 , n24701 );
    xnor g16635 ( n4294 , n6515 , n3282 );
    or g16636 ( n16478 , n5132 , n18146 );
    nor g16637 ( n12743 , n11060 , n25249 );
    not g16638 ( n16611 , n23264 );
    or g16639 ( n13724 , n1265 , n18308 );
    or g16640 ( n24174 , n21281 , n20656 );
    or g16641 ( n1157 , n11393 , n5580 );
    xnor g16642 ( n16183 , n9799 , n414 );
    or g16643 ( n9578 , n11968 , n20958 );
    and g16644 ( n9751 , n24205 , n6069 );
    xnor g16645 ( n9928 , n26234 , n23033 );
    and g16646 ( n16194 , n2707 , n6755 );
    and g16647 ( n20785 , n10221 , n9052 );
    or g16648 ( n936 , n12017 , n15807 );
    or g16649 ( n24971 , n19915 , n21985 );
    not g16650 ( n8477 , n19060 );
    or g16651 ( n23219 , n21113 , n21945 );
    nor g16652 ( n25588 , n22527 , n24032 );
    xnor g16653 ( n3352 , n4384 , n21778 );
    xnor g16654 ( n7891 , n24383 , n6403 );
    and g16655 ( n23110 , n5620 , n23814 );
    xnor g16656 ( n21357 , n14040 , n24711 );
    or g16657 ( n21190 , n12375 , n17003 );
    xnor g16658 ( n26528 , n6429 , n20757 );
    and g16659 ( n15351 , n5670 , n1800 );
    or g16660 ( n4214 , n8419 , n24580 );
    or g16661 ( n22799 , n7019 , n17649 );
    and g16662 ( n2178 , n19551 , n2705 );
    and g16663 ( n16653 , n1776 , n17962 );
    nor g16664 ( n7997 , n19184 , n14661 );
    xnor g16665 ( n409 , n22309 , n19107 );
    or g16666 ( n7542 , n18517 , n15759 );
    and g16667 ( n13820 , n871 , n7412 );
    or g16668 ( n8666 , n8254 , n17874 );
    or g16669 ( n26516 , n940 , n8462 );
    xnor g16670 ( n12880 , n14484 , n21617 );
    and g16671 ( n815 , n11343 , n23618 );
    or g16672 ( n17970 , n488 , n5121 );
    xnor g16673 ( n13625 , n25675 , n21477 );
    and g16674 ( n11372 , n2737 , n24303 );
    nor g16675 ( n14707 , n647 , n26408 );
    xnor g16676 ( n1599 , n6643 , n21252 );
    xnor g16677 ( n19720 , n19789 , n21226 );
    not g16678 ( n5715 , n7841 );
    xnor g16679 ( n2164 , n12457 , n11758 );
    not g16680 ( n14651 , n10093 );
    not g16681 ( n12014 , n23493 );
    and g16682 ( n8063 , n26272 , n3184 );
    not g16683 ( n2060 , n10629 );
    or g16684 ( n25179 , n23345 , n26788 );
    xnor g16685 ( n12194 , n1594 , n762 );
    not g16686 ( n16421 , n16410 );
    or g16687 ( n14662 , n17960 , n7418 );
    xnor g16688 ( n14661 , n24931 , n7890 );
    not g16689 ( n3454 , n14466 );
    xnor g16690 ( n410 , n1510 , n24150 );
    nor g16691 ( n25879 , n11743 , n13301 );
    or g16692 ( n3888 , n19558 , n4648 );
    or g16693 ( n9349 , n23477 , n1334 );
    or g16694 ( n5041 , n1694 , n8206 );
    or g16695 ( n6059 , n2146 , n20216 );
    and g16696 ( n13674 , n21674 , n5090 );
    xnor g16697 ( n11476 , n8696 , n1593 );
    xnor g16698 ( n23366 , n23041 , n6172 );
    xnor g16699 ( n15817 , n18163 , n21784 );
    and g16700 ( n8534 , n24452 , n13528 );
    and g16701 ( n9339 , n370 , n23022 );
    or g16702 ( n17513 , n23244 , n23842 );
    nor g16703 ( n6247 , n15801 , n26047 );
    and g16704 ( n18978 , n2237 , n20475 );
    nor g16705 ( n22271 , n23207 , n15930 );
    or g16706 ( n26772 , n23800 , n3445 );
    xnor g16707 ( n15397 , n7524 , n15967 );
    and g16708 ( n19280 , n18844 , n17107 );
    not g16709 ( n25676 , n25054 );
    xnor g16710 ( n21008 , n18855 , n20218 );
    and g16711 ( n26893 , n8770 , n2286 );
    or g16712 ( n13666 , n27046 , n24125 );
    buf g16713 ( n19313 , n6678 );
    or g16714 ( n25379 , n22365 , n11356 );
    xnor g16715 ( n26006 , n3062 , n11185 );
    or g16716 ( n12794 , n1220 , n13950 );
    not g16717 ( n18257 , n3030 );
    nor g16718 ( n9813 , n22729 , n21698 );
    or g16719 ( n14828 , n6712 , n26501 );
    xnor g16720 ( n5377 , n17412 , n22562 );
    nor g16721 ( n23866 , n9246 , n23120 );
    and g16722 ( n10276 , n25246 , n24728 );
    xnor g16723 ( n7864 , n22571 , n11792 );
    xnor g16724 ( n307 , n18149 , n19103 );
    nor g16725 ( n15856 , n17549 , n4095 );
    xnor g16726 ( n10305 , n21764 , n23900 );
    not g16727 ( n3009 , n13137 );
    not g16728 ( n20145 , n448 );
    nor g16729 ( n19712 , n933 , n5378 );
    or g16730 ( n21835 , n22759 , n19066 );
    not g16731 ( n11919 , n20700 );
    xnor g16732 ( n23587 , n7429 , n9323 );
    or g16733 ( n8872 , n10008 , n27025 );
    not g16734 ( n18785 , n8207 );
    not g16735 ( n5743 , n20176 );
    and g16736 ( n19823 , n6889 , n2648 );
    nor g16737 ( n13992 , n11583 , n17959 );
    xnor g16738 ( n20603 , n15918 , n21735 );
    or g16739 ( n16362 , n19041 , n21006 );
    xnor g16740 ( n20788 , n14279 , n6921 );
    not g16741 ( n14943 , n7568 );
    or g16742 ( n18259 , n24877 , n26549 );
    and g16743 ( n10412 , n22171 , n12283 );
    and g16744 ( n24986 , n11852 , n15037 );
    xnor g16745 ( n8292 , n17924 , n27098 );
    nor g16746 ( n1673 , n11408 , n15787 );
    xnor g16747 ( n11376 , n6262 , n945 );
    nor g16748 ( n25669 , n7692 , n25464 );
    not g16749 ( n10410 , n1050 );
    or g16750 ( n24669 , n21702 , n7815 );
    or g16751 ( n23377 , n7664 , n13678 );
    nor g16752 ( n12698 , n27142 , n9312 );
    xnor g16753 ( n26900 , n12523 , n4454 );
    nor g16754 ( n17014 , n3324 , n4299 );
    and g16755 ( n5043 , n13977 , n14650 );
    and g16756 ( n25790 , n10137 , n26298 );
    or g16757 ( n24094 , n22138 , n10086 );
    and g16758 ( n19034 , n12280 , n24520 );
    xnor g16759 ( n15002 , n24598 , n22326 );
    not g16760 ( n12699 , n18052 );
    nor g16761 ( n24041 , n20542 , n9575 );
    xnor g16762 ( n18532 , n6645 , n7050 );
    xnor g16763 ( n2021 , n22173 , n24032 );
    or g16764 ( n8273 , n24171 , n11671 );
    or g16765 ( n509 , n15973 , n21631 );
    nor g16766 ( n12940 , n19025 , n9655 );
    or g16767 ( n9062 , n14442 , n2634 );
    and g16768 ( n634 , n18214 , n900 );
    and g16769 ( n18789 , n12871 , n8888 );
    xnor g16770 ( n9510 , n455 , n3603 );
    or g16771 ( n20576 , n18452 , n3118 );
    xnor g16772 ( n18181 , n10408 , n14899 );
    xnor g16773 ( n2390 , n21710 , n25237 );
    or g16774 ( n9819 , n16236 , n20019 );
    or g16775 ( n17904 , n25972 , n3707 );
    and g16776 ( n6238 , n8782 , n24561 );
    xnor g16777 ( n15299 , n23114 , n3454 );
    xnor g16778 ( n6891 , n8000 , n22156 );
    and g16779 ( n23847 , n2754 , n9195 );
    not g16780 ( n9107 , n22591 );
    or g16781 ( n2026 , n25156 , n2073 );
    xnor g16782 ( n13846 , n10792 , n19922 );
    xnor g16783 ( n10767 , n4617 , n24261 );
    not g16784 ( n16890 , n1682 );
    and g16785 ( n7673 , n12882 , n3325 );
    xnor g16786 ( n18439 , n4949 , n14170 );
    not g16787 ( n20479 , n24612 );
    or g16788 ( n9644 , n9172 , n10571 );
    or g16789 ( n25788 , n27114 , n3247 );
    not g16790 ( n1062 , n21906 );
    nor g16791 ( n10771 , n23230 , n10053 );
    xnor g16792 ( n9287 , n3859 , n21603 );
    and g16793 ( n4944 , n7912 , n18949 );
    xnor g16794 ( n26860 , n6064 , n4405 );
    xnor g16795 ( n24612 , n3994 , n19228 );
    or g16796 ( n1229 , n24928 , n18187 );
    nor g16797 ( n3927 , n3981 , n24818 );
    or g16798 ( n26737 , n25188 , n1042 );
    or g16799 ( n1874 , n9149 , n23564 );
    or g16800 ( n15208 , n19804 , n13567 );
    nor g16801 ( n5887 , n7693 , n9453 );
    xnor g16802 ( n4300 , n10158 , n3952 );
    xnor g16803 ( n24568 , n5925 , n9058 );
    or g16804 ( n452 , n8192 , n26716 );
    not g16805 ( n2915 , n11481 );
    xnor g16806 ( n6271 , n23439 , n7573 );
    and g16807 ( n10440 , n19689 , n16384 );
    or g16808 ( n2662 , n19797 , n21497 );
    xnor g16809 ( n685 , n1328 , n13987 );
    xnor g16810 ( n4745 , n8915 , n27067 );
    and g16811 ( n9781 , n13838 , n3357 );
    or g16812 ( n8038 , n9326 , n1466 );
    not g16813 ( n6327 , n6283 );
    or g16814 ( n2273 , n16588 , n27047 );
    or g16815 ( n5663 , n23250 , n16856 );
    and g16816 ( n6738 , n17748 , n47 );
    nor g16817 ( n20909 , n22327 , n4559 );
    xnor g16818 ( n407 , n15720 , n18512 );
    or g16819 ( n10752 , n22365 , n20429 );
    xnor g16820 ( n10538 , n21998 , n25779 );
    xnor g16821 ( n9702 , n19366 , n11184 );
    or g16822 ( n2396 , n5794 , n12744 );
    not g16823 ( n27172 , n14386 );
    not g16824 ( n19321 , n12121 );
    and g16825 ( n14192 , n11177 , n10254 );
    or g16826 ( n24173 , n193 , n19415 );
    nor g16827 ( n12238 , n1802 , n7331 );
    not g16828 ( n17938 , n11688 );
    or g16829 ( n9103 , n19161 , n7966 );
    not g16830 ( n15661 , n7940 );
    and g16831 ( n5721 , n2118 , n19960 );
    xnor g16832 ( n5677 , n10763 , n5696 );
    not g16833 ( n22206 , n4714 );
    and g16834 ( n21884 , n8601 , n23815 );
    and g16835 ( n14824 , n15207 , n21787 );
    xnor g16836 ( n10019 , n22806 , n19972 );
    xnor g16837 ( n12659 , n12090 , n12018 );
    xnor g16838 ( n20005 , n7540 , n7944 );
    and g16839 ( n1244 , n238 , n24333 );
    xnor g16840 ( n26609 , n18263 , n12475 );
    xnor g16841 ( n25884 , n8661 , n8496 );
    or g16842 ( n17016 , n16551 , n19166 );
    or g16843 ( n7494 , n12543 , n4934 );
    or g16844 ( n17144 , n4490 , n1949 );
    xnor g16845 ( n27031 , n22564 , n772 );
    xnor g16846 ( n16859 , n23558 , n12421 );
    or g16847 ( n5748 , n5434 , n10074 );
    nor g16848 ( n16168 , n18173 , n5101 );
    not g16849 ( n25942 , n22850 );
    or g16850 ( n21153 , n19 , n26673 );
    and g16851 ( n1911 , n24575 , n15232 );
    or g16852 ( n8263 , n11256 , n745 );
    or g16853 ( n4394 , n2413 , n10449 );
    xnor g16854 ( n16696 , n21058 , n9111 );
    not g16855 ( n4818 , n21361 );
    xnor g16856 ( n7145 , n14016 , n14102 );
    nor g16857 ( n25536 , n16626 , n1998 );
    nor g16858 ( n23640 , n14089 , n15930 );
    and g16859 ( n6526 , n4311 , n11660 );
    or g16860 ( n1614 , n20476 , n6159 );
    nor g16861 ( n14523 , n24475 , n14749 );
    and g16862 ( n21481 , n442 , n6319 );
    or g16863 ( n12588 , n2505 , n6969 );
    nor g16864 ( n24524 , n16091 , n16602 );
    not g16865 ( n2391 , n14091 );
    xnor g16866 ( n5349 , n5563 , n20239 );
    xnor g16867 ( n13235 , n21280 , n24364 );
    or g16868 ( n11265 , n21471 , n22014 );
    and g16869 ( n16005 , n11180 , n20510 );
    and g16870 ( n24878 , n8499 , n8388 );
    not g16871 ( n10258 , n7612 );
    nor g16872 ( n13796 , n12014 , n8405 );
    xnor g16873 ( n11225 , n13494 , n18880 );
    xnor g16874 ( n6128 , n3686 , n21155 );
    and g16875 ( n14836 , n675 , n14934 );
    and g16876 ( n14804 , n16996 , n22025 );
    xnor g16877 ( n7108 , n22428 , n1269 );
    nor g16878 ( n11521 , n6753 , n8779 );
    or g16879 ( n7704 , n9679 , n13405 );
    and g16880 ( n5232 , n4619 , n10901 );
    xnor g16881 ( n12707 , n8817 , n19583 );
    xnor g16882 ( n23731 , n22904 , n19571 );
    and g16883 ( n8287 , n13600 , n14108 );
    nor g16884 ( n15361 , n7785 , n8853 );
    or g16885 ( n15597 , n18253 , n5756 );
    or g16886 ( n18762 , n14344 , n6521 );
    or g16887 ( n8143 , n14569 , n24049 );
    nor g16888 ( n9784 , n9768 , n16276 );
    not g16889 ( n3675 , n4723 );
    xnor g16890 ( n27011 , n24773 , n7492 );
    and g16891 ( n14504 , n11583 , n14085 );
    or g16892 ( n22037 , n20905 , n8670 );
    and g16893 ( n17819 , n23528 , n10852 );
    xnor g16894 ( n16703 , n16722 , n13708 );
    or g16895 ( n7748 , n21213 , n4685 );
    not g16896 ( n1433 , n7002 );
    and g16897 ( n16504 , n19881 , n11532 );
    or g16898 ( n24248 , n8076 , n22031 );
    xnor g16899 ( n14200 , n5559 , n26036 );
    not g16900 ( n6093 , n22435 );
    not g16901 ( n24584 , n13085 );
    not g16902 ( n1890 , n25312 );
    nor g16903 ( n4769 , n21073 , n15975 );
    xnor g16904 ( n13094 , n6632 , n1831 );
    and g16905 ( n21348 , n14123 , n2494 );
    or g16906 ( n16485 , n26312 , n17453 );
    xnor g16907 ( n2758 , n26065 , n13136 );
    xnor g16908 ( n8769 , n8704 , n15596 );
    xnor g16909 ( n9972 , n16737 , n10342 );
    or g16910 ( n10110 , n6709 , n24386 );
    not g16911 ( n11030 , n5028 );
    or g16912 ( n20298 , n23695 , n854 );
    nor g16913 ( n11410 , n22688 , n3474 );
    xnor g16914 ( n26557 , n7336 , n11105 );
    nor g16915 ( n4365 , n26408 , n12477 );
    and g16916 ( n4415 , n4614 , n15132 );
    or g16917 ( n24337 , n25749 , n22082 );
    or g16918 ( n25598 , n18386 , n6689 );
    or g16919 ( n11678 , n2688 , n8163 );
    or g16920 ( n7434 , n16465 , n5709 );
    not g16921 ( n14401 , n20104 );
    xnor g16922 ( n1722 , n13936 , n11201 );
    or g16923 ( n21799 , n23835 , n10947 );
    or g16924 ( n1128 , n23932 , n2606 );
    xnor g16925 ( n13003 , n20754 , n593 );
    not g16926 ( n8071 , n13915 );
    xnor g16927 ( n1195 , n16966 , n14796 );
    or g16928 ( n21411 , n15938 , n5747 );
    or g16929 ( n14896 , n4799 , n11411 );
    and g16930 ( n9288 , n3974 , n717 );
    and g16931 ( n386 , n23281 , n5142 );
    and g16932 ( n25231 , n24687 , n23301 );
    xnor g16933 ( n24728 , n10953 , n2734 );
    nor g16934 ( n20214 , n1118 , n20489 );
    xnor g16935 ( n8025 , n22686 , n15464 );
    or g16936 ( n14990 , n22536 , n22955 );
    or g16937 ( n15207 , n13360 , n16724 );
    or g16938 ( n15459 , n8532 , n22685 );
    and g16939 ( n22754 , n14337 , n24865 );
    or g16940 ( n21149 , n5968 , n5180 );
    nor g16941 ( n10443 , n25119 , n12652 );
    or g16942 ( n24577 , n15890 , n1384 );
    and g16943 ( n11320 , n15235 , n10545 );
    not g16944 ( n25700 , n7538 );
    and g16945 ( n23346 , n11505 , n24352 );
    and g16946 ( n3586 , n20044 , n11835 );
    and g16947 ( n22483 , n4809 , n6114 );
    not g16948 ( n17579 , n1831 );
    not g16949 ( n4017 , n10873 );
    not g16950 ( n17716 , n23820 );
    xnor g16951 ( n25525 , n8455 , n24835 );
    and g16952 ( n23136 , n26342 , n26906 );
    or g16953 ( n26697 , n10840 , n14914 );
    xnor g16954 ( n6013 , n20608 , n6195 );
    or g16955 ( n13864 , n15054 , n25031 );
    not g16956 ( n4032 , n10652 );
    or g16957 ( n26570 , n9526 , n25349 );
    and g16958 ( n17648 , n4200 , n19302 );
    nor g16959 ( n6641 , n14139 , n24152 );
    or g16960 ( n26347 , n10151 , n5324 );
    and g16961 ( n19809 , n716 , n15543 );
    or g16962 ( n26591 , n10090 , n16377 );
    and g16963 ( n30 , n11058 , n14616 );
    nor g16964 ( n10671 , n12375 , n22765 );
    and g16965 ( n2781 , n8574 , n22188 );
    and g16966 ( n8222 , n19327 , n25624 );
    xnor g16967 ( n5940 , n12821 , n5579 );
    xnor g16968 ( n2443 , n17964 , n20651 );
    nor g16969 ( n131 , n1262 , n9557 );
    xnor g16970 ( n7567 , n6037 , n5376 );
    and g16971 ( n6993 , n867 , n11341 );
    xnor g16972 ( n16011 , n11751 , n3245 );
    xnor g16973 ( n13400 , n22965 , n19791 );
    xnor g16974 ( n9867 , n24279 , n3296 );
    and g16975 ( n25549 , n26091 , n17349 );
    nor g16976 ( n18370 , n23686 , n8084 );
    xnor g16977 ( n8826 , n22480 , n7020 );
    and g16978 ( n24516 , n24684 , n12880 );
    xnor g16979 ( n17314 , n14845 , n2274 );
    nor g16980 ( n14717 , n13872 , n14279 );
    xnor g16981 ( n26594 , n24813 , n9396 );
    xnor g16982 ( n2058 , n3123 , n4393 );
    and g16983 ( n26031 , n0 , n22796 );
    or g16984 ( n5089 , n930 , n2638 );
    xnor g16985 ( n8545 , n11336 , n10201 );
    nor g16986 ( n811 , n22375 , n5722 );
    or g16987 ( n7625 , n8979 , n13263 );
    not g16988 ( n22234 , n15384 );
    and g16989 ( n20580 , n22889 , n24790 );
    xnor g16990 ( n12975 , n26056 , n27151 );
    and g16991 ( n23696 , n13335 , n11547 );
    or g16992 ( n6310 , n10964 , n17159 );
    xnor g16993 ( n24916 , n15456 , n18880 );
    xnor g16994 ( n2374 , n7908 , n12723 );
    or g16995 ( n12854 , n24077 , n17615 );
    nor g16996 ( n7423 , n2055 , n17938 );
    and g16997 ( n12613 , n2415 , n8414 );
    xnor g16998 ( n25241 , n25753 , n26018 );
    xnor g16999 ( n8271 , n1731 , n16430 );
    xnor g17000 ( n25561 , n9881 , n12741 );
    nor g17001 ( n19733 , n12153 , n9490 );
    not g17002 ( n24649 , n19608 );
    not g17003 ( n22285 , n12098 );
    or g17004 ( n8758 , n25282 , n10577 );
    or g17005 ( n27085 , n17892 , n3371 );
    not g17006 ( n6170 , n2548 );
    xnor g17007 ( n25602 , n27156 , n3909 );
    not g17008 ( n12416 , n25316 );
    xnor g17009 ( n24518 , n8439 , n3710 );
    xnor g17010 ( n23692 , n2823 , n3630 );
    not g17011 ( n9237 , n9931 );
    and g17012 ( n8278 , n9586 , n12778 );
    or g17013 ( n12372 , n8797 , n23485 );
    not g17014 ( n3280 , n2574 );
    xnor g17015 ( n6149 , n10217 , n11011 );
    xnor g17016 ( n16584 , n3023 , n14320 );
    and g17017 ( n9708 , n10497 , n6656 );
    not g17018 ( n17203 , n17255 );
    not g17019 ( n11039 , n20389 );
    nor g17020 ( n13227 , n10324 , n13719 );
    and g17021 ( n10400 , n15367 , n8350 );
    xnor g17022 ( n25323 , n10593 , n1662 );
    xnor g17023 ( n2101 , n16496 , n17647 );
    not g17024 ( n22987 , n655 );
    or g17025 ( n13634 , n24599 , n12766 );
    xnor g17026 ( n6949 , n5606 , n1698 );
    nor g17027 ( n25634 , n18788 , n15288 );
    or g17028 ( n2493 , n10835 , n7490 );
    xnor g17029 ( n13543 , n14090 , n18962 );
    xnor g17030 ( n19162 , n7530 , n4189 );
    xnor g17031 ( n7069 , n23851 , n4100 );
    or g17032 ( n21443 , n18537 , n10920 );
    and g17033 ( n24747 , n19451 , n25828 );
    or g17034 ( n20846 , n8467 , n4128 );
    or g17035 ( n24893 , n7081 , n24213 );
    xnor g17036 ( n16375 , n10962 , n16789 );
    not g17037 ( n22962 , n6631 );
    nor g17038 ( n16806 , n20365 , n8083 );
    or g17039 ( n22010 , n2590 , n21901 );
    or g17040 ( n11951 , n682 , n5075 );
    xnor g17041 ( n18756 , n20719 , n22918 );
    or g17042 ( n8698 , n20040 , n16555 );
    or g17043 ( n22598 , n20324 , n810 );
    and g17044 ( n18250 , n21977 , n8817 );
    and g17045 ( n12033 , n22500 , n21601 );
    xnor g17046 ( n17592 , n6615 , n22493 );
    nor g17047 ( n2192 , n11958 , n1036 );
    xnor g17048 ( n20691 , n23759 , n13984 );
    and g17049 ( n18334 , n2976 , n10904 );
    not g17050 ( n24074 , n10854 );
    not g17051 ( n7520 , n6834 );
    not g17052 ( n14539 , n14215 );
    not g17053 ( n874 , n3919 );
    not g17054 ( n7933 , n7516 );
    and g17055 ( n23827 , n13153 , n9230 );
    xnor g17056 ( n1431 , n18974 , n26380 );
    not g17057 ( n26805 , n2099 );
    or g17058 ( n16726 , n12551 , n23442 );
    or g17059 ( n11817 , n1999 , n766 );
    xnor g17060 ( n12730 , n23877 , n9830 );
    not g17061 ( n64 , n18815 );
    xnor g17062 ( n16707 , n912 , n5131 );
    not g17063 ( n13960 , n12236 );
    nor g17064 ( n24435 , n10505 , n6925 );
    and g17065 ( n10550 , n13229 , n18670 );
    and g17066 ( n11915 , n20358 , n3960 );
    xnor g17067 ( n10032 , n16038 , n18794 );
    nor g17068 ( n24904 , n15405 , n3940 );
    not g17069 ( n10837 , n19680 );
    xnor g17070 ( n25053 , n12488 , n1437 );
    and g17071 ( n10702 , n22547 , n10428 );
    nor g17072 ( n7504 , n26458 , n6073 );
    nor g17073 ( n20708 , n13915 , n23644 );
    not g17074 ( n2346 , n5899 );
    xnor g17075 ( n8448 , n14291 , n20285 );
    xnor g17076 ( n3263 , n1554 , n21397 );
    xnor g17077 ( n24480 , n7860 , n13719 );
    or g17078 ( n9272 , n2329 , n2753 );
    xnor g17079 ( n14917 , n3990 , n5349 );
    buf g17080 ( n10557 , n12322 );
    xnor g17081 ( n5866 , n20384 , n8008 );
    not g17082 ( n4155 , n13502 );
    xnor g17083 ( n7479 , n19227 , n8381 );
    and g17084 ( n21568 , n25836 , n23569 );
    or g17085 ( n20067 , n24157 , n1910 );
    and g17086 ( n19431 , n25234 , n9405 );
    nor g17087 ( n19880 , n2156 , n5796 );
    xnor g17088 ( n22850 , n21851 , n20868 );
    xnor g17089 ( n15861 , n7339 , n26808 );
    xnor g17090 ( n16923 , n21678 , n24616 );
    xnor g17091 ( n23058 , n6126 , n1420 );
    xnor g17092 ( n14153 , n17876 , n17508 );
    nor g17093 ( n14563 , n27104 , n13317 );
    nor g17094 ( n3518 , n212 , n9928 );
    not g17095 ( n5283 , n26667 );
    not g17096 ( n18114 , n5976 );
    and g17097 ( n7207 , n20568 , n9861 );
    xnor g17098 ( n18553 , n1798 , n8930 );
    or g17099 ( n1930 , n16022 , n1519 );
    xnor g17100 ( n755 , n7574 , n16675 );
    or g17101 ( n26198 , n21450 , n4870 );
    xnor g17102 ( n6179 , n5092 , n19270 );
    or g17103 ( n10481 , n11798 , n7509 );
    xnor g17104 ( n23151 , n2481 , n9477 );
    xnor g17105 ( n9527 , n17022 , n9506 );
    xnor g17106 ( n13654 , n7752 , n12541 );
    not g17107 ( n15109 , n15146 );
    or g17108 ( n15350 , n446 , n13349 );
    or g17109 ( n19801 , n20071 , n12026 );
    not g17110 ( n17366 , n18790 );
    nor g17111 ( n17738 , n5890 , n22838 );
    or g17112 ( n26396 , n10417 , n8362 );
    xnor g17113 ( n21385 , n12474 , n15713 );
    or g17114 ( n25443 , n20921 , n22552 );
    xnor g17115 ( n12313 , n23962 , n2274 );
    xnor g17116 ( n25808 , n21585 , n23146 );
    or g17117 ( n12595 , n2354 , n8940 );
    xnor g17118 ( n7890 , n19282 , n26986 );
    and g17119 ( n7601 , n3285 , n21463 );
    or g17120 ( n3624 , n1665 , n19269 );
    xnor g17121 ( n21093 , n15800 , n3772 );
    or g17122 ( n18490 , n7384 , n6931 );
    or g17123 ( n24308 , n12708 , n9529 );
    and g17124 ( n15754 , n14605 , n22010 );
    not g17125 ( n12111 , n14382 );
    xnor g17126 ( n17854 , n2867 , n20756 );
    not g17127 ( n9584 , n15910 );
    xnor g17128 ( n23748 , n8811 , n645 );
    xnor g17129 ( n3653 , n19155 , n27192 );
    or g17130 ( n22429 , n2372 , n12347 );
    not g17131 ( n198 , n9028 );
    xnor g17132 ( n21189 , n25160 , n18290 );
    nor g17133 ( n25400 , n7818 , n13851 );
    xnor g17134 ( n16166 , n25403 , n22973 );
    not g17135 ( n25509 , n4345 );
    or g17136 ( n13550 , n11144 , n11640 );
    not g17137 ( n7697 , n9527 );
    and g17138 ( n14028 , n25348 , n7153 );
    and g17139 ( n14116 , n17844 , n1962 );
    nor g17140 ( n18099 , n8107 , n18363 );
    or g17141 ( n15163 , n13901 , n4860 );
    not g17142 ( n18841 , n26703 );
    xnor g17143 ( n11451 , n15626 , n5302 );
    or g17144 ( n2439 , n4178 , n16763 );
    or g17145 ( n15731 , n12276 , n22992 );
    xnor g17146 ( n17820 , n8034 , n19724 );
    and g17147 ( n17259 , n9839 , n6754 );
    xnor g17148 ( n5105 , n4599 , n7305 );
    or g17149 ( n14837 , n15643 , n3393 );
    or g17150 ( n10968 , n14132 , n3338 );
    and g17151 ( n13571 , n378 , n5779 );
    and g17152 ( n18264 , n3840 , n24908 );
    and g17153 ( n12750 , n21516 , n26336 );
    and g17154 ( n15076 , n14323 , n12351 );
    not g17155 ( n18100 , n13319 );
    xnor g17156 ( n22017 , n21116 , n1448 );
    xnor g17157 ( n14637 , n21725 , n19283 );
    or g17158 ( n18306 , n9976 , n13702 );
    xnor g17159 ( n14330 , n13006 , n15092 );
    not g17160 ( n4442 , n6037 );
    nor g17161 ( n24462 , n11938 , n8244 );
    nor g17162 ( n10002 , n24244 , n11577 );
    or g17163 ( n15250 , n9826 , n26505 );
    not g17164 ( n8910 , n3925 );
    or g17165 ( n15117 , n7172 , n19806 );
    or g17166 ( n12600 , n9910 , n20342 );
    not g17167 ( n12868 , n4429 );
    nor g17168 ( n15504 , n11303 , n23200 );
    and g17169 ( n19639 , n19340 , n234 );
    xnor g17170 ( n4288 , n10328 , n7579 );
    xnor g17171 ( n21637 , n11206 , n6840 );
    xnor g17172 ( n8338 , n19929 , n23787 );
    or g17173 ( n3087 , n18067 , n2333 );
    not g17174 ( n15502 , n20391 );
    or g17175 ( n24279 , n18852 , n20815 );
    xnor g17176 ( n5351 , n51 , n21513 );
    xnor g17177 ( n18043 , n19591 , n22667 );
    or g17178 ( n8574 , n10159 , n14790 );
    not g17179 ( n7311 , n2088 );
    or g17180 ( n15419 , n11831 , n14777 );
    not g17181 ( n20880 , n7721 );
    and g17182 ( n23781 , n18649 , n11278 );
    and g17183 ( n5944 , n21325 , n27069 );
    and g17184 ( n7161 , n12143 , n20215 );
    or g17185 ( n5896 , n12359 , n22528 );
    and g17186 ( n17358 , n14027 , n23421 );
    xnor g17187 ( n19146 , n6170 , n5115 );
    xnor g17188 ( n10101 , n15510 , n22496 );
    or g17189 ( n23549 , n25218 , n5527 );
    nor g17190 ( n883 , n26951 , n27054 );
    not g17191 ( n6051 , n12341 );
    xnor g17192 ( n21948 , n2720 , n21228 );
    and g17193 ( n24012 , n10040 , n9810 );
    xnor g17194 ( n17470 , n24331 , n24798 );
    xnor g17195 ( n21559 , n21317 , n13110 );
    and g17196 ( n14351 , n8976 , n2466 );
    and g17197 ( n15947 , n2607 , n11687 );
    or g17198 ( n21042 , n8694 , n6900 );
    or g17199 ( n4431 , n13293 , n17388 );
    nor g17200 ( n20466 , n22422 , n13521 );
    xnor g17201 ( n16287 , n5527 , n6551 );
    or g17202 ( n15768 , n16873 , n6591 );
    and g17203 ( n17980 , n16699 , n11621 );
    not g17204 ( n27018 , n16058 );
    or g17205 ( n5698 , n15695 , n18 );
    xnor g17206 ( n18711 , n9399 , n14275 );
    or g17207 ( n6618 , n15101 , n3663 );
    and g17208 ( n3288 , n23105 , n19637 );
    or g17209 ( n22098 , n19777 , n17036 );
    not g17210 ( n16961 , n10869 );
    not g17211 ( n22237 , n4509 );
    not g17212 ( n12902 , n7314 );
    or g17213 ( n21987 , n2175 , n4484 );
    nor g17214 ( n24549 , n11707 , n13643 );
    and g17215 ( n436 , n16053 , n1807 );
    not g17216 ( n4170 , n9489 );
    or g17217 ( n14784 , n26082 , n5210 );
    xnor g17218 ( n25946 , n22176 , n23065 );
    and g17219 ( n18072 , n19669 , n23933 );
    and g17220 ( n20168 , n18120 , n11620 );
    xnor g17221 ( n14231 , n10593 , n19701 );
    and g17222 ( n24817 , n2081 , n8693 );
    or g17223 ( n24396 , n2692 , n21394 );
    xnor g17224 ( n4524 , n4897 , n8772 );
    or g17225 ( n2855 , n26132 , n23184 );
    xnor g17226 ( n15859 , n3191 , n25831 );
    or g17227 ( n8686 , n3927 , n10912 );
    or g17228 ( n16384 , n11913 , n14109 );
    or g17229 ( n9074 , n24277 , n20863 );
    or g17230 ( n8257 , n4969 , n18390 );
    xnor g17231 ( n5626 , n10000 , n6790 );
    xnor g17232 ( n22390 , n21101 , n17779 );
    xnor g17233 ( n3233 , n5320 , n19663 );
    nor g17234 ( n23638 , n8745 , n24278 );
    or g17235 ( n20319 , n23833 , n13558 );
    or g17236 ( n3859 , n17438 , n22490 );
    or g17237 ( n24270 , n11440 , n25111 );
    xnor g17238 ( n18282 , n4217 , n25565 );
    or g17239 ( n13321 , n8975 , n26939 );
    xnor g17240 ( n7211 , n2666 , n14739 );
    not g17241 ( n12780 , n2197 );
    or g17242 ( n16644 , n14646 , n22543 );
    xnor g17243 ( n20694 , n25643 , n21753 );
    xnor g17244 ( n17202 , n26527 , n18686 );
    or g17245 ( n10200 , n20998 , n20250 );
    or g17246 ( n26708 , n2570 , n17239 );
    or g17247 ( n11774 , n12020 , n26447 );
    or g17248 ( n26589 , n18646 , n1140 );
    buf g17249 ( n23099 , n7221 );
    xnor g17250 ( n15675 , n1931 , n9980 );
    and g17251 ( n15088 , n24053 , n2727 );
    and g17252 ( n19509 , n25277 , n21860 );
    nor g17253 ( n1609 , n17726 , n14969 );
    not g17254 ( n6743 , n11435 );
    xnor g17255 ( n4731 , n17148 , n9807 );
    and g17256 ( n2676 , n23210 , n18127 );
    and g17257 ( n20634 , n24305 , n2580 );
    nor g17258 ( n14879 , n8255 , n5625 );
    and g17259 ( n23026 , n13537 , n18285 );
    nor g17260 ( n3749 , n24575 , n15232 );
    not g17261 ( n840 , n11580 );
    xnor g17262 ( n3296 , n18283 , n13400 );
    xnor g17263 ( n16558 , n7364 , n2102 );
    and g17264 ( n21457 , n9601 , n26070 );
    and g17265 ( n24756 , n26167 , n18554 );
    xnor g17266 ( n13133 , n24090 , n13110 );
    xnor g17267 ( n23873 , n27040 , n3711 );
    and g17268 ( n19777 , n15411 , n1079 );
    buf g17269 ( n22083 , n3429 );
    and g17270 ( n9342 , n22384 , n26910 );
    xnor g17271 ( n21561 , n23670 , n23775 );
    xnor g17272 ( n17920 , n16427 , n1807 );
    or g17273 ( n6108 , n24766 , n19529 );
    not g17274 ( n14168 , n26572 );
    xnor g17275 ( n15254 , n23504 , n13940 );
    and g17276 ( n2736 , n9752 , n4467 );
    not g17277 ( n4316 , n9936 );
    and g17278 ( n15745 , n8051 , n25573 );
    nor g17279 ( n10265 , n4040 , n655 );
    or g17280 ( n20375 , n11600 , n2423 );
    xnor g17281 ( n24363 , n22764 , n1536 );
    nor g17282 ( n1479 , n15229 , n8050 );
    and g17283 ( n22233 , n6901 , n23385 );
    or g17284 ( n20063 , n22673 , n16265 );
    or g17285 ( n16920 , n2957 , n19285 );
    not g17286 ( n18498 , n9983 );
    not g17287 ( n14963 , n8067 );
    not g17288 ( n14642 , n3770 );
    or g17289 ( n18809 , n26030 , n3752 );
    xnor g17290 ( n15316 , n17411 , n3915 );
    nor g17291 ( n18361 , n14393 , n26239 );
    xnor g17292 ( n4616 , n5380 , n19296 );
    xnor g17293 ( n1792 , n8879 , n6544 );
    xnor g17294 ( n24311 , n3600 , n12836 );
    xnor g17295 ( n12696 , n20534 , n17131 );
    xnor g17296 ( n23978 , n23266 , n7580 );
    xnor g17297 ( n10624 , n12567 , n12279 );
    xnor g17298 ( n20410 , n16400 , n17561 );
    xnor g17299 ( n10092 , n9923 , n767 );
    or g17300 ( n26916 , n26371 , n2418 );
    xnor g17301 ( n2553 , n16652 , n12141 );
    xnor g17302 ( n26832 , n511 , n703 );
    nor g17303 ( n18328 , n11318 , n2615 );
    and g17304 ( n12881 , n13237 , n1066 );
    or g17305 ( n14997 , n21514 , n7947 );
    xnor g17306 ( n10714 , n14361 , n18511 );
    and g17307 ( n16284 , n23828 , n26346 );
    or g17308 ( n16425 , n23311 , n284 );
    xnor g17309 ( n18858 , n169 , n13934 );
    or g17310 ( n23721 , n19358 , n25302 );
    nor g17311 ( n26543 , n2160 , n7335 );
    and g17312 ( n4261 , n24981 , n4091 );
    or g17313 ( n23138 , n26067 , n6643 );
    or g17314 ( n15540 , n20293 , n22006 );
    xnor g17315 ( n17253 , n12821 , n6596 );
    xnor g17316 ( n24080 , n262 , n4489 );
    and g17317 ( n20877 , n15261 , n14630 );
    or g17318 ( n17918 , n24130 , n4721 );
    and g17319 ( n24541 , n8633 , n22810 );
    not g17320 ( n25915 , n5703 );
    not g17321 ( n5313 , n11737 );
    xnor g17322 ( n2540 , n25625 , n6132 );
    nor g17323 ( n18499 , n5330 , n919 );
    xnor g17324 ( n22643 , n8856 , n8305 );
    or g17325 ( n24027 , n525 , n2501 );
    xnor g17326 ( n21623 , n15257 , n604 );
    or g17327 ( n12309 , n15202 , n25805 );
    xnor g17328 ( n389 , n13944 , n23871 );
    xnor g17329 ( n10551 , n26876 , n1662 );
    xnor g17330 ( n4434 , n13177 , n3164 );
    and g17331 ( n9214 , n4237 , n4495 );
    or g17332 ( n17533 , n13410 , n12564 );
    not g17333 ( n26340 , n13936 );
    and g17334 ( n3562 , n4378 , n23929 );
    not g17335 ( n14739 , n15153 );
    or g17336 ( n25153 , n25928 , n17109 );
    nor g17337 ( n12649 , n19297 , n21248 );
    or g17338 ( n19675 , n7974 , n23369 );
    not g17339 ( n8419 , n15931 );
    xnor g17340 ( n14463 , n19065 , n26232 );
    or g17341 ( n9329 , n14162 , n1947 );
    or g17342 ( n25771 , n12183 , n26017 );
    not g17343 ( n26062 , n6790 );
    and g17344 ( n2325 , n7287 , n20154 );
    and g17345 ( n6420 , n5884 , n26468 );
    not g17346 ( n12692 , n12102 );
    xnor g17347 ( n21885 , n1777 , n4812 );
    xnor g17348 ( n16972 , n25830 , n23897 );
    or g17349 ( n10798 , n3252 , n7637 );
    xnor g17350 ( n26866 , n13267 , n16310 );
    xnor g17351 ( n24746 , n9113 , n25643 );
    nor g17352 ( n9855 , n23173 , n15046 );
    xnor g17353 ( n8272 , n2255 , n12558 );
    or g17354 ( n4778 , n7089 , n16793 );
    or g17355 ( n10294 , n4741 , n17818 );
    xnor g17356 ( n21323 , n1532 , n25426 );
    xnor g17357 ( n17880 , n9069 , n22169 );
    or g17358 ( n20155 , n9099 , n19067 );
    or g17359 ( n24527 , n15334 , n11084 );
    or g17360 ( n3958 , n18205 , n18595 );
    and g17361 ( n22469 , n17451 , n22343 );
    xnor g17362 ( n19261 , n20655 , n23170 );
    not g17363 ( n26521 , n12717 );
    or g17364 ( n26868 , n8869 , n1738 );
    and g17365 ( n3128 , n12073 , n14234 );
    and g17366 ( n25445 , n26186 , n19556 );
    not g17367 ( n22186 , n12426 );
    or g17368 ( n2917 , n7237 , n2813 );
    xnor g17369 ( n4834 , n1329 , n12315 );
    not g17370 ( n17467 , n21353 );
    or g17371 ( n19437 , n25171 , n7946 );
    xnor g17372 ( n16589 , n17025 , n14419 );
    xnor g17373 ( n3716 , n13175 , n9567 );
    xnor g17374 ( n20925 , n9548 , n1885 );
    nor g17375 ( n18175 , n3612 , n21274 );
    nor g17376 ( n12551 , n24862 , n24996 );
    not g17377 ( n14218 , n2575 );
    not g17378 ( n21644 , n25370 );
    not g17379 ( n5812 , n19058 );
    xnor g17380 ( n12816 , n3331 , n1023 );
    or g17381 ( n14295 , n333 , n19017 );
    xnor g17382 ( n22821 , n16812 , n1279 );
    not g17383 ( n18255 , n18108 );
    and g17384 ( n26048 , n10109 , n26742 );
    or g17385 ( n24029 , n7155 , n805 );
    or g17386 ( n445 , n24721 , n863 );
    nor g17387 ( n16241 , n524 , n7566 );
    and g17388 ( n25681 , n18825 , n21866 );
    xnor g17389 ( n4095 , n22405 , n24416 );
    and g17390 ( n18817 , n17413 , n12340 );
    or g17391 ( n21054 , n10274 , n18108 );
    or g17392 ( n12006 , n26997 , n23746 );
    and g17393 ( n24178 , n2368 , n9029 );
    and g17394 ( n10543 , n5900 , n23079 );
    and g17395 ( n17330 , n13031 , n9615 );
    and g17396 ( n6047 , n10957 , n12758 );
    or g17397 ( n25746 , n26897 , n5217 );
    not g17398 ( n14967 , n7788 );
    not g17399 ( n14630 , n16902 );
    and g17400 ( n8789 , n6507 , n9524 );
    and g17401 ( n24390 , n1274 , n17469 );
    not g17402 ( n25110 , n17239 );
    or g17403 ( n15494 , n14730 , n13308 );
    or g17404 ( n15420 , n23073 , n8190 );
    not g17405 ( n553 , n2583 );
    not g17406 ( n23061 , n26332 );
    or g17407 ( n18162 , n7297 , n24102 );
    xnor g17408 ( n11837 , n4353 , n17903 );
    xnor g17409 ( n26764 , n18344 , n2965 );
    or g17410 ( n11604 , n13269 , n13022 );
    xnor g17411 ( n3837 , n15743 , n20658 );
    or g17412 ( n21782 , n23914 , n16501 );
    or g17413 ( n4817 , n13810 , n27024 );
    not g17414 ( n5848 , n4578 );
    not g17415 ( n5378 , n14886 );
    nor g17416 ( n9950 , n22683 , n17553 );
    not g17417 ( n27071 , n11429 );
    xnor g17418 ( n5381 , n22619 , n22043 );
    and g17419 ( n24400 , n20372 , n6434 );
    and g17420 ( n20461 , n22146 , n21709 );
    xnor g17421 ( n13050 , n4184 , n4075 );
    xnor g17422 ( n4123 , n10481 , n15802 );
    nor g17423 ( n22487 , n5834 , n3186 );
    xnor g17424 ( n622 , n23114 , n27009 );
    and g17425 ( n8754 , n19444 , n20689 );
    or g17426 ( n20904 , n26038 , n8473 );
    and g17427 ( n16868 , n69 , n8115 );
    or g17428 ( n11780 , n17607 , n16470 );
    not g17429 ( n1904 , n16183 );
    xnor g17430 ( n12553 , n1789 , n5246 );
    xnor g17431 ( n4108 , n7690 , n1428 );
    xnor g17432 ( n13089 , n4860 , n20248 );
    and g17433 ( n4561 , n14337 , n23211 );
    or g17434 ( n15770 , n9282 , n11962 );
    and g17435 ( n290 , n15589 , n25531 );
    xnor g17436 ( n431 , n2603 , n14917 );
    xnor g17437 ( n2889 , n2813 , n1536 );
    not g17438 ( n27007 , n25948 );
    or g17439 ( n17058 , n26877 , n10440 );
    or g17440 ( n24246 , n20857 , n4808 );
    or g17441 ( n20783 , n14940 , n27029 );
    or g17442 ( n21152 , n27139 , n24560 );
    and g17443 ( n18729 , n11889 , n14249 );
    nor g17444 ( n10555 , n10405 , n13960 );
    and g17445 ( n26871 , n7935 , n18608 );
    xnor g17446 ( n10833 , n8291 , n14459 );
    and g17447 ( n437 , n26689 , n12906 );
    xnor g17448 ( n12959 , n12208 , n27074 );
    or g17449 ( n17618 , n24709 , n9997 );
    not g17450 ( n25049 , n23048 );
    or g17451 ( n23001 , n6393 , n25877 );
    xnor g17452 ( n14157 , n5727 , n6137 );
    not g17453 ( n1642 , n3952 );
    and g17454 ( n939 , n11902 , n10827 );
    or g17455 ( n12578 , n20342 , n8526 );
    xnor g17456 ( n24441 , n2818 , n15536 );
    xnor g17457 ( n24368 , n16896 , n9303 );
    and g17458 ( n9529 , n6627 , n4377 );
    not g17459 ( n1657 , n18338 );
    and g17460 ( n13799 , n10429 , n2627 );
    or g17461 ( n11058 , n9797 , n6095 );
    xnor g17462 ( n7267 , n7193 , n16994 );
    and g17463 ( n17197 , n7948 , n19321 );
    and g17464 ( n5023 , n26320 , n6166 );
    xnor g17465 ( n6867 , n7202 , n11772 );
    or g17466 ( n25425 , n21839 , n19282 );
    xnor g17467 ( n8133 , n6079 , n2483 );
    or g17468 ( n19102 , n20243 , n10015 );
    not g17469 ( n11976 , n25607 );
    not g17470 ( n27121 , n3835 );
    or g17471 ( n13342 , n26123 , n7456 );
    or g17472 ( n27086 , n2453 , n1765 );
    not g17473 ( n13671 , n22359 );
    and g17474 ( n5133 , n17539 , n6377 );
    or g17475 ( n16418 , n13564 , n12612 );
    or g17476 ( n7758 , n18908 , n848 );
    and g17477 ( n23596 , n5203 , n26048 );
    or g17478 ( n19290 , n7582 , n15797 );
    xnor g17479 ( n80 , n22272 , n21654 );
    xnor g17480 ( n21267 , n10377 , n19731 );
    and g17481 ( n10368 , n18678 , n12372 );
    or g17482 ( n1774 , n7140 , n8641 );
    not g17483 ( n20978 , n22607 );
    xnor g17484 ( n26489 , n4338 , n25106 );
    or g17485 ( n13707 , n21269 , n5789 );
    or g17486 ( n380 , n640 , n20227 );
    and g17487 ( n16285 , n19872 , n360 );
    or g17488 ( n21178 , n9143 , n16697 );
    xnor g17489 ( n12515 , n23332 , n2199 );
    and g17490 ( n9682 , n12227 , n26558 );
    and g17491 ( n5241 , n12537 , n283 );
    and g17492 ( n20440 , n20066 , n24295 );
    or g17493 ( n24036 , n296 , n16686 );
    or g17494 ( n18702 , n24044 , n8937 );
    xnor g17495 ( n4009 , n18558 , n10411 );
    and g17496 ( n183 , n8243 , n22190 );
    not g17497 ( n18800 , n23545 );
    xnor g17498 ( n21822 , n9071 , n16071 );
    not g17499 ( n3448 , n2439 );
    and g17500 ( n16906 , n481 , n18111 );
    xnor g17501 ( n9261 , n12097 , n14810 );
    and g17502 ( n25781 , n2235 , n22812 );
    xnor g17503 ( n9753 , n1003 , n23233 );
    or g17504 ( n16237 , n14465 , n15204 );
    and g17505 ( n18927 , n26315 , n9982 );
    or g17506 ( n16735 , n22601 , n25727 );
    or g17507 ( n10458 , n24500 , n10208 );
    or g17508 ( n17011 , n14603 , n15053 );
    and g17509 ( n18623 , n23909 , n3812 );
    or g17510 ( n22742 , n22178 , n25783 );
    xnor g17511 ( n763 , n8507 , n15602 );
    and g17512 ( n17155 , n13011 , n3104 );
    or g17513 ( n25969 , n7373 , n13069 );
    xnor g17514 ( n6673 , n2587 , n21859 );
    xnor g17515 ( n23745 , n27169 , n26940 );
    and g17516 ( n2220 , n1366 , n25084 );
    buf g17517 ( n6435 , n25947 );
    nor g17518 ( n15122 , n16400 , n24907 );
    not g17519 ( n3115 , n4743 );
    or g17520 ( n19054 , n10086 , n20176 );
    xnor g17521 ( n139 , n25946 , n9380 );
    not g17522 ( n20326 , n8292 );
    nor g17523 ( n5508 , n20534 , n13146 );
    or g17524 ( n25803 , n2663 , n7911 );
    xnor g17525 ( n24948 , n14555 , n23912 );
    xnor g17526 ( n7931 , n18749 , n4156 );
    or g17527 ( n6609 , n21487 , n10749 );
    or g17528 ( n11126 , n3906 , n16856 );
    and g17529 ( n22830 , n9693 , n10767 );
    xnor g17530 ( n1082 , n24747 , n14737 );
    xnor g17531 ( n14326 , n9169 , n11304 );
    xnor g17532 ( n2313 , n20822 , n14692 );
    or g17533 ( n16990 , n24844 , n16224 );
    xnor g17534 ( n11308 , n1600 , n5482 );
    nor g17535 ( n11518 , n1578 , n20254 );
    xnor g17536 ( n17157 , n2852 , n1432 );
    and g17537 ( n7842 , n26963 , n22828 );
    nor g17538 ( n8900 , n1352 , n10844 );
    nor g17539 ( n14150 , n2156 , n7402 );
    xnor g17540 ( n20803 , n19413 , n2288 );
    or g17541 ( n10856 , n11909 , n12660 );
    nor g17542 ( n22943 , n5938 , n25071 );
    and g17543 ( n974 , n11342 , n4047 );
    and g17544 ( n15941 , n23679 , n1569 );
    or g17545 ( n26531 , n13227 , n21503 );
    and g17546 ( n15756 , n3740 , n2545 );
    not g17547 ( n27115 , n20618 );
    xnor g17548 ( n564 , n16166 , n14705 );
    nor g17549 ( n24682 , n13 , n23792 );
    nor g17550 ( n11523 , n23428 , n5834 );
    xnor g17551 ( n11482 , n17646 , n24393 );
    xnor g17552 ( n8604 , n21570 , n9598 );
    nor g17553 ( n7661 , n23819 , n22861 );
    nor g17554 ( n11875 , n14904 , n11575 );
    nor g17555 ( n9757 , n4473 , n3798 );
    xnor g17556 ( n24626 , n14043 , n2076 );
    and g17557 ( n7040 , n17122 , n23383 );
    not g17558 ( n13507 , n5038 );
    xnor g17559 ( n6555 , n16755 , n367 );
    not g17560 ( n4087 , n23333 );
    xnor g17561 ( n9106 , n18537 , n5211 );
    and g17562 ( n7043 , n6164 , n25942 );
    and g17563 ( n438 , n21517 , n16972 );
    xnor g17564 ( n16424 , n2854 , n2660 );
    and g17565 ( n20825 , n21582 , n24553 );
    and g17566 ( n13813 , n23472 , n20736 );
    or g17567 ( n18848 , n852 , n13476 );
    not g17568 ( n4315 , n19116 );
    or g17569 ( n9905 , n2219 , n2813 );
    not g17570 ( n24024 , n5737 );
    and g17571 ( n24099 , n14626 , n20843 );
    and g17572 ( n14613 , n21287 , n23705 );
    xnor g17573 ( n9104 , n24653 , n26602 );
    or g17574 ( n5293 , n21869 , n21999 );
    or g17575 ( n23723 , n2369 , n18899 );
    xnor g17576 ( n21396 , n13192 , n18050 );
    or g17577 ( n21921 , n14958 , n5800 );
    xnor g17578 ( n4785 , n11934 , n2094 );
    or g17579 ( n25968 , n6222 , n19378 );
    not g17580 ( n22351 , n8194 );
    xnor g17581 ( n18503 , n1364 , n8256 );
    or g17582 ( n11536 , n12147 , n9485 );
    xnor g17583 ( n13533 , n2225 , n11181 );
    not g17584 ( n19170 , n2923 );
    and g17585 ( n2297 , n16833 , n21910 );
    and g17586 ( n4990 , n6236 , n13160 );
    nor g17587 ( n17753 , n16197 , n24936 );
    xnor g17588 ( n16291 , n6143 , n1689 );
    xnor g17589 ( n4071 , n11247 , n19919 );
    nor g17590 ( n20128 , n21378 , n14584 );
    or g17591 ( n23052 , n3900 , n16202 );
    or g17592 ( n6205 , n26087 , n7243 );
    and g17593 ( n19326 , n27205 , n6858 );
    xnor g17594 ( n17629 , n6191 , n4935 );
    nor g17595 ( n13950 , n10017 , n20349 );
    or g17596 ( n2683 , n24435 , n21179 );
    and g17597 ( n1598 , n21251 , n10830 );
    xnor g17598 ( n10065 , n9259 , n6456 );
    xnor g17599 ( n4529 , n27023 , n10818 );
    or g17600 ( n25860 , n21845 , n8247 );
    not g17601 ( n2896 , n16911 );
    not g17602 ( n11000 , n20925 );
    or g17603 ( n5724 , n25139 , n16696 );
    not g17604 ( n16477 , n14723 );
    or g17605 ( n2707 , n9509 , n6566 );
    xnor g17606 ( n643 , n8300 , n12761 );
    xnor g17607 ( n7402 , n14334 , n23393 );
    xnor g17608 ( n14314 , n2391 , n19647 );
    or g17609 ( n13768 , n23111 , n18536 );
    or g17610 ( n13423 , n4522 , n1579 );
    not g17611 ( n22517 , n20621 );
    xnor g17612 ( n1313 , n21828 , n18227 );
    or g17613 ( n11090 , n8856 , n19768 );
    and g17614 ( n989 , n25931 , n1510 );
    xnor g17615 ( n1391 , n13734 , n18548 );
    or g17616 ( n25587 , n22622 , n16535 );
    xnor g17617 ( n11168 , n1639 , n23842 );
    xnor g17618 ( n27168 , n26935 , n307 );
    or g17619 ( n26750 , n11257 , n24121 );
    xnor g17620 ( n10114 , n18422 , n26816 );
    or g17621 ( n16505 , n8711 , n17318 );
    not g17622 ( n8241 , n13578 );
    xnor g17623 ( n1353 , n20138 , n10372 );
    or g17624 ( n13859 , n2279 , n21232 );
    nor g17625 ( n1841 , n11738 , n24024 );
    and g17626 ( n25837 , n18227 , n21828 );
    not g17627 ( n6139 , n16519 );
    or g17628 ( n25399 , n12051 , n13813 );
    nor g17629 ( n14895 , n26056 , n27151 );
    not g17630 ( n20109 , n21916 );
    xnor g17631 ( n26018 , n12048 , n8210 );
    and g17632 ( n14932 , n14618 , n10370 );
    xnor g17633 ( n12358 , n10001 , n21222 );
    xnor g17634 ( n25057 , n10400 , n15814 );
    and g17635 ( n13091 , n1921 , n20309 );
    nor g17636 ( n5353 , n403 , n509 );
    or g17637 ( n695 , n25579 , n13592 );
    and g17638 ( n22629 , n20257 , n26517 );
    not g17639 ( n3877 , n17902 );
    not g17640 ( n12171 , n4356 );
    nor g17641 ( n8552 , n19270 , n19702 );
    not g17642 ( n14431 , n26443 );
    and g17643 ( n1123 , n23028 , n6539 );
    not g17644 ( n14695 , n4409 );
    and g17645 ( n22088 , n14530 , n19837 );
    or g17646 ( n23993 , n5811 , n13437 );
    xnor g17647 ( n13179 , n13625 , n10989 );
    xnor g17648 ( n496 , n12439 , n15999 );
    not g17649 ( n18676 , n2899 );
    and g17650 ( n22202 , n22435 , n21479 );
    not g17651 ( n16464 , n15636 );
    and g17652 ( n3548 , n14283 , n12782 );
    or g17653 ( n21361 , n26299 , n22535 );
    or g17654 ( n98 , n2422 , n1562 );
    nor g17655 ( n17425 , n16117 , n8891 );
    or g17656 ( n25657 , n22209 , n9896 );
    xnor g17657 ( n23264 , n26978 , n1961 );
    or g17658 ( n26213 , n23660 , n3671 );
    xnor g17659 ( n16954 , n1397 , n7783 );
    or g17660 ( n22657 , n1275 , n7289 );
    not g17661 ( n23436 , n6369 );
    and g17662 ( n908 , n3388 , n18009 );
    nor g17663 ( n7726 , n2247 , n19715 );
    xnor g17664 ( n17228 , n22247 , n19502 );
    or g17665 ( n17990 , n26904 , n17266 );
    nor g17666 ( n8743 , n19531 , n1999 );
    xnor g17667 ( n18758 , n5000 , n18282 );
    xnor g17668 ( n25244 , n20116 , n8245 );
    not g17669 ( n20777 , n19399 );
    xnor g17670 ( n23690 , n23813 , n21968 );
    or g17671 ( n25932 , n16077 , n21210 );
    xnor g17672 ( n18608 , n899 , n3564 );
    xnor g17673 ( n7426 , n1021 , n21604 );
    or g17674 ( n10402 , n14078 , n4583 );
    and g17675 ( n22677 , n26730 , n6823 );
    xnor g17676 ( n2845 , n13206 , n7421 );
    or g17677 ( n7814 , n16053 , n1807 );
    xnor g17678 ( n16847 , n14680 , n16439 );
    and g17679 ( n25907 , n8588 , n23404 );
    and g17680 ( n13811 , n2973 , n19397 );
    xnor g17681 ( n12041 , n5617 , n20734 );
    xnor g17682 ( n4019 , n14254 , n11502 );
    or g17683 ( n21807 , n1009 , n4999 );
    and g17684 ( n5562 , n5401 , n3578 );
    and g17685 ( n18827 , n26578 , n3999 );
    not g17686 ( n24018 , n16482 );
    not g17687 ( n9945 , n3465 );
    xnor g17688 ( n13959 , n11356 , n12587 );
    and g17689 ( n1508 , n15429 , n23723 );
    or g17690 ( n19448 , n4298 , n16290 );
    xnor g17691 ( n26479 , n20231 , n20201 );
    not g17692 ( n10773 , n11455 );
    or g17693 ( n26418 , n22089 , n20139 );
    not g17694 ( n5483 , n16026 );
    or g17695 ( n13716 , n14617 , n9786 );
    xnor g17696 ( n4961 , n2331 , n22879 );
    nor g17697 ( n15629 , n18290 , n9455 );
    xnor g17698 ( n2282 , n25291 , n20558 );
    xnor g17699 ( n3300 , n2939 , n16960 );
    or g17700 ( n4206 , n13910 , n20461 );
    xnor g17701 ( n16915 , n25126 , n21226 );
    nor g17702 ( n10100 , n8694 , n20039 );
    and g17703 ( n19563 , n11760 , n3816 );
    xnor g17704 ( n19020 , n18345 , n25168 );
    and g17705 ( n18738 , n13596 , n10649 );
    and g17706 ( n15557 , n1063 , n15394 );
    not g17707 ( n14140 , n14692 );
    and g17708 ( n22916 , n11635 , n13321 );
    xnor g17709 ( n10234 , n25144 , n11121 );
    or g17710 ( n13431 , n21377 , n13299 );
    or g17711 ( n6225 , n5037 , n17955 );
    not g17712 ( n21322 , n18563 );
    and g17713 ( n24675 , n10180 , n2865 );
    not g17714 ( n9098 , n26972 );
    xnor g17715 ( n3983 , n14824 , n21315 );
    xnor g17716 ( n21155 , n14067 , n7468 );
    xnor g17717 ( n13384 , n20240 , n2845 );
    or g17718 ( n355 , n18477 , n2060 );
    or g17719 ( n23082 , n9733 , n13216 );
    nor g17720 ( n24416 , n9223 , n4055 );
    or g17721 ( n17246 , n14950 , n260 );
    not g17722 ( n20615 , n17188 );
    or g17723 ( n23023 , n9934 , n20290 );
    not g17724 ( n18495 , n11537 );
    or g17725 ( n26950 , n20062 , n6562 );
    or g17726 ( n15107 , n3179 , n12658 );
    xnor g17727 ( n13220 , n3103 , n22471 );
    or g17728 ( n27026 , n11390 , n7970 );
    and g17729 ( n2741 , n22674 , n6378 );
    xnor g17730 ( n21573 , n21352 , n19057 );
    xnor g17731 ( n14533 , n18539 , n16818 );
    and g17732 ( n10776 , n17534 , n19273 );
    xnor g17733 ( n26851 , n9676 , n26771 );
    xnor g17734 ( n8258 , n6403 , n4722 );
    buf g17735 ( n1765 , n5607 );
    nor g17736 ( n7835 , n23005 , n11531 );
    nor g17737 ( n9020 , n14718 , n8820 );
    xnor g17738 ( n16924 , n15591 , n10725 );
    not g17739 ( n26064 , n16247 );
    not g17740 ( n16309 , n2436 );
    xnor g17741 ( n12075 , n12333 , n18863 );
    not g17742 ( n26186 , n7652 );
    or g17743 ( n2393 , n15667 , n1983 );
    or g17744 ( n3941 , n21502 , n5674 );
    nor g17745 ( n15530 , n22491 , n22600 );
    and g17746 ( n5526 , n21802 , n25294 );
    or g17747 ( n11021 , n11566 , n10973 );
    or g17748 ( n7954 , n19770 , n12022 );
    xnor g17749 ( n4446 , n8407 , n13491 );
    and g17750 ( n9904 , n11903 , n14872 );
    or g17751 ( n8446 , n25616 , n23246 );
    xnor g17752 ( n20770 , n5070 , n8734 );
    and g17753 ( n26441 , n2012 , n6960 );
    xnor g17754 ( n11493 , n6115 , n2352 );
    xnor g17755 ( n19623 , n17376 , n7295 );
    or g17756 ( n2183 , n21410 , n5862 );
    xnor g17757 ( n20539 , n5579 , n26054 );
    or g17758 ( n7014 , n19173 , n8483 );
    and g17759 ( n9319 , n24094 , n7922 );
    not g17760 ( n18058 , n15053 );
    or g17761 ( n25313 , n22176 , n19298 );
    not g17762 ( n13159 , n2680 );
    xnor g17763 ( n8085 , n27002 , n18502 );
    or g17764 ( n10656 , n10556 , n13846 );
    xnor g17765 ( n18934 , n23349 , n16759 );
    not g17766 ( n14254 , n21073 );
    or g17767 ( n20066 , n8945 , n16582 );
    and g17768 ( n17646 , n22718 , n22957 );
    and g17769 ( n17767 , n22719 , n24589 );
    and g17770 ( n19257 , n14295 , n2720 );
    or g17771 ( n25601 , n13026 , n13369 );
    xnor g17772 ( n703 , n8657 , n10593 );
    xnor g17773 ( n737 , n13339 , n4623 );
    not g17774 ( n18559 , n26541 );
    not g17775 ( n26212 , n22350 );
    not g17776 ( n13459 , n20036 );
    or g17777 ( n4311 , n12960 , n1344 );
    xnor g17778 ( n19571 , n5374 , n18649 );
    xnor g17779 ( n17237 , n23874 , n23923 );
    xnor g17780 ( n13669 , n24402 , n1230 );
    not g17781 ( n11086 , n21768 );
    xnor g17782 ( n7828 , n12495 , n11479 );
    xnor g17783 ( n5625 , n16976 , n2880 );
    and g17784 ( n25138 , n4887 , n5045 );
    xnor g17785 ( n457 , n23132 , n19204 );
    xnor g17786 ( n3611 , n21998 , n3945 );
    and g17787 ( n17001 , n355 , n27077 );
    xnor g17788 ( n9371 , n16687 , n15213 );
    and g17789 ( n7022 , n21811 , n2571 );
    nor g17790 ( n25085 , n14254 , n6964 );
    and g17791 ( n4866 , n99 , n1399 );
    and g17792 ( n23810 , n26593 , n17374 );
    xnor g17793 ( n20252 , n26705 , n22061 );
    or g17794 ( n18132 , n18774 , n22784 );
    nor g17795 ( n24611 , n12454 , n5714 );
    xnor g17796 ( n6967 , n5492 , n19947 );
    or g17797 ( n26259 , n23843 , n19486 );
    or g17798 ( n213 , n2709 , n1093 );
    and g17799 ( n25048 , n9248 , n14755 );
    xnor g17800 ( n8164 , n15704 , n21308 );
    xnor g17801 ( n15850 , n23533 , n9636 );
    not g17802 ( n10882 , n21324 );
    not g17803 ( n306 , n11201 );
    not g17804 ( n14532 , n24042 );
    and g17805 ( n24293 , n21987 , n8882 );
    nor g17806 ( n5480 , n17906 , n24628 );
    and g17807 ( n6123 , n15354 , n9721 );
    or g17808 ( n3756 , n13172 , n23892 );
    or g17809 ( n14817 , n23269 , n15848 );
    and g17810 ( n17340 , n10376 , n3615 );
    xnor g17811 ( n24935 , n22528 , n20421 );
    xnor g17812 ( n8635 , n7508 , n12438 );
    not g17813 ( n17590 , n4095 );
    not g17814 ( n6486 , n6555 );
    xnor g17815 ( n6669 , n2910 , n19681 );
    and g17816 ( n19419 , n2506 , n4465 );
    or g17817 ( n641 , n21213 , n15392 );
    or g17818 ( n22019 , n15891 , n9319 );
    not g17819 ( n11069 , n20385 );
    and g17820 ( n3994 , n16712 , n3706 );
    or g17821 ( n21954 , n8675 , n18559 );
    or g17822 ( n22572 , n14415 , n26717 );
    not g17823 ( n17617 , n25018 );
    or g17824 ( n21730 , n5338 , n16752 );
    xnor g17825 ( n5614 , n19312 , n24933 );
    xnor g17826 ( n9324 , n26170 , n19884 );
    or g17827 ( n14034 , n19978 , n21111 );
    or g17828 ( n5382 , n22055 , n9184 );
    xnor g17829 ( n1385 , n21949 , n24872 );
    or g17830 ( n12777 , n8636 , n24591 );
    xnor g17831 ( n6911 , n10042 , n2686 );
    not g17832 ( n13027 , n22321 );
    and g17833 ( n22712 , n14060 , n16621 );
    or g17834 ( n4281 , n23448 , n7325 );
    and g17835 ( n6230 , n2080 , n13919 );
    or g17836 ( n18131 , n10720 , n7285 );
    xnor g17837 ( n25719 , n20813 , n10423 );
    xnor g17838 ( n25128 , n5090 , n21674 );
    nor g17839 ( n18340 , n21929 , n485 );
    xnor g17840 ( n50 , n16122 , n9022 );
    and g17841 ( n10556 , n22585 , n23226 );
    xnor g17842 ( n13135 , n14630 , n7270 );
    or g17843 ( n8693 , n5418 , n23847 );
    and g17844 ( n1083 , n20090 , n8811 );
    xnor g17845 ( n3614 , n3205 , n24708 );
    not g17846 ( n15618 , n25688 );
    xnor g17847 ( n21505 , n8959 , n3441 );
    xnor g17848 ( n16280 , n11504 , n752 );
    or g17849 ( n18041 , n18690 , n7685 );
    not g17850 ( n23168 , n11579 );
    and g17851 ( n19915 , n9513 , n23417 );
    xnor g17852 ( n10420 , n4177 , n6545 );
    xnor g17853 ( n4560 , n12616 , n22879 );
    nor g17854 ( n3305 , n2113 , n14345 );
    nor g17855 ( n22994 , n25240 , n6510 );
    or g17856 ( n22056 , n9554 , n9509 );
    nor g17857 ( n13845 , n24600 , n3641 );
    xnor g17858 ( n27164 , n23475 , n13419 );
    nor g17859 ( n23015 , n19940 , n10407 );
    or g17860 ( n23158 , n23750 , n14963 );
    xnor g17861 ( n8896 , n23216 , n1324 );
    nor g17862 ( n1164 , n7360 , n16482 );
    xnor g17863 ( n8681 , n14680 , n25240 );
    and g17864 ( n25440 , n14040 , n8477 );
    or g17865 ( n3732 , n6511 , n13738 );
    xnor g17866 ( n10783 , n15892 , n8448 );
    or g17867 ( n16761 , n23750 , n7678 );
    or g17868 ( n7651 , n52 , n23656 );
    and g17869 ( n9741 , n21434 , n14301 );
    and g17870 ( n23508 , n26474 , n24534 );
    xnor g17871 ( n9042 , n26633 , n20048 );
    xnor g17872 ( n4349 , n8713 , n21300 );
    xnor g17873 ( n12883 , n17600 , n6859 );
    xnor g17874 ( n13834 , n3414 , n20923 );
    xnor g17875 ( n4984 , n4446 , n24551 );
    xnor g17876 ( n11797 , n5055 , n14767 );
    and g17877 ( n25479 , n5282 , n13720 );
    nor g17878 ( n10225 , n2062 , n23191 );
    and g17879 ( n25229 , n2015 , n309 );
    or g17880 ( n24668 , n14897 , n6014 );
    nor g17881 ( n10205 , n11302 , n2146 );
    or g17882 ( n2654 , n23648 , n3646 );
    and g17883 ( n9414 , n12943 , n797 );
    not g17884 ( n6293 , n23882 );
    and g17885 ( n19700 , n25769 , n15776 );
    xnor g17886 ( n186 , n14965 , n25465 );
    xnor g17887 ( n25684 , n13224 , n15041 );
    xnor g17888 ( n11398 , n15287 , n15140 );
    or g17889 ( n6496 , n3403 , n3271 );
    xnor g17890 ( n357 , n23896 , n15909 );
    and g17891 ( n8524 , n10439 , n12139 );
    xnor g17892 ( n26250 , n12331 , n23300 );
    not g17893 ( n17858 , n8724 );
    or g17894 ( n22063 , n20730 , n14453 );
    nor g17895 ( n19304 , n602 , n19971 );
    xnor g17896 ( n14380 , n1489 , n19517 );
    or g17897 ( n10502 , n6830 , n19773 );
    or g17898 ( n25301 , n16009 , n12910 );
    and g17899 ( n22521 , n11457 , n10266 );
    xnor g17900 ( n2923 , n14793 , n25375 );
    and g17901 ( n2691 , n10752 , n21326 );
    and g17902 ( n23661 , n1317 , n5202 );
    xnor g17903 ( n26306 , n13241 , n13998 );
    or g17904 ( n9994 , n13576 , n25165 );
    or g17905 ( n36 , n19472 , n8997 );
    xnor g17906 ( n2197 , n15283 , n8020 );
    xnor g17907 ( n7516 , n4924 , n25230 );
    xor g17908 ( n1177 , n17088 , n18472 );
    xnor g17909 ( n14983 , n21620 , n9404 );
    xnor g17910 ( n8485 , n4289 , n8178 );
    or g17911 ( n23021 , n25674 , n16029 );
    xnor g17912 ( n13436 , n13606 , n7091 );
    xnor g17913 ( n26348 , n11356 , n2999 );
    xnor g17914 ( n4891 , n6906 , n26709 );
    or g17915 ( n13779 , n13704 , n5240 );
    xnor g17916 ( n34 , n5796 , n25856 );
    or g17917 ( n22143 , n9080 , n3609 );
    or g17918 ( n26861 , n17531 , n8592 );
    nor g17919 ( n17957 , n19978 , n24239 );
    or g17920 ( n19395 , n19742 , n4867 );
    or g17921 ( n6856 , n15529 , n11985 );
    or g17922 ( n22663 , n2726 , n23179 );
    or g17923 ( n8907 , n10946 , n18881 );
    or g17924 ( n23777 , n18750 , n11609 );
    nor g17925 ( n20837 , n22736 , n17390 );
    or g17926 ( n5596 , n22919 , n19074 );
    or g17927 ( n12997 , n4130 , n21740 );
    xnor g17928 ( n24953 , n9557 , n21832 );
    and g17929 ( n18778 , n344 , n26205 );
    xnor g17930 ( n7268 , n1567 , n6412 );
    xnor g17931 ( n15376 , n13784 , n17959 );
    nor g17932 ( n4533 , n840 , n7604 );
    or g17933 ( n5175 , n3521 , n8323 );
    nor g17934 ( n2299 , n7827 , n9505 );
    xor g17935 ( n3772 , n10218 , n22612 );
    and g17936 ( n6969 , n17697 , n11599 );
    nor g17937 ( n18853 , n3366 , n23456 );
    xnor g17938 ( n14734 , n7911 , n25983 );
    or g17939 ( n21614 , n4902 , n928 );
    or g17940 ( n16999 , n5611 , n9671 );
    xnor g17941 ( n9854 , n8785 , n14841 );
    not g17942 ( n4353 , n15154 );
    nor g17943 ( n2103 , n21209 , n25001 );
    not g17944 ( n11846 , n4864 );
    xnor g17945 ( n3893 , n26046 , n21246 );
    or g17946 ( n7034 , n1429 , n25555 );
    not g17947 ( n8472 , n4917 );
    xnor g17948 ( n21448 , n19383 , n10422 );
    not g17949 ( n6122 , n152 );
    xnor g17950 ( n20054 , n4588 , n27134 );
    and g17951 ( n14693 , n21687 , n6458 );
    not g17952 ( n7511 , n130 );
    or g17953 ( n19242 , n20751 , n19845 );
    not g17954 ( n8224 , n1138 );
    nor g17955 ( n18990 , n24996 , n24488 );
    xnor g17956 ( n5072 , n15714 , n22364 );
    not g17957 ( n926 , n12436 );
    xnor g17958 ( n18751 , n22356 , n4958 );
    and g17959 ( n22287 , n3914 , n1717 );
    or g17960 ( n4827 , n4974 , n26985 );
    xnor g17961 ( n4459 , n9156 , n9841 );
    xnor g17962 ( n26353 , n6698 , n1086 );
    or g17963 ( n16624 , n8422 , n7100 );
    xnor g17964 ( n25730 , n21125 , n7377 );
    xnor g17965 ( n25223 , n7097 , n9469 );
    or g17966 ( n24300 , n12923 , n23820 );
    or g17967 ( n3372 , n13729 , n21674 );
    and g17968 ( n19179 , n19362 , n15690 );
    or g17969 ( n20738 , n17799 , n13917 );
    or g17970 ( n187 , n24627 , n6374 );
    not g17971 ( n21764 , n9124 );
    or g17972 ( n19945 , n11980 , n9971 );
    or g17973 ( n3088 , n21676 , n5135 );
    or g17974 ( n23521 , n8835 , n2235 );
    xnor g17975 ( n25419 , n8892 , n2313 );
    and g17976 ( n23407 , n9013 , n993 );
    xnor g17977 ( n23602 , n11718 , n13834 );
    and g17978 ( n8537 , n8032 , n1343 );
    or g17979 ( n3032 , n12437 , n17465 );
    and g17980 ( n7911 , n16160 , n7113 );
    or g17981 ( n15436 , n16818 , n13133 );
    xnor g17982 ( n24198 , n7566 , n19357 );
    and g17983 ( n9617 , n3346 , n19311 );
    or g17984 ( n1800 , n734 , n3321 );
    xnor g17985 ( n904 , n13482 , n10686 );
    not g17986 ( n20944 , n19190 );
    and g17987 ( n6907 , n5558 , n7481 );
    xnor g17988 ( n1822 , n14826 , n13549 );
    xnor g17989 ( n15210 , n8948 , n3470 );
    or g17990 ( n24641 , n16842 , n23571 );
    and g17991 ( n1790 , n9490 , n23693 );
    and g17992 ( n13921 , n22892 , n5165 );
    xnor g17993 ( n18611 , n5517 , n21981 );
    or g17994 ( n5290 , n5386 , n24326 );
    nor g17995 ( n9141 , n14818 , n10158 );
    or g17996 ( n16164 , n9098 , n6908 );
    nor g17997 ( n22178 , n21867 , n7948 );
    nor g17998 ( n18294 , n25764 , n17447 );
    xnor g17999 ( n25840 , n16344 , n26454 );
    not g18000 ( n8361 , n19539 );
    and g18001 ( n14689 , n18506 , n3994 );
    xnor g18002 ( n25636 , n21162 , n8614 );
    not g18003 ( n26536 , n25748 );
    xnor g18004 ( n20171 , n363 , n21732 );
    or g18005 ( n15356 , n4140 , n24882 );
    xnor g18006 ( n3271 , n12111 , n12668 );
    or g18007 ( n24467 , n9628 , n21640 );
    xnor g18008 ( n16149 , n3909 , n19081 );
    or g18009 ( n15344 , n18995 , n3614 );
    not g18010 ( n6685 , n13300 );
    or g18011 ( n2392 , n14992 , n22764 );
    and g18012 ( n19795 , n9977 , n14956 );
    nor g18013 ( n14402 , n6321 , n20349 );
    nor g18014 ( n16720 , n22558 , n8155 );
    and g18015 ( n10742 , n14978 , n26455 );
    xnor g18016 ( n9954 , n20127 , n13650 );
    buf g18017 ( n905 , n15723 );
    or g18018 ( n17964 , n5316 , n7152 );
    or g18019 ( n19043 , n23187 , n20833 );
    xnor g18020 ( n23954 , n7909 , n18636 );
    or g18021 ( n25734 , n14374 , n8652 );
    or g18022 ( n4196 , n9134 , n19412 );
    xnor g18023 ( n12012 , n27144 , n14692 );
    nor g18024 ( n22183 , n17250 , n4409 );
    or g18025 ( n3912 , n5039 , n8380 );
    xnor g18026 ( n19176 , n13415 , n6237 );
    xnor g18027 ( n12756 , n17128 , n21441 );
    or g18028 ( n25305 , n22225 , n21620 );
    buf g18029 ( n3981 , n1913 );
    xnor g18030 ( n22974 , n20929 , n24620 );
    or g18031 ( n25483 , n13865 , n4504 );
    xnor g18032 ( n20790 , n17360 , n14684 );
    or g18033 ( n995 , n19898 , n17645 );
    and g18034 ( n27186 , n20826 , n14532 );
    xnor g18035 ( n18163 , n17224 , n8526 );
    xnor g18036 ( n13968 , n13341 , n11251 );
    not g18037 ( n12714 , n19803 );
    xnor g18038 ( n23434 , n719 , n25561 );
    nor g18039 ( n22834 , n10571 , n9431 );
    or g18040 ( n18136 , n25715 , n8343 );
    xnor g18041 ( n24758 , n10589 , n13698 );
    not g18042 ( n12709 , n3223 );
    or g18043 ( n780 , n10311 , n14713 );
    and g18044 ( n21130 , n7730 , n15043 );
    and g18045 ( n24037 , n11759 , n26836 );
    xnor g18046 ( n19694 , n23923 , n25119 );
    and g18047 ( n2224 , n1901 , n12432 );
    not g18048 ( n3314 , n26104 );
    xnor g18049 ( n2124 , n14078 , n18891 );
    xnor g18050 ( n27132 , n23731 , n5842 );
    xnor g18051 ( n3903 , n13132 , n17253 );
    not g18052 ( n9703 , n3729 );
    xnor g18053 ( n12029 , n3447 , n10669 );
    or g18054 ( n17966 , n8739 , n16693 );
    and g18055 ( n26415 , n14972 , n5354 );
    and g18056 ( n1080 , n26692 , n11015 );
    nor g18057 ( n10085 , n13518 , n5743 );
    xnor g18058 ( n13456 , n9173 , n23148 );
    not g18059 ( n21777 , n8107 );
    or g18060 ( n10972 , n307 , n16046 );
    or g18061 ( n20046 , n20965 , n8207 );
    or g18062 ( n471 , n24285 , n6180 );
    not g18063 ( n25270 , n14633 );
    nor g18064 ( n23737 , n20104 , n15616 );
    not g18065 ( n25000 , n27164 );
    xnor g18066 ( n16108 , n23216 , n15093 );
    xnor g18067 ( n15011 , n14368 , n16305 );
    or g18068 ( n247 , n22196 , n20900 );
    xnor g18069 ( n18935 , n25494 , n6659 );
    or g18070 ( n6018 , n15427 , n10168 );
    and g18071 ( n15528 , n1013 , n25154 );
    nor g18072 ( n22432 , n16476 , n15008 );
    or g18073 ( n9571 , n23502 , n24567 );
    and g18074 ( n18443 , n25857 , n14912 );
    xnor g18075 ( n15232 , n23476 , n19783 );
    xnor g18076 ( n23148 , n16559 , n6872 );
    xnor g18077 ( n13198 , n10708 , n20521 );
    nor g18078 ( n14909 , n17069 , n16608 );
    nor g18079 ( n20114 , n617 , n7798 );
    or g18080 ( n22357 , n18853 , n3175 );
    nor g18081 ( n1677 , n26064 , n10930 );
    and g18082 ( n10735 , n13690 , n22927 );
    and g18083 ( n24856 , n10112 , n21849 );
    nor g18084 ( n3766 , n268 , n19265 );
    not g18085 ( n14926 , n6765 );
    xnor g18086 ( n12430 , n2448 , n13296 );
    and g18087 ( n1297 , n17346 , n13606 );
    or g18088 ( n16341 , n26093 , n20138 );
    xnor g18089 ( n10777 , n22788 , n8427 );
    and g18090 ( n1221 , n5271 , n11478 );
    xnor g18091 ( n12812 , n17686 , n4553 );
    or g18092 ( n26579 , n26966 , n18063 );
    not g18093 ( n21774 , n22552 );
    and g18094 ( n6498 , n18870 , n12867 );
    and g18095 ( n3610 , n12343 , n16357 );
    and g18096 ( n8961 , n7014 , n23557 );
    xnor g18097 ( n13568 , n11382 , n16637 );
    xnor g18098 ( n18865 , n6167 , n13581 );
    xnor g18099 ( n22325 , n24362 , n17625 );
    xnor g18100 ( n14857 , n17600 , n16054 );
    nor g18101 ( n16061 , n26553 , n23775 );
    xnor g18102 ( n24419 , n25877 , n26443 );
    nor g18103 ( n26767 , n274 , n2618 );
    xnor g18104 ( n16207 , n14907 , n25238 );
    or g18105 ( n8915 , n24019 , n24238 );
    and g18106 ( n5114 , n16661 , n25859 );
    or g18107 ( n14915 , n15249 , n19550 );
    and g18108 ( n13025 , n10594 , n9355 );
    not g18109 ( n23443 , n532 );
    xnor g18110 ( n1444 , n10529 , n22498 );
    xnor g18111 ( n7867 , n2849 , n20641 );
    or g18112 ( n13688 , n22809 , n584 );
    and g18113 ( n1910 , n18803 , n5327 );
    xnor g18114 ( n3400 , n12877 , n6094 );
    nor g18115 ( n25775 , n11554 , n20734 );
    nor g18116 ( n1154 , n21997 , n26962 );
    or g18117 ( n1306 , n1804 , n15390 );
    not g18118 ( n9366 , n24896 );
    xnor g18119 ( n26857 , n1445 , n18260 );
    nor g18120 ( n18666 , n26452 , n3783 );
    nor g18121 ( n3666 , n18934 , n9820 );
    xnor g18122 ( n757 , n10824 , n13761 );
    or g18123 ( n18053 , n20530 , n4822 );
    or g18124 ( n26841 , n21613 , n16807 );
    or g18125 ( n25059 , n24638 , n26645 );
    xnor g18126 ( n21976 , n11333 , n11648 );
    or g18127 ( n5563 , n16059 , n12737 );
    not g18128 ( n3053 , n9972 );
    or g18129 ( n19548 , n23590 , n20184 );
    not g18130 ( n867 , n25365 );
    xnor g18131 ( n13906 , n26955 , n3478 );
    not g18132 ( n3779 , n4404 );
    nor g18133 ( n26980 , n252 , n20316 );
    and g18134 ( n13663 , n11492 , n1347 );
    and g18135 ( n19748 , n8108 , n24931 );
    xnor g18136 ( n25016 , n10514 , n4514 );
    or g18137 ( n15668 , n10023 , n7216 );
    not g18138 ( n22773 , n23268 );
    xnor g18139 ( n1277 , n16117 , n9832 );
    not g18140 ( n6632 , n10022 );
    and g18141 ( n23880 , n8227 , n11947 );
    xnor g18142 ( n22026 , n3382 , n18363 );
    not g18143 ( n14634 , n11653 );
    xnor g18144 ( n2265 , n19222 , n1786 );
    xnor g18145 ( n4652 , n15912 , n19896 );
    or g18146 ( n12947 , n6549 , n13108 );
    or g18147 ( n19490 , n2404 , n9931 );
    nor g18148 ( n4412 , n22095 , n713 );
    not g18149 ( n23096 , n7505 );
    and g18150 ( n27161 , n10118 , n2544 );
    xnor g18151 ( n12445 , n9137 , n5513 );
    or g18152 ( n5099 , n18294 , n26383 );
    and g18153 ( n12645 , n270 , n5198 );
    or g18154 ( n1220 , n19074 , n6504 );
    xnor g18155 ( n9266 , n178 , n2042 );
    and g18156 ( n10597 , n22091 , n18861 );
    or g18157 ( n13687 , n18370 , n11289 );
    and g18158 ( n17085 , n22529 , n179 );
    or g18159 ( n26480 , n1437 , n17784 );
    or g18160 ( n19165 , n1742 , n1798 );
    and g18161 ( n14678 , n4511 , n19573 );
    not g18162 ( n23234 , n11486 );
    xnor g18163 ( n2561 , n15044 , n6730 );
    xnor g18164 ( n21062 , n18923 , n22416 );
    and g18165 ( n19487 , n16044 , n10772 );
    or g18166 ( n24865 , n23211 , n14569 );
    and g18167 ( n24078 , n20293 , n22006 );
    xnor g18168 ( n21198 , n3480 , n3136 );
    xnor g18169 ( n2316 , n26089 , n389 );
    and g18170 ( n16893 , n4119 , n24746 );
    or g18171 ( n16288 , n14879 , n16181 );
    not g18172 ( n10602 , n16924 );
    xnor g18173 ( n1721 , n12542 , n25525 );
    nor g18174 ( n12863 , n26312 , n23895 );
    xnor g18175 ( n6246 , n2865 , n21989 );
    xnor g18176 ( n13310 , n2705 , n18926 );
    nor g18177 ( n11790 , n22110 , n25485 );
    or g18178 ( n4806 , n2331 , n5506 );
    or g18179 ( n12154 , n12343 , n16357 );
    not g18180 ( n23704 , n11285 );
    and g18181 ( n20851 , n27176 , n25633 );
    and g18182 ( n7563 , n8680 , n7676 );
    and g18183 ( n11823 , n14262 , n20884 );
    nor g18184 ( n24453 , n13114 , n16283 );
    or g18185 ( n10778 , n23479 , n1383 );
    or g18186 ( n22310 , n3506 , n10658 );
    nor g18187 ( n1797 , n6518 , n6410 );
    not g18188 ( n18662 , n21287 );
    or g18189 ( n26365 , n10164 , n21703 );
    and g18190 ( n903 , n11156 , n595 );
    xnor g18191 ( n13565 , n5760 , n1754 );
    xnor g18192 ( n5288 , n13970 , n5805 );
    nor g18193 ( n7424 , n11467 , n26015 );
    xnor g18194 ( n16963 , n3358 , n7108 );
    and g18195 ( n10176 , n21546 , n24548 );
    and g18196 ( n13521 , n17616 , n9966 );
    or g18197 ( n25290 , n23163 , n10176 );
    or g18198 ( n3068 , n16294 , n1380 );
    xnor g18199 ( n16053 , n3980 , n1716 );
    and g18200 ( n8374 , n8673 , n26623 );
    xnor g18201 ( n26727 , n4789 , n14300 );
    not g18202 ( n16130 , n25241 );
    xnor g18203 ( n13209 , n5861 , n10347 );
    and g18204 ( n5756 , n7201 , n14403 );
    not g18205 ( n23539 , n5905 );
    or g18206 ( n2631 , n6422 , n24217 );
    or g18207 ( n4344 , n23707 , n3730 );
    or g18208 ( n5945 , n8322 , n19634 );
    or g18209 ( n18284 , n4717 , n15813 );
    or g18210 ( n9878 , n18060 , n19738 );
    nor g18211 ( n26043 , n19951 , n20655 );
    nor g18212 ( n22791 , n18926 , n6513 );
    xnor g18213 ( n24259 , n5313 , n24009 );
    xnor g18214 ( n26602 , n42 , n24648 );
    not g18215 ( n3690 , n8507 );
    and g18216 ( n24757 , n23521 , n21347 );
    not g18217 ( n21280 , n24873 );
    or g18218 ( n8512 , n5389 , n17313 );
    xnor g18219 ( n5020 , n2242 , n6225 );
    or g18220 ( n22301 , n14251 , n10349 );
    xnor g18221 ( n6450 , n15659 , n18537 );
    not g18222 ( n7892 , n22002 );
    or g18223 ( n20177 , n3249 , n10936 );
    and g18224 ( n22603 , n12429 , n15029 );
    xnor g18225 ( n20901 , n15468 , n4228 );
    xnor g18226 ( n21459 , n9098 , n25881 );
    xnor g18227 ( n8855 , n21392 , n18105 );
    not g18228 ( n24996 , n3906 );
    not g18229 ( n4555 , n22470 );
    and g18230 ( n10459 , n14232 , n11264 );
    xnor g18231 ( n6888 , n5122 , n13821 );
    xnor g18232 ( n24585 , n13643 , n3038 );
    or g18233 ( n11200 , n9986 , n3112 );
    xnor g18234 ( n11537 , n22429 , n6142 );
    or g18235 ( n17275 , n9198 , n37 );
    xnor g18236 ( n10554 , n21110 , n3270 );
    and g18237 ( n10601 , n25452 , n507 );
    not g18238 ( n12944 , n2446 );
    and g18239 ( n13862 , n8061 , n10972 );
    xnor g18240 ( n24767 , n24907 , n24485 );
    nor g18241 ( n26116 , n20592 , n16833 );
    xnor g18242 ( n12842 , n926 , n21125 );
    or g18243 ( n9092 , n26247 , n18135 );
    and g18244 ( n19692 , n2172 , n17315 );
    xnor g18245 ( n12809 , n6003 , n21547 );
    not g18246 ( n11294 , n12892 );
    nor g18247 ( n25819 , n19630 , n16642 );
    and g18248 ( n712 , n12919 , n3434 );
    and g18249 ( n2759 , n7952 , n1365 );
    not g18250 ( n23644 , n26851 );
    nor g18251 ( n16296 , n25879 , n6295 );
    xnor g18252 ( n20339 , n5402 , n7361 );
    not g18253 ( n13023 , n12209 );
    xnor g18254 ( n25289 , n25921 , n21753 );
    and g18255 ( n9799 , n16775 , n22214 );
    nor g18256 ( n11189 , n12950 , n949 );
    or g18257 ( n17268 , n18994 , n2100 );
    xnor g18258 ( n12275 , n8097 , n17210 );
    xnor g18259 ( n485 , n12824 , n16342 );
    or g18260 ( n1867 , n112 , n26264 );
    and g18261 ( n24605 , n11011 , n16711 );
    xnor g18262 ( n18463 , n23849 , n2289 );
    and g18263 ( n5798 , n5315 , n20387 );
    nor g18264 ( n21598 , n16092 , n24536 );
    not g18265 ( n15572 , n7191 );
    and g18266 ( n529 , n3398 , n164 );
    xnor g18267 ( n20505 , n11042 , n24569 );
    not g18268 ( n4940 , n8259 );
    and g18269 ( n9766 , n13719 , n22342 );
    or g18270 ( n7263 , n17872 , n9881 );
    nor g18271 ( n21844 , n11881 , n10225 );
    or g18272 ( n5635 , n23244 , n1801 );
    or g18273 ( n20528 , n1200 , n15254 );
    xnor g18274 ( n9838 , n15568 , n5928 );
    xnor g18275 ( n10965 , n15784 , n25797 );
    not g18276 ( n13480 , n21839 );
    xnor g18277 ( n26937 , n11734 , n22687 );
    nor g18278 ( n14747 , n21780 , n816 );
    or g18279 ( n15948 , n21292 , n654 );
    or g18280 ( n9607 , n18714 , n24745 );
    xnor g18281 ( n10367 , n24244 , n11577 );
    xnor g18282 ( n16419 , n22233 , n13825 );
    xnor g18283 ( n2968 , n9700 , n9969 );
    or g18284 ( n4483 , n9897 , n26711 );
    and g18285 ( n1439 , n13400 , n18283 );
    or g18286 ( n3339 , n23797 , n257 );
    and g18287 ( n10942 , n21589 , n24075 );
    not g18288 ( n15276 , n22805 );
    not g18289 ( n8838 , n9368 );
    nor g18290 ( n10047 , n19726 , n25583 );
    and g18291 ( n5150 , n10200 , n22777 );
    not g18292 ( n9477 , n24109 );
    xnor g18293 ( n440 , n23290 , n20002 );
    or g18294 ( n8397 , n16939 , n968 );
    not g18295 ( n19541 , n2113 );
    xnor g18296 ( n17325 , n19097 , n5333 );
    xnor g18297 ( n26884 , n24465 , n23647 );
    xnor g18298 ( n3748 , n14532 , n20826 );
    or g18299 ( n23621 , n25318 , n21728 );
    not g18300 ( n18768 , n5428 );
    xnor g18301 ( n16 , n851 , n17047 );
    nor g18302 ( n5280 , n14033 , n22797 );
    not g18303 ( n17517 , n15991 );
    xnor g18304 ( n26427 , n18649 , n3795 );
    or g18305 ( n15075 , n16387 , n507 );
    or g18306 ( n26715 , n3257 , n25243 );
    or g18307 ( n18076 , n7344 , n26147 );
    xnor g18308 ( n24447 , n10614 , n21898 );
    and g18309 ( n24688 , n4663 , n19390 );
    and g18310 ( n24262 , n23440 , n25197 );
    or g18311 ( n15951 , n22038 , n17548 );
    and g18312 ( n5159 , n25946 , n18867 );
    or g18313 ( n25157 , n24660 , n2787 );
    xnor g18314 ( n19585 , n14311 , n19895 );
    and g18315 ( n25186 , n25508 , n10052 );
    and g18316 ( n22769 , n26162 , n23556 );
    not g18317 ( n14794 , n4959 );
    xnor g18318 ( n9012 , n25292 , n8765 );
    xnor g18319 ( n14147 , n19492 , n7145 );
    xnor g18320 ( n8718 , n21875 , n20610 );
    not g18321 ( n18256 , n2518 );
    xnor g18322 ( n1865 , n2732 , n1432 );
    or g18323 ( n6572 , n2003 , n6063 );
    and g18324 ( n10988 , n3953 , n13996 );
    or g18325 ( n26627 , n24537 , n11210 );
    xnor g18326 ( n3222 , n10534 , n9366 );
    xnor g18327 ( n21111 , n4945 , n8482 );
    or g18328 ( n1331 , n11122 , n10849 );
    xnor g18329 ( n18455 , n24237 , n4017 );
    not g18330 ( n20667 , n6356 );
    or g18331 ( n8866 , n17558 , n1855 );
    or g18332 ( n22245 , n14383 , n2107 );
    or g18333 ( n5486 , n12543 , n5220 );
    xnor g18334 ( n24102 , n21672 , n19300 );
    xnor g18335 ( n9943 , n17447 , n25764 );
    nor g18336 ( n11884 , n11056 , n18157 );
    nor g18337 ( n21063 , n22626 , n26986 );
    not g18338 ( n17442 , n3420 );
    nor g18339 ( n16698 , n20700 , n932 );
    xnor g18340 ( n13166 , n26400 , n5453 );
    or g18341 ( n20276 , n18483 , n16314 );
    xnor g18342 ( n24292 , n10925 , n22538 );
    and g18343 ( n23297 , n15627 , n15896 );
    nor g18344 ( n9351 , n9711 , n10980 );
    or g18345 ( n25354 , n63 , n25240 );
    and g18346 ( n13854 , n10282 , n4444 );
    and g18347 ( n23845 , n1152 , n10917 );
    and g18348 ( n6803 , n12160 , n10562 );
    or g18349 ( n5759 , n9433 , n11858 );
    xnor g18350 ( n16185 , n17818 , n20144 );
    not g18351 ( n24923 , n22704 );
    xnor g18352 ( n21409 , n1558 , n11566 );
    not g18353 ( n6809 , n12070 );
    xnor g18354 ( n4205 , n5245 , n2326 );
    and g18355 ( n19175 , n4721 , n13930 );
    nor g18356 ( n6759 , n26834 , n5709 );
    and g18357 ( n3767 , n7081 , n24213 );
    nor g18358 ( n10794 , n21779 , n24392 );
    and g18359 ( n17060 , n18629 , n19964 );
    nor g18360 ( n16668 , n25324 , n14148 );
    or g18361 ( n943 , n1896 , n4542 );
    or g18362 ( n8204 , n6753 , n3220 );
    or g18363 ( n10688 , n6778 , n21214 );
    xnor g18364 ( n12683 , n3591 , n3963 );
    nor g18365 ( n23623 , n25389 , n13339 );
    xnor g18366 ( n19496 , n3497 , n3207 );
    or g18367 ( n24352 , n16195 , n1853 );
    xnor g18368 ( n7478 , n26942 , n22634 );
    and g18369 ( n17788 , n8634 , n893 );
    xnor g18370 ( n25230 , n7242 , n25277 );
    xnor g18371 ( n17255 , n17624 , n12632 );
    or g18372 ( n9724 , n9880 , n1152 );
    xnor g18373 ( n11613 , n25724 , n24503 );
    not g18374 ( n10962 , n20927 );
    not g18375 ( n17189 , n4362 );
    or g18376 ( n23470 , n15695 , n583 );
    nor g18377 ( n6932 , n6154 , n21097 );
    or g18378 ( n3522 , n9035 , n9494 );
    nor g18379 ( n1524 , n6940 , n868 );
    xnor g18380 ( n23460 , n19993 , n10511 );
    xnor g18381 ( n11849 , n27203 , n1550 );
    or g18382 ( n18678 , n14965 , n10389 );
    and g18383 ( n15484 , n17175 , n3558 );
    nor g18384 ( n14554 , n6161 , n21793 );
    nor g18385 ( n8413 , n16600 , n11614 );
    xnor g18386 ( n3593 , n12149 , n7447 );
    or g18387 ( n15776 , n26814 , n934 );
    xnor g18388 ( n2918 , n20275 , n26986 );
    nor g18389 ( n1826 , n25558 , n21 );
    or g18390 ( n21500 , n24733 , n2806 );
    xnor g18391 ( n4660 , n22096 , n20850 );
    nor g18392 ( n5297 , n27142 , n2410 );
    and g18393 ( n6681 , n21169 , n10717 );
    nor g18394 ( n979 , n6841 , n13935 );
    nor g18395 ( n20905 , n17287 , n21287 );
    and g18396 ( n25777 , n10507 , n26205 );
    or g18397 ( n3367 , n2812 , n17645 );
    or g18398 ( n9970 , n14816 , n18318 );
    xnor g18399 ( n6287 , n19097 , n7949 );
    nor g18400 ( n20787 , n16889 , n18105 );
    or g18401 ( n26203 , n17358 , n7994 );
    xnor g18402 ( n16368 , n20542 , n25937 );
    not g18403 ( n8351 , n12637 );
    nor g18404 ( n8396 , n18925 , n25150 );
    not g18405 ( n24217 , n16091 );
    not g18406 ( n9908 , n17302 );
    xnor g18407 ( n13764 , n20204 , n14905 );
    and g18408 ( n1772 , n24621 , n7196 );
    and g18409 ( n22604 , n14044 , n91 );
    or g18410 ( n8506 , n26428 , n1085 );
    not g18411 ( n21246 , n23900 );
    and g18412 ( n7654 , n21887 , n12061 );
    or g18413 ( n11156 , n22865 , n12 );
    or g18414 ( n1087 , n5331 , n24960 );
    not g18415 ( n12049 , n13447 );
    nor g18416 ( n26267 , n21416 , n4773 );
    and g18417 ( n10319 , n12880 , n16229 );
    nor g18418 ( n17328 , n12396 , n24937 );
    or g18419 ( n1133 , n11624 , n14299 );
    xnor g18420 ( n27004 , n25493 , n7372 );
    xnor g18421 ( n4936 , n23697 , n19531 );
    xnor g18422 ( n18635 , n18380 , n22806 );
    xnor g18423 ( n10680 , n20811 , n19047 );
    nor g18424 ( n17125 , n15365 , n1973 );
    or g18425 ( n21725 , n6134 , n1707 );
    and g18426 ( n5277 , n6385 , n23030 );
    xnor g18427 ( n18011 , n8398 , n710 );
    or g18428 ( n5272 , n1406 , n19473 );
    or g18429 ( n1175 , n5934 , n983 );
    and g18430 ( n1953 , n7297 , n24102 );
    not g18431 ( n7915 , n20957 );
    xnor g18432 ( n24051 , n10855 , n671 );
    not g18433 ( n22700 , n2005 );
    xnor g18434 ( n7119 , n587 , n22452 );
    and g18435 ( n16742 , n3393 , n1465 );
    and g18436 ( n19008 , n17096 , n22950 );
    xnor g18437 ( n17291 , n5756 , n7467 );
    xnor g18438 ( n9270 , n20527 , n5880 );
    not g18439 ( n7966 , n6127 );
    not g18440 ( n13474 , n21759 );
    xnor g18441 ( n23142 , n7857 , n5060 );
    or g18442 ( n8912 , n8630 , n18696 );
    xnor g18443 ( n253 , n24948 , n11322 );
    nor g18444 ( n25450 , n10001 , n21263 );
    xnor g18445 ( n21496 , n16278 , n8259 );
    nor g18446 ( n21512 , n16755 , n23493 );
    not g18447 ( n4371 , n7191 );
    or g18448 ( n25072 , n4748 , n21029 );
    or g18449 ( n3399 , n23088 , n4668 );
    not g18450 ( n24044 , n10763 );
    or g18451 ( n20095 , n20205 , n4256 );
    and g18452 ( n17321 , n1374 , n22728 );
    not g18453 ( n2151 , n6686 );
    nor g18454 ( n22196 , n13907 , n12493 );
    or g18455 ( n3838 , n8552 , n17167 );
    xnor g18456 ( n5853 , n19360 , n19042 );
    not g18457 ( n9233 , n19711 );
    xnor g18458 ( n23309 , n25877 , n22619 );
    or g18459 ( n16649 , n14133 , n9570 );
    or g18460 ( n8556 , n5605 , n23587 );
    and g18461 ( n20631 , n15976 , n8093 );
    or g18462 ( n26310 , n24359 , n19319 );
    and g18463 ( n14376 , n5464 , n14065 );
    nor g18464 ( n13340 , n11802 , n11502 );
    xnor g18465 ( n20804 , n2656 , n6851 );
    not g18466 ( n18781 , n25906 );
    nor g18467 ( n16444 , n1594 , n762 );
    and g18468 ( n11484 , n17271 , n7159 );
    or g18469 ( n25960 , n18012 , n10776 );
    xnor g18470 ( n24431 , n13020 , n19114 );
    and g18471 ( n6813 , n11155 , n972 );
    xnor g18472 ( n10895 , n10625 , n11481 );
    and g18473 ( n25599 , n26750 , n19538 );
    not g18474 ( n13349 , n4319 );
    not g18475 ( n7597 , n4872 );
    and g18476 ( n25026 , n5097 , n3394 );
    or g18477 ( n14605 , n21520 , n7536 );
    not g18478 ( n17022 , n24315 );
    xnor g18479 ( n25086 , n21636 , n26107 );
    and g18480 ( n6399 , n1977 , n5878 );
    not g18481 ( n9668 , n25881 );
    or g18482 ( n20798 , n11473 , n27 );
    not g18483 ( n7653 , n18194 );
    and g18484 ( n3458 , n14189 , n14795 );
    xnor g18485 ( n3697 , n8100 , n22211 );
    and g18486 ( n13265 , n10627 , n18913 );
    or g18487 ( n22025 , n18420 , n16532 );
    not g18488 ( n9723 , n20557 );
    not g18489 ( n7578 , n8657 );
    or g18490 ( n26005 , n8579 , n27206 );
    xnor g18491 ( n10174 , n767 , n22793 );
    or g18492 ( n6260 , n7066 , n9413 );
    xnor g18493 ( n11935 , n17409 , n10258 );
    and g18494 ( n25729 , n7320 , n25560 );
    xnor g18495 ( n15268 , n3706 , n15539 );
    xnor g18496 ( n25130 , n8391 , n7917 );
    and g18497 ( n4610 , n18325 , n14219 );
    xnor g18498 ( n10561 , n21689 , n16175 );
    xnor g18499 ( n22552 , n20999 , n24029 );
    xnor g18500 ( n5206 , n17060 , n26206 );
    not g18501 ( n23956 , n25937 );
    xnor g18502 ( n26634 , n17222 , n2598 );
    xnor g18503 ( n2073 , n18821 , n9975 );
    or g18504 ( n13623 , n13000 , n13997 );
    and g18505 ( n16079 , n23800 , n1308 );
    and g18506 ( n6642 , n11673 , n11948 );
    xnor g18507 ( n3451 , n8901 , n409 );
    and g18508 ( n13240 , n24038 , n5894 );
    xnor g18509 ( n15679 , n1541 , n7524 );
    or g18510 ( n6368 , n23529 , n10739 );
    not g18511 ( n18575 , n9160 );
    and g18512 ( n12561 , n2156 , n7402 );
    or g18513 ( n370 , n20662 , n16533 );
    or g18514 ( n23703 , n21420 , n21768 );
    not g18515 ( n8648 , n12492 );
    or g18516 ( n15233 , n5816 , n13981 );
    not g18517 ( n20544 , n19042 );
    xnor g18518 ( n15683 , n6510 , n5031 );
    or g18519 ( n20350 , n20474 , n19871 );
    or g18520 ( n20363 , n26127 , n648 );
    and g18521 ( n16271 , n14068 , n17335 );
    or g18522 ( n22111 , n26197 , n19003 );
    or g18523 ( n22276 , n20121 , n18235 );
    xnor g18524 ( n10432 , n16750 , n16981 );
    xnor g18525 ( n13493 , n8780 , n16479 );
    or g18526 ( n20487 , n3297 , n13143 );
    xnor g18527 ( n13036 , n4388 , n23131 );
    or g18528 ( n6519 , n4430 , n16666 );
    nor g18529 ( n26982 , n15875 , n13352 );
    xnor g18530 ( n7975 , n26095 , n24461 );
    and g18531 ( n2014 , n18777 , n8815 );
    xnor g18532 ( n5399 , n15686 , n5771 );
    xnor g18533 ( n15225 , n14487 , n4330 );
    xnor g18534 ( n1925 , n4755 , n25802 );
    not g18535 ( n17881 , n3319 );
    and g18536 ( n153 , n1437 , n12488 );
    or g18537 ( n17697 , n7644 , n11235 );
    nor g18538 ( n45 , n16476 , n19146 );
    xnor g18539 ( n16851 , n18537 , n4376 );
    xnor g18540 ( n2764 , n14686 , n2433 );
    nor g18541 ( n3438 , n4967 , n26541 );
    or g18542 ( n23584 , n23950 , n23002 );
    not g18543 ( n20181 , n7083 );
    or g18544 ( n25391 , n20338 , n13034 );
    not g18545 ( n19489 , n3173 );
    and g18546 ( n24716 , n2355 , n115 );
    or g18547 ( n19661 , n1188 , n22427 );
    not g18548 ( n15265 , n25073 );
    and g18549 ( n7379 , n12490 , n19824 );
    xnor g18550 ( n26228 , n12991 , n24700 );
    or g18551 ( n9355 , n14481 , n17145 );
    and g18552 ( n11909 , n14936 , n15233 );
    and g18553 ( n22544 , n4784 , n2603 );
    and g18554 ( n15492 , n5869 , n19492 );
    nor g18555 ( n16678 , n3138 , n2829 );
    xnor g18556 ( n19552 , n24420 , n12398 );
    xnor g18557 ( n20331 , n25289 , n5255 );
    xnor g18558 ( n18482 , n19416 , n14983 );
    xnor g18559 ( n24421 , n5045 , n7781 );
    xnor g18560 ( n2061 , n1710 , n23284 );
    nor g18561 ( n3302 , n3266 , n3028 );
    xnor g18562 ( n323 , n26880 , n1693 );
    xnor g18563 ( n17715 , n5244 , n14852 );
    xnor g18564 ( n3056 , n18484 , n23855 );
    or g18565 ( n15563 , n1329 , n1152 );
    not g18566 ( n2096 , n14011 );
    and g18567 ( n23564 , n22823 , n19213 );
    xnor g18568 ( n24465 , n26577 , n1074 );
    and g18569 ( n14910 , n17728 , n18319 );
    and g18570 ( n14272 , n12507 , n15739 );
    or g18571 ( n14026 , n6753 , n3376 );
    and g18572 ( n16736 , n26435 , n14903 );
    or g18573 ( n4993 , n2429 , n15961 );
    or g18574 ( n16124 , n4097 , n8527 );
    xnor g18575 ( n12086 , n5830 , n17288 );
    or g18576 ( n20167 , n20993 , n22648 );
    not g18577 ( n18643 , n19303 );
    not g18578 ( n12143 , n19842 );
    xnor g18579 ( n2457 , n24327 , n4325 );
    xnor g18580 ( n16840 , n15443 , n15397 );
    xnor g18581 ( n20517 , n14871 , n23613 );
    nor g18582 ( n25526 , n421 , n15272 );
    or g18583 ( n20028 , n12735 , n11986 );
    xnor g18584 ( n12749 , n18915 , n6662 );
    nor g18585 ( n19688 , n23645 , n22068 );
    or g18586 ( n14039 , n23056 , n10371 );
    and g18587 ( n4471 , n21517 , n8582 );
    and g18588 ( n21084 , n23518 , n12830 );
    or g18589 ( n10197 , n23213 , n4883 );
    nor g18590 ( n14100 , n25268 , n20883 );
    xnor g18591 ( n14236 , n2886 , n1738 );
    xnor g18592 ( n19252 , n13263 , n21779 );
    xnor g18593 ( n24092 , n7500 , n19266 );
    and g18594 ( n8841 , n11592 , n14003 );
    or g18595 ( n7801 , n22170 , n4007 );
    and g18596 ( n9931 , n12915 , n13012 );
    or g18597 ( n20587 , n21100 , n17445 );
    nor g18598 ( n20083 , n2473 , n20203 );
    not g18599 ( n1404 , n22588 );
    and g18600 ( n4864 , n279 , n9891 );
    nor g18601 ( n15623 , n23849 , n2289 );
    or g18602 ( n15664 , n12328 , n20663 );
    xnor g18603 ( n25358 , n15008 , n16476 );
    xnor g18604 ( n3463 , n11733 , n26789 );
    xnor g18605 ( n20575 , n2781 , n18102 );
    xnor g18606 ( n1884 , n18617 , n18452 );
    or g18607 ( n689 , n10471 , n8600 );
    or g18608 ( n13815 , n4040 , n16009 );
    and g18609 ( n6049 , n15410 , n20969 );
    not g18610 ( n6701 , n12900 );
    nor g18611 ( n786 , n8419 , n17067 );
    xnor g18612 ( n7752 , n7150 , n2229 );
    or g18613 ( n20372 , n6659 , n12991 );
    not g18614 ( n3112 , n17412 );
    xnor g18615 ( n26796 , n5194 , n16743 );
    or g18616 ( n7936 , n1882 , n12311 );
    nor g18617 ( n18677 , n12112 , n9404 );
    nor g18618 ( n16293 , n12426 , n11476 );
    nor g18619 ( n16355 , n24620 , n7099 );
    and g18620 ( n4911 , n14141 , n4827 );
    xnor g18621 ( n20118 , n9770 , n19143 );
    xnor g18622 ( n1660 , n27120 , n23065 );
    not g18623 ( n14614 , n13303 );
    xnor g18624 ( n16407 , n20312 , n12352 );
    or g18625 ( n10676 , n22830 , n7171 );
    xnor g18626 ( n17870 , n17135 , n16441 );
    not g18627 ( n9401 , n7421 );
    and g18628 ( n12574 , n20977 , n18076 );
    xnor g18629 ( n25693 , n96 , n8249 );
    and g18630 ( n2271 , n20793 , n24528 );
    xnor g18631 ( n12886 , n9493 , n3918 );
    or g18632 ( n14626 , n5253 , n20146 );
    and g18633 ( n25304 , n21166 , n10811 );
    or g18634 ( n4589 , n17711 , n8398 );
    nor g18635 ( n18960 , n11542 , n18247 );
    and g18636 ( n14617 , n7172 , n19806 );
    xnor g18637 ( n7002 , n16863 , n24816 );
    and g18638 ( n2222 , n8739 , n23655 );
    xnor g18639 ( n13468 , n21464 , n14092 );
    and g18640 ( n24186 , n2641 , n16036 );
    nor g18641 ( n13239 , n7892 , n2718 );
    or g18642 ( n22758 , n11116 , n7825 );
    nor g18643 ( n16015 , n19472 , n24473 );
    xnor g18644 ( n3062 , n17111 , n6829 );
    or g18645 ( n25678 , n7907 , n6455 );
    not g18646 ( n5465 , n17299 );
    or g18647 ( n17270 , n20216 , n3524 );
    or g18648 ( n19145 , n23159 , n9161 );
    not g18649 ( n9603 , n20595 );
    xnor g18650 ( n13450 , n11220 , n3425 );
    xnor g18651 ( n7366 , n2656 , n16929 );
    not g18652 ( n1334 , n21398 );
    and g18653 ( n6259 , n15060 , n10754 );
    or g18654 ( n118 , n5298 , n2359 );
    or g18655 ( n26655 , n1957 , n5197 );
    or g18656 ( n20136 , n17945 , n5787 );
    not g18657 ( n12592 , n1545 );
    and g18658 ( n24132 , n8651 , n178 );
    nor g18659 ( n13461 , n19061 , n9935 );
    or g18660 ( n23342 , n1923 , n17129 );
    or g18661 ( n13532 , n26988 , n21542 );
    xnor g18662 ( n4401 , n13678 , n1854 );
    and g18663 ( n2767 , n21243 , n12331 );
    not g18664 ( n7743 , n18274 );
    or g18665 ( n8051 , n8361 , n1483 );
    xnor g18666 ( n24145 , n18267 , n17765 );
    or g18667 ( n12460 , n25589 , n16831 );
    not g18668 ( n17909 , n21674 );
    not g18669 ( n18079 , n14809 );
    or g18670 ( n14233 , n20733 , n7330 );
    xnor g18671 ( n911 , n839 , n6139 );
    nor g18672 ( n12140 , n10683 , n23832 );
    and g18673 ( n625 , n20370 , n3401 );
    nor g18674 ( n23711 , n11184 , n19366 );
    and g18675 ( n22264 , n24179 , n7998 );
    not g18676 ( n550 , n9397 );
    not g18677 ( n15906 , n24628 );
    or g18678 ( n17025 , n2250 , n4324 );
    or g18679 ( n27083 , n10552 , n2879 );
    or g18680 ( n9176 , n9513 , n23417 );
    xnor g18681 ( n18830 , n8060 , n1695 );
    xnor g18682 ( n4640 , n10024 , n7347 );
    xnor g18683 ( n14841 , n6963 , n25974 );
    xnor g18684 ( n10899 , n6241 , n17462 );
    nor g18685 ( n21174 , n8381 , n12889 );
    not g18686 ( n24510 , n7765 );
    nor g18687 ( n2640 , n19667 , n4272 );
    xnor g18688 ( n22456 , n20283 , n6939 );
    or g18689 ( n18270 , n22855 , n26410 );
    xnor g18690 ( n8033 , n4930 , n21134 );
    or g18691 ( n13746 , n13890 , n12336 );
    xnor g18692 ( n7579 , n7689 , n25115 );
    or g18693 ( n1290 , n11321 , n3746 );
    and g18694 ( n11628 , n14662 , n13187 );
    or g18695 ( n5487 , n5842 , n13429 );
    or g18696 ( n25754 , n11685 , n3890 );
    or g18697 ( n24241 , n13378 , n13459 );
    and g18698 ( n12471 , n25094 , n3049 );
    not g18699 ( n10634 , n13905 );
    and g18700 ( n2476 , n17351 , n21850 );
    or g18701 ( n841 , n5431 , n13469 );
    not g18702 ( n13831 , n23558 );
    and g18703 ( n5899 , n14230 , n19922 );
    xnor g18704 ( n973 , n280 , n13875 );
    not g18705 ( n1655 , n26011 );
    or g18706 ( n19470 , n22166 , n23607 );
    or g18707 ( n13232 , n18378 , n16504 );
    xnor g18708 ( n23835 , n19198 , n22684 );
    not g18709 ( n10684 , n18322 );
    and g18710 ( n2867 , n22164 , n19188 );
    nor g18711 ( n10655 , n5266 , n11428 );
    xnor g18712 ( n7238 , n5001 , n7693 );
    xnor g18713 ( n2897 , n18360 , n11644 );
    and g18714 ( n20170 , n23486 , n16663 );
    or g18715 ( n21343 , n14337 , n4940 );
    or g18716 ( n18913 , n20242 , n12724 );
    or g18717 ( n11250 , n22656 , n3328 );
    or g18718 ( n21388 , n21380 , n5211 );
    or g18719 ( n13076 , n4376 , n19080 );
    or g18720 ( n22982 , n5060 , n15380 );
    or g18721 ( n10170 , n3709 , n8969 );
    and g18722 ( n21359 , n22841 , n9935 );
    or g18723 ( n16610 , n23910 , n21339 );
    or g18724 ( n11107 , n20323 , n8564 );
    nor g18725 ( n1454 , n48 , n8714 );
    xnor g18726 ( n108 , n17009 , n11376 );
    or g18727 ( n22354 , n1826 , n22505 );
    xnor g18728 ( n17227 , n9125 , n10631 );
    or g18729 ( n16141 , n21015 , n11452 );
    xnor g18730 ( n16433 , n16732 , n13056 );
    or g18731 ( n4992 , n6379 , n10923 );
    and g18732 ( n2998 , n1311 , n24270 );
    or g18733 ( n10559 , n11425 , n19531 );
    not g18734 ( n5714 , n2816 );
    or g18735 ( n23902 , n16320 , n3304 );
    or g18736 ( n16248 , n19850 , n24443 );
    or g18737 ( n11942 , n13752 , n20304 );
    xnor g18738 ( n7753 , n6385 , n16223 );
    buf g18739 ( n22169 , n7725 );
    or g18740 ( n4973 , n23075 , n18566 );
    xnor g18741 ( n13801 , n9476 , n21924 );
    or g18742 ( n4369 , n16232 , n4509 );
    not g18743 ( n22851 , n13677 );
    or g18744 ( n5397 , n10403 , n21668 );
    xnor g18745 ( n7825 , n17520 , n5058 );
    and g18746 ( n16348 , n18161 , n23205 );
    or g18747 ( n11041 , n16211 , n7437 );
    nor g18748 ( n6780 , n4780 , n21922 );
    and g18749 ( n10208 , n13516 , n17761 );
    nor g18750 ( n13901 , n7893 , n5400 );
    or g18751 ( n9639 , n2160 , n27095 );
    xnor g18752 ( n9730 , n24705 , n21460 );
    not g18753 ( n14365 , n8717 );
    or g18754 ( n5257 , n23008 , n17640 );
    and g18755 ( n26403 , n5655 , n26655 );
    nor g18756 ( n25763 , n19868 , n19742 );
    not g18757 ( n2482 , n16359 );
    nor g18758 ( n1139 , n19328 , n16123 );
    or g18759 ( n467 , n1847 , n18240 );
    xnor g18760 ( n3291 , n13696 , n7470 );
    or g18761 ( n6004 , n11758 , n12457 );
    not g18762 ( n17677 , n336 );
    xnor g18763 ( n21231 , n7775 , n6848 );
    not g18764 ( n12512 , n14352 );
    not g18765 ( n7195 , n1255 );
    or g18766 ( n26432 , n1180 , n1206 );
    or g18767 ( n18222 , n11870 , n184 );
    not g18768 ( n14498 , n19475 );
    xnor g18769 ( n510 , n4326 , n3952 );
    or g18770 ( n23017 , n1965 , n6220 );
    and g18771 ( n7862 , n18403 , n18956 );
    not g18772 ( n2135 , n20343 );
    and g18773 ( n10902 , n12792 , n2064 );
    or g18774 ( n6144 , n20913 , n5150 );
    nor g18775 ( n8238 , n4769 , n11176 );
    or g18776 ( n3629 , n12396 , n8297 );
    xnor g18777 ( n1499 , n15502 , n8553 );
    nor g18778 ( n17768 , n9402 , n23209 );
    and g18779 ( n13870 , n8678 , n3882 );
    not g18780 ( n18261 , n25694 );
    xnor g18781 ( n17576 , n7057 , n12956 );
    or g18782 ( n8158 , n19313 , n13354 );
    nor g18783 ( n10387 , n25172 , n16545 );
    not g18784 ( n18016 , n6475 );
    or g18785 ( n5730 , n9187 , n4870 );
    xnor g18786 ( n22283 , n11616 , n18534 );
    not g18787 ( n15010 , n6410 );
    or g18788 ( n1459 , n21984 , n6255 );
    or g18789 ( n14425 , n9588 , n14505 );
    xnor g18790 ( n26771 , n27089 , n12657 );
    and g18791 ( n3521 , n26443 , n10017 );
    not g18792 ( n16792 , n24543 );
    xnor g18793 ( n26024 , n14411 , n18243 );
    or g18794 ( n22516 , n25556 , n7938 );
    or g18795 ( n25055 , n15534 , n23885 );
    xnor g18796 ( n6983 , n22604 , n17589 );
    not g18797 ( n15008 , n25805 );
    xnor g18798 ( n13426 , n25538 , n7305 );
    not g18799 ( n24615 , n4590 );
    or g18800 ( n12213 , n21766 , n9480 );
    or g18801 ( n16352 , n24760 , n26721 );
    and g18802 ( n14844 , n16894 , n25803 );
    xnor g18803 ( n25498 , n9365 , n23541 );
    xnor g18804 ( n27118 , n7854 , n6903 );
    not g18805 ( n22036 , n7552 );
    xnor g18806 ( n24144 , n2815 , n10455 );
    or g18807 ( n15680 , n3169 , n8622 );
    or g18808 ( n17113 , n7109 , n19536 );
    nor g18809 ( n23386 , n11045 , n19282 );
    and g18810 ( n2009 , n2662 , n22969 );
    or g18811 ( n3481 , n752 , n11504 );
    nor g18812 ( n2986 , n23160 , n3570 );
    nor g18813 ( n3796 , n3178 , n10614 );
    and g18814 ( n2882 , n15551 , n25678 );
    not g18815 ( n1547 , n13393 );
    xnor g18816 ( n16199 , n7430 , n11996 );
    not g18817 ( n9241 , n25768 );
    xnor g18818 ( n24643 , n15047 , n8286 );
    or g18819 ( n14741 , n10318 , n18752 );
    or g18820 ( n9745 , n15096 , n10143 );
    xnor g18821 ( n15180 , n8755 , n26406 );
    xnor g18822 ( n5354 , n27137 , n26800 );
    xnor g18823 ( n19899 , n6934 , n14622 );
    and g18824 ( n10415 , n17503 , n15833 );
    not g18825 ( n23525 , n685 );
    and g18826 ( n9744 , n5355 , n19962 );
    or g18827 ( n3412 , n10083 , n18928 );
    and g18828 ( n2450 , n9495 , n10073 );
    and g18829 ( n20119 , n21424 , n1318 );
    not g18830 ( n17122 , n25603 );
    or g18831 ( n23078 , n10088 , n21185 );
    or g18832 ( n11742 , n11394 , n5419 );
    not g18833 ( n9514 , n7285 );
    xnor g18834 ( n12205 , n18027 , n19137 );
    xnor g18835 ( n15721 , n14958 , n17888 );
    not g18836 ( n3848 , n2279 );
    xnor g18837 ( n26371 , n6666 , n10355 );
    nor g18838 ( n8741 , n17323 , n5555 );
    nor g18839 ( n12242 , n20000 , n20665 );
    or g18840 ( n2263 , n24366 , n24695 );
    or g18841 ( n11074 , n11630 , n18504 );
    xnor g18842 ( n22511 , n25035 , n10297 );
    xnor g18843 ( n11462 , n20537 , n21044 );
    or g18844 ( n25817 , n13036 , n23307 );
    and g18845 ( n24814 , n6649 , n17570 );
    xnor g18846 ( n4816 , n18895 , n26318 );
    or g18847 ( n3923 , n15175 , n11098 );
    or g18848 ( n1241 , n6653 , n15569 );
    xnor g18849 ( n19367 , n7687 , n23123 );
    xnor g18850 ( n20477 , n13193 , n5866 );
    xnor g18851 ( n14386 , n9385 , n25131 );
    or g18852 ( n13937 , n14390 , n21684 );
    and g18853 ( n15432 , n8068 , n1128 );
    xnor g18854 ( n9126 , n3625 , n13089 );
    or g18855 ( n4515 , n17579 , n3320 );
    or g18856 ( n4142 , n26915 , n8549 );
    or g18857 ( n9105 , n613 , n8961 );
    or g18858 ( n26336 , n4241 , n11160 );
    or g18859 ( n12369 , n20998 , n2576 );
    nor g18860 ( n14502 , n23144 , n8439 );
    xnor g18861 ( n23222 , n26495 , n23620 );
    and g18862 ( n4062 , n744 , n18630 );
    or g18863 ( n12166 , n5768 , n24988 );
    and g18864 ( n7540 , n2974 , n16031 );
    xnor g18865 ( n21675 , n26797 , n24196 );
    and g18866 ( n18546 , n20429 , n22909 );
    xnor g18867 ( n2693 , n3510 , n464 );
    and g18868 ( n2333 , n13619 , n11886 );
    xnor g18869 ( n13753 , n24851 , n9251 );
    or g18870 ( n2270 , n22566 , n19317 );
    and g18871 ( n6363 , n26911 , n16566 );
    xnor g18872 ( n2965 , n5970 , n12570 );
    xnor g18873 ( n12367 , n2873 , n17813 );
    nor g18874 ( n16417 , n18326 , n1230 );
    xnor g18875 ( n21544 , n15233 , n11920 );
    or g18876 ( n8216 , n20599 , n2562 );
    nor g18877 ( n10211 , n1293 , n25413 );
    or g18878 ( n25002 , n20119 , n3168 );
    or g18879 ( n11616 , n19704 , n6469 );
    xnor g18880 ( n24342 , n1556 , n15835 );
    or g18881 ( n7265 , n24114 , n22067 );
    and g18882 ( n22582 , n16624 , n9408 );
    or g18883 ( n10370 , n27136 , n26270 );
    or g18884 ( n26338 , n18818 , n24874 );
    not g18885 ( n12190 , n7289 );
    not g18886 ( n10333 , n5582 );
    xnor g18887 ( n24200 , n5038 , n20483 );
    not g18888 ( n1577 , n13895 );
    or g18889 ( n9563 , n9908 , n19843 );
    nor g18890 ( n85 , n14465 , n15426 );
    xnor g18891 ( n14304 , n22626 , n8856 );
    and g18892 ( n2798 , n9469 , n3237 );
    xnor g18893 ( n9422 , n25119 , n23529 );
    and g18894 ( n4222 , n11501 , n22852 );
    not g18895 ( n6566 , n26857 );
    not g18896 ( n10734 , n2893 );
    xnor g18897 ( n19802 , n19331 , n23910 );
    xnor g18898 ( n15666 , n468 , n1255 );
    or g18899 ( n14842 , n2514 , n26883 );
    and g18900 ( n1592 , n21371 , n18106 );
    or g18901 ( n17007 , n512 , n11571 );
    not g18902 ( n16229 , n18446 );
    and g18903 ( n14591 , n4823 , n10939 );
    or g18904 ( n9369 , n22204 , n13589 );
    or g18905 ( n10724 , n19970 , n3106 );
    not g18906 ( n25014 , n1481 );
    or g18907 ( n9562 , n8576 , n26243 );
    not g18908 ( n12343 , n9140 );
    xnor g18909 ( n4014 , n14592 , n15278 );
    nor g18910 ( n22710 , n2658 , n23172 );
    and g18911 ( n9425 , n7184 , n20564 );
    and g18912 ( n15203 , n14426 , n25159 );
    xnor g18913 ( n9043 , n23005 , n11531 );
    xnor g18914 ( n17478 , n23271 , n7670 );
    or g18915 ( n27059 , n21386 , n23697 );
    and g18916 ( n20000 , n6353 , n12391 );
    and g18917 ( n2405 , n21156 , n24124 );
    nor g18918 ( n718 , n8032 , n12161 );
    not g18919 ( n14881 , n6679 );
    xnor g18920 ( n14216 , n15932 , n16163 );
    nor g18921 ( n26813 , n20588 , n16131 );
    or g18922 ( n26906 , n18954 , n23600 );
    and g18923 ( n19662 , n26180 , n24700 );
    xnor g18924 ( n6362 , n7243 , n20963 );
    xnor g18925 ( n4257 , n2731 , n4376 );
    or g18926 ( n2866 , n791 , n11322 );
    xnor g18927 ( n5929 , n23746 , n7269 );
    or g18928 ( n24220 , n11583 , n1138 );
    nor g18929 ( n11226 , n161 , n12780 );
    nor g18930 ( n5189 , n7777 , n23751 );
    or g18931 ( n9811 , n7807 , n13846 );
    or g18932 ( n27094 , n8252 , n11850 );
    and g18933 ( n17324 , n3059 , n17361 );
    xnor g18934 ( n9370 , n11600 , n16843 );
    or g18935 ( n3715 , n7517 , n24318 );
    or g18936 ( n697 , n15841 , n24808 );
    and g18937 ( n13196 , n18380 , n25645 );
    or g18938 ( n19653 , n6446 , n20060 );
    and g18939 ( n15520 , n16935 , n16691 );
    or g18940 ( n5444 , n12224 , n25829 );
    and g18941 ( n3646 , n5554 , n21461 );
    or g18942 ( n8223 , n7670 , n3253 );
    nor g18943 ( n14309 , n21846 , n25370 );
    xnor g18944 ( n1913 , n24999 , n23594 );
    xnor g18945 ( n21115 , n5171 , n3550 );
    xnor g18946 ( n13685 , n26952 , n17504 );
    nor g18947 ( n17209 , n22432 , n14808 );
    and g18948 ( n19655 , n7969 , n9640 );
    and g18949 ( n21953 , n22803 , n26873 );
    or g18950 ( n6901 , n24226 , n3112 );
    xnor g18951 ( n23653 , n27164 , n7868 );
    or g18952 ( n17214 , n17470 , n25998 );
    or g18953 ( n26643 , n4041 , n3378 );
    and g18954 ( n2925 , n408 , n19853 );
    nor g18955 ( n19347 , n17198 , n2923 );
    or g18956 ( n7222 , n4622 , n27089 );
    or g18957 ( n19243 , n4542 , n2586 );
    and g18958 ( n23928 , n6454 , n5476 );
    xnor g18959 ( n1357 , n3762 , n1862 );
    or g18960 ( n3775 , n4897 , n26819 );
    or g18961 ( n27034 , n16444 , n16284 );
    and g18962 ( n27038 , n7841 , n4941 );
    or g18963 ( n14611 , n436 , n13464 );
    or g18964 ( n12584 , n13523 , n6917 );
    and g18965 ( n26777 , n19531 , n21322 );
    or g18966 ( n19348 , n9987 , n4094 );
    not g18967 ( n15482 , n25210 );
    or g18968 ( n19861 , n9053 , n8974 );
    not g18969 ( n11088 , n9993 );
    or g18970 ( n15589 , n22527 , n2268 );
    xnor g18971 ( n1214 , n3632 , n682 );
    xnor g18972 ( n14622 , n21997 , n19701 );
    and g18973 ( n11430 , n2195 , n21197 );
    xnor g18974 ( n2971 , n12374 , n7695 );
    xnor g18975 ( n17225 , n6356 , n12956 );
    and g18976 ( n19110 , n24131 , n1088 );
    or g18977 ( n24532 , n20489 , n21693 );
    or g18978 ( n2276 , n24762 , n21862 );
    and g18979 ( n16114 , n14239 , n23672 );
    or g18980 ( n8161 , n12543 , n23793 );
    and g18981 ( n16620 , n4613 , n6561 );
    not g18982 ( n13523 , n27015 );
    xnor g18983 ( n19572 , n11871 , n987 );
    not g18984 ( n15400 , n14298 );
    xnor g18985 ( n9946 , n12993 , n23987 );
    or g18986 ( n26262 , n23189 , n26535 );
    or g18987 ( n24831 , n17678 , n12065 );
    xnor g18988 ( n6975 , n26595 , n22717 );
    or g18989 ( n26223 , n1272 , n14247 );
    xnor g18990 ( n2536 , n23715 , n19584 );
    and g18991 ( n14333 , n17778 , n17072 );
    xnor g18992 ( n13204 , n16352 , n9943 );
    not g18993 ( n6039 , n1171 );
    and g18994 ( n21889 , n1165 , n18342 );
    nor g18995 ( n1203 , n13172 , n1881 );
    nor g18996 ( n25259 , n14391 , n6293 );
    and g18997 ( n4829 , n24995 , n3866 );
    xnor g18998 ( n19203 , n15636 , n24618 );
    and g18999 ( n25648 , n3364 , n19199 );
    xnor g19000 ( n12627 , n10712 , n26512 );
    xnor g19001 ( n7006 , n2243 , n7658 );
    not g19002 ( n23412 , n22878 );
    xnor g19003 ( n16175 , n24343 , n15767 );
    or g19004 ( n12934 , n3857 , n3761 );
    and g19005 ( n27143 , n20358 , n21379 );
    or g19006 ( n24702 , n14864 , n6667 );
    xnor g19007 ( n13273 , n1828 , n14305 );
    and g19008 ( n12452 , n3009 , n21729 );
    or g19009 ( n2932 , n25507 , n14340 );
    or g19010 ( n25830 , n15015 , n11216 );
    and g19011 ( n220 , n3717 , n19031 );
    and g19012 ( n26966 , n11454 , n19364 );
    not g19013 ( n13237 , n25872 );
    nor g19014 ( n26319 , n13152 , n15053 );
    nor g19015 ( n11020 , n22061 , n26705 );
    nor g19016 ( n7584 , n6265 , n1336 );
    or g19017 ( n16039 , n26322 , n9962 );
    or g19018 ( n5334 , n2511 , n21714 );
    xnor g19019 ( n11947 , n6301 , n6626 );
    and g19020 ( n5478 , n8104 , n899 );
    or g19021 ( n6649 , n3253 , n21021 );
    or g19022 ( n8921 , n25586 , n23525 );
    or g19023 ( n15151 , n12795 , n13315 );
    not g19024 ( n6241 , n2128 );
    xnor g19025 ( n26969 , n26135 , n8119 );
    xnor g19026 ( n13562 , n11323 , n24504 );
    or g19027 ( n10226 , n16669 , n13656 );
    nor g19028 ( n3604 , n23254 , n27008 );
    or g19029 ( n9343 , n12513 , n25568 );
    or g19030 ( n16643 , n13460 , n5156 );
    xnor g19031 ( n9966 , n7353 , n20620 );
    and g19032 ( n25689 , n6107 , n8725 );
    not g19033 ( n17871 , n18075 );
    nor g19034 ( n24471 , n16158 , n10204 );
    or g19035 ( n27180 , n346 , n27138 );
    not g19036 ( n9363 , n22201 );
    xnor g19037 ( n25439 , n14018 , n7735 );
    or g19038 ( n6608 , n4520 , n1694 );
    nor g19039 ( n12320 , n4061 , n9557 );
    or g19040 ( n1276 , n21140 , n10241 );
    and g19041 ( n25651 , n26810 , n12797 );
    or g19042 ( n18042 , n5258 , n10415 );
    not g19043 ( n26711 , n12456 );
    nor g19044 ( n16770 , n20970 , n12961 );
    or g19045 ( n2542 , n1458 , n19494 );
    nor g19046 ( n16192 , n18371 , n21151 );
    or g19047 ( n23518 , n20229 , n1936 );
    and g19048 ( n2255 , n9436 , n3905 );
    xnor g19049 ( n16657 , n2035 , n26823 );
    not g19050 ( n12232 , n23488 );
    xnor g19051 ( n9687 , n21321 , n1750 );
    nor g19052 ( n4577 , n24355 , n11220 );
    xnor g19053 ( n24201 , n5031 , n11926 );
    and g19054 ( n24007 , n4435 , n8533 );
    or g19055 ( n22297 , n14226 , n23217 );
    xnor g19056 ( n1573 , n2276 , n9937 );
    and g19057 ( n6810 , n3982 , n6439 );
    xnor g19058 ( n6525 , n10620 , n10255 );
    and g19059 ( n4732 , n7866 , n13676 );
    xnor g19060 ( n1120 , n25065 , n6500 );
    and g19061 ( n26644 , n7759 , n725 );
    and g19062 ( n4136 , n15363 , n11704 );
    xnor g19063 ( n21750 , n16191 , n11296 );
    or g19064 ( n4825 , n18652 , n11574 );
    or g19065 ( n14197 , n12591 , n24254 );
    xnor g19066 ( n26733 , n22057 , n1523 );
    or g19067 ( n5359 , n123 , n11130 );
    not g19068 ( n17026 , n21998 );
    nor g19069 ( n3416 , n19399 , n13848 );
    nor g19070 ( n19173 , n528 , n17556 );
    xor g19071 ( n22211 , n2481 , n13650 );
    not g19072 ( n11258 , n8165 );
    and g19073 ( n20464 , n26822 , n5475 );
    not g19074 ( n26672 , n10967 );
    or g19075 ( n17772 , n12876 , n3287 );
    nor g19076 ( n12701 , n4335 , n21544 );
    nor g19077 ( n24656 , n17423 , n5101 );
    or g19078 ( n6337 , n4684 , n16942 );
    or g19079 ( n15982 , n4458 , n3415 );
    xnor g19080 ( n1183 , n25285 , n8293 );
    and g19081 ( n6820 , n4844 , n16723 );
    or g19082 ( n17404 , n16901 , n26171 );
    or g19083 ( n11227 , n1458 , n21372 );
    or g19084 ( n13969 , n4904 , n13829 );
    not g19085 ( n8186 , n2978 );
    or g19086 ( n14146 , n12149 , n19045 );
    nor g19087 ( n26475 , n15190 , n182 );
    or g19088 ( n1511 , n1155 , n11688 );
    or g19089 ( n9128 , n26335 , n24099 );
    nor g19090 ( n1833 , n19138 , n21114 );
    or g19091 ( n10529 , n24851 , n2636 );
    xnor g19092 ( n8508 , n6599 , n19608 );
    xnor g19093 ( n3502 , n3254 , n14418 );
    or g19094 ( n22889 , n7561 , n10797 );
    nor g19095 ( n614 , n144 , n18290 );
    xnor g19096 ( n8103 , n14934 , n13881 );
    not g19097 ( n20209 , n16520 );
    nor g19098 ( n7980 , n9376 , n3045 );
    or g19099 ( n17760 , n13638 , n22798 );
    and g19100 ( n14142 , n6252 , n19329 );
    not g19101 ( n6518 , n9961 );
    xnor g19102 ( n19730 , n18578 , n9090 );
    or g19103 ( n8503 , n21432 , n26994 );
    or g19104 ( n13344 , n5773 , n20464 );
    or g19105 ( n24895 , n2339 , n908 );
    or g19106 ( n11573 , n9206 , n24682 );
    or g19107 ( n15990 , n26085 , n1245 );
    and g19108 ( n6156 , n21125 , n926 );
    xnor g19109 ( n2005 , n13904 , n18463 );
    not g19110 ( n20897 , n1339 );
    xnor g19111 ( n5800 , n6657 , n3513 );
    and g19112 ( n25789 , n8603 , n18469 );
    or g19113 ( n23501 , n6855 , n17217 );
    not g19114 ( n9910 , n25120 );
    or g19115 ( n26701 , n17316 , n1893 );
    and g19116 ( n2958 , n4735 , n25811 );
    or g19117 ( n26207 , n6094 , n12877 );
    not g19118 ( n16399 , n24721 );
    nor g19119 ( n5885 , n13297 , n11165 );
    or g19120 ( n3598 , n2063 , n9621 );
    xnor g19121 ( n9111 , n23369 , n26572 );
    or g19122 ( n18062 , n25913 , n10230 );
    not g19123 ( n18991 , n5329 );
    not g19124 ( n25394 , n2429 );
    nor g19125 ( n19558 , n26673 , n19911 );
    xnor g19126 ( n7147 , n21442 , n8891 );
    xnor g19127 ( n24194 , n8469 , n5367 );
    or g19128 ( n5872 , n10758 , n1717 );
    xnor g19129 ( n6826 , n22984 , n25173 );
    and g19130 ( n22612 , n21672 , n19300 );
    xnor g19131 ( n18459 , n11970 , n1757 );
    xnor g19132 ( n11794 , n27104 , n19005 );
    or g19133 ( n14382 , n13494 , n14031 );
    nor g19134 ( n13809 , n5031 , n11926 );
    buf g19135 ( n6352 , n10795 );
    or g19136 ( n8918 , n24823 , n20886 );
    xnor g19137 ( n14464 , n3357 , n20772 );
    xnor g19138 ( n8473 , n17308 , n8751 );
    not g19139 ( n3674 , n23993 );
    or g19140 ( n4193 , n16209 , n15836 );
    or g19141 ( n19451 , n15761 , n11535 );
    and g19142 ( n16636 , n25728 , n11629 );
    or g19143 ( n10889 , n18504 , n17483 );
    and g19144 ( n25372 , n24657 , n114 );
    and g19145 ( n21503 , n8914 , n4666 );
    xnor g19146 ( n26722 , n4 , n23544 );
    xnor g19147 ( n4499 , n7196 , n1778 );
    and g19148 ( n20643 , n1195 , n21412 );
    and g19149 ( n13143 , n4274 , n20177 );
    or g19150 ( n12497 , n10145 , n7846 );
    and g19151 ( n16190 , n10995 , n1082 );
    xnor g19152 ( n15991 , n15372 , n17857 );
    or g19153 ( n21651 , n18510 , n9888 );
    xnor g19154 ( n7077 , n12702 , n18105 );
    xnor g19155 ( n12766 , n8193 , n9914 );
    xnor g19156 ( n6233 , n23356 , n11129 );
    or g19157 ( n19745 , n16720 , n23510 );
    xnor g19158 ( n3218 , n17789 , n10915 );
    and g19159 ( n13417 , n25291 , n7061 );
    xnor g19160 ( n23433 , n22210 , n21149 );
    not g19161 ( n2453 , n12875 );
    nor g19162 ( n3290 , n22554 , n26318 );
    and g19163 ( n5335 , n9040 , n26799 );
    and g19164 ( n1758 , n26354 , n11873 );
    xnor g19165 ( n1522 , n16266 , n22458 );
    not g19166 ( n13925 , n11335 );
    and g19167 ( n25609 , n22920 , n11715 );
    nor g19168 ( n8989 , n19890 , n6449 );
    xnor g19169 ( n16909 , n11486 , n18409 );
    nor g19170 ( n5356 , n16633 , n22793 );
    xnor g19171 ( n14418 , n728 , n12029 );
    and g19172 ( n1978 , n24358 , n20951 );
    xnor g19173 ( n13452 , n5512 , n16217 );
    xnor g19174 ( n9072 , n7755 , n21097 );
    xnor g19175 ( n24376 , n6255 , n6658 );
    and g19176 ( n7741 , n2160 , n27095 );
    nor g19177 ( n4711 , n16399 , n11603 );
    and g19178 ( n16131 , n25207 , n1101 );
    nor g19179 ( n26094 , n19634 , n19228 );
    and g19180 ( n12332 , n3899 , n15263 );
    not g19181 ( n21506 , n10472 );
    not g19182 ( n265 , n501 );
    nor g19183 ( n12046 , n1314 , n20967 );
    xnor g19184 ( n24160 , n7603 , n15111 );
    xnor g19185 ( n19916 , n18402 , n21816 );
    or g19186 ( n3368 , n12640 , n18274 );
    xnor g19187 ( n8317 , n2739 , n4865 );
    or g19188 ( n22129 , n10757 , n13811 );
    or g19189 ( n4465 , n21598 , n10161 );
    nor g19190 ( n21292 , n5559 , n7697 );
    xnor g19191 ( n23882 , n9355 , n3844 );
    xnor g19192 ( n7658 , n987 , n626 );
    or g19193 ( n8814 , n17514 , n20960 );
    or g19194 ( n16240 , n26625 , n14230 );
    not g19195 ( n19295 , n1167 );
    not g19196 ( n17164 , n23326 );
    xnor g19197 ( n23295 , n6631 , n12209 );
    xnor g19198 ( n11109 , n16401 , n7861 );
    not g19199 ( n23016 , n24202 );
    xnor g19200 ( n15488 , n19978 , n4240 );
    xnor g19201 ( n10359 , n2813 , n23272 );
    or g19202 ( n17477 , n18057 , n9362 );
    or g19203 ( n23403 , n20638 , n5296 );
    nor g19204 ( n11443 , n9215 , n15616 );
    and g19205 ( n12172 , n4117 , n14188 );
    not g19206 ( n19758 , n4368 );
    and g19207 ( n26886 , n19541 , n14182 );
    or g19208 ( n4292 , n4543 , n18860 );
    xnor g19209 ( n21718 , n1798 , n1742 );
    xnor g19210 ( n13048 , n394 , n18005 );
    or g19211 ( n21594 , n1660 , n23634 );
    not g19212 ( n10831 , n2651 );
    not g19213 ( n16928 , n9700 );
    xnor g19214 ( n18961 , n14514 , n2279 );
    or g19215 ( n7121 , n7876 , n11479 );
    and g19216 ( n6953 , n24768 , n1019 );
    or g19217 ( n25417 , n17365 , n6000 );
    not g19218 ( n24484 , n12291 );
    or g19219 ( n17525 , n604 , n13318 );
    not g19220 ( n7213 , n13665 );
    and g19221 ( n3428 , n3260 , n20512 );
    nor g19222 ( n23758 , n15440 , n3147 );
    or g19223 ( n7509 , n6206 , n11529 );
    xnor g19224 ( n9971 , n5754 , n27032 );
    and g19225 ( n5380 , n3788 , n5920 );
    and g19226 ( n18212 , n18451 , n27034 );
    and g19227 ( n17821 , n6103 , n15211 );
    nor g19228 ( n10983 , n10184 , n12366 );
    and g19229 ( n15256 , n5519 , n20934 );
    and g19230 ( n1159 , n17970 , n15250 );
    or g19231 ( n627 , n7472 , n3288 );
    and g19232 ( n10070 , n15202 , n17124 );
    xnor g19233 ( n25555 , n3032 , n11911 );
    or g19234 ( n16661 , n22087 , n4824 );
    nor g19235 ( n16931 , n10989 , n19017 );
    or g19236 ( n26434 , n7893 , n20205 );
    and g19237 ( n26783 , n13088 , n18987 );
    xnor g19238 ( n16140 , n25974 , n8399 );
    or g19239 ( n18299 , n20684 , n16518 );
    xnor g19240 ( n21444 , n8190 , n19714 );
    and g19241 ( n18941 , n25642 , n1133 );
    nor g19242 ( n240 , n1205 , n8568 );
    nor g19243 ( n3519 , n9851 , n10389 );
    and g19244 ( n15227 , n24220 , n14191 );
    or g19245 ( n8726 , n14766 , n8808 );
    nor g19246 ( n5766 , n21749 , n919 );
    xnor g19247 ( n14277 , n10526 , n8665 );
    not g19248 ( n17173 , n10405 );
    nor g19249 ( n2777 , n2780 , n4665 );
    or g19250 ( n24583 , n7818 , n18139 );
    or g19251 ( n1763 , n18119 , n23827 );
    or g19252 ( n16783 , n19175 , n12343 );
    or g19253 ( n4960 , n15820 , n21824 );
    or g19254 ( n5573 , n13920 , n5839 );
    and g19255 ( n26587 , n24384 , n10528 );
    xnor g19256 ( n1695 , n4194 , n14643 );
    or g19257 ( n22796 , n435 , n14494 );
    nor g19258 ( n15317 , n14386 , n24051 );
    and g19259 ( n9449 , n6877 , n17155 );
    or g19260 ( n5153 , n2797 , n17742 );
    not g19261 ( n7639 , n8876 );
    or g19262 ( n2824 , n23772 , n23106 );
    xnor g19263 ( n24896 , n1038 , n15342 );
    nor g19264 ( n8998 , n24202 , n9595 );
    and g19265 ( n6301 , n6317 , n2670 );
    nor g19266 ( n13563 , n5516 , n24085 );
    or g19267 ( n16033 , n23211 , n24665 );
    or g19268 ( n8812 , n8865 , n12946 );
    or g19269 ( n14806 , n21924 , n9476 );
    and g19270 ( n16728 , n3591 , n3963 );
    xnor g19271 ( n11196 , n3280 , n2038 );
    not g19272 ( n11989 , n10051 );
    or g19273 ( n15592 , n9880 , n13714 );
    xnor g19274 ( n2468 , n7107 , n26582 );
    and g19275 ( n23409 , n17356 , n11716 );
    nor g19276 ( n8576 , n8097 , n17210 );
    xnor g19277 ( n13112 , n2068 , n12219 );
    and g19278 ( n24496 , n12210 , n17085 );
    or g19279 ( n451 , n19557 , n9040 );
    or g19280 ( n2720 , n11637 , n27058 );
    or g19281 ( n5965 , n16751 , n27082 );
    xnor g19282 ( n9321 , n14996 , n7678 );
    not g19283 ( n15940 , n9318 );
    xnor g19284 ( n245 , n8399 , n13708 );
    xnor g19285 ( n60 , n16364 , n7680 );
    xnor g19286 ( n19401 , n15708 , n16969 );
    not g19287 ( n19868 , n1304 );
    nor g19288 ( n24899 , n3694 , n14514 );
    xnor g19289 ( n12731 , n24112 , n15077 );
    and g19290 ( n2200 , n26014 , n14144 );
    xnor g19291 ( n984 , n3321 , n14888 );
    xnor g19292 ( n17640 , n1075 , n24016 );
    xnor g19293 ( n21643 , n95 , n3851 );
    not g19294 ( n25835 , n9362 );
    xnor g19295 ( n8596 , n25435 , n18 );
    or g19296 ( n19890 , n9356 , n17373 );
    xnor g19297 ( n13039 , n11253 , n9208 );
    xnor g19298 ( n11565 , n20751 , n24593 );
    xnor g19299 ( n16196 , n23154 , n13788 );
    and g19300 ( n16144 , n2088 , n6414 );
    not g19301 ( n22104 , n10004 );
    nor g19302 ( n19716 , n8067 , n3319 );
    not g19303 ( n11228 , n12573 );
    or g19304 ( n3184 , n4070 , n15479 );
    or g19305 ( n10693 , n12991 , n24700 );
    xnor g19306 ( n20480 , n18759 , n16244 );
    xnor g19307 ( n19940 , n13101 , n19817 );
    xnor g19308 ( n13034 , n3944 , n941 );
    not g19309 ( n25330 , n22138 );
    not g19310 ( n910 , n3016 );
    nor g19311 ( n18612 , n7769 , n25316 );
    and g19312 ( n13103 , n25940 , n22325 );
    or g19313 ( n121 , n4058 , n19534 );
    nor g19314 ( n8580 , n15546 , n5629 );
    xnor g19315 ( n4623 , n20597 , n20055 );
    nor g19316 ( n6664 , n5715 , n22918 );
    xnor g19317 ( n13139 , n20075 , n14386 );
    and g19318 ( n9446 , n3348 , n202 );
    xnor g19319 ( n9915 , n1509 , n2517 );
    xnor g19320 ( n23450 , n6865 , n16378 );
    xnor g19321 ( n21315 , n18797 , n25799 );
    or g19322 ( n20174 , n15864 , n1455 );
    or g19323 ( n18819 , n20752 , n5458 );
    and g19324 ( n4035 , n13775 , n8389 );
    or g19325 ( n6964 , n4926 , n4517 );
    or g19326 ( n6986 , n19650 , n21616 );
    and g19327 ( n12310 , n16237 , n23003 );
    xnor g19328 ( n5513 , n13490 , n12446 );
    and g19329 ( n19759 , n2038 , n2574 );
    and g19330 ( n18297 , n6393 , n2028 );
    xnor g19331 ( n18187 , n15770 , n22881 );
    and g19332 ( n24799 , n21634 , n16007 );
    or g19333 ( n7015 , n11978 , n1194 );
    or g19334 ( n9140 , n9681 , n16475 );
    not g19335 ( n26962 , n7634 );
    not g19336 ( n26211 , n7049 );
    not g19337 ( n7252 , n5188 );
    not g19338 ( n15998 , n2696 );
    xnor g19339 ( n765 , n9793 , n10250 );
    and g19340 ( n16489 , n267 , n16317 );
    xnor g19341 ( n23287 , n24948 , n10514 );
    xnor g19342 ( n13328 , n7749 , n8681 );
    not g19343 ( n13897 , n17035 );
    not g19344 ( n24925 , n287 );
    xnor g19345 ( n7872 , n13633 , n19039 );
    or g19346 ( n15099 , n25844 , n15552 );
    and g19347 ( n15124 , n1330 , n14077 );
    or g19348 ( n7545 , n22781 , n20394 );
    or g19349 ( n12568 , n13481 , n11238 );
    xnor g19350 ( n10272 , n14510 , n16988 );
    and g19351 ( n3042 , n6920 , n1286 );
    xnor g19352 ( n6939 , n15903 , n13468 );
    not g19353 ( n2780 , n8309 );
    and g19354 ( n19237 , n10171 , n10348 );
    xnor g19355 ( n2755 , n11207 , n22358 );
    xnor g19356 ( n4713 , n2420 , n22201 );
    or g19357 ( n5248 , n9899 , n26952 );
    and g19358 ( n4900 , n19894 , n22517 );
    or g19359 ( n2006 , n9600 , n17870 );
    not g19360 ( n25982 , n7707 );
    and g19361 ( n5270 , n15554 , n66 );
    or g19362 ( n11046 , n24044 , n22379 );
    xnor g19363 ( n19244 , n19654 , n21642 );
    not g19364 ( n26524 , n22898 );
    nor g19365 ( n12038 , n13089 , n3625 );
    or g19366 ( n25493 , n13428 , n1368 );
    not g19367 ( n17869 , n914 );
    and g19368 ( n17633 , n2814 , n7651 );
    and g19369 ( n5528 , n21051 , n16035 );
    nor g19370 ( n27003 , n22874 , n9492 );
    xnor g19371 ( n110 , n333 , n15268 );
    not g19372 ( n13944 , n10479 );
    or g19373 ( n3322 , n17848 , n5863 );
    nor g19374 ( n24267 , n20378 , n9493 );
    not g19375 ( n8925 , n11254 );
    or g19376 ( n15310 , n12894 , n25646 );
    or g19377 ( n12611 , n25450 , n2128 );
    xnor g19378 ( n8427 , n16555 , n20040 );
    and g19379 ( n14208 , n13159 , n15924 );
    or g19380 ( n12492 , n1190 , n14721 );
    or g19381 ( n8200 , n9496 , n22515 );
    xnor g19382 ( n27019 , n10110 , n22669 );
    xnor g19383 ( n17130 , n23507 , n16871 );
    nor g19384 ( n19139 , n1163 , n2675 );
    or g19385 ( n26527 , n17908 , n21550 );
    xnor g19386 ( n18720 , n26637 , n19866 );
    and g19387 ( n24874 , n16372 , n10845 );
    nor g19388 ( n7035 , n19789 , n21226 );
    and g19389 ( n24655 , n13059 , n22913 );
    xnor g19390 ( n21956 , n23793 , n18 );
    nor g19391 ( n19705 , n14444 , n1780 );
    xnor g19392 ( n15654 , n7428 , n19107 );
    xnor g19393 ( n1426 , n21079 , n369 );
    or g19394 ( n25300 , n16770 , n12032 );
    not g19395 ( n9113 , n27141 );
    and g19396 ( n8894 , n6804 , n11768 );
    or g19397 ( n8548 , n18666 , n26575 );
    buf g19398 ( n10023 , n23310 );
    not g19399 ( n25122 , n7335 );
    nor g19400 ( n25844 , n14736 , n22139 );
    xnor g19401 ( n14797 , n17122 , n23383 );
    xnor g19402 ( n17765 , n874 , n16949 );
    and g19403 ( n19411 , n22320 , n6563 );
    or g19404 ( n16579 , n9805 , n19055 );
    not g19405 ( n20437 , n18416 );
    buf g19406 ( n21547 , n17152 );
    not g19407 ( n1421 , n10039 );
    xnor g19408 ( n3131 , n6072 , n11706 );
    xnor g19409 ( n23833 , n8712 , n26620 );
    and g19410 ( n2984 , n18074 , n26476 );
    and g19411 ( n22269 , n23000 , n24908 );
    not g19412 ( n3378 , n2965 );
    or g19413 ( n23404 , n1250 , n8413 );
    xnor g19414 ( n20626 , n8672 , n26224 );
    xnor g19415 ( n2869 , n21948 , n20840 );
    not g19416 ( n4282 , n21908 );
    not g19417 ( n21060 , n14482 );
    xnor g19418 ( n26651 , n20700 , n932 );
    nor g19419 ( n14988 , n18295 , n25974 );
    and g19420 ( n10351 , n23141 , n3238 );
    not g19421 ( n14555 , n25601 );
    xnor g19422 ( n2963 , n23895 , n5101 );
    or g19423 ( n16606 , n19731 , n23993 );
    and g19424 ( n1411 , n18379 , n21285 );
    xnor g19425 ( n5880 , n24624 , n23517 );
    or g19426 ( n18457 , n15711 , n27124 );
    or g19427 ( n22146 , n9373 , n7765 );
    xnor g19428 ( n4153 , n18640 , n3814 );
    or g19429 ( n1551 , n9825 , n18612 );
    xnor g19430 ( n14728 , n9751 , n17353 );
    xnor g19431 ( n24919 , n26083 , n22734 );
    or g19432 ( n17127 , n1937 , n1310 );
    or g19433 ( n26844 , n7421 , n20044 );
    not g19434 ( n17511 , n3509 );
    or g19435 ( n17457 , n25156 , n2784 );
    or g19436 ( n24943 , n6369 , n527 );
    or g19437 ( n19136 , n4820 , n7745 );
    or g19438 ( n15068 , n2976 , n10904 );
    and g19439 ( n20593 , n17453 , n26783 );
    and g19440 ( n21875 , n17464 , n4536 );
    nor g19441 ( n1635 , n13422 , n685 );
    nor g19442 ( n12800 , n24327 , n2768 );
    and g19443 ( n17986 , n10175 , n22129 );
    nor g19444 ( n15697 , n6750 , n63 );
    or g19445 ( n276 , n3062 , n18047 );
    or g19446 ( n22057 , n13756 , n7244 );
    xnor g19447 ( n1001 , n4625 , n20835 );
    nor g19448 ( n13386 , n19515 , n10651 );
    not g19449 ( n2995 , n13475 );
    xnor g19450 ( n6834 , n5488 , n7149 );
    or g19451 ( n9255 , n13195 , n12217 );
    xnor g19452 ( n20546 , n20323 , n8564 );
    xnor g19453 ( n23778 , n23353 , n12702 );
    and g19454 ( n6490 , n8325 , n13866 );
    or g19455 ( n7896 , n25058 , n15487 );
    not g19456 ( n26658 , n10053 );
    or g19457 ( n2701 , n7681 , n2338 );
    nor g19458 ( n25922 , n16795 , n17498 );
    nor g19459 ( n14861 , n22281 , n18157 );
    not g19460 ( n10720 , n1685 );
    xnor g19461 ( n20354 , n1478 , n12731 );
    and g19462 ( n7637 , n26121 , n1409 );
    and g19463 ( n18129 , n20228 , n8717 );
    xnor g19464 ( n8765 , n7430 , n18218 );
    and g19465 ( n13833 , n23887 , n18989 );
    xnor g19466 ( n25576 , n23180 , n18690 );
    or g19467 ( n18324 , n23097 , n7399 );
    or g19468 ( n21648 , n9407 , n9109 );
    xnor g19469 ( n24512 , n2492 , n22175 );
    xnor g19470 ( n14070 , n9108 , n6877 );
    nor g19471 ( n21128 , n21489 , n11062 );
    xnor g19472 ( n15960 , n18 , n22843 );
    and g19473 ( n21985 , n9176 , n4907 );
    xnor g19474 ( n6634 , n9029 , n22711 );
    and g19475 ( n4921 , n15785 , n16953 );
    nor g19476 ( n21369 , n6187 , n25641 );
    not g19477 ( n26056 , n14125 );
    nor g19478 ( n9985 , n20151 , n19042 );
    nor g19479 ( n9834 , n14472 , n26821 );
    nor g19480 ( n1039 , n16396 , n8399 );
    xnor g19481 ( n5857 , n21101 , n16722 );
    nor g19482 ( n22887 , n13941 , n6025 );
    xnor g19483 ( n8874 , n9003 , n6369 );
    xnor g19484 ( n19190 , n10919 , n8943 );
    or g19485 ( n33 , n1557 , n5892 );
    and g19486 ( n4348 , n23553 , n12643 );
    not g19487 ( n24043 , n5733 );
    xnor g19488 ( n5392 , n3809 , n8719 );
    and g19489 ( n4485 , n25242 , n8868 );
    and g19490 ( n11411 , n23223 , n13785 );
    or g19491 ( n831 , n20638 , n22986 );
    and g19492 ( n3533 , n21201 , n26242 );
    xnor g19493 ( n15764 , n19990 , n18313 );
    or g19494 ( n8400 , n25424 , n14432 );
    or g19495 ( n21463 , n25510 , n4504 );
    or g19496 ( n2823 , n16512 , n11340 );
    xnor g19497 ( n25322 , n16334 , n21784 );
    xnor g19498 ( n24975 , n17835 , n7026 );
    nor g19499 ( n14864 , n20470 , n3366 );
    xnor g19500 ( n6471 , n17498 , n24989 );
    xnor g19501 ( n8911 , n27047 , n23698 );
    and g19502 ( n16634 , n3959 , n25917 );
    xnor g19503 ( n9500 , n11802 , n15975 );
    and g19504 ( n13182 , n17916 , n21624 );
    xnor g19505 ( n18705 , n19302 , n18875 );
    not g19506 ( n26350 , n2954 );
    and g19507 ( n17489 , n23998 , n17043 );
    or g19508 ( n24429 , n11865 , n10876 );
    xnor g19509 ( n9011 , n246 , n17401 );
    or g19510 ( n15968 , n18929 , n22036 );
    xnor g19511 ( n27072 , n25720 , n19834 );
    and g19512 ( n4458 , n3199 , n3373 );
    xnor g19513 ( n2881 , n13958 , n15586 );
    nor g19514 ( n5069 , n2470 , n10496 );
    xnor g19515 ( n17012 , n14886 , n17639 );
    xnor g19516 ( n26439 , n10128 , n16340 );
    xnor g19517 ( n3234 , n12508 , n22850 );
    xnor g19518 ( n7735 , n12379 , n8067 );
    or g19519 ( n17239 , n19033 , n20724 );
    not g19520 ( n10788 , n3968 );
    and g19521 ( n21550 , n18879 , n25011 );
    and g19522 ( n8057 , n23579 , n26223 );
    buf g19523 ( n19227 , n4956 );
    nor g19524 ( n9080 , n16359 , n26149 );
    and g19525 ( n5207 , n25248 , n13931 );
    or g19526 ( n13086 , n13596 , n10649 );
    nor g19527 ( n7623 , n26717 , n7963 );
    xnor g19528 ( n14636 , n1548 , n18661 );
    or g19529 ( n1872 , n14684 , n21952 );
    and g19530 ( n4018 , n9664 , n20122 );
    xnor g19531 ( n22607 , n13583 , n2963 );
    xnor g19532 ( n14003 , n24061 , n128 );
    or g19533 ( n21345 , n26145 , n20360 );
    xnor g19534 ( n10929 , n13668 , n20923 );
    xnor g19535 ( n22627 , n26023 , n4692 );
    xnor g19536 ( n23048 , n14770 , n15234 );
    nor g19537 ( n3594 , n3968 , n13980 );
    or g19538 ( n27174 , n19862 , n16722 );
    or g19539 ( n22719 , n3739 , n15892 );
    or g19540 ( n14820 , n65 , n22464 );
    and g19541 ( n10795 , n12779 , n18329 );
    xnor g19542 ( n8070 , n17221 , n6491 );
    or g19543 ( n24434 , n19361 , n20060 );
    not g19544 ( n15269 , n23784 );
    and g19545 ( n1643 , n725 , n24804 );
    nor g19546 ( n21865 , n19926 , n21295 );
    or g19547 ( n12853 , n19869 , n20092 );
    or g19548 ( n748 , n4913 , n13489 );
    xnor g19549 ( n1851 , n6486 , n15077 );
    xnor g19550 ( n20447 , n11589 , n4518 );
    not g19551 ( n16052 , n21405 );
    xnor g19552 ( n19793 , n12657 , n23697 );
    not g19553 ( n13164 , n4207 );
    or g19554 ( n270 , n20249 , n9736 );
    xnor g19555 ( n19224 , n19754 , n20611 );
    and g19556 ( n5192 , n17264 , n9128 );
    and g19557 ( n10945 , n16474 , n15491 );
    or g19558 ( n14098 , n14654 , n18519 );
    or g19559 ( n1211 , n5055 , n1318 );
    and g19560 ( n19620 , n23169 , n2823 );
    xnor g19561 ( n23883 , n2097 , n2869 );
    and g19562 ( n24414 , n19144 , n5496 );
    and g19563 ( n7530 , n25745 , n5291 );
    or g19564 ( n340 , n19003 , n24475 );
    xnor g19565 ( n4403 , n12088 , n16029 );
    and g19566 ( n5659 , n6796 , n1032 );
    not g19567 ( n21672 , n18672 );
    or g19568 ( n25702 , n19264 , n22088 );
    or g19569 ( n6663 , n24098 , n23250 );
    and g19570 ( n26017 , n16010 , n7984 );
    xnor g19571 ( n2700 , n3164 , n268 );
    not g19572 ( n23098 , n7407 );
    xnor g19573 ( n17756 , n18191 , n21993 );
    or g19574 ( n2081 , n13420 , n19337 );
    xnor g19575 ( n16768 , n16482 , n13074 );
    xnor g19576 ( n3986 , n26251 , n1630 );
    and g19577 ( n21766 , n1742 , n25394 );
    not g19578 ( n1624 , n7755 );
    and g19579 ( n25096 , n17333 , n19247 );
    and g19580 ( n19840 , n14963 , n19112 );
    xnor g19581 ( n18576 , n14935 , n9256 );
    and g19582 ( n16771 , n1319 , n6864 );
    or g19583 ( n21653 , n7215 , n23493 );
    or g19584 ( n2670 , n10707 , n6535 );
    or g19585 ( n25709 , n1812 , n15172 );
    xnor g19586 ( n9077 , n14652 , n9742 );
    not g19587 ( n4077 , n6107 );
    not g19588 ( n22222 , n1429 );
    not g19589 ( n9600 , n10593 );
    and g19590 ( n13588 , n10138 , n10105 );
    nor g19591 ( n888 , n22824 , n23686 );
    xnor g19592 ( n26694 , n24868 , n13044 );
    and g19593 ( n16523 , n18764 , n14175 );
    and g19594 ( n3051 , n23094 , n24658 );
    and g19595 ( n20861 , n6386 , n3501 );
    nor g19596 ( n13910 , n18125 , n15131 );
    xnor g19597 ( n25465 , n19766 , n11557 );
    not g19598 ( n27065 , n13476 );
    nor g19599 ( n23808 , n8431 , n21547 );
    nor g19600 ( n2613 , n26007 , n5621 );
    and g19601 ( n10254 , n22071 , n26291 );
    or g19602 ( n27166 , n8259 , n16551 );
    and g19603 ( n20347 , n11645 , n17807 );
    or g19604 ( n3255 , n2048 , n2607 );
    or g19605 ( n25859 , n23030 , n4333 );
    and g19606 ( n21737 , n25469 , n20631 );
    and g19607 ( n316 , n11219 , n3088 );
    or g19608 ( n11358 , n24012 , n12109 );
    or g19609 ( n160 , n26408 , n1186 );
    xnor g19610 ( n646 , n14987 , n12959 );
    or g19611 ( n18629 , n16474 , n18302 );
    nor g19612 ( n1280 , n20667 , n26066 );
    or g19613 ( n3374 , n3633 , n23389 );
    and g19614 ( n24238 , n9255 , n7513 );
    and g19615 ( n6469 , n5257 , n6876 );
    or g19616 ( n10583 , n16159 , n22378 );
    xnor g19617 ( n27194 , n6114 , n1671 );
    or g19618 ( n3163 , n17456 , n25653 );
    not g19619 ( n20655 , n16907 );
    not g19620 ( n9964 , n1451 );
    xnor g19621 ( n13611 , n21842 , n3828 );
    xnor g19622 ( n13940 , n15780 , n2387 );
    xnor g19623 ( n25966 , n25197 , n23498 );
    and g19624 ( n25273 , n6554 , n25060 );
    or g19625 ( n11526 , n15998 , n5142 );
    xnor g19626 ( n9622 , n21618 , n26337 );
    xnor g19627 ( n8573 , n24736 , n14603 );
    or g19628 ( n25895 , n5245 , n11259 );
    nor g19629 ( n4398 , n7249 , n10441 );
    and g19630 ( n8236 , n3254 , n2738 );
    not g19631 ( n12968 , n16264 );
    xnor g19632 ( n1840 , n18634 , n20470 );
    xnor g19633 ( n13560 , n1694 , n9909 );
    not g19634 ( n4721 , n6105 );
    not g19635 ( n24559 , n22314 );
    or g19636 ( n24984 , n20325 , n5515 );
    xnor g19637 ( n17236 , n22263 , n9581 );
    nor g19638 ( n24005 , n665 , n17599 );
    xor g19639 ( n3602 , n7973 , n8381 );
    xnor g19640 ( n1007 , n22349 , n13493 );
    and g19641 ( n3857 , n16054 , n17600 );
    or g19642 ( n14246 , n17598 , n17926 );
    xnor g19643 ( n7157 , n18255 , n23369 );
    and g19644 ( n25594 , n21554 , n25158 );
    xnor g19645 ( n26765 , n11098 , n13912 );
    nor g19646 ( n3685 , n12048 , n8210 );
    nor g19647 ( n17877 , n9960 , n21482 );
    or g19648 ( n6163 , n536 , n4848 );
    and g19649 ( n4512 , n12006 , n21806 );
    not g19650 ( n18510 , n11314 );
    not g19651 ( n23710 , n8206 );
    or g19652 ( n12397 , n3153 , n23459 );
    xnor g19653 ( n266 , n21591 , n13612 );
    or g19654 ( n16919 , n20728 , n11483 );
    or g19655 ( n6627 , n14514 , n3848 );
    or g19656 ( n11436 , n26184 , n316 );
    nor g19657 ( n17293 , n15265 , n12152 );
    xnor g19658 ( n2356 , n21014 , n8958 );
    and g19659 ( n15858 , n109 , n6503 );
    xnor g19660 ( n10039 , n17979 , n22659 );
    or g19661 ( n7839 , n10969 , n16470 );
    or g19662 ( n2554 , n5586 , n19522 );
    or g19663 ( n9258 , n524 , n25069 );
    or g19664 ( n23391 , n25558 , n3414 );
    nor g19665 ( n18353 , n24312 , n10847 );
    and g19666 ( n14083 , n19043 , n1087 );
    xnor g19667 ( n9581 , n17953 , n12971 );
    and g19668 ( n10074 , n340 , n700 );
    not g19669 ( n14875 , n3019 );
    not g19670 ( n12249 , n280 );
    and g19671 ( n4895 , n13081 , n18729 );
    xnor g19672 ( n21828 , n13449 , n6381 );
    not g19673 ( n21796 , n15126 );
    not g19674 ( n25036 , n16173 );
    xnor g19675 ( n13412 , n7546 , n25846 );
    xnor g19676 ( n15931 , n15710 , n23309 );
    nor g19677 ( n23202 , n20920 , n26851 );
    or g19678 ( n6958 , n27104 , n15618 );
    or g19679 ( n2592 , n3921 , n1894 );
    not g19680 ( n850 , n12100 );
    or g19681 ( n18747 , n13889 , n12123 );
    and g19682 ( n3696 , n1438 , n11527 );
    and g19683 ( n17701 , n17925 , n2270 );
    and g19684 ( n3885 , n26683 , n16087 );
    or g19685 ( n21454 , n7455 , n27200 );
    or g19686 ( n18246 , n12277 , n10454 );
    xnor g19687 ( n9793 , n25683 , n15014 );
    or g19688 ( n19538 , n26475 , n25364 );
    and g19689 ( n4643 , n23126 , n10781 );
    xnor g19690 ( n6850 , n8006 , n15289 );
    xnor g19691 ( n15281 , n22492 , n9372 );
    xnor g19692 ( n12860 , n20876 , n24335 );
    not g19693 ( n13448 , n21150 );
    or g19694 ( n22174 , n20973 , n13539 );
    xnor g19695 ( n5053 , n16544 , n2160 );
    or g19696 ( n17492 , n6026 , n8531 );
    or g19697 ( n4678 , n11303 , n5948 );
    or g19698 ( n22707 , n9378 , n10833 );
    nor g19699 ( n10365 , n24897 , n24040 );
    not g19700 ( n19549 , n25602 );
    and g19701 ( n23510 , n13586 , n26950 );
    xnor g19702 ( n188 , n26522 , n1553 );
    xnor g19703 ( n3963 , n5644 , n827 );
    nor g19704 ( n1059 , n25794 , n6944 );
    not g19705 ( n3203 , n13195 );
    or g19706 ( n16259 , n22727 , n17411 );
    or g19707 ( n6804 , n7041 , n1924 );
    xnor g19708 ( n4925 , n21466 , n8598 );
    not g19709 ( n7320 , n13914 );
    or g19710 ( n25761 , n15888 , n1398 );
    and g19711 ( n22212 , n2903 , n27041 );
    or g19712 ( n21526 , n23337 , n16213 );
    or g19713 ( n4655 , n3780 , n26311 );
    or g19714 ( n21925 , n13443 , n10739 );
    or g19715 ( n2847 , n8741 , n23919 );
    or g19716 ( n6546 , n15274 , n16514 );
    xnor g19717 ( n14004 , n25789 , n2198 );
    xnor g19718 ( n3346 , n25275 , n18271 );
    and g19719 ( n24244 , n15137 , n1305 );
    and g19720 ( n21738 , n7956 , n4563 );
    xnor g19721 ( n1632 , n7561 , n8714 );
    or g19722 ( n4592 , n11669 , n26523 );
    xnor g19723 ( n22858 , n4106 , n22398 );
    nor g19724 ( n20881 , n2780 , n7910 );
    xnor g19725 ( n2942 , n8195 , n23757 );
    not g19726 ( n15041 , n26109 );
    xnor g19727 ( n22939 , n15067 , n18075 );
    xnor g19728 ( n16230 , n27202 , n24482 );
    xnor g19729 ( n7809 , n1546 , n21532 );
    and g19730 ( n18293 , n21213 , n4685 );
    or g19731 ( n4573 , n21659 , n24914 );
    not g19732 ( n15217 , n17250 );
    xnor g19733 ( n3679 , n11108 , n16794 );
    and g19734 ( n20942 , n2863 , n21043 );
    xnor g19735 ( n17309 , n13286 , n14341 );
    not g19736 ( n32 , n2127 );
    or g19737 ( n13402 , n6764 , n2088 );
    and g19738 ( n15732 , n9289 , n23152 );
    xnor g19739 ( n24047 , n22139 , n10343 );
    or g19740 ( n19669 , n24671 , n10431 );
    xnor g19741 ( n4758 , n21839 , n22270 );
    nor g19742 ( n7662 , n8492 , n8695 );
    xnor g19743 ( n15285 , n12049 , n9392 );
    and g19744 ( n5473 , n14325 , n20063 );
    nor g19745 ( n13704 , n9259 , n6456 );
    or g19746 ( n12506 , n22230 , n20005 );
    and g19747 ( n14161 , n23721 , n15849 );
    not g19748 ( n23805 , n13277 );
    xnor g19749 ( n19747 , n27102 , n20250 );
    xnor g19750 ( n17804 , n17029 , n1416 );
    not g19751 ( n25246 , n24161 );
    xnor g19752 ( n27146 , n16437 , n1129 );
    nor g19753 ( n7551 , n9908 , n4576 );
    xnor g19754 ( n22113 , n2810 , n4929 );
    xnor g19755 ( n23192 , n18290 , n23529 );
    or g19756 ( n8939 , n1178 , n1148 );
    and g19757 ( n15046 , n13312 , n21706 );
    not g19758 ( n962 , n1022 );
    and g19759 ( n5858 , n2752 , n3678 );
    nor g19760 ( n10716 , n349 , n12456 );
    or g19761 ( n2664 , n6509 , n6080 );
    and g19762 ( n1504 , n22901 , n16861 );
    nor g19763 ( n3996 , n1205 , n13319 );
    or g19764 ( n15899 , n22604 , n2093 );
    and g19765 ( n5233 , n1186 , n12317 );
    nor g19766 ( n968 , n10799 , n19326 );
    not g19767 ( n2230 , n8381 );
    xnor g19768 ( n12230 , n18575 , n10430 );
    xnor g19769 ( n19792 , n13232 , n5507 );
    or g19770 ( n24725 , n13339 , n13178 );
    nor g19771 ( n1843 , n14265 , n15906 );
    xnor g19772 ( n10537 , n593 , n20036 );
    not g19773 ( n8094 , n342 );
    nor g19774 ( n3385 , n5095 , n24134 );
    and g19775 ( n10727 , n25183 , n26531 );
    and g19776 ( n459 , n17946 , n26697 );
    not g19777 ( n26477 , n3196 );
    xnor g19778 ( n26940 , n16544 , n4319 );
    xnor g19779 ( n7884 , n14956 , n13622 );
    or g19780 ( n11385 , n15265 , n9911 );
    xnor g19781 ( n19560 , n4921 , n15649 );
    and g19782 ( n1817 , n12974 , n4332 );
    buf g19783 ( n8875 , n19162 );
    or g19784 ( n19167 , n15522 , n21852 );
    or g19785 ( n16018 , n18228 , n23651 );
    xnor g19786 ( n11018 , n25898 , n21674 );
    xnor g19787 ( n8358 , n17424 , n2370 );
    xnor g19788 ( n12011 , n16114 , n12195 );
    nor g19789 ( n11953 , n4514 , n21698 );
    not g19790 ( n14652 , n2020 );
    or g19791 ( n11922 , n25178 , n9150 );
    or g19792 ( n8919 , n2091 , n1940 );
    and g19793 ( n25671 , n16386 , n5739 );
    or g19794 ( n3246 , n5899 , n16567 );
    xnor g19795 ( n16099 , n24949 , n6199 );
    not g19796 ( n14615 , n19683 );
    nor g19797 ( n23603 , n8331 , n26216 );
    not g19798 ( n6857 , n9851 );
    or g19799 ( n17665 , n20249 , n26292 );
    not g19800 ( n1749 , n9701 );
    xnor g19801 ( n259 , n20549 , n10551 );
    xnor g19802 ( n24558 , n6073 , n11344 );
    not g19803 ( n18355 , n25617 );
    or g19804 ( n9939 , n20290 , n21577 );
    or g19805 ( n26610 , n22460 , n15788 );
    not g19806 ( n23983 , n11351 );
    xnor g19807 ( n21521 , n26235 , n8146 );
    or g19808 ( n19612 , n3440 , n6028 );
    xnor g19809 ( n1448 , n16482 , n5400 );
    xnor g19810 ( n18427 , n4858 , n23586 );
    not g19811 ( n12481 , n9494 );
    xnor g19812 ( n5603 , n26558 , n23551 );
    xnor g19813 ( n15094 , n2075 , n11713 );
    and g19814 ( n6361 , n16632 , n8460 );
    not g19815 ( n2906 , n7162 );
    xnor g19816 ( n25778 , n16200 , n2743 );
    nor g19817 ( n15981 , n12472 , n10397 );
    xnor g19818 ( n16299 , n4288 , n14902 );
    buf g19819 ( n6202 , n20014 );
    nor g19820 ( n20400 , n8101 , n15109 );
    nor g19821 ( n12764 , n6209 , n9507 );
    xnor g19822 ( n3891 , n10171 , n14499 );
    or g19823 ( n6821 , n9988 , n21667 );
    and g19824 ( n19811 , n23089 , n9830 );
    and g19825 ( n24729 , n25316 , n8068 );
    nor g19826 ( n25920 , n20957 , n25939 );
    not g19827 ( n1896 , n18295 );
    or g19828 ( n22189 , n8796 , n13833 );
    xnor g19829 ( n21626 , n16357 , n27187 );
    or g19830 ( n15702 , n2985 , n13578 );
    and g19831 ( n11260 , n7127 , n22013 );
    xnor g19832 ( n5169 , n2406 , n23251 );
    xnor g19833 ( n4661 , n21698 , n4514 );
    xnor g19834 ( n13383 , n8285 , n9323 );
    not g19835 ( n6805 , n20384 );
    and g19836 ( n21407 , n8575 , n5653 );
    xnor g19837 ( n21240 , n21028 , n4037 );
    or g19838 ( n3815 , n6321 , n9802 );
    and g19839 ( n12834 , n6227 , n14938 );
    or g19840 ( n12745 , n15198 , n10848 );
    or g19841 ( n4314 , n14858 , n12127 );
    nor g19842 ( n25390 , n8589 , n3619 );
    or g19843 ( n8115 , n323 , n5416 );
    and g19844 ( n12391 , n9031 , n26430 );
    and g19845 ( n25224 , n20085 , n13132 );
    or g19846 ( n24361 , n25514 , n6254 );
    xnor g19847 ( n7746 , n13783 , n25119 );
    not g19848 ( n2300 , n21529 );
    and g19849 ( n3175 , n16790 , n26 );
    or g19850 ( n7969 , n9425 , n22886 );
    or g19851 ( n17657 , n25132 , n11546 );
    and g19852 ( n9666 , n22982 , n1213 );
    and g19853 ( n10145 , n20393 , n26832 );
    xnor g19854 ( n7230 , n6758 , n19585 );
    xnor g19855 ( n6481 , n3053 , n5436 );
    or g19856 ( n23041 , n236 , n6540 );
    xnor g19857 ( n13004 , n23053 , n8612 );
    and g19858 ( n12115 , n10514 , n24806 );
    xnor g19859 ( n17815 , n5052 , n21670 );
    and g19860 ( n3684 , n15222 , n26579 );
    not g19861 ( n13292 , n21733 );
    not g19862 ( n13282 , n25442 );
    and g19863 ( n2983 , n17895 , n4197 );
    xnor g19864 ( n5275 , n6789 , n26417 );
    or g19865 ( n10796 , n21749 , n11676 );
    nor g19866 ( n20747 , n24375 , n14625 );
    xnor g19867 ( n19919 , n24266 , n10493 );
    and g19868 ( n24360 , n7909 , n16864 );
    xnor g19869 ( n5764 , n22895 , n17203 );
    xnor g19870 ( n3843 , n26051 , n18967 );
    xnor g19871 ( n26972 , n14166 , n25045 );
    nor g19872 ( n23768 , n13237 , n12921 );
    xnor g19873 ( n11640 , n17174 , n26144 );
    or g19874 ( n20601 , n20666 , n24251 );
    and g19875 ( n21747 , n9211 , n24394 );
    xnor g19876 ( n13617 , n13899 , n21037 );
    xnor g19877 ( n3072 , n5175 , n15322 );
    nor g19878 ( n14961 , n12960 , n6131 );
    xnor g19879 ( n15917 , n4222 , n25446 );
    and g19880 ( n5135 , n18779 , n17905 );
    not g19881 ( n14991 , n442 );
    xnor g19882 ( n20328 , n22660 , n26823 );
    xnor g19883 ( n11472 , n15177 , n13478 );
    not g19884 ( n7094 , n18345 );
    and g19885 ( n27184 , n26673 , n6820 );
    or g19886 ( n17844 , n2141 , n5790 );
    or g19887 ( n21625 , n25075 , n15564 );
    nor g19888 ( n24127 , n19277 , n5213 );
    and g19889 ( n17742 , n7736 , n18739 );
    xnor g19890 ( n25232 , n647 , n19941 );
    xnor g19891 ( n12771 , n11627 , n7593 );
    or g19892 ( n16578 , n15832 , n19889 );
    not g19893 ( n17641 , n2985 );
    buf g19894 ( n15901 , n5956 );
    not g19895 ( n10722 , n1889 );
    and g19896 ( n2969 , n9930 , n1062 );
    and g19897 ( n20663 , n26537 , n25162 );
    or g19898 ( n2844 , n10334 , n7557 );
    or g19899 ( n13971 , n1461 , n5996 );
    xnor g19900 ( n12987 , n1983 , n622 );
    nor g19901 ( n11115 , n4872 , n24009 );
    or g19902 ( n6739 , n13039 , n6043 );
    and g19903 ( n13304 , n4031 , n11697 );
    or g19904 ( n6153 , n14492 , n1125 );
    and g19905 ( n11571 , n21799 , n7620 );
    xnor g19906 ( n21349 , n23571 , n25104 );
    not g19907 ( n5449 , n13069 );
    xnor g19908 ( n12541 , n14641 , n13499 );
    xnor g19909 ( n7940 , n23600 , n25887 );
    not g19910 ( n8819 , n2698 );
    or g19911 ( n23934 , n21663 , n11323 );
    or g19912 ( n25833 , n12282 , n11003 );
    and g19913 ( n16122 , n21814 , n19073 );
    not g19914 ( n7056 , n14720 );
    or g19915 ( n19833 , n16744 , n24383 );
    and g19916 ( n24543 , n6712 , n15028 );
    and g19917 ( n15898 , n26041 , n19135 );
    or g19918 ( n15290 , n25663 , n9586 );
    or g19919 ( n11421 , n5106 , n9666 );
    or g19920 ( n18449 , n10947 , n23354 );
    xnor g19921 ( n19394 , n3044 , n23453 );
    or g19922 ( n13253 , n14620 , n26914 );
    xnor g19923 ( n19912 , n15930 , n23207 );
    or g19924 ( n11549 , n25466 , n16876 );
    not g19925 ( n15294 , n24072 );
    or g19926 ( n8493 , n18883 , n25146 );
    xnor g19927 ( n7937 , n2969 , n24742 );
    or g19928 ( n7446 , n24521 , n35 );
    and g19929 ( n2205 , n230 , n27109 );
    and g19930 ( n22932 , n12909 , n12173 );
    or g19931 ( n9338 , n13983 , n59 );
    not g19932 ( n3790 , n11377 );
    xnor g19933 ( n6893 , n9507 , n10158 );
    xnor g19934 ( n4429 , n4825 , n22383 );
    or g19935 ( n20625 , n17077 , n14620 );
    xnor g19936 ( n3235 , n22896 , n8848 );
    xnor g19937 ( n18592 , n1483 , n19539 );
    or g19938 ( n4406 , n20654 , n5362 );
    and g19939 ( n13323 , n7656 , n10104 );
    nor g19940 ( n14559 , n19236 , n21930 );
    and g19941 ( n7171 , n15638 , n11636 );
    not g19942 ( n21543 , n9247 );
    or g19943 ( n16212 , n11064 , n23524 );
    not g19944 ( n977 , n17455 );
    xnor g19945 ( n25470 , n19009 , n4927 );
    and g19946 ( n16471 , n16599 , n21202 );
    xnor g19947 ( n10915 , n15612 , n25884 );
    nor g19948 ( n18750 , n23200 , n8391 );
    xnor g19949 ( n14716 , n6501 , n623 );
    and g19950 ( n25616 , n12351 , n6503 );
    and g19951 ( n8318 , n1502 , n22128 );
    not g19952 ( n8344 , n2387 );
    not g19953 ( n17381 , n5842 );
    nor g19954 ( n21034 , n4951 , n26653 );
    and g19955 ( n22485 , n18341 , n18262 );
    not g19956 ( n16559 , n18826 );
    or g19957 ( n7837 , n6907 , n23280 );
    or g19958 ( n15016 , n8439 , n11106 );
    and g19959 ( n1542 , n4011 , n26002 );
    or g19960 ( n10031 , n16190 , n23696 );
    xnor g19961 ( n21809 , n2371 , n19255 );
    not g19962 ( n9586 , n10577 );
    xnor g19963 ( n12827 , n2377 , n19633 );
    or g19964 ( n19463 , n5986 , n23907 );
    nor g19965 ( n12117 , n25877 , n5026 );
    or g19966 ( n14682 , n5146 , n8957 );
    or g19967 ( n7493 , n979 , n6968 );
    not g19968 ( n8853 , n21858 );
    and g19969 ( n11019 , n1284 , n8876 );
    and g19970 ( n25070 , n21918 , n18974 );
    or g19971 ( n14863 , n5826 , n23597 );
    or g19972 ( n1569 , n16537 , n11783 );
    xnor g19973 ( n26522 , n24984 , n7275 );
    xnor g19974 ( n4168 , n2729 , n22298 );
    xnor g19975 ( n12385 , n22330 , n17913 );
    or g19976 ( n7550 , n14790 , n5105 );
    or g19977 ( n19388 , n22793 , n15016 );
    and g19978 ( n19341 , n4841 , n2714 );
    and g19979 ( n11081 , n14728 , n8570 );
    xnor g19980 ( n7792 , n7407 , n3030 );
    or g19981 ( n26476 , n24963 , n10412 );
    xnor g19982 ( n21316 , n18409 , n5704 );
    nor g19983 ( n1781 , n25049 , n23451 );
    nor g19984 ( n1095 , n22892 , n5165 );
    nor g19985 ( n8370 , n19762 , n9789 );
    or g19986 ( n13777 , n18649 , n13968 );
    xnor g19987 ( n14620 , n4036 , n7330 );
    and g19988 ( n15995 , n1558 , n17305 );
    xnor g19989 ( n17997 , n15236 , n23692 );
    nor g19990 ( n20612 , n17047 , n851 );
    and g19991 ( n23416 , n6924 , n18283 );
    or g19992 ( n26308 , n23711 , n16785 );
    or g19993 ( n20765 , n24457 , n19181 );
    xnor g19994 ( n15206 , n23061 , n21276 );
    nor g19995 ( n11417 , n16712 , n10053 );
    or g19996 ( n20949 , n1051 , n18365 );
    xnor g19997 ( n27051 , n18917 , n16368 );
    and g19998 ( n18435 , n14338 , n18422 );
    or g19999 ( n19512 , n10490 , n13324 );
    xnor g20000 ( n10263 , n10763 , n22379 );
    nor g20001 ( n3904 , n6218 , n19652 );
    or g20002 ( n23679 , n22879 , n12616 );
    xnor g20003 ( n25979 , n26264 , n21905 );
    nor g20004 ( n16380 , n10501 , n5914 );
    xnor g20005 ( n26058 , n22935 , n4407 );
    not g20006 ( n25827 , n10709 );
    or g20007 ( n15510 , n16670 , n17247 );
    not g20008 ( n21982 , n15652 );
    nor g20009 ( n24162 , n20959 , n26947 );
    not g20010 ( n13269 , n12385 );
    xnor g20011 ( n19923 , n9123 , n1632 );
    or g20012 ( n19140 , n9490 , n4955 );
    or g20013 ( n12925 , n18639 , n22399 );
    not g20014 ( n13907 , n8319 );
    xnor g20015 ( n20915 , n18389 , n11401 );
    xnor g20016 ( n15362 , n3324 , n2272 );
    not g20017 ( n2165 , n18638 );
    or g20018 ( n11778 , n17061 , n25419 );
    xnor g20019 ( n27006 , n11486 , n13781 );
    nor g20020 ( n5079 , n18934 , n11086 );
    nor g20021 ( n25529 , n23677 , n19717 );
    xnor g20022 ( n15588 , n5773 , n20012 );
    or g20023 ( n17884 , n17173 , n12236 );
    or g20024 ( n22560 , n22313 , n761 );
    not g20025 ( n18846 , n10785 );
    xnor g20026 ( n4770 , n24287 , n1225 );
    xnor g20027 ( n195 , n23878 , n1163 );
    or g20028 ( n11332 , n24662 , n23046 );
    xnor g20029 ( n15139 , n5892 , n1231 );
    or g20030 ( n10016 , n22971 , n20827 );
    xnor g20031 ( n2291 , n8602 , n3387 );
    and g20032 ( n16956 , n8121 , n7723 );
    nor g20033 ( n1264 , n1406 , n10372 );
    xnor g20034 ( n19459 , n23932 , n4939 );
    xnor g20035 ( n4523 , n25700 , n16803 );
    xnor g20036 ( n24826 , n13836 , n25652 );
    xnor g20037 ( n22406 , n15167 , n20036 );
    and g20038 ( n21447 , n19026 , n20473 );
    and g20039 ( n8471 , n2119 , n12982 );
    xnor g20040 ( n11600 , n10384 , n19575 );
    xnor g20041 ( n8251 , n25889 , n7885 );
    xnor g20042 ( n22395 , n21769 , n14779 );
    xnor g20043 ( n2728 , n26979 , n1152 );
    xnor g20044 ( n1092 , n21810 , n10235 );
    and g20045 ( n18638 , n22720 , n1158 );
    or g20046 ( n15720 , n13165 , n12689 );
    xnor g20047 ( n16765 , n12994 , n15594 );
    or g20048 ( n13763 , n2045 , n9992 );
    or g20049 ( n372 , n7204 , n19426 );
    xnor g20050 ( n22822 , n6309 , n15661 );
    xnor g20051 ( n15873 , n12956 , n1118 );
    and g20052 ( n22085 , n3744 , n12248 );
    and g20053 ( n6934 , n6228 , n16248 );
    nor g20054 ( n10687 , n12070 , n3496 );
    or g20055 ( n7074 , n5816 , n1329 );
    not g20056 ( n21743 , n2813 );
    not g20057 ( n13873 , n12702 );
    not g20058 ( n20006 , n26463 );
    xnor g20059 ( n22945 , n13317 , n27104 );
    or g20060 ( n17694 , n4028 , n21187 );
    not g20061 ( n24933 , n19317 );
    and g20062 ( n8209 , n12272 , n16709 );
    or g20063 ( n6806 , n17710 , n3531 );
    or g20064 ( n20490 , n2927 , n26677 );
    xnor g20065 ( n26055 , n20338 , n2756 );
    xnor g20066 ( n6248 , n9016 , n9120 );
    or g20067 ( n12792 , n10037 , n678 );
    xnor g20068 ( n3565 , n17626 , n25241 );
    xnor g20069 ( n4166 , n11840 , n23059 );
    or g20070 ( n15195 , n18773 , n1645 );
    and g20071 ( n16540 , n771 , n23383 );
    xnor g20072 ( n6711 , n14997 , n8461 );
    nor g20073 ( n9857 , n26882 , n19618 );
    not g20074 ( n15125 , n26744 );
    not g20075 ( n21162 , n513 );
    and g20076 ( n5815 , n5127 , n21110 );
    or g20077 ( n16042 , n2302 , n14535 );
    nor g20078 ( n11055 , n5617 , n22414 );
    nor g20079 ( n13243 , n20570 , n23962 );
    not g20080 ( n9736 , n24684 );
    xnor g20081 ( n10626 , n17762 , n16247 );
    or g20082 ( n17048 , n16658 , n20740 );
    not g20083 ( n17536 , n14366 );
    or g20084 ( n1710 , n19996 , n10421 );
    or g20085 ( n2465 , n9068 , n24319 );
    and g20086 ( n10755 , n25969 , n2447 );
    xnor g20087 ( n15428 , n17211 , n25509 );
    xnor g20088 ( n12621 , n10616 , n13060 );
    or g20089 ( n25736 , n4878 , n2477 );
    or g20090 ( n5148 , n22169 , n23783 );
    nor g20091 ( n7261 , n1662 , n20946 );
    or g20092 ( n11545 , n3455 , n14549 );
    or g20093 ( n20387 , n17802 , n16487 );
    not g20094 ( n21701 , n16249 );
    and g20095 ( n17763 , n26633 , n2900 );
    or g20096 ( n2888 , n2875 , n601 );
    and g20097 ( n11383 , n4362 , n8514 );
    and g20098 ( n8445 , n16048 , n7843 );
    nor g20099 ( n16133 , n7071 , n14848 );
    xnor g20100 ( n5984 , n4484 , n2175 );
    or g20101 ( n10981 , n13679 , n11811 );
    or g20102 ( n25741 , n15138 , n26318 );
    not g20103 ( n12837 , n3697 );
    nor g20104 ( n22733 , n15905 , n23160 );
    not g20105 ( n21937 , n27037 );
    xnor g20106 ( n24213 , n12233 , n2552 );
    not g20107 ( n15715 , n11749 );
    or g20108 ( n12428 , n8015 , n20255 );
    and g20109 ( n26700 , n19382 , n26362 );
    nor g20110 ( n1275 , n9076 , n704 );
    and g20111 ( n26238 , n17396 , n19185 );
    or g20112 ( n6978 , n25271 , n7566 );
    and g20113 ( n27047 , n8764 , n5755 );
    and g20114 ( n11585 , n631 , n12734 );
    and g20115 ( n9658 , n21971 , n3640 );
    xnor g20116 ( n26705 , n9276 , n23199 );
    or g20117 ( n21589 , n19488 , n2462 );
    or g20118 ( n9735 , n18345 , n6179 );
    xnor g20119 ( n19158 , n16648 , n9602 );
    and g20120 ( n14565 , n5611 , n20600 );
    and g20121 ( n3936 , n18444 , n17028 );
    nor g20122 ( n5986 , n17351 , n16468 );
    or g20123 ( n14019 , n21543 , n3663 );
    and g20124 ( n11923 , n20256 , n15567 );
    or g20125 ( n5476 , n4020 , n4789 );
    and g20126 ( n13566 , n5971 , n4742 );
    not g20127 ( n1571 , n25736 );
    nor g20128 ( n4807 , n15967 , n2783 );
    or g20129 ( n4912 , n23225 , n3500 );
    xnor g20130 ( n20756 , n22442 , n3324 );
    xnor g20131 ( n21854 , n23974 , n24879 );
    or g20132 ( n1226 , n13088 , n7674 );
    xnor g20133 ( n24873 , n5448 , n4026 );
    xnor g20134 ( n3186 , n10087 , n23534 );
    xnor g20135 ( n13923 , n11204 , n3806 );
    or g20136 ( n22931 , n19616 , n8309 );
    or g20137 ( n11925 , n9904 , n22921 );
    and g20138 ( n11164 , n11369 , n17113 );
    and g20139 ( n24550 , n17452 , n5683 );
    and g20140 ( n14290 , n8216 , n10703 );
    or g20141 ( n5307 , n21289 , n13418 );
    not g20142 ( n21951 , n15023 );
    not g20143 ( n16822 , n19184 );
    xnor g20144 ( n4334 , n1941 , n2659 );
    nor g20145 ( n16512 , n1896 , n16396 );
    xnor g20146 ( n26921 , n24064 , n7764 );
    xnor g20147 ( n15128 , n20203 , n10705 );
    and g20148 ( n17874 , n12321 , n21145 );
    xnor g20149 ( n11506 , n26987 , n23917 );
    xnor g20150 ( n16107 , n20423 , n13093 );
    and g20151 ( n12489 , n13100 , n412 );
    and g20152 ( n25239 , n13114 , n16641 );
    nor g20153 ( n2428 , n14981 , n2718 );
    or g20154 ( n9009 , n19298 , n22843 );
    and g20155 ( n6624 , n26424 , n841 );
    or g20156 ( n5864 , n21428 , n10550 );
    or g20157 ( n17262 , n6396 , n22402 );
    or g20158 ( n15669 , n371 , n25196 );
    or g20159 ( n5033 , n7902 , n13926 );
    and g20160 ( n19647 , n16762 , n1726 );
    xnor g20161 ( n15019 , n26485 , n14506 );
    and g20162 ( n19072 , n3966 , n23077 );
    xnor g20163 ( n5408 , n5176 , n21771 );
    or g20164 ( n378 , n16122 , n23050 );
    and g20165 ( n2107 , n8536 , n13236 );
    and g20166 ( n10498 , n26480 , n1546 );
    or g20167 ( n9688 , n2060 , n6371 );
    xnor g20168 ( n15516 , n14790 , n604 );
    xnor g20169 ( n13356 , n17233 , n686 );
    not g20170 ( n25898 , n5791 );
    xnor g20171 ( n2191 , n7409 , n21755 );
    or g20172 ( n7368 , n20297 , n13603 );
    or g20173 ( n7926 , n11144 , n23166 );
    or g20174 ( n3847 , n22208 , n10902 );
    not g20175 ( n3744 , n1696 );
    not g20176 ( n25914 , n25240 );
    or g20177 ( n8494 , n26582 , n7107 );
    xnor g20178 ( n10020 , n7785 , n1558 );
    or g20179 ( n2452 , n3759 , n22682 );
    and g20180 ( n5346 , n8611 , n10729 );
    and g20181 ( n9852 , n14965 , n10389 );
    or g20182 ( n20272 , n4033 , n8170 );
    xnor g20183 ( n18687 , n20585 , n21144 );
    and g20184 ( n6680 , n155 , n22140 );
    xnor g20185 ( n20703 , n7678 , n11579 );
    or g20186 ( n8486 , n26094 , n19735 );
    or g20187 ( n26345 , n15901 , n21751 );
    or g20188 ( n21597 , n6545 , n12271 );
    and g20189 ( n22221 , n26207 , n6757 );
    or g20190 ( n1131 , n8498 , n3656 );
    or g20191 ( n15020 , n15880 , n10434 );
    and g20192 ( n14014 , n6115 , n7385 );
    and g20193 ( n3171 , n17287 , n16852 );
    xnor g20194 ( n17038 , n23307 , n13495 );
    nor g20195 ( n25742 , n6356 , n1449 );
    xnor g20196 ( n15534 , n11940 , n9860 );
    or g20197 ( n2605 , n5498 , n16886 );
    or g20198 ( n22984 , n13513 , n5537 );
    xnor g20199 ( n22574 , n3468 , n15289 );
    and g20200 ( n14390 , n17993 , n23145 );
    or g20201 ( n25329 , n24245 , n3138 );
    or g20202 ( n24763 , n16509 , n14945 );
    not g20203 ( n22012 , n2489 );
    xnor g20204 ( n6606 , n6773 , n583 );
    or g20205 ( n3777 , n23283 , n529 );
    and g20206 ( n8830 , n12384 , n4667 );
    or g20207 ( n20086 , n11131 , n21022 );
    and g20208 ( n1995 , n21443 , n27014 );
    xnor g20209 ( n18454 , n8363 , n1222 );
    or g20210 ( n15396 , n9961 , n15010 );
    and g20211 ( n19796 , n2959 , n25493 );
    and g20212 ( n11253 , n9951 , n19093 );
    not g20213 ( n4570 , n8898 );
    or g20214 ( n9280 , n26194 , n12299 );
    or g20215 ( n3703 , n6304 , n14290 );
    or g20216 ( n8617 , n18849 , n11066 );
    and g20217 ( n4704 , n11993 , n8541 );
    not g20218 ( n24383 , n21537 );
    xnor g20219 ( n391 , n6104 , n3945 );
    xnor g20220 ( n3668 , n19580 , n26829 );
    nor g20221 ( n3589 , n189 , n5685 );
    xnor g20222 ( n11412 , n21232 , n2279 );
    not g20223 ( n18947 , n16221 );
    xnor g20224 ( n5343 , n9114 , n27104 );
    xnor g20225 ( n4112 , n5048 , n25843 );
    or g20226 ( n17188 , n4514 , n4122 );
    xnor g20227 ( n3390 , n22873 , n18760 );
    nor g20228 ( n25458 , n8910 , n25018 );
    not g20229 ( n9820 , n26573 );
    not g20230 ( n15730 , n4587 );
    not g20231 ( n19074 , n3618 );
    or g20232 ( n2543 , n19429 , n14610 );
    not g20233 ( n15191 , n5777 );
    or g20234 ( n12953 , n25515 , n6949 );
    and g20235 ( n9411 , n26255 , n14210 );
    and g20236 ( n1093 , n10197 , n8800 );
    nor g20237 ( n15373 , n3072 , n20145 );
    nor g20238 ( n842 , n4923 , n14042 );
    or g20239 ( n3466 , n20131 , n224 );
    not g20240 ( n1952 , n1915 );
    xnor g20241 ( n10080 , n9598 , n7759 );
    not g20242 ( n3284 , n8087 );
    or g20243 ( n7641 , n15707 , n12174 );
    and g20244 ( n5592 , n6616 , n17009 );
    or g20245 ( n12958 , n6138 , n16965 );
    or g20246 ( n23908 , n20768 , n25609 );
    nor g20247 ( n18073 , n63 , n22359 );
    not g20248 ( n8083 , n19210 );
    and g20249 ( n19320 , n25534 , n5100 );
    or g20250 ( n23402 , n19588 , n5211 );
    xnor g20251 ( n20728 , n10781 , n26512 );
    xnor g20252 ( n27153 , n8308 , n12522 );
    and g20253 ( n14756 , n24300 , n21408 );
    xnor g20254 ( n6517 , n17212 , n16627 );
    and g20255 ( n20649 , n20091 , n27050 );
    and g20256 ( n19889 , n9292 , n14039 );
    or g20257 ( n21073 , n6824 , n7624 );
    xnor g20258 ( n10241 , n25562 , n12216 );
    or g20259 ( n25056 , n26878 , n6213 );
    and g20260 ( n7244 , n3715 , n291 );
    xnor g20261 ( n4746 , n11382 , n20250 );
    not g20262 ( n15760 , n11578 );
    nor g20263 ( n21327 , n20826 , n18068 );
    and g20264 ( n918 , n3276 , n13177 );
    and g20265 ( n18336 , n20773 , n4750 );
    xnor g20266 ( n23215 , n4719 , n5822 );
    or g20267 ( n8107 , n15364 , n10054 );
    nor g20268 ( n17248 , n3306 , n21567 );
    not g20269 ( n7677 , n18187 );
    xnor g20270 ( n25617 , n10678 , n25166 );
    xnor g20271 ( n19863 , n4317 , n22332 );
    nor g20272 ( n5434 , n17902 , n20249 );
    and g20273 ( n4210 , n20904 , n11573 );
    nor g20274 ( n2131 , n1994 , n16559 );
    xnor g20275 ( n25607 , n4787 , n17405 );
    or g20276 ( n7732 , n24827 , n297 );
    or g20277 ( n23994 , n9948 , n308 );
    not g20278 ( n6779 , n3603 );
    not g20279 ( n6464 , n4410 );
    not g20280 ( n9570 , n2783 );
    not g20281 ( n10353 , n15305 );
    xnor g20282 ( n19974 , n20928 , n18315 );
    and g20283 ( n1312 , n9038 , n13232 );
    xnor g20284 ( n23649 , n17902 , n337 );
    and g20285 ( n17331 , n12341 , n13945 );
    xnor g20286 ( n819 , n14460 , n22026 );
    nor g20287 ( n14913 , n19604 , n7359 );
    or g20288 ( n412 , n11033 , n5699 );
    or g20289 ( n10473 , n23016 , n25515 );
    xnor g20290 ( n18343 , n15270 , n11488 );
    xnor g20291 ( n20402 , n21901 , n5660 );
    xnor g20292 ( n26137 , n15271 , n12161 );
    xnor g20293 ( n6679 , n7978 , n10202 );
    and g20294 ( n5052 , n20584 , n11795 );
    or g20295 ( n15467 , n11143 , n8646 );
    and g20296 ( n16648 , n1506 , n8039 );
    xnor g20297 ( n8276 , n8643 , n27168 );
    and g20298 ( n15390 , n16385 , n25484 );
    or g20299 ( n25325 , n22768 , n18915 );
    xnor g20300 ( n13832 , n13784 , n17302 );
    and g20301 ( n10674 , n6332 , n12374 );
    xnor g20302 ( n20690 , n8526 , n17458 );
    xnor g20303 ( n4506 , n8647 , n18973 );
    or g20304 ( n17424 , n22731 , n9087 );
    or g20305 ( n14755 , n22925 , n13854 );
    and g20306 ( n13046 , n8968 , n4126 );
    xnor g20307 ( n4275 , n3534 , n18756 );
    xnor g20308 ( n23203 , n19526 , n17863 );
    xnor g20309 ( n11054 , n788 , n16573 );
    and g20310 ( n23706 , n3481 , n14054 );
    xnor g20311 ( n12186 , n12366 , n11736 );
    nor g20312 ( n8840 , n25413 , n152 );
    not g20313 ( n13534 , n24600 );
    xnor g20314 ( n19736 , n24190 , n20804 );
    or g20315 ( n18757 , n25740 , n12045 );
    xnor g20316 ( n7497 , n10682 , n10234 );
    xnor g20317 ( n19377 , n5198 , n25501 );
    not g20318 ( n12576 , n25345 );
    xnor g20319 ( n23796 , n18113 , n1467 );
    or g20320 ( n22565 , n14685 , n13282 );
    or g20321 ( n22409 , n25020 , n24385 );
    or g20322 ( n12284 , n21462 , n19872 );
    xnor g20323 ( n11838 , n5405 , n23834 );
    xnor g20324 ( n20291 , n19665 , n10065 );
    or g20325 ( n20983 , n16324 , n23688 );
    and g20326 ( n17426 , n7068 , n2353 );
    xnor g20327 ( n1225 , n6471 , n10448 );
    xnor g20328 ( n7780 , n4968 , n500 );
    nor g20329 ( n1706 , n11615 , n23779 );
    xnor g20330 ( n21067 , n13708 , n23775 );
    not g20331 ( n17601 , n13367 );
    xnor g20332 ( n3543 , n7092 , n24486 );
    xnor g20333 ( n18003 , n20587 , n16457 );
    or g20334 ( n15819 , n21605 , n21898 );
    xnor g20335 ( n4646 , n11833 , n4019 );
    not g20336 ( n15445 , n4372 );
    and g20337 ( n14207 , n1736 , n12243 );
    and g20338 ( n21716 , n6204 , n23254 );
    or g20339 ( n16096 , n16084 , n9557 );
    and g20340 ( n2717 , n26382 , n1217 );
    xnor g20341 ( n14580 , n9892 , n23911 );
    not g20342 ( n2498 , n18003 );
    or g20343 ( n10808 , n23469 , n17666 );
    and g20344 ( n26181 , n19710 , n7965 );
    and g20345 ( n18289 , n22018 , n5979 );
    not g20346 ( n14519 , n2547 );
    not g20347 ( n16637 , n22537 );
    xnor g20348 ( n26222 , n15592 , n25009 );
    or g20349 ( n19052 , n25004 , n1630 );
    and g20350 ( n22747 , n25437 , n15098 );
    nor g20351 ( n22599 , n2659 , n11926 );
    and g20352 ( n17488 , n8851 , n4087 );
    or g20353 ( n24792 , n1956 , n3877 );
    xnor g20354 ( n17500 , n24413 , n11054 );
    xnor g20355 ( n23544 , n6541 , n329 );
    not g20356 ( n23030 , n8869 );
    or g20357 ( n22810 , n7194 , n12180 );
    xnor g20358 ( n14493 , n26222 , n6944 );
    xnor g20359 ( n20868 , n1465 , n23304 );
    xnor g20360 ( n17873 , n11266 , n9926 );
    not g20361 ( n26471 , n11910 );
    and g20362 ( n2158 , n9870 , n4171 );
    and g20363 ( n13221 , n14863 , n16578 );
    xnor g20364 ( n5739 , n11012 , n20118 );
    xnor g20365 ( n1055 , n15776 , n14009 );
    or g20366 ( n20313 , n5475 , n3834 );
    or g20367 ( n491 , n26116 , n1497 );
    or g20368 ( n7309 , n10601 , n5845 );
    or g20369 ( n12193 , n2257 , n21666 );
    not g20370 ( n15944 , n1667 );
    xnor g20371 ( n11933 , n20434 , n3692 );
    not g20372 ( n7365 , n1386 );
    xnor g20373 ( n1509 , n25565 , n21993 );
    xnor g20374 ( n16239 , n17048 , n22624 );
    xnor g20375 ( n11556 , n14397 , n16812 );
    not g20376 ( n18598 , n4256 );
    and g20377 ( n2773 , n4858 , n6895 );
    nor g20378 ( n17365 , n1881 , n26857 );
    and g20379 ( n4098 , n7991 , n4805 );
    xnor g20380 ( n25516 , n20548 , n4813 );
    xnor g20381 ( n19540 , n18076 , n19920 );
    and g20382 ( n22930 , n24650 , n23729 );
    xnor g20383 ( n26970 , n22678 , n783 );
    nor g20384 ( n4530 , n18295 , n23313 );
    or g20385 ( n1538 , n22978 , n15228 );
    or g20386 ( n14928 , n11477 , n22207 );
    and g20387 ( n1100 , n11598 , n10042 );
    or g20388 ( n23115 , n22105 , n5465 );
    not g20389 ( n11740 , n647 );
    and g20390 ( n11173 , n19883 , n21468 );
    not g20391 ( n12855 , n20663 );
    xnor g20392 ( n11127 , n18648 , n23782 );
    xnor g20393 ( n21291 , n26130 , n16909 );
    and g20394 ( n10403 , n18642 , n1899 );
    or g20395 ( n411 , n19393 , n16982 );
    not g20396 ( n15218 , n20950 );
    nor g20397 ( n13641 , n22511 , n10251 );
    or g20398 ( n20296 , n7343 , n11108 );
    nor g20399 ( n12825 , n23476 , n12410 );
    not g20400 ( n5498 , n12650 );
    nor g20401 ( n3402 , n10250 , n13976 );
    or g20402 ( n20038 , n16133 , n10675 );
    or g20403 ( n1699 , n24 , n2876 );
    and g20404 ( n12414 , n5942 , n7023 );
    xnor g20405 ( n20442 , n9462 , n17251 );
    or g20406 ( n13574 , n11417 , n19700 );
    or g20407 ( n26983 , n6186 , n2134 );
    or g20408 ( n17761 , n12784 , n12887 );
    xnor g20409 ( n10354 , n16822 , n14661 );
    not g20410 ( n9187 , n1350 );
    and g20411 ( n21656 , n17473 , n24463 );
    nor g20412 ( n3335 , n4859 , n2570 );
    and g20413 ( n26278 , n6720 , n5396 );
    xor g20414 ( n10392 , n4239 , n11034 );
    or g20415 ( n9281 , n4752 , n13114 );
    nor g20416 ( n14646 , n25900 , n12697 );
    not g20417 ( n6962 , n23253 );
    or g20418 ( n8995 , n16186 , n2643 );
    or g20419 ( n11773 , n24535 , n20052 );
    or g20420 ( n19998 , n12760 , n20295 );
    or g20421 ( n13229 , n10831 , n18500 );
    not g20422 ( n19633 , n19309 );
    or g20423 ( n13482 , n21057 , n13742 );
    xnor g20424 ( n1560 , n25637 , n19540 );
    not g20425 ( n13995 , n5517 );
    not g20426 ( n21575 , n13336 );
    and g20427 ( n3943 , n19952 , n10178 );
    not g20428 ( n10389 , n2599 );
    or g20429 ( n14239 , n9494 , n21723 );
    nor g20430 ( n20993 , n17549 , n20506 );
    not g20431 ( n15144 , n23692 );
    not g20432 ( n26252 , n11650 );
    xnor g20433 ( n26386 , n8391 , n23200 );
    or g20434 ( n469 , n11303 , n10037 );
    xnor g20435 ( n20148 , n7769 , n26625 );
    not g20436 ( n7713 , n25670 );
    or g20437 ( n11015 , n19705 , n16021 );
    not g20438 ( n12788 , n4160 );
    nor g20439 ( n5898 , n14254 , n11502 );
    xnor g20440 ( n14468 , n17938 , n20966 );
    and g20441 ( n18769 , n19165 , n41 );
    or g20442 ( n21220 , n20643 , n12082 );
    or g20443 ( n15971 , n5494 , n1487 );
    and g20444 ( n15169 , n7007 , n8699 );
    or g20445 ( n16986 , n24608 , n26016 );
    or g20446 ( n9353 , n10597 , n10126 );
    not g20447 ( n24940 , n5305 );
    nor g20448 ( n10495 , n16349 , n604 );
    xnor g20449 ( n7587 , n22274 , n24129 );
    xnor g20450 ( n15590 , n25154 , n12323 );
    xnor g20451 ( n15160 , n12650 , n11220 );
    and g20452 ( n204 , n6251 , n5092 );
    or g20453 ( n6350 , n5205 , n6065 );
    or g20454 ( n20555 , n7612 , n20883 );
    xnor g20455 ( n18347 , n20929 , n23068 );
    not g20456 ( n350 , n22154 );
    xnor g20457 ( n11080 , n19823 , n2611 );
    or g20458 ( n1021 , n26747 , n7923 );
    and g20459 ( n5267 , n14826 , n20342 );
    or g20460 ( n1442 , n26513 , n20902 );
    or g20461 ( n15028 , n12125 , n7828 );
    xnor g20462 ( n3692 , n7809 , n25100 );
    or g20463 ( n18080 , n23775 , n4601 );
    or g20464 ( n10058 , n26140 , n843 );
    xnor g20465 ( n25667 , n8541 , n12826 );
    not g20466 ( n19949 , n2659 );
    not g20467 ( n6731 , n23602 );
    xnor g20468 ( n23900 , n4439 , n15281 );
    xnor g20469 ( n22480 , n15388 , n8046 );
    xnor g20470 ( n1887 , n27104 , n18295 );
    not g20471 ( n6698 , n3937 );
    or g20472 ( n8096 , n9514 , n17204 );
    xnor g20473 ( n8403 , n27107 , n7518 );
    xnor g20474 ( n1516 , n9017 , n25647 );
    or g20475 ( n24770 , n6024 , n24334 );
    nor g20476 ( n5531 , n4938 , n14130 );
    and g20477 ( n14893 , n10805 , n247 );
    and g20478 ( n16718 , n8101 , n3019 );
    and g20479 ( n1402 , n15918 , n21021 );
    xnor g20480 ( n20201 , n16721 , n19941 );
    or g20481 ( n9568 , n443 , n4797 );
    xnor g20482 ( n18906 , n2952 , n1639 );
    nor g20483 ( n24322 , n15856 , n14357 );
    xnor g20484 ( n14305 , n182 , n15190 );
    xnor g20485 ( n1044 , n7965 , n6290 );
    and g20486 ( n16730 , n1406 , n19473 );
    xnor g20487 ( n9448 , n16357 , n16880 );
    and g20488 ( n9998 , n15365 , n1973 );
    or g20489 ( n4107 , n4600 , n2264 );
    xnor g20490 ( n800 , n2995 , n18281 );
    and g20491 ( n4840 , n12513 , n14106 );
    or g20492 ( n9132 , n13985 , n12155 );
    and g20493 ( n4308 , n18051 , n8124 );
    or g20494 ( n2737 , n2895 , n16972 );
    xnor g20495 ( n807 , n11650 , n7750 );
    nor g20496 ( n21845 , n2559 , n2117 );
    not g20497 ( n12477 , n8649 );
    nor g20498 ( n23225 , n2659 , n23704 );
    or g20499 ( n20451 , n23413 , n14491 );
    or g20500 ( n15197 , n16192 , n19795 );
    and g20501 ( n17669 , n13876 , n9582 );
    xnor g20502 ( n26229 , n13585 , n9051 );
    or g20503 ( n13686 , n22585 , n22527 );
    xnor g20504 ( n8871 , n17388 , n4242 );
    or g20505 ( n3788 , n8571 , n11285 );
    or g20506 ( n1268 , n26986 , n16832 );
    not g20507 ( n26326 , n23851 );
    or g20508 ( n21314 , n21380 , n16210 );
    nor g20509 ( n22594 , n22895 , n17845 );
    xnor g20510 ( n1970 , n10057 , n8920 );
    xnor g20511 ( n17898 , n16267 , n9240 );
    xnor g20512 ( n3038 , n7082 , n21782 );
    nor g20513 ( n17588 , n3734 , n14257 );
    or g20514 ( n2262 , n17166 , n25989 );
    and g20515 ( n22532 , n25135 , n20136 );
    and g20516 ( n13741 , n24683 , n25801 );
    and g20517 ( n2075 , n26772 , n15718 );
    or g20518 ( n21356 , n25320 , n18836 );
    and g20519 ( n2529 , n22041 , n5099 );
    xnor g20520 ( n21850 , n25117 , n25629 );
    nor g20521 ( n9612 , n20132 , n2810 );
    and g20522 ( n20457 , n748 , n7070 );
    xnor g20523 ( n17583 , n17324 , n23875 );
    xnor g20524 ( n7515 , n10275 , n25240 );
    not g20525 ( n10993 , n13463 );
    nor g20526 ( n6212 , n22607 , n15512 );
    or g20527 ( n3997 , n13099 , n17545 );
    nor g20528 ( n12933 , n15109 , n5532 );
    xnor g20529 ( n24714 , n16432 , n1667 );
    xnor g20530 ( n16305 , n15007 , n12281 );
    xnor g20531 ( n4180 , n1449 , n6356 );
    xnor g20532 ( n13082 , n10940 , n2240 );
    not g20533 ( n9826 , n17970 );
    xnor g20534 ( n12566 , n11872 , n2532 );
    xnor g20535 ( n20494 , n5077 , n13914 );
    xnor g20536 ( n27181 , n11982 , n7931 );
    xnor g20537 ( n9213 , n19393 , n16982 );
    nor g20538 ( n16781 , n16722 , n21101 );
    xnor g20539 ( n11274 , n12398 , n25694 );
    and g20540 ( n12456 , n311 , n12721 );
    xnor g20541 ( n9345 , n14276 , n18035 );
    or g20542 ( n26837 , n22176 , n10666 );
    or g20543 ( n24570 , n16879 , n24235 );
    or g20544 ( n7675 , n24325 , n23913 );
    or g20545 ( n5457 , n7261 , n26601 );
    xnor g20546 ( n12999 , n11908 , n24538 );
    nor g20547 ( n12287 , n8687 , n966 );
    nor g20548 ( n8056 , n22436 , n11146 );
    and g20549 ( n5901 , n21152 , n25496 );
    and g20550 ( n23193 , n7279 , n23378 );
    or g20551 ( n19251 , n3536 , n3109 );
    or g20552 ( n14483 , n3116 , n16696 );
    or g20553 ( n8870 , n15134 , n5179 );
    nor g20554 ( n9540 , n23528 , n9099 );
    or g20555 ( n25401 , n6581 , n17781 );
    or g20556 ( n7442 , n7311 , n19944 );
    not g20557 ( n6300 , n19524 );
    xnor g20558 ( n26454 , n2057 , n19603 );
    xnor g20559 ( n18288 , n25662 , n1482 );
    and g20560 ( n20885 , n21741 , n6926 );
    not g20561 ( n17685 , n11892 );
    or g20562 ( n24489 , n23030 , n6385 );
    xnor g20563 ( n16398 , n22726 , n16451 );
    nor g20564 ( n6689 , n26178 , n21290 );
    and g20565 ( n20217 , n9518 , n14509 );
    not g20566 ( n6466 , n3038 );
    xnor g20567 ( n16426 , n24630 , n6775 );
    nor g20568 ( n5501 , n20796 , n21460 );
    and g20569 ( n13454 , n15875 , n13352 );
    and g20570 ( n18468 , n23195 , n8666 );
    xnor g20571 ( n21404 , n22437 , n5788 );
    and g20572 ( n22437 , n5323 , n22258 );
    or g20573 ( n24653 , n20260 , n18205 );
    xnor g20574 ( n14999 , n18607 , n22159 );
    xnor g20575 ( n19617 , n1068 , n7608 );
    not g20576 ( n20716 , n18398 );
    or g20577 ( n7877 , n4801 , n11970 );
    not g20578 ( n12530 , n23035 );
    nor g20579 ( n17449 , n16319 , n6293 );
    xnor g20580 ( n22503 , n12889 , n24298 );
    nor g20581 ( n10456 , n3750 , n24397 );
    or g20582 ( n17574 , n883 , n5452 );
    nor g20583 ( n6421 , n3069 , n15289 );
    xnor g20584 ( n10437 , n21515 , n25000 );
    nor g20585 ( n25733 , n9969 , n14705 );
    or g20586 ( n8377 , n2192 , n12897 );
    and g20587 ( n15471 , n486 , n18042 );
    not g20588 ( n10369 , n17256 );
    not g20589 ( n2960 , n14981 );
    not g20590 ( n4531 , n24578 );
    and g20591 ( n3887 , n26908 , n21552 );
    xnor g20592 ( n15165 , n12260 , n20997 );
    or g20593 ( n14495 , n20841 , n13528 );
    nor g20594 ( n2766 , n24608 , n428 );
    nor g20595 ( n21686 , n21004 , n18265 );
    or g20596 ( n10476 , n17596 , n22469 );
    xnor g20597 ( n9228 , n11749 , n14954 );
    or g20598 ( n7739 , n22091 , n18861 );
    xnor g20599 ( n8166 , n10727 , n20932 );
    or g20600 ( n13636 , n11521 , n22735 );
    or g20601 ( n24082 , n13605 , n16365 );
    xnor g20602 ( n8234 , n12430 , n17780 );
    xnor g20603 ( n12300 , n20384 , n6659 );
    xnor g20604 ( n7285 , n24930 , n15515 );
    or g20605 ( n16646 , n20572 , n21877 );
    xnor g20606 ( n24139 , n21222 , n26752 );
    xnor g20607 ( n16724 , n20816 , n6772 );
    not g20608 ( n22636 , n15600 );
    xnor g20609 ( n2747 , n7164 , n17193 );
    and g20610 ( n8009 , n18261 , n6413 );
    nor g20611 ( n3745 , n26553 , n15041 );
    xnor g20612 ( n2065 , n1433 , n26344 );
    or g20613 ( n6754 , n3130 , n5983 );
    not g20614 ( n21406 , n13297 );
    or g20615 ( n19481 , n16477 , n11697 );
    xnor g20616 ( n22079 , n25865 , n4403 );
    or g20617 ( n19799 , n26162 , n6814 );
    xnor g20618 ( n11822 , n16702 , n7793 );
    and g20619 ( n6360 , n7180 , n3333 );
    xnor g20620 ( n12426 , n7200 , n19307 );
    and g20621 ( n26577 , n8493 , n865 );
    nor g20622 ( n6451 , n25629 , n3795 );
    xnor g20623 ( n14457 , n940 , n17694 );
    nor g20624 ( n14129 , n25376 , n18617 );
    xnor g20625 ( n21705 , n23068 , n18907 );
    xnor g20626 ( n3316 , n5083 , n4640 );
    and g20627 ( n7173 , n23850 , n9101 );
    and g20628 ( n6940 , n1406 , n1978 );
    xnor g20629 ( n6500 , n8773 , n18599 );
    nor g20630 ( n6617 , n7260 , n13368 );
    and g20631 ( n16095 , n4216 , n24069 );
    xnor g20632 ( n12295 , n23967 , n17251 );
    or g20633 ( n13355 , n9284 , n25683 );
    xnor g20634 ( n14668 , n350 , n18004 );
    or g20635 ( n8145 , n7772 , n10671 );
    nor g20636 ( n22346 , n7963 , n6590 );
    xnor g20637 ( n11469 , n8224 , n20151 );
    and g20638 ( n24389 , n5427 , n19633 );
    xnor g20639 ( n24452 , n10666 , n8656 );
    or g20640 ( n21382 , n15530 , n2739 );
    not g20641 ( n23094 , n13240 );
    or g20642 ( n24046 , n14861 , n24697 );
    or g20643 ( n11441 , n19962 , n22426 );
    or g20644 ( n9417 , n9944 , n23842 );
    and g20645 ( n4894 , n15442 , n18450 );
    nor g20646 ( n23617 , n10593 , n4792 );
    or g20647 ( n10604 , n2628 , n14345 );
    and g20648 ( n9923 , n6841 , n4036 );
    or g20649 ( n13964 , n23923 , n16608 );
    not g20650 ( n25701 , n1869 );
    or g20651 ( n24232 , n6574 , n14351 );
    and g20652 ( n18209 , n21140 , n10241 );
    or g20653 ( n25626 , n1089 , n5094 );
    xnor g20654 ( n16428 , n3034 , n16207 );
    xnor g20655 ( n16753 , n20326 , n5916 );
    or g20656 ( n26071 , n20829 , n18171 );
    nor g20657 ( n10436 , n24305 , n5012 );
    not g20658 ( n23686 , n1047 );
    nor g20659 ( n16389 , n6692 , n21249 );
    or g20660 ( n11369 , n3078 , n15698 );
    or g20661 ( n25772 , n11957 , n3873 );
    xnor g20662 ( n11447 , n7330 , n8439 );
    not g20663 ( n10075 , n23310 );
    or g20664 ( n18309 , n2230 , n16722 );
    xnor g20665 ( n5956 , n19893 , n15171 );
    nor g20666 ( n7632 , n18398 , n25807 );
    not g20667 ( n24959 , n1550 );
    not g20668 ( n22382 , n18726 );
    and g20669 ( n9115 , n3111 , n19671 );
    xnor g20670 ( n16174 , n11089 , n972 );
    and g20671 ( n19101 , n13966 , n17441 );
    xnor g20672 ( n10774 , n15389 , n24468 );
    xnor g20673 ( n21488 , n3136 , n26913 );
    buf g20674 ( n26876 , n7634 );
    nor g20675 ( n11145 , n1612 , n728 );
    not g20676 ( n8779 , n26888 );
    nor g20677 ( n22802 , n18880 , n2978 );
    xnor g20678 ( n2177 , n20192 , n21649 );
    xnor g20679 ( n22050 , n21821 , n10257 );
    or g20680 ( n6478 , n3817 , n8761 );
    xnor g20681 ( n26816 , n14880 , n8210 );
    xnor g20682 ( n5584 , n16439 , n10275 );
    xnor g20683 ( n19783 , n8721 , n1040 );
    or g20684 ( n4419 , n14514 , n26187 );
    xnor g20685 ( n13486 , n8726 , n24911 );
    and g20686 ( n5292 , n2597 , n10682 );
    and g20687 ( n23106 , n13675 , n12010 );
    and g20688 ( n1247 , n3404 , n11943 );
    xnor g20689 ( n16009 , n14313 , n25180 );
    and g20690 ( n26613 , n19429 , n23519 );
    or g20691 ( n9604 , n5154 , n4138 );
    and g20692 ( n4082 , n17878 , n7920 );
    xnor g20693 ( n8139 , n18250 , n7235 );
    not g20694 ( n20536 , n25464 );
    xnor g20695 ( n9124 , n14558 , n12479 );
    xnor g20696 ( n5247 , n20948 , n1658 );
    and g20697 ( n18356 , n7715 , n19528 );
    xnor g20698 ( n3789 , n1831 , n3320 );
    xnor g20699 ( n2528 , n6082 , n3228 );
    not g20700 ( n4050 , n763 );
    xnor g20701 ( n7253 , n16750 , n20819 );
    nor g20702 ( n5651 , n2858 , n26486 );
    xnor g20703 ( n15179 , n67 , n11494 );
    or g20704 ( n4169 , n14628 , n16846 );
    and g20705 ( n15518 , n23356 , n17801 );
    and g20706 ( n199 , n3035 , n24997 );
    nor g20707 ( n2930 , n8220 , n7361 );
    xnor g20708 ( n15671 , n19614 , n21222 );
    and g20709 ( n17468 , n11666 , n17750 );
    and g20710 ( n6654 , n8565 , n16363 );
    xnor g20711 ( n6223 , n22065 , n17865 );
    not g20712 ( n14848 , n26016 );
    xnor g20713 ( n17508 , n3719 , n25119 );
    or g20714 ( n25945 , n18560 , n2958 );
    nor g20715 ( n7245 , n19849 , n18421 );
    and g20716 ( n13288 , n2632 , n7368 );
    xnor g20717 ( n6593 , n27037 , n23913 );
    not g20718 ( n15385 , n11769 );
    and g20719 ( n7226 , n1577 , n22885 );
    not g20720 ( n2607 , n11333 );
    nor g20721 ( n740 , n11220 , n3425 );
    xnor g20722 ( n16925 , n22964 , n21060 );
    or g20723 ( n18186 , n3591 , n3963 );
    xnor g20724 ( n20722 , n24054 , n10723 );
    and g20725 ( n17199 , n25329 , n12676 );
    xnor g20726 ( n17186 , n8857 , n19578 );
    xnor g20727 ( n11169 , n26912 , n12895 );
    and g20728 ( n21748 , n6318 , n96 );
    and g20729 ( n11675 , n23910 , n21339 );
    or g20730 ( n8369 , n2318 , n19038 );
    nor g20731 ( n4951 , n26000 , n14725 );
    and g20732 ( n14296 , n7206 , n6530 );
    or g20733 ( n1393 , n18829 , n27090 );
    xnor g20734 ( n23918 , n15113 , n21957 );
    or g20735 ( n6687 , n13577 , n26691 );
    xnor g20736 ( n4794 , n6104 , n24048 );
    xnor g20737 ( n23823 , n1451 , n16217 );
    xnor g20738 ( n18887 , n5646 , n2367 );
    xnor g20739 ( n18958 , n8244 , n6513 );
    or g20740 ( n7009 , n1365 , n12315 );
    and g20741 ( n23129 , n2331 , n13748 );
    or g20742 ( n490 , n24653 , n10746 );
    xnor g20743 ( n9602 , n16707 , n13037 );
    and g20744 ( n23167 , n6614 , n21305 );
    nor g20745 ( n15375 , n3919 , n26105 );
    and g20746 ( n7972 , n10657 , n1440 );
    not g20747 ( n11975 , n26069 );
    not g20748 ( n16028 , n24070 );
    or g20749 ( n20833 , n8348 , n12625 );
    and g20750 ( n5792 , n22401 , n17594 );
    or g20751 ( n24498 , n24729 , n1846 );
    not g20752 ( n25276 , n5727 );
    xnor g20753 ( n645 , n15930 , n14089 );
    xnor g20754 ( n20515 , n24312 , n5032 );
    or g20755 ( n9582 , n2617 , n13911 );
    xnor g20756 ( n23677 , n25007 , n14083 );
    nor g20757 ( n1912 , n22562 , n17412 );
    or g20758 ( n13118 , n7292 , n14510 );
    not g20759 ( n12138 , n24112 );
    or g20760 ( n18180 , n18431 , n11295 );
    and g20761 ( n6815 , n7692 , n16793 );
    or g20762 ( n15741 , n25744 , n15218 );
    and g20763 ( n15143 , n16827 , n7262 );
    or g20764 ( n18110 , n1192 , n5569 );
    not g20765 ( n24766 , n15440 );
    not g20766 ( n5816 , n6611 );
    nor g20767 ( n25283 , n20384 , n8008 );
    and g20768 ( n12865 , n3820 , n3684 );
    xnor g20769 ( n19104 , n6990 , n26449 );
    or g20770 ( n19810 , n7424 , n4052 );
    nor g20771 ( n22682 , n14302 , n12837 );
    or g20772 ( n21217 , n21846 , n24161 );
    nor g20773 ( n16904 , n3472 , n25085 );
    or g20774 ( n26182 , n11691 , n11073 );
    not g20775 ( n10128 , n8387 );
    not g20776 ( n16147 , n12241 );
    not g20777 ( n15474 , n22270 );
    xnor g20778 ( n13409 , n10106 , n26072 );
    nor g20779 ( n24276 , n4490 , n5261 );
    xnor g20780 ( n11739 , n11011 , n20179 );
    nor g20781 ( n11315 , n5060 , n2808 );
    xnor g20782 ( n2765 , n22318 , n21626 );
    or g20783 ( n9798 , n9003 , n1735 );
    nor g20784 ( n12918 , n8008 , n14516 );
    xnor g20785 ( n20726 , n2160 , n11220 );
    xnor g20786 ( n6602 , n9666 , n6747 );
    not g20787 ( n12402 , n12648 );
    or g20788 ( n15533 , n21517 , n8582 );
    and g20789 ( n630 , n22174 , n22277 );
    not g20790 ( n13451 , n11792 );
    or g20791 ( n24678 , n21016 , n21668 );
    xnor g20792 ( n21960 , n855 , n12234 );
    and g20793 ( n21995 , n15850 , n22206 );
    and g20794 ( n1847 , n7242 , n16123 );
    xnor g20795 ( n1066 , n14678 , n10938 );
    xnor g20796 ( n18143 , n18222 , n26518 );
    not g20797 ( n23877 , n7134 );
    nor g20798 ( n5298 , n5226 , n26724 );
    or g20799 ( n13701 , n20169 , n8718 );
    and g20800 ( n17550 , n13036 , n23307 );
    not g20801 ( n22558 , n10201 );
    nor g20802 ( n24193 , n17542 , n15146 );
    or g20803 ( n9158 , n1715 , n15490 );
    nor g20804 ( n9073 , n20032 , n4844 );
    or g20805 ( n1407 , n11559 , n22861 );
    xnor g20806 ( n13168 , n22555 , n16287 );
    and g20807 ( n6305 , n10519 , n11310 );
    or g20808 ( n4386 , n11745 , n18249 );
    xnor g20809 ( n19308 , n9701 , n6076 );
    xnor g20810 ( n11407 , n20986 , n25471 );
    not g20811 ( n5796 , n1204 );
    and g20812 ( n21214 , n10264 , n21039 );
    xnor g20813 ( n11314 , n14689 , n20179 );
    xnor g20814 ( n18714 , n1337 , n26073 );
    or g20815 ( n9722 , n8447 , n26254 );
    or g20816 ( n3534 , n4493 , n768 );
    not g20817 ( n23798 , n8769 );
    or g20818 ( n18441 , n19827 , n17297 );
    xnor g20819 ( n24266 , n20041 , n7257 );
    xnor g20820 ( n20839 , n11649 , n9872 );
    not g20821 ( n22613 , n2698 );
    or g20822 ( n19278 , n5511 , n12270 );
    not g20823 ( n12543 , n20658 );
    nor g20824 ( n5838 , n9180 , n1262 );
    or g20825 ( n20309 , n12841 , n16361 );
    nor g20826 ( n23554 , n12561 , n11305 );
    or g20827 ( n21837 , n3346 , n19311 );
    xnor g20828 ( n10917 , n2088 , n26979 );
    not g20829 ( n15309 , n15127 );
    and g20830 ( n26663 , n11292 , n3146 );
    not g20831 ( n5039 , n11408 );
    xnor g20832 ( n14694 , n26452 , n5098 );
    and g20833 ( n24999 , n10536 , n17650 );
    or g20834 ( n21815 , n9770 , n26100 );
    or g20835 ( n21669 , n11043 , n1252 );
    and g20836 ( n16463 , n4910 , n1638 );
    or g20837 ( n9861 , n7967 , n19154 );
    and g20838 ( n23447 , n25822 , n13047 );
    xnor g20839 ( n6774 , n16726 , n20068 );
    or g20840 ( n4302 , n25651 , n5921 );
    xnor g20841 ( n2771 , n22207 , n26851 );
    xnor g20842 ( n1034 , n21249 , n6692 );
    and g20843 ( n955 , n1426 , n10105 );
    and g20844 ( n25913 , n24565 , n3729 );
    or g20845 ( n8882 , n7617 , n23706 );
    not g20846 ( n6599 , n2730 );
    xnor g20847 ( n11929 , n13250 , n10685 );
    nor g20848 ( n1037 , n22370 , n6034 );
    or g20849 ( n21043 , n1643 , n20460 );
    or g20850 ( n12037 , n22532 , n2260 );
    not g20851 ( n8295 , n9313 );
    and g20852 ( n26328 , n10558 , n18832 );
    xnor g20853 ( n11832 , n20099 , n3541 );
    and g20854 ( n14602 , n1146 , n8469 );
    xnor g20855 ( n13421 , n17660 , n19758 );
    not g20856 ( n15582 , n11448 );
    nor g20857 ( n3419 , n15572 , n2989 );
    xnor g20858 ( n10262 , n47 , n12230 );
    and g20859 ( n8777 , n18345 , n6179 );
    or g20860 ( n6614 , n6321 , n5026 );
    or g20861 ( n1713 , n13863 , n20134 );
    nor g20862 ( n5919 , n22422 , n18648 );
    not g20863 ( n23608 , n14984 );
    and g20864 ( n11319 , n19380 , n13134 );
    or g20865 ( n11049 , n25004 , n10158 );
    not g20866 ( n25268 , n26000 );
    nor g20867 ( n5316 , n1765 , n21309 );
    xnor g20868 ( n2599 , n11636 , n23673 );
    not g20869 ( n23415 , n2778 );
    not g20870 ( n25582 , n1872 );
    or g20871 ( n26682 , n26914 , n26962 );
    xnor g20872 ( n22711 , n2729 , n9210 );
    and g20873 ( n8247 , n26567 , n9385 );
    xnor g20874 ( n1413 , n9745 , n14900 );
    nor g20875 ( n3085 , n7088 , n3132 );
    xnor g20876 ( n18333 , n2310 , n16769 );
    nor g20877 ( n20782 , n19313 , n5974 );
    xnor g20878 ( n25100 , n16505 , n10080 );
    or g20879 ( n7264 , n13419 , n14937 );
    and g20880 ( n6933 , n15201 , n22705 );
    or g20881 ( n5312 , n6790 , n10000 );
    xnor g20882 ( n25076 , n10083 , n13654 );
    xnor g20883 ( n13158 , n19295 , n22631 );
    xnor g20884 ( n2043 , n10109 , n26742 );
    and g20885 ( n1150 , n533 , n24858 );
    or g20886 ( n18017 , n18548 , n12239 );
    xnor g20887 ( n26001 , n25674 , n5585 );
    xnor g20888 ( n10793 , n18806 , n14518 );
    xnor g20889 ( n5833 , n16121 , n7366 );
    nor g20890 ( n3409 , n21871 , n1314 );
    xnor g20891 ( n10516 , n23200 , n19116 );
    or g20892 ( n22248 , n8910 , n22392 );
    or g20893 ( n21147 , n22329 , n26369 );
    xnor g20894 ( n20713 , n15774 , n13947 );
    or g20895 ( n13011 , n10514 , n24806 );
    buf g20896 ( n5924 , n9054 );
    or g20897 ( n7007 , n13621 , n10114 );
    not g20898 ( n15204 , n11824 );
    xnor g20899 ( n11053 , n17430 , n24311 );
    not g20900 ( n18004 , n21636 );
    xor g20901 ( n5454 , n1398 , n9507 );
    and g20902 ( n25875 , n19514 , n2415 );
    not g20903 ( n1759 , n2189 );
    and g20904 ( n10238 , n14285 , n2934 );
    xnor g20905 ( n12050 , n4742 , n870 );
    and g20906 ( n24941 , n26643 , n383 );
    and g20907 ( n19002 , n7126 , n24120 );
    xnor g20908 ( n18034 , n21222 , n26565 );
    or g20909 ( n3487 , n17198 , n23882 );
    or g20910 ( n18948 , n21437 , n3242 );
    or g20911 ( n8699 , n21790 , n18815 );
    not g20912 ( n21436 , n5462 );
    or g20913 ( n14822 , n25237 , n21710 );
    or g20914 ( n10588 , n11638 , n18382 );
    xnor g20915 ( n16786 , n25749 , n2113 );
    xnor g20916 ( n4999 , n21394 , n894 );
    or g20917 ( n18845 , n25752 , n8173 );
    not g20918 ( n15266 , n10658 );
    or g20919 ( n26279 , n15229 , n20029 );
    or g20920 ( n11553 , n17757 , n1150 );
    and g20921 ( n25806 , n17368 , n2539 );
    not g20922 ( n8650 , n17326 );
    nor g20923 ( n15311 , n11559 , n2328 );
    xnor g20924 ( n15407 , n23928 , n8692 );
    nor g20925 ( n21435 , n144 , n10710 );
    or g20926 ( n10932 , n23736 , n8702 );
    nor g20927 ( n15887 , n11898 , n23166 );
    nor g20928 ( n25424 , n15766 , n6105 );
    nor g20929 ( n8082 , n26961 , n864 );
    nor g20930 ( n11232 , n6387 , n455 );
    or g20931 ( n16302 , n17211 , n4345 );
    and g20932 ( n16552 , n26279 , n23902 );
    or g20933 ( n10221 , n9802 , n10017 );
    xnor g20934 ( n9350 , n8319 , n12493 );
    xnor g20935 ( n3002 , n2622 , n19500 );
    xnor g20936 ( n3049 , n8128 , n23766 );
    nor g20937 ( n11665 , n8513 , n10709 );
    or g20938 ( n23382 , n16698 , n26881 );
    or g20939 ( n6781 , n2517 , n9194 );
    and g20940 ( n1029 , n13293 , n17388 );
    or g20941 ( n23794 , n10193 , n4755 );
    nor g20942 ( n1250 , n13989 , n20138 );
    not g20943 ( n18798 , n618 );
    not g20944 ( n18931 , n25538 );
    and g20945 ( n13274 , n17784 , n725 );
    xnor g20946 ( n4865 , n25115 , n22491 );
    and g20947 ( n13615 , n14886 , n17639 );
    and g20948 ( n11850 , n21855 , n13395 );
    xnor g20949 ( n21665 , n17242 , n24926 );
    or g20950 ( n15212 , n1365 , n4087 );
    or g20951 ( n1977 , n14431 , n8906 );
    nor g20952 ( n9712 , n5719 , n7195 );
    not g20953 ( n417 , n25289 );
    and g20954 ( n24735 , n26380 , n18974 );
    xnor g20955 ( n20941 , n2462 , n19488 );
    xnor g20956 ( n12851 , n24069 , n13684 );
    or g20957 ( n8393 , n24524 , n4069 );
    or g20958 ( n11821 , n15682 , n4080 );
    not g20959 ( n22125 , n26399 );
    and g20960 ( n3321 , n26563 , n10809 );
    xnor g20961 ( n16522 , n26211 , n21219 );
    or g20962 ( n21558 , n602 , n16963 );
    xnor g20963 ( n19015 , n16547 , n4085 );
    or g20964 ( n8710 , n4285 , n16119 );
    and g20965 ( n12274 , n21370 , n16083 );
    and g20966 ( n8990 , n11745 , n6825 );
    xnor g20967 ( n5156 , n25377 , n16482 );
    xnor g20968 ( n97 , n11802 , n11502 );
    and g20969 ( n19161 , n21541 , n16177 );
    or g20970 ( n10062 , n22286 , n199 );
    not g20971 ( n8612 , n23745 );
    and g20972 ( n9890 , n13918 , n21595 );
    nor g20973 ( n25082 , n14588 , n942 );
    xnor g20974 ( n657 , n10758 , n13562 );
    or g20975 ( n18422 , n17550 , n14022 );
    xnor g20976 ( n19301 , n24898 , n22861 );
    xnor g20977 ( n14354 , n23616 , n18444 );
    xnor g20978 ( n23060 , n15135 , n18204 );
    not g20979 ( n11608 , n14756 );
    or g20980 ( n3763 , n3796 , n4416 );
    xnor g20981 ( n150 , n18066 , n20111 );
    nor g20982 ( n10740 , n12366 , n23071 );
    not g20983 ( n14410 , n3132 );
    or g20984 ( n9174 , n378 , n5779 );
    xnor g20985 ( n5564 , n22011 , n17042 );
    and g20986 ( n22330 , n11761 , n23496 );
    not g20987 ( n20550 , n9625 );
    or g20988 ( n19300 , n8504 , n24400 );
    or g20989 ( n4427 , n11583 , n3190 );
    or g20990 ( n1417 , n16748 , n14959 );
    xnor g20991 ( n24049 , n12543 , n15508 );
    nor g20992 ( n26188 , n9240 , n16267 );
    nor g20993 ( n22313 , n8367 , n2113 );
    xnor g20994 ( n15801 , n21478 , n833 );
    xnor g20995 ( n7754 , n23486 , n11734 );
    not g20996 ( n656 , n9906 );
    xnor g20997 ( n10340 , n21690 , n9409 );
    and g20998 ( n8658 , n3945 , n21998 );
    or g20999 ( n15778 , n11322 , n26098 );
    or g21000 ( n26200 , n10117 , n19825 );
    or g21001 ( n11966 , n2926 , n25520 );
    and g21002 ( n18516 , n4957 , n14979 );
    and g21003 ( n13867 , n10877 , n8560 );
    xnor g21004 ( n14669 , n6262 , n11258 );
    xnor g21005 ( n17530 , n8816 , n21679 );
    and g21006 ( n6264 , n19393 , n16982 );
    xnor g21007 ( n16734 , n20043 , n11071 );
    or g21008 ( n10525 , n5631 , n13381 );
    xor g21009 ( n12629 , n6743 , n7713 );
    or g21010 ( n5034 , n7524 , n8799 );
    not g21011 ( n1458 , n20077 );
    xnor g21012 ( n21768 , n11716 , n12775 );
    xnor g21013 ( n3075 , n19656 , n16456 );
    or g21014 ( n21204 , n9921 , n2736 );
    nor g21015 ( n18419 , n3744 , n12248 );
    xnor g21016 ( n6848 , n18052 , n16073 );
    nor g21017 ( n17887 , n1340 , n1099 );
    and g21018 ( n19606 , n9127 , n8390 );
    or g21019 ( n26632 , n10274 , n14168 );
    and g21020 ( n13728 , n9701 , n6076 );
    xnor g21021 ( n18626 , n18171 , n1738 );
    or g21022 ( n9515 , n21406 , n10034 );
    and g21023 ( n16191 , n22369 , n11358 );
    or g21024 ( n1146 , n13775 , n8389 );
    or g21025 ( n11796 , n9942 , n2210 );
    or g21026 ( n17482 , n17543 , n10445 );
    or g21027 ( n26190 , n635 , n22415 );
    not g21028 ( n17423 , n23895 );
    and g21029 ( n9439 , n22585 , n26837 );
    xnor g21030 ( n3835 , n2859 , n608 );
    nor g21031 ( n27131 , n19196 , n6122 );
    or g21032 ( n3350 , n7778 , n4083 );
    xnor g21033 ( n22910 , n14105 , n1001 );
    not g21034 ( n12454 , n8363 );
    or g21035 ( n7274 , n22554 , n21890 );
    xnor g21036 ( n11185 , n1998 , n13230 );
    or g21037 ( n18989 , n12715 , n10303 );
    or g21038 ( n845 , n10990 , n2834 );
    and g21039 ( n6531 , n795 , n10857 );
    or g21040 ( n2589 , n246 , n8763 );
    nor g21041 ( n12844 , n21380 , n24170 );
    nor g21042 ( n4720 , n8236 , n728 );
    or g21043 ( n17136 , n8244 , n8431 );
    xnor g21044 ( n3141 , n11697 , n19711 );
    xnor g21045 ( n22753 , n16401 , n9259 );
    or g21046 ( n16621 , n7949 , n15562 );
    or g21047 ( n4355 , n25432 , n21447 );
    nor g21048 ( n10598 , n15268 , n333 );
    not g21049 ( n21928 , n7710 );
    not g21050 ( n2231 , n20631 );
    or g21051 ( n12909 , n4342 , n9401 );
    xnor g21052 ( n17481 , n15693 , n24701 );
    and g21053 ( n15312 , n16164 , n14221 );
    or g21054 ( n7723 , n12965 , n17571 );
    or g21055 ( n24753 , n20486 , n22556 );
    or g21056 ( n18620 , n11087 , n16437 );
    xnor g21057 ( n15322 , n5822 , n7963 );
    xnor g21058 ( n17201 , n5055 , n3827 );
    not g21059 ( n10152 , n16576 );
    nor g21060 ( n3046 , n167 , n1339 );
    or g21061 ( n22419 , n21125 , n926 );
    xnor g21062 ( n21685 , n14893 , n15919 );
    and g21063 ( n3529 , n21644 , n18555 );
    xnor g21064 ( n19725 , n2109 , n963 );
    not g21065 ( n17995 , n13189 );
    or g21066 ( n22051 , n14963 , n10620 );
    or g21067 ( n13059 , n16762 , n22662 );
    not g21068 ( n950 , n1608 );
    and g21069 ( n9221 , n4983 , n24045 );
    not g21070 ( n25071 , n7212 );
    not g21071 ( n20921 , n3839 );
    xnor g21072 ( n19497 , n16364 , n18891 );
    or g21073 ( n26559 , n1558 , n17305 );
    nor g21074 ( n902 , n14465 , n25074 );
    xnor g21075 ( n10672 , n23277 , n11975 );
    nor g21076 ( n22360 , n12554 , n22871 );
    not g21077 ( n22849 , n10096 );
    or g21078 ( n499 , n19760 , n19994 );
    and g21079 ( n17949 , n24705 , n26444 );
    or g21080 ( n19183 , n21052 , n21576 );
    not g21081 ( n19186 , n11945 );
    or g21082 ( n20093 , n8202 , n14209 );
    and g21083 ( n4728 , n7238 , n14923 );
    xnor g21084 ( n24648 , n17556 , n6896 );
    and g21085 ( n1815 , n13951 , n24355 );
    xnor g21086 ( n1693 , n18649 , n3984 );
    xnor g21087 ( n7820 , n25289 , n4195 );
    nor g21088 ( n14904 , n16722 , n13708 );
    nor g21089 ( n26322 , n13333 , n15681 );
    and g21090 ( n1209 , n16166 , n10407 );
    xnor g21091 ( n11221 , n17433 , n15574 );
    and g21092 ( n13248 , n21462 , n19872 );
    or g21093 ( n22343 , n5867 , n11930 );
    xnor g21094 ( n9245 , n14581 , n19187 );
    and g21095 ( n22045 , n6992 , n2824 );
    or g21096 ( n9548 , n11294 , n20608 );
    xnor g21097 ( n2574 , n8452 , n3141 );
    not g21098 ( n18279 , n14061 );
    or g21099 ( n13242 , n23886 , n13245 );
    xnor g21100 ( n23959 , n23589 , n12891 );
    and g21101 ( n22008 , n17144 , n15641 );
    not g21102 ( n11013 , n11651 );
    not g21103 ( n16762 , n5048 );
    xnor g21104 ( n18689 , n22110 , n11378 );
    and g21105 ( n20741 , n19878 , n20888 );
    nor g21106 ( n10863 , n11381 , n4294 );
    xnor g21107 ( n15753 , n1118 , n4665 );
    xnor g21108 ( n12744 , n5425 , n1081 );
    xnor g21109 ( n8352 , n7482 , n16382 );
    xnor g21110 ( n26323 , n26580 , n13485 );
    or g21111 ( n18856 , n9901 , n13447 );
    nor g21112 ( n10707 , n20826 , n626 );
    and g21113 ( n26294 , n20023 , n12734 );
    and g21114 ( n19086 , n18811 , n21330 );
    not g21115 ( n8176 , n23892 );
    not g21116 ( n12418 , n24863 );
    not g21117 ( n7059 , n20029 );
    and g21118 ( n13399 , n338 , n10806 );
    or g21119 ( n13871 , n6819 , n11671 );
    not g21120 ( n16679 , n13425 );
    or g21121 ( n8121 , n10527 , n5387 );
    and g21122 ( n11543 , n19256 , n16941 );
    or g21123 ( n21706 , n22042 , n6808 );
    nor g21124 ( n5908 , n4149 , n22454 );
    nor g21125 ( n15121 , n1222 , n8292 );
    not g21126 ( n7088 , n21957 );
    xnor g21127 ( n1020 , n23633 , n24284 );
    and g21128 ( n13723 , n2069 , n25315 );
    and g21129 ( n15692 , n20614 , n8141 );
    or g21130 ( n12979 , n20064 , n14345 );
    buf g21131 ( n9291 , n22002 );
    xnor g21132 ( n12998 , n12198 , n10405 );
    or g21133 ( n9977 , n13844 , n19394 );
    and g21134 ( n17531 , n24004 , n21081 );
    and g21135 ( n13381 , n18191 , n18188 );
    xnor g21136 ( n5081 , n25738 , n6861 );
    or g21137 ( n9772 , n12455 , n974 );
    xnor g21138 ( n17852 , n23568 , n27120 );
    and g21139 ( n6208 , n10786 , n22922 );
    or g21140 ( n14013 , n8244 , n22820 );
    or g21141 ( n23077 , n191 , n18072 );
    nor g21142 ( n2811 , n25872 , n2994 );
    not g21143 ( n15581 , n15918 );
    xnor g21144 ( n252 , n26728 , n25655 );
    xnor g21145 ( n19121 , n17911 , n6814 );
    or g21146 ( n16916 , n4999 , n27017 );
    nor g21147 ( n12952 , n9249 , n14732 );
    nor g21148 ( n17445 , n21843 , n20659 );
    and g21149 ( n792 , n5710 , n4439 );
    not g21150 ( n21370 , n22516 );
    not g21151 ( n22836 , n9656 );
    or g21152 ( n9995 , n11045 , n11220 );
    nor g21153 ( n11731 , n9392 , n12049 );
    not g21154 ( n24717 , n24764 );
    not g21155 ( n13308 , n2964 );
    not g21156 ( n19895 , n6254 );
    xnor g21157 ( n6523 , n1670 , n25087 );
    xnor g21158 ( n16394 , n3359 , n14570 );
    xnor g21159 ( n7506 , n3460 , n19477 );
    or g21160 ( n20712 , n17975 , n4202 );
    xnor g21161 ( n4067 , n19 , n13803 );
    xnor g21162 ( n6603 , n11124 , n11469 );
    xnor g21163 ( n10647 , n18388 , n19851 );
    nor g21164 ( n17817 , n17909 , n24650 );
    xnor g21165 ( n4432 , n7559 , n12484 );
    xnor g21166 ( n20704 , n8684 , n6783 );
    nor g21167 ( n292 , n26443 , n23807 );
    xnor g21168 ( n16989 , n12016 , n14921 );
    nor g21169 ( n836 , n5611 , n24420 );
    xnor g21170 ( n23014 , n3145 , n6745 );
    and g21171 ( n24707 , n23360 , n12785 );
    xnor g21172 ( n19044 , n14980 , n9822 );
    not g21173 ( n2248 , n15681 );
    xnor g21174 ( n7734 , n19441 , n26796 );
    or g21175 ( n10382 , n17826 , n24620 );
    not g21176 ( n4687 , n18909 );
    xnor g21177 ( n17070 , n16572 , n22385 );
    not g21178 ( n13443 , n9942 );
    xnor g21179 ( n13277 , n15978 , n11949 );
    xnor g21180 ( n10064 , n15616 , n20104 );
    or g21181 ( n15052 , n20228 , n13856 );
    xnor g21182 ( n6751 , n21997 , n18483 );
    or g21183 ( n17582 , n23540 , n11923 );
    or g21184 ( n13531 , n1792 , n19521 );
    xnor g21185 ( n2732 , n2851 , n4835 );
    xnor g21186 ( n22484 , n12629 , n10232 );
    or g21187 ( n10579 , n323 , n8403 );
    not g21188 ( n1205 , n15743 );
    xnor g21189 ( n6276 , n6343 , n9842 );
    or g21190 ( n0 , n8660 , n8328 );
    xnor g21191 ( n11155 , n1974 , n17576 );
    and g21192 ( n3488 , n19963 , n3432 );
    and g21193 ( n19750 , n6836 , n23517 );
    xnor g21194 ( n23825 , n23166 , n4306 );
    not g21195 ( n18426 , n17094 );
    not g21196 ( n12962 , n13912 );
    or g21197 ( n18141 , n18882 , n8856 );
    xnor g21198 ( n6587 , n4733 , n2699 );
    xnor g21199 ( n7349 , n14681 , n188 );
    nor g21200 ( n19695 , n1531 , n7302 );
    not g21201 ( n20205 , n18483 );
    not g21202 ( n11457 , n16223 );
    and g21203 ( n215 , n16848 , n19628 );
    xnor g21204 ( n10024 , n6074 , n15556 );
    not g21205 ( n23417 , n24801 );
    xnor g21206 ( n16896 , n4831 , n21266 );
    xnor g21207 ( n8019 , n101 , n8416 );
    and g21208 ( n23736 , n22808 , n7824 );
    or g21209 ( n23531 , n4445 , n12574 );
    xnor g21210 ( n25254 , n16318 , n26118 );
    and g21211 ( n13067 , n6695 , n499 );
    xnor g21212 ( n14055 , n15271 , n26748 );
    or g21213 ( n14067 , n9363 , n11088 );
    xnor g21214 ( n12790 , n729 , n25692 );
    xnor g21215 ( n55 , n22776 , n2499 );
    not g21216 ( n5220 , n6307 );
    not g21217 ( n16663 , n6774 );
    xnor g21218 ( n18534 , n26211 , n15583 );
    or g21219 ( n12221 , n21634 , n2035 );
    or g21220 ( n10461 , n8948 , n9242 );
    xnor g21221 ( n6414 , n1152 , n25023 );
    not g21222 ( n26488 , n18951 );
    and g21223 ( n967 , n19911 , n26658 );
    or g21224 ( n4079 , n16593 , n25191 );
    or g21225 ( n4690 , n23455 , n25285 );
    or g21226 ( n13153 , n15560 , n7006 );
    or g21227 ( n10860 , n16695 , n6365 );
    xnor g21228 ( n8778 , n8241 , n2985 );
    and g21229 ( n27020 , n4469 , n7212 );
    or g21230 ( n23348 , n5144 , n5862 );
    xnor g21231 ( n22172 , n26216 , n8331 );
    and g21232 ( n23179 , n15829 , n7690 );
    or g21233 ( n26151 , n11921 , n1324 );
    and g21234 ( n13681 , n22918 , n20719 );
    not g21235 ( n10923 , n16948 );
    nor g21236 ( n1086 , n21715 , n25615 );
    or g21237 ( n7279 , n26695 , n23890 );
    not g21238 ( n16628 , n5558 );
    and g21239 ( n1434 , n3414 , n21465 );
    not g21240 ( n20015 , n20003 );
    not g21241 ( n26013 , n947 );
    xnor g21242 ( n4953 , n22206 , n5030 );
    or g21243 ( n2639 , n9431 , n7592 );
    xnor g21244 ( n24749 , n22985 , n20182 );
    not g21245 ( n24243 , n23344 );
    xnor g21246 ( n9142 , n22022 , n13832 );
    xnor g21247 ( n9743 , n13286 , n7096 );
    or g21248 ( n24149 , n14751 , n7927 );
    xnor g21249 ( n10534 , n9041 , n7117 );
    nor g21250 ( n4586 , n26318 , n18895 );
    or g21251 ( n25567 , n14099 , n13526 );
    nor g21252 ( n2196 , n6169 , n26302 );
    xnor g21253 ( n2301 , n6351 , n7731 );
    xnor g21254 ( n20623 , n22759 , n5435 );
    xnor g21255 ( n26156 , n1475 , n18694 );
    and g21256 ( n3044 , n17942 , n17059 );
    and g21257 ( n21376 , n26715 , n12690 );
    not g21258 ( n22197 , n17900 );
    or g21259 ( n23591 , n17933 , n25003 );
    and g21260 ( n12025 , n27174 , n9866 );
    xnor g21261 ( n17638 , n7874 , n15399 );
    xnor g21262 ( n7725 , n26811 , n3895 );
    nor g21263 ( n16405 , n2252 , n16672 );
    not g21264 ( n11374 , n19876 );
    or g21265 ( n14509 , n20541 , n21754 );
    xnor g21266 ( n22806 , n12513 , n8395 );
    or g21267 ( n12434 , n26170 , n8635 );
    xnor g21268 ( n15252 , n7689 , n3827 );
    or g21269 ( n10853 , n20427 , n13281 );
    xnor g21270 ( n27165 , n8176 , n9554 );
    and g21271 ( n6639 , n9798 , n17672 );
    and g21272 ( n21255 , n19684 , n14877 );
    not g21273 ( n7750 , n20901 );
    not g21274 ( n3411 , n19393 );
    xnor g21275 ( n909 , n17250 , n4409 );
    and g21276 ( n21221 , n21982 , n2606 );
    and g21277 ( n14473 , n11400 , n20130 );
    nor g21278 ( n10799 , n7640 , n3509 );
    xnor g21279 ( n3019 , n22280 , n18522 );
    xnor g21280 ( n6736 , n6297 , n7272 );
    not g21281 ( n8420 , n6456 );
    or g21282 ( n16402 , n14336 , n18149 );
    nor g21283 ( n11026 , n17579 , n6632 );
    or g21284 ( n10558 , n24417 , n4719 );
    or g21285 ( n9664 , n24417 , n24907 );
    and g21286 ( n26254 , n5967 , n21835 );
    and g21287 ( n15837 , n8732 , n4651 );
    and g21288 ( n20230 , n3362 , n21695 );
    xnor g21289 ( n16898 , n18974 , n21918 );
    or g21290 ( n8141 , n16668 , n5982 );
    or g21291 ( n26561 , n522 , n20432 );
    nor g21292 ( n16003 , n1205 , n7494 );
    and g21293 ( n10061 , n26634 , n7314 );
    xnor g21294 ( n5946 , n26549 , n4482 );
    and g21295 ( n7352 , n20395 , n11604 );
    or g21296 ( n25769 , n26658 , n15539 );
    or g21297 ( n10615 , n24231 , n9305 );
    or g21298 ( n24010 , n10555 , n23291 );
    not g21299 ( n21380 , n18537 );
    and g21300 ( n4743 , n23615 , n4521 );
    xnor g21301 ( n19707 , n6566 , n10875 );
    xnor g21302 ( n6127 , n12824 , n7545 );
    not g21303 ( n7621 , n8324 );
    nor g21304 ( n22602 , n26963 , n22828 );
    or g21305 ( n19346 , n11901 , n24044 );
    xnor g21306 ( n12895 , n10649 , n6289 );
    and g21307 ( n8954 , n10726 , n124 );
    and g21308 ( n13524 , n2411 , n9062 );
    and g21309 ( n24803 , n3494 , n6211 );
    or g21310 ( n5219 , n14723 , n12086 );
    or g21311 ( n9059 , n27160 , n13948 );
    xnor g21312 ( n18323 , n64 , n5851 );
    or g21313 ( n9795 , n10744 , n23243 );
    xnor g21314 ( n23984 , n24494 , n24359 );
    and g21315 ( n14776 , n10883 , n19778 );
    and g21316 ( n17386 , n2357 , n6008 );
    nor g21317 ( n20261 , n23428 , n25282 );
    nor g21318 ( n17273 , n27074 , n12208 );
    and g21319 ( n5016 , n11758 , n12457 );
    xnor g21320 ( n11830 , n3574 , n10246 );
    xnor g21321 ( n5507 , n7297 , n304 );
    xnor g21322 ( n25454 , n16667 , n3460 );
    or g21323 ( n24917 , n23974 , n26085 );
    xor g21324 ( n4791 , n25405 , n21627 );
    not g21325 ( n24115 , n11018 );
    or g21326 ( n23971 , n4815 , n22655 );
    not g21327 ( n21455 , n2055 );
    or g21328 ( n4528 , n12844 , n2158 );
    not g21329 ( n22981 , n21907 );
    xnor g21330 ( n15307 , n23079 , n16040 );
    or g21331 ( n465 , n23612 , n3906 );
    xnor g21332 ( n13116 , n13200 , n6147 );
    not g21333 ( n7096 , n17758 );
    and g21334 ( n4702 , n22752 , n16857 );
    xnor g21335 ( n12098 , n4314 , n15001 );
    xnor g21336 ( n26265 , n20030 , n337 );
    not g21337 ( n8549 , n8438 );
    nor g21338 ( n23668 , n9058 , n5925 );
    nor g21339 ( n15155 , n2902 , n19809 );
    or g21340 ( n16404 , n1358 , n12339 );
    not g21341 ( n20608 , n12289 );
    or g21342 ( n15247 , n15104 , n11123 );
    or g21343 ( n20779 , n17354 , n23265 );
    xnor g21344 ( n679 , n9090 , n19107 );
    and g21345 ( n16876 , n25105 , n10925 );
    or g21346 ( n25174 , n25682 , n15457 );
    not g21347 ( n6591 , n8730 );
    and g21348 ( n6048 , n12199 , n14712 );
    xnor g21349 ( n8810 , n4957 , n25797 );
    or g21350 ( n6598 , n11808 , n5645 );
    nor g21351 ( n18453 , n5342 , n26919 );
    or g21352 ( n6405 , n11583 , n18416 );
    or g21353 ( n12711 , n4381 , n26809 );
    or g21354 ( n2398 , n15129 , n541 );
    or g21355 ( n16777 , n20675 , n18778 );
    or g21356 ( n105 , n7142 , n3860 );
    nor g21357 ( n12876 , n14603 , n24736 );
    or g21358 ( n6113 , n16633 , n22379 );
    not g21359 ( n15536 , n21390 );
    nor g21360 ( n954 , n1099 , n6381 );
    and g21361 ( n2502 , n11273 , n23086 );
    not g21362 ( n24665 , n11479 );
    or g21363 ( n25392 , n11737 , n14274 );
    or g21364 ( n23185 , n22198 , n14424 );
    or g21365 ( n24222 , n14633 , n2886 );
    or g21366 ( n13847 , n15125 , n23587 );
    or g21367 ( n26909 , n2121 , n10625 );
    xnor g21368 ( n11860 , n767 , n8806 );
    xnor g21369 ( n13255 , n12088 , n26483 );
    or g21370 ( n26158 , n11919 , n12875 );
    or g21371 ( n16323 , n1096 , n19879 );
    not g21372 ( n25674 , n1777 );
    xnor g21373 ( n4346 , n7437 , n13367 );
    nor g21374 ( n3819 , n23353 , n14881 );
    or g21375 ( n15323 , n26677 , n21745 );
    nor g21376 ( n1335 , n8546 , n10855 );
    or g21377 ( n14234 , n8606 , n16282 );
    or g21378 ( n21591 , n18264 , n14373 );
    xnor g21379 ( n24444 , n7525 , n11900 );
    and g21380 ( n6990 , n20739 , n3864 );
    and g21381 ( n8558 , n16498 , n13342 );
    xnor g21382 ( n13993 , n12928 , n12650 );
    xnor g21383 ( n22717 , n15132 , n4614 );
    nor g21384 ( n24838 , n15655 , n12415 );
    buf g21385 ( n2194 , n13879 );
    or g21386 ( n23598 , n3945 , n3393 );
    and g21387 ( n2330 , n4256 , n20205 );
    xnor g21388 ( n18601 , n21086 , n2861 );
    not g21389 ( n7215 , n8405 );
    and g21390 ( n21560 , n19832 , n3201 );
    not g21391 ( n5916 , n5694 );
    xnor g21392 ( n21295 , n11119 , n22279 );
    nor g21393 ( n6511 , n13897 , n19515 );
    not g21394 ( n19962 , n21993 );
    not g21395 ( n1025 , n18250 );
    or g21396 ( n12220 , n8372 , n17979 );
    nor g21397 ( n25188 , n18438 , n26672 );
    not g21398 ( n3990 , n2937 );
    nor g21399 ( n10971 , n17485 , n17555 );
    xnor g21400 ( n10653 , n1303 , n4425 );
    nor g21401 ( n17118 , n2815 , n4492 );
    or g21402 ( n24944 , n3413 , n17762 );
    and g21403 ( n2424 , n11487 , n2082 );
    or g21404 ( n21783 , n15696 , n13071 );
    and g21405 ( n3055 , n1561 , n13130 );
    xnor g21406 ( n690 , n10208 , n2290 );
    or g21407 ( n4313 , n15121 , n4724 );
    or g21408 ( n24790 , n1454 , n9123 );
    not g21409 ( n15769 , n4836 );
    xnor g21410 ( n27185 , n9025 , n11032 );
    nor g21411 ( n14821 , n10135 , n24863 );
    or g21412 ( n4358 , n14404 , n25479 );
    or g21413 ( n5061 , n25318 , n3955 );
    and g21414 ( n12411 , n936 , n2584 );
    xnor g21415 ( n161 , n2359 , n25213 );
    not g21416 ( n20045 , n21649 );
    and g21417 ( n3275 , n3440 , n6028 );
    or g21418 ( n3812 , n3553 , n5116 );
    not g21419 ( n24272 , n686 );
    and g21420 ( n6180 , n24492 , n17619 );
    xnor g21421 ( n11387 , n25523 , n26318 );
    xnor g21422 ( n21980 , n17467 , n16376 );
    not g21423 ( n20841 , n4417 );
    xnor g21424 ( n15440 , n18733 , n565 );
    xnor g21425 ( n5022 , n13109 , n7731 );
    or g21426 ( n25484 , n27093 , n6056 );
    or g21427 ( n9601 , n22962 , n10567 );
    or g21428 ( n4199 , n13951 , n19388 );
    not g21429 ( n19874 , n13533 );
    xnor g21430 ( n13827 , n6847 , n2051 );
    and g21431 ( n10126 , n24651 , n27162 );
    and g21432 ( n18540 , n13964 , n26576 );
    or g21433 ( n15394 , n12442 , n12677 );
    xnor g21434 ( n13347 , n7365 , n8495 );
    not g21435 ( n5580 , n14570 );
    xnor g21436 ( n15158 , n17109 , n9686 );
    xnor g21437 ( n10202 , n25318 , n2645 );
    xnor g21438 ( n7050 , n8402 , n8589 );
    or g21439 ( n4105 , n1611 , n21763 );
    xnor g21440 ( n23782 , n4856 , n3653 );
    and g21441 ( n13393 , n926 , n14498 );
    and g21442 ( n8279 , n5623 , n13181 );
    or g21443 ( n9894 , n16331 , n5443 );
    and g21444 ( n11468 , n994 , n19503 );
    or g21445 ( n5100 , n21431 , n5529 );
    xnor g21446 ( n7313 , n25672 , n14280 );
    and g21447 ( n16814 , n7739 , n9353 );
    and g21448 ( n15791 , n11212 , n26033 );
    not g21449 ( n394 , n15169 );
    and g21450 ( n21714 , n3621 , n13002 );
    or g21451 ( n6069 , n1918 , n16653 );
    or g21452 ( n10453 , n9004 , n21014 );
    or g21453 ( n21619 , n5825 , n8788 );
    xnor g21454 ( n6250 , n16822 , n17415 );
    nor g21455 ( n16601 , n10882 , n8719 );
    or g21456 ( n3626 , n13195 , n16051 );
    xnor g21457 ( n14046 , n12797 , n26810 );
    and g21458 ( n11865 , n18171 , n24529 );
    and g21459 ( n13582 , n5151 , n3191 );
    or g21460 ( n23615 , n2960 , n1413 );
    or g21461 ( n17556 , n21804 , n22272 );
    and g21462 ( n5218 , n14281 , n8043 );
    xnor g21463 ( n8679 , n19199 , n3166 );
    not g21464 ( n546 , n20442 );
    nor g21465 ( n25897 , n14323 , n14071 );
    or g21466 ( n21403 , n6320 , n8956 );
    not g21467 ( n10375 , n17174 );
    xnor g21468 ( n861 , n3968 , n13980 );
    or g21469 ( n7073 , n19880 , n2405 );
    or g21470 ( n10005 , n20552 , n7841 );
    xnor g21471 ( n5593 , n20688 , n13421 );
    or g21472 ( n5018 , n15025 , n23080 );
    nor g21473 ( n366 , n16800 , n14678 );
    xnor g21474 ( n1731 , n11411 , n25195 );
    xnor g21475 ( n16609 , n258 , n7524 );
    xnor g21476 ( n18326 , n18457 , n9750 );
    xnor g21477 ( n22902 , n21517 , n16972 );
    and g21478 ( n25124 , n9030 , n1789 );
    not g21479 ( n15451 , n1400 );
    xnor g21480 ( n6311 , n6757 , n3400 );
    or g21481 ( n12103 , n20809 , n7560 );
    xnor g21482 ( n19366 , n10115 , n17342 );
    or g21483 ( n21102 , n18476 , n27042 );
    not g21484 ( n4320 , n25848 );
    and g21485 ( n13040 , n7170 , n19186 );
    and g21486 ( n5344 , n14013 , n19656 );
    or g21487 ( n460 , n26691 , n9496 );
    and g21488 ( n8055 , n21487 , n10749 );
    xnor g21489 ( n4374 , n24012 , n18993 );
    not g21490 ( n6319 , n18400 );
    and g21491 ( n24882 , n19007 , n25002 );
    nor g21492 ( n9777 , n9797 , n4240 );
    or g21493 ( n24413 , n16405 , n1729 );
    or g21494 ( n19788 , n7737 , n14218 );
    and g21495 ( n358 , n19054 , n13331 );
    or g21496 ( n392 , n9141 , n12533 );
    or g21497 ( n3491 , n16713 , n17497 );
    not g21498 ( n1464 , n1629 );
    xnor g21499 ( n9256 , n11428 , n5266 );
    not g21500 ( n16725 , n5197 );
    xnor g21501 ( n22144 , n25118 , n3222 );
    xnor g21502 ( n2922 , n10077 , n4651 );
    not g21503 ( n15603 , n9418 );
    not g21504 ( n13894 , n11830 );
    xnor g21505 ( n6346 , n23843 , n25505 );
    xnor g21506 ( n18685 , n10761 , n14384 );
    and g21507 ( n7033 , n19336 , n17111 );
    xnor g21508 ( n13472 , n1017 , n1011 );
    not g21509 ( n23290 , n10603 );
    and g21510 ( n12496 , n16980 , n5390 );
    nor g21511 ( n16879 , n10125 , n7619 );
    xnor g21512 ( n20087 , n10124 , n1893 );
    xnor g21513 ( n13014 , n4119 , n5255 );
    not g21514 ( n8414 , n6988 );
    or g21515 ( n26485 , n1591 , n17621 );
    xnor g21516 ( n13054 , n19031 , n21142 );
    xnor g21517 ( n10229 , n17091 , n20288 );
    xnor g21518 ( n6256 , n19837 , n19686 );
    xnor g21519 ( n15986 , n13391 , n5193 );
    not g21520 ( n6442 , n23773 );
    xnor g21521 ( n19230 , n7740 , n20429 );
    and g21522 ( n2704 , n15572 , n27143 );
    nor g21523 ( n21297 , n24116 , n1163 );
    and g21524 ( n20854 , n4327 , n27045 );
    or g21525 ( n14831 , n25494 , n10713 );
    and g21526 ( n5418 , n13420 , n19337 );
    or g21527 ( n12080 , n15847 , n24017 );
    or g21528 ( n23326 , n12125 , n21224 );
    not g21529 ( n12514 , n1855 );
    nor g21530 ( n5491 , n5376 , n6037 );
    and g21531 ( n5181 , n18921 , n1028 );
    or g21532 ( n15188 , n4623 , n373 );
    xnor g21533 ( n14124 , n19146 , n16476 );
    and g21534 ( n22035 , n6663 , n24253 );
    and g21535 ( n1914 , n2874 , n25960 );
    xnor g21536 ( n15240 , n3917 , n23503 );
    or g21537 ( n17606 , n9764 , n20082 );
    or g21538 ( n17027 , n16929 , n1708 );
    or g21539 ( n6317 , n15560 , n246 );
    and g21540 ( n20834 , n25481 , n16323 );
    and g21541 ( n23130 , n8449 , n14817 );
    or g21542 ( n9014 , n6764 , n9964 );
    nor g21543 ( n15939 , n9680 , n25360 );
    or g21544 ( n1767 , n14972 , n5354 );
    and g21545 ( n15248 , n5243 , n24961 );
    or g21546 ( n17759 , n5445 , n17497 );
    xnor g21547 ( n6021 , n2750 , n25393 );
    not g21548 ( n8261 , n21740 );
    nor g21549 ( n7810 , n16429 , n6607 );
    not g21550 ( n17727 , n1697 );
    and g21551 ( n24422 , n4938 , n10999 );
    or g21552 ( n6386 , n13190 , n15769 );
    or g21553 ( n3988 , n18798 , n4723 );
    or g21554 ( n8515 , n14887 , n4610 );
    not g21555 ( n8277 , n8889 );
    not g21556 ( n23792 , n8473 );
    or g21557 ( n17315 , n7095 , n22665 );
    not g21558 ( n3007 , n20233 );
    or g21559 ( n22046 , n5711 , n26378 );
    or g21560 ( n12706 , n23647 , n24465 );
    and g21561 ( n5441 , n5926 , n2419 );
    xnor g21562 ( n18322 , n5203 , n26048 );
    xnor g21563 ( n19435 , n9814 , n12145 );
    or g21564 ( n16599 , n3791 , n3710 );
    not g21565 ( n5067 , n16217 );
    or g21566 ( n23081 , n19652 , n22610 );
    or g21567 ( n20475 , n3731 , n6176 );
    xnor g21568 ( n1575 , n7402 , n24367 );
    not g21569 ( n6489 , n16875 );
    xnor g21570 ( n6076 , n24336 , n8986 );
    xnor g21571 ( n9377 , n16765 , n11650 );
    xnor g21572 ( n14256 , n23844 , n6328 );
    not g21573 ( n11981 , n10833 );
    xnor g21574 ( n24297 , n17463 , n7210 );
    and g21575 ( n9123 , n9484 , n18641 );
    nor g21576 ( n24065 , n19406 , n2121 );
    or g21577 ( n2458 , n17586 , n11295 );
    xnor g21578 ( n6985 , n17315 , n18489 );
    not g21579 ( n15079 , n14071 );
    or g21580 ( n19096 , n3312 , n2786 );
    and g21581 ( n13572 , n3491 , n20677 );
    and g21582 ( n7489 , n23646 , n17624 );
    or g21583 ( n11 , n1950 , n17809 );
    xnor g21584 ( n23822 , n1153 , n24242 );
    and g21585 ( n17506 , n22709 , n24895 );
    not g21586 ( n20641 , n48 );
    and g21587 ( n24291 , n18091 , n2400 );
    or g21588 ( n19637 , n24904 , n2676 );
    nor g21589 ( n11171 , n16544 , n1835 );
    or g21590 ( n25673 , n23486 , n16663 );
    and g21591 ( n1185 , n22232 , n4316 );
    and g21592 ( n2308 , n12699 , n8688 );
    nor g21593 ( n14284 , n1646 , n16638 );
    xnor g21594 ( n25170 , n16311 , n3356 );
    or g21595 ( n3876 , n14150 , n23554 );
    not g21596 ( n7974 , n8052 );
    and g21597 ( n539 , n8004 , n26485 );
    xnor g21598 ( n19111 , n4328 , n9391 );
    and g21599 ( n5910 , n22461 , n9074 );
    xnor g21600 ( n6633 , n15884 , n5211 );
    and g21601 ( n26785 , n3883 , n4991 );
    nor g21602 ( n24277 , n11048 , n3714 );
    not g21603 ( n8050 , n2366 );
    xnor g21604 ( n580 , n2988 , n14769 );
    and g21605 ( n8593 , n23437 , n16100 );
    xnor g21606 ( n16490 , n7600 , n5627 );
    xnor g21607 ( n13195 , n4534 , n10654 );
    or g21608 ( n922 , n20517 , n16744 );
    or g21609 ( n14283 , n5673 , n16146 );
    not g21610 ( n19971 , n17000 );
    or g21611 ( n5235 , n11378 , n853 );
    nor g21612 ( n13605 , n4149 , n25523 );
    xnor g21613 ( n17380 , n24557 , n26820 );
    and g21614 ( n17178 , n12404 , n7855 );
    xnor g21615 ( n26096 , n18623 , n10298 );
    xnor g21616 ( n18362 , n22373 , n25170 );
    xnor g21617 ( n26168 , n3640 , n20027 );
    nor g21618 ( n14645 , n24517 , n26327 );
    or g21619 ( n5656 , n18528 , n22544 );
    nor g21620 ( n137 , n18745 , n11976 );
    or g21621 ( n24045 , n12557 , n16489 );
    or g21622 ( n2748 , n3753 , n11438 );
    and g21623 ( n7204 , n13367 , n13074 );
    or g21624 ( n11445 , n25376 , n4040 );
    and g21625 ( n10178 , n19610 , n9159 );
    or g21626 ( n14906 , n1234 , n15994 );
    xnor g21627 ( n11737 , n4416 , n24447 );
    or g21628 ( n7154 , n8056 , n6358 );
    nor g21629 ( n3619 , n6645 , n17379 );
    and g21630 ( n2879 , n16169 , n25865 );
    and g21631 ( n5251 , n16613 , n17783 );
    nor g21632 ( n19525 , n13912 , n10684 );
    xnor g21633 ( n25245 , n1112 , n13190 );
    xnor g21634 ( n1834 , n1315 , n25635 );
    not g21635 ( n19978 , n9797 );
    or g21636 ( n18712 , n3230 , n589 );
    nor g21637 ( n2250 , n5072 , n1132 );
    xnor g21638 ( n16547 , n18016 , n647 );
    xnor g21639 ( n7861 , n26171 , n4247 );
    nor g21640 ( n8966 , n7731 , n23509 );
    or g21641 ( n24557 , n25528 , n18556 );
    xnor g21642 ( n10818 , n5205 , n6065 );
    and g21643 ( n15497 , n23732 , n17875 );
    or g21644 ( n19129 , n16822 , n5963 );
    not g21645 ( n9150 , n38 );
    or g21646 ( n6041 , n4350 , n17216 );
    xnor g21647 ( n2094 , n22517 , n19894 );
    or g21648 ( n7762 , n4878 , n15654 );
    nor g21649 ( n1954 , n20213 , n7092 );
    not g21650 ( n26912 , n7001 );
    not g21651 ( n2445 , n17261 );
    nor g21652 ( n22561 , n14563 , n23508 );
    nor g21653 ( n7051 , n655 , n5386 );
    and g21654 ( n7525 , n943 , n23811 );
    xnor g21655 ( n26709 , n14872 , n12553 );
    xnor g21656 ( n9689 , n21391 , n81 );
    nor g21657 ( n1362 , n17771 , n14762 );
    xnor g21658 ( n13973 , n16022 , n18575 );
    not g21659 ( n13789 , n24319 );
    xnor g21660 ( n10257 , n15498 , n16562 );
    or g21661 ( n23795 , n23218 , n22266 );
    nor g21662 ( n7025 , n2377 , n19633 );
    not g21663 ( n12293 , n6184 );
    not g21664 ( n446 , n16544 );
    not g21665 ( n25637 , n12605 );
    nor g21666 ( n26548 , n24301 , n2289 );
    or g21667 ( n10939 , n16480 , n17001 );
    or g21668 ( n22705 , n24595 , n17614 );
    and g21669 ( n9033 , n5152 , n2097 );
    nor g21670 ( n17717 , n20811 , n19047 );
    or g21671 ( n830 , n25872 , n19262 );
    not g21672 ( n3659 , n23754 );
    not g21673 ( n22273 , n19222 );
    not g21674 ( n808 , n11424 );
    or g21675 ( n18025 , n8534 , n24550 );
    not g21676 ( n14111 , n19236 );
    or g21677 ( n20531 , n8472 , n23318 );
    not g21678 ( n15709 , n4811 );
    or g21679 ( n5669 , n19410 , n14035 );
    xnor g21680 ( n3010 , n13866 , n3973 );
    or g21681 ( n5309 , n19150 , n25074 );
    and g21682 ( n17376 , n6260 , n18448 );
    and g21683 ( n8531 , n11992 , n11821 );
    nor g21684 ( n16607 , n13960 , n12990 );
    and g21685 ( n1665 , n5205 , n6065 );
    nor g21686 ( n26390 , n20593 , n4174 );
    nor g21687 ( n11770 , n7385 , n20241 );
    nor g21688 ( n21936 , n11936 , n2756 );
    or g21689 ( n1787 , n11585 , n5023 );
    and g21690 ( n24357 , n11774 , n7250 );
    xnor g21691 ( n19636 , n7465 , n22550 );
    not g21692 ( n10861 , n21726 );
    or g21693 ( n23227 , n19902 , n15125 );
    xnor g21694 ( n6542 , n6187 , n25641 );
    not g21695 ( n12898 , n16176 );
    and g21696 ( n17040 , n2945 , n24946 );
    and g21697 ( n13733 , n1211 , n16050 );
    and g21698 ( n20019 , n15609 , n15915 );
    and g21699 ( n18022 , n3576 , n26712 );
    and g21700 ( n14562 , n2442 , n9041 );
    or g21701 ( n25363 , n11020 , n24225 );
    and g21702 ( n26877 , n20455 , n25099 );
    or g21703 ( n18325 , n4315 , n3945 );
    xnor g21704 ( n16146 , n6166 , n22581 );
    and g21705 ( n21270 , n17607 , n16470 );
    or g21706 ( n23904 , n4359 , n10465 );
    and g21707 ( n25226 , n8494 , n20762 );
    xnor g21708 ( n2046 , n13643 , n11707 );
    and g21709 ( n19900 , n1473 , n7336 );
    not g21710 ( n14076 , n409 );
    or g21711 ( n13055 , n1439 , n13699 );
    and g21712 ( n11498 , n18907 , n13033 );
    or g21713 ( n1502 , n11745 , n10057 );
    and g21714 ( n23154 , n21320 , n23785 );
    xnor g21715 ( n10603 , n22248 , n23567 );
    or g21716 ( n15937 , n7335 , n11578 );
    xnor g21717 ( n3301 , n24017 , n10210 );
    nor g21718 ( n24348 , n11321 , n964 );
    xnor g21719 ( n3125 , n23381 , n24679 );
    and g21720 ( n308 , n21096 , n22044 );
    nor g21721 ( n15950 , n23592 , n14226 );
    xnor g21722 ( n2111 , n27029 , n27028 );
    or g21723 ( n23172 , n17187 , n17985 );
    or g21724 ( n23387 , n1951 , n27008 );
    or g21725 ( n7483 , n5280 , n19774 );
    and g21726 ( n16306 , n21611 , n14585 );
    or g21727 ( n2411 , n6692 , n10897 );
    and g21728 ( n13645 , n5820 , n24445 );
    xnor g21729 ( n7491 , n2244 , n3465 );
    and g21730 ( n20827 , n5041 , n7202 );
    nor g21731 ( n25314 , n9259 , n16401 );
    xnor g21732 ( n22266 , n23977 , n2760 );
    or g21733 ( n9295 , n2454 , n4970 );
    nor g21734 ( n25263 , n16637 , n2776 );
    xnor g21735 ( n19221 , n19782 , n3565 );
    xnor g21736 ( n4651 , n21758 , n11461 );
    and g21737 ( n1616 , n9790 , n3060 );
    or g21738 ( n6370 , n13544 , n13570 );
    not g21739 ( n24851 , n7428 );
    and g21740 ( n23492 , n14685 , n13282 );
    or g21741 ( n9173 , n15340 , n3048 );
    xnor g21742 ( n8042 , n10362 , n12498 );
    nor g21743 ( n18916 , n14465 , n7057 );
    nor g21744 ( n346 , n1055 , n12592 );
    or g21745 ( n5326 , n10184 , n6284 );
    xnor g21746 ( n1917 , n2025 , n5053 );
    or g21747 ( n5136 , n20106 , n4472 );
    xnor g21748 ( n3274 , n11819 , n6583 );
    nor g21749 ( n12557 , n16890 , n3318 );
    or g21750 ( n11059 , n7692 , n16793 );
    xnor g21751 ( n1690 , n7394 , n5579 );
    nor g21752 ( n6578 , n16127 , n18918 );
    and g21753 ( n2459 , n3460 , n24774 );
    nor g21754 ( n20821 , n5065 , n12018 );
    or g21755 ( n4795 , n7101 , n6990 );
    or g21756 ( n14568 , n9592 , n19860 );
    xnor g21757 ( n23829 , n1078 , n13170 );
    not g21758 ( n11198 , n21778 );
    or g21759 ( n24179 , n6859 , n17600 );
    or g21760 ( n4475 , n9725 , n19526 );
    xnor g21761 ( n7588 , n18716 , n26025 );
    or g21762 ( n16315 , n11075 , n5858 );
    and g21763 ( n13522 , n12159 , n23078 );
    xnor g21764 ( n21693 , n6820 , n24278 );
    xnor g21765 ( n24837 , n3354 , n12078 );
    xnor g21766 ( n19930 , n17807 , n8065 );
    xnor g21767 ( n11105 , n21674 , n22597 );
    xnor g21768 ( n9996 , n10684 , n13912 );
    and g21769 ( n9876 , n11526 , n15199 );
    and g21770 ( n853 , n15937 , n3704 );
    or g21771 ( n12170 , n10317 , n23928 );
    nor g21772 ( n793 , n5145 , n3675 );
    not g21773 ( n11714 , n23873 );
    xnor g21774 ( n6897 , n22325 , n25940 );
    xnor g21775 ( n17681 , n25781 , n9469 );
    xnor g21776 ( n20963 , n22610 , n19652 );
    nor g21777 ( n12448 , n20079 , n11406 );
    xnor g21778 ( n1016 , n10015 , n16262 );
    or g21779 ( n22967 , n11633 , n14178 );
    or g21780 ( n26440 , n25199 , n13955 );
    and g21781 ( n11214 , n16081 , n21135 );
    xnor g21782 ( n21300 , n15320 , n245 );
    and g21783 ( n26165 , n22837 , n18033 );
    not g21784 ( n24507 , n25681 );
    xnor g21785 ( n906 , n26066 , n6356 );
    xnor g21786 ( n19698 , n10763 , n12657 );
    xnor g21787 ( n14981 , n22067 , n10516 );
    xnor g21788 ( n21143 , n15459 , n10585 );
    not g21789 ( n12638 , n21165 );
    xnor g21790 ( n8453 , n2980 , n20601 );
    nor g21791 ( n17475 , n23705 , n1759 );
    or g21792 ( n24026 , n8599 , n10954 );
    xnor g21793 ( n17344 , n16172 , n21233 );
    or g21794 ( n26941 , n2725 , n6389 );
    and g21795 ( n5845 , n14435 , n1666 );
    xnor g21796 ( n21390 , n21348 , n21586 );
    not g21797 ( n27025 , n14354 );
    and g21798 ( n12539 , n5148 , n15412 );
    or g21799 ( n22188 , n10495 , n8942 );
    and g21800 ( n19013 , n4681 , n22037 );
    xnor g21801 ( n25490 , n7401 , n15964 );
    xnor g21802 ( n16714 , n17444 , n27037 );
    not g21803 ( n26295 , n15625 );
    or g21804 ( n24377 , n17173 , n4468 );
    xnor g21805 ( n18998 , n24134 , n5095 );
    or g21806 ( n9719 , n1657 , n21672 );
    and g21807 ( n25428 , n24699 , n17406 );
    nor g21808 ( n9112 , n25621 , n6930 );
    and g21809 ( n5027 , n21519 , n25709 );
    or g21810 ( n3388 , n15883 , n14381 );
    or g21811 ( n9941 , n16178 , n3955 );
    and g21812 ( n8428 , n14487 , n27022 );
    xnor g21813 ( n7976 , n2482 , n7448 );
    xnor g21814 ( n20103 , n25269 , n24368 );
    and g21815 ( n21888 , n11056 , n10181 );
    xnor g21816 ( n6339 , n7663 , n12790 );
    and g21817 ( n4491 , n16569 , n19189 );
    and g21818 ( n10916 , n23304 , n17069 );
    not g21819 ( n1997 , n4042 );
    and g21820 ( n3071 , n9560 , n14608 );
    not g21821 ( n24832 , n19762 );
    and g21822 ( n2062 , n24557 , n15630 );
    and g21823 ( n15612 , n12492 , n21594 );
    xnor g21824 ( n6474 , n5998 , n12384 );
    xnor g21825 ( n23990 , n7510 , n13438 );
    xnor g21826 ( n16929 , n3585 , n6207 );
    or g21827 ( n23127 , n19452 , n3527 );
    or g21828 ( n12782 , n14803 , n1115 );
    xnor g21829 ( n2657 , n10988 , n3669 );
    xnor g21830 ( n24472 , n10163 , n20458 );
    or g21831 ( n19906 , n11668 , n7332 );
    or g21832 ( n19188 , n10958 , n19580 );
    nor g21833 ( n976 , n14388 , n21575 );
    xnor g21834 ( n10582 , n1421 , n15378 );
    nor g21835 ( n24324 , n27075 , n16239 );
    xnor g21836 ( n7838 , n23456 , n8964 );
    not g21837 ( n2908 , n14762 );
    not g21838 ( n27111 , n12713 );
    or g21839 ( n4470 , n10892 , n419 );
    nor g21840 ( n23269 , n17847 , n11394 );
    or g21841 ( n7624 , n16515 , n9824 );
    nor g21842 ( n5384 , n3276 , n2547 );
    xnor g21843 ( n15903 , n26576 , n5636 );
    and g21844 ( n18384 , n25797 , n15784 );
    xnor g21845 ( n19420 , n9455 , n18290 );
    xnor g21846 ( n23680 , n10577 , n3279 );
    not g21847 ( n7546 , n27046 );
    and g21848 ( n24061 , n4662 , n25091 );
    xnor g21849 ( n159 , n19683 , n24048 );
    or g21850 ( n5726 , n13277 , n19869 );
    or g21851 ( n7248 , n23943 , n18723 );
    or g21852 ( n4726 , n3248 , n11568 );
    xnor g21853 ( n9521 , n19377 , n17780 );
    nor g21854 ( n7232 , n10631 , n9125 );
    and g21855 ( n9161 , n20348 , n9724 );
    xnor g21856 ( n18252 , n7991 , n3133 );
    not g21857 ( n3498 , n8974 );
    nor g21858 ( n24849 , n22755 , n310 );
    xnor g21859 ( n9240 , n22108 , n22626 );
    and g21860 ( n22075 , n17282 , n169 );
    not g21861 ( n18797 , n9827 );
    and g21862 ( n18224 , n5355 , n17659 );
    xnor g21863 ( n15807 , n439 , n16304 );
    not g21864 ( n16697 , n22006 );
    or g21865 ( n4251 , n4270 , n4438 );
    or g21866 ( n18176 , n24654 , n22340 );
    xnor g21867 ( n11213 , n20196 , n25872 );
    xnor g21868 ( n17160 , n26270 , n19495 );
    or g21869 ( n8854 , n26086 , n7149 );
    xnor g21870 ( n15719 , n21043 , n25963 );
    xnor g21871 ( n10903 , n14109 , n12357 );
    not g21872 ( n26066 , n4067 );
    nor g21873 ( n19567 , n22375 , n24815 );
    and g21874 ( n21523 , n5119 , n6070 );
    or g21875 ( n13900 , n13534 , n15500 );
    or g21876 ( n7357 , n3840 , n24908 );
    xnor g21877 ( n16860 , n25164 , n16490 );
    and g21878 ( n6176 , n25284 , n17823 );
    and g21879 ( n20675 , n19754 , n11308 );
    or g21880 ( n1270 , n9770 , n25676 );
    or g21881 ( n18834 , n614 , n19075 );
    and g21882 ( n2530 , n17532 , n1334 );
    or g21883 ( n17304 , n14007 , n23144 );
    xnor g21884 ( n11241 , n557 , n19390 );
    xnor g21885 ( n3166 , n19914 , n23895 );
    and g21886 ( n10835 , n16812 , n24402 );
    xnor g21887 ( n17866 , n24638 , n19327 );
    not g21888 ( n22254 , n3570 );
    or g21889 ( n26973 , n12058 , n285 );
    xnor g21890 ( n11326 , n8730 , n6130 );
    or g21891 ( n5566 , n4278 , n15074 );
    or g21892 ( n449 , n7676 , n9380 );
    nor g21893 ( n16944 , n19471 , n11491 );
    or g21894 ( n17631 , n5400 , n3149 );
    xnor g21895 ( n4917 , n20381 , n17218 );
    nor g21896 ( n17939 , n985 , n19218 );
    or g21897 ( n23194 , n26746 , n2224 );
    xnor g21898 ( n26076 , n8295 , n13037 );
    or g21899 ( n1920 , n14785 , n480 );
    not g21900 ( n3317 , n27181 );
    xnor g21901 ( n1855 , n16725 , n11973 );
    xnor g21902 ( n22542 , n14510 , n21649 );
    or g21903 ( n10052 , n3417 , n12986 );
    not g21904 ( n26312 , n8614 );
    xnor g21905 ( n5162 , n8472 , n6150 );
    or g21906 ( n17399 , n504 , n26135 );
    and g21907 ( n6438 , n16743 , n24081 );
    and g21908 ( n26618 , n26611 , n4235 );
    or g21909 ( n892 , n24081 , n16743 );
    and g21910 ( n10764 , n7203 , n3989 );
    nor g21911 ( n10123 , n1009 , n1293 );
    xnor g21912 ( n2880 , n2328 , n18274 );
    nor g21913 ( n17799 , n24417 , n11363 );
    nor g21914 ( n6306 , n19106 , n24879 );
    not g21915 ( n17454 , n1418 );
    not g21916 ( n17953 , n11116 );
    or g21917 ( n17434 , n7030 , n23752 );
    not g21918 ( n25936 , n16476 );
    xnor g21919 ( n7369 , n22820 , n7693 );
    xnor g21920 ( n11348 , n2047 , n19485 );
    and g21921 ( n17573 , n25134 , n10865 );
    xnor g21922 ( n5439 , n17970 , n14324 );
    or g21923 ( n14177 , n15463 , n13820 );
    or g21924 ( n20547 , n17992 , n25137 );
    xnor g21925 ( n2076 , n16924 , n10984 );
    and g21926 ( n7385 , n25483 , n1062 );
    or g21927 ( n8723 , n1912 , n1160 );
    not g21928 ( n5066 , n820 );
    or g21929 ( n2962 , n19084 , n28 );
    not g21930 ( n7198 , n14680 );
    and g21931 ( n11677 , n4628 , n21769 );
    nor g21932 ( n22745 , n20192 , n12481 );
    or g21933 ( n6441 , n16380 , n886 );
    not g21934 ( n25393 , n2023 );
    nor g21935 ( n10248 , n22585 , n20986 );
    not g21936 ( n23580 , n22215 );
    or g21937 ( n20878 , n14293 , n2914 );
    not g21938 ( n2787 , n12993 );
    and g21939 ( n511 , n14026 , n15853 );
    or g21940 ( n124 , n609 , n18070 );
    not g21941 ( n22865 , n13489 );
    or g21942 ( n26818 , n25029 , n10089 );
    or g21943 ( n7602 , n24031 , n25261 );
    and g21944 ( n20699 , n22102 , n3560 );
    xnor g21945 ( n5075 , n13062 , n21230 );
    or g21946 ( n24087 , n23202 , n10813 );
    or g21947 ( n7037 , n1191 , n14513 );
    not g21948 ( n16873 , n5751 );
    xnor g21949 ( n7181 , n20925 , n23791 );
    xnor g21950 ( n1684 , n3883 , n18225 );
    xnor g21951 ( n7873 , n8856 , n4319 );
    or g21952 ( n24113 , n18669 , n13891 );
    xnor g21953 ( n17427 , n11428 , n1181 );
    xnor g21954 ( n24835 , n25294 , n22474 );
    not g21955 ( n14974 , n21309 );
    or g21956 ( n5009 , n17660 , n26520 );
    or g21957 ( n19012 , n10116 , n20485 );
    not g21958 ( n8795 , n19111 );
    or g21959 ( n19413 , n2321 , n11950 );
    xnor g21960 ( n9143 , n8531 , n5731 );
    or g21961 ( n24140 , n25939 , n26947 );
    or g21962 ( n19253 , n10940 , n1362 );
    and g21963 ( n21188 , n13460 , n5156 );
    and g21964 ( n9328 , n8412 , n12200 );
    not g21965 ( n14152 , n18478 );
    nor g21966 ( n3091 , n17835 , n8166 );
    nor g21967 ( n26746 , n15918 , n21735 );
    not g21968 ( n14936 , n27188 );
    nor g21969 ( n25347 , n15979 , n15008 );
    and g21970 ( n7441 , n15391 , n20816 );
    and g21971 ( n23937 , n13912 , n11098 );
    xnor g21972 ( n13262 , n18369 , n21319 );
    and g21973 ( n7400 , n2822 , n13090 );
    and g21974 ( n20637 , n7301 , n26115 );
    nor g21975 ( n15461 , n7734 , n5163 );
    nor g21976 ( n24370 , n4859 , n5140 );
    not g21977 ( n16738 , n23752 );
    not g21978 ( n21412 , n11838 );
    xnor g21979 ( n11461 , n15998 , n5142 );
    xnor g21980 ( n6162 , n12875 , n26318 );
    nor g21981 ( n699 , n17647 , n20146 );
    or g21982 ( n8275 , n16427 , n1807 );
    not g21983 ( n25066 , n26142 );
    xnor g21984 ( n2630 , n5673 , n19337 );
    and g21985 ( n23340 , n22839 , n21419 );
    nor g21986 ( n5883 , n5793 , n2782 );
    xnor g21987 ( n2992 , n14152 , n25987 );
    xnor g21988 ( n13291 , n26336 , n3264 );
    or g21989 ( n22668 , n12893 , n2463 );
    and g21990 ( n4283 , n4593 , n7694 );
    xor g21991 ( n26917 , n13918 , n26462 );
    or g21992 ( n18155 , n15696 , n18800 );
    xnor g21993 ( n610 , n13783 , n22332 );
    or g21994 ( n8561 , n12149 , n1915 );
    not g21995 ( n24551 , n4734 );
    xnor g21996 ( n14223 , n16547 , n12900 );
    xnor g21997 ( n26195 , n18558 , n6556 );
    xnor g21998 ( n11564 , n26802 , n22172 );
    xnor g21999 ( n18307 , n20512 , n25726 );
    and g22000 ( n27058 , n15729 , n24831 );
    or g22001 ( n19067 , n18078 , n12543 );
    and g22002 ( n9229 , n14660 , n14929 );
    not g22003 ( n11963 , n20411 );
    or g22004 ( n9066 , n3672 , n14886 );
    and g22005 ( n7401 , n10559 , n10182 );
    and g22006 ( n2136 , n11065 , n23334 );
    xnor g22007 ( n3479 , n1018 , n25808 );
    or g22008 ( n17034 , n10374 , n22389 );
    and g22009 ( n12661 , n9121 , n25343 );
    xnor g22010 ( n20279 , n5433 , n8807 );
    and g22011 ( n23947 , n9739 , n4262 );
    or g22012 ( n3920 , n15224 , n8877 );
    and g22013 ( n26060 , n7796 , n13878 );
    and g22014 ( n21961 , n16929 , n1708 );
    and g22015 ( n17935 , n20357 , n998 );
    xnor g22016 ( n2147 , n3212 , n16251 );
    or g22017 ( n26712 , n25553 , n2882 );
    or g22018 ( n17329 , n12218 , n26637 );
    or g22019 ( n5032 , n18353 , n24206 );
    or g22020 ( n9315 , n3636 , n24889 );
    or g22021 ( n16977 , n13575 , n19305 );
    and g22022 ( n9962 , n3108 , n13805 );
    xnor g22023 ( n4766 , n10186 , n1539 );
    or g22024 ( n5005 , n6353 , n12391 );
    or g22025 ( n25732 , n9297 , n2767 );
    or g22026 ( n5467 , n6032 , n15596 );
    and g22027 ( n20262 , n6605 , n20322 );
    and g22028 ( n8190 , n26526 , n7135 );
    or g22029 ( n10959 , n15034 , n19408 );
    and g22030 ( n731 , n24938 , n21618 );
    xnor g22031 ( n20669 , n26986 , n3425 );
    nor g22032 ( n5684 , n24902 , n8623 );
    or g22033 ( n2120 , n11155 , n972 );
    or g22034 ( n23003 , n13306 , n7525 );
    xnor g22035 ( n12226 , n12592 , n1055 );
    or g22036 ( n11199 , n2058 , n10112 );
    or g22037 ( n7866 , n2169 , n7393 );
    nor g22038 ( n17446 , n19895 , n14311 );
    or g22039 ( n6151 , n53 , n18197 );
    xnor g22040 ( n26867 , n13708 , n24618 );
    or g22041 ( n1878 , n3335 , n8057 );
    not g22042 ( n455 , n14463 );
    and g22043 ( n13520 , n17393 , n18457 );
    and g22044 ( n21530 , n18180 , n5861 );
    xnor g22045 ( n13548 , n6806 , n2065 );
    xnor g22046 ( n11510 , n13651 , n20727 );
    or g22047 ( n18942 , n3083 , n1564 );
    nor g22048 ( n23274 , n18995 , n19357 );
    xnor g22049 ( n1700 , n6434 , n25956 );
    and g22050 ( n14664 , n23108 , n17604 );
    and g22051 ( n19821 , n21499 , n25753 );
    or g22052 ( n1975 , n2868 , n881 );
    and g22053 ( n23311 , n24828 , n19368 );
    or g22054 ( n5869 , n25436 , n8395 );
    xnor g22055 ( n17277 , n25401 , n391 );
    xnor g22056 ( n18863 , n26789 , n342 );
    not g22057 ( n20160 , n23889 );
    or g22058 ( n10715 , n7652 , n18826 );
    or g22059 ( n24983 , n26363 , n22047 );
    and g22060 ( n2505 , n10947 , n23354 );
    xnor g22061 ( n20530 , n26792 , n21584 );
    and g22062 ( n7978 , n9918 , n15420 );
    or g22063 ( n12168 , n10712 , n14467 );
    xnor g22064 ( n18061 , n14817 , n13560 );
    nor g22065 ( n14708 , n2568 , n13625 );
    xnor g22066 ( n3478 , n7439 , n3984 );
    and g22067 ( n4357 , n11233 , n1990 );
    xnor g22068 ( n6334 , n966 , n8687 );
    xnor g22069 ( n21816 , n19974 , n23435 );
    or g22070 ( n18285 , n26550 , n4768 );
    not g22071 ( n10966 , n15424 );
    or g22072 ( n4639 , n10826 , n16381 );
    xnor g22073 ( n18438 , n12415 , n16984 );
    not g22074 ( n23254 , n19432 );
    xnor g22075 ( n7235 , n18046 , n14969 );
    or g22076 ( n22922 , n3305 , n6538 );
    nor g22077 ( n17100 , n7305 , n25538 );
    nor g22078 ( n22134 , n24196 , n22049 );
    xnor g22079 ( n21670 , n9832 , n6513 );
    or g22080 ( n12781 , n15658 , n1312 );
    and g22081 ( n11853 , n24822 , n2772 );
    xnor g22082 ( n24491 , n8194 , n24093 );
    not g22083 ( n5960 , n10739 );
    xnor g22084 ( n12723 , n15135 , n25712 );
    xnor g22085 ( n17947 , n8540 , n2146 );
    nor g22086 ( n12053 , n14528 , n6713 );
    xnor g22087 ( n26719 , n8393 , n11298 );
    not g22088 ( n1839 , n26141 );
    or g22089 ( n26455 , n12847 , n2255 );
    nor g22090 ( n1811 , n24475 , n19568 );
    nor g22091 ( n18659 , n1960 , n18749 );
    and g22092 ( n5149 , n11435 , n25670 );
    or g22093 ( n11292 , n3284 , n2041 );
    not g22094 ( n17779 , n2586 );
    and g22095 ( n21076 , n6312 , n27083 );
    xnor g22096 ( n8299 , n25312 , n9206 );
    and g22097 ( n1477 , n4801 , n9723 );
    xnor g22098 ( n16681 , n3298 , n26443 );
    nor g22099 ( n13102 , n10378 , n2312 );
    xnor g22100 ( n12939 , n10031 , n23578 );
    xnor g22101 ( n11224 , n17211 , n20054 );
    and g22102 ( n22875 , n23158 , n10880 );
    xnor g22103 ( n22568 , n22613 , n22631 );
    xnor g22104 ( n19220 , n3115 , n4523 );
    xnor g22105 ( n24418 , n17444 , n19652 );
    nor g22106 ( n11238 , n1136 , n11667 );
    not g22107 ( n17211 , n25498 );
    xnor g22108 ( n12102 , n8344 , n16217 );
    and g22109 ( n16156 , n4760 , n24711 );
    xnor g22110 ( n17829 , n3161 , n21134 );
    or g22111 ( n11465 , n19 , n26913 );
    and g22112 ( n16946 , n24987 , n15584 );
    xnor g22113 ( n3809 , n2158 , n13830 );
    and g22114 ( n23786 , n21021 , n18355 );
    not g22115 ( n7170 , n20446 );
    xnor g22116 ( n2828 , n6341 , n13783 );
    or g22117 ( n18603 , n25008 , n6501 );
    nor g22118 ( n24405 , n9519 , n22330 );
    xnor g22119 ( n3616 , n14033 , n22554 );
    or g22120 ( n11906 , n26530 , n25465 );
    not g22121 ( n16633 , n767 );
    xnor g22122 ( n16801 , n13186 , n11611 );
    xnor g22123 ( n11996 , n18579 , n2177 );
    or g22124 ( n25266 , n24892 , n8859 );
    or g22125 ( n15102 , n10602 , n10984 );
    not g22126 ( n13379 , n16526 );
    or g22127 ( n24430 , n9673 , n13799 );
    or g22128 ( n15718 , n9115 , n15461 );
    xnor g22129 ( n11843 , n8172 , n9086 );
    nor g22130 ( n5317 , n23373 , n16732 );
    not g22131 ( n23085 , n10179 );
    xnor g22132 ( n13372 , n7311 , n25023 );
    nor g22133 ( n3083 , n19589 , n8935 );
    xnor g22134 ( n14095 , n850 , n6585 );
    and g22135 ( n4267 , n26502 , n23332 );
    nor g22136 ( n10881 , n24969 , n26544 );
    not g22137 ( n23152 , n5969 );
    xnor g22138 ( n24529 , n10179 , n13708 );
    or g22139 ( n17422 , n10425 , n18337 );
    not g22140 ( n25318 , n1835 );
    and g22141 ( n16078 , n17547 , n15524 );
    nor g22142 ( n19830 , n14684 , n17360 );
    or g22143 ( n22147 , n15240 , n14111 );
    nor g22144 ( n21566 , n4602 , n12402 );
    not g22145 ( n15189 , n8256 );
    xnor g22146 ( n8881 , n6656 , n9787 );
    xnor g22147 ( n15333 , n12759 , n26192 );
    and g22148 ( n20082 , n3269 , n26843 );
    nor g22149 ( n21148 , n27104 , n9114 );
    or g22150 ( n9746 , n19644 , n25552 );
    not g22151 ( n20378 , n3918 );
    xnor g22152 ( n9164 , n13913 , n5357 );
    xnor g22153 ( n10851 , n3342 , n11866 );
    or g22154 ( n2427 , n1553 , n13774 );
    and g22155 ( n25137 , n22890 , n23041 );
    nor g22156 ( n2369 , n22077 , n26351 );
    not g22157 ( n7452 , n23513 );
    or g22158 ( n2245 , n9958 , n16538 );
    and g22159 ( n14494 , n26850 , n213 );
    or g22160 ( n23713 , n7747 , n9331 );
    and g22161 ( n2321 , n4304 , n23876 );
    xnor g22162 ( n5847 , n20077 , n6794 );
    nor g22163 ( n24924 , n10096 , n24511 );
    nor g22164 ( n2590 , n24493 , n19200 );
    or g22165 ( n6548 , n26613 , n4771 );
    xnor g22166 ( n22697 , n1126 , n7420 );
    not g22167 ( n2089 , n24586 );
    or g22168 ( n26305 , n14195 , n19874 );
    xnor g22169 ( n3934 , n17580 , n9760 );
    nor g22170 ( n19668 , n8943 , n10919 );
    xnor g22171 ( n12942 , n26589 , n4647 );
    xnor g22172 ( n4435 , n12678 , n2700 );
    nor g22173 ( n25408 , n12002 , n16890 );
    or g22174 ( n1529 , n25257 , n24132 );
    xnor g22175 ( n4092 , n3472 , n10477 );
    or g22176 ( n16930 , n14189 , n14795 );
    nor g22177 ( n5371 , n25322 , n23329 );
    or g22178 ( n15235 , n2389 , n20233 );
    xnor g22179 ( n14081 , n7044 , n6302 );
    nor g22180 ( n8202 , n15415 , n12875 );
    or g22181 ( n3818 , n3606 , n24643 );
    not g22182 ( n7417 , n1243 );
    not g22183 ( n13154 , n9493 );
    or g22184 ( n11961 , n319 , n23032 );
    xnor g22185 ( n17193 , n22626 , n26986 );
    xnor g22186 ( n23647 , n22525 , n6121 );
    xnor g22187 ( n13735 , n115 , n22859 );
    xnor g22188 ( n9993 , n23477 , n21398 );
    and g22189 ( n10552 , n16029 , n12088 );
    or g22190 ( n3394 , n25882 , n19078 );
    or g22191 ( n18567 , n7444 , n17076 );
    not g22192 ( n23678 , n13354 );
    or g22193 ( n24369 , n6259 , n14838 );
    xnor g22194 ( n17969 , n4722 , n14323 );
    xnor g22195 ( n16324 , n25842 , n13736 );
    or g22196 ( n15296 , n18794 , n16038 );
    or g22197 ( n1805 , n25629 , n2291 );
    or g22198 ( n10515 , n3327 , n13120 );
    xnor g22199 ( n25083 , n24149 , n15965 );
    or g22200 ( n11781 , n12511 , n4590 );
    and g22201 ( n11247 , n25319 , n11250 );
    and g22202 ( n761 , n20701 , n4447 );
    xnor g22203 ( n10669 , n5411 , n6729 );
    nor g22204 ( n8909 , n1610 , n1500 );
    or g22205 ( n12031 , n17826 , n13033 );
    and g22206 ( n869 , n16722 , n2230 );
    not g22207 ( n6789 , n5424 );
    and g22208 ( n1534 , n2995 , n15678 );
    or g22209 ( n3523 , n19547 , n12781 );
    nor g22210 ( n5511 , n6352 , n424 );
    nor g22211 ( n1461 , n3228 , n6082 );
    and g22212 ( n12305 , n11921 , n1324 );
    xnor g22213 ( n10817 , n2717 , n5259 );
    and g22214 ( n14670 , n25941 , n13958 );
    or g22215 ( n13790 , n16211 , n2289 );
    xnor g22216 ( n6257 , n15132 , n23514 );
    and g22217 ( n15660 , n3253 , n21021 );
    not g22218 ( n8431 , n24744 );
    xnor g22219 ( n2608 , n3723 , n16823 );
    nor g22220 ( n4815 , n16572 , n22012 );
    or g22221 ( n1294 , n812 , n15498 );
    or g22222 ( n17005 , n9196 , n13731 );
    or g22223 ( n16238 , n7331 , n4356 );
    xnor g22224 ( n14779 , n18765 , n22626 );
    or g22225 ( n15638 , n9693 , n10767 );
    xnor g22226 ( n13567 , n15486 , n11149 );
    xnor g22227 ( n10858 , n25637 , n27100 );
    buf g22228 ( n5793 , n4616 );
    not g22229 ( n15500 , n3641 );
    or g22230 ( n10925 , n25933 , n1323 );
    or g22231 ( n19065 , n17208 , n12182 );
    and g22232 ( n22296 , n653 , n13883 );
    or g22233 ( n15865 , n21662 , n7568 );
    or g22234 ( n16342 , n6547 , n4611 );
    xnor g22235 ( n10352 , n26397 , n13179 );
    xnor g22236 ( n17630 , n19565 , n10867 );
    and g22237 ( n13479 , n17990 , n7037 );
    xnor g22238 ( n16493 , n27177 , n12005 );
    nor g22239 ( n15071 , n17584 , n19282 );
    not g22240 ( n5949 , n25966 );
    and g22241 ( n3194 , n23662 , n22512 );
    not g22242 ( n8457 , n7274 );
    and g22243 ( n23358 , n11766 , n9530 );
    xnor g22244 ( n9302 , n7963 , n12161 );
    or g22245 ( n875 , n7423 , n156 );
    not g22246 ( n20342 , n17458 );
    nor g22247 ( n353 , n24714 , n22501 );
    or g22248 ( n18922 , n1587 , n1685 );
    xnor g22249 ( n16275 , n9604 , n16174 );
    xnor g22250 ( n3556 , n11485 , n19147 );
    or g22251 ( n20781 , n15133 , n4289 );
    and g22252 ( n953 , n21794 , n10332 );
    xnor g22253 ( n19187 , n7177 , n21828 );
    and g22254 ( n17063 , n8416 , n101 );
    nor g22255 ( n11031 , n20138 , n25073 );
    not g22256 ( n1934 , n13562 );
    or g22257 ( n11836 , n6451 , n10988 );
    and g22258 ( n24168 , n3805 , n24159 );
    xnor g22259 ( n23969 , n5111 , n4514 );
    or g22260 ( n11422 , n17642 , n26256 );
    not g22261 ( n8514 , n26080 );
    and g22262 ( n15315 , n4859 , n9793 );
    or g22263 ( n17609 , n14818 , n17532 );
    or g22264 ( n26366 , n18183 , n18466 );
    or g22265 ( n8559 , n19938 , n11623 );
    not g22266 ( n524 , n7693 );
    or g22267 ( n17086 , n22754 , n13569 );
    xnor g22268 ( n9308 , n5444 , n8756 );
    or g22269 ( n21331 , n20312 , n19567 );
    not g22270 ( n5604 , n14899 );
    xnor g22271 ( n7323 , n3379 , n1099 );
    or g22272 ( n24190 , n17272 , n13929 );
    xnor g22273 ( n17555 , n127 , n273 );
    xnor g22274 ( n19482 , n26556 , n12495 );
    and g22275 ( n10613 , n4101 , n16435 );
    nor g22276 ( n25721 , n19469 , n20235 );
    not g22277 ( n16830 , n27104 );
    or g22278 ( n26275 , n25959 , n20392 );
    not g22279 ( n24727 , n4277 );
    or g22280 ( n19475 , n7436 , n4606 );
    xnor g22281 ( n13115 , n715 , n9591 );
    or g22282 ( n18684 , n21016 , n7966 );
    xnor g22283 ( n6125 , n11841 , n19701 );
    not g22284 ( n16882 , n8441 );
    not g22285 ( n8322 , n5213 );
    nor g22286 ( n15841 , n4426 , n25246 );
    or g22287 ( n6926 , n14789 , n3790 );
    or g22288 ( n14743 , n11854 , n19807 );
    or g22289 ( n7128 , n3634 , n9263 );
    or g22290 ( n14166 , n22730 , n8235 );
    and g22291 ( n15056 , n14830 , n6468 );
    and g22292 ( n21466 , n16985 , n8833 );
    and g22293 ( n14317 , n14133 , n7293 );
    xnor g22294 ( n4139 , n25739 , n8419 );
    xnor g22295 ( n12252 , n7334 , n20961 );
    and g22296 ( n5201 , n11898 , n25063 );
    xnor g22297 ( n327 , n23898 , n15182 );
    not g22298 ( n24479 , n8437 );
    not g22299 ( n11060 , n12020 );
    not g22300 ( n19610 , n16818 );
    xnor g22301 ( n17430 , n21362 , n25812 );
    xnor g22302 ( n16201 , n20390 , n12842 );
    or g22303 ( n9008 , n5461 , n20529 );
    xnor g22304 ( n25164 , n23563 , n24979 );
    xnor g22305 ( n20661 , n594 , n9199 );
    or g22306 ( n20573 , n17831 , n15475 );
    or g22307 ( n22524 , n442 , n6319 );
    or g22308 ( n4190 , n7689 , n22600 );
    xnor g22309 ( n24600 , n9701 , n19431 );
    nor g22310 ( n22240 , n14907 , n26522 );
    or g22311 ( n23887 , n14818 , n26491 );
    xnor g22312 ( n31 , n24305 , n2580 );
    xnor g22313 ( n10326 , n7199 , n10386 );
    or g22314 ( n11057 , n21643 , n101 );
    or g22315 ( n25095 , n14886 , n17639 );
    or g22316 ( n21296 , n2556 , n8893 );
    nor g22317 ( n6638 , n22198 , n5337 );
    nor g22318 ( n24942 , n16713 , n15808 );
    nor g22319 ( n20725 , n14272 , n1929 );
    nor g22320 ( n14814 , n9108 , n530 );
    or g22321 ( n14179 , n17385 , n27073 );
    xnor g22322 ( n14666 , n3324 , n16544 );
    not g22323 ( n23451 , n5795 );
    or g22324 ( n6740 , n23274 , n23689 );
    or g22325 ( n21741 , n658 , n25339 );
    xnor g22326 ( n21000 , n9373 , n7677 );
    or g22327 ( n20586 , n420 , n12535 );
    and g22328 ( n22785 , n19353 , n6784 );
    or g22329 ( n6447 , n8150 , n1328 );
    or g22330 ( n12604 , n6691 , n19222 );
    or g22331 ( n8177 , n2967 , n7099 );
    not g22332 ( n507 , n3673 );
    or g22333 ( n14108 , n13999 , n14376 );
    nor g22334 ( n12688 , n1654 , n4256 );
    and g22335 ( n15893 , n22991 , n467 );
    and g22336 ( n4381 , n14923 , n12050 );
    and g22337 ( n5551 , n16096 , n6952 );
    and g22338 ( n319 , n5091 , n9743 );
    and g22339 ( n14438 , n6691 , n21753 );
    or g22340 ( n17786 , n12287 , n20299 );
    not g22341 ( n16178 , n8182 );
    xnor g22342 ( n25632 , n11144 , n25500 );
    xnor g22343 ( n26126 , n22031 , n20824 );
    not g22344 ( n9395 , n21195 );
    or g22345 ( n10953 , n7548 , n9339 );
    not g22346 ( n23837 , n21778 );
    or g22347 ( n8062 , n22845 , n1655 );
    xnor g22348 ( n6388 , n23160 , n3570 );
    and g22349 ( n13810 , n8713 , n6071 );
    xnor g22350 ( n11844 , n15546 , n14702 );
    and g22351 ( n22086 , n24748 , n16170 );
    or g22352 ( n21075 , n6291 , n5693 );
    or g22353 ( n3213 , n25435 , n19527 );
    xnor g22354 ( n9919 , n5716 , n10280 );
    xnor g22355 ( n16484 , n23268 , n15282 );
    nor g22356 ( n13508 , n18891 , n14078 );
    not g22357 ( n3890 , n19575 );
    xnor g22358 ( n17723 , n21317 , n19196 );
    not g22359 ( n16401 , n21577 );
    and g22360 ( n19536 , n3855 , n1193 );
    or g22361 ( n12027 , n3907 , n16586 );
    or g22362 ( n3680 , n21271 , n15772 );
    not g22363 ( n25142 , n20455 );
    or g22364 ( n13210 , n16789 , n10962 );
    not g22365 ( n6193 , n26483 );
    xnor g22366 ( n14827 , n8919 , n5819 );
    nor g22367 ( n6096 , n3967 , n27054 );
    or g22368 ( n7228 , n10181 , n5796 );
    or g22369 ( n6236 , n7566 , n2389 );
    not g22370 ( n18527 , n17854 );
    xnor g22371 ( n1590 , n4109 , n12827 );
    nor g22372 ( n19050 , n18046 , n1025 );
    not g22373 ( n10847 , n5171 );
    or g22374 ( n12243 , n12666 , n7218 );
    or g22375 ( n23635 , n24158 , n24785 );
    xnor g22376 ( n14927 , n20359 , n25240 );
    or g22377 ( n23759 , n13559 , n4250 );
    and g22378 ( n4249 , n22100 , n23482 );
    xnor g22379 ( n5470 , n23631 , n3365 );
    not g22380 ( n4767 , n25076 );
    and g22381 ( n1085 , n9055 , n21990 );
    not g22382 ( n3443 , n1309 );
    and g22383 ( n21006 , n23821 , n17769 );
    xnor g22384 ( n13208 , n17212 , n26725 );
    xnor g22385 ( n12555 , n11209 , n23250 );
    not g22386 ( n14507 , n14603 );
    not g22387 ( n3090 , n7822 );
    not g22388 ( n26235 , n5285 );
    xnor g22389 ( n25963 , n21021 , n18355 );
    nor g22390 ( n707 , n2776 , n4853 );
    xnor g22391 ( n10000 , n19957 , n26954 );
    not g22392 ( n16672 , n22105 );
    not g22393 ( n27122 , n4913 );
    nor g22394 ( n24304 , n9988 , n17824 );
    and g22395 ( n24567 , n27119 , n10656 );
    or g22396 ( n21855 , n840 , n21001 );
    xnor g22397 ( n10289 , n19682 , n9133 );
    or g22398 ( n5423 , n20852 , n26283 );
    xnor g22399 ( n17114 , n24802 , n19108 );
    not g22400 ( n978 , n21964 );
    xnor g22401 ( n15910 , n11527 , n24365 );
    not g22402 ( n22232 , n14045 );
    and g22403 ( n23375 , n1511 , n19690 );
    xnor g22404 ( n8109 , n5979 , n18455 );
    or g22405 ( n15341 , n2576 , n21276 );
    or g22406 ( n9078 , n11650 , n20901 );
    not g22407 ( n13088 , n21915 );
    xnor g22408 ( n25312 , n599 , n22888 );
    xnor g22409 ( n7138 , n10454 , n21856 );
    or g22410 ( n16996 , n1458 , n22433 );
    xnor g22411 ( n2323 , n7601 , n4656 );
    not g22412 ( n6865 , n6613 );
    nor g22413 ( n1067 , n1843 , n25667 );
    xnor g22414 ( n22899 , n16882 , n16683 );
    and g22415 ( n5171 , n25819 , n1050 );
    not g22416 ( n1132 , n5200 );
    not g22417 ( n11045 , n2160 );
    or g22418 ( n26029 , n23923 , n23874 );
    or g22419 ( n23025 , n22519 , n10734 );
    or g22420 ( n26759 , n8605 , n8668 );
    nor g22421 ( n9526 , n19108 , n24802 );
    not g22422 ( n13234 , n6109 );
    not g22423 ( n10048 , n224 );
    or g22424 ( n18239 , n5238 , n26193 );
    xnor g22425 ( n21014 , n9746 , n22391 );
    not g22426 ( n10998 , n15016 );
    nor g22427 ( n9231 , n5420 , n14554 );
    xnor g22428 ( n17285 , n6343 , n25798 );
    or g22429 ( n24003 , n16812 , n1279 );
    not g22430 ( n19055 , n14918 );
    not g22431 ( n3940 , n13455 );
    or g22432 ( n4379 , n21563 , n8365 );
    and g22433 ( n10765 , n13550 , n12062 );
    not g22434 ( n7360 , n1654 );
    or g22435 ( n25294 , n15763 , n5662 );
    xnor g22436 ( n10383 , n26991 , n1354 );
    nor g22437 ( n1424 , n7057 , n7823 );
    xnor g22438 ( n3244 , n20309 , n14194 );
    or g22439 ( n20283 , n21536 , n16491 );
    or g22440 ( n21843 , n19201 , n23211 );
    not g22441 ( n5342 , n24451 );
    xnor g22442 ( n12938 , n5072 , n1132 );
    not g22443 ( n17505 , n22020 );
    and g22444 ( n13165 , n19770 , n11451 );
    or g22445 ( n24888 , n15542 , n8221 );
    and g22446 ( n15781 , n26781 , n20738 );
    xnor g22447 ( n25624 , n14182 , n2113 );
    xnor g22448 ( n25679 , n14984 , n17954 );
    and g22449 ( n22706 , n6393 , n19082 );
    or g22450 ( n22696 , n26104 , n10527 );
    xnor g22451 ( n4959 , n1190 , n20353 );
    and g22452 ( n25129 , n8773 , n11657 );
    xnor g22453 ( n24504 , n6834 , n8399 );
    and g22454 ( n9669 , n23095 , n21704 );
    xnor g22455 ( n20391 , n21311 , n6216 );
    or g22456 ( n21167 , n20570 , n1934 );
    nor g22457 ( n3807 , n8875 , n19215 );
    or g22458 ( n6187 , n24849 , n26785 );
    nor g22459 ( n21377 , n18710 , n21796 );
    or g22460 ( n12634 , n1624 , n23829 );
    xnor g22461 ( n12824 , n18338 , n17549 );
    or g22462 ( n11561 , n18257 , n19905 );
    nor g22463 ( n8878 , n8614 , n24705 );
    nor g22464 ( n20037 , n24550 , n25405 );
    or g22465 ( n3757 , n14988 , n8201 );
    xnor g22466 ( n15999 , n18735 , n14393 );
    nor g22467 ( n3661 , n11486 , n18409 );
    xnor g22468 ( n20850 , n5296 , n8672 );
    or g22469 ( n4378 , n2314 , n1163 );
    nor g22470 ( n25279 , n8152 , n19695 );
    xnor g22471 ( n25423 , n26264 , n19454 );
    nor g22472 ( n17899 , n6168 , n12151 );
    not g22473 ( n16665 , n18584 );
    and g22474 ( n19068 , n18150 , n21440 );
    or g22475 ( n18338 , n20202 , n24633 );
    and g22476 ( n7214 , n1031 , n8443 );
    xnor g22477 ( n387 , n3201 , n9085 );
    and g22478 ( n2047 , n11861 , n22641 );
    nor g22479 ( n6982 , n978 , n26946 );
    xnor g22480 ( n6457 , n14453 , n16860 );
    or g22481 ( n18093 , n20612 , n21264 );
    not g22482 ( n4752 , n19033 );
    or g22483 ( n20994 , n26717 , n26748 );
    not g22484 ( n15930 , n7684 );
    not g22485 ( n1396 , n4024 );
    or g22486 ( n10877 , n16711 , n2059 );
    xnor g22487 ( n17560 , n2289 , n18345 );
    or g22488 ( n12656 , n18090 , n12474 );
    and g22489 ( n21108 , n21643 , n101 );
    or g22490 ( n8903 , n8106 , n10904 );
    xnor g22491 ( n10346 , n18480 , n9499 );
    or g22492 ( n11700 , n25246 , n24728 );
    xnor g22493 ( n17798 , n16443 , n23996 );
    or g22494 ( n9776 , n605 , n8691 );
    xnor g22495 ( n25501 , n20249 , n24684 );
    xnor g22496 ( n4263 , n26720 , n11832 );
    and g22497 ( n3181 , n2465 , n13101 );
    or g22498 ( n6324 , n20140 , n4308 );
    xnor g22499 ( n22213 , n4209 , n21212 );
    or g22500 ( n21273 , n6341 , n21246 );
    or g22501 ( n10786 , n19541 , n23863 );
    nor g22502 ( n958 , n8420 , n10406 );
    xnor g22503 ( n16310 , n23983 , n20040 );
    and g22504 ( n19122 , n15579 , n293 );
    nor g22505 ( n10992 , n2915 , n12014 );
    and g22506 ( n6562 , n7469 , n12608 );
    and g22507 ( n15270 , n11951 , n18713 );
    xnor g22508 ( n26803 , n6696 , n23423 );
    not g22509 ( n23005 , n23102 );
    xnor g22510 ( n23752 , n11150 , n4063 );
    not g22511 ( n1401 , n14830 );
    not g22512 ( n20323 , n23102 );
    xnor g22513 ( n6851 , n5551 , n22078 );
    not g22514 ( n22729 , n10018 );
    xnor g22515 ( n9047 , n21714 , n14868 );
    xnor g22516 ( n6686 , n23141 , n20792 );
    and g22517 ( n8877 , n11388 , n17161 );
    nor g22518 ( n23431 , n10106 , n17379 );
    or g22519 ( n24566 , n2719 , n15229 );
    xnor g22520 ( n19450 , n8686 , n25585 );
    or g22521 ( n16914 , n23563 , n2434 );
    not g22522 ( n456 , n6523 );
    xnor g22523 ( n19152 , n19494 , n2387 );
    not g22524 ( n12311 , n2167 );
    or g22525 ( n230 , n5065 , n8487 );
    and g22526 ( n27129 , n23023 , n23520 );
    not g22527 ( n17932 , n19820 );
    xnor g22528 ( n26449 , n10885 , n19276 );
    and g22529 ( n24523 , n19531 , n11425 );
    nor g22530 ( n20424 , n2969 , n3066 );
    or g22531 ( n4793 , n19331 , n11675 );
    xnor g22532 ( n15955 , n2899 , n6485 );
    not g22533 ( n7604 , n1469 );
    and g22534 ( n3609 , n10670 , n19232 );
    or g22535 ( n12020 , n10914 , n17685 );
    or g22536 ( n8341 , n23492 , n22307 );
    xnor g22537 ( n14352 , n24129 , n9380 );
    xnor g22538 ( n4631 , n7532 , n17664 );
    and g22539 ( n20845 , n13057 , n12391 );
    or g22540 ( n19319 , n26420 , n21694 );
    and g22541 ( n19980 , n19077 , n23149 );
    nor g22542 ( n14953 , n22962 , n1715 );
    or g22543 ( n21892 , n11178 , n1079 );
    or g22544 ( n607 , n10948 , n10243 );
    or g22545 ( n13264 , n20986 , n12212 );
    and g22546 ( n22415 , n15184 , n16605 );
    and g22547 ( n25117 , n13389 , n17695 );
    or g22548 ( n11873 , n11456 , n25118 );
    buf g22549 ( n8891 , n22079 );
    or g22550 ( n14846 , n20716 , n6708 );
    or g22551 ( n8316 , n21222 , n18820 );
    or g22552 ( n15849 , n16047 , n14167 );
    nor g22553 ( n18134 , n3324 , n2272 );
    and g22554 ( n23533 , n9235 , n24667 );
    xnor g22555 ( n17889 , n19744 , n24955 );
    nor g22556 ( n14363 , n4293 , n5739 );
    not g22557 ( n10832 , n115 );
    xnor g22558 ( n22272 , n6775 , n3925 );
    xnor g22559 ( n17485 , n10842 , n18571 );
    and g22560 ( n26243 , n6966 , n27128 );
    nor g22561 ( n9138 , n692 , n26015 );
    xnor g22562 ( n12832 , n8539 , n15975 );
    or g22563 ( n14448 , n26264 , n5661 );
    or g22564 ( n16784 , n7726 , n3550 );
    and g22565 ( n5873 , n10325 , n8544 );
    or g22566 ( n6980 , n2330 , n9188 );
    not g22567 ( n24091 , n26927 );
    xnor g22568 ( n1860 , n2921 , n362 );
    not g22569 ( n6648 , n14649 );
    and g22570 ( n15904 , n16867 , n9173 );
    xnor g22571 ( n16874 , n11747 , n23400 );
    xnor g22572 ( n22592 , n20179 , n26823 );
    and g22573 ( n8260 , n21646 , n22098 );
    xnor g22574 ( n14096 , n20153 , n13308 );
    and g22575 ( n9758 , n24950 , n13416 );
    and g22576 ( n8768 , n7016 , n12584 );
    xnor g22577 ( n24473 , n13433 , n16915 );
    or g22578 ( n22347 , n53 , n14487 );
    not g22579 ( n9096 , n21016 );
    or g22580 ( n9139 , n21341 , n23780 );
    and g22581 ( n3820 , n23516 , n17258 );
    xnor g22582 ( n23006 , n25906 , n22832 );
    xnor g22583 ( n5073 , n23509 , n23755 );
    nor g22584 ( n3345 , n14826 , n13549 );
    xnor g22585 ( n3878 , n25862 , n9996 );
    or g22586 ( n6146 , n5238 , n7351 );
    and g22587 ( n24545 , n24383 , n6403 );
    xnor g22588 ( n14063 , n5320 , n24330 );
    or g22589 ( n18411 , n15358 , n6182 );
    not g22590 ( n23097 , n24475 );
    nor g22591 ( n18000 , n20040 , n9396 );
    and g22592 ( n5413 , n14859 , n3039 );
    xnor g22593 ( n1074 , n10086 , n25330 );
    xnor g22594 ( n11607 , n5558 , n7791 );
    xnor g22595 ( n9975 , n5065 , n6204 );
    xnor g22596 ( n13425 , n4677 , n3918 );
    and g22597 ( n25823 , n1705 , n9456 );
    or g22598 ( n13260 , n18159 , n8887 );
    not g22599 ( n14705 , n10407 );
    xnor g22600 ( n4476 , n21440 , n17833 );
    and g22601 ( n22029 , n13367 , n20970 );
    nor g22602 ( n7836 , n23784 , n4127 );
    or g22603 ( n25640 , n10452 , n22723 );
    or g22604 ( n25661 , n16711 , n21753 );
    and g22605 ( n3103 , n3129 , n26365 );
    nor g22606 ( n25740 , n20751 , n24593 );
    not g22607 ( n1365 , n18962 );
    xnor g22608 ( n15327 , n12340 , n16659 );
    or g22609 ( n14023 , n25742 , n7312 );
    xnor g22610 ( n13860 , n24161 , n4426 );
    or g22611 ( n22616 , n19466 , n25594 );
    or g22612 ( n7301 , n21918 , n18974 );
    or g22613 ( n18095 , n14119 , n7963 );
    xnor g22614 ( n7008 , n9395 , n7144 );
    xnor g22615 ( n5776 , n3624 , n10905 );
    and g22616 ( n6415 , n24073 , n12170 );
    xnor g22617 ( n22734 , n19033 , n7674 );
    or g22618 ( n4761 , n5226 , n11223 );
    xnor g22619 ( n24412 , n19143 , n5891 );
    and g22620 ( n12633 , n18117 , n6997 );
    buf g22621 ( n11322 , n24451 );
    and g22622 ( n19268 , n21924 , n9476 );
    xnor g22623 ( n10138 , n26185 , n4573 );
    and g22624 ( n4988 , n2795 , n12796 );
    nor g22625 ( n2115 , n2576 , n1682 );
    and g22626 ( n14396 , n927 , n17165 );
    nor g22627 ( n23054 , n9631 , n22879 );
    not g22628 ( n20554 , n9445 );
    not g22629 ( n3393 , n22972 );
    xnor g22630 ( n25665 , n5669 , n4358 );
    or g22631 ( n19430 , n2850 , n14482 );
    xnor g22632 ( n24482 , n5934 , n23636 );
    and g22633 ( n15479 , n10636 , n16362 );
    xnor g22634 ( n824 , n23559 , n21455 );
    or g22635 ( n10729 , n10738 , n6934 );
    nor g22636 ( n9407 , n23586 , n17728 );
    and g22637 ( n10926 , n17435 , n2905 );
    or g22638 ( n16317 , n2637 , n4248 );
    xnor g22639 ( n5503 , n25967 , n24327 );
    and g22640 ( n5640 , n17579 , n12452 );
    xnor g22641 ( n14419 , n9605 , n11806 );
    not g22642 ( n20273 , n6414 );
    and g22643 ( n12042 , n21956 , n16076 );
    nor g22644 ( n9000 , n22859 , n12859 );
    not g22645 ( n25931 , n24150 );
    or g22646 ( n17345 , n10480 , n23840 );
    not g22647 ( n7868 , n17614 );
    or g22648 ( n26493 , n6422 , n13503 );
    xnor g22649 ( n8461 , n22631 , n21078 );
    xnor g22650 ( n18753 , n17978 , n6456 );
    or g22651 ( n5303 , n5255 , n6446 );
    not g22652 ( n3258 , n3793 );
    nor g22653 ( n22323 , n13152 , n2688 );
    nor g22654 ( n1768 , n15602 , n8507 );
    and g22655 ( n6072 , n25420 , n14807 );
    or g22656 ( n20889 , n17449 , n568 );
    xnor g22657 ( n24326 , n16111 , n20109 );
    or g22658 ( n26424 , n16029 , n4322 );
    not g22659 ( n8873 , n18589 );
    nor g22660 ( n21790 , n17626 , n2246 );
    xnor g22661 ( n19727 , n17098 , n11096 );
    or g22662 ( n89 , n5427 , n19633 );
    or g22663 ( n4962 , n11740 , n11816 );
    or g22664 ( n5504 , n23718 , n17221 );
    or g22665 ( n1056 , n12575 , n19325 );
    or g22666 ( n17031 , n13529 , n20594 );
    not g22667 ( n17184 , n21510 );
    or g22668 ( n26858 , n18123 , n1697 );
    not g22669 ( n15422 , n17771 );
    nor g22670 ( n24341 , n18787 , n5944 );
    or g22671 ( n533 , n3721 , n26403 );
    xnor g22672 ( n17903 , n5682 , n10468 );
    xnor g22673 ( n21918 , n12559 , n6620 );
    nor g22674 ( n10050 , n20045 , n19357 );
    xnor g22675 ( n15087 , n17363 , n4758 );
    or g22676 ( n17603 , n16496 , n17647 );
    or g22677 ( n25315 , n15136 , n13051 );
    or g22678 ( n2179 , n16128 , n1002 );
    and g22679 ( n15587 , n116 , n16069 );
    and g22680 ( n6494 , n6259 , n14838 );
    or g22681 ( n5202 , n27140 , n19028 );
    not g22682 ( n13 , n26038 );
    xnor g22683 ( n25940 , n1487 , n22928 );
    not g22684 ( n1340 , n20409 );
    and g22685 ( n13927 , n16983 , n14411 );
    xnor g22686 ( n5695 , n9711 , n11317 );
    or g22687 ( n8464 , n20342 , n26830 );
    xnor g22688 ( n16562 , n5985 , n22514 );
    or g22689 ( n13101 , n19688 , n7024 );
    or g22690 ( n9520 , n14306 , n14400 );
    nor g22691 ( n9913 , n395 , n19215 );
    xnor g22692 ( n9695 , n20943 , n17526 );
    xnor g22693 ( n20197 , n3257 , n3677 );
    or g22694 ( n9625 , n10651 , n23639 );
    not g22695 ( n24939 , n26565 );
    or g22696 ( n26863 , n7997 , n15851 );
    xnor g22697 ( n12908 , n7241 , n10592 );
    or g22698 ( n18447 , n483 , n8827 );
    not g22699 ( n14477 , n19138 );
    nor g22700 ( n14897 , n14878 , n16213 );
    nor g22701 ( n4819 , n12956 , n1118 );
    xnor g22702 ( n18763 , n22219 , n4781 );
    xnor g22703 ( n464 , n17734 , n16900 );
    or g22704 ( n9312 , n15505 , n5264 );
    and g22705 ( n7409 , n17179 , n6035 );
    or g22706 ( n16160 , n15127 , n26680 );
    not g22707 ( n4093 , n4105 );
    not g22708 ( n2342 , n3468 );
    xnor g22709 ( n22300 , n11824 , n5709 );
    not g22710 ( n21037 , n26523 );
    and g22711 ( n18976 , n13023 , n9548 );
    or g22712 ( n17822 , n21268 , n14899 );
    xnor g22713 ( n23709 , n18111 , n2944 );
    and g22714 ( n4755 , n24893 , n174 );
    xnor g22715 ( n9483 , n25345 , n23463 );
    xnor g22716 ( n16136 , n15099 , n8825 );
    xnor g22717 ( n12420 , n11397 , n12043 );
    or g22718 ( n2034 , n21767 , n23985 );
    and g22719 ( n22749 , n11611 , n13186 );
    xnor g22720 ( n12201 , n26947 , n4467 );
    nor g22721 ( n5426 , n8000 , n13035 );
    xnor g22722 ( n8001 , n2186 , n19148 );
    nor g22723 ( n7080 , n25512 , n23132 );
    not g22724 ( n17789 , n16430 );
    or g22725 ( n702 , n16820 , n18944 );
    xnor g22726 ( n22150 , n187 , n10549 );
    or g22727 ( n3145 , n24735 , n26339 );
    not g22728 ( n13875 , n16214 );
    or g22729 ( n18379 , n22198 , n24493 );
    and g22730 ( n1326 , n331 , n684 );
    xor g22731 ( n7905 , n25913 , n5490 );
    or g22732 ( n5595 , n6288 , n14333 );
    xnor g22733 ( n142 , n20911 , n11576 );
    not g22734 ( n3276 , n3164 );
    and g22735 ( n26010 , n8175 , n13423 );
    not g22736 ( n4490 , n20169 );
    xnor g22737 ( n7277 , n10462 , n25630 );
    xnor g22738 ( n14977 , n14655 , n13258 );
    xnor g22739 ( n3245 , n4557 , n3573 );
    not g22740 ( n8597 , n24093 );
    or g22741 ( n14460 , n18293 , n11444 );
    not g22742 ( n405 , n26553 );
    and g22743 ( n10517 , n1964 , n21387 );
    or g22744 ( n17284 , n26997 , n6185 );
    xnor g22745 ( n18434 , n20679 , n15624 );
    and g22746 ( n13656 , n22645 , n12711 );
    nor g22747 ( n22434 , n26445 , n3881 );
    and g22748 ( n10941 , n8363 , n2812 );
    nor g22749 ( n5013 , n2659 , n9957 );
    not g22750 ( n17418 , n4670 );
    buf g22751 ( n25514 , n11414 );
    not g22752 ( n25194 , n2073 );
    not g22753 ( n4004 , n25905 );
    and g22754 ( n13702 , n2702 , n22863 );
    and g22755 ( n10329 , n5076 , n22438 );
    and g22756 ( n15531 , n23335 , n12678 );
    not g22757 ( n19952 , n3541 );
    not g22758 ( n4330 , n27022 );
    xnor g22759 ( n22610 , n22629 , n23735 );
    not g22760 ( n9387 , n20822 );
    buf g22761 ( n25846 , n24932 );
    xnor g22762 ( n18596 , n8612 , n3324 );
    nor g22763 ( n12819 , n10343 , n8997 );
    not g22764 ( n2588 , n2425 );
    and g22765 ( n6295 , n17182 , n21625 );
    or g22766 ( n10107 , n15077 , n23412 );
    and g22767 ( n20541 , n4893 , n21451 );
    not g22768 ( n5222 , n19069 );
    not g22769 ( n12878 , n11733 );
    and g22770 ( n14348 , n14205 , n19998 );
    or g22771 ( n6188 , n11055 , n9162 );
    not g22772 ( n23769 , n8845 );
    not g22773 ( n26963 , n379 );
    and g22774 ( n13593 , n13900 , n19744 );
    xnor g22775 ( n18680 , n3968 , n16900 );
    not g22776 ( n23804 , n15506 );
    nor g22777 ( n16135 , n5172 , n16948 );
    and g22778 ( n14199 , n7386 , n13242 );
    xnor g22779 ( n4674 , n26346 , n12194 );
    xnor g22780 ( n6154 , n17709 , n23747 );
    or g22781 ( n25248 , n5498 , n16294 );
    xnor g22782 ( n6554 , n24067 , n20221 );
    not g22783 ( n8451 , n6168 );
    or g22784 ( n20773 , n14899 , n18496 );
    xnor g22785 ( n27105 , n8363 , n2145 );
    or g22786 ( n14616 , n10488 , n2649 );
    xnor g22787 ( n20406 , n21283 , n20859 );
    and g22788 ( n7013 , n18649 , n13968 );
    or g22789 ( n5718 , n15950 , n4399 );
    or g22790 ( n11099 , n6307 , n13079 );
    xnor g22791 ( n11159 , n10358 , n8484 );
    xnor g22792 ( n11845 , n18715 , n9247 );
    and g22793 ( n23651 , n21090 , n1241 );
    or g22794 ( n11839 , n19733 , n21338 );
    and g22795 ( n18701 , n18095 , n18697 );
    xnor g22796 ( n13487 , n24120 , n24446 );
    xnor g22797 ( n24191 , n4887 , n15861 );
    or g22798 ( n3930 , n1967 , n17334 );
    nor g22799 ( n296 , n2857 , n13282 );
    or g22800 ( n21330 , n10704 , n11908 );
    xnor g22801 ( n4585 , n4800 , n25846 );
    not g22802 ( n9594 , n9323 );
    xnor g22803 ( n22940 , n3479 , n22386 );
    xnor g22804 ( n1109 , n5302 , n19116 );
    xnor g22805 ( n25925 , n20444 , n19313 );
    or g22806 ( n5571 , n11027 , n7904 );
    or g22807 ( n13364 , n24324 , n9437 );
    xnor g22808 ( n17215 , n6043 , n13039 );
    not g22809 ( n2509 , n22654 );
    xnor g22810 ( n2900 , n21372 , n13276 );
    or g22811 ( n20520 , n3931 , n20076 );
    not g22812 ( n5668 , n10554 );
    and g22813 ( n16303 , n8394 , n10801 );
    xnor g22814 ( n1723 , n6239 , n20209 );
    xnor g22815 ( n25261 , n2956 , n8985 );
    or g22816 ( n2353 , n19596 , n15191 );
    or g22817 ( n595 , n20605 , n1756 );
    or g22818 ( n1801 , n26793 , n26470 );
    xnor g22819 ( n17749 , n10991 , n6463 );
    nor g22820 ( n1198 , n400 , n2322 );
    or g22821 ( n5311 , n25402 , n21084 );
    or g22822 ( n2796 , n22909 , n19524 );
    xnor g22823 ( n6991 , n19514 , n2731 );
    or g22824 ( n21136 , n7071 , n22122 );
    not g22825 ( n8690 , n2420 );
    xnor g22826 ( n2861 , n5140 , n10250 );
    or g22827 ( n15418 , n4469 , n7212 );
    xnor g22828 ( n11752 , n10041 , n10514 );
    not g22829 ( n1346 , n24638 );
    and g22830 ( n22447 , n7319 , n17224 );
    nor g22831 ( n475 , n8451 , n17047 );
    and g22832 ( n14237 , n22825 , n22689 );
    or g22833 ( n9478 , n3092 , n18645 );
    xnor g22834 ( n3187 , n24129 , n26167 );
    nor g22835 ( n7705 , n18514 , n16507 );
    and g22836 ( n12017 , n18456 , n23530 );
    xnor g22837 ( n9075 , n16058 , n4846 );
    and g22838 ( n3951 , n828 , n25757 );
    xor g22839 ( n22530 , n13918 , n11672 );
    not g22840 ( n12360 , n15800 );
    xnor g22841 ( n26647 , n25624 , n19327 );
    or g22842 ( n7715 , n21263 , n7376 );
    or g22843 ( n11203 , n1734 , n5218 );
    or g22844 ( n8833 , n7419 , n1126 );
    and g22845 ( n16148 , n26436 , n15459 );
    or g22846 ( n7782 , n7111 , n15546 );
    not g22847 ( n15239 , n27042 );
    or g22848 ( n20414 , n6769 , n3852 );
    xnor g22849 ( n21405 , n10642 , n23142 );
    or g22850 ( n6292 , n11000 , n18037 );
    xnor g22851 ( n18350 , n20995 , n12680 );
    not g22852 ( n7133 , n19491 );
    and g22853 ( n20141 , n9574 , n1980 );
    nor g22854 ( n5040 , n11355 , n12596 );
    xnor g22855 ( n5300 , n2806 , n4688 );
    or g22856 ( n19279 , n25923 , n24184 );
    or g22857 ( n11264 , n23431 , n25449 );
    buf g22858 ( n682 , n7636 );
    or g22859 ( n24775 , n8228 , n5570 );
    and g22860 ( n3240 , n8758 , n7591 );
    xnor g22861 ( n20791 , n5101 , n6659 );
    xnor g22862 ( n13070 , n8398 , n17711 );
    not g22863 ( n20639 , n5874 );
    nor g22864 ( n17628 , n617 , n20982 );
    xnor g22865 ( n4228 , n20354 , n18097 );
    xnor g22866 ( n12195 , n4499 , n21671 );
    or g22867 ( n17393 , n15241 , n15146 );
    and g22868 ( n67 , n1968 , n20223 );
    xnor g22869 ( n8584 , n25302 , n3440 );
    and g22870 ( n4162 , n3773 , n6294 );
    not g22871 ( n21269 , n24897 );
    xnor g22872 ( n16104 , n22413 , n18265 );
    or g22873 ( n25642 , n10804 , n20901 );
    or g22874 ( n26657 , n9985 , n14142 );
    xnor g22875 ( n25547 , n13006 , n6933 );
    or g22876 ( n96 , n15727 , n16685 );
    or g22877 ( n26210 , n26565 , n9142 );
    and g22878 ( n1980 , n15700 , n5828 );
    and g22879 ( n9506 , n10802 , n1719 );
    or g22880 ( n16153 , n22808 , n7824 );
    not g22881 ( n17539 , n987 );
    nor g22882 ( n19706 , n3254 , n2738 );
    xnor g22883 ( n4576 , n21640 , n3492 );
    not g22884 ( n5557 , n21622 );
    xnor g22885 ( n13710 , n6512 , n1723 );
    or g22886 ( n23150 , n5505 , n27018 );
    not g22887 ( n11676 , n16707 );
    or g22888 ( n19963 , n25038 , n1380 );
    or g22889 ( n11042 , n2476 , n25414 );
    or g22890 ( n17740 , n25914 , n9242 );
    xnor g22891 ( n16373 , n1641 , n5093 );
    nor g22892 ( n20780 , n2230 , n7973 );
    xnor g22893 ( n3861 , n443 , n18903 );
    nor g22894 ( n14260 , n18662 , n12657 );
    xnor g22895 ( n3823 , n9279 , n5769 );
    and g22896 ( n6181 , n17610 , n11327 );
    and g22897 ( n1751 , n19061 , n13436 );
    and g22898 ( n21002 , n7659 , n15563 );
    xnor g22899 ( n21050 , n5382 , n16226 );
    not g22900 ( n16627 , n11653 );
    and g22901 ( n1928 , n21277 , n1908 );
    or g22902 ( n21166 , n18569 , n14635 );
    or g22903 ( n12340 , n13807 , n301 );
    xnor g22904 ( n15698 , n5136 , n23388 );
    xnor g22905 ( n24887 , n7786 , n14446 );
    xnor g22906 ( n3814 , n12381 , n10557 );
    and g22907 ( n25562 , n14250 , n25714 );
    and g22908 ( n12182 , n26260 , n4214 );
    or g22909 ( n22280 , n17851 , n2691 );
    xnor g22910 ( n18283 , n19167 , n26228 );
    and g22911 ( n22011 , n22929 , n21844 );
    and g22912 ( n9471 , n25629 , n2291 );
    not g22913 ( n1730 , n6373 );
    nor g22914 ( n3130 , n19222 , n1786 );
    or g22915 ( n18939 , n3551 , n17259 );
    xnor g22916 ( n21275 , n23013 , n21622 );
    not g22917 ( n1704 , n26860 );
    xnor g22918 ( n13438 , n17251 , n26107 );
    not g22919 ( n9100 , n5661 );
    xnor g22920 ( n2059 , n16810 , n11739 );
    or g22921 ( n1171 , n4918 , n5235 );
    and g22922 ( n15083 , n23913 , n24325 );
    or g22923 ( n8667 , n16213 , n6468 );
    and g22924 ( n17050 , n20813 , n8290 );
    and g22925 ( n18881 , n12656 , n26869 );
    xnor g22926 ( n24499 , n11871 , n18809 );
    xnor g22927 ( n27127 , n17728 , n22652 );
    not g22928 ( n16094 , n3232 );
    or g22929 ( n2953 , n16122 , n6522 );
    or g22930 ( n10649 , n15695 , n11088 );
    and g22931 ( n11188 , n15265 , n9911 );
    and g22932 ( n5047 , n22003 , n7414 );
    or g22933 ( n14115 , n11346 , n8902 );
    or g22934 ( n12879 , n24125 , n15719 );
    or g22935 ( n21971 , n6456 , n8881 );
    xnor g22936 ( n23766 , n9453 , n3959 );
    not g22937 ( n26093 , n10372 );
    and g22938 ( n8957 , n4992 , n26736 );
    nor g22939 ( n12609 , n4325 , n21941 );
    nor g22940 ( n25432 , n25915 , n13745 );
    and g22941 ( n21028 , n21518 , n16338 );
    and g22942 ( n8613 , n627 , n10579 );
    xnor g22943 ( n14471 , n15197 , n911 );
    and g22944 ( n2749 , n24615 , n6181 );
    not g22945 ( n20516 , n13115 );
    or g22946 ( n26412 , n5646 , n16079 );
    or g22947 ( n14235 , n21423 , n19781 );
    or g22948 ( n4013 , n25347 , n20627 );
    and g22949 ( n22459 , n22597 , n16473 );
    nor g22950 ( n20334 , n656 , n3143 );
    or g22951 ( n10042 , n14821 , n7714 );
    nor g22952 ( n5106 , n1215 , n10486 );
    or g22953 ( n19601 , n18518 , n8733 );
    xnor g22954 ( n1186 , n12778 , n10577 );
    xnor g22955 ( n12383 , n9714 , n8112 );
    or g22956 ( n2652 , n26120 , n4116 );
    not g22957 ( n12797 , n3903 );
    or g22958 ( n20943 , n4223 , n4364 );
    xnor g22959 ( n12043 , n17911 , n25331 );
    xnor g22960 ( n4120 , n21316 , n25073 );
    not g22961 ( n11516 , n14387 );
    not g22962 ( n16111 , n19652 );
    or g22963 ( n21103 , n3011 , n220 );
    and g22964 ( n17666 , n12604 , n20766 );
    xnor g22965 ( n335 , n24612 , n21471 );
    or g22966 ( n2153 , n11901 , n2281 );
    or g22967 ( n19960 , n12764 , n26846 );
    nor g22968 ( n8288 , n8836 , n22853 );
    or g22969 ( n1813 , n13796 , n24740 );
    xnor g22970 ( n18481 , n8745 , n16476 );
    and g22971 ( n15911 , n18269 , n10784 );
    xnor g22972 ( n592 , n22663 , n10737 );
    or g22973 ( n4229 , n26421 , n25359 );
    xnor g22974 ( n3040 , n25229 , n25079 );
    not g22975 ( n15415 , n26318 );
    or g22976 ( n2973 , n7198 , n25914 );
    xnor g22977 ( n24076 , n26085 , n23974 );
    xnor g22978 ( n21228 , n333 , n13625 );
    xnor g22979 ( n1457 , n23160 , n2421 );
    nor g22980 ( n15989 , n23141 , n5579 );
    or g22981 ( n8610 , n15261 , n14630 );
    xnor g22982 ( n5727 , n14029 , n19203 );
    nor g22983 ( n18646 , n15404 , n10610 );
    xnor g22984 ( n22960 , n16785 , n9702 );
    xnor g22985 ( n22364 , n461 , n8678 );
    xnor g22986 ( n12806 , n8414 , n17679 );
    xnor g22987 ( n15872 , n18 , n26808 );
    or g22988 ( n8664 , n11694 , n18040 );
    or g22989 ( n9306 , n22877 , n6582 );
    nor g22990 ( n15943 , n6935 , n13249 );
    xnor g22991 ( n4782 , n15365 , n26545 );
    and g22992 ( n13200 , n7459 , n19253 );
    or g22993 ( n19135 , n17448 , n25167 );
    xnor g22994 ( n17984 , n8363 , n11481 );
    and g22995 ( n9674 , n6091 , n11813 );
    not g22996 ( n24355 , n12507 );
    xnor g22997 ( n21367 , n21099 , n17704 );
    or g22998 ( n18023 , n4697 , n9311 );
    xnor g22999 ( n20027 , n10406 , n6456 );
    or g23000 ( n13320 , n12543 , n25435 );
    not g23001 ( n23962 , n1717 );
    or g23002 ( n4117 , n24609 , n8044 );
    nor g23003 ( n7590 , n11039 , n12679 );
    not g23004 ( n23489 , n22198 );
    or g23005 ( n16580 , n7198 , n8571 );
    xnor g23006 ( n8760 , n23686 , n7523 );
    and g23007 ( n26422 , n8092 , n25278 );
    and g23008 ( n16184 , n19599 , n24055 );
    not g23009 ( n23996 , n13166 );
    xnor g23010 ( n20417 , n19145 , n14050 );
    not g23011 ( n24804 , n25100 );
    nor g23012 ( n11702 , n10637 , n4226 );
    or g23013 ( n12007 , n25953 , n4429 );
    or g23014 ( n10569 , n20732 , n23236 );
    xnor g23015 ( n1764 , n3078 , n26161 );
    nor g23016 ( n6136 , n3623 , n22517 );
    and g23017 ( n24762 , n9172 , n10571 );
    or g23018 ( n15656 , n19692 , n4840 );
    or g23019 ( n25757 , n12459 , n19324 );
    xnor g23020 ( n15336 , n4304 , n23876 );
    not g23021 ( n2171 , n9509 );
    or g23022 ( n21959 , n12004 , n12289 );
    nor g23023 ( n3185 , n17276 , n3780 );
    not g23024 ( n27068 , n12153 );
    or g23025 ( n10391 , n25336 , n20433 );
    and g23026 ( n21290 , n8351 , n11066 );
    and g23027 ( n13099 , n1587 , n14008 );
    and g23028 ( n18135 , n8627 , n9543 );
    and g23029 ( n10956 , n5617 , n22414 );
    and g23030 ( n15403 , n2684 , n3680 );
    or g23031 ( n25965 , n10771 , n7033 );
    or g23032 ( n4200 , n8678 , n16500 );
    not g23033 ( n1686 , n3825 );
    xnor g23034 ( n23374 , n13529 , n7056 );
    xnor g23035 ( n24268 , n8570 , n14728 );
    and g23036 ( n13778 , n20156 , n26440 );
    and g23037 ( n4006 , n8839 , n22758 );
    or g23038 ( n5894 , n22802 , n27087 );
    nor g23039 ( n8180 , n456 , n15400 );
    xnor g23040 ( n8619 , n17630 , n18263 );
    not g23041 ( n21268 , n7026 );
    xnor g23042 ( n6296 , n17122 , n14389 );
    and g23043 ( n25480 , n14254 , n6964 );
    and g23044 ( n1963 , n9004 , n21014 );
    and g23045 ( n19953 , n9804 , n8663 );
    not g23046 ( n19429 , n10477 );
    xnor g23047 ( n7354 , n19331 , n24187 );
    not g23048 ( n16913 , n2517 );
    or g23049 ( n11934 , n20871 , n9612 );
    not g23050 ( n20009 , n14437 );
    xnor g23051 ( n1943 , n14713 , n10311 );
    not g23052 ( n11901 , n6814 );
    not g23053 ( n14852 , n24340 );
    nor g23054 ( n15748 , n13044 , n8845 );
    xnor g23055 ( n16058 , n16231 , n17754 );
    nor g23056 ( n1191 , n2570 , n7569 );
    xnor g23057 ( n7702 , n932 , n10739 );
    xnor g23058 ( n19772 , n27111 , n25265 );
    and g23059 ( n6083 , n10491 , n22103 );
    nor g23060 ( n7389 , n18558 , n6556 );
    xnor g23061 ( n10511 , n20442 , n16988 );
    or g23062 ( n6629 , n18413 , n15591 );
    or g23063 ( n23846 , n13239 , n22356 );
    and g23064 ( n7799 , n212 , n17150 );
    and g23065 ( n12946 , n8012 , n20870 );
    or g23066 ( n23368 , n9756 , n24820 );
    or g23067 ( n7956 , n13023 , n6631 );
    not g23068 ( n6173 , n12113 );
    nor g23069 ( n5455 , n339 , n11266 );
    and g23070 ( n19452 , n25370 , n11603 );
    or g23071 ( n3839 , n5763 , n23548 );
    or g23072 ( n12856 , n2268 , n22417 );
    not g23073 ( n12151 , n7555 );
    and g23074 ( n5837 , n9537 , n4832 );
    nor g23075 ( n2239 , n3506 , n9934 );
    or g23076 ( n7500 , n3385 , n11990 );
    or g23077 ( n18911 , n14572 , n25185 );
    nor g23078 ( n1531 , n21739 , n24805 );
    xnor g23079 ( n8936 , n1807 , n16053 );
    or g23080 ( n8114 , n1905 , n4618 );
    or g23081 ( n6036 , n5516 , n20125 );
    not g23082 ( n18078 , n9090 );
    xnor g23083 ( n1469 , n16711 , n14378 );
    or g23084 ( n11621 , n11791 , n16255 );
    xnor g23085 ( n20718 , n7057 , n14570 );
    and g23086 ( n1889 , n26855 , n23908 );
    xnor g23087 ( n23220 , n23044 , n1681 );
    or g23088 ( n13672 , n26797 , n18234 );
    xnor g23089 ( n9922 , n6477 , n1118 );
    or g23090 ( n16409 , n21700 , n1024 );
    or g23091 ( n16604 , n18841 , n20183 );
    xnor g23092 ( n1708 , n17490 , n7053 );
    or g23093 ( n7724 , n18058 , n12341 );
    xnor g23094 ( n10591 , n26216 , n16339 );
    or g23095 ( n26836 , n5651 , n17683 );
    xnor g23096 ( n26518 , n19489 , n12405 );
    not g23097 ( n19805 , n2723 );
    or g23098 ( n23155 , n203 , n8035 );
    not g23099 ( n10394 , n23224 );
    xnor g23100 ( n26927 , n18022 , n16746 );
    xnor g23101 ( n26380 , n11683 , n19015 );
    nor g23102 ( n7296 , n13590 , n23923 );
    or g23103 ( n556 , n5384 , n16899 );
    and g23104 ( n20312 , n8664 , n22616 );
    xnor g23105 ( n20253 , n9507 , n18409 );
    xnor g23106 ( n14657 , n19985 , n6104 );
    and g23107 ( n7803 , n14690 , n25399 );
    xnor g23108 ( n1541 , n21074 , n1470 );
    and g23109 ( n12804 , n11107 , n17657 );
    or g23110 ( n326 , n23860 , n18179 );
    xnor g23111 ( n10701 , n21660 , n23964 );
    not g23112 ( n27054 , n1819 );
    nor g23113 ( n5394 , n17610 , n4858 );
    or g23114 ( n23143 , n5229 , n18889 );
    or g23115 ( n5456 , n16057 , n12101 );
    or g23116 ( n19443 , n14856 , n9107 );
    not g23117 ( n18973 , n23454 );
    not g23118 ( n20638 , n20213 );
    not g23119 ( n24824 , n21508 );
    not g23120 ( n23313 , n1238 );
    xnor g23121 ( n21344 , n14354 , n22335 );
    xnor g23122 ( n8339 , n12710 , n17149 );
    and g23123 ( n9621 , n6087 , n13364 );
    or g23124 ( n4237 , n468 , n1255 );
    xnor g23125 ( n4481 , n12477 , n26408 );
    nor g23126 ( n983 , n8037 , n23636 );
    and g23127 ( n6910 , n1705 , n5354 );
    xnor g23128 ( n25905 , n8344 , n21654 );
    or g23129 ( n9267 , n932 , n2666 );
    xnor g23130 ( n3971 , n11941 , n8299 );
    or g23131 ( n15370 , n7013 , n7803 );
    and g23132 ( n5107 , n9677 , n12370 );
    not g23133 ( n26241 , n11356 );
    xnor g23134 ( n1004 , n16524 , n13668 );
    not g23135 ( n13339 , n23978 );
    xnor g23136 ( n18040 , n12255 , n14181 );
    nor g23137 ( n9118 , n25914 , n10275 );
    or g23138 ( n20640 , n162 , n20509 );
    and g23139 ( n734 , n22912 , n7484 );
    not g23140 ( n2056 , n24048 );
    xnor g23141 ( n7822 , n1451 , n26979 );
    xnor g23142 ( n19115 , n329 , n1163 );
    and g23143 ( n16138 , n26297 , n18948 );
    xnor g23144 ( n13612 , n4801 , n11970 );
    not g23145 ( n19742 , n3429 );
    nor g23146 ( n8908 , n24487 , n17184 );
    and g23147 ( n13948 , n5119 , n10639 );
    or g23148 ( n5951 , n1329 , n1898 );
    xnor g23149 ( n11375 , n6913 , n9500 );
    and g23150 ( n21133 , n10441 , n6727 );
    or g23151 ( n15811 , n16156 , n18997 );
    or g23152 ( n3170 , n15546 , n14702 );
    nor g23153 ( n2774 , n14632 , n1507 );
    xnor g23154 ( n109 , n9336 , n17969 );
    or g23155 ( n5038 , n20881 , n20492 );
    xnor g23156 ( n3472 , n11022 , n1955 );
    and g23157 ( n26607 , n16743 , n20020 );
    and g23158 ( n2877 , n4913 , n13489 );
    not g23159 ( n26215 , n4867 );
    or g23160 ( n1075 , n15647 , n13660 );
    xnor g23161 ( n2614 , n22173 , n12593 );
    xnor g23162 ( n13858 , n21974 , n22284 );
    or g23163 ( n22980 , n13783 , n6341 );
    or g23164 ( n26978 , n173 , n9380 );
    nor g23165 ( n15923 , n5751 , n8730 );
    xnor g23166 ( n5582 , n26176 , n423 );
    not g23167 ( n5652 , n19459 );
    or g23168 ( n7916 , n15309 , n1934 );
    not g23169 ( n17826 , n1163 );
    and g23170 ( n11124 , n23532 , n16716 );
    nor g23171 ( n2769 , n615 , n6944 );
    xnor g23172 ( n22047 , n19512 , n23984 );
    not g23173 ( n14764 , n25652 );
    and g23174 ( n21473 , n19831 , n15750 );
    xnor g23175 ( n4454 , n19926 , n21295 );
    and g23176 ( n12573 , n27117 , n8725 );
    not g23177 ( n6150 , n13841 );
    xnor g23178 ( n16499 , n13108 , n15258 );
    or g23179 ( n17406 , n24189 , n13217 );
    xnor g23180 ( n13984 , n17606 , n24936 );
    or g23181 ( n878 , n15138 , n22492 );
    and g23182 ( n2022 , n18409 , n25004 );
    xnor g23183 ( n3849 , n25924 , n18962 );
    and g23184 ( n16172 , n15357 , n14470 );
    xnor g23185 ( n22489 , n9795 , n2112 );
    not g23186 ( n14569 , n25435 );
    not g23187 ( n6273 , n9093 );
    and g23188 ( n1048 , n1066 , n9502 );
    and g23189 ( n15836 , n10056 , n20830 );
    nor g23190 ( n8066 , n18145 , n26191 );
    nor g23191 ( n15608 , n9398 , n24599 );
    and g23192 ( n22350 , n8313 , n13371 );
    or g23193 ( n2015 , n25888 , n24615 );
    or g23194 ( n22894 , n19712 , n21080 );
    buf g23195 ( n14289 , n23411 );
    and g23196 ( n22735 , n24958 , n10673 );
    xnor g23197 ( n2055 , n12901 , n27105 );
    xnor g23198 ( n19193 , n24143 , n12420 );
    not g23199 ( n17198 , n16319 );
    or g23200 ( n12608 , n18236 , n14069 );
    or g23201 ( n21712 , n20422 , n12335 );
    or g23202 ( n15097 , n19944 , n18962 );
    not g23203 ( n14654 , n24196 );
    or g23204 ( n16716 , n20496 , n15478 );
    xnor g23205 ( n7278 , n25302 , n19358 );
    or g23206 ( n11588 , n6124 , n26236 );
    xnor g23207 ( n2884 , n13979 , n6385 );
    xnor g23208 ( n7492 , n17088 , n17832 );
    or g23209 ( n2119 , n25324 , n12593 );
    xnor g23210 ( n6636 , n1630 , n9507 );
    or g23211 ( n18801 , n18659 , n3929 );
    xnor g23212 ( n26523 , n21379 , n19731 );
    nor g23213 ( n15727 , n2896 , n7773 );
    and g23214 ( n18716 , n19022 , n875 );
    xnor g23215 ( n8144 , n5747 , n9963 );
    or g23216 ( n16358 , n402 , n14380 );
    and g23217 ( n18590 , n14862 , n16442 );
    or g23218 ( n13385 , n10184 , n18006 );
    or g23219 ( n24958 , n11580 , n1469 );
    and g23220 ( n6411 , n23745 , n23053 );
    xnor g23221 ( n13257 , n24940 , n7719 );
    and g23222 ( n1490 , n26789 , n11733 );
    not g23223 ( n8568 , n2809 );
    xnor g23224 ( n5274 , n25114 , n16125 );
    not g23225 ( n22478 , n26584 );
    xnor g23226 ( n6734 , n26960 , n1394 );
    or g23227 ( n22312 , n13343 , n21286 );
    and g23228 ( n25961 , n8555 , n19021 );
    xnor g23229 ( n16615 , n22433 , n10158 );
    or g23230 ( n20672 , n10661 , n7076 );
    not g23231 ( n17295 , n16807 );
    xnor g23232 ( n687 , n12068 , n4558 );
    not g23233 ( n12 , n20575 );
    xnor g23234 ( n20629 , n23418 , n17207 );
    xnor g23235 ( n9032 , n22698 , n25147 );
    and g23236 ( n21218 , n11630 , n18504 );
    or g23237 ( n163 , n15122 , n16850 );
    or g23238 ( n23385 , n13446 , n5676 );
    xnor g23239 ( n25054 , n9530 , n7596 );
    or g23240 ( n8917 , n4100 , n26326 );
    xnor g23241 ( n19001 , n22554 , n26318 );
    xnor g23242 ( n4537 , n7699 , n4370 );
    xnor g23243 ( n23475 , n8102 , n20791 );
    xnor g23244 ( n23671 , n16203 , n12406 );
    or g23245 ( n10570 , n21479 , n22435 );
    or g23246 ( n7234 , n22347 , n24925 );
    or g23247 ( n21087 , n15952 , n24986 );
    not g23248 ( n2729 , n19751 );
    xnor g23249 ( n133 , n7769 , n25316 );
    xnor g23250 ( n4173 , n10980 , n5695 );
    xnor g23251 ( n8657 , n8457 , n23913 );
    or g23252 ( n6942 , n4418 , n21018 );
    or g23253 ( n2838 , n7048 , n13908 );
    xnor g23254 ( n13104 , n1836 , n5803 );
    xnor g23255 ( n4909 , n24939 , n24880 );
    nor g23256 ( n24562 , n8067 , n11243 );
    not g23257 ( n11596 , n8026 );
    nor g23258 ( n21703 , n17090 , n27120 );
    and g23259 ( n10781 , n3890 , n10384 );
    or g23260 ( n19768 , n14130 , n1097 );
    and g23261 ( n14855 , n20760 , n16151 );
    or g23262 ( n18564 , n6444 , n4404 );
    or g23263 ( n25865 , n23809 , n17209 );
    or g23264 ( n17914 , n18381 , n22073 );
    xnor g23265 ( n25622 , n1875 , n21258 );
    not g23266 ( n25486 , n11997 );
    and g23267 ( n16001 , n8883 , n9624 );
    xnor g23268 ( n25917 , n17548 , n1620 );
    or g23269 ( n25664 , n21517 , n16972 );
    and g23270 ( n14409 , n14195 , n19874 );
    and g23271 ( n22768 , n3984 , n22153 );
    xnor g23272 ( n9220 , n16804 , n22872 );
    nor g23273 ( n22256 , n18925 , n15185 );
    xnor g23274 ( n25288 , n24557 , n15630 );
    or g23275 ( n6228 , n13590 , n23529 );
    xnor g23276 ( n19882 , n17620 , n5330 );
    not g23277 ( n14276 , n92 );
    not g23278 ( n27074 , n4459 );
    xnor g23279 ( n18585 , n8830 , n11407 );
    or g23280 ( n24764 , n647 , n6475 );
    and g23281 ( n2221 , n18969 , n12206 );
    xnor g23282 ( n11070 , n24528 , n17487 );
    or g23283 ( n7461 , n13367 , n20970 );
    or g23284 ( n23350 , n24613 , n5269 );
    xnor g23285 ( n15108 , n20847 , n9415 );
    nor g23286 ( n5977 , n24796 , n15536 );
    or g23287 ( n267 , n1682 , n6427 );
    and g23288 ( n18342 , n222 , n13396 );
    xnor g23289 ( n5090 , n427 , n22198 );
    xnor g23290 ( n6558 , n7993 , n23232 );
    or g23291 ( n15704 , n5829 , n12344 );
    not g23292 ( n18360 , n24756 );
    or g23293 ( n14435 , n21678 , n684 );
    or g23294 ( n1747 , n22232 , n19271 );
    or g23295 ( n17714 , n19858 , n1984 );
    xnor g23296 ( n11347 , n10613 , n15721 );
    not g23297 ( n16211 , n17077 );
    xnor g23298 ( n949 , n5209 , n21358 );
    and g23299 ( n21088 , n21340 , n24266 );
    not g23300 ( n15442 , n5207 );
    and g23301 ( n21271 , n12562 , n12351 );
    and g23302 ( n13994 , n18324 , n24308 );
    and g23303 ( n25077 , n12840 , n26040 );
    not g23304 ( n4280 , n4916 );
    xnor g23305 ( n15889 , n3550 , n2652 );
    or g23306 ( n9660 , n24832 , n21050 );
    xnor g23307 ( n7679 , n23143 , n15783 );
    xnor g23308 ( n26136 , n21509 , n26090 );
    not g23309 ( n20127 , n10141 );
    not g23310 ( n17066 , n15282 );
    or g23311 ( n26560 , n22537 , n15902 );
    or g23312 ( n12624 , n26450 , n13088 );
    or g23313 ( n23210 , n2868 , n13455 );
    xnor g23314 ( n19383 , n26244 , n17051 );
    xnor g23315 ( n26141 , n1569 , n4560 );
    or g23316 ( n21952 , n6631 , n24732 );
    or g23317 ( n19100 , n13748 , n22704 );
    not g23318 ( n25150 , n23783 );
    and g23319 ( n8938 , n24489 , n7848 );
    or g23320 ( n26525 , n3813 , n8303 );
    xnor g23321 ( n23393 , n12878 , n22290 );
    xnor g23322 ( n14801 , n23944 , n2931 );
    and g23323 ( n16121 , n4881 , n24888 );
    and g23324 ( n16195 , n24646 , n4288 );
    not g23325 ( n20896 , n8485 );
    and g23326 ( n6214 , n18038 , n19627 );
    xnor g23327 ( n7466 , n7179 , n3229 );
    and g23328 ( n1452 , n17747 , n21364 );
    or g23329 ( n8388 , n20570 , n18474 );
    and g23330 ( n4705 , n12416 , n11069 );
    or g23331 ( n3991 , n23048 , n5795 );
    xnor g23332 ( n26600 , n7523 , n14440 );
    and g23333 ( n15059 , n1587 , n13303 );
    not g23334 ( n11309 , n21025 );
    or g23335 ( n17450 , n9368 , n2297 );
    and g23336 ( n23033 , n3815 , n12794 );
    nor g23337 ( n12651 , n22335 , n14354 );
    xnor g23338 ( n5028 , n7188 , n21237 );
    xnor g23339 ( n18398 , n13201 , n1353 );
    xnor g23340 ( n24271 , n25913 , n15568 );
    and g23341 ( n12628 , n16371 , n12523 );
    xnor g23342 ( n4519 , n10086 , n6175 );
    or g23343 ( n12970 , n20708 , n1608 );
    xnor g23344 ( n5749 , n23506 , n19789 );
    xnor g23345 ( n17780 , n14427 , n78 );
    xnor g23346 ( n21235 , n4879 , n6460 );
    and g23347 ( n4931 , n11157 , n8341 );
    not g23348 ( n9930 , n21002 );
    not g23349 ( n2557 , n16683 );
    or g23350 ( n3294 , n144 , n21764 );
    not g23351 ( n8016 , n19457 );
    not g23352 ( n5063 , n5739 );
    or g23353 ( n13586 , n10201 , n22379 );
    nor g23354 ( n23111 , n23048 , n2872 );
    xnor g23355 ( n5771 , n3744 , n13990 );
    xnor g23356 ( n18572 , n8445 , n8488 );
    xnor g23357 ( n15965 , n1171 , n3407 );
    xnor g23358 ( n5260 , n14485 , n9483 );
    xnor g23359 ( n23894 , n8663 , n3708 );
    and g23360 ( n17419 , n23436 , n21172 );
    xnor g23361 ( n5942 , n20766 , n21919 );
    and g23362 ( n18235 , n1166 , n4187 );
    not g23363 ( n2100 , n13216 );
    nor g23364 ( n5193 , n26774 , n22177 );
    xnor g23365 ( n17958 , n20053 , n24984 );
    xnor g23366 ( n5819 , n12709 , n3776 );
    nor g23367 ( n24540 , n7470 , n13696 );
    or g23368 ( n12318 , n1182 , n11652 );
    and g23369 ( n1830 , n4598 , n6771 );
    and g23370 ( n26532 , n4999 , n27017 );
    xnor g23371 ( n2198 , n15850 , n4714 );
    or g23372 ( n18640 , n20399 , n12695 );
    xnor g23373 ( n8770 , n17188 , n20225 );
    not g23374 ( n21306 , n494 );
    xnor g23375 ( n7572 , n20228 , n27154 );
    nor g23376 ( n13920 , n12464 , n20179 );
    xnor g23377 ( n24146 , n11453 , n21786 );
    nor g23378 ( n3868 , n7334 , n5925 );
    or g23379 ( n20830 , n9020 , n24957 );
    not g23380 ( n537 , n5605 );
    xnor g23381 ( n15171 , n16696 , n8638 );
    not g23382 ( n13975 , n15087 );
    or g23383 ( n6190 , n5313 , n17156 );
    xnor g23384 ( n3786 , n9331 , n13794 );
    xnor g23385 ( n423 , n2090 , n11926 );
    or g23386 ( n18273 , n6432 , n1045 );
    or g23387 ( n1038 , n4035 , n14602 );
    xnor g23388 ( n17885 , n19230 , n11580 );
    xnor g23389 ( n27175 , n19778 , n6423 );
    xnor g23390 ( n21430 , n4732 , n5286 );
    nor g23391 ( n10815 , n13349 , n13494 );
    xnor g23392 ( n3875 , n15271 , n26882 );
    xnor g23393 ( n17154 , n17835 , n8166 );
    nor g23394 ( n22740 , n8088 , n8624 );
    xnor g23395 ( n11998 , n23209 , n4485 );
    buf g23396 ( n4692 , n15277 );
    or g23397 ( n21414 , n5244 , n24340 );
    xnor g23398 ( n17891 , n725 , n17784 );
    or g23399 ( n318 , n21438 , n2291 );
    and g23400 ( n20600 , n832 , n19046 );
    nor g23401 ( n20988 , n3984 , n7439 );
    not g23402 ( n20065 , n23109 );
    or g23403 ( n2831 , n23039 , n12734 );
    nor g23404 ( n25870 , n11192 , n19805 );
    or g23405 ( n1664 , n16728 , n21884 );
    nor g23406 ( n13306 , n12956 , n11824 );
    or g23407 ( n25217 , n26599 , n4343 );
    and g23408 ( n20254 , n18603 , n13260 );
    xnor g23409 ( n20263 , n5668 , n1163 );
    or g23410 ( n1998 , n17484 , n25141 );
    and g23411 ( n17943 , n25282 , n25729 );
    or g23412 ( n3585 , n9065 , n3667 );
    or g23413 ( n9844 , n5624 , n14469 );
    xnor g23414 ( n2388 , n20310 , n551 );
    nor g23415 ( n17370 , n16824 , n26295 );
    not g23416 ( n19128 , n15250 );
    nor g23417 ( n176 , n2886 , n1738 );
    not g23418 ( n10455 , n13556 );
    or g23419 ( n15733 , n8841 , n14780 );
    xnor g23420 ( n132 , n12762 , n3349 );
    xnor g23421 ( n24187 , n19765 , n19081 );
    xnor g23422 ( n3770 , n14497 , n23593 );
    not g23423 ( n14754 , n17856 );
    xnor g23424 ( n7190 , n19491 , n6918 );
    and g23425 ( n23961 , n13404 , n14169 );
    and g23426 ( n8691 , n18122 , n6272 );
    xnor g23427 ( n7081 , n12855 , n13383 );
    and g23428 ( n17420 , n23570 , n9265 );
    not g23429 ( n16967 , n16739 );
    or g23430 ( n25774 , n17273 , n26392 );
    or g23431 ( n17624 , n17537 , n19280 );
    and g23432 ( n3462 , n20313 , n11641 );
    or g23433 ( n7103 , n19134 , n14385 );
    nor g23434 ( n9987 , n18729 , n13081 );
    xnor g23435 ( n20153 , n11051 , n342 );
    or g23436 ( n5554 , n6353 , n8434 );
    or g23437 ( n12618 , n8068 , n4466 );
    xnor g23438 ( n19210 , n21339 , n19802 );
    xnor g23439 ( n16862 , n8732 , n9285 );
    xnor g23440 ( n26226 , n24750 , n7872 );
    or g23441 ( n8004 , n2261 , n23653 );
    and g23442 ( n15685 , n7902 , n13926 );
    xnor g23443 ( n8418 , n17310 , n23974 );
    or g23444 ( n7909 , n14014 , n5189 );
    xnor g23445 ( n25503 , n8540 , n2399 );
    or g23446 ( n6795 , n7893 , n26876 );
    not g23447 ( n14598 , n17928 );
    xnor g23448 ( n13021 , n11044 , n4325 );
    or g23449 ( n3660 , n4132 , n23849 );
    xnor g23450 ( n23123 , n14306 , n10389 );
    or g23451 ( n16861 , n10788 , n21451 );
    xnor g23452 ( n2161 , n23700 , n26765 );
    nor g23453 ( n9627 , n6385 , n18171 );
    xnor g23454 ( n20382 , n13246 , n15039 );
    or g23455 ( n7220 , n11885 , n5361 );
    and g23456 ( n6186 , n2146 , n20216 );
    and g23457 ( n24830 , n21773 , n3375 );
    not g23458 ( n18300 , n12546 );
    or g23459 ( n17349 , n10903 , n20271 );
    and g23460 ( n25436 , n9995 , n21677 );
    or g23461 ( n7984 , n24516 , n2448 );
    xnor g23462 ( n11619 , n6502 , n19494 );
    and g23463 ( n11691 , n22554 , n2628 );
    not g23464 ( n21213 , n3382 );
    or g23465 ( n3254 , n4684 , n7183 );
    xnor g23466 ( n8947 , n3134 , n16285 );
    and g23467 ( n7771 , n18529 , n3858 );
    and g23468 ( n26139 , n23244 , n1801 );
    or g23469 ( n21554 , n25291 , n7061 );
    or g23470 ( n23458 , n10598 , n26360 );
    or g23471 ( n13782 , n18100 , n14155 );
    xnor g23472 ( n12419 , n19345 , n25574 );
    or g23473 ( n19582 , n6568 , n7055 );
    xnor g23474 ( n7805 , n9349 , n15547 );
    and g23475 ( n12333 , n24234 , n15460 );
    not g23476 ( n12859 , n22960 );
    not g23477 ( n19090 , n10903 );
    not g23478 ( n1605 , n14384 );
    or g23479 ( n680 , n16711 , n11011 );
    or g23480 ( n24997 , n18172 , n26278 );
    xnor g23481 ( n1450 , n12057 , n24638 );
    xnor g23482 ( n17388 , n20636 , n5214 );
    and g23483 ( n15569 , n14332 , n7916 );
    or g23484 ( n4137 , n4242 , n17388 );
    xnor g23485 ( n14599 , n22470 , n11455 );
    not g23486 ( n2808 , n8918 );
    nor g23487 ( n4796 , n21997 , n18483 );
    or g23488 ( n14892 , n141 , n7245 );
    not g23489 ( n3134 , n20291 );
    xnor g23490 ( n11949 , n13976 , n23895 );
    or g23491 ( n14065 , n3766 , n6074 );
    and g23492 ( n17389 , n25821 , n15510 );
    or g23493 ( n21551 , n88 , n14447 );
    or g23494 ( n15700 , n9574 , n13623 );
    xnor g23495 ( n21142 , n2782 , n1387 );
    and g23496 ( n20277 , n2371 , n14713 );
    not g23497 ( n19469 , n6502 );
    or g23498 ( n21958 , n13290 , n10730 );
    xnor g23499 ( n10638 , n3260 , n21832 );
    or g23500 ( n14262 , n2407 , n7538 );
    xnor g23501 ( n8825 , n10785 , n19042 );
    nor g23502 ( n26899 , n16803 , n25700 );
    xnor g23503 ( n16481 , n25488 , n17215 );
    not g23504 ( n3347 , n20055 );
    xnor g23505 ( n14274 , n2748 , n13808 );
    and g23506 ( n2538 , n13686 , n20034 );
    and g23507 ( n534 , n26732 , n19434 );
    and g23508 ( n9253 , n1718 , n20735 );
    and g23509 ( n9480 , n7766 , n5992 );
    nor g23510 ( n4505 , n5196 , n1878 );
    nor g23511 ( n13327 , n19184 , n14580 );
    and g23512 ( n2580 , n20638 , n10512 );
    not g23513 ( n14469 , n6553 );
    or g23514 ( n9618 , n24649 , n4426 );
    or g23515 ( n10560 , n9979 , n25948 );
    xnor g23516 ( n22444 , n21840 , n1555 );
    or g23517 ( n10103 , n21607 , n12726 );
    xnor g23518 ( n1705 , n16404 , n7323 );
    or g23519 ( n10662 , n20214 , n23241 );
    or g23520 ( n27061 , n25324 , n5951 );
    not g23521 ( n18759 , n22380 );
    xnor g23522 ( n17845 , n25046 , n23473 );
    and g23523 ( n24215 , n22436 , n100 );
    and g23524 ( n17850 , n1975 , n26527 );
    xnor g23525 ( n1757 , n3894 , n14993 );
    xnor g23526 ( n8848 , n20059 , n216 );
    xnor g23527 ( n15152 , n19175 , n16880 );
    xnor g23528 ( n5057 , n17578 , n8653 );
    xnor g23529 ( n14225 , n17613 , n10593 );
    nor g23530 ( n20297 , n19144 , n20210 );
    or g23531 ( n281 , n2146 , n22455 );
    not g23532 ( n7137 , n22092 );
    or g23533 ( n25857 , n6230 , n25235 );
    or g23534 ( n8476 , n27091 , n19317 );
    or g23535 ( n2029 , n22506 , n6047 );
    or g23536 ( n21265 , n14323 , n12351 );
    not g23537 ( n7879 , n14192 );
    xnor g23538 ( n6299 , n12354 , n12121 );
    or g23539 ( n13250 , n12134 , n21092 );
    or g23540 ( n11948 , n5950 , n17893 );
    and g23541 ( n19994 , n21454 , n4838 );
    xnor g23542 ( n12985 , n17242 , n336 );
    or g23543 ( n11683 , n11522 , n9327 );
    not g23544 ( n27189 , n23120 );
    not g23545 ( n12697 , n4045 );
    xnor g23546 ( n22375 , n9703 , n25871 );
    or g23547 ( n3095 , n17542 , n24402 );
    nor g23548 ( n13268 , n25738 , n11314 );
    and g23549 ( n11329 , n13986 , n23093 );
    not g23550 ( n8385 , n1047 );
    xnor g23551 ( n19296 , n26486 , n2816 );
    or g23552 ( n3892 , n3124 , n21832 );
    or g23553 ( n16592 , n15923 , n9817 );
    or g23554 ( n26456 , n23786 , n20942 );
    or g23555 ( n9949 , n18000 , n4732 );
    or g23556 ( n6723 , n13844 , n7516 );
    nor g23557 ( n26848 , n3140 , n14103 );
    nor g23558 ( n3957 , n7939 , n2925 );
    or g23559 ( n17222 , n5262 , n22712 );
    or g23560 ( n19189 , n3879 , n15978 );
    nor g23561 ( n14887 , n22194 , n19116 );
    xnor g23562 ( n17612 , n5050 , n1558 );
    and g23563 ( n3569 , n25491 , n26389 );
    or g23564 ( n18170 , n5360 , n21340 );
    xnor g23565 ( n12104 , n11248 , n26318 );
    and g23566 ( n25495 , n12150 , n11699 );
    xnor g23567 ( n24100 , n12098 , n21522 );
    and g23568 ( n18944 , n19910 , n18822 );
    and g23569 ( n12187 , n22324 , n18532 );
    and g23570 ( n15430 , n26582 , n7107 );
    or g23571 ( n21922 , n21127 , n20244 );
    xnor g23572 ( n5943 , n2701 , n9005 );
    not g23573 ( n23092 , n9747 );
    not g23574 ( n13042 , n24095 );
    not g23575 ( n22880 , n23331 );
    or g23576 ( n26611 , n13479 , n20343 );
    not g23577 ( n27 , n17308 );
    or g23578 ( n5691 , n12712 , n3003 );
    xnor g23579 ( n8229 , n14514 , n3694 );
    xnor g23580 ( n11239 , n21021 , n3253 );
    xnor g23581 ( n14110 , n26268 , n26285 );
    or g23582 ( n3047 , n23099 , n24444 );
    or g23583 ( n24163 , n21038 , n24645 );
    and g23584 ( n26172 , n3136 , n11542 );
    or g23585 ( n2109 , n15071 , n19748 );
    xnor g23586 ( n13936 , n26202 , n10712 );
    nor g23587 ( n22792 , n27060 , n25543 );
    xnor g23588 ( n5862 , n19839 , n19979 );
    not g23589 ( n5299 , n24922 );
    and g23590 ( n6213 , n16892 , n14686 );
    nor g23591 ( n3599 , n16544 , n4319 );
    not g23592 ( n18971 , n801 );
    nor g23593 ( n4073 , n10024 , n7347 );
    xnor g23594 ( n8535 , n1333 , n15927 );
    nor g23595 ( n1212 , n17090 , n22173 );
    xnor g23596 ( n18133 , n914 , n26167 );
    and g23597 ( n7293 , n18100 , n14569 );
    xnor g23598 ( n15081 , n13425 , n23580 );
    and g23599 ( n25148 , n17027 , n23206 );
    not g23600 ( n9924 , n16339 );
    or g23601 ( n2988 , n23010 , n11139 );
    or g23602 ( n23031 , n24078 , n21130 );
    not g23603 ( n12160 , n16521 );
    xnor g23604 ( n5416 , n19841 , n25140 );
    nor g23605 ( n24659 , n22588 , n13112 );
    nor g23606 ( n12631 , n25038 , n22442 );
    not g23607 ( n5621 , n15355 );
    xnor g23608 ( n10906 , n24042 , n17635 );
    not g23609 ( n14133 , n15967 );
    or g23610 ( n8800 , n22834 , n903 );
    xnor g23611 ( n22393 , n20409 , n18227 );
    or g23612 ( n21124 , n3909 , n24200 );
    nor g23613 ( n17494 , n11321 , n6703 );
    xnor g23614 ( n12324 , n24882 , n17312 );
    xnor g23615 ( n5011 , n18342 , n23045 );
    xnor g23616 ( n13881 , n25106 , n20921 );
    xnor g23617 ( n6576 , n25116 , n9346 );
    nor g23618 ( n951 , n8964 , n1293 );
    or g23619 ( n15347 , n7102 , n280 );
    not g23620 ( n1540 , n23831 );
    and g23621 ( n10374 , n26483 , n12088 );
    or g23622 ( n2451 , n4462 , n26286 );
    xnor g23623 ( n15064 , n24058 , n21287 );
    nor g23624 ( n14858 , n8155 , n767 );
    and g23625 ( n12032 , n6376 , n18939 );
    or g23626 ( n11343 , n13822 , n15077 );
    not g23627 ( n16468 , n25261 );
    or g23628 ( n6167 , n22713 , n7738 );
    xnor g23629 ( n11471 , n23018 , n11615 );
    xnor g23630 ( n18793 , n26818 , n14164 );
    and g23631 ( n20369 , n8722 , n10791 );
    nor g23632 ( n10587 , n18171 , n24529 );
    and g23633 ( n2317 , n1254 , n9056 );
    or g23634 ( n9902 , n20208 , n6732 );
    and g23635 ( n13570 , n25272 , n9785 );
    not g23636 ( n13057 , n3014 );
    and g23637 ( n18997 , n5953 , n13211 );
    not g23638 ( n19037 , n932 );
    and g23639 ( n15238 , n18148 , n12906 );
    not g23640 ( n11711 , n11473 );
    or g23641 ( n4843 , n26552 , n3337 );
    not g23642 ( n5998 , n25946 );
    not g23643 ( n15805 , n1227 );
    or g23644 ( n21557 , n12576 , n23463 );
    or g23645 ( n12755 , n23489 , n22766 );
    and g23646 ( n7371 , n19554 , n4281 );
    xnor g23647 ( n7388 , n12398 , n23586 );
    nor g23648 ( n22731 , n26241 , n12587 );
    xnor g23649 ( n15036 , n11989 , n14087 );
    or g23650 ( n6987 , n24862 , n14488 );
    or g23651 ( n14908 , n25875 , n4852 );
    xnor g23652 ( n4872 , n14315 , n18626 );
    xnor g23653 ( n162 , n25430 , n8116 );
    or g23654 ( n27081 , n6 , n21040 );
    xnor g23655 ( n21522 , n24087 , n20364 );
    and g23656 ( n20985 , n18569 , n14635 );
    and g23657 ( n1610 , n3090 , n16792 );
    or g23658 ( n9912 , n10050 , n17669 );
    xnor g23659 ( n16656 , n8817 , n12440 );
    or g23660 ( n26526 , n26495 , n26853 );
    not g23661 ( n483 , n1881 );
    or g23662 ( n8005 , n1444 , n3898 );
    or g23663 ( n18821 , n545 , n519 );
    xnor g23664 ( n11120 , n19786 , n22448 );
    or g23665 ( n1361 , n14714 , n3583 );
    or g23666 ( n26850 , n18400 , n6270 );
    buf g23667 ( n26417 , n26303 );
    or g23668 ( n17133 , n17632 , n16702 );
    or g23669 ( n5345 , n15474 , n21839 );
    xnor g23670 ( n18724 , n11614 , n9454 );
    xnor g23671 ( n16214 , n16661 , n23410 );
    xnor g23672 ( n23546 , n4385 , n25814 );
    or g23673 ( n17823 , n1443 , n7673 );
    not g23674 ( n125 , n16619 );
    or g23675 ( n9911 , n733 , n25067 );
    xnor g23676 ( n8380 , n8691 , n22546 );
    not g23677 ( n24821 , n18337 );
    xnor g23678 ( n16969 , n18869 , n10741 );
    or g23679 ( n10845 , n18986 , n2523 );
    or g23680 ( n20035 , n5696 , n7871 );
    not g23681 ( n17495 , n9269 );
    nor g23682 ( n8781 , n23369 , n26572 );
    or g23683 ( n22883 , n9840 , n20939 );
    or g23684 ( n1078 , n17974 , n13025 );
    xnor g23685 ( n7711 , n25074 , n6556 );
    and g23686 ( n25378 , n11678 , n6428 );
    xnor g23687 ( n3337 , n11767 , n18553 );
    or g23688 ( n5536 , n24341 , n6848 );
    xnor g23689 ( n15033 , n24883 , n21696 );
    or g23690 ( n22605 , n9671 , n12964 );
    xnor g23691 ( n25861 , n22515 , n12341 );
    xnor g23692 ( n1750 , n20408 , n23543 );
    xnor g23693 ( n14399 , n11736 , n22470 );
    xnor g23694 ( n5500 , n23697 , n9967 );
    not g23695 ( n12565 , n3631 );
    and g23696 ( n10521 , n24917 , n26983 );
    and g23697 ( n22257 , n22800 , n8075 );
    or g23698 ( n16391 , n10252 , n6102 );
    or g23699 ( n6812 , n19298 , n21038 );
    and g23700 ( n21484 , n3720 , n17262 );
    not g23701 ( n12396 , n15546 );
    xnor g23702 ( n14986 , n4278 , n18687 );
    or g23703 ( n13481 , n9365 , n1334 );
    nor g23704 ( n2709 , n6319 , n19836 );
    nor g23705 ( n19903 , n21972 , n9942 );
    and g23706 ( n1950 , n21649 , n20192 );
    or g23707 ( n4516 , n10576 , n11664 );
    xnor g23708 ( n6480 , n4685 , n21777 );
    xnor g23709 ( n12413 , n26722 , n18687 );
    nor g23710 ( n3058 , n5201 , n9932 );
    nor g23711 ( n22814 , n4719 , n12453 );
    and g23712 ( n6396 , n582 , n3163 );
    and g23713 ( n519 , n19288 , n12213 );
    xnor g23714 ( n12036 , n15008 , n15979 );
    not g23715 ( n24208 , n24154 );
    xnor g23716 ( n6138 , n22032 , n17866 );
    and g23717 ( n20968 , n6193 , n10070 );
    not g23718 ( n10659 , n10712 );
    not g23719 ( n12002 , n20250 );
    xnor g23720 ( n26194 , n9880 , n13714 );
    or g23721 ( n1254 , n2818 , n21390 );
    xnor g23722 ( n14738 , n24907 , n5822 );
    xnor g23723 ( n19263 , n3277 , n13628 );
    xnor g23724 ( n23089 , n2727 , n12214 );
    nor g23725 ( n22042 , n25475 , n13463 );
    xnor g23726 ( n24476 , n16526 , n4310 );
    or g23727 ( n21949 , n17688 , n17389 );
    and g23728 ( n23938 , n3047 , n10724 );
    or g23729 ( n10891 , n15298 , n14855 );
    xnor g23730 ( n9694 , n26797 , n15077 );
    or g23731 ( n8516 , n21101 , n13301 );
    xnor g23732 ( n13941 , n26379 , n19363 );
    nor g23733 ( n10438 , n3299 , n17141 );
    xnor g23734 ( n1266 , n24868 , n13747 );
    and g23735 ( n25196 , n12599 , n23777 );
    not g23736 ( n11784 , n21286 );
    not g23737 ( n11043 , n25629 );
    or g23738 ( n16789 , n25570 , n21747 );
    or g23739 ( n20286 , n23668 , n11769 );
    xnor g23740 ( n10347 , n22862 , n17663 );
    xnor g23741 ( n14763 , n10997 , n26619 );
    and g23742 ( n14287 , n694 , n6217 );
    xnor g23743 ( n5581 , n22034 , n7476 );
    nor g23744 ( n22971 , n5793 , n23710 );
    or g23745 ( n21600 , n1720 , n26212 );
    or g23746 ( n23224 , n7010 , n1547 );
    nor g23747 ( n22770 , n15636 , n24618 );
    not g23748 ( n16325 , n21240 );
    xnor g23749 ( n2051 , n23712 , n16753 );
    xnor g23750 ( n5200 , n19190 , n223 );
    xnor g23751 ( n9879 , n20146 , n5253 );
    or g23752 ( n19126 , n3396 , n9397 );
    xnor g23753 ( n4045 , n11850 , n21189 );
    and g23754 ( n27063 , n14633 , n2886 );
    not g23755 ( n5657 , n13781 );
    xnor g23756 ( n6443 , n10451 , n13677 );
    and g23757 ( n16966 , n2455 , n16564 );
    xnor g23758 ( n13788 , n2436 , n20391 );
    not g23759 ( n6682 , n3253 );
    nor g23760 ( n21483 , n14241 , n7418 );
    xnor g23761 ( n23180 , n10978 , n25126 );
    and g23762 ( n6762 , n21632 , n19423 );
    xnor g23763 ( n22448 , n11714 , n10861 );
    not g23764 ( n21929 , n21016 );
    and g23765 ( n22250 , n22017 , n22671 );
    xnor g23766 ( n3020 , n24430 , n19908 );
    xnor g23767 ( n9547 , n15291 , n13401 );
    not g23768 ( n3318 , n6427 );
    not g23769 ( n22295 , n13241 );
    not g23770 ( n8002 , n1483 );
    xnor g23771 ( n6065 , n18783 , n25908 );
    nor g23772 ( n26067 , n23253 , n26641 );
    xnor g23773 ( n16630 , n11984 , n25815 );
    and g23774 ( n25466 , n20411 , n17212 );
    and g23775 ( n7993 , n26626 , n3073 );
    xnor g23776 ( n14310 , n13305 , n5377 );
    or g23777 ( n9596 , n22065 , n9234 );
    nor g23778 ( n8566 , n17826 , n329 );
    or g23779 ( n13322 , n26294 , n15587 );
    or g23780 ( n21408 , n9828 , n11979 );
    or g23781 ( n25005 , n20142 , n17506 );
    and g23782 ( n568 , n25912 , n18104 );
    xnor g23783 ( n6302 , n8378 , n10633 );
    xnor g23784 ( n14074 , n21739 , n704 );
    and g23785 ( n9260 , n24054 , n14032 );
    not g23786 ( n4177 , n12271 );
    or g23787 ( n4814 , n739 , n4385 );
    not g23788 ( n3363 , n16029 );
    not g23789 ( n3707 , n12733 );
    or g23790 ( n3348 , n20425 , n15498 );
    xnor g23791 ( n18301 , n26638 , n18933 );
    not g23792 ( n21941 , n13161 );
    nor g23793 ( n7306 , n2858 , n13907 );
    or g23794 ( n20622 , n18662 , n9967 );
    not g23795 ( n19048 , n20833 );
    xnor g23796 ( n16583 , n16833 , n18963 );
    or g23797 ( n10154 , n9782 , n17520 );
    xnor g23798 ( n18478 , n13853 , n12274 );
    xnor g23799 ( n6207 , n7099 , n23068 );
    not g23800 ( n20482 , n17541 );
    xnor g23801 ( n14366 , n10524 , n58 );
    xnor g23802 ( n7474 , n7170 , n11945 );
    nor g23803 ( n5846 , n21929 , n6127 );
    xnor g23804 ( n19521 , n22735 , n21244 );
    and g23805 ( n8513 , n16233 , n25566 );
    and g23806 ( n11282 , n26996 , n6657 );
    not g23807 ( n14052 , n9069 );
    nor g23808 ( n19579 , n8614 , n12702 );
    not g23809 ( n17597 , n24213 );
    or g23810 ( n6570 , n13547 , n15601 );
    and g23811 ( n3889 , n24945 , n1516 );
    or g23812 ( n20423 , n19298 , n5816 );
    or g23813 ( n7629 , n8878 , n19122 );
    and g23814 ( n12668 , n4630 , n1073 );
    or g23815 ( n21939 , n22281 , n26332 );
    or g23816 ( n13258 , n20645 , n22577 );
    xnor g23817 ( n24353 , n5206 , n3990 );
    and g23818 ( n8199 , n2217 , n15038 );
    nor g23819 ( n6024 , n7893 , n18569 );
    and g23820 ( n1397 , n5872 , n7945 );
    and g23821 ( n17558 , n15156 , n21048 );
    xnor g23822 ( n3651 , n11890 , n27127 );
    xnor g23823 ( n27005 , n22173 , n583 );
    or g23824 ( n9936 , n24315 , n8268 );
    or g23825 ( n21776 , n22664 , n13524 );
    nor g23826 ( n6728 , n5509 , n21363 );
    buf g23827 ( n22861 , n21900 );
    or g23828 ( n14862 , n8568 , n13140 );
    and g23829 ( n11879 , n2745 , n4637 );
    xnor g23830 ( n26109 , n14133 , n7293 );
    xnor g23831 ( n12877 , n10170 , n19217 );
    nor g23832 ( n25863 , n3909 , n19081 );
    or g23833 ( n25491 , n5119 , n6070 );
    xnor g23834 ( n12835 , n22379 , n15077 );
    not g23835 ( n15456 , n21430 );
    and g23836 ( n1827 , n25673 , n7512 );
    xnor g23837 ( n15822 , n12351 , n12562 );
    xnor g23838 ( n22078 , n25643 , n329 );
    or g23839 ( n11883 , n17384 , n21077 );
    or g23840 ( n17464 , n13577 , n19229 );
    or g23841 ( n7541 , n2056 , n6104 );
    or g23842 ( n19299 , n27006 , n7197 );
    not g23843 ( n5505 , n15732 );
    or g23844 ( n8125 , n17826 , n26660 );
    or g23845 ( n19199 , n4286 , n14562 );
    xnor g23846 ( n21604 , n6729 , n11192 );
    xor g23847 ( n20570 , n11491 , n13826 );
    and g23848 ( n20460 , n12326 , n8446 );
    xnor g23849 ( n9051 , n24102 , n860 );
    xnor g23850 ( n2686 , n18262 , n18341 );
    xnor g23851 ( n12622 , n5992 , n2456 );
    xnor g23852 ( n10187 , n9402 , n2439 );
    or g23853 ( n22039 , n19898 , n17455 );
    xnor g23854 ( n21755 , n506 , n5386 );
    and g23855 ( n13029 , n25559 , n15714 );
    xnor g23856 ( n8661 , n3287 , n8573 );
    xnor g23857 ( n90 , n6442 , n25265 );
    xnor g23858 ( n2283 , n13649 , n5842 );
    xnor g23859 ( n18317 , n7532 , n8745 );
    or g23860 ( n11141 , n16054 , n17600 );
    not g23861 ( n26292 , n21352 );
    xnor g23862 ( n3590 , n25064 , n26427 );
    buf g23863 ( n20462 , n7387 );
    xnor g23864 ( n9430 , n19787 , n10643 );
    not g23865 ( n26030 , n13853 );
    xnor g23866 ( n1023 , n18495 , n2252 );
    and g23867 ( n5372 , n24192 , n929 );
    xnor g23868 ( n15535 , n2385 , n7130 );
    or g23869 ( n7445 , n9172 , n13665 );
    not g23870 ( n9988 , n25336 );
    and g23871 ( n5452 , n5966 , n13394 );
    not g23872 ( n3639 , n6474 );
    not g23873 ( n19094 , n24374 );
    xnor g23874 ( n8809 , n21376 , n4649 );
    xnor g23875 ( n5435 , n17255 , n17597 );
    and g23876 ( n462 , n11501 , n25509 );
    and g23877 ( n26373 , n11631 , n7398 );
    or g23878 ( n11590 , n24828 , n19368 );
    xnor g23879 ( n19307 , n2409 , n7057 );
    or g23880 ( n20992 , n1933 , n21200 );
    or g23881 ( n2627 , n9438 , n22192 );
    and g23882 ( n4926 , n8539 , n14610 );
    xnor g23883 ( n24119 , n8502 , n15488 );
    not g23884 ( n11363 , n7963 );
    or g23885 ( n9386 , n18995 , n7693 );
    xnor g23886 ( n14120 , n1403 , n5284 );
    xnor g23887 ( n10327 , n22184 , n11426 );
    or g23888 ( n15670 , n26565 , n10787 );
    nor g23889 ( n11690 , n5006 , n21117 );
    xnor g23890 ( n11022 , n23209 , n1319 );
    xnor g23891 ( n16098 , n23547 , n25569 );
    and g23892 ( n11614 , n9251 , n8344 );
    not g23893 ( n5407 , n21735 );
    or g23894 ( n13852 , n320 , n4906 );
    and g23895 ( n1384 , n1142 , n10294 );
    xnor g23896 ( n12516 , n24466 , n13595 );
    or g23897 ( n11231 , n11828 , n14032 );
    xnor g23898 ( n14810 , n8352 , n12859 );
    or g23899 ( n16100 , n4012 , n14264 );
    nor g23900 ( n25654 , n5143 , n9337 );
    xnor g23901 ( n24511 , n18615 , n25872 );
    buf g23902 ( n7361 , n26866 );
    nor g23903 ( n15703 , n19967 , n8245 );
    or g23904 ( n24710 , n4022 , n1009 );
    or g23905 ( n23357 , n8310 , n10309 );
    or g23906 ( n18460 , n18077 , n11782 );
    or g23907 ( n17861 , n6851 , n2656 );
    not g23908 ( n19592 , n18793 );
    xnor g23909 ( n502 , n8481 , n11998 );
    xnor g23910 ( n21132 , n13490 , n10739 );
    not g23911 ( n8411 , n11525 );
    or g23912 ( n2825 , n7832 , n9527 );
    not g23913 ( n1106 , n3447 );
    and g23914 ( n16515 , n9259 , n12423 );
    xnor g23915 ( n10295 , n25657 , n11091 );
    or g23916 ( n19826 , n8520 , n4375 );
    or g23917 ( n8449 , n5793 , n20361 );
    and g23918 ( n4055 , n19092 , n23734 );
    xnor g23919 ( n6460 , n7335 , n4319 );
    or g23920 ( n7082 , n15913 , n2037 );
    xor g23921 ( n17720 , n25101 , n27075 );
    and g23922 ( n13465 , n11748 , n7009 );
    and g23923 ( n1343 , n18269 , n12354 );
    or g23924 ( n25569 , n13049 , n5463 );
    not g23925 ( n23854 , n20898 );
    xnor g23926 ( n16447 , n22110 , n25485 );
    or g23927 ( n18937 , n8163 , n7173 );
    or g23928 ( n1235 , n13912 , n11098 );
    xnor g23929 ( n2964 , n24429 , n8314 );
    and g23930 ( n26301 , n7303 , n22946 );
    nor g23931 ( n4383 , n4160 , n12770 );
    or g23932 ( n20995 , n23351 , n24833 );
    nor g23933 ( n6697 , n5689 , n11864 );
    not g23934 ( n11303 , n8964 );
    or g23935 ( n21415 , n17347 , n13939 );
    not g23936 ( n14760 , n19404 );
    or g23937 ( n24968 , n6882 , n719 );
    and g23938 ( n23384 , n20420 , n23761 );
    or g23939 ( n7850 , n16722 , n16165 );
    xnor g23940 ( n25221 , n3583 , n20328 );
    nor g23941 ( n1526 , n8425 , n16184 );
    nor g23942 ( n24535 , n20687 , n8415 );
    xnor g23943 ( n4448 , n17795 , n15051 );
    xnor g23944 ( n8313 , n9036 , n18878 );
    nor g23945 ( n3907 , n7593 , n5101 );
    or g23946 ( n26057 , n16085 , n14160 );
    and g23947 ( n11782 , n753 , n20026 );
    or g23948 ( n21720 , n4347 , n22916 );
    nor g23949 ( n6919 , n12650 , n14765 );
    xnor g23950 ( n12355 , n18749 , n11980 );
    or g23951 ( n21241 , n7348 , n4435 );
    nor g23952 ( n24647 , n19062 , n14105 );
    or g23953 ( n22853 , n2798 , n2319 );
    not g23954 ( n5990 , n7338 );
    xnor g23955 ( n19709 , n20895 , n13373 );
    and g23956 ( n15637 , n26841 , n7011 );
    xnor g23957 ( n7372 , n16672 , n302 );
    xnor g23958 ( n4024 , n26695 , n3742 );
    or g23959 ( n24033 , n15503 , n8128 );
    nor g23960 ( n17052 , n15442 , n17382 );
    and g23961 ( n22192 , n18374 , n22966 );
    nor g23962 ( n26749 , n14265 , n15445 );
    xnor g23963 ( n1418 , n7953 , n20908 );
    xnor g23964 ( n19728 , n6718 , n1611 );
    not g23965 ( n19192 , n25261 );
    xnor g23966 ( n22099 , n12880 , n18446 );
    not g23967 ( n26499 , n12973 );
    or g23968 ( n19954 , n6726 , n18202 );
    xnor g23969 ( n5782 , n18009 , n13466 );
    nor g23970 ( n10413 , n23878 , n5139 );
    not g23971 ( n14415 , n15271 );
    and g23972 ( n10449 , n10825 , n9304 );
    not g23973 ( n17734 , n26641 );
    or g23974 ( n22890 , n19875 , n9737 );
    and g23975 ( n8832 , n24369 , n25894 );
    xnor g23976 ( n19517 , n7082 , n20593 );
    not g23977 ( n17770 , n10232 );
    or g23978 ( n14638 , n5159 , n11377 );
    and g23979 ( n25497 , n20805 , n16289 );
    xnor g23980 ( n27100 , n12854 , n26867 );
    or g23981 ( n1282 , n13719 , n22342 );
    or g23982 ( n24442 , n9294 , n17568 );
    or g23983 ( n21010 , n17098 , n12622 );
    xnor g23984 ( n21860 , n23952 , n4631 );
    nor g23985 ( n14596 , n27203 , n24959 );
    or g23986 ( n16395 , n353 , n22119 );
    or g23987 ( n15871 , n25122 , n13349 );
    nor g23988 ( n22204 , n5112 , n20954 );
    xnor g23989 ( n1819 , n22305 , n17102 );
    not g23990 ( n104 , n17380 );
    or g23991 ( n2186 , n16620 , n15599 );
    xnor g23992 ( n14170 , n7824 , n16654 );
    or g23993 ( n22718 , n14718 , n20920 );
    not g23994 ( n12586 , n21293 );
    or g23995 ( n12969 , n1018 , n22306 );
    or g23996 ( n26379 , n23560 , n21069 );
    or g23997 ( n341 , n407 , n9717 );
    not g23998 ( n19849 , n19163 );
    nor g23999 ( n15676 , n24018 , n5400 );
    xnor g24000 ( n24105 , n11571 , n4725 );
    nor g24001 ( n19927 , n7184 , n20564 );
    or g24002 ( n2569 , n11628 , n2166 );
    or g24003 ( n12752 , n15925 , n1123 );
    xnor g24004 ( n619 , n4348 , n13157 );
    not g24005 ( n19298 , n583 );
    or g24006 ( n6615 , n11581 , n14994 );
    or g24007 ( n7123 , n23602 , n820 );
    or g24008 ( n25814 , n26402 , n11879 );
    and g24009 ( n10960 , n7185 , n5698 );
    or g24010 ( n26991 , n5067 , n8344 );
    and g24011 ( n21069 , n8081 , n21619 );
    or g24012 ( n26616 , n14873 , n3644 );
    or g24013 ( n12599 , n12258 , n1626 );
    nor g24014 ( n5952 , n23566 , n9457 );
    and g24015 ( n23931 , n612 , n17329 );
    or g24016 ( n8864 , n6953 , n7282 );
    or g24017 ( n20742 , n26180 , n24700 );
    or g24018 ( n11153 , n22977 , n20923 );
    and g24019 ( n22338 , n13892 , n16974 );
    and g24020 ( n10318 , n5226 , n21205 );
    not g24021 ( n9814 , n4675 );
    xnor g24022 ( n9210 , n12491 , n8154 );
    xnor g24023 ( n21570 , n20468 , n13453 );
    or g24024 ( n16953 , n25463 , n20526 );
    or g24025 ( n24505 , n15378 , n10039 );
    and g24026 ( n11707 , n13349 , n24422 );
    xnor g24027 ( n23471 , n9629 , n1431 );
    or g24028 ( n26034 , n3094 , n6284 );
    and g24029 ( n24137 , n14647 , n23381 );
    nor g24030 ( n6721 , n22644 , n10642 );
    not g24031 ( n20032 , n19005 );
    xnor g24032 ( n26681 , n20580 , n19727 );
    nor g24033 ( n17385 , n23863 , n25381 );
    xnor g24034 ( n5263 , n13130 , n24491 );
    xnor g24035 ( n1857 , n15404 , n18599 );
    xnor g24036 ( n25375 , n5443 , n1320 );
    and g24037 ( n10708 , n8096 , n14748 );
    xnor g24038 ( n14135 , n17881 , n8067 );
    xnor g24039 ( n9289 , n14569 , n24732 );
    or g24040 ( n15357 , n5122 , n12395 );
    or g24041 ( n8460 , n12524 , n1287 );
    not g24042 ( n4574 , n26180 );
    or g24043 ( n6796 , n212 , n2783 );
    and g24044 ( n8128 , n8967 , n26533 );
    xnor g24045 ( n2083 , n20970 , n12961 );
    not g24046 ( n10220 , n17671 );
    and g24047 ( n15308 , n25447 , n770 );
    xnor g24048 ( n20244 , n4588 , n22201 );
    and g24049 ( n25285 , n16772 , n14286 );
    xnor g24050 ( n4596 , n23832 , n19238 );
    nor g24051 ( n14441 , n7421 , n13206 );
    or g24052 ( n9848 , n24357 , n3699 );
    nor g24053 ( n9546 , n8614 , n21698 );
    not g24054 ( n8609 , n24499 );
    not g24055 ( n24420 , n25696 );
    nor g24056 ( n16932 , n11802 , n7627 );
    not g24057 ( n25724 , n26866 );
    nor g24058 ( n11679 , n14774 , n26300 );
    and g24059 ( n236 , n7973 , n15179 );
    nor g24060 ( n6192 , n20036 , n22515 );
    xnor g24061 ( n21425 , n6865 , n6703 );
    not g24062 ( n684 , n24616 );
    xnor g24063 ( n26718 , n22828 , n379 );
    nor g24064 ( n16429 , n25772 , n21596 );
    xnor g24065 ( n23341 , n10270 , n13801 );
    and g24066 ( n24776 , n3579 , n5667 );
    or g24067 ( n17608 , n328 , n19387 );
    nor g24068 ( n9592 , n1831 , n10250 );
    xnor g24069 ( n5844 , n16846 , n24101 );
    or g24070 ( n4546 , n708 , n2781 );
    xnor g24071 ( n14181 , n3707 , n12802 );
    or g24072 ( n19428 , n21272 , n8769 );
    xnor g24073 ( n12980 , n8725 , n15065 );
    and g24074 ( n11815 , n13868 , n6441 );
    and g24075 ( n25167 , n11612 , n27085 );
    and g24076 ( n23891 , n12521 , n3787 );
    or g24077 ( n18169 , n12091 , n25076 );
    and g24078 ( n20776 , n2849 , n20641 );
    and g24079 ( n3004 , n11001 , n22611 );
    xnor g24080 ( n24998 , n23933 , n17269 );
    xnor g24081 ( n18046 , n15097 , n6893 );
    xnor g24082 ( n946 , n13633 , n13171 );
    and g24083 ( n12480 , n22515 , n10467 );
    nor g24084 ( n8562 , n26695 , n22588 );
    not g24085 ( n8528 , n6333 );
    or g24086 ( n25950 , n26633 , n2900 );
    nor g24087 ( n8348 , n13172 , n16252 );
    xnor g24088 ( n25412 , n5099 , n14216 );
    or g24089 ( n4557 , n22396 , n17980 );
    xnor g24090 ( n13596 , n24032 , n22843 );
    or g24091 ( n26051 , n19214 , n13705 );
    not g24092 ( n24850 , n26882 );
    and g24093 ( n12984 , n24890 , n18303 );
    not g24094 ( n6131 , n18487 );
    not g24095 ( n5938 , n6229 );
    or g24096 ( n5755 , n5666 , n5232 );
    and g24097 ( n22921 , n7381 , n16198 );
    and g24098 ( n11689 , n6534 , n7009 );
    and g24099 ( n11867 , n6854 , n26702 );
    xnor g24100 ( n19663 , n14060 , n6287 );
    xnor g24101 ( n5285 , n1544 , n7052 );
    nor g24102 ( n6023 , n21226 , n586 );
    xnor g24103 ( n22779 , n6472 , n12938 );
    nor g24104 ( n21883 , n3356 , n16311 );
    not g24105 ( n1403 , n25470 );
    and g24106 ( n6690 , n22001 , n3886 );
    xnor g24107 ( n20484 , n4665 , n8309 );
    not g24108 ( n21337 , n8250 );
    xnor g24109 ( n19174 , n1607 , n3234 );
    nor g24110 ( n24470 , n23572 , n18474 );
    or g24111 ( n6868 , n25610 , n10984 );
    xnor g24112 ( n3673 , n26861 , n22160 );
    xnor g24113 ( n7585 , n627 , n4166 );
    or g24114 ( n21773 , n21134 , n4930 );
    xnor g24115 ( n22427 , n8918 , n19365 );
    and g24116 ( n1762 , n3346 , n8044 );
    and g24117 ( n20654 , n7524 , n14133 );
    not g24118 ( n2242 , n6498 );
    or g24119 ( n22438 , n26391 , n2009 );
    or g24120 ( n17896 , n16427 , n17888 );
    xnor g24121 ( n24973 , n18539 , n3366 );
    not g24122 ( n23832 , n18201 );
    xnor g24123 ( n1835 , n19745 , n15160 );
    or g24124 ( n26272 , n22197 , n21164 );
    and g24125 ( n6830 , n5471 , n2864 );
    not g24126 ( n832 , n19789 );
    or g24127 ( n23042 , n26670 , n2206 );
    or g24128 ( n1017 , n6177 , n22833 );
    not g24129 ( n10758 , n20570 );
    nor g24130 ( n5276 , n11011 , n20179 );
    xnor g24131 ( n1301 , n4873 , n23272 );
    or g24132 ( n3701 , n2777 , n11517 );
    nor g24133 ( n23474 , n342 , n26789 );
    xnor g24134 ( n9806 , n20735 , n3463 );
    xnor g24135 ( n16682 , n13342 , n25660 );
    or g24136 ( n5121 , n25903 , n9659 );
    nor g24137 ( n787 , n2383 , n15236 );
    nor g24138 ( n22622 , n18452 , n6397 );
    nor g24139 ( n1725 , n4844 , n13708 );
    or g24140 ( n21582 , n13026 , n13906 );
    and g24141 ( n4074 , n24236 , n19289 );
    xnor g24142 ( n303 , n832 , n19046 );
    and g24143 ( n21427 , n23708 , n6013 );
    or g24144 ( n7663 , n22223 , n731 );
    or g24145 ( n8914 , n14991 , n24638 );
    nor g24146 ( n1383 , n7389 , n7531 );
    not g24147 ( n17266 , n7569 );
    and g24148 ( n4571 , n7458 , n4763 );
    nor g24149 ( n16472 , n11560 , n7080 );
    or g24150 ( n8984 , n8166 , n7554 );
    xnor g24151 ( n22130 , n14103 , n19402 );
    and g24152 ( n2180 , n13976 , n25419 );
    or g24153 ( n10607 , n1224 , n10727 );
    or g24154 ( n20686 , n26107 , n21636 );
    not g24155 ( n23642 , n19240 );
    or g24156 ( n814 , n889 , n13874 );
    nor g24157 ( n26314 , n19457 , n1753 );
    not g24158 ( n19545 , n18507 );
    xnor g24159 ( n4634 , n3480 , n19911 );
    xnor g24160 ( n12330 , n7173 , n13511 );
    or g24161 ( n8555 , n17690 , n17235 );
    xnor g24162 ( n24840 , n14667 , n804 );
    not g24163 ( n8979 , n21779 );
    xnor g24164 ( n7467 , n10406 , n8947 );
    xnor g24165 ( n26665 , n18737 , n2328 );
    xnor g24166 ( n14809 , n17579 , n12452 );
    or g24167 ( n25242 , n3740 , n23683 );
    nor g24168 ( n1273 , n25915 , n8024 );
    xor g24169 ( n25251 , n10930 , n10626 );
    nor g24170 ( n14228 , n18690 , n1183 );
    xnor g24171 ( n20207 , n3498 , n3740 );
    xnor g24172 ( n16082 , n2291 , n21438 );
    xnor g24173 ( n11459 , n8064 , n1240 );
    and g24174 ( n10160 , n21651 , n18460 );
    xnor g24175 ( n2518 , n11327 , n26752 );
    xnor g24176 ( n6433 , n13926 , n25864 );
    xnor g24177 ( n58 , n22660 , n11011 );
    xnor g24178 ( n15404 , n21109 , n5224 );
    or g24179 ( n6957 , n8990 , n13108 );
    nor g24180 ( n4871 , n19157 , n22793 );
    not g24181 ( n623 , n25008 );
    not g24182 ( n126 , n23801 );
    nor g24183 ( n18818 , n16205 , n23068 );
    not g24184 ( n5675 , n26303 );
    and g24185 ( n8353 , n3386 , n22742 );
    and g24186 ( n4648 , n15945 , n25824 );
    xnor g24187 ( n24433 , n21420 , n11086 );
    xnor g24188 ( n21017 , n26115 , n16898 );
    nor g24189 ( n20642 , n9003 , n13453 );
    or g24190 ( n22746 , n5766 , n12382 );
    nor g24191 ( n20211 , n23273 , n10435 );
    or g24192 ( n7710 , n5115 , n2548 );
    and g24193 ( n4328 , n17921 , n4402 );
    nor g24194 ( n13999 , n12587 , n10608 );
    or g24195 ( n19091 , n12649 , n7865 );
    xnor g24196 ( n16870 , n9934 , n2272 );
    not g24197 ( n19265 , n24156 );
    xnor g24198 ( n3143 , n24865 , n11040 );
    and g24199 ( n24789 , n13238 , n17058 );
    xnor g24200 ( n12423 , n26039 , n9554 );
    not g24201 ( n1574 , n8661 );
    not g24202 ( n19025 , n13074 );
    or g24203 ( n4511 , n5355 , n5000 );
    not g24204 ( n8343 , n22253 );
    nor g24205 ( n4081 , n9655 , n22700 );
    and g24206 ( n3759 , n12042 , n11308 );
    xnor g24207 ( n10549 , n21737 , n24020 );
    xnor g24208 ( n2719 , n13357 , n11077 );
    nor g24209 ( n16877 , n1095 , n1367 );
    or g24210 ( n13868 , n9550 , n16203 );
    and g24211 ( n1487 , n14329 , n26157 );
    not g24212 ( n11452 , n20179 );
    nor g24213 ( n4683 , n18754 , n19245 );
    or g24214 ( n23700 , n26448 , n2200 );
    xnor g24215 ( n25513 , n5965 , n11241 );
    or g24216 ( n20183 , n6743 , n5969 );
    not g24217 ( n17013 , n24879 );
    xnor g24218 ( n11245 , n16749 , n20418 );
    and g24219 ( n8201 , n23049 , n10621 );
    and g24220 ( n4399 , n1661 , n15106 );
    and g24221 ( n541 , n10862 , n26005 );
    or g24222 ( n24871 , n22959 , n2529 );
    not g24223 ( n12675 , n6894 );
    xnor g24224 ( n24592 , n27053 , n19501 );
    or g24225 ( n12904 , n4208 , n20083 );
    and g24226 ( n23101 , n21531 , n25098 );
    nor g24227 ( n6871 , n9535 , n11846 );
    not g24228 ( n15562 , n19097 );
    xnor g24229 ( n9961 , n21305 , n7544 );
    xnor g24230 ( n16273 , n11694 , n25810 );
    xnor g24231 ( n10287 , n9743 , n10296 );
    and g24232 ( n23204 , n6190 , n21870 );
    xnor g24233 ( n19311 , n23906 , n8846 );
    not g24234 ( n111 , n22738 );
    or g24235 ( n8102 , n8501 , n25809 );
    nor g24236 ( n25527 , n27199 , n6861 );
    nor g24237 ( n9899 , n17458 , n20687 );
    xnor g24238 ( n10919 , n9582 , n299 );
    and g24239 ( n7125 , n13682 , n22357 );
    and g24240 ( n7178 , n7995 , n18917 );
    and g24241 ( n20591 , n10189 , n23975 );
    or g24242 ( n21453 , n157 , n16235 );
    or g24243 ( n19519 , n859 , n24982 );
    xnor g24244 ( n13703 , n21567 , n3306 );
    xnor g24245 ( n8632 , n7524 , n19680 );
    not g24246 ( n7205 , n4314 );
    not g24247 ( n27066 , n6949 );
    nor g24248 ( n19024 , n27037 , n13775 );
    and g24249 ( n6665 , n22786 , n2921 );
    nor g24250 ( n11847 , n21733 , n1753 );
    or g24251 ( n9801 , n19157 , n6555 );
    or g24252 ( n13639 , n13126 , n25103 );
    or g24253 ( n19684 , n17115 , n2418 );
    or g24254 ( n19957 , n22252 , n15256 );
    not g24255 ( n13301 , n2586 );
    xnor g24256 ( n20485 , n21624 , n20944 );
    not g24257 ( n2820 , n15124 );
    or g24258 ( n3353 , n17292 , n5078 );
    not g24259 ( n11118 , n21284 );
    or g24260 ( n19022 , n12048 , n11688 );
    xnor g24261 ( n18571 , n12875 , n22492 );
    and g24262 ( n2128 , n15419 , n12087 );
    or g24263 ( n12244 , n11579 , n3962 );
    or g24264 ( n8116 , n12933 , n4987 );
    or g24265 ( n6404 , n25068 , n10620 );
    not g24266 ( n8897 , n1893 );
    nor g24267 ( n26370 , n20150 , n26187 );
    not g24268 ( n20907 , n4748 );
    xnor g24269 ( n8382 , n6083 , n9922 );
    or g24270 ( n16987 , n3959 , n25917 );
    or g24271 ( n10530 , n16839 , n19030 );
    and g24272 ( n24408 , n20615 , n20225 );
    or g24273 ( n22127 , n12116 , n10742 );
    or g24274 ( n11932 , n25698 , n10674 );
    not g24275 ( n20972 , n5324 );
    not g24276 ( n2926 , n1092 );
    nor g24277 ( n23347 , n4894 , n2566 );
    or g24278 ( n8433 , n19469 , n25625 );
    nor g24279 ( n5645 , n23110 , n7058 );
    nor g24280 ( n23753 , n9586 , n3279 );
    xnor g24281 ( n16449 , n5080 , n11262 );
    or g24282 ( n4453 , n8455 , n24835 );
    or g24283 ( n16981 , n12259 , n7197 );
    or g24284 ( n26011 , n1127 , n17528 );
    xnor g24285 ( n2429 , n4111 , n17723 );
    xnor g24286 ( n8371 , n2749 , n25464 );
    nor g24287 ( n23184 , n17819 , n23970 );
    xnor g24288 ( n10612 , n4256 , n18483 );
    xnor g24289 ( n26800 , n7787 , n10333 );
    xnor g24290 ( n17625 , n167 , n3554 );
    xnor g24291 ( n12836 , n17993 , n7674 );
    and g24292 ( n15596 , n3068 , n17521 );
    and g24293 ( n23840 , n11642 , n16042 );
    or g24294 ( n13398 , n10276 , n23654 );
    nor g24295 ( n20324 , n17454 , n8389 );
    or g24296 ( n22495 , n83 , n13663 );
    buf g24297 ( n17635 , n18024 );
    or g24298 ( n1692 , n5263 , n9160 );
    or g24299 ( n18083 , n19310 , n7499 );
    or g24300 ( n931 , n920 , n11618 );
    not g24301 ( n11062 , n8823 );
    xnor g24302 ( n23910 , n24296 , n6174 );
    xnor g24303 ( n16455 , n7727 , n24363 );
    not g24304 ( n24560 , n12086 );
    nor g24305 ( n12348 , n5587 , n111 );
    xnor g24306 ( n13915 , n5947 , n14440 );
    and g24307 ( n12277 , n21856 , n24163 );
    and g24308 ( n7152 , n25212 , n127 );
    or g24309 ( n261 , n8538 , n20971 );
    or g24310 ( n21763 , n25094 , n24586 );
    not g24311 ( n23218 , n1183 );
    and g24312 ( n4820 , n3320 , n17579 );
    xnor g24313 ( n9378 , n5573 , n2201 );
    or g24314 ( n23397 , n9872 , n26726 );
    or g24315 ( n1788 , n6309 , n14999 );
    or g24316 ( n5447 , n12446 , n966 );
    not g24317 ( n1898 , n26556 );
    nor g24318 ( n20165 , n25886 , n8399 );
    nor g24319 ( n22062 , n10372 , n12152 );
    or g24320 ( n20569 , n6086 , n3197 );
    xnor g24321 ( n6160 , n4786 , n25222 );
    or g24322 ( n9533 , n16825 , n17703 );
    or g24323 ( n12370 , n2299 , n5792 );
    and g24324 ( n11073 , n6878 , n22280 );
    xnor g24325 ( n21262 , n21460 , n18079 );
    nor g24326 ( n18776 , n15000 , n16106 );
    not g24327 ( n18032 , n3299 );
    not g24328 ( n12810 , n20906 );
    and g24329 ( n16917 , n4897 , n26819 );
    and g24330 ( n4096 , n15702 , n26500 );
    and g24331 ( n19349 , n22522 , n17876 );
    or g24332 ( n14712 , n26615 , n4025 );
    xnor g24333 ( n10169 , n23137 , n11617 );
    xnor g24334 ( n17298 , n25276 , n12341 );
    xnor g24335 ( n18840 , n21537 , n18031 );
    xnor g24336 ( n19866 , n13190 , n9318 );
    xnor g24337 ( n13171 , n16007 , n12821 );
    or g24338 ( n11208 , n20329 , n6397 );
    not g24339 ( n9332 , n9886 );
    xnor g24340 ( n11148 , n7437 , n1662 );
    nor g24341 ( n8983 , n6877 , n874 );
    xnor g24342 ( n10984 , n21274 , n19191 );
    and g24343 ( n22137 , n3660 , n8040 );
    or g24344 ( n2754 , n21261 , n18204 );
    or g24345 ( n13861 , n15796 , n12446 );
    not g24346 ( n19722 , n5176 );
    xnor g24347 ( n2552 , n5313 , n14274 );
    xnor g24348 ( n4467 , n14134 , n20253 );
    not g24349 ( n17674 , n8820 );
    not g24350 ( n2606 , n4939 );
    or g24351 ( n11454 , n13517 , n9522 );
    and g24352 ( n15977 , n25926 , n9646 );
    xnor g24353 ( n17476 , n5938 , n7212 );
    nor g24354 ( n11913 , n23244 , n5128 );
    xnor g24355 ( n12214 , n9345 , n19941 );
    nor g24356 ( n24627 , n22755 , n7503 );
    xnor g24357 ( n10219 , n21211 , n917 );
    xnor g24358 ( n1410 , n20249 , n17902 );
    or g24359 ( n26751 , n7353 , n19730 );
    xnor g24360 ( n8669 , n26660 , n18907 );
    not g24361 ( n21386 , n12657 );
    or g24362 ( n3386 , n25872 , n19618 );
    not g24363 ( n17586 , n16543 );
    not g24364 ( n10527 , n7276 );
    xnor g24365 ( n20917 , n12679 , n11039 );
    or g24366 ( n22901 , n8960 , n12187 );
    xnor g24367 ( n24801 , n22757 , n24870 );
    and g24368 ( n19769 , n8049 , n7446 );
    xnor g24369 ( n8079 , n19860 , n2785 );
    nor g24370 ( n16186 , n26417 , n10509 );
    not g24371 ( n16561 , n18227 );
    and g24372 ( n2638 , n16161 , n2093 );
    or g24373 ( n23813 , n2196 , n1059 );
    or g24374 ( n23465 , n2669 , n347 );
    or g24375 ( n19710 , n2187 , n5832 );
    nor g24376 ( n6592 , n13590 , n1792 );
    xnor g24377 ( n8706 , n13960 , n9493 );
    or g24378 ( n16927 , n1036 , n10967 );
    xnor g24379 ( n9889 , n10666 , n9489 );
    or g24380 ( n3272 , n7017 , n1889 );
    and g24381 ( n13509 , n3310 , n18627 );
    xnor g24382 ( n26870 , n26278 , n5042 );
    xnor g24383 ( n18487 , n23824 , n9730 );
    and g24384 ( n16933 , n20984 , n250 );
    nor g24385 ( n8191 , n23034 , n24684 );
    xnor g24386 ( n21579 , n14187 , n7162 );
    xnor g24387 ( n3471 , n17683 , n5552 );
    or g24388 ( n20522 , n10565 , n23806 );
    and g24389 ( n1126 , n6310 , n20672 );
    and g24390 ( n17775 , n19344 , n14497 );
    xnor g24391 ( n14501 , n21162 , n10018 );
    and g24392 ( n22520 , n26210 , n20380 );
    or g24393 ( n8640 , n9600 , n7578 );
    xnor g24394 ( n11986 , n19693 , n20197 );
    xnor g24395 ( n2623 , n1662 , n3710 );
    and g24396 ( n8996 , n22764 , n26830 );
    or g24397 ( n5544 , n7238 , n14923 );
    xnor g24398 ( n3845 , n5342 , n17559 );
    not g24399 ( n7481 , n7028 );
    xnor g24400 ( n26196 , n18183 , n23071 );
    not g24401 ( n5624 , n12446 );
    nor g24402 ( n17334 , n20077 , n3952 );
    and g24403 ( n3860 , n25909 , n9153 );
    not g24404 ( n12563 , n21725 );
    and g24405 ( n8245 , n24983 , n19278 );
    or g24406 ( n1877 , n4315 , n23200 );
    or g24407 ( n16964 , n12038 , n22070 );
    xnor g24408 ( n22684 , n11822 , n12811 );
    nor g24409 ( n11829 , n20455 , n2884 );
    xnor g24410 ( n14868 , n10097 , n9564 );
    xnor g24411 ( n19648 , n26275 , n26937 );
    xnor g24412 ( n11390 , n10902 , n9952 );
    not g24413 ( n25021 , n19701 );
    or g24414 ( n9541 , n22762 , n24846 );
    xnor g24415 ( n19500 , n5211 , n12811 );
    xnor g24416 ( n2209 , n23817 , n15299 );
    xnor g24417 ( n20621 , n15733 , n18692 );
    xnor g24418 ( n24128 , n5976 , n2694 );
    nor g24419 ( n14933 , n23755 , n23509 );
    or g24420 ( n23929 , n8566 , n24619 );
    and g24421 ( n8956 , n26839 , n9667 );
    xnor g24422 ( n19542 , n3780 , n17276 );
    xnor g24423 ( n18231 , n13696 , n25514 );
    and g24424 ( n5598 , n882 , n26097 );
    xnor g24425 ( n6925 , n13030 , n71 );
    xnor g24426 ( n791 , n19122 , n23632 );
    nor g24427 ( n21181 , n10893 , n9817 );
    xnor g24428 ( n3846 , n4196 , n11415 );
    or g24429 ( n6053 , n4871 , n815 );
    xnor g24430 ( n18972 , n23931 , n19020 );
    and g24431 ( n10358 , n6773 , n20089 );
    nor g24432 ( n18018 , n11630 , n3783 );
    not g24433 ( n880 , n1513 );
    and g24434 ( n23128 , n12541 , n3412 );
    or g24435 ( n22929 , n20883 , n5859 );
    xnor g24436 ( n18634 , n23340 , n7570 );
    not g24437 ( n17926 , n9218 );
    or g24438 ( n16253 , n23981 , n17709 );
    xnor g24439 ( n17232 , n12026 , n10672 );
    nor g24440 ( n15295 , n10405 , n8241 );
    or g24441 ( n8307 , n17087 , n16092 );
    or g24442 ( n17777 , n6325 , n27161 );
    and g24443 ( n24225 , n14227 , n15968 );
    not g24444 ( n17087 , n3694 );
    and g24445 ( n7574 , n7724 , n3322 );
    nor g24446 ( n24760 , n216 , n20059 );
    or g24447 ( n7367 , n25139 , n7974 );
    or g24448 ( n2410 , n18017 , n15582 );
    and g24449 ( n11064 , n15766 , n7465 );
    xnor g24450 ( n23727 , n21393 , n3935 );
    and g24451 ( n3532 , n5444 , n18748 );
    nor g24452 ( n17507 , n25846 , n7546 );
    xnor g24453 ( n13691 , n10611 , n2680 );
    xnor g24454 ( n26007 , n21338 , n27010 );
    and g24455 ( n11205 , n7099 , n18888 );
    xnor g24456 ( n21717 , n3609 , n24148 );
    not g24457 ( n8859 , n17294 );
    xnor g24458 ( n3810 , n2161 , n5924 );
    xnor g24459 ( n10279 , n2410 , n6230 );
    xnor g24460 ( n4520 , n26535 , n4198 );
    xnor g24461 ( n11910 , n21033 , n9441 );
    or g24462 ( n5151 , n16529 , n20005 );
    xnor g24463 ( n1414 , n474 , n12104 );
    or g24464 ( n16985 , n3981 , n1741 );
    and g24465 ( n12185 , n19056 , n22854 );
    xnor g24466 ( n22744 , n23155 , n14456 );
    or g24467 ( n25849 , n20652 , n2890 );
    nor g24468 ( n942 , n15258 , n2420 );
    or g24469 ( n23476 , n22123 , n18078 );
    not g24470 ( n26437 , n264 );
    or g24471 ( n13538 , n7693 , n15644 );
    or g24472 ( n9731 , n23629 , n25648 );
    nor g24473 ( n2212 , n23234 , n20138 );
    buf g24474 ( n15659 , n3002 );
    not g24475 ( n788 , n14816 );
    xnor g24476 ( n24464 , n26857 , n1881 );
    or g24477 ( n18675 , n6915 , n15996 );
    or g24478 ( n26612 , n212 , n2146 );
    xnor g24479 ( n25264 , n17716 , n25475 );
    or g24480 ( n12796 , n25440 , n20644 );
    nor g24481 ( n20113 , n15271 , n26748 );
    and g24482 ( n14722 , n24638 , n19327 );
    or g24483 ( n23893 , n15086 , n13927 );
    and g24484 ( n15095 , n523 , n9912 );
    xnor g24485 ( n9206 , n20551 , n8283 );
    xnor g24486 ( n17538 , n21527 , n26174 );
    or g24487 ( n18366 , n20544 , n22652 );
    and g24488 ( n24088 , n1767 , n3250 );
    xnor g24489 ( n18765 , n22769 , n21839 );
    and g24490 ( n21882 , n9657 , n19275 );
    and g24491 ( n4341 , n19110 , n26753 );
    and g24492 ( n8733 , n7225 , n26352 );
    or g24493 ( n12517 , n2131 , n11809 );
    or g24494 ( n4091 , n27092 , n2052 );
    not g24495 ( n5203 , n7377 );
    or g24496 ( n7473 , n14790 , n26075 );
    xnor g24497 ( n2078 , n24165 , n15842 );
    and g24498 ( n16715 , n12309 , n4013 );
    xnor g24499 ( n26160 , n14487 , n53 );
    and g24500 ( n7110 , n25544 , n18184 );
    and g24501 ( n11003 , n18842 , n26487 );
    or g24502 ( n4021 , n3025 , n9137 );
    nor g24503 ( n10928 , n9570 , n1667 );
    not g24504 ( n14385 , n9748 );
    nor g24505 ( n14785 , n23863 , n14702 );
    and g24506 ( n16658 , n10405 , n12198 );
    and g24507 ( n26266 , n21652 , n5225 );
    nor g24508 ( n321 , n16846 , n24101 );
    nor g24509 ( n22794 , n9416 , n17587 );
    xnor g24510 ( n3524 , n12316 , n20340 );
    and g24511 ( n18823 , n4085 , n16547 );
    and g24512 ( n23306 , n9493 , n15507 );
    nor g24513 ( n10754 , n11534 , n8659 );
    xnor g24514 ( n9110 , n25935 , n15817 );
    xnor g24515 ( n26515 , n26973 , n24533 );
    xnor g24516 ( n1498 , n7078 , n17012 );
    nor g24517 ( n23173 , n18880 , n26594 );
    or g24518 ( n10814 , n13326 , n2293 );
    and g24519 ( n5922 , n16029 , n4322 );
    and g24520 ( n23294 , n21558 , n18783 );
    not g24521 ( n16213 , n18429 );
    xnor g24522 ( n24203 , n2576 , n15532 );
    and g24523 ( n21236 , n6446 , n20060 );
    xnor g24524 ( n21479 , n347 , n4346 );
    nor g24525 ( n21663 , n8399 , n6834 );
    not g24526 ( n9856 , n24392 );
    xnor g24527 ( n3377 , n26667 , n16183 );
    and g24528 ( n4677 , n12535 , n4705 );
    xnor g24529 ( n7031 , n4326 , n14148 );
    not g24530 ( n10378 , n1090 );
    or g24531 ( n6007 , n9018 , n18047 );
    xnor g24532 ( n4927 , n5330 , n919 );
    xnor g24533 ( n19314 , n6719 , n11967 );
    not g24534 ( n18995 , n7566 );
    xnor g24535 ( n1351 , n10160 , n8229 );
    xnor g24536 ( n3289 , n14844 , n16862 );
    or g24537 ( n6770 , n27202 , n15085 );
    xnor g24538 ( n4393 , n27095 , n2160 );
    xnor g24539 ( n17243 , n9408 , n11431 );
    xnor g24540 ( n22385 , n22012 , n13387 );
    and g24541 ( n17992 , n19875 , n9737 );
    not g24542 ( n13214 , n9170 );
    or g24543 ( n16461 , n26370 , n10782 );
    and g24544 ( n24067 , n15780 , n24358 );
    and g24545 ( n16487 , n8880 , n5975 );
    not g24546 ( n14870 , n12470 );
    xnor g24547 ( n18549 , n18799 , n10763 );
    or g24548 ( n25992 , n15186 , n26928 );
    or g24549 ( n25780 , n15712 , n12571 );
    xnor g24550 ( n17115 , n21185 , n27165 );
    nor g24551 ( n15371 , n17790 , n9651 );
    xnor g24552 ( n25467 , n20411 , n9512 );
    nor g24553 ( n13814 , n24116 , n23408 );
    or g24554 ( n14520 , n20137 , n1662 );
    and g24555 ( n22336 , n17162 , n868 );
    not g24556 ( n23359 , n2979 );
    or g24557 ( n13289 , n10323 , n25785 );
    xnor g24558 ( n14174 , n16425 , n19356 );
    xnor g24559 ( n22667 , n13249 , n25156 );
    and g24560 ( n2448 , n12590 , n16270 );
    not g24561 ( n26090 , n25608 );
    xnor g24562 ( n22903 , n20439 , n17114 );
    xnor g24563 ( n8716 , n4830 , n19740 );
    or g24564 ( n10811 , n9791 , n13462 );
    and g24565 ( n19479 , n25535 , n16546 );
    or g24566 ( n26354 , n10534 , n24896 );
    xnor g24567 ( n17808 , n22748 , n24128 );
    xnor g24568 ( n3121 , n18888 , n7099 );
    nor g24569 ( n7224 , n10124 , n8897 );
    xnor g24570 ( n5876 , n2036 , n23630 );
    xnor g24571 ( n1240 , n27120 , n11192 );
    xnor g24572 ( n16215 , n19637 , n11297 );
    nor g24573 ( n19445 , n5682 , n10468 );
    or g24574 ( n6920 , n22454 , n10710 );
    or g24575 ( n1142 , n10191 , n15792 );
    and g24576 ( n26574 , n14040 , n24711 );
    not g24577 ( n10849 , n18551 );
    or g24578 ( n19939 , n20032 , n19144 );
    xnor g24579 ( n19060 , n21387 , n12487 );
    xnor g24580 ( n12141 , n18438 , n26672 );
    or g24581 ( n1395 , n22843 , n4155 );
    xnor g24582 ( n19752 , n835 , n13668 );
    not g24583 ( n18090 , n18649 );
    xnor g24584 ( n27154 , n14365 , n2804 );
    or g24585 ( n13211 , n26153 , n11372 );
    not g24586 ( n20537 , n4597 );
    xnor g24587 ( n7787 , n21453 , n4273 );
    and g24588 ( n810 , n3107 , n26941 );
    not g24589 ( n10097 , n19589 );
    and g24590 ( n20656 , n12007 , n23377 );
    and g24591 ( n16113 , n4498 , n19766 );
    and g24592 ( n5010 , n14012 , n7774 );
    nor g24593 ( n15196 , n22240 , n2375 );
    xnor g24594 ( n25140 , n910 , n12891 );
    nor g24595 ( n14698 , n1307 , n25219 );
    xnor g24596 ( n6216 , n19886 , n14091 );
    not g24597 ( n2312 , n12687 );
    or g24598 ( n23622 , n17137 , n11689 );
    not g24599 ( n22009 , n24458 );
    and g24600 ( n21635 , n14538 , n23862 );
    nor g24601 ( n15667 , n10751 , n27009 );
    nor g24602 ( n17642 , n21915 , n24919 );
    or g24603 ( n1488 , n22559 , n19995 );
    not g24604 ( n6284 , n2320 );
    or g24605 ( n8655 , n16594 , n17351 );
    or g24606 ( n13598 , n15026 , n5063 );
    xnor g24607 ( n10834 , n10187 , n26331 );
    xnor g24608 ( n24517 , n22840 , n11765 );
    and g24609 ( n11491 , n13380 , n2067 );
    or g24610 ( n19353 , n6543 , n1720 );
    xnor g24611 ( n1348 , n5220 , n6948 );
    xnor g24612 ( n9005 , n4572 , n23581 );
    not g24613 ( n22015 , n21784 );
    not g24614 ( n12128 , n25623 );
    not g24615 ( n16529 , n16536 );
    and g24616 ( n6644 , n7463 , n16821 );
    not g24617 ( n4143 , n17415 );
    or g24618 ( n10072 , n11805 , n20426 );
    and g24619 ( n13298 , n16401 , n7861 );
    not g24620 ( n5194 , n3072 );
    not g24621 ( n21230 , n14058 );
    nor g24622 ( n21057 , n25692 , n729 );
    xnor g24623 ( n2326 , n25052 , n25895 );
    nor g24624 ( n10071 , n10267 , n12592 );
    or g24625 ( n13697 , n8963 , n24041 );
    or g24626 ( n4171 , n13337 , n7200 );
    or g24627 ( n16566 , n23419 , n22951 );
    or g24628 ( n11359 , n20410 , n7365 );
    and g24629 ( n10143 , n937 , n15733 );
    xnor g24630 ( n21897 , n23920 , n5231 );
    nor g24631 ( n4902 , n16524 , n20923 );
    xnor g24632 ( n21707 , n586 , n15274 );
    and g24633 ( n15154 , n19019 , n16408 );
    or g24634 ( n15472 , n3682 , n5339 );
    nor g24635 ( n2511 , n19589 , n9564 );
    not g24636 ( n21975 , n3955 );
    not g24637 ( n10610 , n18599 );
    or g24638 ( n21667 , n4087 , n808 );
    xnor g24639 ( n17524 , n3167 , n6001 );
    not g24640 ( n6240 , n13090 );
    and g24641 ( n5210 , n24598 , n14006 );
    or g24642 ( n15870 , n3877 , n23034 );
    or g24643 ( n19677 , n1573 , n4652 );
    and g24644 ( n6732 , n22499 , n3331 );
    not g24645 ( n2713 , n21471 );
    xnor g24646 ( n17696 , n18409 , n3952 );
    or g24647 ( n23732 , n18027 , n4866 );
    not g24648 ( n9974 , n5910 );
    or g24649 ( n9573 , n17741 , n10451 );
    xnor g24650 ( n20340 , n16345 , n4542 );
    and g24651 ( n23977 , n24891 , n7878 );
    xnor g24652 ( n14811 , n15442 , n6015 );
    not g24653 ( n15935 , n5587 );
    nor g24654 ( n19511 , n19646 , n8277 );
    not g24655 ( n20771 , n8085 );
    xnor g24656 ( n24533 , n15236 , n2383 );
    not g24657 ( n12815 , n3976 );
    and g24658 ( n20031 , n22056 , n20817 );
    not g24659 ( n13114 , n17037 );
    xnor g24660 ( n25655 , n26986 , n2272 );
    xnor g24661 ( n9742 , n13783 , n9942 );
    or g24662 ( n10206 , n20365 , n14127 );
    nor g24663 ( n26469 , n13898 , n25004 );
    and g24664 ( n18268 , n5360 , n21340 );
    and g24665 ( n19016 , n22976 , n21958 );
    and g24666 ( n22059 , n9793 , n22361 );
    and g24667 ( n12647 , n2933 , n372 );
    or g24668 ( n25284 , n13044 , n4038 );
    and g24669 ( n20394 , n5489 , n16342 );
    not g24670 ( n7353 , n6307 );
    and g24671 ( n26009 , n20346 , n9315 );
    and g24672 ( n6406 , n543 , n2244 );
    not g24673 ( n12258 , n23200 );
    or g24674 ( n4046 , n22271 , n19417 );
    and g24675 ( n13620 , n21265 , n23266 );
    or g24676 ( n19991 , n14718 , n6814 );
    and g24677 ( n13592 , n14955 , n13098 );
    xnor g24678 ( n17731 , n12875 , n7751 );
    nor g24679 ( n22055 , n1685 , n9514 );
    xnor g24680 ( n5383 , n11056 , n20478 );
    and g24681 ( n20321 , n22962 , n10567 );
    or g24682 ( n24652 , n13967 , n18972 );
    or g24683 ( n19369 , n1215 , n23715 );
    xnor g24684 ( n14064 , n5506 , n2331 );
    not g24685 ( n5180 , n22698 );
    and g24686 ( n7104 , n23836 , n7562 );
    xnor g24687 ( n19365 , n390 , n5060 );
    and g24688 ( n22653 , n7763 , n1627 );
    xnor g24689 ( n16797 , n20437 , n26565 );
    and g24690 ( n21283 , n9880 , n20273 );
    xnor g24691 ( n11741 , n24243 , n26044 );
    and g24692 ( n588 , n16089 , n9316 );
    nor g24693 ( n27093 , n144 , n5960 );
    xnor g24694 ( n20774 , n11588 , n21098 );
    nor g24695 ( n4133 , n4194 , n8795 );
    xnor g24696 ( n16886 , n14287 , n585 );
    and g24697 ( n13559 , n13117 , n20084 );
    not g24698 ( n25697 , n2989 );
    and g24699 ( n1619 , n22687 , n11734 );
    xnor g24700 ( n16895 , n22197 , n5927 );
    and g24701 ( n21862 , n9644 , n17894 );
    nor g24702 ( n5688 , n22379 , n22207 );
    nor g24703 ( n14950 , n12137 , n10258 );
    xnor g24704 ( n23871 , n25100 , n23765 );
    xnor g24705 ( n19845 , n23604 , n15328 );
    nor g24706 ( n203 , n21759 , n5445 );
    and g24707 ( n26397 , n22331 , n9203 );
    xnor g24708 ( n24857 , n6002 , n20107 );
    or g24709 ( n26739 , n25558 , n13668 );
    or g24710 ( n24354 , n15995 , n516 );
    and g24711 ( n6080 , n19799 , n15112 );
    xnor g24712 ( n19877 , n2783 , n6785 );
    not g24713 ( n4941 , n20707 );
    or g24714 ( n15916 , n7952 , n1136 );
    or g24715 ( n3640 , n1300 , n14567 );
    or g24716 ( n18777 , n13171 , n13633 );
    or g24717 ( n3507 , n10147 , n15169 );
    or g24718 ( n20306 , n16086 , n7105 );
    not g24719 ( n1687 , n679 );
    or g24720 ( n24123 , n25112 , n18084 );
    nor g24721 ( n19703 , n1202 , n4246 );
    or g24722 ( n11760 , n23920 , n23344 );
    or g24723 ( n23604 , n20676 , n19400 );
    and g24724 ( n20493 , n10693 , n19167 );
    xnor g24725 ( n23575 , n20409 , n1099 );
    xnor g24726 ( n7270 , n19123 , n18208 );
    xnor g24727 ( n8626 , n19508 , n21234 );
    xnor g24728 ( n11591 , n2654 , n10979 );
    not g24729 ( n2718 , n1413 );
    xnor g24730 ( n18698 , n16793 , n18428 );
    xnor g24731 ( n21759 , n806 , n4051 );
    xnor g24732 ( n14597 , n23655 , n23755 );
    xnor g24733 ( n9293 , n4467 , n9752 );
    xnor g24734 ( n14534 , n2966 , n19627 );
    xnor g24735 ( n11888 , n18861 , n22091 );
    xnor g24736 ( n14319 , n7105 , n3543 );
    and g24737 ( n6776 , n21089 , n13224 );
    and g24738 ( n26385 , n16316 , n9279 );
    nor g24739 ( n24754 , n25733 , n19498 );
    xnor g24740 ( n9346 , n7824 , n22808 );
    xnor g24741 ( n17652 , n2447 , n9089 );
    not g24742 ( n21249 , n14999 );
    xnor g24743 ( n19276 , n16627 , n6765 );
    xnor g24744 ( n13194 , n3239 , n6648 );
    or g24745 ( n14650 , n21138 , n14230 );
    xnor g24746 ( n2132 , n2939 , n6366 );
    or g24747 ( n217 , n5719 , n14130 );
    not g24748 ( n2628 , n25381 );
    xnor g24749 ( n2244 , n1496 , n7502 );
    xnor g24750 ( n7314 , n18785 , n14096 );
    nor g24751 ( n3525 , n2858 , n5521 );
    or g24752 ( n16745 , n8381 , n20382 );
    not g24753 ( n25220 , n24988 );
    xnor g24754 ( n25585 , n3675 , n5145 );
    and g24755 ( n2658 , n10522 , n23024 );
    xnor g24756 ( n26463 , n163 , n13015 );
    xnor g24757 ( n22870 , n26761 , n22080 );
    xnor g24758 ( n10001 , n22774 , n1611 );
    xnor g24759 ( n21585 , n11558 , n2280 );
    or g24760 ( n11861 , n1923 , n9200 );
    xnor g24761 ( n25952 , n25015 , n15131 );
    and g24762 ( n512 , n10565 , n23806 );
    and g24763 ( n24275 , n3482 , n25374 );
    xnor g24764 ( n23799 , n11858 , n17885 );
    xnor g24765 ( n19767 , n16878 , n19835 );
    nor g24766 ( n24966 , n18976 , n15090 );
    or g24767 ( n19965 , n23867 , n12296 );
    xnor g24768 ( n19132 , n6165 , n12201 );
    and g24769 ( n6782 , n1437 , n17784 );
    xnor g24770 ( n17743 , n115 , n2355 );
    or g24771 ( n25306 , n19355 , n8153 );
    or g24772 ( n6755 , n5233 , n7214 );
    xnor g24773 ( n894 , n1742 , n4590 );
    xnor g24774 ( n11997 , n5196 , n4491 );
    xnor g24775 ( n19233 , n20024 , n6088 );
    xnor g24776 ( n18799 , n7869 , n14968 );
    not g24777 ( n2412 , n8041 );
    and g24778 ( n25683 , n13644 , n3712 );
    xnor g24779 ( n18263 , n1148 , n17810 );
    xnor g24780 ( n9550 , n19952 , n10178 );
    not g24781 ( n424 , n22047 );
    and g24782 ( n11333 , n6394 , n9273 );
    xnor g24783 ( n21517 , n5959 , n9835 );
    or g24784 ( n20463 , n2281 , n1047 );
    xnor g24785 ( n19089 , n12495 , n15780 );
    nor g24786 ( n15213 , n8989 , n12162 );
    not g24787 ( n3376 , n9455 );
    not g24788 ( n25103 , n10229 );
    xnor g24789 ( n6168 , n16403 , n13008 );
    xnor g24790 ( n2651 , n9283 , n6633 );
    or g24791 ( n15060 , n7593 , n25317 );
    or g24792 ( n26623 , n5013 , n5305 );
    xnor g24793 ( n11488 , n15294 , n5538 );
    not g24794 ( n11178 , n17485 );
    or g24795 ( n2955 , n3161 , n18201 );
    xnor g24796 ( n6835 , n11931 , n17229 );
    or g24797 ( n15466 , n4692 , n15775 );
    or g24798 ( n13954 , n120 , n4939 );
    or g24799 ( n25976 , n8891 , n7406 );
    xnor g24800 ( n7212 , n13554 , n7004 );
    and g24801 ( n22826 , n6081 , n15434 );
    and g24802 ( n8659 , n17776 , n8512 );
    or g24803 ( n3237 , n793 , n12736 );
    or g24804 ( n25319 , n11030 , n6141 );
    nor g24805 ( n10757 , n8363 , n1222 );
    and g24806 ( n5644 , n12365 , n20306 );
    xnor g24807 ( n12767 , n13378 , n10444 );
    or g24808 ( n5775 , n1705 , n9456 );
    or g24809 ( n7912 , n7391 , n24134 );
    nor g24810 ( n3312 , n12522 , n8308 );
    xnor g24811 ( n7610 , n14929 , n2132 );
    or g24812 ( n14439 , n1404 , n14684 );
    and g24813 ( n5425 , n20893 , n18128 );
    or g24814 ( n5127 , n24620 , n21753 );
    or g24815 ( n20186 , n12398 , n25696 );
    xnor g24816 ( n8753 , n21138 , n20385 );
    and g24817 ( n10753 , n5313 , n17156 );
    xnor g24818 ( n94 , n24808 , n13860 );
    xnor g24819 ( n24483 , n24034 , n26885 );
    nor g24820 ( n17484 , n26471 , n22382 );
    or g24821 ( n25717 , n21566 , n14343 );
    or g24822 ( n717 , n8368 , n7504 );
    xnor g24823 ( n7547 , n6861 , n5255 );
    xnor g24824 ( n23903 , n17700 , n1728 );
    xnor g24825 ( n6020 , n8853 , n23036 );
    or g24826 ( n5177 , n20120 , n9313 );
    or g24827 ( n6272 , n7639 , n11703 );
    or g24828 ( n3883 , n22288 , n24023 );
    or g24829 ( n14263 , n14051 , n290 );
    nor g24830 ( n846 , n13494 , n3425 );
    xnor g24831 ( n14952 , n22634 , n17816 );
    xnor g24832 ( n6175 , n10888 , n14176 );
    not g24833 ( n6393 , n22619 );
    and g24834 ( n23674 , n9773 , n26163 );
    nor g24835 ( n13629 , n3659 , n17635 );
    xnor g24836 ( n26504 , n11694 , n18040 );
    xnor g24837 ( n5126 , n7935 , n18608 );
    xnor g24838 ( n3870 , n2462 , n21150 );
    or g24839 ( n23836 , n16439 , n10275 );
    xnor g24840 ( n772 , n2498 , n14185 );
    and g24841 ( n4741 , n10191 , n15792 );
    nor g24842 ( n20042 , n5938 , n960 );
    and g24843 ( n2154 , n25047 , n1381 );
    xnor g24844 ( n22488 , n27037 , n13775 );
    xnor g24845 ( n2510 , n21326 , n12623 );
    xor g24846 ( n9252 , n25855 , n24714 );
    xnor g24847 ( n8962 , n11146 , n17095 );
    and g24848 ( n9473 , n21091 , n13415 );
    xnor g24849 ( n25087 , n14790 , n342 );
    xnor g24850 ( n9714 , n17590 , n17549 );
    or g24851 ( n4757 , n13300 , n17000 );
    xnor g24852 ( n13352 , n652 , n16181 );
    nor g24853 ( n17973 , n24187 , n19331 );
    or g24854 ( n6563 , n8966 , n12128 );
    xnor g24855 ( n4436 , n769 , n16280 );
    or g24856 ( n13068 , n23932 , n9380 );
    xnor g24857 ( n19798 , n10630 , n18876 );
    or g24858 ( n12791 , n1838 , n14127 );
    or g24859 ( n16134 , n5292 , n25144 );
    or g24860 ( n1035 , n20853 , n10238 );
    or g24861 ( n9155 , n19138 , n13066 );
    not g24862 ( n5119 , n26641 );
    or g24863 ( n21895 , n18345 , n22700 );
    not g24864 ( n11366 , n8233 );
    and g24865 ( n23019 , n16157 , n16343 );
    or g24866 ( n22869 , n22775 , n20895 );
    not g24867 ( n7447 , n19045 );
    or g24868 ( n11956 , n18430 , n10764 );
    or g24869 ( n11916 , n9654 , n23057 );
    not g24870 ( n5261 , n8718 );
    or g24871 ( n12520 , n22003 , n23705 );
    and g24872 ( n16883 , n20319 , n25046 );
    xnor g24873 ( n20351 , n20049 , n12610 );
    not g24874 ( n23573 , n7260 );
    and g24875 ( n22506 , n7523 , n23686 );
    xnor g24876 ( n24646 , n8486 , n22592 );
    xnor g24877 ( n1231 , n4602 , n21337 );
    xnor g24878 ( n25332 , n23152 , n1909 );
    xnor g24879 ( n16808 , n19757 , n8126 );
    xnor g24880 ( n19425 , n6360 , n15970 );
    or g24881 ( n1595 , n11186 , n23878 );
    or g24882 ( n8747 , n15932 , n8728 );
    xnor g24883 ( n18864 , n25845 , n18497 );
    not g24884 ( n14306 , n9851 );
    xor g24885 ( n12700 , n3790 , n11192 );
    and g24886 ( n5051 , n1251 , n23595 );
    not g24887 ( n19084 , n22154 );
    and g24888 ( n6413 , n10966 , n3420 );
    and g24889 ( n24218 , n24411 , n6957 );
    or g24890 ( n1043 , n10414 , n23193 );
    xnor g24891 ( n24165 , n11948 , n652 );
    nor g24892 ( n24172 , n2033 , n13706 );
    or g24893 ( n14450 , n472 , n26752 );
    xnor g24894 ( n3220 , n5873 , n19001 );
    nor g24895 ( n6288 , n21593 , n20972 );
    or g24896 ( n23699 , n9048 , n14951 );
    and g24897 ( n11546 , n18292 , n2029 );
    nor g24898 ( n2318 , n18004 , n350 );
    and g24899 ( n2834 , n8640 , n13065 );
    not g24900 ( n10541 , n17048 );
    and g24901 ( n9168 , n18523 , n9774 );
    xnor g24902 ( n19352 , n15258 , n4588 );
    not g24903 ( n7341 , n22215 );
    or g24904 ( n19657 , n14507 , n23208 );
    nor g24905 ( n3970 , n9222 , n19143 );
    or g24906 ( n8565 , n12924 , n23597 );
    or g24907 ( n2740 , n9832 , n21240 );
    or g24908 ( n20843 , n24783 , n5199 );
    nor g24909 ( n4833 , n8856 , n8305 );
    and g24910 ( n10063 , n2517 , n9194 );
    not g24911 ( n14346 , n18234 );
    nor g24912 ( n16127 , n8363 , n2816 );
    or g24913 ( n19972 , n23362 , n13196 );
    and g24914 ( n25029 , n16473 , n2111 );
    and g24915 ( n4691 , n2371 , n19255 );
    nor g24916 ( n249 , n10341 , n9855 );
    xnor g24917 ( n25398 , n7546 , n6831 );
    and g24918 ( n21058 , n17609 , n12568 );
    or g24919 ( n15714 , n7090 , n16855 );
    not g24920 ( n9402 , n24692 );
    xnor g24921 ( n19913 , n23591 , n19465 );
    xnor g24922 ( n16340 , n252 , n20316 );
    xnor g24923 ( n24086 , n2146 , n19144 );
    nor g24924 ( n25690 , n19469 , n27188 );
    and g24925 ( n23548 , n1644 , n21612 );
    xnor g24926 ( n25310 , n7973 , n15179 );
    and g24927 ( n13145 , n23522 , n7500 );
    xnor g24928 ( n13695 , n13376 , n4643 );
    not g24929 ( n14783 , n13472 );
    nor g24930 ( n1816 , n17568 , n26986 );
    xnor g24931 ( n650 , n23256 , n23287 );
    xnor g24932 ( n10836 , n9793 , n22361 );
    nor g24933 ( n22460 , n24031 , n21915 );
    and g24934 ( n19269 , n6350 , n27023 );
    xnor g24935 ( n12814 , n17993 , n23145 );
    and g24936 ( n8152 , n21739 , n24805 );
    buf g24937 ( n11669 , n26208 );
    xnor g24938 ( n26853 , n9242 , n17541 );
    xnor g24939 ( n24632 , n8331 , n5743 );
    xnor g24940 ( n26726 , n7815 , n18210 );
    or g24941 ( n2064 , n10211 , n19565 );
    or g24942 ( n18410 , n16755 , n2816 );
    and g24943 ( n5736 , n8948 , n3470 );
    xnor g24944 ( n14648 , n2984 , n25867 );
    not g24945 ( n17581 , n14487 );
    and g24946 ( n20465 , n2796 , n18984 );
    and g24947 ( n13806 , n19373 , n23381 );
    not g24948 ( n19106 , n10611 );
    nor g24949 ( n18394 , n15959 , n10075 );
    and g24950 ( n6540 , n15431 , n21105 );
    or g24951 ( n23169 , n23487 , n12956 );
    and g24952 ( n25834 , n4671 , n7128 );
    xnor g24953 ( n17913 , n13152 , n2688 );
    xnor g24954 ( n10278 , n151 , n21405 );
    nor g24955 ( n13653 , n6351 , n354 );
    nor g24956 ( n11402 , n23160 , n8067 );
    not g24957 ( n15274 , n24473 );
    nor g24958 ( n15684 , n6658 , n6255 );
    xnor g24959 ( n18782 , n1382 , n2356 );
    and g24960 ( n11962 , n19697 , n11890 );
    or g24961 ( n11427 , n7189 , n11255 );
    not g24962 ( n3742 , n21952 );
    xnor g24963 ( n23188 , n11207 , n20986 );
    or g24964 ( n26757 , n7026 , n17835 );
    or g24965 ( n986 , n16045 , n7321 );
    xnor g24966 ( n14600 , n194 , n24696 );
    not g24967 ( n1799 , n21001 );
    and g24968 ( n10675 , n21917 , n16986 );
    xnor g24969 ( n12483 , n14573 , n25381 );
    not g24970 ( n5094 , n474 );
    nor g24971 ( n17528 , n2263 , n13857 );
    xnor g24972 ( n4247 , n3740 , n21784 );
    xnor g24973 ( n9455 , n10868 , n22554 );
    not g24974 ( n2077 , n14954 );
    or g24975 ( n9283 , n14203 , n26554 );
    not g24976 ( n24325 , n16376 );
    not g24977 ( n11259 , n26893 );
    or g24978 ( n23520 , n14525 , n6818 );
    not g24979 ( n6182 , n23357 );
    nor g24980 ( n11978 , n2657 , n13073 );
    or g24981 ( n16773 , n16443 , n23829 );
    nor g24982 ( n8192 , n4040 , n13775 );
    xnor g24983 ( n12552 , n4329 , n8019 );
    xnor g24984 ( n691 , n17936 , n11971 );
    and g24985 ( n5130 , n1681 , n9196 );
    xnor g24986 ( n10388 , n9271 , n21893 );
    not g24987 ( n14699 , n1844 );
    and g24988 ( n11370 , n19094 , n19156 );
    or g24989 ( n11446 , n17479 , n26054 );
    not g24990 ( n21007 , n9185 );
    xnor g24991 ( n7484 , n16037 , n18291 );
    nor g24992 ( n19211 , n22557 , n7447 );
    or g24993 ( n22649 , n19716 , n10269 );
    nor g24994 ( n3206 , n13480 , n22270 );
    xnor g24995 ( n12679 , n10415 , n11299 );
    not g24996 ( n3672 , n933 );
    nor g24997 ( n19986 , n25043 , n25612 );
    or g24998 ( n10646 , n17230 , n658 );
    xnor g24999 ( n6853 , n7248 , n12099 );
    or g25000 ( n14054 , n22990 , n769 );
    or g25001 ( n1284 , n5328 , n20273 );
    and g25002 ( n20548 , n24366 , n14395 );
    xnor g25003 ( n26556 , n6764 , n1451 );
    and g25004 ( n17465 , n1930 , n5681 );
    nor g25005 ( n10421 , n18412 , n1837 );
    nor g25006 ( n17187 , n2935 , n3203 );
    xnor g25007 ( n2010 , n7761 , n22222 );
    nor g25008 ( n10548 , n446 , n3324 );
    or g25009 ( n11093 , n12066 , n7788 );
    nor g25010 ( n6161 , n11198 , n4384 );
    xnor g25011 ( n3662 , n13562 , n15127 );
    and g25012 ( n16220 , n11389 , n9369 );
    buf g25013 ( n6068 , n25607 );
    or g25014 ( n5097 , n4061 , n18473 );
    nor g25015 ( n2202 , n19926 , n1243 );
    and g25016 ( n25349 , n20272 , n20439 );
    xnor g25017 ( n19485 , n1066 , n21565 );
    or g25018 ( n25280 , n4650 , n19008 );
    nor g25019 ( n25409 , n2436 , n15502 );
    or g25020 ( n16250 , n16931 , n26397 );
    xnor g25021 ( n12558 , n20179 , n3460 );
    and g25022 ( n5002 , n23387 , n701 );
    not g25023 ( n2514 , n12811 );
    xnor g25024 ( n18630 , n22919 , n3618 );
    nor g25025 ( n15298 , n15897 , n24217 );
    or g25026 ( n18376 , n7035 , n8529 );
    xnor g25027 ( n25641 , n7400 , n2124 );
    nor g25028 ( n4321 , n17088 , n17832 );
    xnor g25029 ( n3746 , n2162 , n3486 );
    nor g25030 ( n18986 , n18473 , n19514 );
    or g25031 ( n11904 , n13088 , n12720 );
    not g25032 ( n16163 , n3075 );
    and g25033 ( n4845 , n8068 , n4466 );
    xnor g25034 ( n8148 , n16112 , n1034 );
    or g25035 ( n14729 , n2563 , n19381 );
    xnor g25036 ( n18373 , n20289 , n12293 );
    xnor g25037 ( n10874 , n6973 , n21049 );
    not g25038 ( n14318 , n219 );
    not g25039 ( n11685 , n25126 );
    nor g25040 ( n10946 , n10514 , n4514 );
    or g25041 ( n14232 , n7883 , n8402 );
    or g25042 ( n4578 , n16971 , n15600 );
    nor g25043 ( n2821 , n21492 , n7776 );
    nor g25044 ( n22924 , n8002 , n19539 );
    xnor g25045 ( n19177 , n1174 , n1109 );
    or g25046 ( n19934 , n17013 , n18674 );
    or g25047 ( n514 , n5802 , n19368 );
    xnor g25048 ( n14656 , n22342 , n13719 );
    or g25049 ( n21801 , n10406 , n8947 );
    xnor g25050 ( n5802 , n10419 , n765 );
    or g25051 ( n5913 , n16244 , n16264 );
    xnor g25052 ( n19309 , n893 , n13439 );
    or g25053 ( n8110 , n8648 , n13287 );
    or g25054 ( n5540 , n24325 , n6381 );
    xnor g25055 ( n16038 , n7851 , n10045 );
    xnor g25056 ( n15140 , n4294 , n11381 );
    and g25057 ( n9896 , n15003 , n8995 );
    not g25058 ( n18220 , n9259 );
    xnor g25059 ( n13010 , n20826 , n626 );
    or g25060 ( n19473 , n24358 , n1898 );
    or g25061 ( n21439 , n1154 , n20854 );
    or g25062 ( n21553 , n10719 , n19958 );
    not g25063 ( n9505 , n9266 );
    and g25064 ( n8356 , n17682 , n3546 );
    or g25065 ( n17778 , n15062 , n15985 );
    and g25066 ( n22142 , n20974 , n2932 );
    and g25067 ( n19643 , n17304 , n19212 );
    nor g25068 ( n24231 , n16084 , n21691 );
    xnor g25069 ( n1945 , n10201 , n22379 );
    xnor g25070 ( n19641 , n10187 , n17165 );
    or g25071 ( n11475 , n13283 , n24296 );
    or g25072 ( n26710 , n27020 , n1567 );
    or g25073 ( n9536 , n26857 , n13739 );
    not g25074 ( n24695 , n25023 );
    not g25075 ( n10191 , n3832 );
    xnor g25076 ( n16226 , n14996 , n9226 );
    or g25077 ( n13325 , n7769 , n21436 );
    or g25078 ( n9475 , n22333 , n5072 );
    and g25079 ( n10299 , n16269 , n6314 );
    and g25080 ( n15924 , n15944 , n16432 );
    xnor g25081 ( n22494 , n13741 , n15728 );
    or g25082 ( n3539 , n7027 , n24436 );
    and g25083 ( n7521 , n1720 , n6543 );
    xnor g25084 ( n24481 , n11332 , n25423 );
    xnor g25085 ( n12235 , n17869 , n4183 );
    or g25086 ( n6106 , n13400 , n18283 );
    and g25087 ( n16677 , n15778 , n18588 );
    xnor g25088 ( n7834 , n5870 , n6752 );
    or g25089 ( n19099 , n17475 , n23262 );
    xnor g25090 ( n21319 , n8888 , n12871 );
    xnor g25091 ( n3369 , n1753 , n21733 );
    not g25092 ( n25324 , n4326 );
    not g25093 ( n9576 , n4762 );
    or g25094 ( n25997 , n19806 , n5737 );
    and g25095 ( n285 , n9016 , n26842 );
    xnor g25096 ( n5643 , n18568 , n674 );
    and g25097 ( n3631 , n26194 , n12299 );
    xnor g25098 ( n23053 , n3433 , n13993 );
    nor g25099 ( n896 , n17780 , n19377 );
    xnor g25100 ( n11277 , n2371 , n14713 );
    or g25101 ( n13749 , n27199 , n19843 );
    xnor g25102 ( n21682 , n24868 , n23268 );
    not g25103 ( n5366 , n27169 );
    and g25104 ( n23648 , n6353 , n8434 );
    not g25105 ( n3069 , n8006 );
    and g25106 ( n11524 , n14220 , n24678 );
    and g25107 ( n11895 , n420 , n18219 );
    not g25108 ( n2163 , n26425 );
    nor g25109 ( n24077 , n1642 , n18409 );
    or g25110 ( n13275 , n13353 , n18035 );
    xnor g25111 ( n23047 , n3688 , n11206 );
    and g25112 ( n4265 , n13960 , n19785 );
    not g25113 ( n22702 , n20238 );
    and g25114 ( n18451 , n20314 , n13348 );
    xnor g25115 ( n19696 , n8695 , n8492 );
    nor g25116 ( n21994 , n23321 , n6300 );
    and g25117 ( n18985 , n6036 , n20892 );
    xnor g25118 ( n9803 , n21838 , n25489 );
    nor g25119 ( n16308 , n12249 , n13875 );
    nor g25120 ( n19850 , n144 , n25119 );
    and g25121 ( n2643 , n16912 , n7315 );
    xnor g25122 ( n11149 , n10027 , n5822 );
    and g25123 ( n7614 , n21343 , n9710 );
    and g25124 ( n9019 , n15187 , n5995 );
    xnor g25125 ( n21384 , n16524 , n20923 );
    or g25126 ( n20990 , n26822 , n5475 );
    and g25127 ( n21480 , n4030 , n13636 );
    nor g25128 ( n15952 , n20517 , n26239 );
    nor g25129 ( n21022 , n2704 , n7732 );
    nor g25130 ( n14823 , n13291 , n2443 );
    or g25131 ( n6333 , n22660 , n1596 );
    or g25132 ( n17886 , n26296 , n25372 );
    xnor g25133 ( n2023 , n6000 , n24464 );
    xnor g25134 ( n15511 , n22556 , n7069 );
    nor g25135 ( n20496 , n7693 , n22820 );
    or g25136 ( n19598 , n22558 , n6814 );
    or g25137 ( n12107 , n22118 , n7058 );
    xnor g25138 ( n21998 , n17830 , n10739 );
    xnor g25139 ( n15874 , n8052 , n23369 );
    or g25140 ( n12846 , n7893 , n1654 );
    or g25141 ( n18579 , n18896 , n3101 );
    and g25142 ( n2406 , n12031 , n14752 );
    or g25143 ( n3695 , n15507 , n19785 );
    xnor g25144 ( n11800 , n26947 , n12612 );
    or g25145 ( n6858 , n18361 , n12439 );
    or g25146 ( n9892 , n5356 , n5639 );
    xnor g25147 ( n4322 , n21928 , n11223 );
    or g25148 ( n1041 , n1090 , n12687 );
    and g25149 ( n3961 , n4041 , n3378 );
    or g25150 ( n9530 , n17185 , n12747 );
    nor g25151 ( n20472 , n23034 , n21352 );
    and g25152 ( n9553 , n2567 , n4525 );
    xnor g25153 ( n17207 , n15242 , n11669 );
    or g25154 ( n6688 , n25558 , n13748 );
    nor g25155 ( n5406 , n6337 , n3686 );
    xnor g25156 ( n535 , n22114 , n268 );
    nor g25157 ( n2403 , n21846 , n9493 );
    or g25158 ( n8551 , n6528 , n16194 );
    xnor g25159 ( n6652 , n26254 , n8826 );
    and g25160 ( n2143 , n315 , n25804 );
    not g25161 ( n25139 , n11615 );
    nor g25162 ( n26971 , n8272 , n17888 );
    xnor g25163 ( n1924 , n19418 , n3901 );
    or g25164 ( n24693 , n3260 , n21832 );
    xnor g25165 ( n18486 , n9294 , n26022 );
    or g25166 ( n10567 , n26661 , n8596 );
    xnor g25167 ( n23783 , n4302 , n3872 );
    xnor g25168 ( n2050 , n10097 , n8935 );
    and g25169 ( n22066 , n9563 , n9903 );
    and g25170 ( n1068 , n4188 , n12922 );
    not g25171 ( n2017 , n9872 );
    and g25172 ( n23776 , n17097 , n24909 );
    and g25173 ( n21562 , n22442 , n25038 );
    xnor g25174 ( n14713 , n18093 , n25427 );
    or g25175 ( n23444 , n3069 , n5211 );
    or g25176 ( n12139 , n15076 , n13620 );
    xnor g25177 ( n23743 , n26028 , n17867 );
    and g25178 ( n44 , n22115 , n22163 );
    xnor g25179 ( n12146 , n10299 , n24353 );
    xnor g25180 ( n21237 , n14749 , n856 );
    not g25181 ( n23466 , n21782 );
    not g25182 ( n12207 , n2226 );
    buf g25183 ( n10505 , n17653 );
    not g25184 ( n17369 , n4909 );
    and g25185 ( n10609 , n20758 , n5308 );
    and g25186 ( n24697 , n15341 , n226 );
    not g25187 ( n182 , n6445 );
    nor g25188 ( n15830 , n27167 , n14804 );
    not g25189 ( n17390 , n25113 );
    nor g25190 ( n23055 , n19588 , n8322 );
    nor g25191 ( n3410 , n17316 , n14750 );
    not g25192 ( n3178 , n21898 );
    or g25193 ( n594 , n1806 , n22185 );
    and g25194 ( n18910 , n20712 , n12896 );
    and g25195 ( n16224 , n22184 , n5962 );
    or g25196 ( n17534 , n20929 , n23068 );
    xnor g25197 ( n18215 , n12657 , n21287 );
    not g25198 ( n14002 , n22871 );
    and g25199 ( n2810 , n7839 , n23363 );
    or g25200 ( n1989 , n12871 , n8888 );
    or g25201 ( n3720 , n6501 , n14941 );
    xnor g25202 ( n12131 , n2683 , n19071 );
    and g25203 ( n430 , n4369 , n4336 );
    xnor g25204 ( n1823 , n16701 , n25144 );
    not g25205 ( n26078 , n12860 );
    and g25206 ( n16537 , n2117 , n6711 );
    or g25207 ( n19528 , n20717 , n482 );
    xnor g25208 ( n91 , n25556 , n5328 );
    nor g25209 ( n20588 , n10077 , n9285 );
    not g25210 ( n26544 , n16724 );
    nor g25211 ( n15712 , n4042 , n10833 );
    and g25212 ( n17135 , n17839 , n2294 );
    xnor g25213 ( n1854 , n25953 , n12868 );
    or g25214 ( n23437 , n7143 , n10728 );
    xnor g25215 ( n4189 , n23704 , n20359 );
    or g25216 ( n25357 , n16742 , n12285 );
    xnor g25217 ( n8974 , n10157 , n22753 );
    xnor g25218 ( n6373 , n15988 , n5343 );
    or g25219 ( n8014 , n8087 , n15643 );
    or g25220 ( n22553 , n3046 , n19655 );
    xnor g25221 ( n16457 , n10096 , n26553 );
    or g25222 ( n6077 , n3384 , n6244 );
    or g25223 ( n10636 , n17122 , n26177 );
    xnor g25224 ( n10631 , n22037 , n20669 );
    and g25225 ( n13599 , n9533 , n23794 );
    xnor g25226 ( n8146 , n25374 , n6532 );
    xnor g25227 ( n2418 , n12185 , n1301 );
    nor g25228 ( n24864 , n399 , n13949 );
    or g25229 ( n24362 , n18217 , n12718 );
    nor g25230 ( n22577 , n7676 , n12512 );
    and g25231 ( n18465 , n20532 , n7416 );
    or g25232 ( n26756 , n11278 , n2815 );
    or g25233 ( n14581 , n6156 , n19859 );
    or g25234 ( n19197 , n776 , n21430 );
    xnor g25235 ( n17733 , n350 , n1882 );
    or g25236 ( n24773 , n10119 , n2526 );
    or g25237 ( n18140 , n9679 , n22626 );
    or g25238 ( n16763 , n25760 , n18330 );
    xnor g25239 ( n26667 , n20855 , n5827 );
    xnor g25240 ( n23170 , n3888 , n2993 );
    or g25241 ( n25143 , n4713 , n14067 );
    or g25242 ( n19999 , n25772 , n22047 );
    or g25243 ( n559 , n12160 , n10562 );
    and g25244 ( n13840 , n12482 , n19441 );
    xnor g25245 ( n16304 , n17382 , n5207 );
    not g25246 ( n277 , n10001 );
    not g25247 ( n5728 , n23372 );
    or g25248 ( n7016 , n11896 , n9384 );
    xnor g25249 ( n6863 , n4304 , n1563 );
    or g25250 ( n13440 , n14437 , n16663 );
    not g25251 ( n21694 , n1185 );
    or g25252 ( n18825 , n24051 , n15996 );
    or g25253 ( n1897 , n5641 , n1430 );
    xnor g25254 ( n12850 , n16325 , n9832 );
    or g25255 ( n25472 , n543 , n2244 );
    xnor g25256 ( n22004 , n8933 , n6865 );
    or g25257 ( n20320 , n7380 , n3226 );
    not g25258 ( n15113 , n14156 );
    and g25259 ( n11437 , n8436 , n16076 );
    or g25260 ( n16622 , n16294 , n17568 );
    not g25261 ( n6917 , n22993 );
    xnor g25262 ( n7555 , n8902 , n5902 );
    xnor g25263 ( n17183 , n6440 , n23420 );
    nor g25264 ( n9162 , n10956 , n1598 );
    xnor g25265 ( n1339 , n12935 , n22162 );
    or g25266 ( n738 , n7320 , n6381 );
    or g25267 ( n2789 , n18280 , n5937 );
    and g25268 ( n23265 , n26852 , n13213 );
    xnor g25269 ( n2002 , n1339 , n14633 );
    xnor g25270 ( n14126 , n10750 , n2086 );
    or g25271 ( n4363 , n20667 , n12956 );
    and g25272 ( n3230 , n19127 , n18200 );
    nor g25273 ( n23073 , n8084 , n18755 );
    or g25274 ( n27137 , n14422 , n16113 );
    xnor g25275 ( n19951 , n12745 , n22542 );
    or g25276 ( n1063 , n20544 , n23586 );
    or g25277 ( n1711 , n19606 , n14578 );
    and g25278 ( n746 , n10470 , n4062 );
    not g25279 ( n23059 , n8403 );
    or g25280 ( n17991 , n10248 , n10358 );
    or g25281 ( n14417 , n24611 , n6578 );
    xnor g25282 ( n16091 , n10765 , n2337 );
    not g25283 ( n12301 , n17968 );
    and g25284 ( n15938 , n23144 , n10306 );
    or g25285 ( n591 , n12320 , n194 );
    nor g25286 ( n1868 , n24327 , n4325 );
    xnor g25287 ( n12665 , n27069 , n4937 );
    xnor g25288 ( n15379 , n5226 , n11223 );
    or g25289 ( n14556 , n12160 , n16994 );
    and g25290 ( n20682 , n15425 , n19870 );
    xnor g25291 ( n3270 , n24620 , n21753 );
    xnor g25292 ( n15573 , n9862 , n19308 );
    buf g25293 ( n17549 , n7856 );
    xnor g25294 ( n16907 , n9390 , n11730 );
    xnor g25295 ( n1991 , n11163 , n19642 );
    or g25296 ( n2188 , n9118 , n13661 );
    xnor g25297 ( n26419 , n16009 , n12910 );
    not g25298 ( n3921 , n152 );
    or g25299 ( n20914 , n16084 , n18537 );
    xnor g25300 ( n22888 , n23517 , n10369 );
    and g25301 ( n22952 , n5622 , n12077 );
    xnor g25302 ( n25687 , n11454 , n19364 );
    or g25303 ( n8136 , n15144 , n25359 );
    or g25304 ( n17919 , n13109 , n24898 );
    and g25305 ( n25438 , n3655 , n17924 );
    xnor g25306 ( n7793 , n26107 , n4376 );
    xnor g25307 ( n22105 , n12684 , n21683 );
    and g25308 ( n15072 , n26925 , n9394 );
    xnor g25309 ( n873 , n22647 , n6402 );
    not g25310 ( n6595 , n24949 );
    not g25311 ( n12639 , n2272 );
    and g25312 ( n10576 , n4338 , n24430 );
    xnor g25313 ( n5184 , n4754 , n13648 );
    and g25314 ( n4111 , n16999 , n7370 );
    xnor g25315 ( n13684 , n24320 , n8256 );
    or g25316 ( n2934 , n8802 , n16191 );
    and g25317 ( n10503 , n11742 , n19600 );
    xnor g25318 ( n24726 , n17371 , n15506 );
    or g25319 ( n20565 , n23144 , n22125 );
    and g25320 ( n22431 , n7675 , n26182 );
    xnor g25321 ( n9938 , n21183 , n23364 );
    and g25322 ( n14792 , n1076 , n5678 );
    and g25323 ( n17042 , n33 , n999 );
    and g25324 ( n4028 , n7923 , n11458 );
    or g25325 ( n14726 , n5714 , n12531 );
    or g25326 ( n14266 , n11026 , n13441 );
    nor g25327 ( n25589 , n14719 , n1421 );
    xnor g25328 ( n24796 , n14674 , n10733 );
    or g25329 ( n12124 , n24480 , n16627 );
    or g25330 ( n20810 , n26462 , n2208 );
    xnor g25331 ( n17569 , n19805 , n11192 );
    not g25332 ( n21556 , n7099 );
    not g25333 ( n4642 , n19161 );
    xnor g25334 ( n9986 , n12336 , n11752 );
    nor g25335 ( n21978 , n16665 , n19803 );
    not g25336 ( n15693 , n9850 );
    nor g25337 ( n19006 , n18105 , n21392 );
    xnor g25338 ( n6422 , n19048 , n16955 );
    xnor g25339 ( n317 , n24912 , n8490 );
    or g25340 ( n444 , n26264 , n12911 );
    or g25341 ( n26676 , n13013 , n14591 );
    xnor g25342 ( n10938 , n13224 , n11273 );
    not g25343 ( n22281 , n21276 );
    not g25344 ( n13495 , n13036 );
    and g25345 ( n12981 , n24328 , n13616 );
    xnor g25346 ( n8219 , n456 , n15400 );
    or g25347 ( n23051 , n7462 , n6524 );
    nor g25348 ( n305 , n18737 , n15268 );
    nor g25349 ( n15984 , n22425 , n14984 );
    nor g25350 ( n11291 , n8138 , n21656 );
    xnor g25351 ( n18037 , n19387 , n14229 );
    xnor g25352 ( n6807 , n26536 , n19607 );
    xnor g25353 ( n11973 , n5207 , n21284 );
    or g25354 ( n3805 , n16878 , n17883 );
    xnor g25355 ( n11893 , n14308 , n25979 );
    xnor g25356 ( n15175 , n26791 , n2457 );
    and g25357 ( n14347 , n2120 , n877 );
    nor g25358 ( n24877 , n537 , n8456 );
    or g25359 ( n6191 , n12237 , n6639 );
    and g25360 ( n6000 , n16598 , n2373 );
    xnor g25361 ( n17730 , n21941 , n4325 );
    or g25362 ( n15214 , n10918 , n12105 );
    and g25363 ( n21482 , n25717 , n26608 );
    nor g25364 ( n22595 , n25475 , n17716 );
    and g25365 ( n11072 , n15442 , n17382 );
    and g25366 ( n19666 , n8671 , n17181 );
    xnor g25367 ( n25934 , n13541 , n12832 );
    or g25368 ( n22479 , n21420 , n26573 );
    and g25369 ( n19794 , n3909 , n13591 );
    or g25370 ( n18969 , n20056 , n13356 );
    nor g25371 ( n22238 , n14440 , n21287 );
    or g25372 ( n18641 , n9177 , n18233 );
    or g25373 ( n18374 , n1105 , n21175 );
    or g25374 ( n13330 , n5480 , n1067 );
    and g25375 ( n19739 , n17280 , n8312 );
    not g25376 ( n7396 , n10529 );
    or g25377 ( n4351 , n7341 , n2954 );
    or g25378 ( n10789 , n6924 , n18283 );
    xnor g25379 ( n23355 , n8107 , n19891 );
    xnor g25380 ( n6323 , n261 , n12538 );
    not g25381 ( n286 , n15360 );
    not g25382 ( n8032 , n26748 );
    xnor g25383 ( n1398 , n14148 , n1152 );
    and g25384 ( n11721 , n5799 , n20067 );
    nor g25385 ( n9065 , n2514 , n19514 );
    or g25386 ( n25990 , n644 , n154 );
    xnor g25387 ( n7871 , n16852 , n9967 );
    xnor g25388 ( n14454 , n14777 , n3236 );
    and g25389 ( n19374 , n8337 , n2493 );
    xnor g25390 ( n1005 , n23847 , n2630 );
    not g25391 ( n25610 , n8088 );
    and g25392 ( n12127 , n6113 , n18733 );
    and g25393 ( n23469 , n6691 , n19222 );
    xnor g25394 ( n22361 , n19937 , n20162 );
    or g25395 ( n19699 , n9502 , n1066 );
    xnor g25396 ( n6343 , n24805 , n11321 );
    xnor g25397 ( n6082 , n6762 , n2289 );
    or g25398 ( n20614 , n16937 , n19005 );
    and g25399 ( n17591 , n18812 , n22408 );
    not g25400 ( n22034 , n16582 );
    and g25401 ( n19638 , n11562 , n2635 );
    and g25402 ( n20902 , n9246 , n12955 );
    or g25403 ( n5398 , n22468 , n5679 );
    and g25404 ( n14082 , n11269 , n17025 );
    xnor g25405 ( n5161 , n21772 , n626 );
    xnor g25406 ( n26801 , n2824 , n13827 );
    or g25407 ( n16556 , n2269 , n21689 );
    not g25408 ( n4508 , n10750 );
    xnor g25409 ( n7887 , n25345 , n25475 );
    and g25410 ( n23526 , n18345 , n20964 );
    and g25411 ( n768 , n19279 , n6041 );
    and g25412 ( n14491 , n9154 , n3658 );
    or g25413 ( n10930 , n9095 , n7913 );
    or g25414 ( n2419 , n13992 , n11722 );
    or g25415 ( n17394 , n2915 , n10625 );
    not g25416 ( n42 , n10746 );
    not g25417 ( n5974 , n20933 );
    not g25418 ( n1349 , n27055 );
    xnor g25419 ( n9057 , n3582 , n21784 );
    not g25420 ( n22666 , n4108 );
    xnor g25421 ( n4801 , n21027 , n13555 );
    and g25422 ( n1006 , n2483 , n6079 );
    xnor g25423 ( n8250 , n23191 , n25288 );
    and g25424 ( n13904 , n11490 , n6856 );
    and g25425 ( n16329 , n14490 , n2803 );
    and g25426 ( n1002 , n9380 , n7676 );
    nor g25427 ( n16453 , n17171 , n182 );
    or g25428 ( n16710 , n5684 , n8558 );
    nor g25429 ( n4579 , n10593 , n8657 );
    not g25430 ( n23217 , n15064 );
    xnor g25431 ( n22157 , n13862 , n4015 );
    nor g25432 ( n24631 , n6731 , n5066 );
    xnor g25433 ( n24596 , n8302 , n14545 );
    and g25434 ( n23930 , n25371 , n17565 );
    and g25435 ( n7854 , n18871 , n21614 );
    or g25436 ( n14558 , n6398 , n5251 );
    xnor g25437 ( n8195 , n22615 , n14015 );
    xnor g25438 ( n3405 , n25361 , n5187 );
    or g25439 ( n6537 , n2391 , n19886 );
    or g25440 ( n13302 , n2967 , n20179 );
    and g25441 ( n6645 , n6299 , n14341 );
    nor g25442 ( n24387 , n19081 , n21400 );
    nor g25443 ( n22817 , n7917 , n8391 );
    not g25444 ( n11217 , n12668 );
    xnor g25445 ( n22058 , n17938 , n21455 );
    xnor g25446 ( n22620 , n4842 , n24634 );
    xnor g25447 ( n18719 , n17692 , n4877 );
    and g25448 ( n7340 , n12600 , n3210 );
    xnor g25449 ( n20618 , n2167 , n17733 );
    not g25450 ( n13191 , n25185 );
    and g25451 ( n20426 , n5447 , n26811 );
    or g25452 ( n3201 , n7898 , n27103 );
    and g25453 ( n8865 , n13708 , n13842 );
    not g25454 ( n20751 , n14153 );
    and g25455 ( n8527 , n22707 , n7852 );
    or g25456 ( n6211 , n13887 , n7786 );
    and g25457 ( n18211 , n17031 , n11868 );
    nor g25458 ( n24252 , n12762 , n25533 );
    xnor g25459 ( n5707 , n376 , n7721 );
    xnor g25460 ( n26511 , n14003 , n10920 );
    or g25461 ( n14220 , n23153 , n16523 );
    or g25462 ( n21638 , n8082 , n24864 );
    xnor g25463 ( n19988 , n9478 , n10032 );
    or g25464 ( n10857 , n8055 , n12527 );
    xnor g25465 ( n14900 , n19521 , n3719 );
    and g25466 ( n12646 , n22811 , n15485 );
    and g25467 ( n10179 , n7682 , n733 );
    or g25468 ( n16016 , n17869 , n24664 );
    and g25469 ( n14105 , n13608 , n3768 );
    not g25470 ( n13073 , n22548 );
    or g25471 ( n14586 , n6498 , n5319 );
    and g25472 ( n11651 , n6307 , n477 );
    or g25473 ( n21025 , n19905 , n21501 );
    or g25474 ( n24038 , n776 , n8186 );
    or g25475 ( n23334 , n17856 , n21280 );
    or g25476 ( n18709 , n12554 , n18295 );
    nor g25477 ( n23056 , n6178 , n18715 );
    not g25478 ( n25505 , n7435 );
    not g25479 ( n9202 , n26075 );
    and g25480 ( n11286 , n25591 , n23759 );
    not g25481 ( n25502 , n10267 );
    xnor g25482 ( n7650 , n18444 , n26224 );
    not g25483 ( n13633 , n5139 );
    xnor g25484 ( n3800 , n14111 , n14114 );
    and g25485 ( n10309 , n9939 , n6899 );
    nor g25486 ( n8099 , n7143 , n3625 );
    and g25487 ( n20362 , n5673 , n16146 );
    and g25488 ( n2757 , n15350 , n22451 );
    nor g25489 ( n7586 , n3480 , n19911 );
    and g25490 ( n23394 , n21650 , n7411 );
    and g25491 ( n11572 , n12858 , n1436 );
    xnor g25492 ( n16492 , n21674 , n9172 );
    xnor g25493 ( n8985 , n15182 , n21915 );
    not g25494 ( n688 , n6204 );
    xnor g25495 ( n3067 , n5497 , n15226 );
    and g25496 ( n9786 , n19771 , n3910 );
    xnor g25497 ( n25032 , n19605 , n16448 );
    xnor g25498 ( n23578 , n15511 , n19192 );
    or g25499 ( n3286 , n14288 , n6900 );
    nor g25500 ( n4039 , n15967 , n1396 );
    nor g25501 ( n18508 , n20715 , n25065 );
    or g25502 ( n22923 , n1709 , n24961 );
    or g25503 ( n10320 , n10038 , n23409 );
    or g25504 ( n21478 , n9049 , n18524 );
    and g25505 ( n14715 , n25335 , n20041 );
    xnor g25506 ( n20248 , n5400 , n21997 );
    nor g25507 ( n7898 , n8509 , n4315 );
    not g25508 ( n19907 , n19924 );
    or g25509 ( n20648 , n22961 , n8342 );
    nor g25510 ( n8122 , n8495 , n1386 );
    or g25511 ( n21201 , n9603 , n10728 );
    or g25512 ( n19832 , n3228 , n22470 );
    or g25513 ( n17828 , n26725 , n17212 );
    not g25514 ( n7324 , n3834 );
    nor g25515 ( n9264 , n17143 , n3007 );
    nor g25516 ( n17471 , n25345 , n9967 );
    xnor g25517 ( n5722 , n16410 , n13652 );
    xnor g25518 ( n448 , n13112 , n7707 );
    nor g25519 ( n17596 , n22724 , n10001 );
    xnor g25520 ( n6752 , n25700 , n7281 );
    nor g25521 ( n17945 , n2723 , n15650 );
    xnor g25522 ( n22993 , n25598 , n22503 );
    xnor g25523 ( n18802 , n3382 , n1668 );
    or g25524 ( n8175 , n7940 , n6309 );
    and g25525 ( n14758 , n5613 , n25193 );
    xnor g25526 ( n19202 , n24329 , n12683 );
    xnor g25527 ( n16667 , n20968 , n24768 );
    and g25528 ( n11609 , n13749 , n15741 );
    and g25529 ( n19565 , n18366 , n25580 );
    xnor g25530 ( n1992 , n20429 , n26054 );
    xnor g25531 ( n13338 , n23730 , n24900 );
    nor g25532 ( n22403 , n26162 , n8806 );
    xnor g25533 ( n4723 , n21633 , n24376 );
    xnor g25534 ( n11744 , n3474 , n12075 );
    xnor g25535 ( n23310 , n13315 , n5503 );
    or g25536 ( n10901 , n12849 , n25755 );
    and g25537 ( n13819 , n20035 , n12559 );
    not g25538 ( n3238 , n20792 );
    or g25539 ( n25600 , n26252 , n16765 );
    not g25540 ( n6251 , n19270 );
    and g25541 ( n10616 , n5566 , n26676 );
    or g25542 ( n4620 , n21644 , n20562 );
    and g25543 ( n670 , n5906 , n21851 );
    or g25544 ( n13866 , n7980 , n3065 );
    nor g25545 ( n1180 , n8101 , n17250 );
    not g25546 ( n19976 , n12395 );
    or g25547 ( n291 , n2222 , n8567 );
    nor g25548 ( n5931 , n2498 , n14185 );
    and g25549 ( n23298 , n4764 , n6043 );
    not g25550 ( n24825 , n13110 );
    or g25551 ( n9400 , n21267 , n16874 );
    or g25552 ( n26588 , n7452 , n21 );
    and g25553 ( n11289 , n7700 , n13758 );
    xnor g25554 ( n26874 , n19215 , n8875 );
    and g25555 ( n10419 , n18397 , n7720 );
    and g25556 ( n21742 , n12164 , n4817 );
    xnor g25557 ( n10360 , n27114 , n17727 );
    nor g25558 ( n11581 , n26951 , n22477 );
    and g25559 ( n25297 , n26632 , n17049 );
    xnor g25560 ( n13607 , n17803 , n10201 );
    nor g25561 ( n7987 , n22764 , n1536 );
    and g25562 ( n24903 , n23089 , n12877 );
    not g25563 ( n27151 , n25971 );
    and g25564 ( n11937 , n15110 , n16701 );
    or g25565 ( n7129 , n17846 , n12488 );
    or g25566 ( n21578 , n11045 , n25122 );
    and g25567 ( n23406 , n22604 , n2093 );
    not g25568 ( n10324 , n18444 );
    and g25569 ( n2649 , n16835 , n18757 );
    and g25570 ( n11878 , n26473 , n16478 );
    and g25571 ( n1853 , n19966 , n17281 );
    xnor g25572 ( n20017 , n6505 , n6249 );
    nor g25573 ( n25973 , n15506 , n3246 );
    xnor g25574 ( n27095 , n10922 , n16870 );
    xnor g25575 ( n8497 , n2588 , n1654 );
    or g25576 ( n11519 , n11393 , n3480 );
    nor g25577 ( n11560 , n6478 , n17590 );
    or g25578 ( n7760 , n26731 , n17764 );
    xnor g25579 ( n26311 , n8551 , n17071 );
    xnor g25580 ( n10130 , n10885 , n26725 );
    or g25581 ( n22608 , n26374 , n14028 );
    xnor g25582 ( n17976 , n17606 , n9590 );
    xnor g25583 ( n14206 , n26629 , n22266 );
    or g25584 ( n23716 , n19566 , n10300 );
    and g25585 ( n16202 , n26898 , n1149 );
    and g25586 ( n8342 , n12833 , n21009 );
    or g25587 ( n25397 , n343 , n22302 );
    not g25588 ( n15647 , n16167 );
    and g25589 ( n8893 , n14019 , n651 );
    xnor g25590 ( n14976 , n1584 , n17690 );
    or g25591 ( n20453 , n16711 , n12464 );
    nor g25592 ( n21823 , n2446 , n2439 );
    or g25593 ( n2770 , n3480 , n7373 );
    xnor g25594 ( n23212 , n3618 , n8581 );
    xnor g25595 ( n11419 , n25109 , n24514 );
    or g25596 ( n10539 , n1322 , n17194 );
    nor g25597 ( n7664 , n25490 , n12868 );
    and g25598 ( n2334 , n14790 , n5105 );
    or g25599 ( n4041 , n3652 , n22210 );
    or g25600 ( n9903 , n15452 , n22022 );
    nor g25601 ( n20222 , n18651 , n5855 );
    and g25602 ( n244 , n5347 , n14663 );
    xnor g25603 ( n19291 , n3506 , n2743 );
    xor g25604 ( n5187 , n19875 , n7057 );
    xnor g25605 ( n13015 , n27102 , n21078 );
    xnor g25606 ( n20218 , n20925 , n17311 );
    or g25607 ( n2506 , n23097 , n11365 );
    or g25608 ( n15886 , n1401 , n22478 );
    not g25609 ( n420 , n5330 );
    xnor g25610 ( n17857 , n11835 , n20044 );
    or g25611 ( n26075 , n10096 , n22345 );
    or g25612 ( n7070 , n11004 , n18081 );
    or g25613 ( n7594 , n967 , n23511 );
    and g25614 ( n473 , n22605 , n21648 );
    xnor g25615 ( n14965 , n13942 , n10222 );
    and g25616 ( n19629 , n4567 , n19723 );
    xnor g25617 ( n15556 , n19265 , n268 );
    xnor g25618 ( n18843 , n9181 , n6928 );
    and g25619 ( n19059 , n13863 , n5133 );
    nor g25620 ( n15209 , n10156 , n20551 );
    and g25621 ( n536 , n9003 , n23436 );
    not g25622 ( n21085 , n21459 );
    not g25623 ( n3577 , n8070 );
    or g25624 ( n8108 , n11544 , n26986 );
    not g25625 ( n9294 , n13494 );
    xnor g25626 ( n14769 , n15636 , n16223 );
    or g25627 ( n12676 , n16256 , n12079 );
    not g25628 ( n20064 , n14702 );
    nor g25629 ( n14508 , n9093 , n17599 );
    not g25630 ( n24025 , n23504 );
    not g25631 ( n11764 , n2429 );
    not g25632 ( n23095 , n7751 );
    xnor g25633 ( n13478 , n14830 , n6468 );
    or g25634 ( n19441 , n12067 , n6067 );
    nor g25635 ( n8625 , n4613 , n6561 );
    or g25636 ( n23214 , n14707 , n6049 );
    or g25637 ( n799 , n18872 , n5254 );
    or g25638 ( n1842 , n11653 , n14926 );
    xnor g25639 ( n789 , n3196 , n2046 );
    xnor g25640 ( n22027 , n10238 , n3300 );
    xnor g25641 ( n11701 , n12142 , n6787 );
    nor g25642 ( n17137 , n1642 , n10158 );
    xnor g25643 ( n9783 , n25456 , n4408 );
    and g25644 ( n18049 , n20305 , n2179 );
    or g25645 ( n14529 , n11159 , n10186 );
    nor g25646 ( n19763 , n23966 , n13925 );
    and g25647 ( n25698 , n26892 , n11623 );
    and g25648 ( n9466 , n4514 , n5111 );
    or g25649 ( n25169 , n13033 , n18907 );
    nor g25650 ( n3329 , n2342 , n23430 );
    not g25651 ( n13497 , n2117 );
    and g25652 ( n19591 , n1663 , n3777 );
    nor g25653 ( n18413 , n7237 , n25120 );
    or g25654 ( n5347 , n1994 , n19556 );
    and g25655 ( n25125 , n5589 , n7934 );
    and g25656 ( n8134 , n14936 , n20423 );
    xnor g25657 ( n18826 , n20763 , n12013 );
    and g25658 ( n18217 , n10335 , n10141 );
    and g25659 ( n19505 , n11059 , n23948 );
    or g25660 ( n9704 , n19461 , n6440 );
    or g25661 ( n19687 , n13870 , n13029 );
    and g25662 ( n6524 , n1157 , n20765 );
    not g25663 ( n21151 , n19394 );
    nor g25664 ( n10252 , n20462 , n7086 );
    xnor g25665 ( n26205 , n10335 , n9954 );
    or g25666 ( n1644 , n16252 , n23166 );
    or g25667 ( n3530 , n6927 , n5344 );
    xnor g25668 ( n10745 , n8614 , n12702 );
    xnor g25669 ( n13072 , n15497 , n26509 );
    or g25670 ( n114 , n9325 , n17633 );
    or g25671 ( n8181 , n19236 , n4275 );
    or g25672 ( n23739 , n8068 , n25316 );
    or g25673 ( n2830 , n12447 , n23599 );
    xnor g25674 ( n6189 , n14938 , n22497 );
    or g25675 ( n770 , n13809 , n4512 );
    and g25676 ( n23870 , n8158 , n2475 );
    nor g25677 ( n12435 , n7882 , n24727 );
    xnor g25678 ( n4115 , n1173 , n583 );
    xnor g25679 ( n3902 , n7910 , n8309 );
    xnor g25680 ( n15304 , n23068 , n20179 );
    or g25681 ( n478 , n8853 , n17652 );
    or g25682 ( n11902 , n6379 , n3040 );
    or g25683 ( n1342 , n25743 , n17751 );
    not g25684 ( n9678 , n25426 );
    xnor g25685 ( n1111 , n8912 , n9474 );
    xnor g25686 ( n10838 , n7305 , n1204 );
    nor g25687 ( n13802 , n26807 , n9273 );
    or g25688 ( n19007 , n21424 , n1318 );
    and g25689 ( n22464 , n7549 , n15247 );
    or g25690 ( n7728 , n12420 , n24143 );
    xnor g25691 ( n12674 , n6810 , n9375 );
    buf g25692 ( n10964 , n7276 );
    and g25693 ( n3328 , n5033 , n3177 );
    xnor g25694 ( n11300 , n19836 , n27121 );
    nor g25695 ( n24264 , n20542 , n25937 );
    xnor g25696 ( n23216 , n518 , n18619 );
    xnor g25697 ( n12158 , n4262 , n20786 );
    or g25698 ( n5589 , n13154 , n4426 );
    or g25699 ( n221 , n12871 , n20411 );
    and g25700 ( n23457 , n11144 , n25500 );
    or g25701 ( n17565 , n26166 , n2106 );
    xnor g25702 ( n4441 , n6793 , n18459 );
    nor g25703 ( n7487 , n14486 , n18031 );
    not g25704 ( n11483 , n18438 );
    and g25705 ( n13446 , n24226 , n3112 );
    xnor g25706 ( n7420 , n676 , n3981 );
    and g25707 ( n15161 , n24869 , n1392 );
    nor g25708 ( n6778 , n22170 , n5098 );
    not g25709 ( n856 , n6129 );
    or g25710 ( n21531 , n26227 , n21284 );
    not g25711 ( n13651 , n18927 );
    xnor g25712 ( n4088 , n11065 , n13869 );
    or g25713 ( n3437 , n24453 , n23844 );
    not g25714 ( n12371 , n11209 );
    or g25715 ( n26787 , n22591 , n24756 );
    xnor g25716 ( n11717 , n21140 , n10241 );
    and g25717 ( n25791 , n19941 , n9345 );
    xnor g25718 ( n10165 , n17825 , n20574 );
    and g25719 ( n1194 , n5881 , n4206 );
    or g25720 ( n3146 , n18892 , n25482 );
    xnor g25721 ( n9691 , n18742 , n20409 );
    or g25722 ( n17274 , n9383 , n21283 );
    xnor g25723 ( n13222 , n25915 , n8024 );
    nor g25724 ( n26828 , n11615 , n8052 );
    or g25725 ( n20831 , n18103 , n5182 );
    nor g25726 ( n23656 , n11829 , n12935 );
    or g25727 ( n18956 , n6623 , n2837 );
    or g25728 ( n1506 , n9040 , n26799 );
    not g25729 ( n22422 , n4856 );
    xnor g25730 ( n14583 , n15967 , n2783 );
    nor g25731 ( n25962 , n12956 , n26913 );
    and g25732 ( n26153 , n2895 , n16972 );
    not g25733 ( n8689 , n10183 );
    nor g25734 ( n7870 , n19905 , n14733 );
    not g25735 ( n13528 , n17452 );
    not g25736 ( n14736 , n19472 );
    not g25737 ( n19427 , n17739 );
    or g25738 ( n6981 , n20338 , n20477 );
    and g25739 ( n373 , n16438 , n2569 );
    or g25740 ( n10133 , n13715 , n10634 );
    and g25741 ( n12564 , n7114 , n9746 );
    and g25742 ( n9720 , n26802 , n18110 );
    xnor g25743 ( n25947 , n17987 , n15683 );
    xnor g25744 ( n21879 , n23291 , n14201 );
    or g25745 ( n13644 , n688 , n3795 );
    or g25746 ( n1908 , n26482 , n26089 );
    xnor g25747 ( n15255 , n12573 , n5614 );
    and g25748 ( n20900 , n6198 , n9544 );
    or g25749 ( n20855 , n8191 , n12645 );
    xnor g25750 ( n21909 , n21205 , n5226 );
    or g25751 ( n7562 , n20400 , n13520 );
    and g25752 ( n21689 , n17459 , n5216 );
    not g25753 ( n11113 , n17233 );
    xnor g25754 ( n10493 , n17134 , n21573 );
    and g25755 ( n12681 , n7255 , n22598 );
    xnor g25756 ( n1709 , n8951 , n9775 );
    and g25757 ( n26147 , n17513 , n26490 );
    not g25758 ( n22723 , n13668 );
    xnor g25759 ( n8233 , n13164 , n12060 );
    xnor g25760 ( n5803 , n22442 , n22253 );
    not g25761 ( n24686 , n11458 );
    and g25762 ( n17033 , n1743 , n25598 );
    xnor g25763 ( n6328 , n16283 , n17037 );
    xnor g25764 ( n19141 , n18393 , n5336 );
    not g25765 ( n11111 , n7234 );
    xnor g25766 ( n24964 , n14761 , n6218 );
    xnor g25767 ( n7345 , n24599 , n9398 );
    or g25768 ( n24454 , n4500 , n855 );
    xnor g25769 ( n25891 , n2463 , n5677 );
    not g25770 ( n13405 , n8305 );
    or g25771 ( n18642 , n25038 , n16544 );
    xnor g25772 ( n11987 , n10749 , n21487 );
    and g25773 ( n5520 , n7960 , n7015 );
    and g25774 ( n14590 , n26366 , n17080 );
    and g25775 ( n19410 , n6659 , n20384 );
    xnor g25776 ( n20935 , n13057 , n17032 );
    or g25777 ( n8583 , n14440 , n3504 );
    xnor g25778 ( n10260 , n22755 , n7503 );
    nor g25779 ( n782 , n26437 , n25415 );
    not g25780 ( n14185 , n26058 );
    or g25781 ( n8404 , n7880 , n3389 );
    xnor g25782 ( n22586 , n19701 , n13074 );
    or g25783 ( n18096 , n4468 , n2780 );
    or g25784 ( n17161 , n9073 , n17044 );
    or g25785 ( n25714 , n26995 , n25344 );
    nor g25786 ( n17737 , n3890 , n12465 );
    nor g25787 ( n10028 , n23865 , n19200 );
    or g25788 ( n19764 , n19050 , n19130 );
    xnor g25789 ( n27158 , n10196 , n2234 );
    nor g25790 ( n5890 , n20323 , n7835 );
    or g25791 ( n10136 , n5580 , n19911 );
    and g25792 ( n6194 , n16866 , n18066 );
    and g25793 ( n19032 , n7524 , n10314 );
    or g25794 ( n1663 , n18639 , n16097 );
    not g25795 ( n23537 , n17183 );
    and g25796 ( n2310 , n15063 , n16253 );
    or g25797 ( n24598 , n25138 , n19784 );
    or g25798 ( n21711 , n10109 , n4007 );
    or g25799 ( n23734 , n26640 , n18175 );
    not g25800 ( n27076 , n7592 );
    not g25801 ( n1449 , n21927 );
    xnor g25802 ( n16940 , n4041 , n3378 );
    nor g25803 ( n11112 , n17453 , n10250 );
    xnor g25804 ( n12508 , n11923 , n17237 );
    xnor g25805 ( n8518 , n16968 , n23120 );
    and g25806 ( n4350 , n6790 , n10000 );
    xnor g25807 ( n25758 , n16197 , n9381 );
    or g25808 ( n24950 , n25724 , n2173 );
    xnor g25809 ( n6130 , n5751 , n25184 );
    nor g25810 ( n25680 , n20409 , n18227 );
    not g25811 ( n762 , n25575 );
    xnor g25812 ( n22639 , n2058 , n5954 );
    xnor g25813 ( n9485 , n9311 , n12829 );
    xnor g25814 ( n12775 , n2510 , n8324 );
    xnor g25815 ( n16279 , n6326 , n2211 );
    and g25816 ( n21374 , n11577 , n24244 );
    or g25817 ( n25236 , n9823 , n25842 );
    nor g25818 ( n26273 , n19039 , n13633 );
    and g25819 ( n8941 , n14439 , n11661 );
    xnor g25820 ( n11812 , n8382 , n10352 );
    and g25821 ( n3167 , n1766 , n25280 );
    nor g25822 ( n17151 , n13453 , n14733 );
    or g25823 ( n23339 , n2126 , n20624 );
    xnor g25824 ( n1324 , n26650 , n23422 );
    or g25825 ( n24674 , n14336 , n9349 );
    not g25826 ( n26095 , n24517 );
    xnor g25827 ( n6733 , n11572 , n23259 );
    xnor g25828 ( n4933 , n2518 , n1637 );
    not g25829 ( n21593 , n23722 );
    nor g25830 ( n26817 , n3737 , n25367 );
    and g25831 ( n21394 , n14450 , n22866 );
    or g25832 ( n4679 , n20289 , n25192 );
    and g25833 ( n12803 , n20571 , n5595 );
    xnor g25834 ( n8314 , n22780 , n5752 );
    not g25835 ( n5993 , n26420 );
    xnor g25836 ( n6536 , n8166 , n26413 );
    xnor g25837 ( n12000 , n13226 , n9324 );
    nor g25838 ( n13924 , n23369 , n18255 );
    nor g25839 ( n23860 , n25929 , n10013 );
    xnor g25840 ( n21266 , n10096 , n16824 );
    not g25841 ( n26951 , n19709 );
    and g25842 ( n6749 , n19530 , n23992 );
    and g25843 ( n21493 , n8204 , n27094 );
    not g25844 ( n22387 , n4112 );
    xnor g25845 ( n9459 , n23972 , n22004 );
    nor g25846 ( n26061 , n21257 , n25935 );
    xnor g25847 ( n18878 , n14440 , n21287 );
    xnor g25848 ( n7946 , n26456 , n14973 );
    or g25849 ( n1666 , n8360 , n18396 );
    not g25850 ( n23408 , n21753 );
    xnor g25851 ( n25605 , n333 , n22091 );
    and g25852 ( n25383 , n5487 , n14682 );
    nor g25853 ( n1796 , n19852 , n23035 );
    xnor g25854 ( n21723 , n23127 , n22908 );
    and g25855 ( n2417 , n12124 , n22429 );
    and g25856 ( n21474 , n19555 , n21655 );
    or g25857 ( n667 , n20044 , n11835 );
    or g25858 ( n18739 , n13248 , n15219 );
    xnor g25859 ( n13069 , n7531 , n26195 );
    not g25860 ( n7429 , n5915 );
    not g25861 ( n16687 , n19890 );
    and g25862 ( n8475 , n9267 , n10808 );
    or g25863 ( n5653 , n15866 , n16552 );
    or g25864 ( n16910 , n21562 , n3865 );
    and g25865 ( n11950 , n7847 , n20195 );
    and g25866 ( n9109 , n4420 , n26975 );
    and g25867 ( n17278 , n5352 , n24339 );
    or g25868 ( n5935 , n21867 , n8557 );
    or g25869 ( n26352 , n17205 , n3042 );
    not g25870 ( n18097 , n7134 );
    or g25871 ( n11067 , n11680 , n24378 );
    not g25872 ( n18357 , n14106 );
    not g25873 ( n23063 , n20138 );
    xnor g25874 ( n1545 , n25051 , n13642 );
    xnor g25875 ( n9841 , n11918 , n20250 );
    xnor g25876 ( n1640 , n7058 , n22625 );
    xnor g25877 ( n5123 , n26994 , n4257 );
    nor g25878 ( n9863 , n23612 , n8167 );
    or g25879 ( n3446 , n21380 , n3018 );
    xnor g25880 ( n2426 , n8964 , n23200 );
    and g25881 ( n18480 , n14842 , n11475 );
    nor g25882 ( n16842 , n22933 , n11185 );
    or g25883 ( n4617 , n23627 , n12165 );
    xnor g25884 ( n6245 , n3109 , n25786 );
    or g25885 ( n893 , n2495 , n18804 );
    or g25886 ( n25084 , n6780 , n961 );
    not g25887 ( n19616 , n4665 );
    or g25888 ( n10439 , n17784 , n725 );
    nor g25889 ( n25414 , n18385 , n22840 );
    or g25890 ( n14793 , n21978 , n19953 );
    or g25891 ( n7844 , n21937 , n9219 );
    xnor g25892 ( n82 , n9251 , n16968 );
    or g25893 ( n11429 , n17824 , n5955 );
    not g25894 ( n7832 , n5559 );
    xnor g25895 ( n4089 , n6259 , n14665 );
    or g25896 ( n25047 , n12762 , n4263 );
    or g25897 ( n22645 , n13447 , n2072 );
    not g25898 ( n1694 , n4616 );
    xnor g25899 ( n11706 , n20967 , n1314 );
    or g25900 ( n18525 , n24625 , n11497 );
    xnor g25901 ( n5252 , n10135 , n552 );
    xnor g25902 ( n15399 , n2060 , n6660 );
    and g25903 ( n25807 , n13753 , n16792 );
    xnor g25904 ( n17771 , n5863 , n20838 );
    not g25905 ( n13368 , n6637 );
    and g25906 ( n11150 , n9882 , n23338 );
    xnor g25907 ( n11071 , n17547 , n13755 );
    xnor g25908 ( n4075 , n12184 , n17322 );
    nor g25909 ( n15722 , n2035 , n26823 );
    and g25910 ( n18614 , n11999 , n5759 );
    not g25911 ( n2891 , n12391 );
    and g25912 ( n24644 , n20866 , n13574 );
    nor g25913 ( n15513 , n6175 , n17967 );
    nor g25914 ( n2617 , n7743 , n2328 );
    and g25915 ( n22680 , n25123 , n15283 );
    and g25916 ( n14210 , n16400 , n17561 );
    or g25917 ( n701 , n11236 , n15231 );
    or g25918 ( n18245 , n2743 , n1584 );
    not g25919 ( n25235 , n9312 );
    and g25920 ( n14867 , n22524 , n2276 );
    or g25921 ( n15545 , n5929 , n24536 );
    xnor g25922 ( n12412 , n13368 , n7260 );
    or g25923 ( n26040 , n68 , n25677 );
    and g25924 ( n16571 , n922 , n13030 );
    xnor g25925 ( n7004 , n16642 , n8386 );
    not g25926 ( n22670 , n2764 );
    xnor g25927 ( n11504 , n3175 , n24973 );
    or g25928 ( n19883 , n25674 , n9992 );
    xnor g25929 ( n12399 , n10372 , n20235 );
    or g25930 ( n1661 , n14130 , n12861 );
    nor g25931 ( n7048 , n26695 , n15944 );
    xnor g25932 ( n14547 , n7615 , n6586 );
    or g25933 ( n24034 , n11443 , n17303 );
    or g25934 ( n24987 , n3506 , n26414 );
    and g25935 ( n8542 , n8895 , n13727 );
    or g25936 ( n2744 , n13159 , n10611 );
    xnor g25937 ( n661 , n16353 , n3485 );
    xnor g25938 ( n18272 , n3687 , n24879 );
    xnor g25939 ( n6371 , n12716 , n18862 );
    nor g25940 ( n3867 , n7442 , n12485 );
    or g25941 ( n23538 , n11349 , n20160 );
    xnor g25942 ( n17068 , n13381 , n6746 );
    nor g25943 ( n27187 , n3610 , n25546 );
    xnor g25944 ( n24404 , n25998 , n17470 );
    nor g25945 ( n635 , n6682 , n23084 );
    and g25946 ( n26742 , n21853 , n20468 );
    and g25947 ( n25768 , n19861 , n13397 );
    not g25948 ( n7465 , n24399 );
    and g25949 ( n4534 , n988 , n24642 );
    or g25950 ( n15080 , n11380 , n5411 );
    xnor g25951 ( n20187 , n5653 , n23959 );
    and g25952 ( n969 , n5544 , n1296 );
    xnor g25953 ( n24318 , n7744 , n2266 );
    xnor g25954 ( n10645 , n21412 , n1195 );
    or g25955 ( n18117 , n2156 , n26332 );
    not g25956 ( n1026 , n22640 );
    not g25957 ( n24974 , n22068 );
    xnor g25958 ( n17653 , n5188 , n18481 );
    or g25959 ( n16563 , n5123 , n15482 );
    not g25960 ( n5948 , n22554 );
    xnor g25961 ( n1604 , n25164 , n9270 );
    xnor g25962 ( n20446 , n14240 , n5865 );
    or g25963 ( n22911 , n17122 , n23383 );
    xnor g25964 ( n1698 , n863 , n25370 );
    and g25965 ( n2786 , n9491 , n8392 );
    xnor g25966 ( n26025 , n15512 , n15147 );
    or g25967 ( n11418 , n21083 , n8052 );
    nor g25968 ( n20852 , n6750 , n14680 );
    xnor g25969 ( n7144 , n7146 , n3549 );
    and g25970 ( n6455 , n9481 , n16741 );
    xnor g25971 ( n8319 , n11551 , n15393 );
    or g25972 ( n16655 , n7689 , n10807 );
    and g25973 ( n22073 , n15455 , n20310 );
    xnor g25974 ( n15278 , n154 , n7722 );
    or g25975 ( n12637 , n26556 , n10917 );
    and g25976 ( n859 , n19911 , n5580 );
    xnor g25977 ( n4407 , n1066 , n25872 );
    or g25978 ( n24885 , n21997 , n15773 );
    xnor g25979 ( n26696 , n56 , n16472 );
    nor g25980 ( n6672 , n8838 , n1987 );
    or g25981 ( n6710 , n442 , n7445 );
    or g25982 ( n7656 , n426 , n19943 );
    or g25983 ( n23869 , n21632 , n13190 );
    and g25984 ( n8712 , n6417 , n21899 );
    xnor g25985 ( n9440 , n22200 , n17805 );
    or g25986 ( n4976 , n15901 , n9418 );
    and g25987 ( n24949 , n18762 , n12027 );
    xnor g25988 ( n5058 , n16083 , n12161 );
    or g25989 ( n3505 , n9465 , n4074 );
    and g25990 ( n17830 , n23408 , n25921 );
    xnor g25991 ( n26562 , n162 , n19568 );
    xnor g25992 ( n13895 , n13781 , n9251 );
    not g25993 ( n7535 , n11876 );
    nor g25994 ( n21781 , n19090 , n17166 );
    xnor g25995 ( n23632 , n6705 , n8614 );
    or g25996 ( n11331 , n6218 , n9296 );
    or g25997 ( n17079 , n15767 , n26733 );
    and g25998 ( n2463 , n26569 , n23465 );
    and g25999 ( n9421 , n15826 , n21585 );
    or g26000 ( n15789 , n8847 , n3651 );
    xnor g26001 ( n22721 , n25974 , n2355 );
    or g26002 ( n11280 , n13340 , n24186 );
    xnor g26003 ( n20678 , n529 , n2488 );
    not g26004 ( n8564 , n21284 );
    or g26005 ( n16980 , n25738 , n6861 );
    xnor g26006 ( n18204 , n3949 , n5961 );
    not g26007 ( n6504 , n15936 );
    xnor g26008 ( n19660 , n16933 , n15672 );
    or g26009 ( n6758 , n13903 , n14073 );
    xnor g26010 ( n1528 , n17573 , n11029 );
    xnor g26011 ( n15593 , n15087 , n23272 );
    or g26012 ( n18658 , n13546 , n9831 );
    not g26013 ( n23681 , n789 );
    or g26014 ( n4367 , n16462 , n10135 );
    and g26015 ( n10937 , n2628 , n8786 );
    nor g26016 ( n4312 , n14830 , n26584 );
    xnor g26017 ( n24307 , n12020 , n5164 );
    xnor g26018 ( n4774 , n15185 , n22169 );
    or g26019 ( n22813 , n5221 , n2157 );
    xnor g26020 ( n18125 , n1453 , n27179 );
    not g26021 ( n6521 , n5101 );
    nor g26022 ( n19557 , n19673 , n5678 );
    xnor g26023 ( n11557 , n10767 , n4031 );
    or g26024 ( n13432 , n15238 , n4571 );
    or g26025 ( n7609 , n24665 , n1687 );
    or g26026 ( n5672 , n20206 , n10250 );
    and g26027 ( n21200 , n6621 , n10062 );
    not g26028 ( n2597 , n11121 );
    nor g26029 ( n25530 , n16562 , n15170 );
    or g26030 ( n26692 , n12422 , n19087 );
    xnor g26031 ( n20933 , n5153 , n12548 );
    not g26032 ( n26100 , n19143 );
    nor g26033 ( n16475 , n15012 , n7401 );
    and g26034 ( n13604 , n8177 , n3585 );
    or g26035 ( n17416 , n23709 , n16267 );
    or g26036 ( n22424 , n483 , n6566 );
    xnor g26037 ( n20802 , n2608 , n13553 );
    xnor g26038 ( n12852 , n4459 , n19391 );
    or g26039 ( n2793 , n24876 , n24037 );
    xnor g26040 ( n13466 , n26289 , n14273 );
    xnor g26041 ( n4242 , n11361 , n13208 );
    xnor g26042 ( n1802 , n1456 , n10405 );
    or g26043 ( n16316 , n2355 , n16223 );
    and g26044 ( n25856 , n12921 , n17197 );
    not g26045 ( n6070 , n16900 );
    nor g26046 ( n6244 , n21880 , n9007 );
    xnor g26047 ( n725 , n7535 , n9003 );
    xnor g26048 ( n1845 , n20538 , n17873 );
    nor g26049 ( n5518 , n14777 , n21442 );
    or g26050 ( n1832 , n27202 , n15949 );
    or g26051 ( n25175 , n25050 , n23281 );
    and g26052 ( n4213 , n20554 , n25806 );
    or g26053 ( n16143 , n364 , n6083 );
    xnor g26054 ( n11414 , n22916 , n11213 );
    xnor g26055 ( n9199 , n10861 , n21857 );
    or g26056 ( n19079 , n12800 , n26498 );
    xnor g26057 ( n12273 , n19429 , n14610 );
    xnor g26058 ( n21683 , n17397 , n18227 );
    xnor g26059 ( n18950 , n6960 , n10150 );
    or g26060 ( n12432 , n566 , n374 );
    or g26061 ( n9041 , n10983 , n23562 );
    xnor g26062 ( n21567 , n23536 , n14899 );
    and g26063 ( n10652 , n20232 , n12970 );
    xnor g26064 ( n8823 , n11816 , n24954 );
    not g26065 ( n12354 , n8920 );
    or g26066 ( n25146 , n2606 , n17211 );
    xnor g26067 ( n16719 , n20920 , n17911 );
    xnor g26068 ( n21740 , n9769 , n15955 );
    and g26069 ( n20744 , n24255 , n9604 );
    not g26070 ( n310 , n8729 );
    or g26071 ( n23183 , n26947 , n15639 );
    xnor g26072 ( n11733 , n26924 , n24861 );
    not g26073 ( n19588 , n15884 );
    and g26074 ( n9701 , n23665 , n13355 );
    xnor g26075 ( n19143 , n7594 , n6991 );
    nor g26076 ( n21767 , n23512 , n9124 );
    xnor g26077 ( n15135 , n16700 , n9321 );
    or g26078 ( n3108 , n6580 , n11350 );
    or g26079 ( n4034 , n11665 , n20211 );
    not g26080 ( n3045 , n4618 );
    xnor g26081 ( n14222 , n20812 , n24596 );
    or g26082 ( n17238 , n14117 , n5824 );
    nor g26083 ( n24469 , n9502 , n2168 );
    or g26084 ( n837 , n8745 , n8479 );
    xnor g26085 ( n25773 , n16076 , n1728 );
    xnor g26086 ( n7583 , n11841 , n17077 );
    xnor g26087 ( n4293 , n7451 , n8874 );
    and g26088 ( n241 , n24426 , n3574 );
    and g26089 ( n10977 , n3627 , n9367 );
    and g26090 ( n21416 , n25494 , n10713 );
    or g26091 ( n2974 , n26324 , n6359 );
    nor g26092 ( n7000 , n23141 , n1370 );
    xnor g26093 ( n5064 , n568 , n14865 );
    and g26094 ( n11729 , n11035 , n25266 );
    nor g26095 ( n3977 , n25475 , n23697 );
    or g26096 ( n14641 , n26793 , n25067 );
    and g26097 ( n23072 , n921 , n10590 );
    or g26098 ( n21811 , n12713 , n180 );
    xnor g26099 ( n16659 , n21613 , n6242 );
    not g26100 ( n26467 , n560 );
    or g26101 ( n11629 , n6234 , n14384 );
    xnor g26102 ( n9797 , n24770 , n13445 );
    xnor g26103 ( n13869 , n14754 , n26344 );
    nor g26104 ( n4876 , n15182 , n26797 );
    or g26105 ( n6116 , n20159 , n10884 );
    not g26106 ( n21450 , n9110 );
    or g26107 ( n21569 , n10578 , n5901 );
    not g26108 ( n15826 , n23146 );
    or g26109 ( n20348 , n13561 , n14148 );
    not g26110 ( n26677 , n4335 );
    or g26111 ( n12197 , n17128 , n26912 );
    xnor g26112 ( n24829 , n3131 , n22442 );
    xnor g26113 ( n3151 , n10057 , n5026 );
    or g26114 ( n19901 , n11452 , n26823 );
    xnor g26115 ( n4150 , n13394 , n5997 );
    not g26116 ( n24417 , n5822 );
    or g26117 ( n8860 , n16755 , n20326 );
    xnor g26118 ( n2938 , n26799 , n12059 );
    or g26119 ( n23535 , n2331 , n4587 );
    or g26120 ( n11495 , n20133 , n5255 );
    xnor g26121 ( n638 , n2224 , n20603 );
    or g26122 ( n6064 , n13351 , n7622 );
    nor g26123 ( n25320 , n6724 , n6127 );
    not g26124 ( n10711 , n19107 );
    or g26125 ( n8187 , n5446 , n22647 );
    nor g26126 ( n25644 , n811 , n13609 );
    or g26127 ( n17387 , n18855 , n8787 );
    xnor g26128 ( n8523 , n3173 , n25393 );
    and g26129 ( n1679 , n22290 , n12878 );
    xnor g26130 ( n3097 , n24350 , n6062 );
    xnor g26131 ( n4356 , n26773 , n19301 );
    nor g26132 ( n23245 , n16687 , n20906 );
    and g26133 ( n5405 , n18955 , n11887 );
    or g26134 ( n6976 , n4471 , n8168 );
    or g26135 ( n1124 , n14895 , n24409 );
    or g26136 ( n15833 , n11622 , n9276 );
    and g26137 ( n16538 , n20194 , n12089 );
    or g26138 ( n25333 , n7953 , n13894 );
    nor g26139 ( n12614 , n21823 , n11702 );
    or g26140 ( n9999 , n26380 , n18974 );
    or g26141 ( n13957 , n6898 , n6448 );
    xnor g26142 ( n22972 , n17656 , n25267 );
    not g26143 ( n26307 , n14366 );
    nor g26144 ( n844 , n11302 , n24786 );
    or g26145 ( n21490 , n11339 , n5870 );
    or g26146 ( n24066 , n2137 , n11085 );
    or g26147 ( n3537 , n25674 , n21832 );
    xnor g26148 ( n26541 , n1010 , n9238 );
    not g26149 ( n2080 , n8708 );
    and g26150 ( n10654 , n3756 , n4354 );
    xnor g26151 ( n9006 , n3909 , n268 );
    or g26152 ( n1649 , n20530 , n11394 );
    or g26153 ( n11857 , n11544 , n2160 );
    or g26154 ( n9117 , n4435 , n8533 );
    and g26155 ( n19721 , n7804 , n4716 );
    not g26156 ( n23036 , n21879 );
    or g26157 ( n1208 , n21148 , n15988 );
    xnor g26158 ( n17643 , n3837 , n1040 );
    nor g26159 ( n18119 , n22198 , n575 );
    xnor g26160 ( n16337 , n11580 , n2035 );
    not g26161 ( n20146 , n4851 );
    xnor g26162 ( n3344 , n1370 , n26054 );
    not g26163 ( n23865 , n24106 );
    xnor g26164 ( n9648 , n10871 , n17637 );
    or g26165 ( n22168 , n10097 , n11974 );
    xnor g26166 ( n17754 , n19534 , n13319 );
    xnor g26167 ( n18610 , n1497 , n433 );
    or g26168 ( n18740 , n10802 , n15903 );
    nor g26169 ( n263 , n20311 , n20741 );
    and g26170 ( n22630 , n2504 , n25860 );
    nor g26171 ( n17537 , n15715 , n14954 );
    or g26172 ( n24586 , n21538 , n6725 );
    or g26173 ( n14060 , n13017 , n21483 );
    xnor g26174 ( n16441 , n23913 , n3710 );
    and g26175 ( n16381 , n4761 , n8683 );
    xnor g26176 ( n10448 , n4018 , n19747 );
    or g26177 ( n18354 , n10963 , n12969 );
    not g26178 ( n24666 , n6606 );
    or g26179 ( n660 , n17580 , n11008 );
    and g26180 ( n24525 , n5888 , n4653 );
    and g26181 ( n20452 , n14806 , n10270 );
    and g26182 ( n18893 , n24494 , n14080 );
    or g26183 ( n5778 , n21972 , n17120 );
    xnor g26184 ( n1982 , n10571 , n9172 );
    not g26185 ( n23441 , n11266 );
    and g26186 ( n8890 , n6611 , n26895 );
    xnor g26187 ( n24117 , n17564 , n26196 );
    not g26188 ( n7071 , n24608 );
    xnor g26189 ( n4714 , n7488 , n13310 );
    xnor g26190 ( n17395 , n27170 , n1136 );
    xnor g26191 ( n12663 , n25691 , n13783 );
    xnor g26192 ( n2742 , n21912 , n9291 );
    xnor g26193 ( n4804 , n15267 , n2010 );
    xnor g26194 ( n2841 , n21075 , n16828 );
    xnor g26195 ( n7791 , n23280 , n4162 );
    nor g26196 ( n5514 , n7130 , n2044 );
    and g26197 ( n10 , n20201 , n20231 );
    xnor g26198 ( n17342 , n15053 , n3828 );
    not g26199 ( n20945 , n12445 );
    or g26200 ( n26331 , n3972 , n14396 );
    xnor g26201 ( n8622 , n2231 , n14070 );
    nor g26202 ( n24623 , n12713 , n24701 );
    xnor g26203 ( n13595 , n5938 , n5987 );
    xnor g26204 ( n3474 , n3560 , n8863 );
    xnor g26205 ( n17690 , n272 , n19291 );
    xnor g26206 ( n330 , n6340 , n23667 );
    nor g26207 ( n9823 , n7377 , n5629 );
    or g26208 ( n1445 , n20261 , n13632 );
    and g26209 ( n12747 , n24531 , n13852 );
    xnor g26210 ( n13354 , n8704 , n3488 );
    or g26211 ( n7176 , n25342 , n16662 );
    xnor g26212 ( n10298 , n18601 , n13533 );
    or g26213 ( n10648 , n11393 , n13359 );
    not g26214 ( n1780 , n19087 );
    xnor g26215 ( n25735 , n9700 , n25210 );
    not g26216 ( n18607 , n22826 );
    xnor g26217 ( n9532 , n23722 , n20972 );
    xnor g26218 ( n1249 , n12075 , n4957 );
    xnor g26219 ( n19711 , n22930 , n19327 );
    nor g26220 ( n21052 , n24825 , n21317 );
    xnor g26221 ( n14184 , n3876 , n3748 );
    or g26222 ( n22324 , n20820 , n16058 );
    not g26223 ( n21613 , n23411 );
    or g26224 ( n20819 , n10194 , n9597 );
    xnor g26225 ( n20999 , n2080 , n1319 );
    not g26226 ( n8582 , n19904 );
    not g26227 ( n4575 , n9545 );
    nor g26228 ( n22855 , n21957 , n14156 );
    and g26229 ( n12368 , n490 , n26755 );
    nor g26230 ( n13106 , n25126 , n19575 );
    or g26231 ( n8091 , n5044 , n10635 );
    nor g26232 ( n9249 , n25797 , n15784 );
    or g26233 ( n14812 , n25762 , n15612 );
    and g26234 ( n17303 , n11362 , n6326 );
    or g26235 ( n22320 , n11559 , n16693 );
    or g26236 ( n8755 , n19706 , n4720 );
    and g26237 ( n7318 , n4973 , n16815 );
    xnor g26238 ( n9219 , n17923 , n1752 );
    xnor g26239 ( n11824 , n20007 , n11799 );
    or g26240 ( n6605 , n13898 , n6502 );
    and g26241 ( n22848 , n19598 , n4251 );
    xnor g26242 ( n19947 , n10833 , n4042 );
    xnor g26243 ( n9344 , n14413 , n9175 );
    or g26244 ( n11478 , n18224 , n6640 );
    or g26245 ( n22957 , n8749 , n12972 );
    or g26246 ( n6573 , n12022 , n8889 );
    xnor g26247 ( n4103 , n11164 , n22251 );
    xnor g26248 ( n6915 , n14876 , n2472 );
    xnor g26249 ( n6458 , n22176 , n19922 );
    nor g26250 ( n6201 , n19439 , n22747 );
    xnor g26251 ( n22531 , n1690 , n1000 );
    and g26252 ( n4803 , n3018 , n21380 );
    xnor g26253 ( n21462 , n12638 , n7026 );
    xnor g26254 ( n22546 , n23313 , n2586 );
    and g26255 ( n24296 , n13128 , n10662 );
    not g26256 ( n10314 , n1541 );
    nor g26257 ( n1179 , n17705 , n22421 );
    or g26258 ( n2940 , n23234 , n7682 );
    or g26259 ( n18147 , n7290 , n18758 );
    not g26260 ( n7529 , n2646 );
    and g26261 ( n16032 , n2710 , n1124 );
    or g26262 ( n18251 , n19652 , n21916 );
    xnor g26263 ( n15300 , n13599 , n564 );
    or g26264 ( n19787 , n200 , n25247 );
    and g26265 ( n17955 , n14586 , n14729 );
    nor g26266 ( n15200 , n25041 , n25643 );
    xnor g26267 ( n3332 , n16123 , n497 );
    or g26268 ( n11859 , n678 , n3921 );
    xnor g26269 ( n2211 , n15616 , n9215 );
    xnor g26270 ( n3209 , n6703 , n11321 );
    or g26271 ( n26624 , n13406 , n8471 );
    or g26272 ( n8671 , n21293 , n2926 );
    nor g26273 ( n6929 , n10966 , n19789 );
    nor g26274 ( n27182 , n20840 , n21948 );
    not g26275 ( n10691 , n20210 );
    not g26276 ( n2872 , n20731 );
    not g26277 ( n15131 , n4890 );
    xnor g26278 ( n2327 , n17321 , n1053 );
    and g26279 ( n25699 , n6222 , n9744 );
    nor g26280 ( n18560 , n642 , n21194 );
    and g26281 ( n1400 , n9594 , n5915 );
    xnor g26282 ( n21940 , n725 , n24804 );
    not g26283 ( n25403 , n22008 );
    xnor g26284 ( n13276 , n19520 , n20077 );
    and g26285 ( n5138 , n17457 , n10828 );
    nor g26286 ( n8932 , n6915 , n9748 );
    or g26287 ( n12994 , n1263 , n9885 );
    xnor g26288 ( n6884 , n4479 , n11986 );
    not g26289 ( n12184 , n16494 );
    xnor g26290 ( n2989 , n4199 , n23101 );
    or g26291 ( n12199 , n18511 , n14361 );
    xnor g26292 ( n2578 , n6761 , n7122 );
    or g26293 ( n23062 , n2027 , n26942 );
    xnor g26294 ( n16846 , n5100 , n14200 );
    or g26295 ( n9352 , n19836 , n3835 );
    not g26296 ( n13249 , n2784 );
    nor g26297 ( n7939 , n4801 , n9723 );
    or g26298 ( n18469 , n15260 , n26148 );
    or g26299 ( n4466 , n23932 , n10666 );
    not g26300 ( n9572 , n16201 );
    or g26301 ( n22018 , n10873 , n25250 );
    xnor g26302 ( n15831 , n20657 , n3799 );
    or g26303 ( n749 , n24330 , n5320 );
    and g26304 ( n12387 , n26565 , n9142 );
    xnor g26305 ( n7310 , n23921 , n11302 );
    xnor g26306 ( n14835 , n6011 , n13137 );
    or g26307 ( n20310 , n18085 , n5157 );
    xnor g26308 ( n19724 , n1405 , n3317 );
    not g26309 ( n7327 , n18988 );
    xnor g26310 ( n11696 , n16396 , n8399 );
    or g26311 ( n9271 , n27155 , n10803 );
    xnor g26312 ( n10027 , n1123 , n26137 );
    or g26313 ( n659 , n24755 , n22295 );
    nor g26314 ( n15453 , n26363 , n1553 );
    or g26315 ( n21346 , n25324 , n1642 );
    xnor g26316 ( n12648 , n5075 , n9241 );
    or g26317 ( n675 , n20921 , n25106 );
    xnor g26318 ( n2666 , n21704 , n7751 );
    xnor g26319 ( n10573 , n19978 , n24239 );
    xnor g26320 ( n9645 , n2705 , n19551 );
    or g26321 ( n226 , n718 , n7158 );
    nor g26322 ( n18386 , n8351 , n11066 );
    nor g26323 ( n25176 , n3382 , n18363 );
    not g26324 ( n5719 , n468 );
    xnor g26325 ( n11129 , n455 , n6387 );
    not g26326 ( n16937 , n7149 );
    xnor g26327 ( n23801 , n11579 , n3962 );
    or g26328 ( n1615 , n11393 , n12956 );
    xnor g26329 ( n22215 , n1645 , n3978 );
    xnor g26330 ( n11945 , n20177 , n14946 );
    or g26331 ( n18320 , n19905 , n2547 );
    not g26332 ( n8367 , n25749 );
    and g26333 ( n25537 , n18996 , n23461 );
    xnor g26334 ( n7526 , n19633 , n5427 );
    nor g26335 ( n16497 , n677 , n24243 );
    and g26336 ( n25262 , n24852 , n20487 );
    or g26337 ( n13314 , n19042 , n18846 );
    xnor g26338 ( n23550 , n17602 , n14843 );
    or g26339 ( n25151 , n12371 , n10534 );
    not g26340 ( n9490 , n17653 );
    xnor g26341 ( n5750 , n13616 , n20263 );
    or g26342 ( n22504 , n16309 , n20391 );
    or g26343 ( n17093 , n22741 , n3944 );
    not g26344 ( n5065 , n6819 );
    xnor g26345 ( n12265 , n21197 , n6125 );
    xnor g26346 ( n13155 , n10312 , n10013 );
    or g26347 ( n26487 , n14079 , n5758 );
    or g26348 ( n8992 , n14292 , n9876 );
    xnor g26349 ( n7060 , n5390 , n5081 );
    xnor g26350 ( n6278 , n14254 , n14610 );
    and g26351 ( n5996 , n4179 , n10959 );
    xnor g26352 ( n26509 , n5852 , n19971 );
    or g26353 ( n17153 , n26139 , n2952 );
    xnor g26354 ( n4266 , n17724 , n22633 );
    xnor g26355 ( n22787 , n7422 , n20917 );
    xnor g26356 ( n13075 , n23097 , n19568 );
    or g26357 ( n22103 , n17551 , n8785 );
    or g26358 ( n13105 , n19673 , n12416 );
    not g26359 ( n3778 , n3859 );
    nor g26360 ( n23452 , n17223 , n4488 );
    or g26361 ( n12504 , n9766 , n16918 );
    or g26362 ( n12787 , n10201 , n19691 );
    not g26363 ( n3840 , n7797 );
    xnor g26364 ( n15927 , n5143 , n19625 );
    xnor g26365 ( n26931 , n23331 , n20604 );
    and g26366 ( n20745 , n17088 , n5241 );
endmodule
