// Benchmark "top" written by ABC on Sun Dec 21 18:07:32 2025

module top ( 
    n1, n9, n67, n69, n84, n96, n107, n120, n128, n135, n137, n145, n147,
    n182, n184, n198, n209, n220, n222, n230, n233, n268, n283, n289, n290,
    n293, n296, n325, n330, n342, n356, n362, n365, n373, n386, n403, n415,
    n418, n421, n432, n468, n478, n481, n490, n507, n514, n526, n532, n574,
    n576, n579, n588, n596, n605, n615, n629, n635, n646, n654, n664, n677,
    n704, n710, n716, n726, n727, n737, n750, n751, n765, n769, n793, n794,
    n797, n818, n824, n829, n835, n837, n842, n848, n851, n857, n859, n869,
    n877, n901, n909, n923, n933, n934, n938, n950, n956, n973, n974, n989,
    n990, n1013, n1014, n1025, n1030, n1042, n1049, n1052, n1058, n1065,
    n1070, n1091, n1093, n1098, n1099, n1108, n1121, n1131, n1134, n1143,
    n1146, n1150, n1161, n1162, n1165, n1170, n1184, n1187, n1189, n1223,
    n1240, n1243, n1251, n1253, n1255, n1276, n1280, n1303, n1310, n1311,
    n1331, n1335, n1339, n1361, n1366, n1373, n1378, n1389, n1396, n1398,
    n1407, n1409, n1412, n1413, n1418, n1422, n1425, n1438, n1475, n1479,
    n1485, n1508, n1511, n1515, n1518, n1530, n1545, n1549, n1551, n1555,
    n1562, n1575, n1580, n1581, n1596, n1606, n1620, n1630, n1648, n1655,
    n1676,
    n8, n21, n24, n32, n54, n61, n64, n76, n83, n97, n110, n117, n142,
    n150, n154, n167, n170, n172, n190, n204, n210, n231, n232, n240, n253,
    n265, n269, n291, n292, n313, n324, n336, n347, n350, n363, n364, n368,
    n383, n388, n427, n434, n476, n480, n489, n506, n524, n543, n565, n598,
    n608, n614, n618, n623, n633, n640, n656, n663, n675, n676, n678, n691,
    n693, n717, n722, n740, n785, n786, n790, n800, n814, n821, n836, n840,
    n845, n887, n894, n928, n964, n1019, n1021, n1023, n1026, n1032, n1036,
    n1039, n1043, n1117, n1122, n1138, n1151, n1157, n1160, n1177, n1192,
    n1194, n1198, n1239, n1275, n1314, n1375, n1392, n1411, n1442, n1454,
    n1474, n1478, n1512, n1531, n1542, n1547, n1552, n1556, n1574, n1589,
    n1594, n1601, n1604, n1628, n1629, n1631, n1645, n1665, n1671  );
  input  n1, n9, n67, n69, n84, n96, n107, n120, n128, n135, n137, n145,
    n147, n182, n184, n198, n209, n220, n222, n230, n233, n268, n283, n289,
    n290, n293, n296, n325, n330, n342, n356, n362, n365, n373, n386, n403,
    n415, n418, n421, n432, n468, n478, n481, n490, n507, n514, n526, n532,
    n574, n576, n579, n588, n596, n605, n615, n629, n635, n646, n654, n664,
    n677, n704, n710, n716, n726, n727, n737, n750, n751, n765, n769, n793,
    n794, n797, n818, n824, n829, n835, n837, n842, n848, n851, n857, n859,
    n869, n877, n901, n909, n923, n933, n934, n938, n950, n956, n973, n974,
    n989, n990, n1013, n1014, n1025, n1030, n1042, n1049, n1052, n1058,
    n1065, n1070, n1091, n1093, n1098, n1099, n1108, n1121, n1131, n1134,
    n1143, n1146, n1150, n1161, n1162, n1165, n1170, n1184, n1187, n1189,
    n1223, n1240, n1243, n1251, n1253, n1255, n1276, n1280, n1303, n1310,
    n1311, n1331, n1335, n1339, n1361, n1366, n1373, n1378, n1389, n1396,
    n1398, n1407, n1409, n1412, n1413, n1418, n1422, n1425, n1438, n1475,
    n1479, n1485, n1508, n1511, n1515, n1518, n1530, n1545, n1549, n1551,
    n1555, n1562, n1575, n1580, n1581, n1596, n1606, n1620, n1630, n1648,
    n1655, n1676;
  output n8, n21, n24, n32, n54, n61, n64, n76, n83, n97, n110, n117, n142,
    n150, n154, n167, n170, n172, n190, n204, n210, n231, n232, n240, n253,
    n265, n269, n291, n292, n313, n324, n336, n347, n350, n363, n364, n368,
    n383, n388, n427, n434, n476, n480, n489, n506, n524, n543, n565, n598,
    n608, n614, n618, n623, n633, n640, n656, n663, n675, n676, n678, n691,
    n693, n717, n722, n740, n785, n786, n790, n800, n814, n821, n836, n840,
    n845, n887, n894, n928, n964, n1019, n1021, n1023, n1026, n1032, n1036,
    n1039, n1043, n1117, n1122, n1138, n1151, n1157, n1160, n1177, n1192,
    n1194, n1198, n1239, n1275, n1314, n1375, n1392, n1411, n1442, n1454,
    n1474, n1478, n1512, n1531, n1542, n1547, n1552, n1556, n1574, n1589,
    n1594, n1601, n1604, n1628, n1629, n1631, n1645, n1665, n1671;
  wire new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313_1, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324_1, new_n325_1, new_n326, new_n327, new_n328,
    new_n329, new_n330_1, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336_1, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342_1, new_n343, new_n344, new_n345, new_n346, new_n347_1,
    new_n348, new_n349, new_n350_1, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356_1, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362_1, new_n363_1, new_n364_1, new_n365_1, new_n366, new_n367,
    new_n368_1, new_n369, new_n370, new_n371, new_n372, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n384, new_n385, new_n386_1, new_n387, new_n388_1, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403_1,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415_1, new_n416, new_n417,
    new_n418_1, new_n419, new_n420, new_n421_1, new_n422, new_n423,
    new_n424, new_n425, new_n426, new_n427_1, new_n428, new_n429, new_n430,
    new_n431, new_n432_1, new_n433, new_n434_1, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468_1, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n476_1, new_n477, new_n478_1,
    new_n479, new_n480_1, new_n481_1, new_n482, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489_1, new_n490_1, new_n491,
    new_n492, new_n493, new_n494, new_n495, new_n496, new_n497, new_n498,
    new_n499, new_n500, new_n501, new_n503, new_n504, new_n505, new_n506_1,
    new_n507_1, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514_1, new_n515, new_n516, new_n517, new_n519, new_n520, new_n521,
    new_n522, new_n523, new_n524_1, new_n525, new_n526_1, new_n528,
    new_n529, new_n530, new_n531, new_n532_1, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543_1, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565_1, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574_1, new_n575, new_n576_1,
    new_n577, new_n578, new_n579_1, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588_1, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596_1, new_n597,
    new_n598_1, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605_1, new_n606, new_n607, new_n608_1, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614_1, new_n615_1, new_n616,
    new_n617, new_n618_1, new_n619, new_n620, new_n621, new_n622,
    new_n623_1, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629_1, new_n630, new_n631, new_n632, new_n633_1, new_n634,
    new_n635_1, new_n636, new_n637, new_n638, new_n639, new_n640_1,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646_1, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654_1,
    new_n655, new_n656_1, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663_1, new_n664_1, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675_1, new_n676_1, new_n677_1, new_n678_1, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691_1, new_n692, new_n693_1,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704_1, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710_1, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716_1, new_n717_1, new_n718, new_n719, new_n720,
    new_n721, new_n722_1, new_n723, new_n724, new_n725, new_n726_1,
    new_n727_1, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737_1, new_n738, new_n739,
    new_n740_1, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750_1, new_n751_1, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765_1, new_n766,
    new_n767, new_n768, new_n769_1, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785_1, new_n786_1,
    new_n787, new_n788, new_n789, new_n790_1, new_n791, new_n792,
    new_n793_1, new_n794_1, new_n795, new_n796, new_n797_1, new_n798,
    new_n799, new_n800_1, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814_1, new_n815, new_n816, new_n817, new_n818_1,
    new_n819, new_n820, new_n821_1, new_n822, new_n823, new_n824_1,
    new_n825, new_n826, new_n827, new_n828, new_n829_1, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835_1, new_n836_1, new_n837_1,
    new_n838, new_n839, new_n840_1, new_n841, new_n842_1, new_n843,
    new_n844, new_n845_1, new_n846, new_n847, new_n848_1, new_n849,
    new_n850, new_n851_1, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857_1, new_n858, new_n859_1, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869_1,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877_1, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887_1, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894_1, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901_1, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909_1, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923_1, new_n924, new_n925, new_n926, new_n927,
    new_n928_1, new_n929, new_n930, new_n931, new_n932, new_n933_1,
    new_n934_1, new_n935, new_n936, new_n937, new_n938_1, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950_1, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956_1, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974_1, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989_1, new_n990_1, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013_1,
    new_n1014_1, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019_1,
    new_n1020, new_n1021_1, new_n1022, new_n1023_1, new_n1024, new_n1025_1,
    new_n1026_1, new_n1027, new_n1028, new_n1029, new_n1030_1, new_n1031,
    new_n1032_1, new_n1033, new_n1034, new_n1035, new_n1036_1, new_n1038,
    new_n1040, new_n1041, new_n1042_1, new_n1043_1, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049_1, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1062, new_n1063, new_n1064, new_n1065_1, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070_1, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091_1,
    new_n1093_1, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098_1,
    new_n1099_1, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108_1, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1117_1,
    new_n1118, new_n1119, new_n1120, new_n1121_1, new_n1122_1, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1132, new_n1133, new_n1134_1, new_n1135, new_n1136, new_n1138_1,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143_1, new_n1144,
    new_n1146_1, new_n1147, new_n1149, new_n1150_1, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1157_1, new_n1158, new_n1159, new_n1160_1,
    new_n1161_1, new_n1163, new_n1164, new_n1165_1, new_n1166, new_n1167,
    new_n1168, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1178, new_n1179, new_n1180, new_n1181, new_n1183,
    new_n1184_1, new_n1185, new_n1186, new_n1187_1, new_n1188, new_n1189_1,
    new_n1191, new_n1192_1, new_n1193, new_n1194_1, new_n1196, new_n1197,
    new_n1198_1, new_n1199, new_n1200, new_n1201, new_n1202, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223_1, new_n1224,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239_1, new_n1241, new_n1242, new_n1243_1, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1249, new_n1250, new_n1251_1, new_n1252,
    new_n1253_1, new_n1254, new_n1255_1, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275_1, new_n1276_1, new_n1277, new_n1278, new_n1279, new_n1280_1,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303_1, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310_1, new_n1311_1,
    new_n1312, new_n1313, new_n1314_1, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1327, new_n1328, new_n1329, new_n1330,
    new_n1332, new_n1333, new_n1334, new_n1335_1, new_n1336, new_n1337,
    new_n1339_1, new_n1340, new_n1341, new_n1342, new_n1344, new_n1345,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361_1, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366_1, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1375_1, new_n1376, new_n1377, new_n1378_1,
    new_n1380, new_n1381, new_n1382, new_n1383, new_n1384, new_n1385,
    new_n1387, new_n1389_1, new_n1390, new_n1391, new_n1393, new_n1394,
    new_n1395, new_n1396_1, new_n1397, new_n1398_1, new_n1399, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406, new_n1407_1,
    new_n1409_1, new_n1411_1, new_n1412_1, new_n1413_1, new_n1414,
    new_n1415, new_n1416, new_n1417, new_n1418_1, new_n1419, new_n1420,
    new_n1421, new_n1422_1, new_n1423, new_n1424, new_n1425_1, new_n1426,
    new_n1427, new_n1428, new_n1429, new_n1430, new_n1431, new_n1432,
    new_n1433, new_n1436, new_n1437, new_n1438_1, new_n1439, new_n1440,
    new_n1442_1, new_n1443, new_n1444, new_n1446, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1453, new_n1454_1, new_n1455,
    new_n1456, new_n1457, new_n1458, new_n1459, new_n1461, new_n1462,
    new_n1463, new_n1464, new_n1465, new_n1466, new_n1468, new_n1469,
    new_n1470, new_n1471, new_n1472, new_n1473, new_n1474_1, new_n1476,
    new_n1477, new_n1478_1, new_n1479_1, new_n1480, new_n1481, new_n1483,
    new_n1484, new_n1485_1, new_n1486, new_n1487, new_n1488, new_n1489,
    new_n1491, new_n1492, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1499, new_n1500, new_n1501, new_n1502, new_n1503,
    new_n1504, new_n1506, new_n1507, new_n1508_1, new_n1510, new_n1511_1,
    new_n1512_1, new_n1513, new_n1514, new_n1515_1, new_n1517, new_n1518_1,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1524, new_n1525,
    new_n1526, new_n1527, new_n1528, new_n1529, new_n1530_1, new_n1532,
    new_n1533, new_n1534, new_n1535, new_n1536, new_n1537, new_n1540,
    new_n1541, new_n1542_1, new_n1543, new_n1544, new_n1545_1, new_n1546,
    new_n1548, new_n1549_1, new_n1550, new_n1551_1, new_n1552_1, new_n1553,
    new_n1555_1, new_n1556_1, new_n1557, new_n1560, new_n1561, new_n1562_1,
    new_n1563, new_n1564, new_n1565, new_n1567, new_n1568, new_n1569,
    new_n1570, new_n1571, new_n1572, new_n1573, new_n1576, new_n1577,
    new_n1578, new_n1579, new_n1580_1, new_n1581_1;
  assign new_n302 = ~n1551 & ~n1655;
  assign new_n303 = n532 & ~n1065;
  assign new_n304 = n1170 & n1606;
  assign new_n305 = n1335 & ~n1606;
  assign new_n306 = ~new_n304 & ~new_n305;
  assign new_n307 = n842 & n1606;
  assign new_n308 = n629 & ~n1606;
  assign new_n309 = ~new_n307 & ~new_n308;
  assign new_n310 = new_n306 & new_n309;
  assign new_n311 = n1223 & n1606;
  assign new_n312 = n490 & ~n1606;
  assign new_n313_1 = ~new_n311 & ~new_n312;
  assign new_n314 = n1165 & ~new_n313_1;
  assign new_n315 = n1025 & n1606;
  assign new_n316 = n654 & ~n1606;
  assign new_n317 = ~new_n315 & ~new_n316;
  assign new_n318 = n1389 & ~new_n317;
  assign new_n319 = ~n1165 & new_n313_1;
  assign new_n320 = ~new_n314 & ~new_n319;
  assign new_n321 = new_n318 & new_n320;
  assign new_n322 = ~new_n314 & ~new_n321;
  assign new_n323 = n727 & n1606;
  assign new_n324_1 = n1058 & ~n1606;
  assign new_n325_1 = ~new_n323 & ~new_n324_1;
  assign new_n326 = n403 & ~new_n325_1;
  assign new_n327 = ~n403 & new_n325_1;
  assign new_n328 = ~n574 & n1606;
  assign new_n329 = n1545 & ~new_n328;
  assign new_n330_1 = n1013 & n1606;
  assign new_n331 = n1161 & ~n1606;
  assign new_n332 = ~new_n330_1 & ~new_n331;
  assign new_n333 = n1596 & n1606;
  assign new_n334 = n1518 & ~n1606;
  assign new_n335 = ~new_n333 & ~new_n334;
  assign new_n336_1 = ~n769 & new_n335;
  assign new_n337 = n481 & n1606;
  assign new_n338 = n646 & ~n1606;
  assign new_n339 = ~new_n337 & ~new_n338;
  assign new_n340 = n1378 & ~new_n339;
  assign new_n341 = n769 & ~new_n335;
  assign new_n342_1 = ~new_n340 & ~new_n341;
  assign new_n343 = ~new_n336_1 & ~new_n342_1;
  assign new_n344 = new_n332 & ~new_n343;
  assign new_n345 = ~n1545 & new_n328;
  assign new_n346 = ~n1378 & new_n339;
  assign new_n347_1 = ~new_n340 & ~new_n346;
  assign new_n348 = ~new_n336_1 & ~new_n341;
  assign new_n349 = new_n347_1 & new_n348;
  assign new_n350_1 = ~new_n343 & ~new_n349;
  assign new_n351 = ~new_n345 & ~new_n350_1;
  assign new_n352 = ~new_n344 & new_n351;
  assign new_n353 = ~new_n329 & ~new_n352;
  assign new_n354 = ~new_n327 & ~new_n353;
  assign new_n355 = ~new_n326 & ~new_n354;
  assign new_n356_1 = ~new_n329 & ~new_n345;
  assign new_n357 = new_n349 & new_n356_1;
  assign new_n358 = ~new_n326 & ~new_n327;
  assign new_n359 = new_n332 & new_n358;
  assign new_n360 = new_n357 & new_n359;
  assign new_n361 = n1555 & new_n360;
  assign new_n362_1 = new_n355 & ~new_n361;
  assign new_n363_1 = ~n1389 & new_n317;
  assign new_n364_1 = ~new_n318 & ~new_n363_1;
  assign new_n365_1 = ~new_n362_1 & new_n364_1;
  assign new_n366 = new_n320 & new_n365_1;
  assign new_n367 = new_n322 & ~new_n366;
  assign new_n368_1 = new_n310 & ~new_n367;
  assign new_n369 = new_n306 & ~new_n367;
  assign new_n370 = ~new_n306 & ~new_n309;
  assign new_n371 = ~new_n310 & ~new_n370;
  assign new_n372 = ~new_n369 & new_n371;
  assign n693 = ~new_n368_1 & ~new_n372;
  assign new_n374 = new_n303 & n693;
  assign new_n375 = ~n532 & n1065;
  assign new_n376 = n664 & new_n375;
  assign new_n377 = ~n532 & ~n1065;
  assign new_n378 = n325 & n629;
  assign new_n379 = n507 & ~n629;
  assign new_n380 = ~new_n378 & ~new_n379;
  assign new_n381 = new_n377 & ~new_n380;
  assign new_n382 = ~new_n376 & ~new_n381;
  assign n1478 = new_n374 | ~new_n382;
  assign new_n384 = new_n302 & ~n1478;
  assign new_n385 = ~n1551 & n1655;
  assign new_n386_1 = n373 & n1243;
  assign new_n387 = n677 & ~n1243;
  assign new_n388_1 = ~new_n386_1 & ~new_n387;
  assign new_n389 = n1240 & ~new_n388_1;
  assign new_n390 = ~n1240 & new_n388_1;
  assign new_n391 = ~new_n389 & ~new_n390;
  assign new_n392 = n137 & n1243;
  assign new_n393 = n859 & ~n1243;
  assign new_n394 = ~new_n392 & ~new_n393;
  assign new_n395 = n184 & ~new_n394;
  assign new_n396 = ~n184 & new_n394;
  assign new_n397 = n1243 & n1331;
  assign new_n398 = n824 & ~n1243;
  assign new_n399 = ~new_n397 & ~new_n398;
  assign new_n400 = n1530 & ~new_n399;
  assign new_n401 = ~n1530 & new_n399;
  assign new_n402 = ~new_n400 & ~new_n401;
  assign new_n403_1 = n737 & n1243;
  assign new_n404 = n135 & ~n1243;
  assign new_n405 = ~new_n403_1 & ~new_n404;
  assign new_n406 = n765 & ~new_n405;
  assign new_n407 = new_n402 & new_n406;
  assign new_n408 = ~new_n400 & ~new_n407;
  assign new_n409 = ~new_n396 & ~new_n408;
  assign new_n410 = ~new_n395 & ~new_n409;
  assign new_n411 = ~new_n395 & ~new_n396;
  assign new_n412 = ~n765 & new_n405;
  assign new_n413 = new_n402 & ~new_n412;
  assign new_n414 = ~new_n406 & new_n413;
  assign new_n415_1 = new_n411 & new_n414;
  assign new_n416 = n579 & n1243;
  assign new_n417 = n1143 & ~n1243;
  assign new_n418_1 = ~new_n416 & ~new_n417;
  assign new_n419 = n1108 & ~new_n418_1;
  assign new_n420 = ~n1108 & new_n418_1;
  assign new_n421_1 = ~new_n419 & ~new_n420;
  assign new_n422 = n1243 & n1407;
  assign new_n423 = n956 & ~n1243;
  assign new_n424 = ~new_n422 & ~new_n423;
  assign new_n425 = ~n1479 & new_n424;
  assign new_n426 = n1479 & ~new_n424;
  assign new_n427_1 = n69 & n1243;
  assign new_n428 = ~n1243 & n1251;
  assign new_n429 = ~new_n427_1 & ~new_n428;
  assign new_n430 = ~n147 & new_n429;
  assign new_n431 = n147 & ~new_n429;
  assign new_n432_1 = n356 & n1243;
  assign new_n433 = n1030 & ~n1243;
  assign new_n434_1 = ~new_n432_1 & ~new_n433;
  assign new_n435 = ~n938 & new_n434_1;
  assign new_n436 = n938 & ~new_n434_1;
  assign new_n437 = n107 & n1243;
  assign new_n438 = n209 & ~n1243;
  assign new_n439 = ~new_n437 & ~new_n438;
  assign new_n440 = n950 & ~new_n439;
  assign new_n441 = ~new_n436 & ~new_n440;
  assign new_n442 = ~new_n435 & ~new_n441;
  assign new_n443 = ~new_n431 & ~new_n442;
  assign new_n444 = ~new_n430 & ~new_n443;
  assign new_n445 = ~new_n435 & ~new_n436;
  assign new_n446 = ~new_n430 & ~new_n431;
  assign new_n447 = new_n445 & new_n446;
  assign new_n448 = ~n950 & new_n439;
  assign new_n449 = ~new_n440 & ~new_n448;
  assign new_n450 = n857 & new_n449;
  assign new_n451 = new_n447 & new_n450;
  assign new_n452 = ~new_n444 & ~new_n451;
  assign new_n453 = ~new_n426 & new_n452;
  assign new_n454 = ~new_n425 & ~new_n453;
  assign new_n455 = new_n421_1 & new_n454;
  assign new_n456 = ~new_n419 & ~new_n455;
  assign new_n457 = new_n415_1 & ~new_n456;
  assign new_n458 = new_n410 & ~new_n457;
  assign new_n459 = new_n391 & new_n458;
  assign new_n460 = ~new_n391 & ~new_n458;
  assign new_n461 = ~new_n459 & ~new_n460;
  assign new_n462 = new_n303 & ~new_n461;
  assign new_n463 = n198 & n677;
  assign new_n464 = ~n677 & n1311;
  assign new_n465 = n1240 & ~new_n464;
  assign new_n466 = ~new_n463 & new_n465;
  assign new_n467 = ~n507 & ~n677;
  assign new_n468_1 = ~n325 & n677;
  assign new_n469 = ~new_n467 & ~new_n468_1;
  assign new_n470 = ~n1240 & new_n469;
  assign new_n471 = ~new_n466 & ~new_n470;
  assign new_n472 = new_n377 & ~new_n471;
  assign new_n473 = n1475 & new_n375;
  assign new_n474 = ~new_n472 & ~new_n473;
  assign n1645 = new_n462 | ~new_n474;
  assign new_n476_1 = new_n385 & ~n1645;
  assign new_n477 = n1551 & n1655;
  assign new_n478_1 = ~n526 & new_n477;
  assign new_n479 = n1551 & ~n1655;
  assign new_n480_1 = ~n362 & new_n479;
  assign new_n481_1 = ~new_n478_1 & ~new_n480_1;
  assign new_n482 = ~new_n476_1 & new_n481_1;
  assign n21 = new_n384 | ~new_n482;
  assign new_n484 = n84 & ~n726;
  assign new_n485 = ~new_n425 & ~new_n426;
  assign new_n486 = new_n452 & new_n485;
  assign new_n487 = ~new_n452 & ~new_n485;
  assign new_n488 = ~new_n486 & ~new_n487;
  assign new_n489_1 = new_n303 & ~new_n488;
  assign new_n490_1 = n751 & new_n375;
  assign new_n491 = ~n365 & ~n956;
  assign new_n492 = ~n230 & n956;
  assign new_n493 = n1479 & ~new_n492;
  assign new_n494 = ~new_n491 & new_n493;
  assign new_n495 = n956 & n1425;
  assign new_n496 = ~n956 & n1255;
  assign new_n497 = ~new_n495 & ~new_n496;
  assign new_n498 = ~n1479 & new_n497;
  assign new_n499 = ~new_n494 & ~new_n498;
  assign new_n500 = new_n377 & ~new_n499;
  assign new_n501 = ~new_n490_1 & ~new_n500;
  assign n928 = new_n489_1 | ~new_n501;
  assign new_n503 = new_n484 & ~n928;
  assign new_n504 = ~n84 & ~n726;
  assign new_n505 = ~n1555 & new_n332;
  assign new_n506_1 = ~new_n343 & new_n505;
  assign new_n507_1 = ~new_n350_1 & ~new_n506_1;
  assign new_n508 = ~new_n356_1 & new_n507_1;
  assign new_n509 = new_n356_1 & ~new_n507_1;
  assign new_n510 = ~new_n508 & ~new_n509;
  assign new_n511 = new_n303 & ~new_n510;
  assign new_n512 = n1189 & new_n375;
  assign new_n513 = n230 & n1545;
  assign new_n514_1 = ~n1425 & ~n1545;
  assign new_n515 = ~new_n513 & ~new_n514_1;
  assign new_n516 = new_n377 & ~new_n515;
  assign new_n517 = ~new_n512 & ~new_n516;
  assign n1157 = new_n511 | ~new_n517;
  assign new_n519 = new_n504 & ~n1157;
  assign new_n520 = ~n84 & n726;
  assign new_n521 = ~n468 & new_n520;
  assign new_n522 = n84 & n726;
  assign new_n523 = ~n934 & new_n522;
  assign new_n524_1 = ~new_n521 & ~new_n523;
  assign new_n525 = n1310 & new_n524_1;
  assign new_n526_1 = ~new_n519 & new_n525;
  assign n24 = new_n503 | ~new_n526_1;
  assign new_n528 = n901 & n1065;
  assign new_n529 = new_n421_1 & new_n440;
  assign new_n530 = ~new_n421_1 & ~new_n440;
  assign new_n531 = ~new_n529 & ~new_n530;
  assign new_n532_1 = ~new_n430 & new_n442;
  assign new_n533 = ~new_n443 & ~new_n532_1;
  assign new_n534 = new_n485 & new_n533;
  assign new_n535 = ~new_n485 & ~new_n533;
  assign new_n536 = ~new_n534 & ~new_n535;
  assign new_n537 = new_n531 & ~new_n536;
  assign new_n538 = ~new_n531 & new_n536;
  assign new_n539 = ~new_n537 & ~new_n538;
  assign new_n540 = ~new_n445 & ~new_n446;
  assign new_n541 = ~new_n447 & ~new_n540;
  assign new_n542 = ~new_n426 & ~new_n444;
  assign new_n543_1 = ~new_n425 & ~new_n542;
  assign new_n544 = new_n449 & new_n543_1;
  assign new_n545 = ~new_n449 & ~new_n543_1;
  assign new_n546 = ~new_n544 & ~new_n545;
  assign new_n547 = ~new_n541 & new_n546;
  assign new_n548 = new_n541 & ~new_n546;
  assign new_n549 = ~new_n547 & ~new_n548;
  assign new_n550 = ~new_n539 & ~new_n549;
  assign new_n551 = new_n539 & new_n549;
  assign new_n552 = ~n283 & ~new_n551;
  assign new_n553 = ~new_n550 & new_n552;
  assign new_n554 = new_n447 & new_n449;
  assign new_n555 = new_n485 & new_n554;
  assign new_n556 = new_n445 & new_n485;
  assign new_n557 = ~new_n445 & ~new_n485;
  assign new_n558 = ~new_n556 & ~new_n557;
  assign new_n559 = ~new_n555 & ~new_n558;
  assign new_n560 = new_n546 & ~new_n559;
  assign new_n561 = ~new_n546 & ~new_n558;
  assign new_n562 = ~new_n560 & ~new_n561;
  assign new_n563 = ~new_n436 & new_n448;
  assign new_n564 = ~new_n435 & ~new_n563;
  assign new_n565_1 = ~new_n421_1 & new_n446;
  assign new_n566 = new_n421_1 & ~new_n446;
  assign new_n567 = ~new_n565_1 & ~new_n566;
  assign new_n568 = new_n564 & new_n567;
  assign new_n569 = ~new_n564 & ~new_n567;
  assign new_n570 = ~new_n568 & ~new_n569;
  assign new_n571 = new_n444 & new_n448;
  assign new_n572 = ~new_n448 & ~new_n554;
  assign new_n573 = ~new_n444 & new_n572;
  assign new_n574_1 = ~new_n571 & ~new_n573;
  assign new_n575 = ~new_n570 & new_n574_1;
  assign new_n576_1 = new_n570 & ~new_n574_1;
  assign new_n577 = ~new_n575 & ~new_n576_1;
  assign new_n578 = ~new_n562 & new_n577;
  assign new_n579_1 = new_n562 & ~new_n577;
  assign new_n580 = ~new_n578 & ~new_n579_1;
  assign new_n581 = n283 & ~new_n580;
  assign new_n582 = ~new_n553 & ~new_n581;
  assign new_n583 = new_n421_1 & new_n555;
  assign new_n584 = n283 & new_n583;
  assign new_n585 = ~new_n419 & ~new_n543_1;
  assign new_n586 = ~new_n420 & ~new_n585;
  assign new_n587 = ~new_n584 & ~new_n586;
  assign new_n588_1 = new_n410 & ~new_n415_1;
  assign new_n589 = ~new_n402 & ~new_n406;
  assign new_n590 = ~new_n407 & ~new_n589;
  assign new_n591 = ~new_n400 & ~new_n413;
  assign new_n592 = new_n391 & new_n411;
  assign new_n593 = ~new_n391 & ~new_n411;
  assign new_n594 = ~new_n592 & ~new_n593;
  assign new_n595 = new_n591 & new_n594;
  assign new_n596_1 = ~new_n591 & ~new_n594;
  assign new_n597 = ~new_n595 & ~new_n596_1;
  assign new_n598_1 = ~new_n590 & new_n597;
  assign new_n599 = new_n590 & ~new_n597;
  assign new_n600 = ~new_n598_1 & ~new_n599;
  assign new_n601 = ~new_n588_1 & new_n600;
  assign new_n602 = new_n588_1 & ~new_n600;
  assign new_n603 = ~new_n601 & ~new_n602;
  assign new_n604 = ~new_n587 & ~new_n603;
  assign new_n605_1 = ~new_n395 & new_n408;
  assign new_n606 = ~new_n409 & ~new_n605_1;
  assign new_n607 = ~new_n402 & new_n412;
  assign new_n608_1 = ~new_n413 & ~new_n607;
  assign new_n609 = ~new_n594 & ~new_n608_1;
  assign new_n610 = new_n594 & new_n608_1;
  assign new_n611 = ~new_n609 & ~new_n610;
  assign new_n612 = new_n606 & new_n611;
  assign new_n613 = ~new_n606 & ~new_n611;
  assign new_n614_1 = ~new_n612 & ~new_n613;
  assign new_n615_1 = new_n587 & new_n614_1;
  assign new_n616 = ~new_n604 & ~new_n615_1;
  assign new_n617 = ~new_n582 & new_n616;
  assign new_n618_1 = new_n582 & ~new_n616;
  assign new_n619 = new_n303 & ~new_n618_1;
  assign new_n620 = ~new_n617 & new_n619;
  assign new_n621 = n198 & n1251;
  assign new_n622 = ~n1251 & n1311;
  assign new_n623_1 = n147 & ~new_n622;
  assign new_n624 = ~new_n621 & new_n623_1;
  assign new_n625 = ~n507 & ~n1251;
  assign new_n626 = ~n325 & n1251;
  assign new_n627 = ~new_n625 & ~new_n626;
  assign new_n628 = ~n147 & new_n627;
  assign new_n629_1 = ~new_n624 & ~new_n628;
  assign new_n630 = n198 & n824;
  assign new_n631 = ~n824 & n1311;
  assign new_n632 = n1530 & ~new_n631;
  assign new_n633_1 = ~new_n630 & new_n632;
  assign new_n634 = ~n507 & ~n824;
  assign new_n635_1 = ~n325 & n824;
  assign new_n636 = ~new_n634 & ~new_n635_1;
  assign new_n637 = ~n1530 & new_n636;
  assign new_n638 = ~new_n633_1 & ~new_n637;
  assign new_n639 = new_n629_1 & new_n638;
  assign new_n640_1 = ~new_n629_1 & ~new_n638;
  assign new_n641 = ~new_n639 & ~new_n640_1;
  assign new_n642 = n198 & n859;
  assign new_n643 = ~n859 & n1311;
  assign new_n644 = n184 & ~new_n643;
  assign new_n645 = ~new_n642 & new_n644;
  assign new_n646_1 = ~n507 & ~n859;
  assign new_n647 = ~n325 & n859;
  assign new_n648 = ~new_n646_1 & ~new_n647;
  assign new_n649 = ~n184 & new_n648;
  assign new_n650 = ~new_n645 & ~new_n649;
  assign new_n651 = n198 & n209;
  assign new_n652 = ~n209 & n1311;
  assign new_n653 = n950 & ~new_n652;
  assign new_n654_1 = ~new_n651 & new_n653;
  assign new_n655 = ~n209 & ~n507;
  assign new_n656_1 = n209 & ~n325;
  assign new_n657 = ~new_n655 & ~new_n656_1;
  assign new_n658 = ~n950 & new_n657;
  assign new_n659 = ~new_n654_1 & ~new_n658;
  assign new_n660 = new_n650 & new_n659;
  assign new_n661 = ~new_n650 & ~new_n659;
  assign new_n662 = ~new_n660 & ~new_n661;
  assign new_n663_1 = new_n641 & ~new_n662;
  assign new_n664_1 = ~new_n641 & new_n662;
  assign new_n665 = ~new_n663_1 & ~new_n664_1;
  assign new_n666 = n135 & n198;
  assign new_n667 = ~n135 & n1311;
  assign new_n668 = n765 & ~new_n667;
  assign new_n669 = ~new_n666 & new_n668;
  assign new_n670 = ~n135 & ~n507;
  assign new_n671 = n135 & ~n325;
  assign new_n672 = ~new_n670 & ~new_n671;
  assign new_n673 = ~n765 & new_n672;
  assign new_n674 = ~new_n669 & ~new_n673;
  assign new_n675_1 = new_n471 & new_n674;
  assign new_n676_1 = ~new_n471 & ~new_n674;
  assign new_n677_1 = ~new_n675_1 & ~new_n676_1;
  assign new_n678_1 = n198 & n1143;
  assign new_n679 = ~n1143 & n1311;
  assign new_n680 = n1108 & ~new_n679;
  assign new_n681 = ~new_n678_1 & new_n680;
  assign new_n682 = ~n507 & ~n1143;
  assign new_n683 = ~n325 & n1143;
  assign new_n684 = ~new_n682 & ~new_n683;
  assign new_n685 = ~n1108 & new_n684;
  assign new_n686 = ~new_n681 & ~new_n685;
  assign new_n687 = n198 & n956;
  assign new_n688 = ~n956 & n1311;
  assign new_n689 = n1479 & ~new_n688;
  assign new_n690 = ~new_n687 & new_n689;
  assign new_n691_1 = ~n507 & ~n956;
  assign new_n692 = ~n325 & n956;
  assign new_n693_1 = ~new_n691_1 & ~new_n692;
  assign new_n694 = ~n1479 & new_n693_1;
  assign new_n695 = ~new_n690 & ~new_n694;
  assign new_n696 = n198 & n1030;
  assign new_n697 = ~n1030 & n1311;
  assign new_n698 = n938 & ~new_n697;
  assign new_n699 = ~new_n696 & new_n698;
  assign new_n700 = ~n507 & ~n1030;
  assign new_n701 = ~n325 & n1030;
  assign new_n702 = ~new_n700 & ~new_n701;
  assign new_n703 = ~n938 & new_n702;
  assign new_n704_1 = ~new_n699 & ~new_n703;
  assign new_n705 = ~new_n695 & ~new_n704_1;
  assign new_n706 = new_n695 & new_n704_1;
  assign new_n707 = ~new_n705 & ~new_n706;
  assign new_n708 = new_n686 & new_n707;
  assign new_n709 = ~new_n686 & ~new_n707;
  assign new_n710_1 = ~new_n708 & ~new_n709;
  assign new_n711 = new_n677_1 & ~new_n710_1;
  assign new_n712 = ~new_n677_1 & new_n710_1;
  assign new_n713 = ~new_n711 & ~new_n712;
  assign new_n714 = new_n665 & new_n713;
  assign new_n715 = ~new_n665 & ~new_n713;
  assign new_n716_1 = new_n377 & ~new_n715;
  assign new_n717_1 = ~new_n714 & new_n716_1;
  assign new_n718 = ~new_n620 & ~new_n717_1;
  assign new_n719 = ~new_n528 & new_n718;
  assign new_n720 = n989 & ~n1413;
  assign new_n721 = ~new_n719 & new_n720;
  assign new_n722_1 = n989 & n1413;
  assign new_n723 = n1515 & new_n722_1;
  assign new_n724 = ~n989 & n1413;
  assign new_n725 = n1121 & new_n724;
  assign new_n726_1 = n837 & n1065;
  assign new_n727_1 = n198 & n654;
  assign new_n728 = ~n654 & n1311;
  assign new_n729 = n1389 & ~new_n728;
  assign new_n730 = ~new_n727_1 & new_n729;
  assign new_n731 = ~n507 & ~n654;
  assign new_n732 = ~n325 & n654;
  assign new_n733 = ~new_n731 & ~new_n732;
  assign new_n734 = ~n1389 & new_n733;
  assign new_n735 = ~new_n730 & ~new_n734;
  assign new_n736 = n198 & n1161;
  assign new_n737_1 = ~n1161 & n1311;
  assign new_n738 = ~new_n736 & ~new_n737_1;
  assign new_n739 = ~new_n735 & new_n738;
  assign new_n740_1 = new_n735 & ~new_n738;
  assign new_n741 = ~new_n739 & ~new_n740_1;
  assign new_n742 = n198 & n1518;
  assign new_n743 = n1311 & ~n1518;
  assign new_n744 = n769 & ~new_n743;
  assign new_n745 = ~new_n742 & new_n744;
  assign new_n746 = ~n507 & ~n1518;
  assign new_n747 = ~n325 & n1518;
  assign new_n748 = ~new_n746 & ~new_n747;
  assign new_n749 = ~n769 & new_n748;
  assign new_n750_1 = ~new_n745 & ~new_n749;
  assign new_n751_1 = n198 & n1335;
  assign new_n752 = n1311 & ~n1335;
  assign new_n753 = ~new_n751_1 & ~new_n752;
  assign new_n754 = ~new_n380 & new_n753;
  assign new_n755 = new_n380 & ~new_n753;
  assign new_n756 = ~new_n754 & ~new_n755;
  assign new_n757 = n198 & n490;
  assign new_n758 = ~n490 & n1311;
  assign new_n759 = n1165 & ~new_n758;
  assign new_n760 = ~new_n757 & new_n759;
  assign new_n761 = ~n490 & ~n507;
  assign new_n762 = ~n325 & n490;
  assign new_n763 = ~new_n761 & ~new_n762;
  assign new_n764 = ~n1165 & new_n763;
  assign new_n765_1 = ~new_n760 & ~new_n764;
  assign new_n766 = new_n756 & new_n765_1;
  assign new_n767 = ~new_n756 & ~new_n765_1;
  assign new_n768 = ~new_n766 & ~new_n767;
  assign new_n769_1 = new_n750_1 & new_n768;
  assign new_n770 = ~new_n750_1 & ~new_n768;
  assign new_n771 = ~new_n769_1 & ~new_n770;
  assign new_n772 = ~new_n741 & new_n771;
  assign new_n773 = new_n741 & ~new_n771;
  assign new_n774 = ~new_n772 & ~new_n773;
  assign new_n775 = n198 & n1058;
  assign new_n776 = ~n1058 & n1311;
  assign new_n777 = n403 & ~new_n776;
  assign new_n778 = ~new_n775 & new_n777;
  assign new_n779 = ~n507 & ~n1058;
  assign new_n780 = ~n325 & n1058;
  assign new_n781 = ~new_n779 & ~new_n780;
  assign new_n782 = ~n403 & new_n781;
  assign new_n783 = ~new_n778 & ~new_n782;
  assign new_n784 = n198 & n646;
  assign new_n785_1 = ~n646 & n1311;
  assign new_n786_1 = n1378 & ~new_n785_1;
  assign new_n787 = ~new_n784 & new_n786_1;
  assign new_n788 = ~n507 & ~n646;
  assign new_n789 = ~n325 & n646;
  assign new_n790_1 = ~new_n788 & ~new_n789;
  assign new_n791 = ~n1378 & new_n790_1;
  assign new_n792 = ~new_n787 & ~new_n791;
  assign new_n793_1 = n198 & n1545;
  assign new_n794_1 = ~n325 & ~n1545;
  assign new_n795 = ~new_n793_1 & ~new_n794_1;
  assign new_n796 = ~new_n792 & new_n795;
  assign new_n797_1 = new_n792 & ~new_n795;
  assign new_n798 = ~new_n796 & ~new_n797_1;
  assign new_n799 = new_n783 & ~new_n798;
  assign new_n800_1 = ~new_n783 & new_n798;
  assign new_n801 = ~new_n799 & ~new_n800_1;
  assign new_n802 = new_n774 & new_n801;
  assign new_n803 = ~new_n774 & ~new_n801;
  assign new_n804 = new_n377 & ~new_n803;
  assign new_n805 = ~new_n802 & new_n804;
  assign new_n806 = ~new_n347_1 & ~new_n348;
  assign new_n807 = ~new_n349 & ~new_n806;
  assign new_n808 = new_n332 & new_n807;
  assign new_n809 = ~new_n332 & ~new_n807;
  assign new_n810 = ~new_n808 & ~new_n809;
  assign new_n811 = new_n356_1 & new_n358;
  assign new_n812 = ~new_n356_1 & ~new_n358;
  assign new_n813 = ~new_n811 & ~new_n812;
  assign new_n814_1 = new_n332 & ~new_n340;
  assign new_n815 = ~new_n346 & ~new_n814_1;
  assign new_n816 = ~new_n813 & new_n815;
  assign new_n817 = new_n813 & ~new_n815;
  assign new_n818_1 = ~new_n816 & ~new_n817;
  assign new_n819 = ~new_n810 & new_n818_1;
  assign new_n820 = new_n810 & ~new_n818_1;
  assign new_n821_1 = ~new_n819 & ~new_n820;
  assign new_n822 = ~new_n332 & ~new_n350_1;
  assign new_n823 = ~new_n344 & ~new_n822;
  assign new_n824_1 = new_n353 & new_n823;
  assign new_n825 = ~new_n353 & ~new_n823;
  assign new_n826 = ~new_n824_1 & ~new_n825;
  assign new_n827 = ~new_n821_1 & new_n826;
  assign new_n828 = new_n821_1 & ~new_n826;
  assign new_n829_1 = ~new_n827 & ~new_n828;
  assign new_n830 = ~n1 & new_n829_1;
  assign new_n831 = ~new_n329 & new_n350_1;
  assign new_n832 = ~new_n351 & ~new_n831;
  assign new_n833 = ~new_n813 & new_n832;
  assign new_n834 = new_n813 & ~new_n832;
  assign new_n835_1 = ~new_n833 & ~new_n834;
  assign new_n836_1 = ~new_n346 & ~new_n810;
  assign new_n837_1 = new_n346 & new_n810;
  assign new_n838 = ~new_n836_1 & ~new_n837_1;
  assign new_n839 = ~new_n835_1 & ~new_n838;
  assign new_n840_1 = new_n835_1 & new_n838;
  assign new_n841 = ~new_n839 & ~new_n840_1;
  assign new_n842_1 = n1 & new_n841;
  assign new_n843 = ~new_n830 & ~new_n842_1;
  assign new_n844 = n1 & new_n360;
  assign new_n845_1 = new_n355 & ~new_n844;
  assign new_n846 = new_n306 & new_n319;
  assign new_n847 = new_n306 & ~new_n318;
  assign new_n848_1 = new_n320 & ~new_n847;
  assign new_n849 = ~new_n846 & ~new_n848_1;
  assign new_n850 = ~new_n371 & new_n849;
  assign new_n851_1 = new_n371 & ~new_n849;
  assign new_n852 = ~new_n850 & ~new_n851_1;
  assign new_n853 = new_n322 & new_n363_1;
  assign new_n854 = ~new_n322 & ~new_n363_1;
  assign new_n855 = ~new_n853 & ~new_n854;
  assign new_n856 = new_n852 & ~new_n855;
  assign new_n857_1 = ~new_n852 & new_n855;
  assign new_n858 = ~new_n856 & ~new_n857_1;
  assign new_n859_1 = new_n845_1 & ~new_n858;
  assign new_n860 = ~new_n318 & ~new_n320;
  assign new_n861 = ~new_n321 & ~new_n860;
  assign new_n862 = new_n320 & new_n364_1;
  assign new_n863 = ~new_n306 & new_n322;
  assign new_n864 = ~new_n862 & new_n863;
  assign new_n865 = new_n371 & ~new_n864;
  assign new_n866 = ~new_n309 & new_n864;
  assign new_n867 = ~new_n865 & ~new_n866;
  assign new_n868 = new_n861 & new_n867;
  assign new_n869_1 = ~new_n861 & ~new_n867;
  assign new_n870 = ~new_n868 & ~new_n869_1;
  assign new_n871 = ~new_n845_1 & ~new_n870;
  assign new_n872 = ~new_n859_1 & ~new_n871;
  assign new_n873 = new_n843 & new_n872;
  assign new_n874 = ~new_n843 & ~new_n872;
  assign new_n875 = new_n303 & ~new_n874;
  assign new_n876 = ~new_n873 & new_n875;
  assign new_n877_1 = ~new_n805 & ~new_n876;
  assign new_n878 = ~new_n726_1 & new_n877_1;
  assign new_n879 = ~n989 & ~n1413;
  assign new_n880 = ~new_n878 & new_n879;
  assign new_n881 = ~new_n725 & ~new_n880;
  assign new_n882 = ~new_n723 & new_n881;
  assign new_n883 = ~new_n721 & new_n882;
  assign n32 = n1310 & ~new_n883;
  assign new_n885 = ~new_n365_1 & new_n860;
  assign new_n886 = ~new_n321 & ~new_n885;
  assign new_n887_1 = ~new_n366 & new_n886;
  assign new_n888 = new_n347_1 & ~new_n887_1;
  assign new_n889 = n1555 & ~new_n332;
  assign new_n890 = ~new_n505 & ~new_n889;
  assign new_n891 = n1555 & new_n357;
  assign new_n892 = new_n353 & ~new_n891;
  assign new_n893 = ~new_n358 & new_n892;
  assign new_n894_1 = new_n358 & ~new_n892;
  assign new_n895 = ~new_n893 & ~new_n894_1;
  assign new_n896 = new_n890 & ~new_n895;
  assign new_n897 = new_n888 & new_n896;
  assign new_n898 = ~new_n306 & new_n367;
  assign new_n899 = ~new_n369 & ~new_n898;
  assign new_n900 = new_n362_1 & ~new_n364_1;
  assign new_n901_1 = ~new_n365_1 & ~new_n900;
  assign new_n902 = ~new_n340 & new_n505;
  assign new_n903 = ~new_n346 & ~new_n902;
  assign new_n904 = ~new_n348 & new_n903;
  assign new_n905 = new_n348 & ~new_n903;
  assign new_n906 = ~new_n904 & ~new_n905;
  assign new_n907 = ~new_n901_1 & new_n906;
  assign new_n908 = new_n510 & new_n907;
  assign new_n909_1 = ~new_n899 & new_n908;
  assign new_n910 = ~n693 & new_n909_1;
  assign n54 = ~new_n897 | ~new_n910;
  assign new_n912 = n182 & ~n877;
  assign new_n913 = new_n719 & new_n912;
  assign new_n914 = ~n182 & ~n877;
  assign new_n915 = new_n878 & new_n914;
  assign new_n916 = n182 & n877;
  assign new_n917 = ~n923 & new_n916;
  assign new_n918 = ~n182 & n877;
  assign new_n919 = ~n1280 & new_n918;
  assign new_n920 = ~new_n917 & ~new_n919;
  assign new_n921 = ~new_n915 & new_n920;
  assign n64 = new_n913 | ~new_n921;
  assign new_n923_1 = ~new_n440 & ~new_n450;
  assign new_n924 = new_n445 & ~new_n923_1;
  assign new_n925 = ~new_n436 & ~new_n924;
  assign new_n926 = ~new_n446 & new_n925;
  assign new_n927 = new_n446 & ~new_n925;
  assign new_n928_1 = ~new_n926 & ~new_n927;
  assign new_n929 = new_n303 & new_n928_1;
  assign new_n930 = n1418 & new_n375;
  assign new_n931 = ~n365 & ~n1251;
  assign new_n932 = ~n230 & n1251;
  assign new_n933_1 = n147 & ~new_n932;
  assign new_n934_1 = ~new_n931 & new_n933_1;
  assign new_n935 = n1251 & n1425;
  assign new_n936 = ~n1251 & n1255;
  assign new_n937 = ~new_n935 & ~new_n936;
  assign new_n938_1 = ~n147 & new_n937;
  assign new_n939 = ~new_n934_1 & ~new_n938_1;
  assign new_n940 = new_n377 & ~new_n939;
  assign new_n941 = ~new_n930 & ~new_n940;
  assign n1589 = new_n929 | ~new_n941;
  assign new_n943 = new_n484 & ~n1589;
  assign new_n944 = ~n909 & new_n520;
  assign new_n945 = ~n1511 & new_n522;
  assign new_n946 = n1310 & ~new_n945;
  assign new_n947 = ~new_n944 & new_n946;
  assign new_n948 = new_n303 & ~new_n906;
  assign new_n949 = n1049 & new_n375;
  assign new_n950_1 = ~n365 & ~n1518;
  assign new_n951 = ~n230 & n1518;
  assign new_n952 = n769 & ~new_n951;
  assign new_n953 = ~new_n950_1 & new_n952;
  assign new_n954 = n1425 & n1518;
  assign new_n955 = n1255 & ~n1518;
  assign new_n956_1 = ~new_n954 & ~new_n955;
  assign new_n957 = ~n769 & new_n956_1;
  assign new_n958 = ~new_n953 & ~new_n957;
  assign new_n959 = new_n377 & ~new_n958;
  assign new_n960 = ~new_n949 & ~new_n959;
  assign n1177 = new_n948 | ~new_n960;
  assign new_n962 = new_n504 & ~n1177;
  assign new_n963 = new_n947 & ~new_n962;
  assign n76 = new_n943 | ~new_n963;
  assign n167 = n421 & n1412;
  assign n83 = n415 & n167;
  assign new_n967 = new_n912 & ~n1589;
  assign new_n968 = new_n914 & ~n1177;
  assign new_n969 = ~n933 & new_n918;
  assign new_n970 = ~n1042 & new_n916;
  assign new_n971 = ~new_n969 & ~new_n970;
  assign new_n972 = ~new_n968 & new_n971;
  assign n97 = new_n967 | ~new_n972;
  assign new_n974_1 = new_n310 & new_n360;
  assign n110 = ~new_n862 | ~new_n974_1;
  assign new_n976 = ~n365 & ~n824;
  assign new_n977 = ~n230 & n824;
  assign new_n978 = n1530 & ~new_n977;
  assign new_n979 = ~new_n976 & new_n978;
  assign new_n980 = n824 & n1425;
  assign new_n981 = ~n824 & n1255;
  assign new_n982 = ~new_n980 & ~new_n981;
  assign new_n983 = ~n1530 & new_n982;
  assign new_n984 = ~new_n979 & ~new_n983;
  assign new_n985 = ~n365 & ~n859;
  assign new_n986 = ~n230 & n859;
  assign new_n987 = n184 & ~new_n986;
  assign new_n988 = ~new_n985 & new_n987;
  assign new_n989_1 = n859 & n1425;
  assign new_n990_1 = ~n859 & n1255;
  assign new_n991 = ~new_n989_1 & ~new_n990_1;
  assign new_n992 = ~n184 & new_n991;
  assign new_n993 = ~new_n988 & ~new_n992;
  assign new_n994 = ~n135 & ~n365;
  assign new_n995 = n135 & ~n230;
  assign new_n996 = n765 & ~new_n995;
  assign new_n997 = ~new_n994 & new_n996;
  assign new_n998 = n135 & n1425;
  assign new_n999 = ~n135 & n1255;
  assign new_n1000 = ~new_n998 & ~new_n999;
  assign new_n1001 = ~n765 & new_n1000;
  assign new_n1002 = ~new_n997 & ~new_n1001;
  assign new_n1003 = new_n993 & new_n1002;
  assign new_n1004 = ~n365 & ~n1030;
  assign new_n1005 = ~n230 & n1030;
  assign new_n1006 = n938 & ~new_n1005;
  assign new_n1007 = ~new_n1004 & new_n1006;
  assign new_n1008 = n1030 & n1425;
  assign new_n1009 = ~n1030 & n1255;
  assign new_n1010 = ~new_n1008 & ~new_n1009;
  assign new_n1011 = ~n938 & new_n1010;
  assign new_n1012 = ~new_n1007 & ~new_n1011;
  assign new_n1013_1 = new_n499 & new_n1012;
  assign new_n1014_1 = new_n1003 & new_n1013_1;
  assign new_n1015 = new_n471 & new_n939;
  assign new_n1016 = ~n209 & ~n365;
  assign new_n1017 = n209 & ~n230;
  assign new_n1018 = n950 & ~new_n1017;
  assign new_n1019_1 = ~new_n1016 & new_n1018;
  assign new_n1020 = n209 & n1425;
  assign new_n1021_1 = ~n209 & n1255;
  assign new_n1022 = ~new_n1020 & ~new_n1021_1;
  assign new_n1023_1 = ~n950 & new_n1022;
  assign new_n1024 = ~new_n1019_1 & ~new_n1023_1;
  assign new_n1025_1 = ~n365 & ~n1143;
  assign new_n1026_1 = ~n230 & n1143;
  assign new_n1027 = n1108 & ~new_n1026_1;
  assign new_n1028 = ~new_n1025_1 & new_n1027;
  assign new_n1029 = n1143 & n1425;
  assign new_n1030_1 = ~n1143 & n1255;
  assign new_n1031 = ~new_n1029 & ~new_n1030_1;
  assign new_n1032_1 = ~n1108 & new_n1031;
  assign new_n1033 = ~new_n1028 & ~new_n1032_1;
  assign new_n1034 = new_n1024 & new_n1033;
  assign new_n1035 = new_n1015 & new_n1034;
  assign new_n1036_1 = new_n1014_1 & new_n1035;
  assign n117 = ~new_n984 | ~new_n1036_1;
  assign new_n1038 = new_n414 & new_n592;
  assign n142 = ~new_n583 | ~new_n1038;
  assign new_n1040 = ~n1146 & new_n520;
  assign new_n1041 = ~n1398 & new_n522;
  assign new_n1042_1 = ~new_n1040 & ~new_n1041;
  assign new_n1043_1 = n1310 & new_n1042_1;
  assign new_n1044 = ~new_n406 & ~new_n412;
  assign new_n1045 = ~new_n456 & new_n1044;
  assign new_n1046 = new_n456 & ~new_n1044;
  assign new_n1047 = ~new_n1045 & ~new_n1046;
  assign new_n1048 = new_n303 & new_n1047;
  assign new_n1049_1 = n233 & new_n375;
  assign new_n1050 = new_n377 & ~new_n1002;
  assign new_n1051 = ~new_n1049_1 & ~new_n1050;
  assign n675 = new_n1048 | ~new_n1051;
  assign new_n1053 = new_n484 & ~n675;
  assign new_n1054 = new_n303 & new_n901_1;
  assign new_n1055 = new_n377 & ~new_n735;
  assign new_n1056 = n1580 & new_n375;
  assign new_n1057 = ~new_n1055 & ~new_n1056;
  assign n434 = new_n1054 | ~new_n1057;
  assign new_n1059 = new_n504 & ~n434;
  assign new_n1060 = ~new_n1053 & ~new_n1059;
  assign n150 = ~new_n1043_1 | ~new_n1060;
  assign new_n1062 = ~new_n445 & new_n923_1;
  assign new_n1063 = ~new_n924 & ~new_n1062;
  assign new_n1064 = new_n413 & ~new_n456;
  assign new_n1065_1 = new_n408 & ~new_n1064;
  assign new_n1066 = ~new_n411 & new_n1065_1;
  assign new_n1067 = new_n411 & ~new_n1065_1;
  assign new_n1068 = ~new_n1066 & ~new_n1067;
  assign new_n1069 = ~new_n1063 & ~new_n1068;
  assign new_n1070_1 = new_n589 & ~new_n1045;
  assign new_n1071 = ~new_n406 & new_n456;
  assign new_n1072 = new_n413 & ~new_n1071;
  assign new_n1073 = ~new_n1070_1 & ~new_n1072;
  assign new_n1074 = ~new_n421_1 & ~new_n454;
  assign new_n1075 = ~new_n455 & ~new_n1074;
  assign new_n1076 = ~new_n928_1 & ~new_n1075;
  assign new_n1077 = ~new_n1047 & new_n1076;
  assign new_n1078 = ~new_n1073 & new_n1077;
  assign new_n1079 = ~n857 & ~new_n449;
  assign new_n1080 = ~new_n450 & ~new_n1079;
  assign new_n1081 = new_n488 & ~new_n1080;
  assign new_n1082 = new_n461 & new_n1081;
  assign new_n1083 = new_n1078 & new_n1082;
  assign n170 = ~new_n1069 | ~new_n1083;
  assign new_n1085 = new_n484 & ~new_n719;
  assign new_n1086 = n1515 & new_n522;
  assign new_n1087 = n1121 & new_n520;
  assign new_n1088 = new_n504 & ~new_n878;
  assign new_n1089 = ~new_n1087 & ~new_n1088;
  assign new_n1090 = ~new_n1086 & new_n1089;
  assign new_n1091_1 = ~new_n1085 & new_n1090;
  assign n172 = n1310 & ~new_n1091_1;
  assign new_n1093_1 = ~n365 & ~n1058;
  assign new_n1094 = ~n230 & n1058;
  assign new_n1095 = n403 & ~new_n1094;
  assign new_n1096 = ~new_n1093_1 & new_n1095;
  assign new_n1097 = n1058 & n1425;
  assign new_n1098_1 = ~n1058 & n1255;
  assign new_n1099_1 = ~new_n1097 & ~new_n1098_1;
  assign new_n1100 = ~n403 & new_n1099_1;
  assign new_n1101 = ~new_n1096 & ~new_n1100;
  assign new_n1102 = new_n515 & new_n755;
  assign new_n1103 = new_n958 & new_n1102;
  assign new_n1104 = new_n1101 & new_n1103;
  assign new_n1105 = ~n365 & ~n646;
  assign new_n1106 = ~n230 & n646;
  assign new_n1107 = n1378 & ~new_n1106;
  assign new_n1108_1 = ~new_n1105 & new_n1107;
  assign new_n1109 = n646 & n1425;
  assign new_n1110 = ~n646 & n1255;
  assign new_n1111 = ~new_n1109 & ~new_n1110;
  assign new_n1112 = ~n1378 & new_n1111;
  assign new_n1113 = ~new_n1108_1 & ~new_n1112;
  assign new_n1114 = new_n765_1 & new_n1113;
  assign new_n1115 = new_n740_1 & new_n1114;
  assign n190 = ~new_n1104 | ~new_n1115;
  assign new_n1117_1 = ~n1478 & new_n914;
  assign new_n1118 = ~n1645 & new_n912;
  assign new_n1119 = ~n362 & new_n918;
  assign new_n1120 = ~n526 & new_n916;
  assign new_n1121_1 = ~new_n1119 & ~new_n1120;
  assign new_n1122_1 = ~new_n1118 & new_n1121_1;
  assign n204 = new_n1117_1 | ~new_n1122_1;
  assign new_n1124 = n635 & new_n375;
  assign new_n1125 = new_n377 & ~new_n1113;
  assign new_n1126 = ~new_n1124 & ~new_n1125;
  assign new_n1127 = ~new_n347_1 & new_n505;
  assign new_n1128 = new_n347_1 & ~new_n505;
  assign new_n1129 = new_n303 & ~new_n1128;
  assign new_n1130 = ~new_n1127 & new_n1129;
  assign n210 = ~new_n1126 | new_n1130;
  assign new_n1132 = ~n1014 & new_n916;
  assign new_n1133 = new_n303 & new_n895;
  assign new_n1134_1 = n1620 & new_n375;
  assign new_n1135 = new_n377 & ~new_n1101;
  assign new_n1136 = ~new_n1134_1 & ~new_n1135;
  assign n1665 = new_n1133 | ~new_n1136;
  assign new_n1138_1 = new_n914 & ~n1665;
  assign new_n1139 = ~new_n1132 & ~new_n1138_1;
  assign new_n1140 = ~n596 & new_n918;
  assign new_n1141 = new_n303 & new_n1075;
  assign new_n1142 = n432 & new_n375;
  assign new_n1143_1 = new_n377 & ~new_n1033;
  assign new_n1144 = ~new_n1142 & ~new_n1143_1;
  assign n1039 = new_n1141 | ~new_n1144;
  assign new_n1146_1 = new_n912 & ~n1039;
  assign new_n1147 = ~new_n1140 & ~new_n1146_1;
  assign n231 = ~new_n1139 | ~new_n1147;
  assign new_n1149 = ~new_n355 & new_n862;
  assign new_n1150_1 = new_n322 & ~new_n1149;
  assign n232 = new_n310 & new_n1150_1;
  assign new_n1152 = new_n303 & new_n887_1;
  assign new_n1153 = new_n377 & ~new_n765_1;
  assign new_n1154 = n1131 & new_n375;
  assign new_n1155 = ~new_n1153 & ~new_n1154;
  assign n640 = new_n1152 | ~new_n1155;
  assign new_n1157_1 = new_n504 & ~n640;
  assign new_n1158 = new_n303 & new_n1073;
  assign new_n1159 = new_n377 & ~new_n984;
  assign new_n1160_1 = n973 & new_n375;
  assign new_n1161_1 = ~new_n1159 & ~new_n1160_1;
  assign n964 = new_n1158 | ~new_n1161_1;
  assign new_n1163 = new_n484 & ~n964;
  assign new_n1164 = ~n289 & new_n520;
  assign new_n1165_1 = ~n1485 & new_n522;
  assign new_n1166 = ~new_n1164 & ~new_n1165_1;
  assign new_n1167 = n1310 & new_n1166;
  assign new_n1168 = ~new_n1163 & new_n1167;
  assign n240 = new_n1157_1 | ~new_n1168;
  assign n265 = ~n220 | n797;
  assign new_n1171 = ~n290 & new_n916;
  assign new_n1172 = new_n912 & ~n675;
  assign new_n1173 = ~new_n1171 & ~new_n1172;
  assign new_n1174 = ~n818 & new_n918;
  assign new_n1175 = new_n914 & ~n434;
  assign new_n1176 = ~new_n1174 & ~new_n1175;
  assign n269 = ~new_n1173 | ~new_n1176;
  assign new_n1178 = new_n303 & ~new_n890;
  assign new_n1179 = n716 & new_n375;
  assign new_n1180 = new_n377 & new_n738;
  assign new_n1181 = ~new_n1179 & ~new_n1180;
  assign n291 = new_n1178 | ~new_n1181;
  assign new_n1183 = ~n1146 & new_n724;
  assign new_n1184_1 = ~n1398 & new_n722_1;
  assign new_n1185 = ~new_n1183 & ~new_n1184_1;
  assign new_n1186 = n1310 & new_n1185;
  assign new_n1187_1 = new_n720 & ~n675;
  assign new_n1188 = new_n879 & ~n434;
  assign new_n1189_1 = ~new_n1187_1 & ~new_n1188;
  assign n313 = ~new_n1186 | ~new_n1189_1;
  assign new_n1191 = new_n303 & new_n1068;
  assign new_n1192_1 = n1508 & new_n375;
  assign new_n1193 = new_n377 & ~new_n993;
  assign new_n1194_1 = ~new_n1192_1 & ~new_n1193;
  assign n336 = new_n1191 | ~new_n1194_1;
  assign new_n1196 = ~n386 & new_n520;
  assign new_n1197 = ~n605 & new_n522;
  assign new_n1198_1 = ~new_n1196 & ~new_n1197;
  assign new_n1199 = n1310 & new_n1198_1;
  assign new_n1200 = new_n484 & ~n1039;
  assign new_n1201 = new_n504 & ~n1665;
  assign new_n1202 = ~new_n1200 & ~new_n1201;
  assign n347 = ~new_n1199 | ~new_n1202;
  assign new_n1204 = n1276 & n1396;
  assign new_n1205 = ~n835 & new_n309;
  assign new_n1206 = n835 & ~new_n309;
  assign new_n1207 = ~new_n1205 & ~new_n1206;
  assign new_n1208 = ~n120 & ~new_n1207;
  assign new_n1209 = n120 & n693;
  assign new_n1210 = n869 & ~new_n1209;
  assign new_n1211 = ~new_n1208 & new_n1210;
  assign new_n1212 = ~n120 & ~new_n380;
  assign new_n1213 = n120 & n664;
  assign new_n1214 = ~n869 & ~new_n1213;
  assign new_n1215 = ~new_n1212 & new_n1214;
  assign new_n1216 = ~new_n1211 & ~new_n1215;
  assign n363 = new_n1204 | ~new_n1216;
  assign new_n1218 = ~n693 & ~new_n1207;
  assign new_n1219 = n693 & new_n1207;
  assign n368 = ~new_n1218 & ~new_n1219;
  assign new_n1221 = ~n514 & n167;
  assign new_n1222 = n576 & new_n1221;
  assign new_n1223_1 = n514 & n167;
  assign new_n1224 = n1052 & new_n1223_1;
  assign n383 = new_n1222 | new_n1224;
  assign new_n1226 = new_n385 & ~n928;
  assign new_n1227 = new_n302 & ~n1157;
  assign new_n1228 = ~n9 & new_n479;
  assign new_n1229 = ~n1162 & new_n477;
  assign new_n1230 = ~new_n1228 & ~new_n1229;
  assign new_n1231 = ~new_n1227 & new_n1230;
  assign n427 = new_n1226 | ~new_n1231;
  assign new_n1233 = ~n386 & new_n724;
  assign new_n1234 = ~n605 & new_n722_1;
  assign new_n1235 = ~new_n1233 & ~new_n1234;
  assign new_n1236 = n1310 & new_n1235;
  assign new_n1237 = new_n720 & ~n1039;
  assign new_n1238 = new_n879 & ~n1665;
  assign new_n1239_1 = ~new_n1237 & ~new_n1238;
  assign n506 = ~new_n1236 | ~new_n1239_1;
  assign new_n1241 = ~n1478 & new_n504;
  assign new_n1242 = ~n1645 & new_n484;
  assign new_n1243_1 = ~n1091 & new_n522;
  assign new_n1244 = ~n418 & new_n520;
  assign new_n1245 = ~new_n1243_1 & ~new_n1244;
  assign new_n1246 = ~new_n1242 & new_n1245;
  assign new_n1247 = n1310 & new_n1246;
  assign n524 = new_n1241 | ~new_n1247;
  assign new_n1249 = new_n720 & ~n1589;
  assign new_n1250 = ~n909 & new_n724;
  assign new_n1251_1 = ~n1511 & new_n722_1;
  assign new_n1252 = n1310 & ~new_n1251_1;
  assign new_n1253_1 = ~new_n1250 & new_n1252;
  assign new_n1254 = new_n879 & ~n1177;
  assign new_n1255_1 = new_n1253_1 & ~new_n1254;
  assign n543 = new_n1249 | ~new_n1255_1;
  assign new_n1257 = ~n1366 & new_n375;
  assign n598 = ~new_n718 | new_n1257;
  assign new_n1259 = new_n410 & ~new_n586;
  assign new_n1260 = new_n391 & ~new_n588_1;
  assign new_n1261 = ~new_n1259 & new_n1260;
  assign n623 = ~new_n389 & ~new_n1261;
  assign new_n1263 = ~n596 & new_n479;
  assign new_n1264 = new_n385 & ~n1039;
  assign new_n1265 = ~new_n1263 & ~new_n1264;
  assign new_n1266 = ~n1014 & new_n477;
  assign new_n1267 = new_n302 & ~n1665;
  assign new_n1268 = ~new_n1266 & ~new_n1267;
  assign n633 = ~new_n1265 | ~new_n1268;
  assign new_n1270 = ~n1575 & ~n1606;
  assign new_n1271 = ~n588 & n1606;
  assign new_n1272 = ~new_n1270 & ~new_n1271;
  assign new_n1273 = ~new_n339 & new_n1272;
  assign new_n1274 = new_n339 & ~new_n1272;
  assign new_n1275_1 = ~new_n1273 & ~new_n1274;
  assign new_n1276_1 = new_n325_1 & ~new_n328;
  assign new_n1277 = n727 & new_n328;
  assign new_n1278 = ~new_n1276_1 & ~new_n1277;
  assign new_n1279 = new_n332 & new_n1278;
  assign new_n1280_1 = ~new_n332 & ~new_n1278;
  assign new_n1281 = ~new_n1279 & ~new_n1280_1;
  assign new_n1282 = new_n1275_1 & new_n1281;
  assign new_n1283 = ~new_n1275_1 & ~new_n1281;
  assign new_n1284 = ~new_n1282 & ~new_n1283;
  assign new_n1285 = new_n317 & new_n335;
  assign new_n1286 = ~new_n317 & ~new_n335;
  assign new_n1287 = ~new_n1285 & ~new_n1286;
  assign new_n1288 = new_n313_1 & ~new_n371;
  assign new_n1289 = ~new_n313_1 & new_n371;
  assign new_n1290 = ~new_n1288 & ~new_n1289;
  assign new_n1291 = ~new_n1287 & new_n1290;
  assign new_n1292 = new_n1287 & ~new_n1290;
  assign new_n1293 = ~new_n1291 & ~new_n1292;
  assign new_n1294 = ~new_n1284 & ~new_n1293;
  assign new_n1295 = new_n1284 & new_n1293;
  assign n656 = ~new_n1294 & ~new_n1295;
  assign new_n1297 = ~new_n399 & new_n405;
  assign new_n1298 = new_n399 & ~new_n405;
  assign new_n1299 = ~new_n1297 & ~new_n1298;
  assign new_n1300 = new_n388_1 & new_n394;
  assign new_n1301 = ~new_n388_1 & ~new_n394;
  assign new_n1302 = ~new_n1300 & ~new_n1301;
  assign new_n1303_1 = new_n1299 & ~new_n1302;
  assign new_n1304 = ~new_n1299 & new_n1302;
  assign new_n1305 = ~new_n1303_1 & ~new_n1304;
  assign new_n1306 = new_n429 & new_n1305;
  assign new_n1307 = ~new_n429 & ~new_n1305;
  assign new_n1308 = ~new_n1306 & ~new_n1307;
  assign new_n1309 = new_n418_1 & new_n434_1;
  assign new_n1310_1 = ~new_n418_1 & ~new_n434_1;
  assign new_n1311_1 = ~new_n1309 & ~new_n1310_1;
  assign new_n1312 = new_n439 & new_n1311_1;
  assign new_n1313 = ~new_n439 & ~new_n1311_1;
  assign new_n1314_1 = ~new_n1312 & ~new_n1313;
  assign new_n1315 = ~n268 & ~n1243;
  assign new_n1316 = n1243 & ~n1253;
  assign new_n1317 = ~new_n1315 & ~new_n1316;
  assign new_n1318 = ~new_n424 & new_n1317;
  assign new_n1319 = new_n424 & ~new_n1317;
  assign new_n1320 = ~new_n1318 & ~new_n1319;
  assign new_n1321 = new_n1314_1 & ~new_n1320;
  assign new_n1322 = ~new_n1314_1 & new_n1320;
  assign new_n1323 = ~new_n1321 & ~new_n1322;
  assign new_n1324 = ~new_n1308 & new_n1323;
  assign new_n1325 = new_n1308 & ~new_n1323;
  assign n676 = new_n1324 | new_n1325;
  assign new_n1327 = new_n303 & new_n1080;
  assign new_n1328 = n1339 & new_n375;
  assign new_n1329 = new_n377 & ~new_n1024;
  assign new_n1330 = ~new_n1328 & ~new_n1329;
  assign n1601 = new_n1327 | ~new_n1330;
  assign new_n1332 = new_n385 & ~n1601;
  assign new_n1333 = new_n302 & ~n291;
  assign new_n1334 = ~n1184 & new_n479;
  assign new_n1335_1 = ~n1361 & new_n477;
  assign new_n1336 = ~new_n1334 & ~new_n1335_1;
  assign new_n1337 = ~new_n1333 & new_n1336;
  assign n691 = new_n1332 | ~new_n1337;
  assign new_n1339_1 = new_n303 & new_n899;
  assign new_n1340 = new_n377 & new_n753;
  assign new_n1341 = n145 & new_n375;
  assign new_n1342 = ~new_n1340 & ~new_n1341;
  assign n722 = new_n1339_1 | ~new_n1342;
  assign new_n1344 = n1648 & new_n1221;
  assign new_n1345 = n1549 & new_n1223_1;
  assign n740 = new_n1344 | new_n1345;
  assign new_n1347 = ~n1143 & n1251;
  assign new_n1348 = n1143 & ~n1251;
  assign new_n1349 = ~new_n1347 & ~new_n1348;
  assign new_n1350 = n956 & n1030;
  assign new_n1351 = ~n956 & ~n1030;
  assign new_n1352 = ~new_n1350 & ~new_n1351;
  assign new_n1353 = new_n1349 & new_n1352;
  assign new_n1354 = ~new_n1349 & ~new_n1352;
  assign new_n1355 = ~new_n1353 & ~new_n1354;
  assign new_n1356 = ~n135 & n824;
  assign new_n1357 = n135 & ~n824;
  assign new_n1358 = ~new_n1356 & ~new_n1357;
  assign new_n1359 = new_n1355 & ~new_n1358;
  assign new_n1360 = ~new_n1355 & new_n1358;
  assign new_n1361_1 = ~new_n1359 & ~new_n1360;
  assign new_n1362 = n209 & n268;
  assign new_n1363 = ~n209 & ~n268;
  assign new_n1364 = ~new_n1362 & ~new_n1363;
  assign new_n1365 = n677 & n859;
  assign new_n1366_1 = ~n677 & ~n859;
  assign new_n1367 = ~new_n1365 & ~new_n1366_1;
  assign new_n1368 = new_n1364 & ~new_n1367;
  assign new_n1369 = ~new_n1364 & new_n1367;
  assign new_n1370 = ~new_n1368 & ~new_n1369;
  assign new_n1371 = ~new_n1361_1 & ~new_n1370;
  assign new_n1372 = new_n1361_1 & new_n1370;
  assign n785 = new_n1371 | new_n1372;
  assign n790 = ~n128 | ~n1562;
  assign new_n1375_1 = new_n303 & new_n1063;
  assign new_n1376 = n1303 & new_n375;
  assign new_n1377 = new_n377 & ~new_n1012;
  assign new_n1378_1 = ~new_n1376 & ~new_n1377;
  assign n887 = new_n1375_1 | ~new_n1378_1;
  assign new_n1380 = new_n385 & ~n887;
  assign new_n1381 = new_n302 & ~n210;
  assign new_n1382 = ~n793 & new_n479;
  assign new_n1383 = ~n1676 & new_n477;
  assign new_n1384 = ~new_n1382 & ~new_n1383;
  assign new_n1385 = ~new_n1381 & new_n1384;
  assign n814 = new_n1380 | ~new_n1385;
  assign new_n1387 = ~n222 & new_n375;
  assign n821 = ~new_n877_1 | new_n1387;
  assign new_n1389_1 = ~n1438 & new_n1223_1;
  assign new_n1390 = ~n704 & new_n1221;
  assign new_n1391 = n1150 & ~new_n1390;
  assign n836 = new_n1389_1 | ~new_n1391;
  assign new_n1393 = new_n504 & ~n722;
  assign new_n1394 = new_n484 & ~n336;
  assign new_n1395 = ~n851 & new_n522;
  assign new_n1396_1 = ~n615 & new_n520;
  assign new_n1397 = ~new_n1395 & ~new_n1396_1;
  assign new_n1398_1 = n1310 & new_n1397;
  assign new_n1399 = ~new_n1394 & new_n1398_1;
  assign n840 = new_n1393 | ~new_n1399;
  assign new_n1401 = new_n484 & ~n1601;
  assign new_n1402 = ~n710 & new_n520;
  assign new_n1403 = new_n504 & ~n291;
  assign new_n1404 = ~new_n1402 & ~new_n1403;
  assign new_n1405 = ~n1187 & new_n522;
  assign new_n1406 = n1310 & ~new_n1405;
  assign new_n1407_1 = new_n1404 & new_n1406;
  assign n894 = new_n1401 | ~new_n1407_1;
  assign new_n1409_1 = n676 & n785;
  assign n1032 = ~n293 | ~n750;
  assign new_n1411_1 = ~n1335 & n1575;
  assign new_n1412_1 = n1335 & ~n1575;
  assign new_n1413_1 = ~new_n1411_1 & ~new_n1412_1;
  assign new_n1414 = n629 & n1161;
  assign new_n1415 = ~n629 & ~n1161;
  assign new_n1416 = ~new_n1414 & ~new_n1415;
  assign new_n1417 = new_n1413_1 & new_n1416;
  assign new_n1418_1 = ~new_n1413_1 & ~new_n1416;
  assign new_n1419 = ~new_n1417 & ~new_n1418_1;
  assign new_n1420 = ~n1058 & ~n1518;
  assign new_n1421 = n1058 & n1518;
  assign new_n1422_1 = ~new_n1420 & ~new_n1421;
  assign new_n1423 = n490 & n646;
  assign new_n1424 = ~n490 & ~n646;
  assign new_n1425_1 = ~new_n1423 & ~new_n1424;
  assign new_n1426 = n654 & ~new_n1425_1;
  assign new_n1427 = ~n654 & new_n1425_1;
  assign new_n1428 = ~new_n1426 & ~new_n1427;
  assign new_n1429 = ~new_n1422_1 & new_n1428;
  assign new_n1430 = new_n1422_1 & ~new_n1428;
  assign new_n1431 = ~new_n1429 & ~new_n1430;
  assign new_n1432 = ~new_n1419 & ~new_n1431;
  assign new_n1433 = new_n1419 & new_n1431;
  assign n1411 = new_n1432 | new_n1433;
  assign n1631 = n296 & n1409;
  assign new_n1436 = n829 & n1631;
  assign new_n1437 = n1630 & new_n1436;
  assign new_n1438_1 = n1411 & new_n1437;
  assign new_n1439 = ~n1032 & new_n1438_1;
  assign new_n1440 = n656 & new_n1439;
  assign n1019 = ~new_n1409_1 | ~new_n1440;
  assign new_n1442_1 = ~n990 & new_n1223_1;
  assign new_n1443 = ~n330 & new_n1221;
  assign new_n1444 = n1150 & ~new_n1443;
  assign n1021 = new_n1442_1 | ~new_n1444;
  assign new_n1446 = new_n912 & ~n887;
  assign new_n1447 = new_n914 & ~n210;
  assign new_n1448 = ~n1676 & new_n916;
  assign new_n1449 = ~n793 & new_n918;
  assign new_n1450 = ~new_n1448 & ~new_n1449;
  assign new_n1451 = ~new_n1447 & new_n1450;
  assign n1036 = new_n1446 | ~new_n1451;
  assign new_n1453 = new_n720 & ~n1601;
  assign new_n1454_1 = ~n710 & new_n724;
  assign new_n1455 = new_n879 & ~n291;
  assign new_n1456 = ~new_n1454_1 & ~new_n1455;
  assign new_n1457 = ~n1187 & new_n722_1;
  assign new_n1458 = n1310 & ~new_n1457;
  assign new_n1459 = new_n1456 & new_n1458;
  assign n1043 = new_n1453 | ~new_n1459;
  assign new_n1461 = new_n912 & ~n1601;
  assign new_n1462 = new_n914 & ~n291;
  assign new_n1463 = ~n1361 & new_n916;
  assign new_n1464 = ~n1184 & new_n918;
  assign new_n1465 = ~new_n1463 & ~new_n1464;
  assign new_n1466 = ~new_n1462 & new_n1465;
  assign n1122 = new_n1461 | ~new_n1466;
  assign new_n1468 = new_n484 & ~n887;
  assign new_n1469 = ~n342 & new_n520;
  assign new_n1470 = new_n504 & ~n210;
  assign new_n1471 = ~new_n1469 & ~new_n1470;
  assign new_n1472 = ~n1093 & new_n522;
  assign new_n1473 = n1310 & ~new_n1472;
  assign new_n1474_1 = new_n1471 & new_n1473;
  assign n1138 = new_n1468 | ~new_n1474_1;
  assign new_n1476 = new_n302 & ~n722;
  assign new_n1477 = ~n67 & new_n479;
  assign new_n1478_1 = ~n1373 & new_n477;
  assign new_n1479_1 = new_n385 & ~n336;
  assign new_n1480 = ~new_n1478_1 & ~new_n1479_1;
  assign new_n1481 = ~new_n1477 & new_n1480;
  assign n1151 = new_n1476 | ~new_n1481;
  assign new_n1483 = new_n879 & ~n640;
  assign new_n1484 = new_n720 & ~n964;
  assign new_n1485_1 = ~n289 & new_n724;
  assign new_n1486 = ~n1485 & new_n722_1;
  assign new_n1487 = ~new_n1485_1 & ~new_n1486;
  assign new_n1488 = n1310 & new_n1487;
  assign new_n1489 = ~new_n1484 & new_n1488;
  assign n1160 = new_n1483 | ~new_n1489;
  assign new_n1491 = new_n720 & ~n887;
  assign new_n1492 = ~n342 & new_n724;
  assign new_n1493 = new_n879 & ~n210;
  assign new_n1494 = ~new_n1492 & ~new_n1493;
  assign new_n1495 = ~n1093 & new_n722_1;
  assign new_n1496 = n1310 & ~new_n1495;
  assign new_n1497 = new_n1494 & new_n1496;
  assign n1194 = new_n1491 | ~new_n1497;
  assign new_n1499 = new_n385 & ~n1589;
  assign new_n1500 = new_n302 & ~n1177;
  assign new_n1501 = ~n1042 & new_n477;
  assign new_n1502 = ~n933 & new_n479;
  assign new_n1503 = ~new_n1501 & ~new_n1502;
  assign new_n1504 = ~new_n1500 & new_n1503;
  assign n1198 = new_n1499 | ~new_n1504;
  assign new_n1506 = ~n1422 & new_n1223_1;
  assign new_n1507 = ~n1070 & new_n1221;
  assign new_n1508_1 = n1150 & ~new_n1507;
  assign n1239 = new_n1506 | ~new_n1508_1;
  assign new_n1510 = ~n818 & new_n479;
  assign new_n1511_1 = new_n302 & ~n434;
  assign new_n1512_1 = ~new_n1510 & ~new_n1511_1;
  assign new_n1513 = ~n290 & new_n477;
  assign new_n1514 = new_n385 & ~n675;
  assign new_n1515_1 = ~new_n1513 & ~new_n1514;
  assign n1275 = ~new_n1512_1 | ~new_n1515_1;
  assign new_n1517 = ~n928 & new_n912;
  assign new_n1518_1 = ~n1157 & new_n914;
  assign new_n1519 = ~n1162 & new_n916;
  assign new_n1520 = ~n9 & new_n918;
  assign new_n1521 = ~new_n1519 & ~new_n1520;
  assign new_n1522 = ~new_n1518_1 & new_n1521;
  assign n1314 = new_n1517 | ~new_n1522;
  assign new_n1524 = ~n928 & new_n720;
  assign new_n1525 = ~n1157 & new_n879;
  assign new_n1526 = ~n468 & new_n724;
  assign new_n1527 = ~n934 & new_n722_1;
  assign new_n1528 = ~new_n1526 & ~new_n1527;
  assign new_n1529 = n1310 & new_n1528;
  assign new_n1530_1 = ~new_n1525 & new_n1529;
  assign n1375 = new_n1524 | ~new_n1530_1;
  assign new_n1532 = new_n914 & ~n722;
  assign new_n1533 = ~n1373 & new_n916;
  assign new_n1534 = ~n67 & new_n918;
  assign new_n1535 = new_n912 & ~n336;
  assign new_n1536 = ~new_n1534 & ~new_n1535;
  assign new_n1537 = ~new_n1533 & new_n1536;
  assign n1392 = new_n1532 | ~new_n1537;
  assign n1454 = ~n1099 & n1412;
  assign new_n1540 = ~n1478 & new_n879;
  assign new_n1541 = ~n1645 & new_n720;
  assign new_n1542_1 = ~n1091 & new_n722_1;
  assign new_n1543 = ~n418 & new_n724;
  assign new_n1544 = ~new_n1542_1 & ~new_n1543;
  assign new_n1545_1 = ~new_n1541 & new_n1544;
  assign new_n1546 = n1310 & new_n1545_1;
  assign n1474 = new_n1540 | ~new_n1546;
  assign new_n1548 = new_n914 & ~n640;
  assign new_n1549_1 = new_n912 & ~n964;
  assign new_n1550 = ~n1581 & new_n916;
  assign new_n1551_1 = ~n848 & new_n918;
  assign new_n1552_1 = ~new_n1550 & ~new_n1551_1;
  assign new_n1553 = ~new_n1549_1 & new_n1552_1;
  assign n1512 = new_n1548 | ~new_n1553;
  assign new_n1555_1 = ~n974 & new_n1223_1;
  assign new_n1556_1 = ~n1098 & new_n1221;
  assign new_n1557 = n1150 & ~new_n1556_1;
  assign n1531 = new_n1555_1 | ~new_n1557;
  assign n1574 = ~n96 | ~n1150;
  assign new_n1560 = new_n385 & new_n719;
  assign new_n1561 = new_n302 & new_n878;
  assign new_n1562_1 = ~n1280 & new_n479;
  assign new_n1563 = ~n923 & new_n477;
  assign new_n1564 = ~new_n1562_1 & ~new_n1563;
  assign new_n1565 = ~new_n1561 & new_n1564;
  assign n1594 = new_n1560 | ~new_n1565;
  assign new_n1567 = new_n879 & ~n722;
  assign new_n1568 = new_n720 & ~n336;
  assign new_n1569 = ~n851 & new_n722_1;
  assign new_n1570 = ~n615 & new_n724;
  assign new_n1571 = ~new_n1569 & ~new_n1570;
  assign new_n1572 = n1310 & new_n1571;
  assign new_n1573 = ~new_n1568 & new_n1572;
  assign n1604 = new_n1567 | ~new_n1573;
  assign n1628 = n794 & n167;
  assign new_n1576 = new_n302 & ~n640;
  assign new_n1577 = new_n385 & ~n964;
  assign new_n1578 = ~n848 & new_n479;
  assign new_n1579 = ~n1581 & new_n477;
  assign new_n1580_1 = ~new_n1578 & ~new_n1579;
  assign new_n1581_1 = ~new_n1577 & new_n1580_1;
  assign n1671 = new_n1576 | ~new_n1581_1;
  assign n8 = ~n1150;
  assign n61 = ~n128;
  assign n292 = ~n1134;
  assign n565 = ~n842;
  assign n618 = ~n797;
  assign n800 = ~n629;
  assign n1629 = ~n1310;
  assign n154 = n478;
  assign n253 = n481;
  assign n324 = n293;
  assign n350 = n61;
  assign n364 = n842;
  assign n388 = n1013;
  assign n476 = n8;
  assign n480 = n232;
  assign n489 = n61;
  assign n608 = n1596;
  assign n614 = n142;
  assign n663 = n61;
  assign n678 = n623;
  assign n717 = n1134;
  assign n786 = n478;
  assign n845 = n61;
  assign n1023 = n1630;
  assign n1026 = n740;
  assign n1117 = n110;
  assign n1192 = n1134;
  assign n1442 = n574;
  assign n1542 = n750;
  assign n1547 = n565;
  assign n1552 = n478;
  assign n1556 = n829;
endmodule


