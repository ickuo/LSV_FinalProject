module top( n3 , n4 , n8 , n9 , n11 , n12 , n13 , n16 , n19 , 
n22 , n32 , n38 , n48 , n55 , n56 , n79 , n82 , n84 , n87 , 
n96 , n98 , n102 , n106 , n108 , n113 , n117 , n122 , n125 , n131 , 
n132 , n133 , n138 , n141 , n144 , n164 , n166 , n182 , n183 , n184 , 
n187 , n190 , n194 , n196 , n198 , n199 , n200 , n207 , n211 , n212 , 
n213 , n214 , n215 , n216 , n219 , n222 , n237 , n239 , n241 , n244 , 
n247 , n248 , n258 , n259 , n262 , n271 , n272 , n275 , n279 , n288 , 
n291 , n293 , n303 , n306 );
    input n8 , n12 , n13 , n16 , n19 , n32 , n38 , n48 , n55 , 
n79 , n82 , n102 , n106 , n108 , n113 , n117 , n122 , n132 , n138 , 
n141 , n164 , n166 , n182 , n183 , n184 , n187 , n198 , n200 , n212 , 
n213 , n214 , n219 , n237 , n241 , n244 , n247 , n248 , n271 , n272 , 
n291 , n293 ;
    output n3 , n4 , n9 , n11 , n22 , n56 , n84 , n87 , n96 , 
n98 , n125 , n131 , n133 , n144 , n190 , n194 , n196 , n199 , n207 , 
n211 , n215 , n216 , n222 , n239 , n258 , n259 , n262 , n275 , n279 , 
n288 , n303 , n306 ;
    wire n0 , n1 , n2 , n5 , n6 , n7 , n10 , n14 , n15 , 
n17 , n18 , n20 , n21 , n23 , n24 , n25 , n26 , n27 , n28 , 
n29 , n30 , n31 , n33 , n34 , n35 , n36 , n37 , n39 , n40 , 
n41 , n42 , n43 , n44 , n45 , n46 , n47 , n49 , n50 , n51 , 
n52 , n53 , n54 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , 
n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , 
n74 , n75 , n76 , n77 , n78 , n80 , n81 , n83 , n85 , n86 , 
n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n97 , n99 , 
n100 , n101 , n103 , n104 , n105 , n107 , n109 , n110 , n111 , n112 , 
n114 , n115 , n116 , n118 , n119 , n120 , n121 , n123 , n124 , n126 , 
n127 , n128 , n129 , n130 , n134 , n135 , n136 , n137 , n139 , n140 , 
n142 , n143 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , 
n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , 
n163 , n165 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , 
n175 , n176 , n177 , n178 , n179 , n180 , n181 , n185 , n186 , n188 , 
n189 , n191 , n192 , n193 , n195 , n197 , n201 , n202 , n203 , n204 , 
n205 , n206 , n208 , n209 , n210 , n217 , n218 , n220 , n221 , n223 , 
n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , 
n234 , n235 , n236 , n238 , n240 , n242 , n243 , n245 , n246 , n249 , 
n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n260 , n261 , 
n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n273 , n274 , 
n276 , n277 , n278 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , 
n287 , n289 , n290 , n292 , n294 , n295 , n296 , n297 , n298 , n299 , 
n300 , n301 , n302 , n304 , n305 ;
    not g0 ( n41 , n27 );
    not g1 ( n276 , n188 );
    not g2 ( n265 , n174 );
    not g3 ( n46 , n73 );
    xnor g4 ( n42 , n106 , n19 );
    not g5 ( n60 , n290 );
    xnor g6 ( n190 , n107 , n214 );
    not g7 ( n284 , n128 );
    xnor g8 ( n136 , n64 , n249 );
    xnor g9 ( n254 , n169 , n230 );
    xnor g10 ( n196 , n76 , n247 );
    xnor g11 ( n221 , n214 , n237 );
    or g12 ( n119 , n69 , n251 );
    xnor g13 ( n171 , n241 , n122 );
    xnor g14 ( n9 , n210 , n12 );
    not g15 ( n286 , n296 );
    xnor g16 ( n3 , n165 , n102 );
    or g17 ( n154 , n155 , n91 );
    not g18 ( n180 , n283 );
    not g19 ( n78 , n7 );
    xnor g20 ( n11 , n261 , n132 );
    or g21 ( n23 , n156 , n150 );
    not g22 ( n304 , n167 );
    or g23 ( n91 , n53 , n70 );
    xnor g24 ( n306 , n2 , n166 );
    xnor g25 ( n302 , n187 , n82 );
    or g26 ( n186 , n250 , n111 );
    not g27 ( n188 , n63 );
    nor g28 ( n159 , n272 , n204 );
    not g29 ( n292 , n192 );
    xnor g30 ( n176 , n138 , n247 );
    xnor g31 ( n245 , n249 , n85 );
    xnor g32 ( n234 , n301 , n209 );
    xnor g33 ( n259 , n225 , n122 );
    not g34 ( n218 , n94 );
    not g35 ( n66 , n294 );
    or g36 ( n139 , n74 , n31 );
    xnor g37 ( n118 , n241 , n271 );
    or g38 ( n120 , n24 , n180 );
    or g39 ( n261 , n156 , n186 );
    not g40 ( n130 , n246 );
    xnor g41 ( n275 , n30 , n198 );
    not g42 ( n167 , n97 );
    xnor g43 ( n112 , n129 , n101 );
    or g44 ( n195 , n146 , n298 );
    or g45 ( n142 , n157 , n287 );
    xnor g46 ( n169 , n183 , n291 );
    or g47 ( n127 , n24 , n130 );
    xnor g48 ( n297 , n132 , n19 );
    xnor g49 ( n99 , n189 , n263 );
    xnor g50 ( n273 , n297 , n50 );
    xnor g51 ( n285 , n16 , n166 );
    or g52 ( n172 , n134 , n90 );
    not g53 ( n270 , n224 );
    or g54 ( n149 , n143 , n217 );
    or g55 ( n135 , n157 , n277 );
    not g56 ( n223 , n44 );
    not g57 ( n65 , n61 );
    not g58 ( n228 , n277 );
    not g59 ( n157 , n33 );
    xnor g60 ( n131 , n274 , n241 );
    xnor g61 ( n258 , n154 , n244 );
    xnor g62 ( n128 , n273 , n43 );
    not g63 ( n266 , n304 );
    xnor g64 ( n222 , n137 , n237 );
    or g65 ( n274 , n286 , n150 );
    buf g66 ( n74 , n81 );
    not g67 ( n28 , n63 );
    and g68 ( n27 , n146 , n236 );
    or g69 ( n72 , n267 , n6 );
    or g70 ( n163 , n175 , n115 );
    not g71 ( n88 , n178 );
    not g72 ( n296 , n295 );
    xnor g73 ( n305 , n201 , n254 );
    not g74 ( n295 , n92 );
    not g75 ( n53 , n188 );
    or g76 ( n217 , n236 , n235 );
    xnor g77 ( n93 , n32 , n291 );
    not g78 ( n227 , n128 );
    xnor g79 ( n303 , n142 , n291 );
    xnor g80 ( n239 , n229 , n138 );
    xnor g81 ( n62 , n244 , n187 );
    not g82 ( n155 , n206 );
    xnor g83 ( n301 , n16 , n117 );
    or g84 ( n181 , n69 , n242 );
    xnor g85 ( n199 , n135 , n48 );
    not g86 ( n204 , n212 );
    not g87 ( n25 , n284 );
    not g88 ( n238 , n278 );
    not g89 ( n299 , n97 );
    and g90 ( n235 , n139 , n10 );
    not g91 ( n174 , n186 );
    xnor g92 ( n5 , n12 , n8 );
    xnor g93 ( n279 , n280 , n106 );
    or g94 ( n277 , n147 , n40 );
    nor g95 ( n83 , n182 , n17 );
    or g96 ( n30 , n53 , n90 );
    xnor g97 ( n240 , n243 , n15 );
    not g98 ( n168 , n278 );
    xnor g99 ( n68 , n54 , n62 );
    nor g100 ( n116 , n184 , n114 );
    or g101 ( n280 , n255 , n277 );
    or g102 ( n40 , n185 , n195 );
    xnor g103 ( n1 , n176 , n29 );
    or g104 ( n77 , n155 , n35 );
    xnor g105 ( n243 , n253 , n221 );
    or g106 ( n242 , n103 , n6 );
    or g107 ( n123 , n266 , n35 );
    or g108 ( n193 , n218 , n46 );
    xnor g109 ( n257 , n102 , n132 );
    or g110 ( n80 , n292 , n217 );
    or g111 ( n70 , n75 , n126 );
    xnor g112 ( n129 , n191 , n252 );
    xnor g113 ( n252 , n244 , n213 );
    xnor g114 ( n249 , n220 , n42 );
    buf g115 ( n185 , n240 );
    not g116 ( n18 , n295 );
    xnor g117 ( n211 , n23 , n271 );
    not g118 ( n246 , n289 );
    xnor g119 ( n209 , n198 , n183 );
    not g120 ( n147 , n282 );
    or g121 ( n59 , n203 , n6 );
    xnor g122 ( n153 , n285 , n257 );
    not g123 ( n283 , n71 );
    or g124 ( n229 , n168 , n289 );
    xnor g125 ( n84 , n160 , n200 );
    not g126 ( n205 , n20 );
    nor g127 ( n64 , n248 , n114 );
    or g128 ( n202 , n175 , n265 );
    xnor g129 ( n262 , n14 , n183 );
    buf g130 ( n233 , n92 );
    xnor g131 ( n22 , n202 , n16 );
    xnor g132 ( n85 , n152 , n254 );
    or g133 ( n35 , n233 , n181 );
    xnor g134 ( n109 , n159 , n129 );
    or g135 ( n158 , n233 , n86 );
    or g136 ( n111 , n185 , n47 );
    xnor g137 ( n260 , n153 , n99 );
    xnor g138 ( n4 , n151 , n108 );
    xnor g139 ( n15 , n263 , n305 );
    or g140 ( n71 , n74 , n158 );
    xnor g141 ( n92 , n67 , n112 );
    not g142 ( n236 , n299 );
    not g143 ( n17 , n212 );
    not g144 ( n287 , n205 );
    or g145 ( n107 , n223 , n91 );
    and g146 ( n6 , n45 , n26 );
    nor g147 ( n201 , n141 , n197 );
    xnor g148 ( n49 , n21 , n36 );
    not g149 ( n44 , n290 );
    or g150 ( n148 , n300 , n149 );
    not g151 ( n61 , n49 );
    not g152 ( n115 , n228 );
    not g153 ( n231 , n170 );
    not g154 ( n300 , n60 );
    and g155 ( n224 , n233 , n69 );
    and g156 ( n192 , n250 , n185 );
    or g157 ( n226 , n269 , n71 );
    not g158 ( n175 , n28 );
    or g159 ( n298 , n238 , n235 );
    xnor g160 ( n104 , n145 , n109 );
    xnor g161 ( n125 , n172 , n32 );
    xnor g162 ( n140 , n79 , n8 );
    xnor g163 ( n97 , n1 , n0 );
    xnor g164 ( n100 , n89 , n5 );
    not g165 ( n94 , n231 );
    not g166 ( n267 , n178 );
    not g167 ( n290 , n240 );
    not g168 ( n197 , n212 );
    or g169 ( n37 , n185 , n27 );
    not g170 ( n124 , n65 );
    not g171 ( n114 , n212 );
    or g172 ( n161 , n147 , n66 );
    not g173 ( n75 , n296 );
    buf g174 ( n146 , n105 );
    not g175 ( n24 , n94 );
    and g176 ( n251 , n74 , n203 );
    xnor g177 ( n96 , n127 , n79 );
    xnor g178 ( n264 , n83 , n100 );
    or g179 ( n137 , n223 , n46 );
    or g180 ( n47 , n41 , n235 );
    xnor g181 ( n215 , n232 , n38 );
    xnor g182 ( n216 , n161 , n213 );
    or g183 ( n160 , n78 , n289 );
    or g184 ( n150 , n250 , n148 );
    or g185 ( n173 , n270 , n59 );
    xnor g186 ( n144 , n179 , n219 );
    or g187 ( n232 , n88 , n20 );
    not g188 ( n203 , n227 );
    not g189 ( n282 , n231 );
    xnor g190 ( n208 , n213 , n82 );
    nor g191 ( n189 , n13 , n197 );
    xnor g192 ( n87 , n256 , n19 );
    not g193 ( n63 , n81 );
    xnor g194 ( n43 , n145 , n264 );
    not g195 ( n103 , n251 );
    not g196 ( n73 , n35 );
    xnor g197 ( n98 , n193 , n82 );
    or g198 ( n2 , n134 , n265 );
    not g199 ( n294 , n91 );
    xnor g200 ( n288 , n123 , n55 );
    not g201 ( n39 , n105 );
    xnor g202 ( n253 , n108 , n113 );
    nor g203 ( n58 , n164 , n204 );
    not g204 ( n134 , n65 );
    xnor g205 ( n170 , n34 , n245 );
    xnor g206 ( n50 , n271 , n38 );
    xnor g207 ( n36 , n100 , n281 );
    xnor g208 ( n29 , n219 , n55 );
    xnor g209 ( n67 , n52 , n171 );
    not g210 ( n143 , n7 );
    xnor g211 ( n34 , n140 , n208 );
    xnor g212 ( n162 , n108 , n138 );
    xnor g213 ( n81 , n234 , n104 );
    or g214 ( n76 , n266 , n180 );
    xnor g215 ( n207 , n77 , n187 );
    xnor g216 ( n263 , n177 , n118 );
    or g217 ( n51 , n97 , n192 );
    xnor g218 ( n281 , n116 , n95 );
    or g219 ( n26 , n250 , n37 );
    xnor g220 ( n110 , n200 , n79 );
    or g221 ( n289 , n74 , n173 );
    xnor g222 ( n52 , n102 , n106 );
    or g223 ( n45 , n146 , n51 );
    not g224 ( n269 , n60 );
    or g225 ( n225 , n255 , n20 );
    or g226 ( n151 , n269 , n130 );
    not g227 ( n121 , n150 );
    or g228 ( n165 , n286 , n186 );
    xnor g229 ( n21 , n268 , n93 );
    not g230 ( n156 , n25 );
    xnor g231 ( n101 , n58 , n95 );
    buf g232 ( n250 , n170 );
    xnor g233 ( n191 , n214 , n219 );
    xnor g234 ( n177 , n198 , n32 );
    xnor g235 ( n220 , n117 , n48 );
    or g236 ( n14 , n276 , n287 );
    not g237 ( n7 , n39 );
    xnor g238 ( n57 , n237 , n55 );
    xnor g239 ( n230 , n122 , n38 );
    or g240 ( n210 , n78 , n71 );
    not g241 ( n33 , n61 );
    not g242 ( n90 , n121 );
    xnor g243 ( n145 , n57 , n302 );
    or g244 ( n179 , n168 , n66 );
    nor g245 ( n152 , n293 , n17 );
    or g246 ( n10 , n233 , n119 );
    buf g247 ( n69 , n49 );
    not g248 ( n206 , n39 );
    xnor g249 ( n105 , n68 , n260 );
    or g250 ( n256 , n88 , n115 );
    not g251 ( n178 , n284 );
    or g252 ( n86 , n124 , n72 );
    not g253 ( n278 , n167 );
    xnor g254 ( n0 , n153 , n136 );
    xnor g255 ( n268 , n166 , n48 );
    or g256 ( n20 , n146 , n80 );
    xnor g257 ( n133 , n163 , n117 );
    not g258 ( n255 , n18 );
    xnor g259 ( n95 , n162 , n110 );
    xnor g260 ( n54 , n200 , n12 );
    xnor g261 ( n56 , n226 , n113 );
    xnor g262 ( n194 , n120 , n8 );
    or g263 ( n126 , n69 , n59 );
    xnor g264 ( n89 , n113 , n247 );
    or g265 ( n31 , n128 , n224 );
endmodule
