module top( n1 , n6 , n9 , n24 , n25 , n26 , n27 , n30 , n41 , 
n53 , n66 , n76 , n82 , n86 , n94 , n101 , n102 , n105 , n118 , 
n128 , n136 , n139 , n144 , n148 , n156 , n181 , n186 , n195 , n196 , 
n202 , n203 , n204 , n206 , n213 , n214 , n220 , n239 , n244 , n247 , 
n258 , n266 , n268 , n273 , n277 , n282 , n290 , n291 , n293 , n304 , 
n306 , n307 , n309 , n317 , n326 , n341 , n350 , n371 , n375 , n379 , 
n382 , n388 , n391 , n401 , n403 , n412 , n417 , n423 , n425 , n431 , 
n434 , n441 , n449 , n455 , n481 , n484 , n487 , n494 , n511 , n537 , 
n538 , n541 , n547 , n553 , n557 , n565 , n566 , n581 , n588 , n590 , 
n596 , n602 , n608 , n609 , n615 , n621 , n625 , n642 , n646 , n656 , 
n657 , n677 , n679 , n680 , n684 , n687 , n691 , n698 , n700 , n711 , 
n714 , n715 , n724 , n725 , n727 , n739 , n744 , n745 , n749 , n756 , 
n760 , n778 , n785 , n790 , n792 , n800 , n802 , n807 , n817 , n818 , 
n829 , n837 , n838 , n851 , n857 , n858 , n864 , n867 , n871 , n879 , 
n888 , n897 , n902 , n904 , n916 , n935 , n960 , n961 , n965 , n972 , 
n987 , n989 , n992 , n997 , n1009 , n1013 , n1015 , n1025 , n1039 , n1052 , 
n1057 , n1069 , n1076 , n1077 , n1082 , n1102 , n1125 , n1131 , n1132 , n1147 , 
n1150 , n1172 , n1176 , n1178 , n1194 , n1198 , n1212 , n1227 , n1234 , n1237 , 
n1245 , n1265 , n1267 , n1270 , n1277 , n1280 , n1284 , n1290 , n1295 , n1298 , 
n1305 , n1310 , n1313 , n1320 , n1329 , n1331 , n1335 , n1342 , n1345 , n1348 , 
n1349 , n1355 , n1358 , n1381 , n1386 , n1393 , n1400 , n1403 , n1404 , n1438 , 
n1445 , n1447 , n1449 , n1455 , n1458 , n1472 , n1473 , n1494 , n1504 , n1511 , 
n1515 , n1519 , n1524 , n1539 , n1541 , n1543 , n1558 , n1562 , n1574 , n1580 , 
n1581 , n1595 , n1598 , n1604 , n1605 , n1606 , n1612 , n1613 , n1616 , n1624 , 
n1630 , n1632 , n1639 , n1640 , n1641 , n1646 , n1650 , n1654 , n1655 , n1665 , 
n1666 , n1673 , n1674 , n1677 , n1682 , n1686 , n1688 , n1692 , n1693 , n1695 , 
n1697 , n1705 , n1708 , n1715 , n1719 , n1726 , n1734 , n1735 , n1739 , n1743 , 
n1756 , n1760 );
    input n1 , n66 , n86 , n94 , n118 , n195 , n202 , n204 , n213 , 
n244 , n247 , n306 , n309 , n371 , n375 , n382 , n388 , n403 , n412 , 
n417 , n423 , n425 , n481 , n484 , n487 , n494 , n511 , n547 , n557 , 
n621 , n625 , n656 , n657 , n677 , n680 , n684 , n687 , n725 , n744 , 
n745 , n749 , n807 , n818 , n829 , n857 , n864 , n871 , n897 , n902 , 
n916 , n935 , n960 , n961 , n989 , n997 , n1052 , n1132 , n1147 , n1172 , 
n1198 , n1234 , n1245 , n1265 , n1277 , n1280 , n1284 , n1290 , n1313 , n1320 , 
n1342 , n1345 , n1349 , n1386 , n1455 , n1473 , n1494 , n1562 , n1605 , n1612 , 
n1624 , n1640 , n1646 , n1665 , n1673 , n1682 , n1686 , n1692 , n1735 , n1743 ;
    output n6 , n9 , n24 , n25 , n26 , n27 , n30 , n41 , n53 , 
n76 , n82 , n101 , n102 , n105 , n128 , n136 , n139 , n144 , n148 , 
n156 , n181 , n186 , n196 , n203 , n206 , n214 , n220 , n239 , n258 , 
n266 , n268 , n273 , n277 , n282 , n290 , n291 , n293 , n304 , n307 , 
n317 , n326 , n341 , n350 , n379 , n391 , n401 , n431 , n434 , n441 , 
n449 , n455 , n537 , n538 , n541 , n553 , n565 , n566 , n581 , n588 , 
n590 , n596 , n602 , n608 , n609 , n615 , n642 , n646 , n679 , n691 , 
n698 , n700 , n711 , n714 , n715 , n724 , n727 , n739 , n756 , n760 , 
n778 , n785 , n790 , n792 , n800 , n802 , n817 , n837 , n838 , n851 , 
n858 , n867 , n879 , n888 , n904 , n965 , n972 , n987 , n992 , n1009 , 
n1013 , n1015 , n1025 , n1039 , n1057 , n1069 , n1076 , n1077 , n1082 , n1102 , 
n1125 , n1131 , n1150 , n1176 , n1178 , n1194 , n1212 , n1227 , n1237 , n1267 , 
n1270 , n1295 , n1298 , n1305 , n1310 , n1329 , n1331 , n1335 , n1348 , n1355 , 
n1358 , n1381 , n1393 , n1400 , n1403 , n1404 , n1438 , n1445 , n1447 , n1449 , 
n1458 , n1472 , n1504 , n1511 , n1515 , n1519 , n1524 , n1539 , n1541 , n1543 , 
n1558 , n1574 , n1580 , n1581 , n1595 , n1598 , n1604 , n1606 , n1613 , n1616 , 
n1630 , n1632 , n1639 , n1641 , n1650 , n1654 , n1655 , n1666 , n1674 , n1677 , 
n1688 , n1693 , n1695 , n1697 , n1705 , n1708 , n1715 , n1719 , n1726 , n1734 , 
n1739 , n1756 , n1760 ;
    wire n0 , n2 , n3 , n4 , n5 , n7 , n8 , n10 , n11 , 
n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , 
n22 , n23 , n28 , n29 , n31 , n32 , n33 , n34 , n35 , n36 , 
n37 , n38 , n39 , n40 , n42 , n43 , n44 , n45 , n46 , n47 , 
n48 , n49 , n50 , n51 , n52 , n54 , n55 , n56 , n57 , n58 , 
n59 , n60 , n61 , n62 , n63 , n64 , n65 , n67 , n68 , n69 , 
n70 , n71 , n72 , n73 , n74 , n75 , n77 , n78 , n79 , n80 , 
n81 , n83 , n84 , n85 , n87 , n88 , n89 , n90 , n91 , n92 , 
n93 , n95 , n96 , n97 , n98 , n99 , n100 , n103 , n104 , n106 , 
n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , 
n117 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , 
n129 , n130 , n131 , n132 , n133 , n134 , n135 , n137 , n138 , n140 , 
n141 , n142 , n143 , n145 , n146 , n147 , n149 , n150 , n151 , n152 , 
n153 , n154 , n155 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , 
n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , 
n174 , n175 , n176 , n177 , n178 , n179 , n180 , n182 , n183 , n184 , 
n185 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n197 , 
n198 , n199 , n200 , n201 , n205 , n207 , n208 , n209 , n210 , n211 , 
n212 , n215 , n216 , n217 , n218 , n219 , n221 , n222 , n223 , n224 , 
n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , 
n235 , n236 , n237 , n238 , n240 , n241 , n242 , n243 , n245 , n246 , 
n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , 
n259 , n260 , n261 , n262 , n263 , n264 , n265 , n267 , n269 , n270 , 
n271 , n272 , n274 , n275 , n276 , n278 , n279 , n280 , n281 , n283 , 
n284 , n285 , n286 , n287 , n288 , n289 , n292 , n294 , n295 , n296 , 
n297 , n298 , n299 , n300 , n301 , n302 , n303 , n305 , n308 , n310 , 
n311 , n312 , n313 , n314 , n315 , n316 , n318 , n319 , n320 , n321 , 
n322 , n323 , n324 , n325 , n327 , n328 , n329 , n330 , n331 , n332 , 
n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n342 , n343 , 
n344 , n345 , n346 , n347 , n348 , n349 , n351 , n352 , n353 , n354 , 
n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , 
n365 , n366 , n367 , n368 , n369 , n370 , n372 , n373 , n374 , n376 , 
n377 , n378 , n380 , n381 , n383 , n384 , n385 , n386 , n387 , n389 , 
n390 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , 
n402 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n413 , 
n414 , n415 , n416 , n418 , n419 , n420 , n421 , n422 , n424 , n426 , 
n427 , n428 , n429 , n430 , n432 , n433 , n435 , n436 , n437 , n438 , 
n439 , n440 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n450 , 
n451 , n452 , n453 , n454 , n456 , n457 , n458 , n459 , n460 , n461 , 
n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , 
n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n482 , 
n483 , n485 , n486 , n488 , n489 , n490 , n491 , n492 , n493 , n495 , 
n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , 
n506 , n507 , n508 , n509 , n510 , n512 , n513 , n514 , n515 , n516 , 
n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , 
n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , 
n539 , n540 , n542 , n543 , n544 , n545 , n546 , n548 , n549 , n550 , 
n551 , n552 , n554 , n555 , n556 , n558 , n559 , n560 , n561 , n562 , 
n563 , n564 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
n575 , n576 , n577 , n578 , n579 , n580 , n582 , n583 , n584 , n585 , 
n586 , n587 , n589 , n591 , n592 , n593 , n594 , n595 , n597 , n598 , 
n599 , n600 , n601 , n603 , n604 , n605 , n606 , n607 , n610 , n611 , 
n612 , n613 , n614 , n616 , n617 , n618 , n619 , n620 , n622 , n623 , 
n624 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , 
n635 , n636 , n637 , n638 , n639 , n640 , n641 , n643 , n644 , n645 , 
n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n658 , 
n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , 
n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n678 , n681 , 
n682 , n683 , n685 , n686 , n688 , n689 , n690 , n692 , n693 , n694 , 
n695 , n696 , n697 , n699 , n701 , n702 , n703 , n704 , n705 , n706 , 
n707 , n708 , n709 , n710 , n712 , n713 , n716 , n717 , n718 , n719 , 
n720 , n721 , n722 , n723 , n726 , n728 , n729 , n730 , n731 , n732 , 
n733 , n734 , n735 , n736 , n737 , n738 , n740 , n741 , n742 , n743 , 
n746 , n747 , n748 , n750 , n751 , n752 , n753 , n754 , n755 , n757 , 
n758 , n759 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , 
n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n779 , 
n780 , n781 , n782 , n783 , n784 , n786 , n787 , n788 , n789 , n791 , 
n793 , n794 , n795 , n796 , n797 , n798 , n799 , n801 , n803 , n804 , 
n805 , n806 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , 
n816 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , 
n828 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n839 , n840 , 
n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , 
n852 , n853 , n854 , n855 , n856 , n859 , n860 , n861 , n862 , n863 , 
n865 , n866 , n868 , n869 , n870 , n872 , n873 , n874 , n875 , n876 , 
n877 , n878 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , 
n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n898 , n899 , 
n900 , n901 , n903 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , 
n912 , n913 , n914 , n915 , n917 , n918 , n919 , n920 , n921 , n922 , 
n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , 
n933 , n934 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , 
n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , 
n954 , n955 , n956 , n957 , n958 , n959 , n962 , n963 , n964 , n966 , 
n967 , n968 , n969 , n970 , n971 , n973 , n974 , n975 , n976 , n977 , 
n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n988 , 
n990 , n991 , n993 , n994 , n995 , n996 , n998 , n999 , n1000 , n1001 , 
n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1010 , n1011 , n1012 , 
n1014 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , 
n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , 
n1036 , n1037 , n1038 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , 
n1047 , n1048 , n1049 , n1050 , n1051 , n1053 , n1054 , n1055 , n1056 , n1058 , 
n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , 
n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1078 , n1079 , n1080 , n1081 , 
n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , 
n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1103 , 
n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , 
n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , 
n1124 , n1126 , n1127 , n1128 , n1129 , n1130 , n1133 , n1134 , n1135 , n1136 , 
n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , 
n1148 , n1149 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , 
n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , 
n1169 , n1170 , n1171 , n1173 , n1174 , n1175 , n1177 , n1179 , n1180 , n1181 , 
n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , 
n1192 , n1193 , n1195 , n1196 , n1197 , n1199 , n1200 , n1201 , n1202 , n1203 , 
n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1213 , n1214 , 
n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , 
n1225 , n1226 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1235 , n1236 , 
n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1246 , n1247 , n1248 , 
n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , 
n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1266 , n1268 , n1269 , n1271 , 
n1272 , n1273 , n1274 , n1275 , n1276 , n1278 , n1279 , n1281 , n1282 , n1283 , 
n1285 , n1286 , n1287 , n1288 , n1289 , n1291 , n1292 , n1293 , n1294 , n1296 , 
n1297 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1306 , n1307 , n1308 , 
n1309 , n1311 , n1312 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1321 , 
n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1330 , n1332 , n1333 , 
n1334 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1343 , n1344 , n1346 , 
n1347 , n1350 , n1351 , n1352 , n1353 , n1354 , n1356 , n1357 , n1359 , n1360 , 
n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , 
n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , 
n1382 , n1383 , n1384 , n1385 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , 
n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1401 , n1402 , n1405 , n1406 , 
n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , 
n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , 
n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , 
n1437 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1446 , n1448 , n1450 , 
n1451 , n1452 , n1453 , n1454 , n1456 , n1457 , n1459 , n1460 , n1461 , n1462 , 
n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1474 , 
n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , 
n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1495 , 
n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1505 , n1506 , 
n1507 , n1508 , n1509 , n1510 , n1512 , n1513 , n1514 , n1516 , n1517 , n1518 , 
n1520 , n1521 , n1522 , n1523 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , 
n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1540 , n1542 , 
n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , 
n1554 , n1555 , n1556 , n1557 , n1559 , n1560 , n1561 , n1563 , n1564 , n1565 , 
n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1575 , n1576 , 
n1577 , n1578 , n1579 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , 
n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1596 , n1597 , n1599 , n1600 , 
n1601 , n1602 , n1603 , n1607 , n1608 , n1609 , n1610 , n1611 , n1614 , n1615 , 
n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1625 , n1626 , n1627 , 
n1628 , n1629 , n1631 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1642 , 
n1643 , n1644 , n1645 , n1647 , n1648 , n1649 , n1651 , n1652 , n1653 , n1656 , 
n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1667 , n1668 , 
n1669 , n1670 , n1671 , n1672 , n1675 , n1676 , n1678 , n1679 , n1680 , n1681 , 
n1683 , n1684 , n1685 , n1687 , n1689 , n1690 , n1691 , n1694 , n1696 , n1698 , 
n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1706 , n1707 , n1709 , n1710 , 
n1711 , n1712 , n1713 , n1714 , n1716 , n1717 , n1718 , n1720 , n1721 , n1722 , 
n1723 , n1724 , n1725 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , 
n1736 , n1737 , n1738 , n1740 , n1741 , n1742 , n1744 , n1745 , n1746 , n1747 , 
n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1757 , n1758 , 
n1759 , n1761 , n1762 , n1763 ;
    and g0 ( n501 , n585 , n789 );
    not g1 ( n1369 , n1640 );
    xnor g2 ( n331 , n1663 , n177 );
    or g3 ( n1544 , n299 , n1452 );
    xnor g4 ( n1697 , n1329 , n630 );
    and g5 ( n528 , n741 , n139 );
    nor g6 ( n1397 , n1673 , n184 );
    not g7 ( n1367 , n1172 );
    xnor g8 ( n770 , n444 , n306 );
    or g9 ( n1362 , n520 , n510 );
    xnor g10 ( n422 , n865 , n1514 );
    or g11 ( n1289 , n1211 , n1146 );
    not g12 ( n60 , n135 );
    and g13 ( n1224 , n643 , n979 );
    nor g14 ( n1597 , n1349 , n22 );
    or g15 ( n851 , n1296 , n943 );
    xor g16 ( n837 , n1539 , n528 );
    nor g17 ( n432 , n284 , n1733 );
    nor g18 ( n932 , n1409 , n1111 );
    xnor g19 ( n1543 , n1155 , n1419 );
    xnor g20 ( n265 , n1645 , n523 );
    not g21 ( n694 , n1202 );
    nor g22 ( n940 , n487 , n1349 );
    xnor g23 ( n9 , n1005 , n1423 );
    or g24 ( n814 , n1163 , n1402 );
    not g25 ( n978 , n512 );
    and g26 ( n1296 , n1505 , n1576 );
    xor g27 ( n933 , n1730 , n250 );
    and g28 ( n1196 , n1058 , n1436 );
    nor g29 ( n720 , n1577 , n799 );
    xnor g30 ( n463 , n916 , n1494 );
    and g31 ( n479 , n296 , n762 );
    xor g32 ( n1705 , n1307 , n59 );
    xnor g33 ( n1141 , n1234 , n1052 );
    or g34 ( n1467 , n1518 , n234 );
    xnor g35 ( n192 , n807 , n1052 );
    and g36 ( n2 , n251 , n187 );
    or g37 ( n1112 , n478 , n1089 );
    xnor g38 ( n1161 , n953 , n580 );
    and g39 ( n241 , n521 , n1537 );
    xnor g40 ( n889 , n460 , n902 );
    xnor g41 ( n596 , n252 , n945 );
    xor g42 ( n602 , n1258 , n1004 );
    and g43 ( n915 , n1192 , n322 );
    not g44 ( n828 , n177 );
    not g45 ( n217 , n44 );
    not g46 ( n40 , n1263 );
    nor g47 ( n732 , n1284 , n815 );
    nor g48 ( n1074 , n1121 , n1034 );
    not g49 ( n533 , n393 );
    xnor g50 ( n1595 , n1369 , n72 );
    and g51 ( n906 , n504 , n1019 );
    xnor g52 ( n1403 , n230 , n475 );
    or g53 ( n7 , n1474 , n1221 );
    not g54 ( n145 , n1468 );
    or g55 ( n394 , n354 , n1095 );
    or g56 ( n1649 , n1663 , n536 );
    buf g57 ( n144 , 1'b0 );
    xnor g58 ( n537 , n1190 , n1159 );
    xnor g59 ( n1613 , n466 , n773 );
    not g60 ( n755 , n309 );
    not g61 ( n1430 , n1562 );
    nor g62 ( n1599 , n801 , n907 );
    or g63 ( n976 , n366 , n351 );
    not g64 ( n99 , n1716 );
    xnor g65 ( n1302 , n1536 , n721 );
    not g66 ( n183 , n742 );
    and g67 ( n87 , n1052 , n382 );
    buf g68 ( n711 , 1'b0 );
    nor g69 ( n995 , n791 , n726 );
    and g70 ( n522 , n973 , n1044 );
    not g71 ( n1721 , n119 );
    not g72 ( n1325 , n748 );
    not g73 ( n223 , n133 );
    or g74 ( n1181 , n1520 , n21 );
    and g75 ( n1714 , n1052 , n1265 );
    not g76 ( n29 , n829 );
    and g77 ( n719 , n1395 , n1040 );
    xnor g78 ( n508 , n981 , n1763 );
    not g79 ( n299 , n1345 );
    not g80 ( n1308 , n1042 );
    not g81 ( n1561 , n145 );
    not g82 ( n1481 , n172 );
    not g83 ( n62 , n1475 );
    xnor g84 ( n1311 , n1745 , n1134 );
    xnor g85 ( n421 , n358 , n1614 );
    not g86 ( n1167 , n480 );
    not g87 ( n57 , n1346 );
    and g88 ( n478 , n1349 , n897 );
    xnor g89 ( n475 , n264 , n352 );
    and g90 ( n1095 , n1287 , n985 );
    and g91 ( n984 , n563 , n783 );
    not g92 ( n1529 , n994 );
    and g93 ( n855 , n1081 , n1667 );
    buf g94 ( n879 , 1'b0 );
    not g95 ( n1191 , n1134 );
    not g96 ( n284 , n66 );
    and g97 ( n1089 , n869 , n218 );
    or g98 ( n610 , n1003 , n1037 );
    nor g99 ( n1332 , n452 , n439 );
    xnor g100 ( n673 , n1725 , n1365 );
    not g101 ( n899 , n643 );
    xnor g102 ( n25 , n1196 , n954 );
    nor g103 ( n998 , n1074 , n69 );
    and g104 ( n1327 , n862 , n539 );
    xnor g105 ( n59 , n1589 , n914 );
    not g106 ( n1244 , n592 );
    xnor g107 ( n386 , n1414 , n1313 );
    xnor g108 ( n220 , n1633 , n1169 );
    not g109 ( n28 , n1755 );
    not g110 ( n942 , n768 );
    xnor g111 ( n778 , n1304 , n1178 );
    xnor g112 ( n731 , n1290 , n1349 );
    not g113 ( n527 , n17 );
    or g114 ( n1491 , n1091 , n1139 );
    xnor g115 ( n1039 , n951 , n699 );
    not g116 ( n177 , n536 );
    xor g117 ( n1387 , n298 , n1308 );
    xnor g118 ( n1598 , n1103 , n886 );
    and g119 ( n1601 , n167 , n948 );
    and g120 ( n704 , n1735 , n1284 );
    or g121 ( n1710 , n1367 , n969 );
    not g122 ( n706 , n216 );
    not g123 ( n442 , n1653 );
    not g124 ( n68 , n522 );
    nor g125 ( n1406 , n657 , n1501 );
    xnor g126 ( n1695 , n1736 , n1005 );
    not g127 ( n160 , n1071 );
    or g128 ( n287 , n1553 , n1163 );
    xnor g129 ( n130 , n382 , n1052 );
    and g130 ( n127 , n405 , n483 );
    nor g131 ( n1620 , n749 , n312 );
    or g132 ( n407 , n324 , n1525 );
    and g133 ( n110 , n1551 , n644 );
    or g134 ( n655 , n952 , n629 );
    or g135 ( n222 , n1134 , n957 );
    not g136 ( n1645 , n236 );
    xnor g137 ( n214 , n1287 , n1311 );
    and g138 ( n832 , n1433 , n335 );
    not g139 ( n924 , n205 );
    or g140 ( n1346 , n829 , n1564 );
    or g141 ( n458 , n592 , n964 );
    xnor g142 ( n702 , n1692 , n1494 );
    not g143 ( n911 , n1522 );
    and g144 ( n1538 , n868 , n1735 );
    or g145 ( n733 , n1427 , n1196 );
    and g146 ( n516 , n910 , n314 );
    and g147 ( n1038 , n164 , n824 );
    not g148 ( n672 , n1575 );
    xnor g149 ( n660 , n1188 , n933 );
    and g150 ( n380 , n12 , n705 );
    nor g151 ( n1351 , n766 , n710 );
    nor g152 ( n506 , n644 , n1670 );
    and g153 ( n1051 , n1263 , n68 );
    not g154 ( n667 , n104 );
    or g155 ( n95 , n1110 , n772 );
    nor g156 ( n55 , n518 , n1008 );
    xnor g157 ( n954 , n32 , n1621 );
    not g158 ( n1722 , n1682 );
    not g159 ( n569 , n453 );
    xnor g160 ( n1363 , n1173 , n1208 );
    and g161 ( n325 , n1261 , n1255 );
    or g162 ( n1546 , n949 , n91 );
    xnor g163 ( n461 , n1645 , n1407 );
    xnor g164 ( n216 , n179 , n1326 );
    not g165 ( n1681 , n11 );
    xnor g166 ( n431 , n1162 , n275 );
    not g167 ( n437 , n652 );
    not g168 ( n349 , n1536 );
    not g169 ( n641 , n779 );
    not g170 ( n734 , n557 );
    or g171 ( n647 , n1675 , n428 );
    or g172 ( n579 , n1375 , n861 );
    not g173 ( n1309 , n343 );
    not g174 ( n473 , n1432 );
    or g175 ( n339 , n876 , n496 );
    xnor g176 ( n1209 , n1455 , n1052 );
    and g177 ( n966 , n986 , n243 );
    not g178 ( n147 , n1433 );
    or g179 ( n1328 , n831 , n779 );
    nor g180 ( n1628 , n661 , n1142 );
    nor g181 ( n1482 , n657 , n201 );
    nor g182 ( n1413 , n334 , n1251 );
    not g183 ( n77 , n440 );
    or g184 ( n1587 , n1173 , n830 );
    and g185 ( n1516 , n1167 , n1748 );
    nor g186 ( n825 , n745 , n1245 );
    not g187 ( n20 , n1228 );
    or g188 ( n929 , n378 , n855 );
    and g189 ( n1159 , n874 , n241 );
    xnor g190 ( n1739 , n1618 , n256 );
    not g191 ( n658 , n360 );
    nor g192 ( n359 , n408 , n1622 );
    not g193 ( n294 , n383 );
    xnor g194 ( n793 , n1724 , n1064 );
    xnor g195 ( n1391 , n925 , n1245 );
    and g196 ( n1200 , n210 , n631 );
    not g197 ( n303 , n1508 );
    xor g198 ( n1693 , n60 , n289 );
    xnor g199 ( n773 , n592 , n1003 );
    not g200 ( n593 , n1147 );
    or g201 ( n550 , n483 , n717 );
    xnor g202 ( n1511 , n1712 , n1216 );
    and g203 ( n1317 , n929 , n1301 );
    or g204 ( n1385 , n786 , n1406 );
    and g205 ( n104 , n60 , n289 );
    and g206 ( n1408 , n981 , n47 );
    not g207 ( n1486 , n883 );
    xnor g208 ( n524 , n1112 , n1209 );
    or g209 ( n612 , n1203 , n355 );
    or g210 ( n1276 , n1607 , n474 );
    and g211 ( n1243 , n1245 , n1277 );
    and g212 ( n558 , n584 , n1587 );
    or g213 ( n662 , n1290 , n1349 );
    not g214 ( n881 , n1640 );
    and g215 ( n1020 , n112 , n924 );
    or g216 ( n1168 , n219 , n881 );
    not g217 ( n1356 , n1685 );
    or g218 ( n488 , n1659 , n468 );
    and g219 ( n368 , n706 , n103 );
    nor g220 ( n696 , n1024 , n713 );
    xnor g221 ( n159 , n453 , n247 );
    or g222 ( n1738 , n363 , n1452 );
    not g223 ( n854 , n1114 );
    and g224 ( n100 , n1282 , n98 );
    not g225 ( n64 , n644 );
    xnor g226 ( n1581 , n251 , n320 );
    and g227 ( n1183 , n1068 , n1509 );
    not g228 ( n1745 , n1079 );
    xnor g229 ( n1305 , n365 , n939 );
    or g230 ( n1399 , n428 , n804 );
    not g231 ( n816 , n636 );
    xnor g232 ( n1329 , n387 , n923 );
    nor g233 ( n1373 , n435 , n146 );
    and g234 ( n1563 , n1660 , n1710 );
    or g235 ( n535 , n1324 , n106 );
    not g236 ( n88 , n232 );
    or g237 ( n1501 , n1195 , n29 );
    not g238 ( n639 , n944 );
    and g239 ( n278 , n301 , n152 );
    not g240 ( n1297 , n236 );
    or g241 ( n1321 , n638 , n854 );
    and g242 ( n242 , n1207 , n971 );
    not g243 ( n1017 , n1246 );
    not g244 ( n363 , n487 );
    xnor g245 ( n1674 , n562 , n1761 );
    and g246 ( n936 , n1252 , n678 );
    nor g247 ( n211 , n1409 , n637 );
    and g248 ( n1258 , n827 , n1281 );
    xnor g249 ( n1125 , n1317 , n1582 );
    xnor g250 ( n1515 , n607 , n79 );
    or g251 ( n490 , n524 , n172 );
    xor g252 ( n105 , n767 , n1629 );
    or g253 ( n708 , n1056 , n895 );
    or g254 ( n1184 , n1332 , n383 );
    and g255 ( n1622 , n958 , n1544 );
    or g256 ( n1392 , n1078 , n1151 );
    not g257 ( n748 , n107 );
    xnor g258 ( n588 , n1014 , n842 );
    not g259 ( n281 , n1492 );
    or g260 ( n1699 , n735 , n1568 );
    nor g261 ( n1417 , n1702 , n575 );
    and g262 ( n1569 , n1467 , n1174 );
    or g263 ( n817 , n1504 , n1036 );
    or g264 ( n1436 , n311 , n1328 );
    and g265 ( n1402 , n1215 , n140 );
    xnor g266 ( n435 , n433 , n481 );
    not g267 ( n880 , n1347 );
    nor g268 ( n409 , n1188 , n595 );
    not g269 ( n1754 , n1466 );
    or g270 ( n1711 , n198 , n1718 );
    and g271 ( n852 , n20 , n1318 );
    not g272 ( n730 , n259 );
    or g273 ( n1101 , n116 , n1643 );
    nor g274 ( n874 , n52 , n1353 );
    not g275 ( n1120 , n1241 );
    nor g276 ( n1288 , n1502 , n893 );
    not g277 ( n1670 , n887 );
    not g278 ( n729 , n899 );
    not g279 ( n1553 , n1052 );
    or g280 ( n1434 , n1223 , n1177 );
    or g281 ( n1058 , n240 , n472 );
    or g282 ( n1700 , n426 , n1553 );
    or g283 ( n1458 , n1225 , n471 );
    xnor g284 ( n1003 , n1321 , n1352 );
    and g285 ( n1100 , n908 , n125 );
    not g286 ( n11 , n1279 );
    or g287 ( n882 , n1652 , n1601 );
    not g288 ( n1414 , n644 );
    or g289 ( n973 , n1054 , n1625 );
    nor g290 ( n366 , n1494 , n1488 );
    and g291 ( n1225 , n1015 , n573 );
    not g292 ( n905 , n605 );
    and g293 ( n1720 , n701 , n684 );
    not g294 ( n1464 , n1444 );
    xor g295 ( n30 , n1421 , n434 );
    or g296 ( n199 , n678 , n836 );
    or g297 ( n1044 , n1147 , n71 );
    or g298 ( n323 , n561 , n1093 );
    or g299 ( n404 , n1256 , n938 );
    nor g300 ( n1750 , n1113 , n1273 );
    not g301 ( n8 , n857 );
    nor g302 ( n474 , n109 , n398 );
    or g303 ( n1760 , n1327 , n1117 );
    and g304 ( n1729 , n525 , n616 );
    or g305 ( n493 , n940 , n358 );
    and g306 ( n772 , n976 , n1480 );
    or g307 ( n1725 , n821 , n720 );
    and g308 ( n1086 , n1273 , n352 );
    nor g309 ( n1210 , n1195 , n803 );
    or g310 ( n1326 , n835 , n670 );
    xnor g311 ( n441 , n1190 , n559 );
    not g312 ( n666 , n826 );
    not g313 ( n1653 , n1226 );
    xnor g314 ( n741 , n351 , n151 );
    not g315 ( n1330 , n1061 );
    not g316 ( n1178 , n1382 );
    xnor g317 ( n894 , n1689 , n655 );
    and g318 ( n1600 , n377 , n1269 );
    and g319 ( n949 , n978 , n730 );
    or g320 ( n630 , n1469 , n1464 );
    or g321 ( n1030 , n1092 , n577 );
    not g322 ( n809 , n1701 );
    or g323 ( n1708 , n955 , n559 );
    xnor g324 ( n727 , n1736 , n779 );
    not g325 ( n898 , n438 );
    buf g326 ( n1740 , n693 );
    not g327 ( n385 , n78 );
    and g328 ( n44 , n1540 , n1346 );
    or g329 ( n1073 , n425 , n1245 );
    or g330 ( n751 , n189 , n160 );
    or g331 ( n1246 , n120 , n628 );
    not g332 ( n1576 , n1011 );
    xnor g333 ( n74 , n86 , n1494 );
    xnor g334 ( n790 , n325 , n0 );
    not g335 ( n834 , n605 );
    and g336 ( n492 , n1717 , n46 );
    not g337 ( n1442 , n933 );
    not g338 ( n1488 , n1144 );
    xnor g339 ( n1517 , n165 , n396 );
    or g340 ( n838 , n761 , n1746 );
    not g341 ( n1609 , n259 );
    or g342 ( n914 , n1156 , n433 );
    nor g343 ( n348 , n86 , n1494 );
    not g344 ( n1724 , n829 );
    and g345 ( n1090 , n1392 , n1399 );
    or g346 ( n604 , n182 , n1050 );
    not g347 ( n860 , n1686 );
    xnor g348 ( n1572 , n1151 , n1429 );
    xnor g349 ( n1579 , n1308 , n1121 );
    not g350 ( n38 , n36 );
    not g351 ( n893 , n451 );
    or g352 ( n682 , n64 , n280 );
    xnor g353 ( n1256 , n330 , n1545 );
    and g354 ( n34 , n726 , n1754 );
    not g355 ( n771 , n1513 );
    not g356 ( n340 , n657 );
    not g357 ( n1746 , n856 );
    not g358 ( n1567 , n1005 );
    and g359 ( n358 , n534 , n138 );
    or g360 ( n824 , n926 , n462 );
    and g361 ( n619 , n1383 , n917 );
    and g362 ( n1203 , n830 , n1435 );
    xor g363 ( n536 , n1221 , n611 );
    xnor g364 ( n939 , n1318 , n1107 );
    or g365 ( n1667 , n103 , n843 );
    and g366 ( n1067 , n1522 , n421 );
    not g367 ( n1272 , n627 );
    not g368 ( n947 , n621 );
    nor g369 ( n1520 , n1 , n1706 );
    xor g370 ( n26 , n147 , n335 );
    not g371 ( n1027 , n1716 );
    and g372 ( n606 , n1238 , n1479 );
    or g373 ( n1757 , n1075 , n265 );
    and g374 ( n1570 , n1550 , n154 );
    not g375 ( n428 , n1245 );
    and g376 ( n1453 , n975 , n1138 );
    not g377 ( n1205 , n375 );
    and g378 ( n690 , n121 , n999 );
    or g379 ( n1263 , n1422 , n640 );
    xnor g380 ( n1216 , n1536 , n580 );
    and g381 ( n1687 , n1052 , n1234 );
    xnor g382 ( n992 , n586 , n525 );
    nor g383 ( n472 , n1024 , n1162 );
    and g384 ( n1307 , n392 , n877 );
    xnor g385 ( n1545 , n312 , n749 );
    and g386 ( n1532 , n1507 , n679 );
    or g387 ( n45 , n620 , n158 );
    and g388 ( n319 , n1245 , n425 );
    xnor g389 ( n1271 , n716 , n375 );
    or g390 ( n598 , n284 , n831 );
    xnor g391 ( n1523 , n1139 , n997 );
    not g392 ( n1566 , n706 );
    not g393 ( n17 , n1702 );
    not g394 ( n429 , n1640 );
    not g395 ( n22 , n1115 );
    not g396 ( n1431 , n1555 );
    nor g397 ( n620 , n1147 , n683 );
    not g398 ( n791 , n1466 );
    or g399 ( n981 , n1512 , n798 );
    or g400 ( n381 , n603 , n461 );
    and g401 ( n236 , n193 , n1149 );
    xnor g402 ( n1468 , n1129 , n731 );
    xnor g403 ( n797 , n784 , n1052 );
    not g404 ( n141 , n393 );
    not g405 ( n709 , n796 );
    nor g406 ( n775 , n835 , n1661 );
    and g407 ( n518 , n329 , n1433 );
    not g408 ( n170 , n308 );
    and g409 ( n237 , n1222 , n1478 );
    or g410 ( n1108 , n1570 , n108 );
    or g411 ( n46 , n491 , n915 );
    not g412 ( n257 , n1160 );
    and g413 ( n424 , n1325 , n1070 );
    or g414 ( n1668 , n852 , n365 );
    or g415 ( n384 , n272 , n919 );
    nor g416 ( n890 , n657 , n338 );
    xnor g417 ( n1524 , n1133 , n235 );
    and g418 ( n1103 , n1083 , n1649 );
    nor g419 ( n1751 , n896 , n1085 );
    or g420 ( n330 , n594 , n468 );
    xnor g421 ( n1169 , n88 , n1264 );
    or g422 ( n1540 , n515 , n294 );
    xnor g423 ( n845 , n629 , n202 );
    or g424 ( n1046 , n1062 , n1389 );
    or g425 ( n476 , n781 , n200 );
    nor g426 ( n574 , n306 , n925 );
    not g427 ( n1135 , n260 );
    nor g428 ( n173 , n1210 , n847 );
    not g429 ( n543 , n950 );
    not g430 ( n631 , n1198 );
    and g431 ( n466 , n641 , n648 );
    not g432 ( n3 , n1132 );
    not g433 ( n1137 , n1184 );
    xnor g434 ( n56 , n1184 , n930 );
    or g435 ( n314 , n593 , n947 );
    xor g436 ( n532 , n1653 , n1349 );
    nor g437 ( n1036 , n5 , n399 );
    xnor g438 ( n565 , n616 , n194 );
    or g439 ( n296 , n544 , n1148 );
    and g440 ( n430 , n580 , n1536 );
    not g441 ( n1549 , n693 );
    xnor g442 ( n756 , n355 , n1762 );
    and g443 ( n395 , n1129 , n662 );
    or g444 ( n117 , n529 , n1443 );
    or g445 ( n80 , n406 , n1286 );
    and g446 ( n946 , n523 , n649 );
    not g447 ( n962 , n687 );
    or g448 ( n739 , n1631 , n261 );
    not g449 ( n835 , n442 );
    or g450 ( n288 , n31 , n539 );
    buf g451 ( n1409 , n1468 );
    and g452 ( n477 , n1400 , n469 );
    or g453 ( n1215 , n283 , n492 );
    or g454 ( n218 , n897 , n1349 );
    not g455 ( n1424 , n412 );
    and g456 ( n1304 , n1572 , n1532 );
    or g457 ( n1040 , n1547 , n604 );
    or g458 ( n1656 , n502 , n1219 );
    nor g459 ( n1338 , n1462 , n1068 );
    xnor g460 ( n1348 , n736 , n1608 );
    nor g461 ( n467 , n13 , n906 );
    and g462 ( n548 , n446 , n1415 );
    and g463 ( n378 , n336 , n1063 );
    nor g464 ( n1454 , n1707 , n1065 );
    or g465 ( n671 , n1390 , n255 );
    and g466 ( n1398 , n1661 , n1498 );
    nor g467 ( n1092 , n1052 , n179 );
    nor g468 ( n174 , n599 , n990 );
    or g469 ( n1068 , n45 , n1416 );
    or g470 ( n1129 , n319 , n1527 );
    or g471 ( n269 , n1337 , n405 );
    not g472 ( n502 , n1147 );
    or g473 ( n753 , n883 , n1135 );
    buf g474 ( n644 , n808 );
    not g475 ( n970 , n1605 );
    xnor g476 ( n389 , n412 , n1245 );
    buf g477 ( n1024 , n1696 );
    xnor g478 ( n1127 , n850 , n871 );
    not g479 ( n1223 , n1320 );
    xnor g480 ( n1107 , n310 , n814 );
    not g481 ( n1528 , n554 );
    xnor g482 ( n858 , n822 , n750 );
    not g483 ( n1319 , n1640 );
    xnor g484 ( n957 , n1609 , n512 );
    not g485 ( n5 , n1077 );
    xnor g486 ( n438 , n618 , n833 );
    not g487 ( n1109 , n826 );
    not g488 ( n1727 , n694 );
    and g489 ( n761 , n862 , n288 );
    nor g490 ( n582 , n807 , n1052 );
    xor g491 ( n1076 , n1678 , n1271 );
    xnor g492 ( n136 , n1467 , n1459 );
    xor g493 ( n1190 , n913 , n423 );
    buf g494 ( n698 , 1'b0 );
    and g495 ( n628 , n1633 , n689 );
    and g496 ( n33 , n404 , n685 );
    not g497 ( n665 , n1470 );
    nor g498 ( n1053 , n302 , n262 );
    not g499 ( n1578 , n1012 );
    not g500 ( n109 , n1665 );
    or g501 ( n1602 , n1620 , n330 );
    xnor g502 ( n285 , n949 , n1134 );
    and g503 ( n1251 , n650 , n241 );
    xnor g504 ( n128 , n69 , n1579 );
    or g505 ( n1556 , n683 , n722 );
    not g506 ( n1707 , n652 );
    not g507 ( n1010 , n495 );
    or g508 ( n877 , n1002 , n721 );
    or g509 ( n460 , n1687 , n1554 );
    or g510 ( n1642 , n456 , n1658 );
    xnor g511 ( n750 , n122 , n1486 );
    or g512 ( n975 , n947 , n1740 );
    xnor g513 ( n135 , n1249 , n625 );
    and g514 ( n693 , n1623 , n1198 );
    xnor g515 ( n82 , n712 , n331 );
    nor g516 ( n1499 , n1024 , n1014 );
    xnor g517 ( n651 , n99 , n1557 );
    not g518 ( n1756 , n1303 );
    not g519 ( n1496 , n1034 );
    not g520 ( n1278 , n1473 );
    or g521 ( n1192 , n54 , n1740 );
    not g522 ( n112 , n707 );
    not g523 ( n1374 , n118 );
    not g524 ( n581 , n1744 );
    and g525 ( n1316 , n619 , n274 );
    and g526 ( n252 , n587 , n682 );
    not g527 ( n1643 , n521 );
    not g528 ( n1177 , n1300 );
    not g529 ( n133 , n893 );
    not g530 ( n1238 , n1266 );
    not g531 ( n352 , n1247 );
    not g532 ( n336 , n58 );
    nor g533 ( n1737 , n644 , n1323 );
    xnor g534 ( n1423 , n507 , n403 );
    xor g535 ( n760 , n1360 , n52 );
    xnor g536 ( n956 , n1068 , n1462 );
    and g537 ( n1259 , n10 , n1080 );
    and g538 ( n329 , n1746 , n422 );
    and g539 ( n1025 , n1118 , n423 );
    and g540 ( n120 , n162 , n1264 );
    nor g541 ( n659 , n967 , n1317 );
    xnor g542 ( n291 , n1576 , n1371 );
    not g543 ( n794 , n960 );
    and g544 ( n697 , n610 , n458 );
    not g545 ( n552 , n1536 );
    xnor g546 ( n1063 , n1497 , n1342 );
    not g547 ( n1156 , n481 );
    or g548 ( n1164 , n300 , n64 );
    xor g549 ( n1009 , n641 , n648 );
    and g550 ( n1527 , n1725 , n1073 );
    not g551 ( n270 , n768 );
    nor g552 ( n943 , n28 , n1170 );
    or g553 ( n1531 , n1707 , n1426 );
    not g554 ( n1353 , n626 );
    xor g555 ( n111 , n84 , n1183 );
    and g556 ( n922 , n271 , n213 );
    and g557 ( n1412 , n892 , n891 );
    or g558 ( n1717 , n574 , n65 );
    or g559 ( n603 , n1657 , n372 );
    or g560 ( n10 , n759 , n1671 );
    xnor g561 ( n1102 , n1059 , n1158 );
    xor g562 ( n1604 , n147 , n329 );
    not g563 ( n1299 , n1696 );
    and g564 ( n272 , n1589 , n1611 );
    xor g565 ( n1072 , n1720 , n961 );
    or g566 ( n1552 , n413 , n263 );
    not g567 ( n804 , n1314 );
    or g568 ( n1133 , n1751 , n878 );
    or g569 ( n152 , n333 , n572 );
    and g570 ( n1324 , n373 , n1533 );
    not g571 ( n1314 , n1334 );
    or g572 ( n1480 , n969 , n510 );
    and g573 ( n471 , n1441 , n1683 );
    not g574 ( n1249 , n839 );
    xnor g575 ( n615 , n291 , n117 );
    or g576 ( n1627 , n644 , n1060 );
    and g577 ( n1339 , n721 , n1285 );
    and g578 ( n510 , n663 , n903 );
    xnor g579 ( n333 , n578 , n118 );
    xnor g580 ( n1755 , n37 , n1031 );
    and g581 ( n390 , n671 , n226 );
    and g582 ( n106 , n562 , n795 );
    or g583 ( n892 , n1597 , n180 );
    xnor g584 ( n886 , n421 , n637 );
    and g585 ( n1048 , n1160 , n914 );
    or g586 ( n776 , n443 , n325 );
    not g587 ( n614 , n185 );
    buf g588 ( n1134 , n1368 );
    not g589 ( n653 , n281 );
    xnor g590 ( n151 , n1157 , n1494 );
    not g591 ( n1105 , n388 );
    not g592 ( n1162 , n1328 );
    not g593 ( n500 , n923 );
    xnor g594 ( n464 , n126 , n1665 );
    not g595 ( n1638 , n440 );
    xnor g596 ( n529 , n1276 , n1303 );
    not g597 ( n996 , n1625 );
    nor g598 ( n121 , n704 , n732 );
    not g599 ( n1375 , n749 );
    xnor g600 ( n171 , n488 , n19 );
    not g601 ( n1703 , n515 );
    not g602 ( n1659 , n725 );
    and g603 ( n712 , n197 , n407 );
    xnor g604 ( n1574 , n1022 , n1218 );
    and g605 ( n1490 , n1602 , n579 );
    and g606 ( n774 , n215 , n924 );
    xnor g607 ( n1650 , n1755 , n1170 );
    or g608 ( n1152 , n1318 , n718 );
    not g609 ( n1471 , n1704 );
    not g610 ( n1376 , n1248 );
    xnor g611 ( n317 , n848 , n660 );
    not g612 ( n1384 , n241 );
    or g613 ( n1138 , n1205 , n223 );
    not g614 ( n839 , n72 );
    or g615 ( n453 , n775 , n1398 );
    or g616 ( n400 , n622 , n163 );
    or g617 ( n1281 , n201 , n598 );
    or g618 ( n958 , n410 , n1600 );
    xnor g619 ( n1106 , n1168 , n463 );
    or g620 ( n1301 , n1063 , n360 );
    xnor g621 ( n648 , n507 , n371 );
    not g622 ( n573 , n1683 );
    or g623 ( n1758 , n1193 , n1678 );
    or g624 ( n212 , n396 , n20 );
    nor g625 ( n819 , n913 , n559 );
    not g626 ( n931 , n1479 );
    or g627 ( n1081 , n368 , n479 );
    or g628 ( n742 , n50 , n295 );
    or g629 ( n1261 , n841 , n1017 );
    and g630 ( n84 , n356 , n497 );
    not g631 ( n1116 , n657 );
    or g632 ( n903 , n201 , n880 );
    and g633 ( n1094 , n379 , n541 );
    xnor g634 ( n1069 , n697 , n1723 );
    not g635 ( n509 , n57 );
    xnor g636 ( n1526 , n1259 , n556 );
    not g637 ( n1117 , n143 );
    or g638 ( n1269 , n1032 , n376 );
    xnor g639 ( n266 , n270 , n135 );
    not g640 ( n1136 , n257 );
    not g641 ( n1262 , n889 );
    not g642 ( n1015 , n1441 );
    or g643 ( n318 , n1553 , n237 );
    or g644 ( n1537 , n552 , n1344 );
    xnor g645 ( n972 , n104 , n1204 );
    or g646 ( n301 , n127 , n1242 );
    not g647 ( n934 , n191 );
    not g648 ( n925 , n316 );
    and g649 ( n1625 , n23 , n1735 );
    and g650 ( n999 , n134 , n1140 );
    not g651 ( n311 , n811 );
    or g652 ( n377 , n825 , n1259 );
    nor g653 ( n1451 , n1147 , n1182 );
    not g654 ( n176 , n661 );
    xnor g655 ( n206 , n895 , n150 );
    not g656 ( n1510 , n1681 );
    and g657 ( n1626 , n1727 , n816 );
    not g658 ( n1163 , n784 );
    xnor g659 ( n1352 , n1488 , n94 );
    not g660 ( n361 , n1046 );
    not g661 ( n805 , n1431 );
    not g662 ( n405 , n688 );
    nor g663 ( n1056 , n1470 , n1742 );
    or g664 ( n1230 , n936 , n1100 );
    xnor g665 ( n440 , n65 , n770 );
    or g666 ( n1312 , n1067 , n1103 );
    and g667 ( n1631 , n342 , n1197 );
    xnor g668 ( n18 , n926 , n1111 );
    buf g669 ( n883 , n1354 );
    or g670 ( n623 , n430 , n1217 );
    not g671 ( n447 , n247 );
    or g672 ( n37 , n982 , n963 );
    and g673 ( n670 , n419 , n1684 );
    or g674 ( n123 , n657 , n436 );
    not g675 ( n468 , n809 );
    and g676 ( n1059 , n568 , n764 );
    not g677 ( n445 , n185 );
    nor g678 ( n991 , n655 , n111 );
    nor g679 ( n459 , n1619 , n482 );
    and g680 ( n356 , n1573 , n567 );
    or g681 ( n1155 , n1596 , n597 );
    and g682 ( n194 , n668 , n1465 );
    not g683 ( n1741 , n710 );
    nor g684 ( n546 , n970 , n1116 );
    xnor g685 ( n945 , n934 , n396 );
    not g686 ( n1293 , n45 );
    not g687 ( n1644 , n1484 );
    or g688 ( n124 , n8 , n184 );
    xnor g689 ( n1533 , n1440 , n388 );
    xnor g690 ( n626 , n521 , n464 );
    nor g691 ( n1333 , n340 , n947 );
    not g692 ( n228 , n1013 );
    not g693 ( n803 , n1313 );
    and g694 ( n230 , n1668 , n1152 );
    nor g695 ( n1565 , n1172 , n1494 );
    or g696 ( n1194 , n477 , n1304 );
    nor g697 ( n983 , n744 , n1245 );
    xnor g698 ( n987 , n245 , n1517 );
    or g699 ( n856 , n31 , n143 );
    and g700 ( n1683 , n806 , n528 );
    xnor g701 ( n264 , n1028 , n195 );
    xnor g702 ( n24 , n476 , n581 );
    or g703 ( n1153 , n409 , n1377 );
    buf g704 ( n523 , n1248 );
    not g705 ( n201 , n1132 );
    not g706 ( n950 , n536 );
    or g707 ( n1440 , n1374 , n578 );
    not g708 ( n1747 , n1128 );
    and g709 ( n517 , n7 , n124 );
    or g710 ( n568 , n171 , n1637 );
    not g711 ( n1621 , n927 );
    not g712 ( n1378 , n658 );
    nor g713 ( n841 , n953 , n580 );
    xnor g714 ( n1582 , n1411 , n979 );
    not g715 ( n545 , n280 );
    xnor g716 ( n304 , n1420 , n1534 );
    not g717 ( n843 , n1566 );
    buf g718 ( n184 , n1199 );
    not g719 ( n1675 , n744 );
    and g720 ( n1368 , n1720 , n961 );
    not g721 ( n162 , n232 );
    and g722 ( n227 , n493 , n1738 );
    xnor g723 ( n324 , n1591 , n74 );
    not g724 ( n815 , n829 );
    nor g725 ( n988 , n247 , n453 );
    nor g726 ( n576 , n1320 , n312 );
    and g727 ( n23 , n1605 , n1686 );
    not g728 ( n1492 , n1066 );
    xnor g729 ( n1541 , n726 , n686 );
    not g730 ( n1377 , n848 );
    not g731 ( n205 , n310 );
    not g732 ( n450 , n1241 );
    buf g733 ( n102 , 1'b0 );
    nor g734 ( n161 , n1064 , n1086 );
    nor g735 ( n75 , n832 , n157 );
    xnor g736 ( n498 , n1070 , n617 );
    and g737 ( n365 , n1108 , n884 );
    and g738 ( n904 , n321 , n480 );
    xor g739 ( n570 , n1617 , n709 );
    not g740 ( n1691 , n1314 );
    not g741 ( n594 , n625 );
    or g742 ( n1226 , n1333 , n362 );
    or g743 ( n505 , n132 , n614 );
    not g744 ( n1323 , n664 );
    xnor g745 ( n455 , n1066 , n849 );
    not g746 ( n496 , n1706 );
    xnor g747 ( n592 , n1671 , n83 );
    or g748 ( n743 , n661 , n1241 );
    not g749 ( n451 , n1549 );
    xnor g750 ( n1433 , n100 , n793 );
    xnor g751 ( n1034 , n457 , n703 );
    xnor g752 ( n611 , n184 , n857 );
    or g753 ( n885 , n546 , n1753 );
    not g754 ( n1084 , n280 );
    not g755 ( n376 , n1245 );
    xor g756 ( n1279 , n1226 , n670 );
    not g757 ( n1463 , n1648 );
    or g758 ( n399 , n1240 , n321 );
    or g759 ( n1425 , n1055 , n1136 );
    or g760 ( n446 , n348 , n1591 );
    xnor g761 ( n699 , n1119 , n1187 );
    not g762 ( n1416 , n820 );
    or g763 ( n1359 , n346 , n1321 );
    xnor g764 ( n360 , n885 , n1704 );
    and g765 ( n1273 , n49 , n212 );
    not g766 ( n1610 , n1160 );
    nor g767 ( n873 , n43 , n227 );
    buf g768 ( n831 , n549 );
    not g769 ( n1685 , n1431 );
    or g770 ( n142 , n1006 , n1041 );
    xnor g771 ( n1057 , n855 , n345 );
    not g772 ( n1144 , n448 );
    and g773 ( n313 , n1052 , n807 );
    nor g774 ( n982 , n1364 , n1740 );
    or g775 ( n827 , n533 , n1372 );
    or g776 ( n1715 , n1552 , n669 );
    xnor g777 ( n888 , n270 , n974 );
    xor g778 ( n229 , n1617 , n1411 );
    xnor g779 ( n1583 , n1414 , n1084 );
    and g780 ( n1206 , n543 , n1663 );
    nor g781 ( n1592 , n661 , n617 );
    xnor g782 ( n1639 , n598 , n1214 );
    not g783 ( n1575 , n56 );
    or g784 ( n526 , n87 , n873 );
    or g785 ( n571 , n1361 , n1097 );
    and g786 ( n1292 , n1584 , n437 );
    and g787 ( n1421 , n1043 , n1329 );
    or g788 ( n765 , n169 , n1001 );
    xnor g789 ( n714 , n1360 , n986 );
    xnor g790 ( n1459 , n1285 , n62 );
    and g791 ( n383 , n439 , n170 );
    xnor g792 ( n979 , n166 , n935 );
    xnor g793 ( n1614 , n487 , n1349 );
    not g794 ( n519 , n1612 );
    xnor g795 ( n1558 , n1732 , n856 );
    not g796 ( n51 , n1379 );
    or g797 ( n635 , n1388 , n1294 );
    or g798 ( n1174 , n1536 , n1721 );
    nor g799 ( n798 , n224 , n1168 );
    not g800 ( n977 , n564 );
    not g801 ( n456 , n1743 );
    not g802 ( n12 , n1749 );
    not g803 ( n190 , n1171 );
    not g804 ( n444 , n316 );
    not g805 ( n397 , n324 );
    not g806 ( n341 , n1167 );
    not g807 ( n1337 , n636 );
    not g808 ( n207 , n1020 );
    xnor g809 ( n129 , n678 , n901 );
    not g810 ( n276 , n1494 );
    or g811 ( n781 , n1304 , n1382 );
    and g812 ( n1372 , n598 , n3 );
    not g813 ( n491 , n306 );
    not g814 ( n1669 , n1326 );
    or g815 ( n353 , n1594 , n230 );
    xnor g816 ( n1752 , n364 , n687 );
    xnor g817 ( n779 , n1114 , n1624 );
    xnor g818 ( n862 , n267 , n386 );
    xnor g819 ( n792 , n1370 , n18 );
    xnor g820 ( n292 , n311 , n527 );
    not g821 ( n1285 , n1536 );
    and g822 ( n1128 , n1567 , n1423 );
    not g823 ( n215 , n814 );
    and g824 ( n315 , n1200 , n1605 );
    or g825 ( n985 , n1134 , n1689 );
    xor g826 ( n280 , n1379 , n1402 );
    xnor g827 ( n293 , n1201 , n1306 );
    not g828 ( n1542 , n901 );
    or g829 ( n47 , n1277 , n1245 );
    not g830 ( n185 , n1145 );
    and g831 ( n148 , n1535 , n37 );
    nor g832 ( n224 , n916 , n1494 );
    and g833 ( n531 , n708 , n1229 );
    and g834 ( n245 , n777 , n692 );
    or g835 ( n91 , n1571 , n1220 );
    not g836 ( n595 , n1442 );
    not g837 ( n81 , n989 );
    xnor g838 ( n418 , n1754 , n333 );
    and g839 ( n21 , n513 , n1491 );
    xnor g840 ( n235 , n1551 , n644 );
    nor g841 ( n1041 , n503 , n1316 );
    not g842 ( n452 , n308 );
    not g843 ( n964 , n466 );
    not g844 ( n499 , n172 );
    xnor g845 ( n1381 , n781 , n1630 );
    not g846 ( n1508 , n1279 );
    or g847 ( n1007 , n170 , n591 );
    xnor g848 ( n867 , n724 , n1171 );
    xnor g849 ( n1472 , n91 , n285 );
    not g850 ( n165 , n1378 );
    not g851 ( n307 , n1507 );
    xnor g852 ( n1761 , n373 , n1533 );
    not g853 ( n1617 , n385 );
    not g854 ( n260 , n1272 );
    or g855 ( n36 , n1714 , n359 );
    and g856 ( n168 , n90 , n457 );
    xnor g857 ( n1264 , n1642 , n989 );
    not g858 ( n586 , n616 );
    not g859 ( n638 , n1624 );
    or g860 ( n923 , n1109 , n207 );
    and g861 ( n1678 , n225 , n746 );
    xor g862 ( n1702 , n1460 , n1523 );
    and g863 ( n267 , n1758 , n70 );
    xnor g864 ( n139 , n1114 , n1640 );
    xnor g865 ( n808 , n414 , n1141 );
    and g866 ( n813 , n1127 , n1147 );
    xnor g867 ( n27 , n535 , n1694 );
    and g868 ( n1479 , n846 , n1487 );
    not g869 ( n503 , n385 );
    and g870 ( n701 , n1463 , n547 );
    xnor g871 ( n391 , n1615 , n1439 );
    not g872 ( n131 , n461 );
    xnor g873 ( n154 , n1622 , n859 );
    buf g874 ( n396 , n889 );
    xnor g875 ( n1004 , n32 , n204 );
    and g876 ( n157 , n918 , n1531 );
    xnor g877 ( n1419 , n1552 , n1134 );
    and g878 ( n1437 , n1733 , n1686 );
    not g879 ( n901 , n1252 );
    or g880 ( n758 , n452 , n1471 );
    not g881 ( n232 , n238 );
    and g882 ( n69 , n1023 , n751 );
    nor g883 ( n955 , n626 , n966 );
    or g884 ( n1591 , n645 , n1369 );
    not g885 ( n1555 , n145 );
    or g886 ( n944 , n666 , n1418 );
    xnor g887 ( n275 , n1330 , n240 );
    or g888 ( n663 , n482 , n1740 );
    or g889 ( n703 , n1137 , n1283 );
    or g890 ( n1033 , n1234 , n1052 );
    not g891 ( n1530 , n805 );
    not g892 ( n1550 , n545 );
    not g893 ( n1055 , n1134 );
    xnor g894 ( n1450 , n1495 , n216 );
    xnor g895 ( n1731 , n248 , n1065 );
    not g896 ( n1060 , n499 );
    xnor g897 ( n715 , n390 , n1450 );
    xnor g898 ( n1121 , n1658 , n1743 );
    not g899 ( n210 , n1284 );
    xnor g900 ( n79 , n176 , n1432 );
    and g901 ( n1233 , n818 , n657 );
    or g902 ( n980 , n1435 , n438 );
    xnor g903 ( n823 , n141 , n171 );
    nor g904 ( n1078 , n1245 , n184 );
    nor g905 ( n1006 , n274 , n619 );
    or g906 ( n416 , n946 , n1599 );
    nor g907 ( n1518 , n437 , n627 );
    xnor g908 ( n41 , n558 , n740 );
    or g909 ( n564 , n1728 , n1451 );
    nor g910 ( n305 , n221 , n117 );
    not g911 ( n448 , n510 );
    not g912 ( n182 , n1625 );
    not g913 ( n723 , n495 );
    not g914 ( n539 , n1076 );
    buf g915 ( n580 , n149 );
    or g916 ( n372 , n81 , n1642 );
    and g917 ( n599 , n111 , n655 );
    xnor g918 ( n486 , n614 , n132 );
    not g919 ( n219 , n403 );
    or g920 ( n411 , n1394 , n1498 );
    or g921 ( n900 , n1536 , n580 );
    not g922 ( n1113 , n796 );
    not g923 ( n830 , n560 );
    not g924 ( n836 , n757 );
    xnor g925 ( n327 , n1706 , n1 );
    not g926 ( n248 , n652 );
    and g927 ( n607 , n634 , n632 );
    not g928 ( n1228 , n718 );
    xnor g929 ( n254 , n996 , n1612 );
    or g930 ( n166 , n542 , n374 );
    and g931 ( n1560 , n1181 , n339 );
    xnor g932 ( n19 , n312 , n1320 );
    nor g933 ( n769 , n583 , n482 );
    or g934 ( n1300 , n769 , n1482 );
    not g935 ( n921 , n1662 );
    xor g936 ( n1077 , n1197 , n1516 );
    nor g937 ( n1062 , n1054 , n1430 );
    xnor g938 ( n608 , n1662 , n367 );
    xnor g939 ( n724 , n310 , n707 );
    or g940 ( n251 , n467 , n1053 );
    and g941 ( n821 , n1494 , n1692 );
    or g942 ( n1248 , n1477 , n250 );
    xnor g943 ( n483 , n420 , n1682 );
    and g944 ( n559 , n966 , n334 );
    xnor g945 ( n1719 , n1295 , n738 );
    not g946 ( n1498 , n442 );
    or g947 ( n297 , n1628 , n1059 );
    nor g948 ( n1718 , n1339 , n246 );
    nor g949 ( n1026 , n680 , n1337 );
    xnor g950 ( n367 , n1191 , n99 );
    and g951 ( n1151 , n400 , n1126 );
    xnor g952 ( n875 , n1412 , n797 );
    not g953 ( n119 , n719 );
    and g954 ( n963 , n1740 , n423 );
    not g955 ( n338 , n204 );
    not g956 ( n784 , n51 );
    not g957 ( n1661 , n63 );
    buf g958 ( n642 , n1445 );
    not g959 ( n146 , n1759 );
    and g960 ( n137 , n776 , n381 );
    xnor g961 ( n103 , n540 , n192 );
    or g962 ( n178 , n421 , n462 );
    or g963 ( n1371 , n810 , n1756 );
    not g964 ( n969 , n1494 );
    and g965 ( n231 , n84 , n347 );
    and g966 ( n1217 , n1712 , n900 );
    not g967 ( n298 , n555 );
    or g968 ( n1506 , n844 , n1485 );
    not g969 ( n1422 , n1236 );
    not g970 ( n1115 , n674 );
    or g971 ( n1460 , n794 , n361 );
    and g972 ( n986 , n1008 , n518 );
    xnor g973 ( n39 , n184 , n1673 );
    xnor g974 ( n1514 , n1010 , n680 );
    xnor g975 ( n567 , n606 , n1236 );
    not g976 ( n67 , n526 );
    xnor g977 ( n1763 , n1277 , n1245 );
    not g978 ( n767 , n974 );
    nor g979 ( n1726 , n1119 , n1448 );
    and g980 ( n1426 , n1634 , n1672 );
    not g981 ( n1611 , n1134 );
    not g982 ( n93 , n195 );
    not g983 ( n994 , n1256 );
    not g984 ( n1260 , n672 );
    xnor g985 ( n1393 , n255 , n485 );
    or g986 ( n746 , n338 , n406 );
    xnor g987 ( n1676 , n1345 , n1349 );
    and g988 ( n1513 , n780 , n515 );
    and g989 ( n1185 , n56 , n189 );
    not g990 ( n426 , n1455 );
    not g991 ( n688 , n1202 );
    or g992 ( n98 , n1502 , n396 );
    xnor g993 ( n1404 , n33 , n498 );
    or g994 ( n777 , n506 , n390 );
    not g995 ( n489 , n417 );
    and g996 ( n1148 , n737 , n470 );
    or g997 ( n869 , n1243 , n1408 );
    xnor g998 ( n1666 , n1128 , n937 );
    nor g999 ( n1427 , n661 , n1621 );
    nor g1000 ( n1093 , n1702 , n696 );
    nor g1001 ( n208 , n1605 , n210 );
    not g1002 ( n1493 , n450 );
    not g1003 ( n674 , n1453 );
    nor g1004 ( n346 , n94 , n1157 );
    and g1005 ( n295 , n340 , n423 );
    nor g1006 ( n1651 , n300 , n880 );
    xnor g1007 ( n1534 , n1356 , n1085 );
    or g1008 ( n310 , n315 , n1165 );
    xnor g1009 ( n740 , n1260 , n396 );
    or g1010 ( n1684 , n1096 , n804 );
    or g1011 ( n587 , n1737 , n501 );
    not g1012 ( n1213 , n264 );
    xnor g1013 ( n169 , n905 , n1007 );
    not g1014 ( n1394 , n1349 );
    xnor g1015 ( n1122 , n1493 , n508 );
    not g1016 ( n347 , n1183 );
    or g1017 ( n1483 , n1278 , n1394 );
    and g1018 ( n1606 , n819 , n423 );
    not g1019 ( n1635 , n661 );
    and g1020 ( n1075 , n922 , n1386 );
    xnor g1021 ( n427 , n1486 , n627 );
    or g1022 ( n634 , n1529 , n1499 );
    or g1023 ( n1662 , n73 , n747 );
    and g1024 ( n1500 , n416 , n1757 );
    not g1025 ( n1713 , n1112 );
    not g1026 ( n928 , n1291 );
    xnor g1027 ( n326 , n948 , n1122 );
    nor g1028 ( n763 , n941 , n137 );
    xnor g1029 ( n289 , n1319 , n557 );
    not g1030 ( n153 , n257 );
    or g1031 ( n97 , n376 , n915 );
    not g1032 ( n1239 , n833 );
    xnor g1033 ( n186 , n143 , n1732 );
    xor g1034 ( n643 , n834 , n758 );
    not g1035 ( n1145 , n1085 );
    xnor g1036 ( n1655 , n479 , n1124 );
    or g1037 ( n692 , n1495 , n843 );
    not g1038 ( n1334 , n1199 );
    not g1039 ( n1104 , n1049 );
    not g1040 ( n1505 , n1031 );
    and g1041 ( n1401 , n1266 , n931 );
    xnor g1042 ( n181 , n1038 , n1363 );
    and g1043 ( n1603 , n1578 , n1134 );
    or g1044 ( n585 , n932 , n1370 );
    nor g1045 ( n1389 , n1147 , n436 );
    not g1046 ( n1096 , n1673 );
    xnor g1047 ( n1214 , n141 , n1132 );
    xnor g1048 ( n457 , n905 , n383 );
    or g1049 ( n1130 , n734 , n507 );
    xnor g1050 ( n1331 , n1100 , n129 );
    not g1051 ( n722 , n1134 );
    xnor g1052 ( n1380 , n22 , n1349 );
    or g1053 ( n584 , n454 , n1038 );
    or g1054 ( n948 , n1154 , n1417 );
    not g1055 ( n1589 , n1610 );
    or g1056 ( n402 , n1213 , n1113 );
    xnor g1057 ( n89 , n1568 , n465 );
    not g1058 ( n637 , n676 );
    xnor g1059 ( n806 , n772 , n1391 );
    not g1060 ( n239 , n875 );
    and g1061 ( n1220 , n951 , n222 );
    not g1062 ( n1364 , n871 );
    xnor g1063 ( n800 , n1748 , n480 );
    not g1064 ( n434 , n529 );
    or g1065 ( n789 , n896 , n836 );
    not g1066 ( n1011 , n37 );
    or g1067 ( n164 , n211 , n1618 );
    or g1068 ( n504 , n369 , n245 );
    or g1069 ( n762 , n89 , n1279 );
    or g1070 ( n140 , n962 , n1453 );
    not g1071 ( n1146 , n1741 );
    or g1072 ( n1268 , n766 , n122 );
    xnor g1073 ( n1298 , n713 , n292 );
    xnor g1074 ( n203 , n142 , n1731 );
    and g1075 ( n1087 , n223 , n1562 );
    and g1076 ( n1170 , n1366 , n1250 );
    not g1077 ( n555 , n78 );
    xnor g1078 ( n83 , n417 , n1494 );
    xnor g1079 ( n1310 , n501 , n1583 );
    not g1080 ( n840 , n677 );
    not g1081 ( n1157 , n1144 );
    and g1082 ( n544 , n303 , n89 );
    not g1083 ( n1521 , n822 );
    xnor g1084 ( n556 , n745 , n1245 );
    not g1085 ( n243 , n1384 );
    and g1086 ( n865 , n85 , n1164 );
    xnor g1087 ( n1318 , n36 , n484 );
    not g1088 ( n640 , n606 );
    not g1089 ( n716 , n1561 );
    not g1090 ( n993 , n484 );
    not g1091 ( n710 , n933 );
    not g1092 ( n240 , n1350 );
    and g1093 ( n342 , n332 , n1297 );
    not g1094 ( n1295 , n602 );
    xnor g1095 ( n691 , n906 , n229 );
    xnor g1096 ( n465 , n1473 , n1349 );
    and g1097 ( n1573 , n633 , n870 );
    not g1098 ( n1736 , n1503 );
    or g1099 ( n1047 , n1588 , n1090 );
    not g1100 ( n1050 , n1416 );
    xor g1101 ( n1696 , n799 , n702 );
    and g1102 ( n707 , n1180 , n287 );
    nor g1103 ( n1193 , n375 , n1409 );
    or g1104 ( n1201 , n110 , n782 );
    not g1105 ( n1079 , n415 );
    or g1106 ( n1080 , n489 , n969 );
    not g1107 ( n1247 , n709 );
    or g1108 ( n250 , n834 , n758 );
    nor g1109 ( n801 , n649 , n523 );
    not g1110 ( n811 , n533 );
    xnor g1111 ( n1005 , n1046 , n960 );
    not g1112 ( n1716 , n1410 );
    xnor g1113 ( n268 , n1246 , n1161 );
    and g1114 ( n1636 , n593 , n423 );
    not g1115 ( n718 , n1107 );
    nor g1116 ( n675 , n349 , n1275 );
    and g1117 ( n654 , n1349 , n1290 );
    not g1118 ( n1466 , n1484 );
    or g1119 ( n848 , n1224 , n659 );
    xnor g1120 ( n249 , n1130 , n1343 );
    and g1121 ( n1099 , n572 , n333 );
    and g1122 ( n624 , n623 , n209 );
    not g1123 ( n1197 , n183 );
    or g1124 ( n138 , n1424 , n376 );
    or g1125 ( n1478 , n860 , n1116 );
    and g1126 ( n443 , n461 , n603 );
    not g1127 ( n1733 , n1347 );
    xnor g1128 ( n802 , n1013 , n765 );
    not g1129 ( n780 , n1007 );
    xnor g1130 ( n401 , n1273 , n570 );
    or g1131 ( n629 , n1105 , n1440 );
    or g1132 ( n1465 , n1055 , n1027 );
    not g1133 ( n31 , n602 );
    or g1134 ( n1366 , n1048 , n1307 );
    not g1135 ( n1054 , n1147 );
    not g1136 ( n122 , n1143 );
    or g1137 ( n795 , n1533 , n1135 );
    not g1138 ( n1035 , n618 );
    not g1139 ( n328 , n499 );
    or g1140 ( n1287 , n675 , n1569 );
    not g1141 ( n78 , n343 );
    not g1142 ( n1432 , n107 );
    xor g1143 ( n1484 , n1573 , n567 );
    xnor g1144 ( n859 , n1265 , n1052 );
    xnor g1145 ( n937 , n527 , n1106 );
    not g1146 ( n1753 , n1564 );
    and g1147 ( n561 , n713 , n1024 );
    not g1148 ( n1452 , n1349 );
    xnor g1149 ( n1663 , n548 , n389 );
    not g1150 ( n1443 , n1421 );
    not g1151 ( n48 , n86 );
    and g1152 ( n650 , n157 , n832 );
    and g1153 ( n713 , n1567 , n942 );
    xnor g1154 ( n1694 , n845 , n719 );
    not g1155 ( n583 , n657 );
    and g1156 ( n1097 , n1506 , n490 );
    not g1157 ( n968 , n166 );
    or g1158 ( n321 , n228 , n765 );
    buf g1159 ( n1536 , n1072 );
    or g1160 ( n822 , n1750 , n161 );
    and g1161 ( n1236 , n752 , n1656 );
    or g1162 ( n1031 , n810 , n146 );
    not g1163 ( n436 , n66 );
    and g1164 ( n1088 , n384 , n1425 );
    xnor g1165 ( n1070 , n1563 , n16 );
    or g1166 ( n534 , n788 , n548 );
    buf g1167 ( n1580 , 1'b0 );
    not g1168 ( n332 , n1548 );
    and g1169 ( n820 , n40 , n522 );
    not g1170 ( n155 , n657 );
    buf g1171 ( n1734 , n1639 );
    xnor g1172 ( n842 , n1175 , n1529 );
    nor g1173 ( n116 , n1665 , n1134 );
    or g1174 ( n853 , n1635 , n107 );
    not g1175 ( n1240 , n800 );
    xor g1176 ( n566 , n1444 , n590 );
    or g1177 ( n209 , n1134 , n866 );
    not g1178 ( n810 , n1276 );
    or g1179 ( n870 , n1401 , n606 );
    and g1180 ( n1444 , n724 , n190 );
    and g1181 ( n355 , n1312 , n178 );
    not g1182 ( n1698 , n898 );
    and g1183 ( n540 , n1699 , n1483 );
    xnor g1184 ( n1469 , n826 , n1020 );
    and g1185 ( n1242 , n571 , n550 );
    xnor g1186 ( n1179 , n897 , n1349 );
    or g1187 ( n1171 , n471 , n875 );
    not g1188 ( n1140 , n1200 );
    or g1189 ( n1383 , n1253 , n558 );
    nor g1190 ( n15 , n1052 , n1379 );
    or g1191 ( n197 , n600 , n1021 );
    xnor g1192 ( n912 , n653 , n1134 );
    or g1193 ( n910 , n1147 , n253 );
    not g1194 ( n279 , n460 );
    nor g1195 ( n938 , n286 , n104 );
    not g1196 ( n520 , n94 );
    xnor g1197 ( n1641 , n800 , n321 );
    not g1198 ( n766 , n652 );
    or g1199 ( n1680 , n576 , n488 );
    not g1200 ( n4 , n1297 );
    or g1201 ( n917 , n396 , n160 );
    nor g1202 ( n812 , n204 , n661 );
    nor g1203 ( n1637 , n1024 , n928 );
    not g1204 ( n274 , n1042 );
    not g1205 ( n1730 , n509 );
    and g1206 ( n1022 , n767 , n1629 );
    or g1207 ( n1255 , n1018 , n1407 );
    and g1208 ( n108 , n1230 , n199 );
    not g1209 ( n52 , n650 );
    not g1210 ( n738 , n1076 );
    and g1211 ( n1485 , n882 , n505 );
    not g1212 ( n1173 , n644 );
    nor g1213 ( n1438 , n722 , n1546 );
    not g1214 ( n861 , n1585 );
    xnor g1215 ( n601 , n1686 , n1605 );
    and g1216 ( n263 , n231 , n956 );
    not g1217 ( n1294 , n535 );
    xnor g1218 ( n1336 , n89 , n1510 );
    or g1219 ( n1049 , n459 , n114 );
    xnor g1220 ( n785 , n957 , n137 );
    not g1221 ( n572 , n1644 );
    or g1222 ( n512 , n236 , n580 );
    and g1223 ( n1303 , n500 , n35 );
    not g1224 ( n286 , n249 );
    or g1225 ( n187 , n883 , n595 );
    or g1226 ( n1282 , n1026 , n865 );
    xnor g1227 ( n1237 , n695 , n427 );
    and g1228 ( n786 , n1735 , n657 );
    and g1229 ( n262 , n906 , n13 );
    nor g1230 ( n1154 , n1106 , n1747 );
    or g1231 ( n70 , n253 , n716 );
    and g1232 ( n65 , n1359 , n1362 );
    nor g1233 ( n76 , n1303 , n1421 );
    and g1234 ( n439 , n1398 , n237 );
    not g1235 ( n1410 , n265 );
    and g1236 ( n1652 , n113 , n508 );
    xnor g1237 ( n1343 , n1172 , n1494 );
    not g1238 ( n554 , n237 );
    and g1239 ( n271 , n968 , n935 );
    not g1240 ( n253 , n375 );
    nor g1241 ( n408 , n1265 , n1052 );
    not g1242 ( n1341 , n1049 );
    not g1243 ( n1495 , n644 );
    nor g1244 ( n1728 , n1619 , n54 );
    or g1245 ( n846 , n1147 , n173 );
    and g1246 ( n669 , n849 , n1492 );
    not g1247 ( n259 , n742 );
    nor g1248 ( n410 , n1345 , n1349 );
    not g1249 ( n1411 , n729 );
    not g1250 ( n1211 , n1188 );
    not g1251 ( n72 , n1701 );
    nor g1252 ( n1690 , n1134 , n265 );
    xnor g1253 ( n1470 , n909 , n244 );
    not g1254 ( n941 , n957 );
    or g1255 ( n562 , n1099 , n278 );
    xnor g1256 ( n1632 , n394 , n912 );
    xnor g1257 ( n1082 , n1506 , n920 );
    xnor g1258 ( n282 , n990 , n894 );
    buf g1259 ( n1519 , 1'b0 );
    not g1260 ( n1559 , n242 );
    xnor g1261 ( n1522 , n517 , n159 );
    or g1262 ( n134 , n1623 , n970 );
    and g1263 ( n990 , n635 , n1340 );
    nor g1264 ( n1593 , n997 , n1341 );
    and g1265 ( n1344 , n1426 , n248 );
    and g1266 ( n344 , n100 , n1724 );
    not g1267 ( n563 , n1560 );
    not g1268 ( n926 , n805 );
    not g1269 ( n1407 , n149 );
    not g1270 ( n1187 , n42 );
    and g1271 ( n913 , n1101 , n1556 );
    xor g1272 ( n1241 , n21 , n327 );
    not g1273 ( n1064 , n343 );
    and g1274 ( n1615 , n612 , n980 );
    or g1275 ( n1114 , n1087 , n432 );
    or g1276 ( n188 , n1635 , n543 );
    or g1277 ( n1633 , n233 , n998 );
    or g1278 ( n1648 , n1679 , n279 );
    or g1279 ( n497 , n1051 , n1050 );
    or g1280 ( n193 , n657 , n109 );
    xnor g1281 ( n1150 , n1595 , n307 );
    nor g1282 ( n759 , n417 , n1494 );
    and g1283 ( n591 , n1030 , n318 );
    or g1284 ( n322 , n1182 , n398 );
    and g1285 ( n847 , n803 , n1195 );
    and g1286 ( n1361 , n328 , n524 );
    not g1287 ( n1623 , n1284 );
    or g1288 ( n515 , n1385 , n57 );
    nor g1289 ( n754 , n582 , n540 );
    not g1290 ( n1657 , n1280 );
    not g1291 ( n115 , n1742 );
    or g1292 ( n850 , n519 , n996 );
    not g1293 ( n1548 , n1376 );
    or g1294 ( n156 , n148 , n305 );
    nor g1295 ( n283 , n687 , n364 );
    not g1296 ( n92 , n450 );
    not g1297 ( n1071 , n56 );
    not g1298 ( n1446 , n885 );
    or g1299 ( n167 , n508 , n92 );
    or g1300 ( n1149 , n519 , n155 );
    or g1301 ( n125 , n1526 , n440 );
    or g1302 ( n1083 , n1206 , n712 );
    nor g1303 ( n1474 , n857 , n1691 );
    or g1304 ( n1266 , n1559 , n12 );
    or g1305 ( n1415 , n48 , n276 );
    not g1306 ( n1043 , n630 );
    and g1307 ( n158 , n254 , n1147 );
    or g1308 ( n1647 , n1134 , n653 );
    not g1309 ( n373 , n260 );
    nor g1310 ( n1594 , n264 , n796 );
    or g1311 ( n392 , n1373 , n531 );
    nor g1312 ( n43 , n382 , n1052 );
    xnor g1313 ( n1306 , n723 , n1202 );
    xnor g1314 ( n1706 , n1049 , n564 );
    not g1315 ( n1395 , n84 );
    xnor g1316 ( n1677 , n928 , n823 );
    xnor g1317 ( n1124 , n103 , n1670 );
    xnor g1318 ( n1449 , n1711 , n1586 );
    not g1319 ( n1547 , n1147 );
    or g1320 ( n1180 , n15 , n1412 );
    not g1321 ( n530 , n1522 );
    buf g1322 ( n6 , 1'b0 );
    and g1323 ( n246 , n1709 , n1268 );
    or g1324 ( n891 , n1452 , n1453 );
    xnor g1325 ( n132 , n869 , n1179 );
    or g1326 ( n632 , n1330 , n1186 );
    xor g1327 ( n172 , n984 , n1322 );
    not g1328 ( n927 , n77 );
    not g1329 ( n96 , n1548 );
    xnor g1330 ( n1085 , n380 , n1560 );
    or g1331 ( n85 , n728 , n267 );
    xnor g1332 ( n551 , n1578 , n1134 );
    buf g1333 ( n350 , 1'b0 );
    and g1334 ( n1759 , n639 , n387 );
    xnor g1335 ( n678 , n1600 , n1676 );
    not g1336 ( n1476 , n157 );
    not g1337 ( n179 , n1528 );
    and g1338 ( n1405 , n1286 , n1526 );
    nor g1339 ( n1390 , n1409 , n1510 );
    xnor g1340 ( n965 , n1755 , n1088 );
    or g1341 ( n1660 , n1565 , n1130 );
    or g1342 ( n695 , n34 , n370 );
    nor g1343 ( n1118 , n913 , n1159 );
    and g1344 ( n1618 , n297 , n188 );
    or g1345 ( n1199 , n1233 , n890 );
    and g1346 ( n1568 , n1461 , n647 );
    not g1347 ( n1283 , n930 );
    and g1348 ( n1504 , n1516 , n742 );
    nor g1349 ( n454 , n644 , n1208 );
    and g1350 ( n597 , n394 , n1647 );
    xor g1351 ( n1354 , n701 , n684 );
    not g1352 ( n1525 , n1022 );
    not g1353 ( n768 , n1315 );
    not g1354 ( n379 , n741 );
    or g1355 ( n700 , n1296 , n1257 );
    not g1356 ( n469 , n1532 );
    or g1357 ( n53 , n1094 , n528 );
    xnor g1358 ( n1335 , n882 , n486 );
    buf g1359 ( n721 , n1759 );
    nor g1360 ( n1253 , n816 , n1260 );
    buf g1361 ( n290 , 1'b0 );
    nor g1362 ( n73 , n1285 , n96 );
    not g1363 ( n482 , n656 );
    not g1364 ( n238 , n1065 );
    not g1365 ( n1347 , n1549 );
    xnor g1366 ( n1013 , n1730 , n1513 );
    xnor g1367 ( n920 , n1060 , n524 );
    not g1368 ( n393 , n1299 );
    not g1369 ( n1585 , n1177 );
    nor g1370 ( n50 , n1364 , n155 );
    xor g1371 ( n686 , n298 , n1484 );
    not g1372 ( n600 , n1274 );
    not g1373 ( n1619 , n1147 );
    not g1374 ( n126 , n1134 );
    and g1375 ( n577 , n1047 , n411 );
    xor g1376 ( n1188 , n271 , n213 );
    or g1377 ( n1131 , n55 , n986 );
    nor g1378 ( n1588 , n1349 , n1226 );
    or g1379 ( n226 , n1530 , n303 );
    not g1380 ( n1551 , n1481 );
    nor g1381 ( n728 , n1313 , n644 );
    or g1382 ( n1487 , n601 , n1547 );
    nor g1383 ( n863 , n1455 , n1052 );
    or g1384 ( n971 , n1147 , n1313 );
    and g1385 ( n1370 , n733 , n80 );
    not g1386 ( n541 , n139 );
    not g1387 ( n35 , n690 );
    and g1388 ( n844 , n445 , n132 );
    and g1389 ( n1221 , n1680 , n1434 );
    xnor g1390 ( n1742 , n35 , n944 );
    xnor g1391 ( n1441 , n180 , n1380 );
    not g1392 ( n896 , n1561 );
    or g1393 ( n480 , n1477 , n771 );
    nor g1394 ( n1110 , n1245 , n444 );
    not g1395 ( n876 , n1 );
    or g1396 ( n1509 , n1293 , n820 );
    xnor g1397 ( n549 , n677 , n1640 );
    or g1398 ( n1231 , n1536 , n523 );
    not g1399 ( n90 , n703 );
    or g1400 ( n1229 , n665 , n115 );
    not g1401 ( n1123 , n554 );
    buf g1402 ( n652 , n1354 );
    not g1403 ( n1002 , n435 );
    not g1404 ( n1061 , n1299 );
    or g1405 ( n1000 , n1592 , n607 );
    or g1406 ( n1254 , n863 , n1713 );
    or g1407 ( n726 , n1626 , n1166 );
    or g1408 ( n1098 , n1364 , n787 );
    or g1409 ( n1176 , n75 , n650 );
    nor g1410 ( n1571 , n1611 , n1187 );
    or g1411 ( n578 , n1722 , n420 );
    and g1412 ( n335 , n422 , n1117 );
    xnor g1413 ( n1723 , n1526 , n77 );
    or g1414 ( n826 , n1538 , n690 );
    not g1415 ( n302 , n555 );
    not g1416 ( n952 , n202 );
    not g1417 ( n364 , n1115 );
    not g1418 ( n645 , n864 );
    not g1419 ( n866 , n1012 );
    xnor g1420 ( n1428 , n312 , n1494 );
    not g1421 ( n1689 , n1079 );
    not g1422 ( n1175 , n1061 );
    nor g1423 ( n967 , n979 , n643 );
    and g1424 ( n895 , n353 , n402 );
    and g1425 ( n681 , n1341 , n977 );
    and g1426 ( n354 , n1745 , n1134 );
    not g1427 ( n334 , n1353 );
    or g1428 ( n1028 , n993 , n38 );
    and g1429 ( n420 , n1254 , n1700 );
    not g1430 ( n676 , n530 );
    or g1431 ( n705 , n516 , n681 );
    and g1432 ( n878 , n1420 , n613 );
    xnor g1433 ( n273 , n1077 , n399 );
    or g1434 ( n1420 , n589 , n61 );
    not g1435 ( n783 , n380 );
    or g1436 ( n521 , n1536 , n918 );
    not g1437 ( n1477 , n1346 );
    or g1438 ( n1355 , n1631 , n1729 );
    or g1439 ( n685 , n249 , n667 );
    xnor g1440 ( n1204 , n249 , n1256 );
    xnor g1441 ( n1158 , n176 , n1142 );
    xnor g1442 ( n1219 , n23 , n1735 );
    xnor g1443 ( n1688 , n301 , n418 );
    or g1444 ( n689 , n1264 , n162 );
    or g1445 ( n1340 , n1590 , n62 );
    and g1446 ( n747 , n736 , n1231 );
    or g1447 ( n414 , n654 , n395 );
    not g1448 ( n1142 , n828 );
    or g1449 ( n1497 , n313 , n754 );
    xor g1450 ( n649 , n922 , n1386 );
    or g1451 ( n351 , n881 , n854 );
    not g1452 ( n1232 , n371 );
    or g1453 ( n470 , n1070 , n1325 );
    and g1454 ( n255 , n1000 , n853 );
    nor g1455 ( n1257 , n28 , n1088 );
    nor g1456 ( n1235 , n723 , n934 );
    buf g1457 ( n312 , n1300 );
    not g1458 ( n374 , n1497 );
    or g1459 ( n1379 , n1437 , n1651 );
    or g1460 ( n514 , n447 , n569 );
    xnor g1461 ( n1227 , n619 , n1387 );
    not g1462 ( n1489 , n1123 );
    nor g1463 ( n198 , n552 , n721 );
    not g1464 ( n1032 , n745 );
    or g1465 ( n1222 , n657 , n803 );
    or g1466 ( n908 , n1405 , n697 );
    not g1467 ( n113 , n1120 );
    or g1468 ( n951 , n1603 , n624 );
    not g1469 ( n175 , n915 );
    xnor g1470 ( n646 , n1148 , n1336 );
    xnor g1471 ( n1664 , n1489 , n1052 );
    not g1472 ( n1014 , n1186 );
    not g1473 ( n300 , n1313 );
    xor g1474 ( n616 , n1609 , n342 );
    xnor g1475 ( n1189 , n435 , n721 );
    or g1476 ( n225 , n812 , n1258 );
    or g1477 ( n736 , n1351 , n2 );
    not g1478 ( n918 , n1344 );
    or g1479 ( n787 , n850 , n1338 );
    not g1480 ( n542 , n1342 );
    xnor g1481 ( n101 , n531 , n1189 );
    and g1482 ( n782 , n1133 , n1627 );
    not g1483 ( n221 , n291 );
    xor g1484 ( n1744 , n885 , n591 );
    not g1485 ( n1208 , n1698 );
    and g1486 ( n1554 , n414 , n1033 );
    nor g1487 ( n788 , n412 , n1245 );
    xnor g1488 ( n1629 , n1319 , n864 );
    not g1489 ( n683 , n1665 );
    xnor g1490 ( n953 , n372 , n1280 );
    and g1491 ( n233 , n1034 , n1121 );
    xor g1492 ( n618 , n1123 , n1398 );
    xnor g1493 ( n14 , n154 , n1323 );
    not g1494 ( n1557 , n1075 );
    not g1495 ( n415 , n111 );
    not g1496 ( n757 , n1252 );
    xnor g1497 ( n1429 , n184 , n1245 );
    or g1498 ( n1671 , n1232 , n429 );
    xnor g1499 ( n1322 , n242 , n1749 );
    not g1500 ( n1590 , n845 );
    nor g1501 ( n1021 , n397 , n1022 );
    or g1502 ( n849 , n991 , n174 );
    not g1503 ( n1012 , n131 );
    or g1504 ( n1658 , n755 , n67 );
    not g1505 ( n58 , n360 );
    xnor g1506 ( n320 , n1146 , n1486 );
    xnor g1507 ( n189 , n526 , n309 );
    or g1508 ( n737 , n424 , n33 );
    or g1509 ( n1207 , n1686 , n502 );
    nor g1510 ( n1577 , n1692 , n1494 );
    or g1511 ( n613 , n1409 , n445 );
    not g1512 ( n560 , n438 );
    not g1513 ( n636 , n1262 );
    or g1514 ( n884 , n154 , n1550 );
    xnor g1515 ( n150 , n1584 , n1470 );
    not g1516 ( n1139 , n1104 );
    xnor g1517 ( n1435 , n227 , n130 );
    xnor g1518 ( n1252 , n492 , n1752 );
    and g1519 ( n930 , n1239 , n1035 );
    not g1520 ( n1286 , n1638 );
    xnor g1521 ( n1616 , n623 , n551 );
    not g1522 ( n462 , n911 );
    or g1523 ( n668 , n1690 , n921 );
    xnor g1524 ( n1270 , n108 , n14 );
    and g1525 ( n71 , n847 , n815 );
    and g1526 ( n1701 , n123 , n337 );
    or g1527 ( n752 , n1147 , n1456 );
    xnor g1528 ( n1365 , n425 , n1245 );
    xnor g1529 ( n1382 , n1090 , n532 );
    or g1530 ( n149 , n217 , n1016 );
    and g1531 ( n1749 , n681 , n516 );
    or g1532 ( n525 , n357 , n1500 );
    or g1533 ( n609 , n1413 , n1159 );
    or g1534 ( n799 , n840 , n881 );
    or g1535 ( n419 , n1397 , n1490 );
    not g1536 ( n1042 , n1496 );
    xnor g1537 ( n1160 , n1276 , n721 );
    not g1538 ( n1400 , n1572 );
    nor g1539 ( n1607 , n519 , n1740 );
    xor g1540 ( n256 , n1685 , n530 );
    or g1541 ( n1564 , n657 , n680 );
    not g1542 ( n1630 , n200 );
    xnor g1543 ( n1456 , n847 , n829 );
    or g1544 ( n1462 , n1636 , n813 );
    not g1545 ( n617 , n473 );
    not g1546 ( n1503 , n1315 );
    xnor g1547 ( n1762 , n1435 , n898 );
    not g1548 ( n1018 , n953 );
    or g1549 ( n1019 , n396 , n336 );
    or g1550 ( n959 , n883 , n88 );
    or g1551 ( n1457 , n988 , n517 );
    and g1552 ( n1045 , n142 , n959 );
    or g1553 ( n1291 , n831 , n974 );
    or g1554 ( n49 , n1235 , n252 );
    nor g1555 ( n413 , n593 , n1098 );
    xnor g1556 ( n796 , n666 , n774 );
    or g1557 ( n143 , n738 , n862 );
    not g1558 ( n495 , n1262 );
    and g1559 ( n633 , n984 , n1322 );
    xnor g1560 ( n1507 , n163 , n1428 );
    not g1561 ( n1357 , n244 );
    xnor g1562 ( n974 , n1249 , n725 );
    buf g1563 ( n661 , n673 );
    xnor g1564 ( n1608 , n96 , n349 );
    xnor g1565 ( n1066 , n956 , n231 );
    or g1566 ( n1712 , n1454 , n1045 );
    not g1567 ( n1679 , n902 );
    nor g1568 ( n370 , n1309 , n995 );
    xnor g1569 ( n538 , n416 , n651 );
    and g1570 ( n234 , n695 , n753 );
    or g1571 ( n1461 , n983 , n1563 );
    nor g1572 ( n622 , n1494 , n312 );
    or g1573 ( n1672 , n29 , n100 );
    and g1574 ( n1704 , n1669 , n1489 );
    nor g1575 ( n362 , n657 , n1205 );
    not g1576 ( n679 , n1595 );
    xnor g1577 ( n485 , n1356 , n11 );
    xnor g1578 ( n553 , n239 , n471 );
    not g1579 ( n308 , n1446 );
    not g1580 ( n1584 , n1742 );
    not g1581 ( n1091 , n997 );
    not g1582 ( n1539 , n806 );
    not g1583 ( n717 , n694 );
    not g1584 ( n1535 , n1371 );
    not g1585 ( n919 , n1711 );
    not g1586 ( n868 , n999 );
    not g1587 ( n196 , n169 );
    xnor g1588 ( n107 , n1490 , n39 );
    xnor g1589 ( n1439 , n189 , n1575 );
    not g1590 ( n1111 , n1542 );
    not g1591 ( n1748 , n4 );
    not g1592 ( n63 , n1334 );
    xnor g1593 ( n0 , n866 , n603 );
    not g1594 ( n406 , n661 );
    xnor g1595 ( n1029 , n332 , n649 );
    and g1596 ( n1512 , n1494 , n916 );
    not g1597 ( n507 , n1640 );
    or g1598 ( n1165 , n208 , n1288 );
    xnor g1599 ( n345 , n1063 , n658 );
    or g1600 ( n909 , n93 , n1028 );
    not g1601 ( n1418 , n774 );
    not g1602 ( n590 , n1469 );
    not g1603 ( n32 , n661 );
    xnor g1604 ( n1396 , n1727 , n483 );
    not g1605 ( n1143 , n115 );
    or g1606 ( n1126 , n276 , n861 );
    nor g1607 ( n357 , n1557 , n1027 );
    or g1608 ( n1634 , n1309 , n344 );
    xnor g1609 ( n277 , n246 , n1302 );
    or g1610 ( n433 , n1357 , n909 );
    or g1611 ( n1186 , n831 , n135 );
    xnor g1612 ( n200 , n577 , n1664 );
    xnor g1613 ( n449 , n323 , n872 );
    and g1614 ( n575 , n1747 , n1106 );
    xnor g1615 ( n1445 , n831 , n66 );
    nor g1616 ( n369 , n1010 , n165 );
    or g1617 ( n1709 , n1292 , n1521 );
    and g1618 ( n61 , n743 , n323 );
    xor g1619 ( n1202 , n870 , n633 );
    nor g1620 ( n735 , n1473 , n1349 );
    xnor g1621 ( n1586 , n1136 , n1191 );
    nor g1622 ( n114 , n1147 , n3 );
    and g1623 ( n833 , n1457 , n514 );
    xnor g1624 ( n343 , n1648 , n547 );
    not g1625 ( n1274 , n171 );
    or g1626 ( n1023 , n1185 , n1615 );
    xnor g1627 ( n627 , n497 , n356 );
    xnor g1628 ( n16 , n744 , n1245 );
    not g1629 ( n1275 , n1721 );
    xnor g1630 ( n1218 , n324 , n600 );
    not g1631 ( n605 , n1703 );
    nor g1632 ( n1037 , n1244 , n466 );
    or g1633 ( n1250 , n914 , n153 );
    nor g1634 ( n1388 , n845 , n719 );
    not g1635 ( n316 , n175 );
    not g1636 ( n387 , n690 );
    not g1637 ( n1360 , n1384 );
    not g1638 ( n54 , n818 );
    not g1639 ( n13 , n729 );
    or g1640 ( n337 , n583 , n1430 );
    buf g1641 ( n1654 , 1'b0 );
    not g1642 ( n664 , n1084 );
    not g1643 ( n398 , n451 );
    or g1644 ( n1212 , n949 , n763 );
    not g1645 ( n1195 , n680 );
    not g1646 ( n1475 , n1275 );
    not g1647 ( n887 , n216 );
    and g1648 ( n1166 , n1201 , n269 );
    and g1649 ( n907 , n1153 , n1289 );
    or g1650 ( n163 , n429 , n1701 );
    not g1651 ( n1119 , n1134 );
    and g1652 ( n180 , n95 , n97 );
    buf g1653 ( n1447 , 1'b0 );
    xnor g1654 ( n258 , n907 , n1029 );
    nor g1655 ( n1596 , n126 , n1066 );
    xnor g1656 ( n1267 , n571 , n1396 );
    not g1657 ( n1016 , n168 );
    not g1658 ( n1502 , n680 );
    not g1659 ( n1732 , n422 );
    xnor g1660 ( n1065 , n44 , n168 );
    xnor g1661 ( n872 , n113 , n661 );
    not g1662 ( n1182 , n204 );
    not g1663 ( n1008 , n1476 );
    and g1664 ( n589 , n1493 , n661 );
    or g1665 ( n764 , n1175 , n1291 );
    not g1666 ( n42 , n941 );
    or g1667 ( n1448 , n1552 , n1155 );
    xnor g1668 ( n1358 , n196 , n1001 );
    not g1669 ( n1350 , n1003 );
    not g1670 ( n191 , n1107 );
    nor g1671 ( n261 , n586 , n194 );
    not g1672 ( n1315 , n549 );
    or g1673 ( n513 , n1593 , n1460 );
    or g1674 ( n1001 , n476 , n1744 );
endmodule
