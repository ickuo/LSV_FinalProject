// Benchmark "top" written by ABC on Sun Dec 21 18:10:42 2025

module top ( 
    n9, n22, n103, n124, n287, n353, n389, n401, n411, n443, n469, n497,
    n499, n510, n603, n761, n767, n772, n817, n834, n854, n937, n951,
    n1007, n1084, n1165, n1198, n1231, n1302, n1307, n1364, n1392, n1636,
    n1650, n1709, n1724, n1757, n1912, n1916, n1982, n2057, n2068, n2174,
    n2252, n2295, n2339, n2341, n2458, n2482, n2498, n2590, n2592, n2666,
    n2737, n2758, n2771, n2777, n2882, n3006, n3076, n3085, n3112, n3130,
    n3178, n3311, n3409, n3591, n3641, n3669, n3677, n3769, n3815, n3832,
    n4006, n4075, n4114, n4122, n4141, n4330, n4335, n4357, n4382, n4419,
    n4452, n4470, n4743, n4748, n4862, n4964, n4998, n5031, n5065, n5167,
    n5189, n5214, n5320, n5356, n5427, n5470, n5536, n5548, n5568, n5586,
    n5671, n5684, n5715, n5729, n5758, n5801, n5884, n5920, n5962, n5969,
    n6023, n6085, n6149, n6168, n6333, n6392, n6409, n6655, n6668, n6818,
    n6826, n6843, n6937, n7061, n7113, n7161, n7374, n7411, n7529, n7659,
    n7715, n7720, n7729, n7772, n7812, n7974, n8139, n8163, n8183, n8228,
    n8230, n8233, n8290, n8308, n8332, n8466, n8468, n8506, n8522, n8716,
    n8768, n8820, n8859, n8860, n8940, n9041, n9093, n9187, n9216, n9300,
    n9353, n9475, n9528, n9531, n9570, n9591, n9620, n9669, n9732, n9747,
    n9846, n9887, n9906, n9915, n10063, n10113, n10122, n10142, n10162,
    n10168, n10408, n10416, n10451, n10522, n10560, n10594, n10606, n10642,
    n10657, n10770, n10805, n10866, n10874, n10908, n11030, n11058, n11061,
    n11109, n11111, n11180, n11222, n11236, n11324, n11350, n11396, n11411,
    n11429, n11488, n11537, n11574, n11634, n11665, n11734, n11835, n11891,
    n12003, n12065, n12263, n12284, n12289, n12306, n12348, n12352, n12372,
    n12408, n12482, n12579, n12592, n12605, n12651, n12693, n12750, n12853,
    n12912, n12965, n13058, n13060, n13201,
    n134, n201, n211, n358, n370, n396, n460, n537, n573, n728, n758, n762,
    n777, n800, n831, n846, n922, n927, n985, n1097, n1112, n1181, n1401,
    n1487, n1561, n1806, n1860, n1937, n2061, n2190, n2235, n2549, n2709,
    n2805, n2904, n2934, n3262, n3323, n3362, n3748, n3790, n3946, n4059,
    n4202, n4553, n4777, n4824, n4864, n5003, n5060, n5364, n5549, n5557,
    n5609, n5882, n6019, n6103, n6109, n6297, n6301, n6434, n6586, n6683,
    n6862, n7034, n7111, n7132, n7241, n7553, n7582, n7687, n7755, n7790,
    n7858, n7860, n7968, n8172, n8219, n8265, n8336, n8516, n8701, n9100,
    n9329, n9866, n9872, n10101, n10243, n10453, n10524, n10628, n10736,
    n10797, n11057, n11077, n11140, n11147, n11252, n11264, n11484, n11667,
    n11732, n11778, n11792, n11879, n11882, n11895, n12059, n12067, n12187,
    n12334, n12406, n12463, n12503, n12515, n12616, n12839, n12968, n13002,
    n13035  );
  input  n9, n22, n103, n124, n287, n353, n389, n401, n411, n443, n469,
    n497, n499, n510, n603, n761, n767, n772, n817, n834, n854, n937, n951,
    n1007, n1084, n1165, n1198, n1231, n1302, n1307, n1364, n1392, n1636,
    n1650, n1709, n1724, n1757, n1912, n1916, n1982, n2057, n2068, n2174,
    n2252, n2295, n2339, n2341, n2458, n2482, n2498, n2590, n2592, n2666,
    n2737, n2758, n2771, n2777, n2882, n3006, n3076, n3085, n3112, n3130,
    n3178, n3311, n3409, n3591, n3641, n3669, n3677, n3769, n3815, n3832,
    n4006, n4075, n4114, n4122, n4141, n4330, n4335, n4357, n4382, n4419,
    n4452, n4470, n4743, n4748, n4862, n4964, n4998, n5031, n5065, n5167,
    n5189, n5214, n5320, n5356, n5427, n5470, n5536, n5548, n5568, n5586,
    n5671, n5684, n5715, n5729, n5758, n5801, n5884, n5920, n5962, n5969,
    n6023, n6085, n6149, n6168, n6333, n6392, n6409, n6655, n6668, n6818,
    n6826, n6843, n6937, n7061, n7113, n7161, n7374, n7411, n7529, n7659,
    n7715, n7720, n7729, n7772, n7812, n7974, n8139, n8163, n8183, n8228,
    n8230, n8233, n8290, n8308, n8332, n8466, n8468, n8506, n8522, n8716,
    n8768, n8820, n8859, n8860, n8940, n9041, n9093, n9187, n9216, n9300,
    n9353, n9475, n9528, n9531, n9570, n9591, n9620, n9669, n9732, n9747,
    n9846, n9887, n9906, n9915, n10063, n10113, n10122, n10142, n10162,
    n10168, n10408, n10416, n10451, n10522, n10560, n10594, n10606, n10642,
    n10657, n10770, n10805, n10866, n10874, n10908, n11030, n11058, n11061,
    n11109, n11111, n11180, n11222, n11236, n11324, n11350, n11396, n11411,
    n11429, n11488, n11537, n11574, n11634, n11665, n11734, n11835, n11891,
    n12003, n12065, n12263, n12284, n12289, n12306, n12348, n12352, n12372,
    n12408, n12482, n12579, n12592, n12605, n12651, n12693, n12750, n12853,
    n12912, n12965, n13058, n13060, n13201;
  output n134, n201, n211, n358, n370, n396, n460, n537, n573, n728, n758,
    n762, n777, n800, n831, n846, n922, n927, n985, n1097, n1112, n1181,
    n1401, n1487, n1561, n1806, n1860, n1937, n2061, n2190, n2235, n2549,
    n2709, n2805, n2904, n2934, n3262, n3323, n3362, n3748, n3790, n3946,
    n4059, n4202, n4553, n4777, n4824, n4864, n5003, n5060, n5364, n5549,
    n5557, n5609, n5882, n6019, n6103, n6109, n6297, n6301, n6434, n6586,
    n6683, n6862, n7034, n7111, n7132, n7241, n7553, n7582, n7687, n7755,
    n7790, n7858, n7860, n7968, n8172, n8219, n8265, n8336, n8516, n8701,
    n9100, n9329, n9866, n9872, n10101, n10243, n10453, n10524, n10628,
    n10736, n10797, n11057, n11077, n11140, n11147, n11252, n11264, n11484,
    n11667, n11732, n11778, n11792, n11879, n11882, n11895, n12059, n12067,
    n12187, n12334, n12406, n12463, n12503, n12515, n12616, n12839, n12968,
    n13002, n13035;
  wire new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370_1, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389_1,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396_1,
    new_n397, new_n398, new_n399, new_n400, new_n401_1, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411_1, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443_1, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460_1, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497_1, new_n498, new_n499_1, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510_1, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537_1, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573_1, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603_1, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728_1, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758_1, new_n759, new_n760,
    new_n761_1, new_n762_1, new_n763, new_n764, new_n765, new_n766,
    new_n767_1, new_n768, new_n769, new_n770, new_n771, new_n772_1,
    new_n773, new_n774, new_n775, new_n776, new_n777_1, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800_1,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817_1, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831_1, new_n832, new_n833, new_n834_1,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846_1, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854_1, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922_1, new_n923, new_n924, new_n925,
    new_n926, new_n927_1, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937_1, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951_1, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985_1, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007_1,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084_1, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1097_1,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112_1, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165_1, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181_1,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198_1, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231_1, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302_1, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307_1,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338, new_n1339, new_n1340, new_n1341, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347, new_n1348, new_n1349,
    new_n1350, new_n1351, new_n1352, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363, new_n1364_1, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369, new_n1370, new_n1371, new_n1372, new_n1373,
    new_n1374, new_n1375, new_n1376, new_n1377, new_n1378, new_n1379,
    new_n1380, new_n1381, new_n1382, new_n1383, new_n1384, new_n1385,
    new_n1386, new_n1387, new_n1388, new_n1389, new_n1390, new_n1391,
    new_n1392_1, new_n1393, new_n1394, new_n1395, new_n1396, new_n1397,
    new_n1398, new_n1399, new_n1400, new_n1401_1, new_n1402, new_n1403,
    new_n1404, new_n1405, new_n1406, new_n1407, new_n1408, new_n1409,
    new_n1410, new_n1411, new_n1412, new_n1413, new_n1414, new_n1415,
    new_n1416, new_n1417, new_n1418, new_n1419, new_n1420, new_n1421,
    new_n1422, new_n1423, new_n1424, new_n1425, new_n1426, new_n1427,
    new_n1428, new_n1429, new_n1430, new_n1431, new_n1432, new_n1433,
    new_n1434, new_n1435, new_n1436, new_n1437, new_n1438, new_n1439,
    new_n1440, new_n1441, new_n1442, new_n1443, new_n1444, new_n1445,
    new_n1446, new_n1447, new_n1448, new_n1449, new_n1450, new_n1451,
    new_n1452, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1467, new_n1468, new_n1469, new_n1470, new_n1471,
    new_n1472, new_n1473, new_n1474, new_n1475, new_n1476, new_n1477,
    new_n1478, new_n1479, new_n1480, new_n1481, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1486, new_n1487_1, new_n1488, new_n1489,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1494, new_n1495,
    new_n1496, new_n1497, new_n1498, new_n1499, new_n1500, new_n1501,
    new_n1502, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507,
    new_n1508, new_n1509, new_n1510, new_n1511, new_n1512, new_n1513,
    new_n1514, new_n1515, new_n1516, new_n1517, new_n1518, new_n1519,
    new_n1520, new_n1521, new_n1522, new_n1523, new_n1524, new_n1525,
    new_n1526, new_n1527, new_n1528, new_n1529, new_n1530, new_n1531,
    new_n1532, new_n1533, new_n1534, new_n1535, new_n1536, new_n1537,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1558, new_n1559, new_n1560, new_n1561_1,
    new_n1562, new_n1563, new_n1564, new_n1565, new_n1566, new_n1567,
    new_n1568, new_n1569, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1590, new_n1591,
    new_n1592, new_n1593, new_n1594, new_n1595, new_n1596, new_n1597,
    new_n1598, new_n1599, new_n1600, new_n1601, new_n1602, new_n1603,
    new_n1604, new_n1605, new_n1606, new_n1607, new_n1608, new_n1609,
    new_n1610, new_n1611, new_n1612, new_n1613, new_n1614, new_n1615,
    new_n1616, new_n1617, new_n1618, new_n1619, new_n1620, new_n1621,
    new_n1622, new_n1623, new_n1624, new_n1625, new_n1626, new_n1627,
    new_n1628, new_n1629, new_n1630, new_n1631, new_n1632, new_n1633,
    new_n1634, new_n1635, new_n1636_1, new_n1637, new_n1638, new_n1639,
    new_n1640, new_n1641, new_n1642, new_n1643, new_n1644, new_n1645,
    new_n1646, new_n1647, new_n1648, new_n1649, new_n1650_1, new_n1651,
    new_n1652, new_n1653, new_n1654, new_n1655, new_n1656, new_n1657,
    new_n1658, new_n1659, new_n1660, new_n1661, new_n1662, new_n1663,
    new_n1664, new_n1665, new_n1666, new_n1667, new_n1668, new_n1669,
    new_n1670, new_n1671, new_n1672, new_n1673, new_n1674, new_n1675,
    new_n1676, new_n1677, new_n1678, new_n1679, new_n1680, new_n1681,
    new_n1682, new_n1683, new_n1684, new_n1685, new_n1686, new_n1687,
    new_n1688, new_n1689, new_n1690, new_n1691, new_n1692, new_n1693,
    new_n1694, new_n1695, new_n1696, new_n1697, new_n1698, new_n1699,
    new_n1700, new_n1701, new_n1702, new_n1703, new_n1704, new_n1705,
    new_n1706, new_n1707, new_n1708, new_n1709_1, new_n1710, new_n1711,
    new_n1712, new_n1713, new_n1714, new_n1715, new_n1716, new_n1717,
    new_n1718, new_n1719, new_n1720, new_n1721, new_n1722, new_n1723,
    new_n1724_1, new_n1725, new_n1726, new_n1727, new_n1728, new_n1729,
    new_n1730, new_n1731, new_n1732, new_n1733, new_n1734, new_n1735,
    new_n1736, new_n1737, new_n1738, new_n1739, new_n1740, new_n1741,
    new_n1742, new_n1743, new_n1744, new_n1745, new_n1746, new_n1747,
    new_n1748, new_n1749, new_n1750, new_n1751, new_n1752, new_n1753,
    new_n1754, new_n1755, new_n1756, new_n1757_1, new_n1758, new_n1759,
    new_n1760, new_n1761, new_n1762, new_n1763, new_n1764, new_n1765,
    new_n1766, new_n1767, new_n1768, new_n1769, new_n1770, new_n1771,
    new_n1772, new_n1773, new_n1774, new_n1775, new_n1776, new_n1777,
    new_n1778, new_n1779, new_n1780, new_n1781, new_n1782, new_n1783,
    new_n1784, new_n1785, new_n1786, new_n1787, new_n1788, new_n1789,
    new_n1790, new_n1791, new_n1792, new_n1793, new_n1794, new_n1795,
    new_n1796, new_n1797, new_n1798, new_n1799, new_n1800, new_n1801,
    new_n1802, new_n1803, new_n1804, new_n1805, new_n1806_1, new_n1807,
    new_n1808, new_n1809, new_n1810, new_n1811, new_n1812, new_n1813,
    new_n1814, new_n1815, new_n1816, new_n1817, new_n1818, new_n1819,
    new_n1820, new_n1821, new_n1822, new_n1823, new_n1824, new_n1825,
    new_n1826, new_n1827, new_n1828, new_n1829, new_n1830, new_n1831,
    new_n1832, new_n1833, new_n1834, new_n1835, new_n1836, new_n1837,
    new_n1838, new_n1839, new_n1840, new_n1841, new_n1842, new_n1843,
    new_n1844, new_n1845, new_n1846, new_n1847, new_n1848, new_n1849,
    new_n1850, new_n1851, new_n1852, new_n1853, new_n1854, new_n1855,
    new_n1856, new_n1857, new_n1858, new_n1859, new_n1860_1, new_n1861,
    new_n1862, new_n1863, new_n1864, new_n1865, new_n1866, new_n1867,
    new_n1868, new_n1869, new_n1870, new_n1871, new_n1872, new_n1873,
    new_n1874, new_n1875, new_n1876, new_n1877, new_n1878, new_n1879,
    new_n1880, new_n1881, new_n1882, new_n1883, new_n1884, new_n1885,
    new_n1886, new_n1887, new_n1888, new_n1889, new_n1890, new_n1891,
    new_n1892, new_n1893, new_n1894, new_n1895, new_n1896, new_n1897,
    new_n1898, new_n1899, new_n1900, new_n1901, new_n1902, new_n1903,
    new_n1904, new_n1905, new_n1906, new_n1907, new_n1908, new_n1909,
    new_n1910, new_n1911, new_n1912_1, new_n1913, new_n1914, new_n1915,
    new_n1916_1, new_n1917, new_n1918, new_n1919, new_n1920, new_n1921,
    new_n1922, new_n1923, new_n1924, new_n1925, new_n1926, new_n1927,
    new_n1928, new_n1929, new_n1930, new_n1931, new_n1932, new_n1933,
    new_n1934, new_n1935, new_n1936, new_n1937_1, new_n1938, new_n1939,
    new_n1940, new_n1941, new_n1942, new_n1943, new_n1944, new_n1945,
    new_n1946, new_n1947, new_n1948, new_n1949, new_n1950, new_n1951,
    new_n1952, new_n1953, new_n1954, new_n1955, new_n1956, new_n1957,
    new_n1958, new_n1959, new_n1960, new_n1961, new_n1962, new_n1963,
    new_n1964, new_n1965, new_n1966, new_n1967, new_n1968, new_n1969,
    new_n1970, new_n1971, new_n1972, new_n1973, new_n1974, new_n1975,
    new_n1976, new_n1977, new_n1978, new_n1979, new_n1980, new_n1981,
    new_n1982_1, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2006,
    new_n2007, new_n2008, new_n2009, new_n2010, new_n2011, new_n2012,
    new_n2013, new_n2014, new_n2015, new_n2016, new_n2017, new_n2018,
    new_n2019, new_n2020, new_n2021, new_n2022, new_n2023, new_n2024,
    new_n2025, new_n2026, new_n2027, new_n2028, new_n2029, new_n2030,
    new_n2031, new_n2032, new_n2033, new_n2034, new_n2035, new_n2036,
    new_n2037, new_n2038, new_n2039, new_n2040, new_n2041, new_n2042,
    new_n2043, new_n2044, new_n2045, new_n2046, new_n2047, new_n2048,
    new_n2049, new_n2050, new_n2051, new_n2052, new_n2053, new_n2054,
    new_n2055, new_n2056, new_n2057_1, new_n2058, new_n2059, new_n2060,
    new_n2061_1, new_n2062, new_n2063, new_n2064, new_n2065, new_n2066,
    new_n2067, new_n2068_1, new_n2069, new_n2070, new_n2071, new_n2072,
    new_n2073, new_n2074, new_n2075, new_n2076, new_n2077, new_n2078,
    new_n2079, new_n2080, new_n2081, new_n2082, new_n2083, new_n2084,
    new_n2085, new_n2086, new_n2087, new_n2088, new_n2089, new_n2090,
    new_n2091, new_n2092, new_n2093, new_n2094, new_n2095, new_n2096,
    new_n2097, new_n2098, new_n2099, new_n2100, new_n2101, new_n2102,
    new_n2103, new_n2104, new_n2105, new_n2106, new_n2107, new_n2108,
    new_n2109, new_n2110, new_n2111, new_n2112, new_n2113, new_n2114,
    new_n2115, new_n2116, new_n2117, new_n2118, new_n2119, new_n2120,
    new_n2121, new_n2122, new_n2123, new_n2124, new_n2125, new_n2126,
    new_n2127, new_n2128, new_n2129, new_n2130, new_n2131, new_n2132,
    new_n2133, new_n2134, new_n2135, new_n2136, new_n2137, new_n2138,
    new_n2139, new_n2140, new_n2141, new_n2142, new_n2143, new_n2144,
    new_n2145, new_n2146, new_n2147, new_n2148, new_n2149, new_n2150,
    new_n2151, new_n2152, new_n2153, new_n2154, new_n2155, new_n2156,
    new_n2157, new_n2158, new_n2159, new_n2160, new_n2161, new_n2162,
    new_n2163, new_n2164, new_n2165, new_n2166, new_n2167, new_n2168,
    new_n2169, new_n2170, new_n2171, new_n2172, new_n2173, new_n2174_1,
    new_n2175, new_n2176, new_n2177, new_n2178, new_n2179, new_n2180,
    new_n2181, new_n2182, new_n2183, new_n2184, new_n2185, new_n2186,
    new_n2187, new_n2188, new_n2189, new_n2190_1, new_n2191, new_n2192,
    new_n2193, new_n2194, new_n2195, new_n2196, new_n2197, new_n2198,
    new_n2199, new_n2200, new_n2201, new_n2202, new_n2203, new_n2204,
    new_n2205, new_n2206, new_n2207, new_n2208, new_n2209, new_n2210,
    new_n2211, new_n2212, new_n2213, new_n2214, new_n2215, new_n2216,
    new_n2217, new_n2218, new_n2219, new_n2220, new_n2221, new_n2222,
    new_n2223, new_n2224, new_n2225, new_n2226, new_n2227, new_n2228,
    new_n2229, new_n2230, new_n2231, new_n2232, new_n2233, new_n2234,
    new_n2235_1, new_n2236, new_n2237, new_n2238, new_n2239, new_n2240,
    new_n2241, new_n2242, new_n2243, new_n2244, new_n2245, new_n2246,
    new_n2247, new_n2248, new_n2249, new_n2250, new_n2251, new_n2252_1,
    new_n2253, new_n2254, new_n2255, new_n2256, new_n2257, new_n2258,
    new_n2259, new_n2260, new_n2261, new_n2262, new_n2263, new_n2264,
    new_n2265, new_n2266, new_n2267, new_n2268, new_n2269, new_n2270,
    new_n2271, new_n2272, new_n2273, new_n2274, new_n2275, new_n2276,
    new_n2277, new_n2278, new_n2279, new_n2280, new_n2281, new_n2282,
    new_n2283, new_n2284, new_n2285, new_n2286, new_n2287, new_n2288,
    new_n2289, new_n2290, new_n2291, new_n2292, new_n2293, new_n2294,
    new_n2295_1, new_n2296, new_n2297, new_n2298, new_n2299, new_n2300,
    new_n2301, new_n2302, new_n2303, new_n2304, new_n2305, new_n2306,
    new_n2307, new_n2308, new_n2309, new_n2310, new_n2311, new_n2312,
    new_n2313, new_n2314, new_n2315, new_n2316, new_n2317, new_n2318,
    new_n2319, new_n2320, new_n2321, new_n2322, new_n2323, new_n2324,
    new_n2325, new_n2326, new_n2327, new_n2328, new_n2329, new_n2330,
    new_n2331, new_n2332, new_n2333, new_n2334, new_n2335, new_n2336,
    new_n2337, new_n2338, new_n2339_1, new_n2340, new_n2341_1, new_n2342,
    new_n2343, new_n2344, new_n2345, new_n2346, new_n2347, new_n2348,
    new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361, new_n2362, new_n2363, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416, new_n2417, new_n2418, new_n2419, new_n2420,
    new_n2421, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440, new_n2441, new_n2442, new_n2443, new_n2444,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458_1, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482_1, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498_1,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513, new_n2514, new_n2515, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547, new_n2548, new_n2549_1, new_n2550, new_n2551, new_n2552,
    new_n2553, new_n2554, new_n2555, new_n2556, new_n2557, new_n2558,
    new_n2559, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572, new_n2573, new_n2574, new_n2575, new_n2576,
    new_n2577, new_n2578, new_n2579, new_n2580, new_n2581, new_n2582,
    new_n2583, new_n2584, new_n2585, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590_1, new_n2591, new_n2592_1, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624,
    new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666_1,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696,
    new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702,
    new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708,
    new_n2709_1, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2720,
    new_n2721, new_n2722, new_n2723, new_n2724, new_n2725, new_n2726,
    new_n2727, new_n2728, new_n2729, new_n2730, new_n2731, new_n2732,
    new_n2733, new_n2734, new_n2735, new_n2736, new_n2737_1, new_n2738,
    new_n2739, new_n2740, new_n2741, new_n2742, new_n2743, new_n2744,
    new_n2745, new_n2746, new_n2747, new_n2748, new_n2749, new_n2750,
    new_n2751, new_n2752, new_n2753, new_n2754, new_n2755, new_n2756,
    new_n2757, new_n2758_1, new_n2759, new_n2760, new_n2761, new_n2762,
    new_n2763, new_n2764, new_n2765, new_n2766, new_n2767, new_n2768,
    new_n2769, new_n2770, new_n2771_1, new_n2772, new_n2773, new_n2774,
    new_n2775, new_n2776, new_n2777_1, new_n2778, new_n2779, new_n2780,
    new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792,
    new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2798,
    new_n2799, new_n2800, new_n2801, new_n2802, new_n2803, new_n2804,
    new_n2805_1, new_n2806, new_n2807, new_n2808, new_n2809, new_n2810,
    new_n2811, new_n2812, new_n2813, new_n2814, new_n2815, new_n2816,
    new_n2817, new_n2818, new_n2819, new_n2820, new_n2821, new_n2822,
    new_n2823, new_n2824, new_n2825, new_n2826, new_n2827, new_n2828,
    new_n2829, new_n2830, new_n2831, new_n2832, new_n2833, new_n2834,
    new_n2835, new_n2836, new_n2837, new_n2838, new_n2839, new_n2840,
    new_n2841, new_n2842, new_n2843, new_n2844, new_n2845, new_n2846,
    new_n2847, new_n2848, new_n2849, new_n2850, new_n2851, new_n2852,
    new_n2853, new_n2854, new_n2855, new_n2856, new_n2857, new_n2858,
    new_n2859, new_n2860, new_n2861, new_n2862, new_n2863, new_n2864,
    new_n2865, new_n2866, new_n2867, new_n2868, new_n2869, new_n2871,
    new_n2872, new_n2873, new_n2874, new_n2875, new_n2876, new_n2877,
    new_n2878, new_n2879, new_n2880, new_n2881, new_n2882_1, new_n2883,
    new_n2884, new_n2885, new_n2886, new_n2887, new_n2888, new_n2889,
    new_n2890, new_n2891, new_n2892, new_n2893, new_n2894, new_n2895,
    new_n2896, new_n2897, new_n2898, new_n2899, new_n2900, new_n2901,
    new_n2902, new_n2903, new_n2904_1, new_n2905, new_n2906, new_n2907,
    new_n2908, new_n2909, new_n2910, new_n2911, new_n2912, new_n2913,
    new_n2914, new_n2915, new_n2916, new_n2917, new_n2918, new_n2919,
    new_n2920, new_n2921, new_n2922, new_n2923, new_n2924, new_n2925,
    new_n2926, new_n2927, new_n2928, new_n2929, new_n2930, new_n2931,
    new_n2932, new_n2933, new_n2934_1, new_n2935, new_n2936, new_n2937,
    new_n2938, new_n2939, new_n2940, new_n2941, new_n2942, new_n2943,
    new_n2944, new_n2945, new_n2946, new_n2947, new_n2948, new_n2949,
    new_n2950, new_n2951, new_n2952, new_n2953, new_n2954, new_n2955,
    new_n2956, new_n2957, new_n2958, new_n2959, new_n2960, new_n2961,
    new_n2962, new_n2963, new_n2964, new_n2965, new_n2966, new_n2967,
    new_n2968, new_n2969, new_n2970, new_n2971, new_n2972, new_n2973,
    new_n2974, new_n2975, new_n2976, new_n2977, new_n2978, new_n2979,
    new_n2980, new_n2981, new_n2982, new_n2983, new_n2984, new_n2985,
    new_n2986, new_n2987, new_n2988, new_n2989, new_n2990, new_n2991,
    new_n2992, new_n2993, new_n2994, new_n2995, new_n2996, new_n2997,
    new_n2998, new_n2999, new_n3000, new_n3001, new_n3002, new_n3003,
    new_n3004, new_n3005, new_n3006_1, new_n3007, new_n3008, new_n3009,
    new_n3010, new_n3011, new_n3012, new_n3013, new_n3014, new_n3015,
    new_n3016, new_n3017, new_n3018, new_n3019, new_n3020, new_n3021,
    new_n3022, new_n3023, new_n3024, new_n3025, new_n3026, new_n3027,
    new_n3028, new_n3029, new_n3030, new_n3031, new_n3032, new_n3033,
    new_n3034, new_n3035, new_n3036, new_n3037, new_n3038, new_n3039,
    new_n3040, new_n3041, new_n3042, new_n3043, new_n3044, new_n3045,
    new_n3046, new_n3047, new_n3048, new_n3049, new_n3050, new_n3051,
    new_n3052, new_n3053, new_n3054, new_n3055, new_n3056, new_n3057,
    new_n3058, new_n3059, new_n3060, new_n3061, new_n3062, new_n3063,
    new_n3064, new_n3065, new_n3066, new_n3067, new_n3068, new_n3069,
    new_n3070, new_n3071, new_n3072, new_n3073, new_n3074, new_n3075,
    new_n3076_1, new_n3077, new_n3078, new_n3079, new_n3080, new_n3081,
    new_n3082, new_n3083, new_n3084, new_n3085_1, new_n3086, new_n3087,
    new_n3088, new_n3089, new_n3090, new_n3091, new_n3092, new_n3093,
    new_n3094, new_n3095, new_n3096, new_n3097, new_n3098, new_n3099,
    new_n3100, new_n3101, new_n3102, new_n3103, new_n3104, new_n3105,
    new_n3106, new_n3107, new_n3108, new_n3109, new_n3110, new_n3111,
    new_n3112_1, new_n3113, new_n3114, new_n3115, new_n3116, new_n3117,
    new_n3118, new_n3119, new_n3120, new_n3121, new_n3122, new_n3123,
    new_n3124, new_n3125, new_n3126, new_n3127, new_n3128, new_n3129,
    new_n3130_1, new_n3131, new_n3132, new_n3133, new_n3134, new_n3135,
    new_n3136, new_n3137, new_n3138, new_n3139, new_n3140, new_n3141,
    new_n3142, new_n3143, new_n3144, new_n3145, new_n3146, new_n3147,
    new_n3148, new_n3149, new_n3150, new_n3151, new_n3152, new_n3153,
    new_n3154, new_n3155, new_n3156, new_n3157, new_n3158, new_n3159,
    new_n3160, new_n3161, new_n3162, new_n3163, new_n3164, new_n3165,
    new_n3166, new_n3167, new_n3168, new_n3169, new_n3170, new_n3171,
    new_n3172, new_n3173, new_n3174, new_n3175, new_n3176, new_n3177,
    new_n3178_1, new_n3179, new_n3180, new_n3181, new_n3182, new_n3183,
    new_n3184, new_n3185, new_n3186, new_n3187, new_n3188, new_n3189,
    new_n3190, new_n3191, new_n3192, new_n3193, new_n3194, new_n3195,
    new_n3196, new_n3197, new_n3198, new_n3199, new_n3200, new_n3201,
    new_n3202, new_n3203, new_n3204, new_n3205, new_n3206, new_n3207,
    new_n3208, new_n3209, new_n3210, new_n3211, new_n3212, new_n3213,
    new_n3214, new_n3215, new_n3216, new_n3217, new_n3218, new_n3219,
    new_n3220, new_n3221, new_n3222, new_n3223, new_n3224, new_n3225,
    new_n3226, new_n3227, new_n3228, new_n3229, new_n3230, new_n3231,
    new_n3232, new_n3233, new_n3234, new_n3235, new_n3236, new_n3237,
    new_n3238, new_n3239, new_n3240, new_n3241, new_n3242, new_n3243,
    new_n3244, new_n3245, new_n3246, new_n3247, new_n3248, new_n3249,
    new_n3250, new_n3251, new_n3252, new_n3253, new_n3254, new_n3255,
    new_n3256, new_n3257, new_n3258, new_n3259, new_n3260, new_n3261,
    new_n3262_1, new_n3263, new_n3264, new_n3265, new_n3266, new_n3267,
    new_n3268, new_n3269, new_n3270, new_n3271, new_n3272, new_n3273,
    new_n3274, new_n3275, new_n3276, new_n3277, new_n3278, new_n3279,
    new_n3280, new_n3281, new_n3282, new_n3283, new_n3284, new_n3285,
    new_n3286, new_n3287, new_n3288, new_n3289, new_n3290, new_n3291,
    new_n3292, new_n3293, new_n3294, new_n3295, new_n3296, new_n3297,
    new_n3298, new_n3299, new_n3300, new_n3301, new_n3302, new_n3303,
    new_n3304, new_n3305, new_n3306, new_n3307, new_n3308, new_n3309,
    new_n3310, new_n3311_1, new_n3312, new_n3313, new_n3314, new_n3315,
    new_n3316, new_n3317, new_n3318, new_n3319, new_n3320, new_n3321,
    new_n3322, new_n3323_1, new_n3324, new_n3325, new_n3326, new_n3327,
    new_n3328, new_n3329, new_n3330, new_n3331, new_n3332, new_n3333,
    new_n3334, new_n3335, new_n3336, new_n3337, new_n3338, new_n3339,
    new_n3340, new_n3341, new_n3342, new_n3343, new_n3344, new_n3345,
    new_n3346, new_n3347, new_n3348, new_n3349, new_n3350, new_n3351,
    new_n3352, new_n3353, new_n3354, new_n3355, new_n3356, new_n3357,
    new_n3358, new_n3359, new_n3360, new_n3361, new_n3362_1, new_n3363,
    new_n3364, new_n3365, new_n3366, new_n3367, new_n3368, new_n3369,
    new_n3370, new_n3371, new_n3372, new_n3373, new_n3374, new_n3375,
    new_n3376, new_n3377, new_n3378, new_n3379, new_n3380, new_n3381,
    new_n3382, new_n3383, new_n3384, new_n3385, new_n3386, new_n3387,
    new_n3388, new_n3389, new_n3390, new_n3391, new_n3392, new_n3393,
    new_n3394, new_n3395, new_n3396, new_n3397, new_n3398, new_n3399,
    new_n3400, new_n3401, new_n3402, new_n3403, new_n3404, new_n3405,
    new_n3406, new_n3407, new_n3408, new_n3409_1, new_n3410, new_n3411,
    new_n3412, new_n3413, new_n3414, new_n3415, new_n3416, new_n3417,
    new_n3418, new_n3419, new_n3420, new_n3421, new_n3422, new_n3423,
    new_n3424, new_n3425, new_n3426, new_n3427, new_n3428, new_n3429,
    new_n3430, new_n3431, new_n3432, new_n3433, new_n3434, new_n3435,
    new_n3436, new_n3437, new_n3438, new_n3439, new_n3440, new_n3441,
    new_n3442, new_n3443, new_n3444, new_n3445, new_n3446, new_n3447,
    new_n3448, new_n3449, new_n3450, new_n3451, new_n3452, new_n3453,
    new_n3454, new_n3455, new_n3456, new_n3457, new_n3458, new_n3459,
    new_n3460, new_n3461, new_n3462, new_n3463, new_n3464, new_n3465,
    new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471,
    new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477,
    new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483,
    new_n3484, new_n3485, new_n3486, new_n3487, new_n3488, new_n3489,
    new_n3490, new_n3491, new_n3492, new_n3493, new_n3494, new_n3495,
    new_n3496, new_n3497, new_n3498, new_n3499, new_n3500, new_n3501,
    new_n3502, new_n3503, new_n3504, new_n3505, new_n3506, new_n3507,
    new_n3508, new_n3509, new_n3510, new_n3511, new_n3512, new_n3513,
    new_n3514, new_n3515, new_n3516, new_n3517, new_n3518, new_n3519,
    new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525,
    new_n3526, new_n3527, new_n3528, new_n3529, new_n3530, new_n3531,
    new_n3532, new_n3534, new_n3535, new_n3536, new_n3537, new_n3538,
    new_n3539, new_n3540, new_n3541, new_n3542, new_n3543, new_n3544,
    new_n3545, new_n3546, new_n3547, new_n3548, new_n3549, new_n3550,
    new_n3551, new_n3552, new_n3553, new_n3554, new_n3555, new_n3556,
    new_n3557, new_n3558, new_n3559, new_n3560, new_n3561, new_n3562,
    new_n3563, new_n3564, new_n3565, new_n3566, new_n3567, new_n3568,
    new_n3569, new_n3570, new_n3571, new_n3572, new_n3573, new_n3574,
    new_n3575, new_n3576, new_n3577, new_n3578, new_n3579, new_n3580,
    new_n3581, new_n3582, new_n3583, new_n3584, new_n3585, new_n3586,
    new_n3587, new_n3588, new_n3589, new_n3590, new_n3591_1, new_n3592,
    new_n3593, new_n3594, new_n3595, new_n3596, new_n3597, new_n3598,
    new_n3599, new_n3600, new_n3601, new_n3602, new_n3603, new_n3604,
    new_n3605, new_n3606, new_n3607, new_n3608, new_n3609, new_n3610,
    new_n3611, new_n3612, new_n3613, new_n3614, new_n3615, new_n3616,
    new_n3617, new_n3618, new_n3619, new_n3620, new_n3621, new_n3622,
    new_n3623, new_n3624, new_n3625, new_n3626, new_n3627, new_n3628,
    new_n3629, new_n3630, new_n3631, new_n3632, new_n3633, new_n3634,
    new_n3635, new_n3636, new_n3637, new_n3638, new_n3639, new_n3640,
    new_n3641_1, new_n3642, new_n3643, new_n3644, new_n3645, new_n3646,
    new_n3647, new_n3648, new_n3649, new_n3650, new_n3651, new_n3652,
    new_n3653, new_n3654, new_n3655, new_n3656, new_n3657, new_n3658,
    new_n3659, new_n3660, new_n3661, new_n3662, new_n3663, new_n3664,
    new_n3665, new_n3666, new_n3667, new_n3668, new_n3669_1, new_n3670,
    new_n3671, new_n3672, new_n3673, new_n3674, new_n3675, new_n3676,
    new_n3677_1, new_n3678, new_n3679, new_n3680, new_n3681, new_n3682,
    new_n3683, new_n3684, new_n3685, new_n3686, new_n3687, new_n3688,
    new_n3689, new_n3690, new_n3691, new_n3692, new_n3693, new_n3694,
    new_n3695, new_n3696, new_n3697, new_n3698, new_n3699, new_n3700,
    new_n3701, new_n3702, new_n3703, new_n3704, new_n3705, new_n3706,
    new_n3707, new_n3708, new_n3709, new_n3710, new_n3711, new_n3712,
    new_n3713, new_n3714, new_n3715, new_n3716, new_n3717, new_n3718,
    new_n3719, new_n3720, new_n3721, new_n3722, new_n3723, new_n3724,
    new_n3725, new_n3726, new_n3727, new_n3728, new_n3729, new_n3730,
    new_n3731, new_n3732, new_n3733, new_n3734, new_n3735, new_n3736,
    new_n3737, new_n3738, new_n3739, new_n3740, new_n3741, new_n3742,
    new_n3743, new_n3744, new_n3745, new_n3746, new_n3747, new_n3748_1,
    new_n3749, new_n3750, new_n3751, new_n3752, new_n3754, new_n3755,
    new_n3756, new_n3758, new_n3759, new_n3760, new_n3761, new_n3762,
    new_n3763, new_n3764, new_n3765, new_n3766, new_n3767, new_n3768,
    new_n3769_1, new_n3771, new_n3772, new_n3773, new_n3774, new_n3775,
    new_n3776, new_n3777, new_n3778, new_n3779, new_n3780, new_n3781,
    new_n3782, new_n3783, new_n3784, new_n3785, new_n3786, new_n3787,
    new_n3788, new_n3789, new_n3790_1, new_n3791, new_n3792, new_n3793,
    new_n3794, new_n3795, new_n3796, new_n3797, new_n3798, new_n3799,
    new_n3800, new_n3801, new_n3802, new_n3803, new_n3804, new_n3805,
    new_n3806, new_n3807, new_n3808, new_n3809, new_n3810, new_n3811,
    new_n3812, new_n3813, new_n3814, new_n3815_1, new_n3816, new_n3817,
    new_n3818, new_n3819, new_n3820, new_n3821, new_n3822, new_n3823,
    new_n3824, new_n3825, new_n3826, new_n3827, new_n3828, new_n3829,
    new_n3830, new_n3831, new_n3832_1, new_n3833, new_n3834, new_n3835,
    new_n3836, new_n3837, new_n3838, new_n3839, new_n3840, new_n3841,
    new_n3842, new_n3843, new_n3844, new_n3845, new_n3846, new_n3847,
    new_n3848, new_n3849, new_n3850, new_n3851, new_n3852, new_n3853,
    new_n3854, new_n3855, new_n3856, new_n3857, new_n3858, new_n3859,
    new_n3860, new_n3861, new_n3862, new_n3863, new_n3864, new_n3865,
    new_n3866, new_n3867, new_n3868, new_n3869, new_n3870, new_n3871,
    new_n3872, new_n3873, new_n3874, new_n3875, new_n3876, new_n3877,
    new_n3878, new_n3879, new_n3880, new_n3881, new_n3882, new_n3883,
    new_n3884, new_n3885, new_n3886, new_n3887, new_n3888, new_n3889,
    new_n3890, new_n3891, new_n3892, new_n3893, new_n3894, new_n3895,
    new_n3896, new_n3897, new_n3898, new_n3899, new_n3900, new_n3901,
    new_n3902, new_n3903, new_n3904, new_n3905, new_n3906, new_n3907,
    new_n3908, new_n3909, new_n3910, new_n3911, new_n3912, new_n3913,
    new_n3914, new_n3915, new_n3916, new_n3917, new_n3918, new_n3919,
    new_n3920, new_n3921, new_n3922, new_n3923, new_n3924, new_n3925,
    new_n3926, new_n3927, new_n3928, new_n3929, new_n3930, new_n3931,
    new_n3932, new_n3933, new_n3934, new_n3935, new_n3936, new_n3937,
    new_n3938, new_n3939, new_n3940, new_n3941, new_n3942, new_n3943,
    new_n3944, new_n3945, new_n3946_1, new_n3947, new_n3948, new_n3949,
    new_n3950, new_n3951, new_n3952, new_n3953, new_n3954, new_n3955,
    new_n3956, new_n3957, new_n3958, new_n3959, new_n3960, new_n3961,
    new_n3962, new_n3963, new_n3964, new_n3965, new_n3966, new_n3967,
    new_n3968, new_n3969, new_n3970, new_n3971, new_n3972, new_n3973,
    new_n3974, new_n3975, new_n3976, new_n3977, new_n3978, new_n3979,
    new_n3980, new_n3981, new_n3982, new_n3983, new_n3984, new_n3985,
    new_n3986, new_n3987, new_n3988, new_n3989, new_n3990, new_n3991,
    new_n3992, new_n3994, new_n3995, new_n3996, new_n3997, new_n3998,
    new_n3999, new_n4000, new_n4001, new_n4002, new_n4003, new_n4004,
    new_n4005, new_n4006_1, new_n4007, new_n4008, new_n4009, new_n4010,
    new_n4011, new_n4012, new_n4013, new_n4014, new_n4015, new_n4016,
    new_n4017, new_n4018, new_n4019, new_n4020, new_n4021, new_n4022,
    new_n4023, new_n4024, new_n4025, new_n4026, new_n4027, new_n4028,
    new_n4029, new_n4030, new_n4031, new_n4032, new_n4033, new_n4034,
    new_n4035, new_n4036, new_n4037, new_n4038, new_n4039, new_n4040,
    new_n4041, new_n4042, new_n4043, new_n4044, new_n4045, new_n4046,
    new_n4047, new_n4048, new_n4049, new_n4050, new_n4051, new_n4052,
    new_n4053, new_n4054, new_n4055, new_n4056, new_n4057, new_n4058,
    new_n4059_1, new_n4060, new_n4061, new_n4062, new_n4063, new_n4064,
    new_n4065, new_n4066, new_n4067, new_n4068, new_n4069, new_n4070,
    new_n4071, new_n4072, new_n4073, new_n4074, new_n4075_1, new_n4076,
    new_n4077, new_n4078, new_n4079, new_n4080, new_n4081, new_n4082,
    new_n4083, new_n4084, new_n4085, new_n4086, new_n4087, new_n4088,
    new_n4089, new_n4090, new_n4091, new_n4092, new_n4093, new_n4094,
    new_n4095, new_n4096, new_n4097, new_n4098, new_n4099, new_n4100,
    new_n4101, new_n4102, new_n4103, new_n4104, new_n4105, new_n4106,
    new_n4107, new_n4108, new_n4109, new_n4110, new_n4111, new_n4113,
    new_n4114_1, new_n4115, new_n4116, new_n4117, new_n4118, new_n4119,
    new_n4120, new_n4121, new_n4122_1, new_n4123, new_n4124, new_n4125,
    new_n4126, new_n4127, new_n4128, new_n4129, new_n4130, new_n4131,
    new_n4132, new_n4133, new_n4134, new_n4135, new_n4136, new_n4137,
    new_n4138, new_n4139, new_n4140, new_n4141_1, new_n4142, new_n4143,
    new_n4144, new_n4145, new_n4146, new_n4147, new_n4148, new_n4149,
    new_n4150, new_n4151, new_n4152, new_n4153, new_n4154, new_n4155,
    new_n4156, new_n4157, new_n4158, new_n4159, new_n4160, new_n4161,
    new_n4163, new_n4165, new_n4166, new_n4167, new_n4169, new_n4170,
    new_n4171, new_n4172, new_n4173, new_n4174, new_n4175, new_n4176,
    new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182,
    new_n4183, new_n4184, new_n4185, new_n4186, new_n4187, new_n4188,
    new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194,
    new_n4195, new_n4196, new_n4197, new_n4198, new_n4199, new_n4200,
    new_n4201, new_n4202_1, new_n4203, new_n4204, new_n4205, new_n4206,
    new_n4207, new_n4208, new_n4209, new_n4210, new_n4211, new_n4212,
    new_n4213, new_n4214, new_n4215, new_n4216, new_n4217, new_n4218,
    new_n4219, new_n4220, new_n4221, new_n4222, new_n4223, new_n4224,
    new_n4225, new_n4226, new_n4227, new_n4228, new_n4229, new_n4230,
    new_n4231, new_n4232, new_n4233, new_n4234, new_n4235, new_n4236,
    new_n4237, new_n4238, new_n4239, new_n4240, new_n4241, new_n4242,
    new_n4243, new_n4244, new_n4245, new_n4246, new_n4247, new_n4248,
    new_n4249, new_n4250, new_n4251, new_n4252, new_n4253, new_n4254,
    new_n4255, new_n4256, new_n4257, new_n4258, new_n4259, new_n4260,
    new_n4261, new_n4262, new_n4263, new_n4264, new_n4265, new_n4266,
    new_n4267, new_n4268, new_n4269, new_n4270, new_n4271, new_n4272,
    new_n4273, new_n4274, new_n4275, new_n4276, new_n4277, new_n4278,
    new_n4279, new_n4280, new_n4281, new_n4282, new_n4283, new_n4284,
    new_n4285, new_n4286, new_n4287, new_n4288, new_n4289, new_n4290,
    new_n4291, new_n4292, new_n4293, new_n4294, new_n4295, new_n4296,
    new_n4297, new_n4298, new_n4299, new_n4300, new_n4301, new_n4302,
    new_n4303, new_n4304, new_n4305, new_n4306, new_n4307, new_n4308,
    new_n4309, new_n4310, new_n4311, new_n4312, new_n4313, new_n4314,
    new_n4315, new_n4316, new_n4317, new_n4318, new_n4319, new_n4320,
    new_n4321, new_n4322, new_n4323, new_n4324, new_n4325, new_n4326,
    new_n4327, new_n4328, new_n4329, new_n4330_1, new_n4331, new_n4332,
    new_n4333, new_n4334, new_n4335_1, new_n4336, new_n4337, new_n4338,
    new_n4339, new_n4340, new_n4341, new_n4342, new_n4343, new_n4344,
    new_n4345, new_n4346, new_n4347, new_n4348, new_n4349, new_n4350,
    new_n4351, new_n4352, new_n4353, new_n4354, new_n4355, new_n4356,
    new_n4357_1, new_n4358, new_n4359, new_n4360, new_n4361, new_n4362,
    new_n4363, new_n4364, new_n4365, new_n4366, new_n4367, new_n4368,
    new_n4369, new_n4370, new_n4371, new_n4372, new_n4373, new_n4374,
    new_n4375, new_n4376, new_n4377, new_n4378, new_n4379, new_n4380,
    new_n4381, new_n4382_1, new_n4383, new_n4384, new_n4385, new_n4386,
    new_n4387, new_n4388, new_n4389, new_n4390, new_n4391, new_n4392,
    new_n4393, new_n4394, new_n4395, new_n4396, new_n4397, new_n4398,
    new_n4399, new_n4400, new_n4401, new_n4402, new_n4403, new_n4404,
    new_n4405, new_n4406, new_n4407, new_n4408, new_n4409, new_n4410,
    new_n4411, new_n4412, new_n4413, new_n4414, new_n4415, new_n4416,
    new_n4417, new_n4418, new_n4419_1, new_n4420, new_n4421, new_n4422,
    new_n4423, new_n4424, new_n4425, new_n4426, new_n4427, new_n4428,
    new_n4429, new_n4430, new_n4431, new_n4432, new_n4433, new_n4434,
    new_n4435, new_n4436, new_n4437, new_n4438, new_n4439, new_n4440,
    new_n4441, new_n4442, new_n4443, new_n4444, new_n4445, new_n4446,
    new_n4447, new_n4448, new_n4449, new_n4450, new_n4451, new_n4452_1,
    new_n4453, new_n4454, new_n4455, new_n4456, new_n4457, new_n4458,
    new_n4459, new_n4460, new_n4461, new_n4462, new_n4463, new_n4464,
    new_n4465, new_n4466, new_n4467, new_n4468, new_n4469, new_n4470_1,
    new_n4471, new_n4472, new_n4473, new_n4474, new_n4475, new_n4476,
    new_n4477, new_n4478, new_n4479, new_n4480, new_n4481, new_n4482,
    new_n4483, new_n4484, new_n4485, new_n4486, new_n4487, new_n4488,
    new_n4489, new_n4490, new_n4491, new_n4492, new_n4493, new_n4494,
    new_n4495, new_n4496, new_n4497, new_n4498, new_n4499, new_n4500,
    new_n4501, new_n4502, new_n4503, new_n4504, new_n4505, new_n4506,
    new_n4507, new_n4508, new_n4509, new_n4510, new_n4511, new_n4512,
    new_n4513, new_n4514, new_n4515, new_n4516, new_n4517, new_n4518,
    new_n4519, new_n4520, new_n4521, new_n4522, new_n4523, new_n4524,
    new_n4525, new_n4526, new_n4527, new_n4528, new_n4529, new_n4530,
    new_n4531, new_n4532, new_n4533, new_n4534, new_n4535, new_n4536,
    new_n4537, new_n4538, new_n4539, new_n4540, new_n4541, new_n4542,
    new_n4543, new_n4544, new_n4545, new_n4546, new_n4547, new_n4548,
    new_n4549, new_n4550, new_n4551, new_n4552, new_n4553_1, new_n4554,
    new_n4555, new_n4556, new_n4557, new_n4558, new_n4559, new_n4560,
    new_n4561, new_n4562, new_n4563, new_n4564, new_n4565, new_n4566,
    new_n4567, new_n4568, new_n4569, new_n4570, new_n4571, new_n4572,
    new_n4573, new_n4574, new_n4575, new_n4576, new_n4577, new_n4578,
    new_n4579, new_n4580, new_n4581, new_n4582, new_n4583, new_n4584,
    new_n4585, new_n4586, new_n4587, new_n4588, new_n4589, new_n4590,
    new_n4591, new_n4592, new_n4593, new_n4594, new_n4595, new_n4596,
    new_n4597, new_n4598, new_n4599, new_n4600, new_n4601, new_n4602,
    new_n4603, new_n4604, new_n4605, new_n4606, new_n4607, new_n4608,
    new_n4609, new_n4610, new_n4611, new_n4612, new_n4613, new_n4614,
    new_n4615, new_n4616, new_n4617, new_n4618, new_n4619, new_n4620,
    new_n4621, new_n4622, new_n4623, new_n4624, new_n4625, new_n4626,
    new_n4627, new_n4628, new_n4629, new_n4630, new_n4631, new_n4632,
    new_n4633, new_n4634, new_n4635, new_n4636, new_n4637, new_n4638,
    new_n4639, new_n4640, new_n4641, new_n4642, new_n4643, new_n4644,
    new_n4645, new_n4646, new_n4647, new_n4648, new_n4649, new_n4650,
    new_n4651, new_n4652, new_n4653, new_n4654, new_n4655, new_n4656,
    new_n4657, new_n4658, new_n4659, new_n4660, new_n4661, new_n4662,
    new_n4663, new_n4664, new_n4665, new_n4666, new_n4667, new_n4668,
    new_n4669, new_n4670, new_n4671, new_n4672, new_n4673, new_n4674,
    new_n4675, new_n4676, new_n4677, new_n4678, new_n4679, new_n4680,
    new_n4681, new_n4682, new_n4683, new_n4684, new_n4685, new_n4686,
    new_n4687, new_n4688, new_n4689, new_n4690, new_n4691, new_n4692,
    new_n4693, new_n4694, new_n4695, new_n4696, new_n4697, new_n4698,
    new_n4699, new_n4700, new_n4701, new_n4702, new_n4703, new_n4704,
    new_n4705, new_n4706, new_n4707, new_n4708, new_n4709, new_n4710,
    new_n4711, new_n4712, new_n4713, new_n4714, new_n4715, new_n4716,
    new_n4717, new_n4718, new_n4719, new_n4720, new_n4721, new_n4722,
    new_n4723, new_n4724, new_n4725, new_n4726, new_n4727, new_n4728,
    new_n4729, new_n4730, new_n4731, new_n4732, new_n4733, new_n4734,
    new_n4735, new_n4736, new_n4737, new_n4738, new_n4739, new_n4740,
    new_n4741, new_n4742, new_n4743_1, new_n4744, new_n4745, new_n4746,
    new_n4747, new_n4748_1, new_n4749, new_n4750, new_n4751, new_n4752,
    new_n4753, new_n4754, new_n4755, new_n4756, new_n4757, new_n4758,
    new_n4759, new_n4760, new_n4761, new_n4762, new_n4763, new_n4764,
    new_n4765, new_n4766, new_n4767, new_n4768, new_n4769, new_n4770,
    new_n4771, new_n4772, new_n4773, new_n4774, new_n4775, new_n4776,
    new_n4777_1, new_n4778, new_n4779, new_n4780, new_n4781, new_n4782,
    new_n4783, new_n4784, new_n4785, new_n4786, new_n4787, new_n4788,
    new_n4789, new_n4790, new_n4791, new_n4792, new_n4793, new_n4794,
    new_n4795, new_n4796, new_n4797, new_n4798, new_n4799, new_n4800,
    new_n4801, new_n4802, new_n4803, new_n4804, new_n4805, new_n4806,
    new_n4807, new_n4808, new_n4809, new_n4810, new_n4811, new_n4812,
    new_n4813, new_n4814, new_n4815, new_n4816, new_n4817, new_n4818,
    new_n4819, new_n4820, new_n4821, new_n4822, new_n4823, new_n4824_1,
    new_n4825, new_n4826, new_n4827, new_n4828, new_n4829, new_n4830,
    new_n4831, new_n4832, new_n4833, new_n4834, new_n4835, new_n4836,
    new_n4837, new_n4838, new_n4839, new_n4840, new_n4841, new_n4842,
    new_n4843, new_n4844, new_n4845, new_n4846, new_n4847, new_n4848,
    new_n4849, new_n4850, new_n4851, new_n4852, new_n4853, new_n4854,
    new_n4855, new_n4856, new_n4857, new_n4858, new_n4859, new_n4860,
    new_n4861, new_n4862_1, new_n4863, new_n4864_1, new_n4865, new_n4866,
    new_n4867, new_n4868, new_n4869, new_n4870, new_n4871, new_n4872,
    new_n4873, new_n4874, new_n4875, new_n4876, new_n4877, new_n4878,
    new_n4879, new_n4880, new_n4881, new_n4882, new_n4883, new_n4884,
    new_n4885, new_n4886, new_n4887, new_n4888, new_n4889, new_n4890,
    new_n4891, new_n4892, new_n4893, new_n4894, new_n4895, new_n4896,
    new_n4897, new_n4898, new_n4899, new_n4900, new_n4901, new_n4902,
    new_n4903, new_n4904, new_n4905, new_n4906, new_n4907, new_n4908,
    new_n4909, new_n4910, new_n4911, new_n4912, new_n4913, new_n4914,
    new_n4915, new_n4916, new_n4917, new_n4918, new_n4919, new_n4920,
    new_n4921, new_n4922, new_n4923, new_n4924, new_n4925, new_n4926,
    new_n4927, new_n4928, new_n4929, new_n4930, new_n4931, new_n4932,
    new_n4933, new_n4934, new_n4935, new_n4936, new_n4937, new_n4938,
    new_n4939, new_n4940, new_n4941, new_n4942, new_n4943, new_n4944,
    new_n4945, new_n4946, new_n4947, new_n4948, new_n4949, new_n4950,
    new_n4951, new_n4952, new_n4953, new_n4954, new_n4955, new_n4956,
    new_n4957, new_n4958, new_n4959, new_n4960, new_n4961, new_n4962,
    new_n4963, new_n4964_1, new_n4965, new_n4966, new_n4967, new_n4968,
    new_n4969, new_n4970, new_n4971, new_n4972, new_n4973, new_n4974,
    new_n4975, new_n4976, new_n4977, new_n4978, new_n4979, new_n4980,
    new_n4981, new_n4982, new_n4983, new_n4984, new_n4985, new_n4986,
    new_n4987, new_n4988, new_n4989, new_n4990, new_n4991, new_n4992,
    new_n4993, new_n4994, new_n4995, new_n4996, new_n4997, new_n4998_1,
    new_n4999, new_n5000, new_n5001, new_n5002, new_n5003_1, new_n5004,
    new_n5005, new_n5006, new_n5007, new_n5008, new_n5009, new_n5010,
    new_n5011, new_n5012, new_n5013, new_n5014, new_n5015, new_n5016,
    new_n5017, new_n5018, new_n5019, new_n5020, new_n5021, new_n5022,
    new_n5023, new_n5024, new_n5025, new_n5026, new_n5027, new_n5028,
    new_n5029, new_n5030, new_n5031_1, new_n5032, new_n5033, new_n5034,
    new_n5035, new_n5036, new_n5037, new_n5038, new_n5039, new_n5040,
    new_n5041, new_n5042, new_n5043, new_n5044, new_n5045, new_n5046,
    new_n5047, new_n5048, new_n5049, new_n5050, new_n5051, new_n5052,
    new_n5053, new_n5054, new_n5055, new_n5056, new_n5057, new_n5058,
    new_n5059, new_n5060_1, new_n5061, new_n5062, new_n5063, new_n5064,
    new_n5065_1, new_n5066, new_n5067, new_n5068, new_n5069, new_n5070,
    new_n5071, new_n5072, new_n5073, new_n5074, new_n5075, new_n5076,
    new_n5077, new_n5078, new_n5079, new_n5080, new_n5081, new_n5082,
    new_n5083, new_n5084, new_n5085, new_n5086, new_n5087, new_n5088,
    new_n5089, new_n5090, new_n5091, new_n5092, new_n5093, new_n5094,
    new_n5095, new_n5096, new_n5097, new_n5098, new_n5099, new_n5100,
    new_n5101, new_n5102, new_n5103, new_n5104, new_n5105, new_n5106,
    new_n5107, new_n5108, new_n5109, new_n5110, new_n5111, new_n5112,
    new_n5113, new_n5114, new_n5115, new_n5116, new_n5117, new_n5118,
    new_n5119, new_n5120, new_n5121, new_n5122, new_n5123, new_n5124,
    new_n5125, new_n5126, new_n5127, new_n5128, new_n5129, new_n5130,
    new_n5131, new_n5132, new_n5133, new_n5134, new_n5135, new_n5136,
    new_n5137, new_n5138, new_n5139, new_n5140, new_n5141, new_n5142,
    new_n5143, new_n5144, new_n5145, new_n5146, new_n5147, new_n5148,
    new_n5149, new_n5150, new_n5151, new_n5152, new_n5153, new_n5154,
    new_n5155, new_n5156, new_n5157, new_n5158, new_n5159, new_n5160,
    new_n5161, new_n5162, new_n5163, new_n5164, new_n5165, new_n5166,
    new_n5167_1, new_n5168, new_n5170, new_n5171, new_n5172, new_n5173,
    new_n5174, new_n5175, new_n5176, new_n5177, new_n5178, new_n5179,
    new_n5180, new_n5182, new_n5183, new_n5184, new_n5185, new_n5186,
    new_n5187, new_n5188, new_n5189_1, new_n5190, new_n5191, new_n5192,
    new_n5193, new_n5194, new_n5195, new_n5196, new_n5197, new_n5198,
    new_n5199, new_n5200, new_n5201, new_n5202, new_n5203, new_n5204,
    new_n5205, new_n5206, new_n5207, new_n5208, new_n5209, new_n5210,
    new_n5211, new_n5212, new_n5213, new_n5214_1, new_n5215, new_n5216,
    new_n5217, new_n5218, new_n5219, new_n5220, new_n5221, new_n5222,
    new_n5223, new_n5224, new_n5225, new_n5226, new_n5227, new_n5228,
    new_n5229, new_n5230, new_n5231, new_n5232, new_n5233, new_n5234,
    new_n5235, new_n5236, new_n5237, new_n5238, new_n5239, new_n5240,
    new_n5241, new_n5242, new_n5243, new_n5244, new_n5245, new_n5246,
    new_n5247, new_n5248, new_n5249, new_n5250, new_n5251, new_n5252,
    new_n5253, new_n5254, new_n5255, new_n5256, new_n5257, new_n5258,
    new_n5259, new_n5260, new_n5261, new_n5262, new_n5263, new_n5264,
    new_n5265, new_n5266, new_n5267, new_n5268, new_n5269, new_n5270,
    new_n5271, new_n5272, new_n5273, new_n5274, new_n5275, new_n5276,
    new_n5277, new_n5278, new_n5279, new_n5280, new_n5281, new_n5282,
    new_n5283, new_n5284, new_n5285, new_n5286, new_n5287, new_n5288,
    new_n5289, new_n5290, new_n5291, new_n5292, new_n5293, new_n5294,
    new_n5295, new_n5296, new_n5297, new_n5298, new_n5299, new_n5300,
    new_n5301, new_n5302, new_n5303, new_n5304, new_n5305, new_n5306,
    new_n5307, new_n5308, new_n5309, new_n5310, new_n5311, new_n5312,
    new_n5313, new_n5314, new_n5315, new_n5316, new_n5317, new_n5318,
    new_n5319, new_n5320_1, new_n5321, new_n5322, new_n5323, new_n5324,
    new_n5325, new_n5326, new_n5327, new_n5328, new_n5329, new_n5330,
    new_n5331, new_n5332, new_n5333, new_n5334, new_n5335, new_n5336,
    new_n5337, new_n5338, new_n5339, new_n5340, new_n5341, new_n5342,
    new_n5343, new_n5344, new_n5345, new_n5346, new_n5347, new_n5348,
    new_n5349, new_n5350, new_n5351, new_n5352, new_n5353, new_n5354,
    new_n5355, new_n5356_1, new_n5357, new_n5358, new_n5359, new_n5360,
    new_n5361, new_n5362, new_n5363, new_n5364_1, new_n5365, new_n5366,
    new_n5367, new_n5368, new_n5369, new_n5370, new_n5371, new_n5372,
    new_n5373, new_n5374, new_n5375, new_n5376, new_n5377, new_n5378,
    new_n5379, new_n5380, new_n5381, new_n5382, new_n5383, new_n5384,
    new_n5385, new_n5386, new_n5387, new_n5388, new_n5389, new_n5390,
    new_n5391, new_n5392, new_n5393, new_n5394, new_n5395, new_n5396,
    new_n5397, new_n5398, new_n5399, new_n5400, new_n5401, new_n5403,
    new_n5404, new_n5405, new_n5406, new_n5407, new_n5408, new_n5409,
    new_n5410, new_n5411, new_n5412, new_n5413, new_n5414, new_n5415,
    new_n5416, new_n5417, new_n5418, new_n5419, new_n5420, new_n5421,
    new_n5422, new_n5423, new_n5424, new_n5425, new_n5426, new_n5427_1,
    new_n5428, new_n5429, new_n5430, new_n5431, new_n5432, new_n5433,
    new_n5434, new_n5435, new_n5436, new_n5437, new_n5438, new_n5439,
    new_n5440, new_n5441, new_n5442, new_n5443, new_n5444, new_n5445,
    new_n5446, new_n5447, new_n5448, new_n5449, new_n5450, new_n5451,
    new_n5452, new_n5453, new_n5454, new_n5455, new_n5456, new_n5457,
    new_n5458, new_n5459, new_n5460, new_n5461, new_n5462, new_n5463,
    new_n5464, new_n5465, new_n5466, new_n5467, new_n5468, new_n5469,
    new_n5470_1, new_n5471, new_n5472, new_n5473, new_n5474, new_n5475,
    new_n5476, new_n5477, new_n5478, new_n5479, new_n5480, new_n5481,
    new_n5482, new_n5483, new_n5484, new_n5485, new_n5486, new_n5487,
    new_n5488, new_n5489, new_n5490, new_n5491, new_n5492, new_n5493,
    new_n5494, new_n5495, new_n5496, new_n5497, new_n5498, new_n5499,
    new_n5500, new_n5501, new_n5502, new_n5503, new_n5504, new_n5505,
    new_n5506, new_n5507, new_n5508, new_n5509, new_n5510, new_n5511,
    new_n5512, new_n5513, new_n5514, new_n5515, new_n5516, new_n5517,
    new_n5518, new_n5519, new_n5520, new_n5521, new_n5522, new_n5523,
    new_n5524, new_n5525, new_n5526, new_n5527, new_n5528, new_n5529,
    new_n5530, new_n5531, new_n5532, new_n5533, new_n5534, new_n5535,
    new_n5536_1, new_n5537, new_n5538, new_n5539, new_n5540, new_n5541,
    new_n5542, new_n5543, new_n5544, new_n5545, new_n5546, new_n5547,
    new_n5548_1, new_n5549_1, new_n5550, new_n5551, new_n5552, new_n5553,
    new_n5554, new_n5555, new_n5556, new_n5557_1, new_n5558, new_n5559,
    new_n5560, new_n5561, new_n5562, new_n5563, new_n5564, new_n5565,
    new_n5566, new_n5567, new_n5568_1, new_n5569, new_n5570, new_n5571,
    new_n5572, new_n5573, new_n5574, new_n5575, new_n5576, new_n5577,
    new_n5578, new_n5579, new_n5580, new_n5581, new_n5582, new_n5583,
    new_n5584, new_n5585, new_n5586_1, new_n5587, new_n5588, new_n5589,
    new_n5590, new_n5591, new_n5592, new_n5593, new_n5594, new_n5595,
    new_n5596, new_n5597, new_n5598, new_n5599, new_n5600, new_n5601,
    new_n5602, new_n5603, new_n5604, new_n5605, new_n5606, new_n5607,
    new_n5608, new_n5609_1, new_n5610, new_n5611, new_n5612, new_n5613,
    new_n5614, new_n5615, new_n5616, new_n5617, new_n5618, new_n5619,
    new_n5620, new_n5621, new_n5622, new_n5623, new_n5624, new_n5625,
    new_n5626, new_n5627, new_n5628, new_n5629, new_n5630, new_n5631,
    new_n5632, new_n5633, new_n5634, new_n5635, new_n5636, new_n5637,
    new_n5638, new_n5639, new_n5640, new_n5641, new_n5642, new_n5643,
    new_n5644, new_n5645, new_n5646, new_n5647, new_n5648, new_n5650,
    new_n5651, new_n5652, new_n5653, new_n5654, new_n5655, new_n5656,
    new_n5657, new_n5658, new_n5659, new_n5660, new_n5662, new_n5663,
    new_n5664, new_n5665, new_n5666, new_n5667, new_n5668, new_n5669,
    new_n5670, new_n5671_1, new_n5672, new_n5673, new_n5674, new_n5675,
    new_n5676, new_n5677, new_n5678, new_n5679, new_n5680, new_n5681,
    new_n5682, new_n5683, new_n5684_1, new_n5685, new_n5686, new_n5687,
    new_n5688, new_n5689, new_n5690, new_n5691, new_n5692, new_n5693,
    new_n5694, new_n5695, new_n5696, new_n5697, new_n5698, new_n5699,
    new_n5700, new_n5701, new_n5702, new_n5703, new_n5704, new_n5705,
    new_n5706, new_n5707, new_n5708, new_n5709, new_n5710, new_n5711,
    new_n5712, new_n5713, new_n5714, new_n5715_1, new_n5716, new_n5717,
    new_n5718, new_n5719, new_n5720, new_n5721, new_n5722, new_n5723,
    new_n5724, new_n5725, new_n5726, new_n5727, new_n5728, new_n5729_1,
    new_n5730, new_n5731, new_n5732, new_n5733, new_n5734, new_n5735,
    new_n5736, new_n5737, new_n5738, new_n5739, new_n5740, new_n5741,
    new_n5742, new_n5743, new_n5744, new_n5745, new_n5746, new_n5747,
    new_n5748, new_n5749, new_n5750, new_n5751, new_n5752, new_n5753,
    new_n5754, new_n5755, new_n5756, new_n5757, new_n5758_1, new_n5759,
    new_n5760, new_n5761, new_n5762, new_n5763, new_n5764, new_n5765,
    new_n5766, new_n5767, new_n5768, new_n5769, new_n5770, new_n5771,
    new_n5772, new_n5773, new_n5774, new_n5775, new_n5776, new_n5777,
    new_n5778, new_n5779, new_n5780, new_n5781, new_n5782, new_n5783,
    new_n5784, new_n5785, new_n5786, new_n5787, new_n5788, new_n5789,
    new_n5790, new_n5791, new_n5792, new_n5793, new_n5794, new_n5795,
    new_n5796, new_n5797, new_n5798, new_n5799, new_n5800, new_n5801_1,
    new_n5802, new_n5803, new_n5804, new_n5805, new_n5806, new_n5807,
    new_n5808, new_n5809, new_n5810, new_n5811, new_n5812, new_n5813,
    new_n5814, new_n5815, new_n5816, new_n5817, new_n5818, new_n5819,
    new_n5820, new_n5821, new_n5822, new_n5823, new_n5824, new_n5825,
    new_n5826, new_n5827, new_n5828, new_n5829, new_n5830, new_n5831,
    new_n5832, new_n5833, new_n5834, new_n5835, new_n5836, new_n5837,
    new_n5838, new_n5839, new_n5840, new_n5841, new_n5842, new_n5843,
    new_n5844, new_n5845, new_n5846, new_n5847, new_n5848, new_n5849,
    new_n5850, new_n5851, new_n5852, new_n5853, new_n5854, new_n5855,
    new_n5856, new_n5857, new_n5858, new_n5859, new_n5860, new_n5861,
    new_n5862, new_n5863, new_n5864, new_n5865, new_n5866, new_n5867,
    new_n5868, new_n5869, new_n5870, new_n5871, new_n5872, new_n5873,
    new_n5874, new_n5875, new_n5876, new_n5877, new_n5878, new_n5879,
    new_n5880, new_n5881, new_n5882_1, new_n5883, new_n5884_1, new_n5885,
    new_n5886, new_n5887, new_n5888, new_n5889, new_n5890, new_n5891,
    new_n5892, new_n5893, new_n5894, new_n5895, new_n5896, new_n5897,
    new_n5898, new_n5899, new_n5900, new_n5901, new_n5902, new_n5903,
    new_n5904, new_n5905, new_n5906, new_n5907, new_n5908, new_n5909,
    new_n5910, new_n5911, new_n5912, new_n5913, new_n5914, new_n5915,
    new_n5916, new_n5917, new_n5918, new_n5919, new_n5920_1, new_n5921,
    new_n5922, new_n5923, new_n5924, new_n5925, new_n5926, new_n5927,
    new_n5928, new_n5929, new_n5930, new_n5931, new_n5932, new_n5933,
    new_n5934, new_n5935, new_n5936, new_n5937, new_n5938, new_n5939,
    new_n5940, new_n5941, new_n5942, new_n5943, new_n5944, new_n5945,
    new_n5946, new_n5947, new_n5948, new_n5949, new_n5950, new_n5951,
    new_n5952, new_n5953, new_n5954, new_n5955, new_n5956, new_n5957,
    new_n5958, new_n5959, new_n5960, new_n5961, new_n5962_1, new_n5963,
    new_n5964, new_n5965, new_n5966, new_n5967, new_n5968, new_n5969_1,
    new_n5970, new_n5971, new_n5972, new_n5973, new_n5974, new_n5975,
    new_n5976, new_n5977, new_n5978, new_n5979, new_n5980, new_n5981,
    new_n5982, new_n5983, new_n5984, new_n5985, new_n5986, new_n5987,
    new_n5988, new_n5989, new_n5990, new_n5991, new_n5992, new_n5993,
    new_n5994, new_n5995, new_n5996, new_n5997, new_n5998, new_n5999,
    new_n6000, new_n6001, new_n6002, new_n6003, new_n6004, new_n6005,
    new_n6006, new_n6007, new_n6008, new_n6009, new_n6010, new_n6011,
    new_n6012, new_n6013, new_n6014, new_n6015, new_n6016, new_n6017,
    new_n6018, new_n6019_1, new_n6020, new_n6021, new_n6022, new_n6023_1,
    new_n6024, new_n6025, new_n6026, new_n6027, new_n6028, new_n6029,
    new_n6030, new_n6031, new_n6032, new_n6033, new_n6034, new_n6035,
    new_n6036, new_n6037, new_n6038, new_n6039, new_n6040, new_n6041,
    new_n6042, new_n6043, new_n6044, new_n6045, new_n6046, new_n6047,
    new_n6048, new_n6049, new_n6050, new_n6051, new_n6052, new_n6053,
    new_n6054, new_n6055, new_n6056, new_n6057, new_n6058, new_n6059,
    new_n6060, new_n6061, new_n6062, new_n6063, new_n6064, new_n6065,
    new_n6066, new_n6067, new_n6068, new_n6069, new_n6070, new_n6071,
    new_n6072, new_n6073, new_n6074, new_n6075, new_n6076, new_n6077,
    new_n6078, new_n6079, new_n6080, new_n6081, new_n6082, new_n6083,
    new_n6084, new_n6085_1, new_n6086, new_n6087, new_n6088, new_n6089,
    new_n6090, new_n6091, new_n6092, new_n6093, new_n6094, new_n6095,
    new_n6096, new_n6097, new_n6098, new_n6099, new_n6100, new_n6101,
    new_n6102, new_n6103_1, new_n6104, new_n6105, new_n6106, new_n6107,
    new_n6108, new_n6109_1, new_n6110, new_n6111, new_n6112, new_n6113,
    new_n6114, new_n6115, new_n6116, new_n6117, new_n6118, new_n6119,
    new_n6120, new_n6121, new_n6122, new_n6123, new_n6124, new_n6125,
    new_n6126, new_n6127, new_n6128, new_n6129, new_n6130, new_n6131,
    new_n6132, new_n6133, new_n6134, new_n6135, new_n6136, new_n6137,
    new_n6138, new_n6139, new_n6140, new_n6141, new_n6142, new_n6143,
    new_n6144, new_n6145, new_n6146, new_n6147, new_n6148, new_n6149_1,
    new_n6150, new_n6151, new_n6152, new_n6153, new_n6154, new_n6155,
    new_n6156, new_n6157, new_n6158, new_n6159, new_n6160, new_n6161,
    new_n6162, new_n6163, new_n6164, new_n6165, new_n6166, new_n6167,
    new_n6168_1, new_n6169, new_n6170, new_n6171, new_n6172, new_n6173,
    new_n6174, new_n6175, new_n6176, new_n6177, new_n6178, new_n6179,
    new_n6180, new_n6181, new_n6182, new_n6183, new_n6184, new_n6185,
    new_n6186, new_n6187, new_n6188, new_n6189, new_n6190, new_n6191,
    new_n6192, new_n6193, new_n6194, new_n6195, new_n6196, new_n6197,
    new_n6198, new_n6199, new_n6201, new_n6202, new_n6203, new_n6204,
    new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210,
    new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216,
    new_n6217, new_n6218, new_n6219, new_n6220, new_n6221, new_n6222,
    new_n6223, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246,
    new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254, new_n6255, new_n6256, new_n6257, new_n6258,
    new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264,
    new_n6265, new_n6266, new_n6267, new_n6268, new_n6269, new_n6270,
    new_n6271, new_n6272, new_n6273, new_n6274, new_n6275, new_n6276,
    new_n6277, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282,
    new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294,
    new_n6295, new_n6296, new_n6297_1, new_n6298, new_n6299, new_n6300,
    new_n6301_1, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333_1, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358, new_n6359, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6376, new_n6377, new_n6378,
    new_n6379, new_n6380, new_n6381, new_n6382, new_n6383, new_n6384,
    new_n6385, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390,
    new_n6391, new_n6392_1, new_n6393, new_n6394, new_n6395, new_n6396,
    new_n6397, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402,
    new_n6403, new_n6404, new_n6405, new_n6406, new_n6407, new_n6408,
    new_n6409_1, new_n6410, new_n6411, new_n6412, new_n6413, new_n6414,
    new_n6415, new_n6416, new_n6417, new_n6418, new_n6419, new_n6420,
    new_n6421, new_n6422, new_n6423, new_n6424, new_n6425, new_n6426,
    new_n6427, new_n6428, new_n6429, new_n6430, new_n6431, new_n6432,
    new_n6433, new_n6434_1, new_n6435, new_n6436, new_n6437, new_n6438,
    new_n6439, new_n6440, new_n6441, new_n6442, new_n6443, new_n6444,
    new_n6445, new_n6446, new_n6447, new_n6448, new_n6449, new_n6450,
    new_n6451, new_n6452, new_n6453, new_n6454, new_n6455, new_n6456,
    new_n6457, new_n6458, new_n6459, new_n6460, new_n6461, new_n6462,
    new_n6463, new_n6464, new_n6465, new_n6466, new_n6467, new_n6468,
    new_n6469, new_n6470, new_n6471, new_n6472, new_n6473, new_n6474,
    new_n6475, new_n6476, new_n6477, new_n6478, new_n6479, new_n6480,
    new_n6481, new_n6482, new_n6483, new_n6484, new_n6485, new_n6486,
    new_n6487, new_n6488, new_n6489, new_n6490, new_n6491, new_n6492,
    new_n6493, new_n6494, new_n6495, new_n6496, new_n6497, new_n6498,
    new_n6499, new_n6500, new_n6501, new_n6502, new_n6503, new_n6504,
    new_n6505, new_n6506, new_n6507, new_n6508, new_n6509, new_n6510,
    new_n6511, new_n6512, new_n6513, new_n6514, new_n6515, new_n6516,
    new_n6517, new_n6518, new_n6519, new_n6520, new_n6521, new_n6522,
    new_n6523, new_n6524, new_n6525, new_n6526, new_n6527, new_n6528,
    new_n6529, new_n6530, new_n6531, new_n6532, new_n6533, new_n6534,
    new_n6535, new_n6536, new_n6537, new_n6538, new_n6539, new_n6540,
    new_n6541, new_n6542, new_n6543, new_n6544, new_n6545, new_n6546,
    new_n6547, new_n6548, new_n6549, new_n6550, new_n6551, new_n6552,
    new_n6553, new_n6554, new_n6555, new_n6556, new_n6557, new_n6558,
    new_n6559, new_n6560, new_n6561, new_n6562, new_n6563, new_n6564,
    new_n6565, new_n6566, new_n6567, new_n6568, new_n6569, new_n6570,
    new_n6571, new_n6572, new_n6573, new_n6574, new_n6575, new_n6576,
    new_n6577, new_n6578, new_n6579, new_n6580, new_n6581, new_n6582,
    new_n6583, new_n6584, new_n6585, new_n6586_1, new_n6587, new_n6588,
    new_n6589, new_n6590, new_n6591, new_n6592, new_n6593, new_n6594,
    new_n6595, new_n6596, new_n6597, new_n6598, new_n6599, new_n6600,
    new_n6601, new_n6602, new_n6603, new_n6604, new_n6605, new_n6606,
    new_n6607, new_n6608, new_n6609, new_n6610, new_n6611, new_n6612,
    new_n6613, new_n6614, new_n6615, new_n6616, new_n6617, new_n6618,
    new_n6619, new_n6620, new_n6621, new_n6622, new_n6623, new_n6624,
    new_n6625, new_n6626, new_n6627, new_n6628, new_n6629, new_n6630,
    new_n6631, new_n6632, new_n6633, new_n6634, new_n6635, new_n6636,
    new_n6637, new_n6638, new_n6639, new_n6640, new_n6641, new_n6642,
    new_n6643, new_n6644, new_n6645, new_n6646, new_n6647, new_n6648,
    new_n6649, new_n6650, new_n6651, new_n6652, new_n6653, new_n6654,
    new_n6655_1, new_n6656, new_n6657, new_n6658, new_n6659, new_n6661,
    new_n6662, new_n6663, new_n6664, new_n6665, new_n6666, new_n6667,
    new_n6668_1, new_n6669, new_n6670, new_n6671, new_n6672, new_n6673,
    new_n6674, new_n6675, new_n6676, new_n6677, new_n6678, new_n6679,
    new_n6680, new_n6681, new_n6682, new_n6683_1, new_n6684, new_n6685,
    new_n6686, new_n6687, new_n6688, new_n6689, new_n6690, new_n6691,
    new_n6692, new_n6693, new_n6694, new_n6695, new_n6696, new_n6697,
    new_n6698, new_n6699, new_n6700, new_n6701, new_n6702, new_n6703,
    new_n6704, new_n6705, new_n6706, new_n6707, new_n6708, new_n6709,
    new_n6710, new_n6711, new_n6712, new_n6713, new_n6714, new_n6715,
    new_n6716, new_n6717, new_n6718, new_n6719, new_n6720, new_n6721,
    new_n6722, new_n6723, new_n6724, new_n6725, new_n6726, new_n6727,
    new_n6728, new_n6729, new_n6730, new_n6731, new_n6732, new_n6733,
    new_n6734, new_n6735, new_n6736, new_n6737, new_n6738, new_n6739,
    new_n6740, new_n6741, new_n6742, new_n6743, new_n6744, new_n6745,
    new_n6746, new_n6747, new_n6748, new_n6749, new_n6750, new_n6751,
    new_n6752, new_n6753, new_n6754, new_n6755, new_n6756, new_n6757,
    new_n6758, new_n6759, new_n6760, new_n6761, new_n6762, new_n6763,
    new_n6764, new_n6765, new_n6766, new_n6767, new_n6768, new_n6769,
    new_n6770, new_n6771, new_n6772, new_n6773, new_n6774, new_n6775,
    new_n6776, new_n6777, new_n6778, new_n6779, new_n6780, new_n6781,
    new_n6782, new_n6783, new_n6784, new_n6785, new_n6786, new_n6787,
    new_n6788, new_n6789, new_n6790, new_n6791, new_n6792, new_n6793,
    new_n6794, new_n6795, new_n6796, new_n6797, new_n6798, new_n6799,
    new_n6800, new_n6801, new_n6802, new_n6803, new_n6804, new_n6805,
    new_n6806, new_n6807, new_n6808, new_n6809, new_n6810, new_n6811,
    new_n6812, new_n6813, new_n6814, new_n6815, new_n6816, new_n6817,
    new_n6818_1, new_n6819, new_n6820, new_n6821, new_n6822, new_n6823,
    new_n6824, new_n6825, new_n6826_1, new_n6827, new_n6828, new_n6829,
    new_n6830, new_n6831, new_n6832, new_n6833, new_n6834, new_n6835,
    new_n6836, new_n6837, new_n6838, new_n6839, new_n6840, new_n6841,
    new_n6842, new_n6843_1, new_n6844, new_n6845, new_n6846, new_n6847,
    new_n6848, new_n6849, new_n6850, new_n6851, new_n6852, new_n6853,
    new_n6854, new_n6855, new_n6856, new_n6857, new_n6858, new_n6859,
    new_n6860, new_n6861, new_n6862_1, new_n6863, new_n6864, new_n6865,
    new_n6866, new_n6867, new_n6868, new_n6869, new_n6870, new_n6871,
    new_n6872, new_n6873, new_n6874, new_n6875, new_n6876, new_n6877,
    new_n6878, new_n6879, new_n6880, new_n6881, new_n6882, new_n6883,
    new_n6884, new_n6885, new_n6886, new_n6887, new_n6888, new_n6889,
    new_n6890, new_n6891, new_n6892, new_n6893, new_n6894, new_n6895,
    new_n6896, new_n6897, new_n6898, new_n6899, new_n6900, new_n6901,
    new_n6902, new_n6903, new_n6904, new_n6905, new_n6906, new_n6907,
    new_n6908, new_n6909, new_n6910, new_n6911, new_n6912, new_n6913,
    new_n6914, new_n6915, new_n6916, new_n6917, new_n6918, new_n6919,
    new_n6920, new_n6921, new_n6922, new_n6923, new_n6924, new_n6925,
    new_n6926, new_n6927, new_n6928, new_n6929, new_n6930, new_n6931,
    new_n6932, new_n6933, new_n6934, new_n6935, new_n6936, new_n6937_1,
    new_n6938, new_n6939, new_n6940, new_n6941, new_n6942, new_n6943,
    new_n6944, new_n6945, new_n6946, new_n6947, new_n6948, new_n6949,
    new_n6950, new_n6951, new_n6952, new_n6953, new_n6954, new_n6955,
    new_n6956, new_n6957, new_n6958, new_n6959, new_n6960, new_n6961,
    new_n6962, new_n6963, new_n6964, new_n6965, new_n6966, new_n6967,
    new_n6968, new_n6969, new_n6970, new_n6971, new_n6972, new_n6973,
    new_n6974, new_n6975, new_n6976, new_n6977, new_n6978, new_n6979,
    new_n6980, new_n6981, new_n6982, new_n6983, new_n6984, new_n6985,
    new_n6986, new_n6987, new_n6988, new_n6989, new_n6990, new_n6991,
    new_n6992, new_n6993, new_n6994, new_n6995, new_n6996, new_n6997,
    new_n6998, new_n6999, new_n7000, new_n7001, new_n7002, new_n7003,
    new_n7004, new_n7005, new_n7006, new_n7007, new_n7008, new_n7009,
    new_n7010, new_n7011, new_n7012, new_n7013, new_n7014, new_n7015,
    new_n7016, new_n7017, new_n7018, new_n7019, new_n7020, new_n7021,
    new_n7022, new_n7023, new_n7024, new_n7025, new_n7026, new_n7027,
    new_n7028, new_n7029, new_n7030, new_n7031, new_n7032, new_n7033,
    new_n7034_1, new_n7035, new_n7036, new_n7037, new_n7038, new_n7039,
    new_n7040, new_n7041, new_n7042, new_n7043, new_n7044, new_n7045,
    new_n7046, new_n7047, new_n7048, new_n7049, new_n7050, new_n7051,
    new_n7052, new_n7053, new_n7054, new_n7055, new_n7056, new_n7057,
    new_n7058, new_n7059, new_n7060, new_n7061_1, new_n7062, new_n7063,
    new_n7064, new_n7065, new_n7066, new_n7067, new_n7068, new_n7069,
    new_n7070, new_n7071, new_n7072, new_n7073, new_n7074, new_n7075,
    new_n7076, new_n7077, new_n7078, new_n7079, new_n7080, new_n7081,
    new_n7082, new_n7083, new_n7084, new_n7085, new_n7086, new_n7087,
    new_n7088, new_n7089, new_n7090, new_n7091, new_n7092, new_n7093,
    new_n7094, new_n7095, new_n7096, new_n7097, new_n7098, new_n7099,
    new_n7100, new_n7101, new_n7102, new_n7103, new_n7104, new_n7105,
    new_n7106, new_n7107, new_n7108, new_n7109, new_n7110, new_n7111_1,
    new_n7112, new_n7113_1, new_n7114, new_n7115, new_n7116, new_n7117,
    new_n7118, new_n7119, new_n7120, new_n7121, new_n7122, new_n7123,
    new_n7124, new_n7125, new_n7126, new_n7127, new_n7128, new_n7129,
    new_n7130, new_n7131, new_n7132_1, new_n7133, new_n7134, new_n7135,
    new_n7136, new_n7137, new_n7138, new_n7139, new_n7140, new_n7141,
    new_n7142, new_n7143, new_n7144, new_n7145, new_n7146, new_n7147,
    new_n7148, new_n7149, new_n7150, new_n7151, new_n7152, new_n7153,
    new_n7154, new_n7155, new_n7156, new_n7157, new_n7158, new_n7159,
    new_n7160, new_n7161_1, new_n7162, new_n7163, new_n7164, new_n7165,
    new_n7166, new_n7167, new_n7168, new_n7169, new_n7170, new_n7171,
    new_n7172, new_n7173, new_n7174, new_n7175, new_n7176, new_n7177,
    new_n7178, new_n7179, new_n7180, new_n7181, new_n7182, new_n7183,
    new_n7184, new_n7185, new_n7186, new_n7187, new_n7188, new_n7189,
    new_n7190, new_n7191, new_n7192, new_n7193, new_n7194, new_n7195,
    new_n7196, new_n7197, new_n7198, new_n7199, new_n7200, new_n7201,
    new_n7202, new_n7203, new_n7204, new_n7205, new_n7206, new_n7207,
    new_n7208, new_n7209, new_n7210, new_n7211, new_n7212, new_n7213,
    new_n7214, new_n7215, new_n7216, new_n7217, new_n7218, new_n7219,
    new_n7220, new_n7221, new_n7222, new_n7223, new_n7224, new_n7225,
    new_n7226, new_n7227, new_n7228, new_n7229, new_n7230, new_n7231,
    new_n7232, new_n7233, new_n7234, new_n7235, new_n7236, new_n7237,
    new_n7238, new_n7239, new_n7240, new_n7241_1, new_n7242, new_n7243,
    new_n7244, new_n7245, new_n7246, new_n7247, new_n7248, new_n7249,
    new_n7250, new_n7251, new_n7252, new_n7253, new_n7254, new_n7255,
    new_n7256, new_n7257, new_n7258, new_n7259, new_n7260, new_n7261,
    new_n7262, new_n7263, new_n7264, new_n7265, new_n7266, new_n7267,
    new_n7268, new_n7269, new_n7270, new_n7271, new_n7272, new_n7273,
    new_n7274, new_n7275, new_n7276, new_n7277, new_n7278, new_n7279,
    new_n7280, new_n7281, new_n7282, new_n7283, new_n7284, new_n7285,
    new_n7286, new_n7287, new_n7288, new_n7289, new_n7290, new_n7291,
    new_n7292, new_n7293, new_n7294, new_n7295, new_n7296, new_n7297,
    new_n7298, new_n7299, new_n7300, new_n7301, new_n7302, new_n7303,
    new_n7304, new_n7305, new_n7306, new_n7307, new_n7308, new_n7309,
    new_n7310, new_n7311, new_n7312, new_n7313, new_n7314, new_n7315,
    new_n7316, new_n7317, new_n7318, new_n7319, new_n7320, new_n7321,
    new_n7322, new_n7323, new_n7324, new_n7325, new_n7326, new_n7327,
    new_n7328, new_n7329, new_n7330, new_n7331, new_n7332, new_n7333,
    new_n7334, new_n7335, new_n7336, new_n7337, new_n7338, new_n7339,
    new_n7340, new_n7341, new_n7342, new_n7343, new_n7344, new_n7345,
    new_n7346, new_n7347, new_n7348, new_n7349, new_n7350, new_n7351,
    new_n7352, new_n7353, new_n7354, new_n7355, new_n7356, new_n7357,
    new_n7358, new_n7359, new_n7360, new_n7361, new_n7362, new_n7363,
    new_n7364, new_n7365, new_n7366, new_n7367, new_n7368, new_n7369,
    new_n7370, new_n7371, new_n7372, new_n7373, new_n7374_1, new_n7375,
    new_n7376, new_n7377, new_n7378, new_n7379, new_n7380, new_n7381,
    new_n7382, new_n7383, new_n7384, new_n7385, new_n7386, new_n7387,
    new_n7388, new_n7389, new_n7390, new_n7391, new_n7392, new_n7393,
    new_n7394, new_n7395, new_n7396, new_n7397, new_n7398, new_n7399,
    new_n7400, new_n7401, new_n7402, new_n7403, new_n7404, new_n7405,
    new_n7406, new_n7407, new_n7408, new_n7409, new_n7410, new_n7411_1,
    new_n7412, new_n7413, new_n7414, new_n7415, new_n7416, new_n7417,
    new_n7418, new_n7419, new_n7420, new_n7421, new_n7422, new_n7423,
    new_n7424, new_n7425, new_n7426, new_n7427, new_n7428, new_n7429,
    new_n7430, new_n7431, new_n7432, new_n7433, new_n7435, new_n7437,
    new_n7438, new_n7439, new_n7441, new_n7442, new_n7443, new_n7444,
    new_n7445, new_n7446, new_n7447, new_n7448, new_n7449, new_n7450,
    new_n7451, new_n7452, new_n7453, new_n7454, new_n7455, new_n7456,
    new_n7457, new_n7458, new_n7459, new_n7460, new_n7461, new_n7462,
    new_n7463, new_n7464, new_n7465, new_n7466, new_n7467, new_n7468,
    new_n7469, new_n7470, new_n7471, new_n7472, new_n7473, new_n7474,
    new_n7475, new_n7476, new_n7477, new_n7478, new_n7479, new_n7480,
    new_n7481, new_n7482, new_n7483, new_n7484, new_n7485, new_n7486,
    new_n7487, new_n7488, new_n7489, new_n7490, new_n7491, new_n7492,
    new_n7493, new_n7494, new_n7495, new_n7496, new_n7497, new_n7498,
    new_n7499, new_n7500, new_n7501, new_n7502, new_n7503, new_n7504,
    new_n7505, new_n7506, new_n7507, new_n7508, new_n7509, new_n7510,
    new_n7511, new_n7512, new_n7513, new_n7514, new_n7515, new_n7516,
    new_n7517, new_n7518, new_n7519, new_n7520, new_n7521, new_n7522,
    new_n7523, new_n7524, new_n7525, new_n7526, new_n7527, new_n7528,
    new_n7529_1, new_n7530, new_n7531, new_n7532, new_n7533, new_n7534,
    new_n7535, new_n7536, new_n7537, new_n7538, new_n7539, new_n7540,
    new_n7541, new_n7542, new_n7543, new_n7544, new_n7545, new_n7546,
    new_n7547, new_n7548, new_n7549, new_n7550, new_n7551, new_n7552,
    new_n7553_1, new_n7554, new_n7555, new_n7556, new_n7557, new_n7558,
    new_n7559, new_n7560, new_n7561, new_n7562, new_n7563, new_n7564,
    new_n7565, new_n7566, new_n7567, new_n7568, new_n7569, new_n7570,
    new_n7571, new_n7572, new_n7573, new_n7574, new_n7575, new_n7576,
    new_n7577, new_n7578, new_n7579, new_n7580, new_n7581, new_n7582_1,
    new_n7583, new_n7584, new_n7585, new_n7586, new_n7587, new_n7588,
    new_n7589, new_n7590, new_n7591, new_n7592, new_n7593, new_n7594,
    new_n7595, new_n7596, new_n7597, new_n7598, new_n7599, new_n7600,
    new_n7601, new_n7602, new_n7603, new_n7604, new_n7605, new_n7606,
    new_n7607, new_n7608, new_n7609, new_n7610, new_n7611, new_n7612,
    new_n7613, new_n7614, new_n7615, new_n7616, new_n7617, new_n7618,
    new_n7619, new_n7620, new_n7621, new_n7622, new_n7623, new_n7624,
    new_n7625, new_n7626, new_n7627, new_n7628, new_n7629, new_n7630,
    new_n7631, new_n7632, new_n7633, new_n7634, new_n7635, new_n7636,
    new_n7637, new_n7638, new_n7639, new_n7640, new_n7641, new_n7642,
    new_n7643, new_n7644, new_n7645, new_n7646, new_n7647, new_n7648,
    new_n7649, new_n7650, new_n7651, new_n7652, new_n7653, new_n7654,
    new_n7655, new_n7656, new_n7657, new_n7658, new_n7659_1, new_n7660,
    new_n7661, new_n7662, new_n7663, new_n7664, new_n7665, new_n7666,
    new_n7667, new_n7668, new_n7669, new_n7670, new_n7671, new_n7672,
    new_n7673, new_n7674, new_n7675, new_n7676, new_n7677, new_n7678,
    new_n7679, new_n7680, new_n7681, new_n7682, new_n7683, new_n7684,
    new_n7685, new_n7686, new_n7687_1, new_n7688, new_n7689, new_n7690,
    new_n7691, new_n7692, new_n7693, new_n7694, new_n7695, new_n7696,
    new_n7697, new_n7698, new_n7699, new_n7700, new_n7701, new_n7702,
    new_n7703, new_n7704, new_n7705, new_n7706, new_n7707, new_n7708,
    new_n7709, new_n7710, new_n7711, new_n7712, new_n7713, new_n7714,
    new_n7715_1, new_n7716, new_n7717, new_n7718, new_n7719, new_n7720_1,
    new_n7721, new_n7722, new_n7723, new_n7724, new_n7725, new_n7726,
    new_n7727, new_n7728, new_n7729_1, new_n7730, new_n7731, new_n7732,
    new_n7733, new_n7734, new_n7735, new_n7736, new_n7737, new_n7738,
    new_n7739, new_n7740, new_n7741, new_n7742, new_n7743, new_n7744,
    new_n7745, new_n7746, new_n7747, new_n7748, new_n7749, new_n7750,
    new_n7751, new_n7752, new_n7753, new_n7754, new_n7755_1, new_n7756,
    new_n7757, new_n7758, new_n7759, new_n7760, new_n7761, new_n7762,
    new_n7763, new_n7764, new_n7765, new_n7766, new_n7767, new_n7768,
    new_n7769, new_n7770, new_n7771, new_n7772_1, new_n7773, new_n7774,
    new_n7775, new_n7776, new_n7777, new_n7778, new_n7779, new_n7780,
    new_n7781, new_n7782, new_n7783, new_n7784, new_n7785, new_n7786,
    new_n7787, new_n7788, new_n7789, new_n7790_1, new_n7791, new_n7792,
    new_n7793, new_n7794, new_n7795, new_n7796, new_n7797, new_n7798,
    new_n7799, new_n7800, new_n7801, new_n7802, new_n7803, new_n7804,
    new_n7805, new_n7806, new_n7807, new_n7808, new_n7809, new_n7810,
    new_n7811, new_n7812_1, new_n7813, new_n7814, new_n7815, new_n7816,
    new_n7817, new_n7818, new_n7819, new_n7820, new_n7821, new_n7822,
    new_n7823, new_n7824, new_n7825, new_n7826, new_n7827, new_n7828,
    new_n7829, new_n7830, new_n7831, new_n7832, new_n7833, new_n7834,
    new_n7835, new_n7836, new_n7837, new_n7838, new_n7839, new_n7840,
    new_n7841, new_n7842, new_n7843, new_n7844, new_n7845, new_n7846,
    new_n7847, new_n7848, new_n7849, new_n7850, new_n7851, new_n7852,
    new_n7853, new_n7854, new_n7855, new_n7856, new_n7857, new_n7858_1,
    new_n7859, new_n7860_1, new_n7861, new_n7862, new_n7863, new_n7864,
    new_n7865, new_n7866, new_n7867, new_n7868, new_n7869, new_n7870,
    new_n7871, new_n7872, new_n7873, new_n7874, new_n7875, new_n7876,
    new_n7877, new_n7878, new_n7879, new_n7880, new_n7881, new_n7882,
    new_n7883, new_n7884, new_n7885, new_n7886, new_n7887, new_n7888,
    new_n7889, new_n7890, new_n7891, new_n7892, new_n7893, new_n7894,
    new_n7895, new_n7896, new_n7897, new_n7898, new_n7899, new_n7900,
    new_n7901, new_n7902, new_n7903, new_n7904, new_n7905, new_n7906,
    new_n7907, new_n7908, new_n7909, new_n7910, new_n7911, new_n7912,
    new_n7913, new_n7914, new_n7915, new_n7916, new_n7917, new_n7918,
    new_n7919, new_n7920, new_n7921, new_n7922, new_n7923, new_n7924,
    new_n7925, new_n7926, new_n7927, new_n7928, new_n7929, new_n7930,
    new_n7931, new_n7932, new_n7933, new_n7934, new_n7935, new_n7936,
    new_n7937, new_n7938, new_n7939, new_n7940, new_n7941, new_n7942,
    new_n7943, new_n7944, new_n7945, new_n7946, new_n7947, new_n7948,
    new_n7949, new_n7950, new_n7951, new_n7952, new_n7953, new_n7954,
    new_n7955, new_n7956, new_n7957, new_n7958, new_n7959, new_n7960,
    new_n7961, new_n7962, new_n7963, new_n7964, new_n7965, new_n7966,
    new_n7968_1, new_n7969, new_n7970, new_n7972, new_n7973, new_n7974_1,
    new_n7976, new_n7977, new_n7978, new_n7980, new_n7981, new_n7982,
    new_n7983, new_n7984, new_n7985, new_n7986, new_n7987, new_n7988,
    new_n7989, new_n7990, new_n7991, new_n7992, new_n7993, new_n7994,
    new_n7995, new_n7996, new_n7997, new_n7998, new_n7999, new_n8000,
    new_n8001, new_n8002, new_n8003, new_n8004, new_n8005, new_n8006,
    new_n8007, new_n8008, new_n8009, new_n8010, new_n8011, new_n8012,
    new_n8013, new_n8014, new_n8015, new_n8016, new_n8017, new_n8018,
    new_n8019, new_n8020, new_n8021, new_n8022, new_n8023, new_n8024,
    new_n8025, new_n8026, new_n8027, new_n8028, new_n8029, new_n8030,
    new_n8031, new_n8032, new_n8033, new_n8034, new_n8035, new_n8036,
    new_n8037, new_n8038, new_n8039, new_n8040, new_n8041, new_n8042,
    new_n8043, new_n8044, new_n8045, new_n8046, new_n8047, new_n8048,
    new_n8049, new_n8050, new_n8051, new_n8052, new_n8053, new_n8054,
    new_n8055, new_n8056, new_n8057, new_n8058, new_n8059, new_n8060,
    new_n8061, new_n8062, new_n8063, new_n8064, new_n8065, new_n8066,
    new_n8067, new_n8068, new_n8069, new_n8070, new_n8071, new_n8072,
    new_n8073, new_n8074, new_n8075, new_n8076, new_n8077, new_n8078,
    new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084,
    new_n8085, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090,
    new_n8091, new_n8092, new_n8093, new_n8094, new_n8095, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102,
    new_n8103, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8109, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114,
    new_n8115, new_n8116, new_n8117, new_n8118, new_n8119, new_n8120,
    new_n8121, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126,
    new_n8127, new_n8128, new_n8129, new_n8130, new_n8131, new_n8132,
    new_n8133, new_n8134, new_n8135, new_n8136, new_n8137, new_n8138,
    new_n8139_1, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144,
    new_n8145, new_n8146, new_n8147, new_n8148, new_n8149, new_n8150,
    new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156,
    new_n8157, new_n8158, new_n8159, new_n8160, new_n8161, new_n8162,
    new_n8163_1, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168,
    new_n8169, new_n8170, new_n8171, new_n8172_1, new_n8173, new_n8174,
    new_n8175, new_n8176, new_n8177, new_n8178, new_n8179, new_n8180,
    new_n8181, new_n8182, new_n8183_1, new_n8184, new_n8185, new_n8186,
    new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192,
    new_n8193, new_n8194, new_n8195, new_n8196, new_n8197, new_n8198,
    new_n8199, new_n8200, new_n8201, new_n8202, new_n8203, new_n8204,
    new_n8205, new_n8206, new_n8207, new_n8208, new_n8209, new_n8210,
    new_n8211, new_n8212, new_n8213, new_n8214, new_n8215, new_n8216,
    new_n8217, new_n8218, new_n8219_1, new_n8220, new_n8221, new_n8222,
    new_n8223, new_n8224, new_n8225, new_n8226, new_n8227, new_n8228_1,
    new_n8229, new_n8230_1, new_n8231, new_n8232, new_n8233_1, new_n8234,
    new_n8235, new_n8236, new_n8237, new_n8238, new_n8239, new_n8240,
    new_n8241, new_n8242, new_n8243, new_n8244, new_n8245, new_n8246,
    new_n8247, new_n8248, new_n8249, new_n8250, new_n8251, new_n8252,
    new_n8253, new_n8254, new_n8255, new_n8256, new_n8257, new_n8258,
    new_n8259, new_n8260, new_n8261, new_n8262, new_n8263, new_n8264,
    new_n8265_1, new_n8266, new_n8267, new_n8268, new_n8269, new_n8270,
    new_n8271, new_n8272, new_n8273, new_n8274, new_n8275, new_n8276,
    new_n8277, new_n8278, new_n8279, new_n8280, new_n8281, new_n8282,
    new_n8283, new_n8284, new_n8285, new_n8286, new_n8287, new_n8288,
    new_n8289, new_n8290_1, new_n8291, new_n8292, new_n8293, new_n8294,
    new_n8295, new_n8296, new_n8297, new_n8298, new_n8299, new_n8300,
    new_n8301, new_n8302, new_n8303, new_n8304, new_n8305, new_n8306,
    new_n8307, new_n8308_1, new_n8309, new_n8310, new_n8311, new_n8312,
    new_n8313, new_n8314, new_n8315, new_n8316, new_n8317, new_n8318,
    new_n8319, new_n8320, new_n8321, new_n8322, new_n8323, new_n8324,
    new_n8325, new_n8326, new_n8327, new_n8328, new_n8329, new_n8330,
    new_n8331, new_n8332_1, new_n8333, new_n8334, new_n8335, new_n8336_1,
    new_n8337, new_n8338, new_n8339, new_n8340, new_n8341, new_n8342,
    new_n8343, new_n8344, new_n8345, new_n8346, new_n8347, new_n8348,
    new_n8349, new_n8350, new_n8351, new_n8352, new_n8353, new_n8354,
    new_n8355, new_n8356, new_n8357, new_n8358, new_n8359, new_n8360,
    new_n8361, new_n8362, new_n8363, new_n8364, new_n8365, new_n8366,
    new_n8367, new_n8368, new_n8369, new_n8370, new_n8371, new_n8372,
    new_n8373, new_n8374, new_n8375, new_n8376, new_n8377, new_n8378,
    new_n8379, new_n8380, new_n8381, new_n8382, new_n8383, new_n8384,
    new_n8385, new_n8386, new_n8387, new_n8388, new_n8389, new_n8390,
    new_n8391, new_n8392, new_n8393, new_n8394, new_n8395, new_n8396,
    new_n8397, new_n8398, new_n8399, new_n8400, new_n8401, new_n8402,
    new_n8403, new_n8404, new_n8405, new_n8406, new_n8407, new_n8408,
    new_n8409, new_n8410, new_n8411, new_n8412, new_n8413, new_n8414,
    new_n8415, new_n8416, new_n8417, new_n8418, new_n8419, new_n8420,
    new_n8421, new_n8422, new_n8423, new_n8424, new_n8425, new_n8426,
    new_n8427, new_n8428, new_n8429, new_n8430, new_n8431, new_n8432,
    new_n8433, new_n8434, new_n8435, new_n8436, new_n8437, new_n8438,
    new_n8439, new_n8440, new_n8441, new_n8442, new_n8443, new_n8444,
    new_n8445, new_n8446, new_n8447, new_n8448, new_n8449, new_n8450,
    new_n8451, new_n8452, new_n8453, new_n8454, new_n8455, new_n8456,
    new_n8457, new_n8458, new_n8459, new_n8460, new_n8461, new_n8462,
    new_n8463, new_n8464, new_n8465, new_n8466_1, new_n8467, new_n8468_1,
    new_n8469, new_n8470, new_n8471, new_n8472, new_n8473, new_n8474,
    new_n8475, new_n8476, new_n8477, new_n8478, new_n8479, new_n8480,
    new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486,
    new_n8487, new_n8488, new_n8489, new_n8490, new_n8491, new_n8492,
    new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498,
    new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505, new_n8506_1, new_n8507, new_n8508, new_n8509, new_n8510,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516_1,
    new_n8517, new_n8518, new_n8519, new_n8520, new_n8521, new_n8522_1,
    new_n8523, new_n8524, new_n8525, new_n8526, new_n8527, new_n8528,
    new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534,
    new_n8535, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550, new_n8551, new_n8552,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8574, new_n8575, new_n8576,
    new_n8577, new_n8578, new_n8579, new_n8580, new_n8581, new_n8582,
    new_n8583, new_n8584, new_n8585, new_n8586, new_n8587, new_n8588,
    new_n8589, new_n8590, new_n8591, new_n8592, new_n8593, new_n8594,
    new_n8595, new_n8596, new_n8597, new_n8598, new_n8599, new_n8600,
    new_n8601, new_n8602, new_n8603, new_n8604, new_n8605, new_n8606,
    new_n8607, new_n8608, new_n8609, new_n8610, new_n8611, new_n8612,
    new_n8613, new_n8614, new_n8615, new_n8616, new_n8617, new_n8618,
    new_n8619, new_n8620, new_n8621, new_n8622, new_n8623, new_n8624,
    new_n8625, new_n8626, new_n8627, new_n8628, new_n8629, new_n8630,
    new_n8631, new_n8632, new_n8633, new_n8634, new_n8635, new_n8636,
    new_n8637, new_n8638, new_n8639, new_n8640, new_n8641, new_n8642,
    new_n8643, new_n8644, new_n8645, new_n8646, new_n8647, new_n8648,
    new_n8649, new_n8650, new_n8651, new_n8652, new_n8653, new_n8654,
    new_n8655, new_n8656, new_n8657, new_n8658, new_n8659, new_n8660,
    new_n8661, new_n8662, new_n8663, new_n8664, new_n8665, new_n8666,
    new_n8667, new_n8668, new_n8669, new_n8670, new_n8671, new_n8672,
    new_n8673, new_n8674, new_n8675, new_n8676, new_n8677, new_n8678,
    new_n8679, new_n8680, new_n8681, new_n8682, new_n8683, new_n8684,
    new_n8685, new_n8686, new_n8687, new_n8688, new_n8689, new_n8690,
    new_n8691, new_n8692, new_n8693, new_n8694, new_n8695, new_n8696,
    new_n8697, new_n8698, new_n8699, new_n8700, new_n8701_1, new_n8702,
    new_n8703, new_n8704, new_n8705, new_n8706, new_n8707, new_n8708,
    new_n8709, new_n8710, new_n8711, new_n8712, new_n8713, new_n8714,
    new_n8715, new_n8716_1, new_n8717, new_n8718, new_n8719, new_n8720,
    new_n8721, new_n8722, new_n8723, new_n8724, new_n8725, new_n8726,
    new_n8727, new_n8728, new_n8729, new_n8730, new_n8731, new_n8732,
    new_n8733, new_n8734, new_n8735, new_n8736, new_n8737, new_n8738,
    new_n8739, new_n8740, new_n8741, new_n8742, new_n8743, new_n8744,
    new_n8745, new_n8746, new_n8747, new_n8748, new_n8749, new_n8750,
    new_n8751, new_n8752, new_n8753, new_n8754, new_n8755, new_n8756,
    new_n8757, new_n8758, new_n8759, new_n8760, new_n8761, new_n8762,
    new_n8763, new_n8764, new_n8765, new_n8766, new_n8767, new_n8768_1,
    new_n8769, new_n8770, new_n8771, new_n8772, new_n8773, new_n8774,
    new_n8775, new_n8776, new_n8777, new_n8778, new_n8779, new_n8780,
    new_n8781, new_n8782, new_n8783, new_n8784, new_n8785, new_n8786,
    new_n8787, new_n8788, new_n8789, new_n8790, new_n8791, new_n8792,
    new_n8793, new_n8794, new_n8795, new_n8796, new_n8797, new_n8798,
    new_n8799, new_n8800, new_n8801, new_n8802, new_n8803, new_n8804,
    new_n8805, new_n8806, new_n8807, new_n8808, new_n8809, new_n8810,
    new_n8811, new_n8812, new_n8813, new_n8814, new_n8815, new_n8816,
    new_n8817, new_n8818, new_n8819, new_n8820_1, new_n8821, new_n8822,
    new_n8823, new_n8824, new_n8825, new_n8826, new_n8827, new_n8828,
    new_n8829, new_n8830, new_n8831, new_n8832, new_n8833, new_n8834,
    new_n8835, new_n8836, new_n8837, new_n8838, new_n8839, new_n8840,
    new_n8841, new_n8842, new_n8843, new_n8844, new_n8845, new_n8846,
    new_n8847, new_n8848, new_n8849, new_n8850, new_n8851, new_n8852,
    new_n8853, new_n8854, new_n8855, new_n8856, new_n8857, new_n8858,
    new_n8859_1, new_n8860_1, new_n8861, new_n8862, new_n8863, new_n8864,
    new_n8865, new_n8866, new_n8867, new_n8868, new_n8869, new_n8870,
    new_n8871, new_n8872, new_n8873, new_n8874, new_n8875, new_n8876,
    new_n8877, new_n8878, new_n8879, new_n8880, new_n8881, new_n8882,
    new_n8883, new_n8884, new_n8885, new_n8886, new_n8887, new_n8888,
    new_n8889, new_n8890, new_n8891, new_n8892, new_n8893, new_n8894,
    new_n8895, new_n8896, new_n8897, new_n8898, new_n8899, new_n8900,
    new_n8901, new_n8902, new_n8903, new_n8904, new_n8905, new_n8906,
    new_n8907, new_n8908, new_n8909, new_n8910, new_n8911, new_n8912,
    new_n8913, new_n8914, new_n8915, new_n8916, new_n8917, new_n8918,
    new_n8919, new_n8920, new_n8921, new_n8922, new_n8923, new_n8924,
    new_n8925, new_n8927, new_n8928, new_n8929, new_n8931, new_n8932,
    new_n8933, new_n8934, new_n8935, new_n8936, new_n8937, new_n8938,
    new_n8939, new_n8940_1, new_n8941, new_n8942, new_n8943, new_n8944,
    new_n8945, new_n8946, new_n8947, new_n8948, new_n8949, new_n8950,
    new_n8951, new_n8952, new_n8953, new_n8954, new_n8955, new_n8956,
    new_n8957, new_n8958, new_n8959, new_n8960, new_n8961, new_n8962,
    new_n8963, new_n8964, new_n8965, new_n8966, new_n8967, new_n8968,
    new_n8969, new_n8970, new_n8971, new_n8972, new_n8973, new_n8974,
    new_n8975, new_n8976, new_n8977, new_n8978, new_n8980, new_n8981,
    new_n8982, new_n8984, new_n8985, new_n8986, new_n8988, new_n8990,
    new_n8991, new_n8992, new_n8994, new_n8995, new_n8996, new_n8998,
    new_n8999, new_n9000, new_n9002, new_n9003, new_n9004, new_n9005,
    new_n9006, new_n9007, new_n9008, new_n9009, new_n9010, new_n9011,
    new_n9012, new_n9013, new_n9014, new_n9015, new_n9016, new_n9017,
    new_n9018, new_n9019, new_n9020, new_n9021, new_n9022, new_n9023,
    new_n9024, new_n9025, new_n9026, new_n9027, new_n9028, new_n9029,
    new_n9030, new_n9031, new_n9032, new_n9033, new_n9034, new_n9035,
    new_n9036, new_n9037, new_n9038, new_n9039, new_n9040, new_n9041_1,
    new_n9042, new_n9043, new_n9044, new_n9045, new_n9046, new_n9047,
    new_n9048, new_n9049, new_n9050, new_n9051, new_n9052, new_n9053,
    new_n9054, new_n9055, new_n9056, new_n9057, new_n9058, new_n9059,
    new_n9060, new_n9061, new_n9062, new_n9063, new_n9064, new_n9065,
    new_n9066, new_n9067, new_n9068, new_n9069, new_n9070, new_n9071,
    new_n9072, new_n9073, new_n9074, new_n9075, new_n9076, new_n9077,
    new_n9078, new_n9079, new_n9080, new_n9081, new_n9082, new_n9083,
    new_n9084, new_n9085, new_n9086, new_n9087, new_n9088, new_n9089,
    new_n9090, new_n9091, new_n9092, new_n9093_1, new_n9094, new_n9095,
    new_n9096, new_n9097, new_n9098, new_n9099, new_n9100_1, new_n9101,
    new_n9102, new_n9103, new_n9104, new_n9105, new_n9106, new_n9107,
    new_n9108, new_n9109, new_n9110, new_n9111, new_n9112, new_n9113,
    new_n9114, new_n9115, new_n9116, new_n9117, new_n9118, new_n9119,
    new_n9120, new_n9121, new_n9122, new_n9123, new_n9124, new_n9125,
    new_n9126, new_n9127, new_n9128, new_n9129, new_n9130, new_n9131,
    new_n9132, new_n9133, new_n9134, new_n9135, new_n9136, new_n9137,
    new_n9138, new_n9139, new_n9140, new_n9141, new_n9142, new_n9143,
    new_n9144, new_n9145, new_n9146, new_n9147, new_n9148, new_n9149,
    new_n9150, new_n9151, new_n9152, new_n9153, new_n9154, new_n9155,
    new_n9156, new_n9157, new_n9158, new_n9159, new_n9160, new_n9161,
    new_n9162, new_n9163, new_n9164, new_n9165, new_n9166, new_n9167,
    new_n9168, new_n9169, new_n9170, new_n9171, new_n9172, new_n9173,
    new_n9174, new_n9175, new_n9176, new_n9177, new_n9178, new_n9179,
    new_n9180, new_n9181, new_n9182, new_n9183, new_n9184, new_n9185,
    new_n9186, new_n9187_1, new_n9188, new_n9189, new_n9190, new_n9191,
    new_n9192, new_n9193, new_n9194, new_n9195, new_n9196, new_n9197,
    new_n9198, new_n9199, new_n9200, new_n9201, new_n9202, new_n9203,
    new_n9204, new_n9205, new_n9206, new_n9207, new_n9208, new_n9209,
    new_n9210, new_n9211, new_n9212, new_n9213, new_n9214, new_n9215,
    new_n9216_1, new_n9217, new_n9218, new_n9219, new_n9220, new_n9221,
    new_n9222, new_n9223, new_n9224, new_n9225, new_n9226, new_n9227,
    new_n9228, new_n9229, new_n9230, new_n9231, new_n9232, new_n9233,
    new_n9234, new_n9235, new_n9236, new_n9237, new_n9238, new_n9239,
    new_n9240, new_n9241, new_n9242, new_n9243, new_n9244, new_n9245,
    new_n9246, new_n9247, new_n9248, new_n9249, new_n9250, new_n9251,
    new_n9252, new_n9253, new_n9254, new_n9255, new_n9256, new_n9257,
    new_n9258, new_n9259, new_n9260, new_n9261, new_n9262, new_n9263,
    new_n9264, new_n9265, new_n9266, new_n9267, new_n9268, new_n9269,
    new_n9270, new_n9271, new_n9272, new_n9273, new_n9274, new_n9275,
    new_n9276, new_n9277, new_n9278, new_n9279, new_n9280, new_n9281,
    new_n9282, new_n9283, new_n9284, new_n9285, new_n9286, new_n9287,
    new_n9288, new_n9289, new_n9290, new_n9291, new_n9292, new_n9293,
    new_n9294, new_n9295, new_n9296, new_n9297, new_n9298, new_n9299,
    new_n9300_1, new_n9301, new_n9302, new_n9303, new_n9304, new_n9305,
    new_n9306, new_n9307, new_n9308, new_n9309, new_n9310, new_n9311,
    new_n9312, new_n9313, new_n9314, new_n9315, new_n9316, new_n9317,
    new_n9318, new_n9319, new_n9320, new_n9321, new_n9322, new_n9323,
    new_n9324, new_n9325, new_n9326, new_n9327, new_n9328, new_n9329_1,
    new_n9330, new_n9331, new_n9332, new_n9333, new_n9334, new_n9335,
    new_n9336, new_n9337, new_n9338, new_n9339, new_n9340, new_n9341,
    new_n9342, new_n9343, new_n9344, new_n9345, new_n9346, new_n9347,
    new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353_1,
    new_n9354, new_n9356, new_n9357, new_n9358, new_n9360, new_n9361,
    new_n9362, new_n9364, new_n9365, new_n9366, new_n9368, new_n9369,
    new_n9370, new_n9372, new_n9373, new_n9374, new_n9376, new_n9377,
    new_n9378, new_n9380, new_n9381, new_n9382, new_n9383, new_n9384,
    new_n9385, new_n9386, new_n9387, new_n9388, new_n9389, new_n9390,
    new_n9391, new_n9392, new_n9393, new_n9394, new_n9395, new_n9396,
    new_n9397, new_n9398, new_n9399, new_n9400, new_n9401, new_n9402,
    new_n9403, new_n9404, new_n9405, new_n9406, new_n9407, new_n9408,
    new_n9409, new_n9410, new_n9411, new_n9412, new_n9413, new_n9414,
    new_n9415, new_n9416, new_n9417, new_n9418, new_n9419, new_n9420,
    new_n9421, new_n9422, new_n9423, new_n9424, new_n9425, new_n9426,
    new_n9427, new_n9428, new_n9429, new_n9430, new_n9431, new_n9432,
    new_n9433, new_n9434, new_n9435, new_n9436, new_n9437, new_n9438,
    new_n9439, new_n9440, new_n9441, new_n9442, new_n9443, new_n9444,
    new_n9445, new_n9446, new_n9447, new_n9448, new_n9449, new_n9450,
    new_n9451, new_n9452, new_n9453, new_n9454, new_n9455, new_n9456,
    new_n9457, new_n9458, new_n9459, new_n9460, new_n9461, new_n9462,
    new_n9463, new_n9464, new_n9465, new_n9466, new_n9467, new_n9468,
    new_n9469, new_n9470, new_n9471, new_n9472, new_n9473, new_n9474,
    new_n9475_1, new_n9476, new_n9477, new_n9478, new_n9479, new_n9480,
    new_n9481, new_n9482, new_n9483, new_n9484, new_n9485, new_n9486,
    new_n9487, new_n9488, new_n9489, new_n9490, new_n9491, new_n9492,
    new_n9493, new_n9494, new_n9495, new_n9496, new_n9497, new_n9498,
    new_n9499, new_n9500, new_n9501, new_n9502, new_n9503, new_n9504,
    new_n9505, new_n9506, new_n9507, new_n9508, new_n9509, new_n9510,
    new_n9511, new_n9512, new_n9513, new_n9514, new_n9515, new_n9516,
    new_n9517, new_n9518, new_n9519, new_n9520, new_n9521, new_n9522,
    new_n9523, new_n9524, new_n9525, new_n9526, new_n9527, new_n9528_1,
    new_n9529, new_n9530, new_n9531_1, new_n9532, new_n9533, new_n9534,
    new_n9535, new_n9536, new_n9537, new_n9538, new_n9539, new_n9540,
    new_n9541, new_n9542, new_n9543, new_n9544, new_n9545, new_n9546,
    new_n9547, new_n9548, new_n9549, new_n9550, new_n9551, new_n9552,
    new_n9553, new_n9554, new_n9555, new_n9556, new_n9557, new_n9558,
    new_n9559, new_n9560, new_n9561, new_n9562, new_n9563, new_n9564,
    new_n9565, new_n9566, new_n9567, new_n9568, new_n9569, new_n9570_1,
    new_n9571, new_n9572, new_n9573, new_n9574, new_n9575, new_n9576,
    new_n9577, new_n9578, new_n9579, new_n9580, new_n9581, new_n9582,
    new_n9583, new_n9584, new_n9585, new_n9586, new_n9587, new_n9588,
    new_n9589, new_n9590, new_n9591_1, new_n9592, new_n9593, new_n9594,
    new_n9595, new_n9596, new_n9597, new_n9598, new_n9599, new_n9600,
    new_n9601, new_n9602, new_n9603, new_n9604, new_n9605, new_n9606,
    new_n9607, new_n9608, new_n9609, new_n9610, new_n9611, new_n9612,
    new_n9613, new_n9614, new_n9615, new_n9616, new_n9617, new_n9618,
    new_n9619, new_n9620_1, new_n9621, new_n9622, new_n9623, new_n9624,
    new_n9625, new_n9626, new_n9627, new_n9628, new_n9629, new_n9630,
    new_n9631, new_n9632, new_n9633, new_n9634, new_n9635, new_n9636,
    new_n9637, new_n9638, new_n9639, new_n9640, new_n9641, new_n9642,
    new_n9643, new_n9644, new_n9645, new_n9646, new_n9647, new_n9648,
    new_n9649, new_n9650, new_n9651, new_n9652, new_n9653, new_n9654,
    new_n9655, new_n9656, new_n9657, new_n9658, new_n9659, new_n9660,
    new_n9661, new_n9662, new_n9663, new_n9664, new_n9665, new_n9666,
    new_n9667, new_n9668, new_n9669_1, new_n9670, new_n9671, new_n9672,
    new_n9673, new_n9674, new_n9675, new_n9676, new_n9677, new_n9678,
    new_n9679, new_n9680, new_n9681, new_n9682, new_n9683, new_n9684,
    new_n9685, new_n9686, new_n9687, new_n9688, new_n9689, new_n9690,
    new_n9691, new_n9692, new_n9693, new_n9694, new_n9695, new_n9696,
    new_n9697, new_n9698, new_n9699, new_n9700, new_n9701, new_n9702,
    new_n9703, new_n9704, new_n9705, new_n9706, new_n9707, new_n9708,
    new_n9709, new_n9710, new_n9711, new_n9712, new_n9713, new_n9714,
    new_n9715, new_n9716, new_n9717, new_n9718, new_n9719, new_n9720,
    new_n9721, new_n9722, new_n9723, new_n9724, new_n9725, new_n9726,
    new_n9727, new_n9728, new_n9729, new_n9730, new_n9731, new_n9732_1,
    new_n9733, new_n9734, new_n9735, new_n9736, new_n9737, new_n9738,
    new_n9739, new_n9740, new_n9741, new_n9742, new_n9743, new_n9744,
    new_n9745, new_n9746, new_n9747_1, new_n9748, new_n9749, new_n9750,
    new_n9751, new_n9752, new_n9753, new_n9754, new_n9755, new_n9756,
    new_n9757, new_n9758, new_n9759, new_n9760, new_n9761, new_n9762,
    new_n9763, new_n9764, new_n9765, new_n9766, new_n9767, new_n9768,
    new_n9769, new_n9770, new_n9771, new_n9772, new_n9773, new_n9774,
    new_n9775, new_n9776, new_n9777, new_n9778, new_n9779, new_n9780,
    new_n9781, new_n9782, new_n9783, new_n9784, new_n9785, new_n9786,
    new_n9787, new_n9788, new_n9789, new_n9790, new_n9791, new_n9792,
    new_n9793, new_n9794, new_n9795, new_n9796, new_n9797, new_n9798,
    new_n9799, new_n9800, new_n9801, new_n9802, new_n9803, new_n9804,
    new_n9805, new_n9806, new_n9807, new_n9808, new_n9809, new_n9810,
    new_n9811, new_n9812, new_n9813, new_n9814, new_n9815, new_n9816,
    new_n9817, new_n9818, new_n9819, new_n9820, new_n9822, new_n9823,
    new_n9824, new_n9825, new_n9826, new_n9827, new_n9828, new_n9829,
    new_n9830, new_n9831, new_n9832, new_n9833, new_n9834, new_n9835,
    new_n9836, new_n9837, new_n9838, new_n9839, new_n9840, new_n9841,
    new_n9842, new_n9843, new_n9844, new_n9845, new_n9846_1, new_n9847,
    new_n9848, new_n9849, new_n9850, new_n9851, new_n9852, new_n9853,
    new_n9854, new_n9855, new_n9856, new_n9857, new_n9858, new_n9859,
    new_n9860, new_n9861, new_n9862, new_n9863, new_n9864, new_n9865,
    new_n9866_1, new_n9867, new_n9868, new_n9869, new_n9870, new_n9871,
    new_n9872_1, new_n9873, new_n9874, new_n9875, new_n9876, new_n9877,
    new_n9878, new_n9879, new_n9880, new_n9881, new_n9882, new_n9883,
    new_n9884, new_n9885, new_n9886, new_n9887_1, new_n9888, new_n9889,
    new_n9890, new_n9891, new_n9892, new_n9893, new_n9894, new_n9895,
    new_n9896, new_n9897, new_n9898, new_n9899, new_n9900, new_n9901,
    new_n9902, new_n9903, new_n9904, new_n9905, new_n9906_1, new_n9907,
    new_n9908, new_n9909, new_n9910, new_n9911, new_n9912, new_n9913,
    new_n9914, new_n9915_1, new_n9916, new_n9917, new_n9918, new_n9919,
    new_n9920, new_n9921, new_n9922, new_n9923, new_n9924, new_n9925,
    new_n9926, new_n9927, new_n9928, new_n9929, new_n9930, new_n9931,
    new_n9932, new_n9933, new_n9934, new_n9935, new_n9936, new_n9937,
    new_n9938, new_n9939, new_n9940, new_n9941, new_n9942, new_n9943,
    new_n9944, new_n9945, new_n9946, new_n9947, new_n9948, new_n9949,
    new_n9950, new_n9951, new_n9952, new_n9953, new_n9954, new_n9955,
    new_n9956, new_n9957, new_n9958, new_n9959, new_n9960, new_n9961,
    new_n9962, new_n9963, new_n9964, new_n9965, new_n9966, new_n9967,
    new_n9968, new_n9969, new_n9970, new_n9971, new_n9972, new_n9973,
    new_n9974, new_n9975, new_n9976, new_n9977, new_n9978, new_n9979,
    new_n9980, new_n9981, new_n9982, new_n9983, new_n9984, new_n9985,
    new_n9986, new_n9987, new_n9988, new_n9989, new_n9990, new_n9991,
    new_n9992, new_n9993, new_n9994, new_n9995, new_n9996, new_n9997,
    new_n9998, new_n9999, new_n10000, new_n10001, new_n10002, new_n10003,
    new_n10004, new_n10005, new_n10006, new_n10007, new_n10008, new_n10009,
    new_n10010, new_n10011, new_n10012, new_n10013, new_n10014, new_n10015,
    new_n10016, new_n10017, new_n10018, new_n10019, new_n10020, new_n10021,
    new_n10022, new_n10023, new_n10024, new_n10025, new_n10026, new_n10027,
    new_n10028, new_n10029, new_n10030, new_n10031, new_n10032, new_n10033,
    new_n10034, new_n10035, new_n10036, new_n10037, new_n10038, new_n10039,
    new_n10040, new_n10041, new_n10042, new_n10043, new_n10044, new_n10045,
    new_n10046, new_n10047, new_n10048, new_n10049, new_n10050, new_n10051,
    new_n10052, new_n10053, new_n10054, new_n10055, new_n10056, new_n10057,
    new_n10058, new_n10059, new_n10060, new_n10061, new_n10062,
    new_n10063_1, new_n10064, new_n10065, new_n10067, new_n10069,
    new_n10070, new_n10071, new_n10073, new_n10074, new_n10075, new_n10077,
    new_n10078, new_n10079, new_n10081, new_n10082, new_n10083, new_n10085,
    new_n10086, new_n10087, new_n10089, new_n10090, new_n10091, new_n10092,
    new_n10093, new_n10094, new_n10095, new_n10096, new_n10097, new_n10098,
    new_n10099, new_n10100, new_n10101_1, new_n10102, new_n10103,
    new_n10104, new_n10105, new_n10106, new_n10107, new_n10108, new_n10109,
    new_n10110, new_n10111, new_n10112, new_n10113_1, new_n10114,
    new_n10115, new_n10116, new_n10117, new_n10118, new_n10119, new_n10120,
    new_n10121, new_n10122_1, new_n10123, new_n10124, new_n10125,
    new_n10126, new_n10127, new_n10128, new_n10129, new_n10130, new_n10131,
    new_n10132, new_n10133, new_n10134, new_n10135, new_n10136, new_n10137,
    new_n10138, new_n10139, new_n10140, new_n10141, new_n10142_1,
    new_n10143, new_n10144, new_n10145, new_n10146, new_n10147, new_n10148,
    new_n10149, new_n10150, new_n10151, new_n10152, new_n10153, new_n10154,
    new_n10155, new_n10156, new_n10157, new_n10158, new_n10159, new_n10160,
    new_n10161, new_n10162_1, new_n10163, new_n10164, new_n10165,
    new_n10166, new_n10167, new_n10168_1, new_n10169, new_n10170,
    new_n10171, new_n10172, new_n10173, new_n10174, new_n10175, new_n10176,
    new_n10177, new_n10178, new_n10179, new_n10180, new_n10181, new_n10182,
    new_n10183, new_n10184, new_n10185, new_n10186, new_n10187, new_n10188,
    new_n10189, new_n10190, new_n10191, new_n10192, new_n10193, new_n10194,
    new_n10195, new_n10196, new_n10197, new_n10198, new_n10199, new_n10200,
    new_n10201, new_n10202, new_n10203, new_n10204, new_n10205, new_n10206,
    new_n10207, new_n10208, new_n10209, new_n10210, new_n10211, new_n10212,
    new_n10213, new_n10214, new_n10215, new_n10216, new_n10217, new_n10218,
    new_n10219, new_n10220, new_n10221, new_n10222, new_n10223, new_n10224,
    new_n10225, new_n10226, new_n10227, new_n10228, new_n10229, new_n10230,
    new_n10231, new_n10232, new_n10233, new_n10234, new_n10235, new_n10236,
    new_n10237, new_n10238, new_n10239, new_n10240, new_n10241, new_n10242,
    new_n10243_1, new_n10244, new_n10245, new_n10246, new_n10247,
    new_n10248, new_n10249, new_n10250, new_n10251, new_n10252, new_n10253,
    new_n10254, new_n10255, new_n10256, new_n10257, new_n10258, new_n10259,
    new_n10260, new_n10261, new_n10262, new_n10263, new_n10265, new_n10266,
    new_n10267, new_n10268, new_n10269, new_n10270, new_n10271, new_n10272,
    new_n10273, new_n10274, new_n10275, new_n10276, new_n10277, new_n10278,
    new_n10279, new_n10280, new_n10281, new_n10282, new_n10283, new_n10284,
    new_n10285, new_n10286, new_n10287, new_n10288, new_n10289, new_n10290,
    new_n10291, new_n10292, new_n10293, new_n10294, new_n10295, new_n10296,
    new_n10297, new_n10298, new_n10299, new_n10300, new_n10301, new_n10302,
    new_n10303, new_n10304, new_n10305, new_n10306, new_n10307, new_n10308,
    new_n10309, new_n10310, new_n10311, new_n10312, new_n10313, new_n10314,
    new_n10315, new_n10316, new_n10317, new_n10318, new_n10319, new_n10320,
    new_n10321, new_n10322, new_n10323, new_n10324, new_n10325, new_n10326,
    new_n10327, new_n10328, new_n10329, new_n10330, new_n10331, new_n10332,
    new_n10333, new_n10334, new_n10335, new_n10336, new_n10337, new_n10338,
    new_n10339, new_n10340, new_n10341, new_n10342, new_n10343, new_n10344,
    new_n10345, new_n10346, new_n10347, new_n10348, new_n10349, new_n10350,
    new_n10351, new_n10353, new_n10354, new_n10355, new_n10357, new_n10358,
    new_n10359, new_n10361, new_n10362, new_n10363, new_n10365, new_n10366,
    new_n10367, new_n10369, new_n10370, new_n10371, new_n10372, new_n10373,
    new_n10374, new_n10375, new_n10376, new_n10377, new_n10378, new_n10379,
    new_n10380, new_n10381, new_n10382, new_n10383, new_n10384, new_n10385,
    new_n10386, new_n10387, new_n10388, new_n10389, new_n10390, new_n10391,
    new_n10392, new_n10393, new_n10394, new_n10395, new_n10396, new_n10397,
    new_n10398, new_n10399, new_n10400, new_n10401, new_n10402, new_n10403,
    new_n10404, new_n10405, new_n10406, new_n10407, new_n10408_1,
    new_n10409, new_n10410, new_n10411, new_n10412, new_n10413, new_n10414,
    new_n10415, new_n10416_1, new_n10417, new_n10418, new_n10419,
    new_n10420, new_n10421, new_n10422, new_n10423, new_n10424, new_n10425,
    new_n10426, new_n10427, new_n10428, new_n10429, new_n10430, new_n10431,
    new_n10432, new_n10433, new_n10434, new_n10435, new_n10436, new_n10437,
    new_n10438, new_n10439, new_n10440, new_n10441, new_n10442, new_n10443,
    new_n10444, new_n10445, new_n10446, new_n10447, new_n10448, new_n10449,
    new_n10450, new_n10451_1, new_n10452, new_n10453_1, new_n10454,
    new_n10455, new_n10456, new_n10457, new_n10458, new_n10459, new_n10460,
    new_n10461, new_n10462, new_n10463, new_n10464, new_n10465, new_n10466,
    new_n10467, new_n10468, new_n10469, new_n10470, new_n10471, new_n10472,
    new_n10473, new_n10474, new_n10475, new_n10476, new_n10477, new_n10478,
    new_n10479, new_n10480, new_n10481, new_n10482, new_n10483, new_n10484,
    new_n10485, new_n10486, new_n10487, new_n10488, new_n10489, new_n10490,
    new_n10491, new_n10492, new_n10493, new_n10494, new_n10495, new_n10496,
    new_n10497, new_n10498, new_n10499, new_n10500, new_n10501, new_n10502,
    new_n10503, new_n10504, new_n10505, new_n10506, new_n10507, new_n10508,
    new_n10509, new_n10510, new_n10511, new_n10512, new_n10513, new_n10514,
    new_n10515, new_n10516, new_n10517, new_n10518, new_n10519, new_n10520,
    new_n10521, new_n10522_1, new_n10523, new_n10524_1, new_n10525,
    new_n10526, new_n10527, new_n10528, new_n10529, new_n10530, new_n10531,
    new_n10532, new_n10533, new_n10534, new_n10535, new_n10536, new_n10537,
    new_n10538, new_n10539, new_n10540, new_n10541, new_n10542, new_n10543,
    new_n10544, new_n10545, new_n10546, new_n10547, new_n10548, new_n10549,
    new_n10550, new_n10551, new_n10552, new_n10553, new_n10554, new_n10555,
    new_n10556, new_n10557, new_n10558, new_n10559, new_n10560_1,
    new_n10561, new_n10562, new_n10563, new_n10564, new_n10565, new_n10566,
    new_n10567, new_n10568, new_n10569, new_n10570, new_n10571, new_n10573,
    new_n10574, new_n10575, new_n10577, new_n10578, new_n10579, new_n10581,
    new_n10582, new_n10583, new_n10585, new_n10586, new_n10587, new_n10588,
    new_n10589, new_n10590, new_n10591, new_n10592, new_n10593,
    new_n10594_1, new_n10595, new_n10596, new_n10597, new_n10598,
    new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604,
    new_n10605, new_n10606_1, new_n10607, new_n10608, new_n10609,
    new_n10610, new_n10611, new_n10612, new_n10613, new_n10614, new_n10615,
    new_n10616, new_n10617, new_n10618, new_n10619, new_n10620, new_n10621,
    new_n10622, new_n10623, new_n10624, new_n10625, new_n10626, new_n10627,
    new_n10628_1, new_n10629, new_n10630, new_n10631, new_n10632,
    new_n10633, new_n10634, new_n10635, new_n10636, new_n10637, new_n10638,
    new_n10639, new_n10640, new_n10641, new_n10642_1, new_n10643,
    new_n10644, new_n10645, new_n10646, new_n10647, new_n10648, new_n10649,
    new_n10650, new_n10651, new_n10652, new_n10653, new_n10654, new_n10655,
    new_n10656, new_n10657_1, new_n10658, new_n10659, new_n10660,
    new_n10661, new_n10662, new_n10663, new_n10664, new_n10665, new_n10666,
    new_n10667, new_n10668, new_n10669, new_n10670, new_n10671, new_n10672,
    new_n10673, new_n10674, new_n10675, new_n10676, new_n10677, new_n10678,
    new_n10679, new_n10680, new_n10681, new_n10682, new_n10683, new_n10684,
    new_n10685, new_n10686, new_n10687, new_n10688, new_n10689, new_n10690,
    new_n10691, new_n10692, new_n10693, new_n10694, new_n10695, new_n10696,
    new_n10697, new_n10698, new_n10699, new_n10700, new_n10701, new_n10702,
    new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708,
    new_n10709, new_n10710, new_n10711, new_n10712, new_n10713, new_n10714,
    new_n10715, new_n10716, new_n10717, new_n10718, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736_1, new_n10737,
    new_n10738, new_n10739, new_n10740, new_n10741, new_n10742, new_n10743,
    new_n10744, new_n10745, new_n10746, new_n10747, new_n10748, new_n10749,
    new_n10750, new_n10751, new_n10752, new_n10753, new_n10754, new_n10755,
    new_n10756, new_n10757, new_n10758, new_n10759, new_n10760, new_n10761,
    new_n10762, new_n10763, new_n10764, new_n10765, new_n10766, new_n10767,
    new_n10768, new_n10769, new_n10770_1, new_n10771, new_n10772,
    new_n10773, new_n10774, new_n10775, new_n10776, new_n10777, new_n10778,
    new_n10779, new_n10780, new_n10781, new_n10782, new_n10783, new_n10784,
    new_n10785, new_n10786, new_n10787, new_n10788, new_n10789, new_n10790,
    new_n10791, new_n10792, new_n10793, new_n10794, new_n10795, new_n10796,
    new_n10797_1, new_n10798, new_n10799, new_n10800, new_n10801,
    new_n10802, new_n10803, new_n10804, new_n10805_1, new_n10806,
    new_n10807, new_n10808, new_n10809, new_n10810, new_n10811, new_n10812,
    new_n10813, new_n10814, new_n10815, new_n10816, new_n10817, new_n10818,
    new_n10819, new_n10820, new_n10821, new_n10822, new_n10823, new_n10824,
    new_n10825, new_n10826, new_n10827, new_n10828, new_n10829, new_n10830,
    new_n10831, new_n10832, new_n10833, new_n10834, new_n10835, new_n10836,
    new_n10837, new_n10838, new_n10839, new_n10840, new_n10841, new_n10842,
    new_n10843, new_n10844, new_n10845, new_n10846, new_n10847, new_n10848,
    new_n10849, new_n10850, new_n10851, new_n10852, new_n10853, new_n10854,
    new_n10855, new_n10856, new_n10857, new_n10858, new_n10859, new_n10860,
    new_n10861, new_n10862, new_n10863, new_n10864, new_n10865,
    new_n10866_1, new_n10867, new_n10868, new_n10869, new_n10870,
    new_n10871, new_n10872, new_n10873, new_n10874_1, new_n10875,
    new_n10876, new_n10877, new_n10878, new_n10879, new_n10880, new_n10881,
    new_n10882, new_n10883, new_n10884, new_n10885, new_n10886, new_n10887,
    new_n10888, new_n10889, new_n10890, new_n10891, new_n10892, new_n10893,
    new_n10894, new_n10895, new_n10896, new_n10897, new_n10898, new_n10899,
    new_n10900, new_n10901, new_n10902, new_n10903, new_n10904, new_n10905,
    new_n10906, new_n10907, new_n10908_1, new_n10909, new_n10910,
    new_n10911, new_n10912, new_n10913, new_n10914, new_n10915, new_n10916,
    new_n10917, new_n10918, new_n10919, new_n10920, new_n10921, new_n10922,
    new_n10923, new_n10924, new_n10925, new_n10926, new_n10927, new_n10928,
    new_n10929, new_n10930, new_n10931, new_n10932, new_n10933, new_n10934,
    new_n10935, new_n10936, new_n10937, new_n10938, new_n10939, new_n10940,
    new_n10941, new_n10942, new_n10943, new_n10944, new_n10945, new_n10946,
    new_n10947, new_n10948, new_n10949, new_n10950, new_n10951, new_n10952,
    new_n10953, new_n10954, new_n10955, new_n10956, new_n10957, new_n10958,
    new_n10959, new_n10960, new_n10961, new_n10962, new_n10963, new_n10964,
    new_n10965, new_n10966, new_n10967, new_n10968, new_n10969, new_n10970,
    new_n10971, new_n10972, new_n10973, new_n10974, new_n10975, new_n10976,
    new_n10977, new_n10978, new_n10979, new_n10980, new_n10981, new_n10982,
    new_n10983, new_n10984, new_n10985, new_n10986, new_n10987, new_n10988,
    new_n10989, new_n10990, new_n10991, new_n10992, new_n10993, new_n10994,
    new_n10995, new_n10996, new_n10997, new_n10998, new_n10999, new_n11000,
    new_n11001, new_n11002, new_n11003, new_n11004, new_n11005, new_n11006,
    new_n11007, new_n11008, new_n11009, new_n11010, new_n11011, new_n11012,
    new_n11013, new_n11014, new_n11015, new_n11016, new_n11017, new_n11018,
    new_n11019, new_n11020, new_n11021, new_n11022, new_n11023, new_n11024,
    new_n11025, new_n11026, new_n11027, new_n11028, new_n11029,
    new_n11030_1, new_n11031, new_n11032, new_n11033, new_n11034,
    new_n11035, new_n11036, new_n11037, new_n11038, new_n11039, new_n11040,
    new_n11041, new_n11042, new_n11043, new_n11044, new_n11045, new_n11046,
    new_n11047, new_n11048, new_n11049, new_n11050, new_n11051, new_n11052,
    new_n11053, new_n11054, new_n11055, new_n11056, new_n11057_1,
    new_n11058_1, new_n11059, new_n11060, new_n11061_1, new_n11062,
    new_n11063, new_n11064, new_n11065, new_n11066, new_n11067, new_n11068,
    new_n11069, new_n11070, new_n11071, new_n11072, new_n11073, new_n11074,
    new_n11075, new_n11076, new_n11077_1, new_n11078, new_n11079,
    new_n11080, new_n11081, new_n11082, new_n11083, new_n11084, new_n11085,
    new_n11086, new_n11087, new_n11088, new_n11089, new_n11090, new_n11091,
    new_n11092, new_n11093, new_n11094, new_n11095, new_n11096, new_n11097,
    new_n11098, new_n11099, new_n11100, new_n11101, new_n11102, new_n11103,
    new_n11104, new_n11105, new_n11106, new_n11107, new_n11108,
    new_n11109_1, new_n11110, new_n11111_1, new_n11112, new_n11113,
    new_n11114, new_n11115, new_n11116, new_n11117, new_n11118, new_n11119,
    new_n11120, new_n11121, new_n11122, new_n11123, new_n11124, new_n11125,
    new_n11126, new_n11127, new_n11128, new_n11129, new_n11130, new_n11131,
    new_n11132, new_n11133, new_n11134, new_n11135, new_n11136, new_n11137,
    new_n11138, new_n11139, new_n11140_1, new_n11141, new_n11142,
    new_n11143, new_n11144, new_n11145, new_n11146, new_n11147_1,
    new_n11148, new_n11149, new_n11150, new_n11151, new_n11152, new_n11153,
    new_n11154, new_n11155, new_n11156, new_n11157, new_n11158, new_n11159,
    new_n11160, new_n11161, new_n11162, new_n11163, new_n11164, new_n11165,
    new_n11166, new_n11167, new_n11168, new_n11169, new_n11170, new_n11171,
    new_n11172, new_n11173, new_n11174, new_n11175, new_n11176, new_n11177,
    new_n11178, new_n11179, new_n11180_1, new_n11181, new_n11182,
    new_n11183, new_n11184, new_n11185, new_n11186, new_n11187, new_n11188,
    new_n11189, new_n11190, new_n11191, new_n11192, new_n11193, new_n11194,
    new_n11195, new_n11196, new_n11197, new_n11198, new_n11199, new_n11200,
    new_n11201, new_n11202, new_n11203, new_n11204, new_n11205, new_n11206,
    new_n11207, new_n11208, new_n11209, new_n11210, new_n11211, new_n11212,
    new_n11213, new_n11214, new_n11215, new_n11216, new_n11217, new_n11218,
    new_n11219, new_n11221, new_n11222_1, new_n11223, new_n11224,
    new_n11225, new_n11226, new_n11227, new_n11228, new_n11229, new_n11230,
    new_n11231, new_n11232, new_n11233, new_n11234, new_n11235,
    new_n11236_1, new_n11237, new_n11238, new_n11239, new_n11240,
    new_n11241, new_n11242, new_n11243, new_n11244, new_n11245, new_n11246,
    new_n11247, new_n11248, new_n11249, new_n11250, new_n11251,
    new_n11252_1, new_n11253, new_n11254, new_n11255, new_n11256,
    new_n11257, new_n11258, new_n11259, new_n11260, new_n11261, new_n11262,
    new_n11263, new_n11264_1, new_n11265, new_n11266, new_n11267,
    new_n11268, new_n11269, new_n11270, new_n11271, new_n11272, new_n11273,
    new_n11274, new_n11275, new_n11276, new_n11277, new_n11278, new_n11279,
    new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285,
    new_n11286, new_n11287, new_n11288, new_n11289, new_n11290, new_n11291,
    new_n11292, new_n11293, new_n11294, new_n11295, new_n11296, new_n11297,
    new_n11298, new_n11299, new_n11300, new_n11301, new_n11302, new_n11303,
    new_n11304, new_n11305, new_n11306, new_n11307, new_n11308, new_n11309,
    new_n11310, new_n11311, new_n11312, new_n11313, new_n11314, new_n11315,
    new_n11316, new_n11317, new_n11318, new_n11319, new_n11320, new_n11321,
    new_n11322, new_n11323, new_n11324_1, new_n11325, new_n11326,
    new_n11327, new_n11328, new_n11329, new_n11330, new_n11331, new_n11332,
    new_n11333, new_n11334, new_n11335, new_n11336, new_n11337, new_n11338,
    new_n11339, new_n11340, new_n11341, new_n11342, new_n11343, new_n11344,
    new_n11345, new_n11346, new_n11347, new_n11348, new_n11349,
    new_n11350_1, new_n11351, new_n11352, new_n11353, new_n11354,
    new_n11355, new_n11356, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375, new_n11376, new_n11377, new_n11378,
    new_n11379, new_n11380, new_n11381, new_n11382, new_n11383, new_n11384,
    new_n11385, new_n11386, new_n11387, new_n11388, new_n11389, new_n11390,
    new_n11391, new_n11392, new_n11393, new_n11394, new_n11395,
    new_n11396_1, new_n11397, new_n11398, new_n11399, new_n11400,
    new_n11401, new_n11402, new_n11403, new_n11404, new_n11405, new_n11406,
    new_n11407, new_n11408, new_n11409, new_n11410, new_n11411_1,
    new_n11412, new_n11413, new_n11414, new_n11415, new_n11416, new_n11417,
    new_n11418, new_n11419, new_n11420, new_n11421, new_n11422, new_n11423,
    new_n11424, new_n11425, new_n11426, new_n11427, new_n11428,
    new_n11429_1, new_n11430, new_n11431, new_n11432, new_n11433,
    new_n11434, new_n11435, new_n11436, new_n11437, new_n11438, new_n11439,
    new_n11440, new_n11441, new_n11442, new_n11443, new_n11444, new_n11445,
    new_n11446, new_n11447, new_n11448, new_n11449, new_n11450, new_n11451,
    new_n11452, new_n11453, new_n11454, new_n11455, new_n11456, new_n11457,
    new_n11458, new_n11459, new_n11460, new_n11461, new_n11462, new_n11463,
    new_n11464, new_n11465, new_n11466, new_n11467, new_n11468, new_n11469,
    new_n11470, new_n11471, new_n11472, new_n11473, new_n11474, new_n11475,
    new_n11476, new_n11477, new_n11478, new_n11479, new_n11480, new_n11481,
    new_n11482, new_n11483, new_n11484_1, new_n11485, new_n11486,
    new_n11487, new_n11488_1, new_n11489, new_n11490, new_n11491,
    new_n11492, new_n11493, new_n11494, new_n11495, new_n11496, new_n11497,
    new_n11498, new_n11499, new_n11500, new_n11501, new_n11502, new_n11503,
    new_n11504, new_n11505, new_n11506, new_n11507, new_n11508, new_n11509,
    new_n11510, new_n11511, new_n11512, new_n11513, new_n11514, new_n11515,
    new_n11516, new_n11517, new_n11518, new_n11519, new_n11520, new_n11521,
    new_n11522, new_n11523, new_n11524, new_n11525, new_n11526, new_n11527,
    new_n11528, new_n11529, new_n11530, new_n11531, new_n11532, new_n11533,
    new_n11534, new_n11535, new_n11536, new_n11537_1, new_n11538,
    new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544,
    new_n11545, new_n11546, new_n11547, new_n11548, new_n11549, new_n11550,
    new_n11551, new_n11552, new_n11553, new_n11554, new_n11555, new_n11556,
    new_n11557, new_n11558, new_n11559, new_n11560, new_n11561, new_n11562,
    new_n11563, new_n11564, new_n11565, new_n11566, new_n11567, new_n11568,
    new_n11569, new_n11570, new_n11571, new_n11572, new_n11573,
    new_n11574_1, new_n11575, new_n11576, new_n11577, new_n11578,
    new_n11579, new_n11580, new_n11581, new_n11582, new_n11583, new_n11584,
    new_n11585, new_n11586, new_n11587, new_n11588, new_n11589, new_n11590,
    new_n11591, new_n11592, new_n11593, new_n11594, new_n11595, new_n11596,
    new_n11597, new_n11598, new_n11599, new_n11600, new_n11601, new_n11602,
    new_n11603, new_n11604, new_n11605, new_n11606, new_n11607, new_n11608,
    new_n11609, new_n11610, new_n11611, new_n11612, new_n11613, new_n11614,
    new_n11615, new_n11616, new_n11617, new_n11618, new_n11619, new_n11620,
    new_n11621, new_n11622, new_n11623, new_n11624, new_n11625, new_n11626,
    new_n11627, new_n11628, new_n11629, new_n11630, new_n11631, new_n11632,
    new_n11633, new_n11634_1, new_n11635, new_n11636, new_n11637,
    new_n11638, new_n11639, new_n11640, new_n11641, new_n11642, new_n11643,
    new_n11644, new_n11645, new_n11646, new_n11647, new_n11648, new_n11649,
    new_n11650, new_n11651, new_n11652, new_n11653, new_n11654, new_n11655,
    new_n11656, new_n11657, new_n11658, new_n11659, new_n11660, new_n11661,
    new_n11662, new_n11663, new_n11664, new_n11665_1, new_n11666,
    new_n11667_1, new_n11668, new_n11669, new_n11670, new_n11671,
    new_n11672, new_n11673, new_n11674, new_n11675, new_n11676, new_n11677,
    new_n11678, new_n11679, new_n11680, new_n11681, new_n11682, new_n11683,
    new_n11684, new_n11685, new_n11686, new_n11687, new_n11688, new_n11689,
    new_n11690, new_n11691, new_n11692, new_n11693, new_n11694, new_n11695,
    new_n11696, new_n11697, new_n11698, new_n11699, new_n11700, new_n11702,
    new_n11703, new_n11704, new_n11705, new_n11706, new_n11707, new_n11708,
    new_n11709, new_n11710, new_n11711, new_n11712, new_n11713, new_n11714,
    new_n11715, new_n11716, new_n11717, new_n11718, new_n11719, new_n11720,
    new_n11721, new_n11722, new_n11723, new_n11724, new_n11725, new_n11726,
    new_n11727, new_n11728, new_n11729, new_n11730, new_n11731,
    new_n11732_1, new_n11733, new_n11734_1, new_n11735, new_n11736,
    new_n11737, new_n11738, new_n11739, new_n11740, new_n11741, new_n11742,
    new_n11743, new_n11744, new_n11745, new_n11746, new_n11747, new_n11748,
    new_n11749, new_n11750, new_n11751, new_n11752, new_n11753, new_n11754,
    new_n11755, new_n11756, new_n11757, new_n11758, new_n11759, new_n11760,
    new_n11761, new_n11762, new_n11763, new_n11764, new_n11765, new_n11766,
    new_n11767, new_n11768, new_n11769, new_n11770, new_n11771, new_n11772,
    new_n11773, new_n11774, new_n11775, new_n11776, new_n11777,
    new_n11778_1, new_n11779, new_n11780, new_n11781, new_n11782,
    new_n11783, new_n11784, new_n11785, new_n11786, new_n11787, new_n11788,
    new_n11789, new_n11790, new_n11791, new_n11792_1, new_n11793,
    new_n11794, new_n11795, new_n11796, new_n11797, new_n11798, new_n11799,
    new_n11800, new_n11801, new_n11802, new_n11803, new_n11804, new_n11805,
    new_n11806, new_n11807, new_n11808, new_n11809, new_n11810, new_n11811,
    new_n11812, new_n11813, new_n11814, new_n11815, new_n11816, new_n11817,
    new_n11818, new_n11819, new_n11820, new_n11821, new_n11822, new_n11823,
    new_n11824, new_n11825, new_n11826, new_n11827, new_n11828, new_n11829,
    new_n11830, new_n11831, new_n11832, new_n11833, new_n11834,
    new_n11835_1, new_n11836, new_n11837, new_n11838, new_n11839,
    new_n11840, new_n11841, new_n11842, new_n11843, new_n11844, new_n11845,
    new_n11846, new_n11847, new_n11848, new_n11849, new_n11850, new_n11851,
    new_n11852, new_n11853, new_n11854, new_n11855, new_n11856, new_n11857,
    new_n11858, new_n11859, new_n11860, new_n11861, new_n11862, new_n11863,
    new_n11864, new_n11865, new_n11866, new_n11867, new_n11868, new_n11869,
    new_n11870, new_n11871, new_n11872, new_n11873, new_n11874, new_n11875,
    new_n11876, new_n11877, new_n11878, new_n11879_1, new_n11880,
    new_n11881, new_n11882_1, new_n11883, new_n11884, new_n11885,
    new_n11886, new_n11887, new_n11888, new_n11889, new_n11890,
    new_n11891_1, new_n11892, new_n11893, new_n11894, new_n11895_1,
    new_n11896, new_n11897, new_n11898, new_n11899, new_n11900, new_n11901,
    new_n11902, new_n11903, new_n11904, new_n11905, new_n11906, new_n11907,
    new_n11908, new_n11909, new_n11910, new_n11911, new_n11912, new_n11913,
    new_n11914, new_n11915, new_n11916, new_n11917, new_n11918, new_n11919,
    new_n11920, new_n11921, new_n11922, new_n11923, new_n11924, new_n11925,
    new_n11926, new_n11927, new_n11928, new_n11929, new_n11930, new_n11931,
    new_n11932, new_n11933, new_n11934, new_n11935, new_n11936, new_n11937,
    new_n11938, new_n11939, new_n11940, new_n11941, new_n11942, new_n11943,
    new_n11944, new_n11945, new_n11946, new_n11947, new_n11948, new_n11949,
    new_n11950, new_n11951, new_n11952, new_n11953, new_n11954, new_n11955,
    new_n11956, new_n11957, new_n11958, new_n11959, new_n11960, new_n11961,
    new_n11962, new_n11963, new_n11964, new_n11965, new_n11966, new_n11967,
    new_n11968, new_n11969, new_n11970, new_n11971, new_n11972, new_n11973,
    new_n11974, new_n11975, new_n11976, new_n11977, new_n11978, new_n11979,
    new_n11980, new_n11981, new_n11982, new_n11983, new_n11984, new_n11985,
    new_n11986, new_n11987, new_n11988, new_n11989, new_n11990, new_n11991,
    new_n11992, new_n11993, new_n11994, new_n11995, new_n11996, new_n11997,
    new_n11998, new_n11999, new_n12000, new_n12001, new_n12002,
    new_n12003_1, new_n12004, new_n12005, new_n12006, new_n12007,
    new_n12008, new_n12009, new_n12010, new_n12011, new_n12012, new_n12013,
    new_n12014, new_n12015, new_n12016, new_n12017, new_n12018, new_n12019,
    new_n12020, new_n12021, new_n12022, new_n12023, new_n12024, new_n12025,
    new_n12026, new_n12027, new_n12028, new_n12029, new_n12030, new_n12031,
    new_n12032, new_n12033, new_n12034, new_n12035, new_n12036, new_n12037,
    new_n12038, new_n12039, new_n12040, new_n12041, new_n12042, new_n12043,
    new_n12044, new_n12045, new_n12046, new_n12047, new_n12048, new_n12049,
    new_n12050, new_n12051, new_n12052, new_n12053, new_n12054, new_n12055,
    new_n12056, new_n12057, new_n12058, new_n12059_1, new_n12060,
    new_n12061, new_n12062, new_n12063, new_n12064, new_n12065_1,
    new_n12066, new_n12067_1, new_n12068, new_n12069, new_n12070,
    new_n12071, new_n12072, new_n12073, new_n12074, new_n12075, new_n12076,
    new_n12077, new_n12078, new_n12079, new_n12080, new_n12081, new_n12082,
    new_n12083, new_n12084, new_n12085, new_n12086, new_n12087, new_n12088,
    new_n12089, new_n12090, new_n12091, new_n12092, new_n12093, new_n12094,
    new_n12095, new_n12096, new_n12097, new_n12098, new_n12099, new_n12100,
    new_n12101, new_n12102, new_n12103, new_n12104, new_n12105, new_n12106,
    new_n12107, new_n12108, new_n12109, new_n12110, new_n12111, new_n12112,
    new_n12113, new_n12114, new_n12115, new_n12116, new_n12117, new_n12118,
    new_n12119, new_n12120, new_n12121, new_n12122, new_n12123, new_n12124,
    new_n12125, new_n12126, new_n12127, new_n12128, new_n12129, new_n12130,
    new_n12131, new_n12132, new_n12133, new_n12134, new_n12135, new_n12136,
    new_n12137, new_n12138, new_n12139, new_n12140, new_n12141, new_n12142,
    new_n12143, new_n12144, new_n12145, new_n12146, new_n12147, new_n12148,
    new_n12149, new_n12150, new_n12151, new_n12152, new_n12153, new_n12154,
    new_n12155, new_n12156, new_n12157, new_n12158, new_n12159, new_n12160,
    new_n12161, new_n12162, new_n12163, new_n12164, new_n12165, new_n12166,
    new_n12167, new_n12168, new_n12169, new_n12170, new_n12171, new_n12172,
    new_n12173, new_n12174, new_n12175, new_n12176, new_n12177, new_n12178,
    new_n12179, new_n12180, new_n12181, new_n12182, new_n12183, new_n12184,
    new_n12185, new_n12186, new_n12187_1, new_n12188, new_n12189,
    new_n12190, new_n12191, new_n12192, new_n12193, new_n12194, new_n12195,
    new_n12196, new_n12197, new_n12198, new_n12199, new_n12200, new_n12201,
    new_n12202, new_n12203, new_n12204, new_n12205, new_n12206, new_n12207,
    new_n12208, new_n12209, new_n12210, new_n12211, new_n12212, new_n12213,
    new_n12214, new_n12215, new_n12216, new_n12217, new_n12218, new_n12219,
    new_n12220, new_n12221, new_n12222, new_n12223, new_n12224, new_n12225,
    new_n12226, new_n12227, new_n12228, new_n12229, new_n12230, new_n12231,
    new_n12232, new_n12233, new_n12234, new_n12235, new_n12236, new_n12237,
    new_n12238, new_n12239, new_n12240, new_n12241, new_n12242, new_n12243,
    new_n12244, new_n12245, new_n12246, new_n12247, new_n12248, new_n12249,
    new_n12250, new_n12251, new_n12252, new_n12253, new_n12254, new_n12255,
    new_n12256, new_n12257, new_n12258, new_n12259, new_n12260, new_n12261,
    new_n12262, new_n12263_1, new_n12264, new_n12265, new_n12266,
    new_n12267, new_n12268, new_n12269, new_n12270, new_n12271, new_n12272,
    new_n12273, new_n12274, new_n12275, new_n12276, new_n12277, new_n12278,
    new_n12279, new_n12280, new_n12281, new_n12282, new_n12283,
    new_n12284_1, new_n12285, new_n12286, new_n12287, new_n12288,
    new_n12289_1, new_n12290, new_n12291, new_n12292, new_n12293,
    new_n12294, new_n12295, new_n12296, new_n12297, new_n12298, new_n12299,
    new_n12300, new_n12301, new_n12302, new_n12303, new_n12304, new_n12305,
    new_n12306_1, new_n12307, new_n12308, new_n12309, new_n12310,
    new_n12311, new_n12312, new_n12313, new_n12314, new_n12315, new_n12316,
    new_n12317, new_n12318, new_n12319, new_n12320, new_n12321, new_n12322,
    new_n12323, new_n12324, new_n12325, new_n12326, new_n12327, new_n12328,
    new_n12329, new_n12330, new_n12331, new_n12332, new_n12333,
    new_n12334_1, new_n12335, new_n12336, new_n12337, new_n12338,
    new_n12339, new_n12340, new_n12341, new_n12342, new_n12343, new_n12344,
    new_n12345, new_n12346, new_n12347, new_n12348_1, new_n12349,
    new_n12350, new_n12351, new_n12352_1, new_n12353, new_n12354,
    new_n12355, new_n12356, new_n12357, new_n12358, new_n12359, new_n12360,
    new_n12361, new_n12362, new_n12363, new_n12364, new_n12365, new_n12366,
    new_n12367, new_n12368, new_n12369, new_n12370, new_n12371,
    new_n12372_1, new_n12373, new_n12374, new_n12375, new_n12376,
    new_n12377, new_n12378, new_n12379, new_n12380, new_n12381, new_n12382,
    new_n12383, new_n12384, new_n12385, new_n12386, new_n12387, new_n12388,
    new_n12389, new_n12390, new_n12391, new_n12392, new_n12393, new_n12394,
    new_n12395, new_n12396, new_n12397, new_n12398, new_n12399, new_n12400,
    new_n12401, new_n12402, new_n12403, new_n12404, new_n12405,
    new_n12406_1, new_n12407, new_n12408_1, new_n12409, new_n12410,
    new_n12411, new_n12412, new_n12413, new_n12414, new_n12415, new_n12416,
    new_n12417, new_n12418, new_n12419, new_n12420, new_n12421, new_n12422,
    new_n12423, new_n12424, new_n12425, new_n12426, new_n12427, new_n12428,
    new_n12429, new_n12430, new_n12431, new_n12432, new_n12433, new_n12434,
    new_n12435, new_n12436, new_n12437, new_n12438, new_n12439, new_n12440,
    new_n12441, new_n12442, new_n12443, new_n12444, new_n12445, new_n12446,
    new_n12447, new_n12448, new_n12449, new_n12450, new_n12451, new_n12452,
    new_n12453, new_n12454, new_n12455, new_n12456, new_n12457, new_n12458,
    new_n12459, new_n12460, new_n12461, new_n12462, new_n12463_1,
    new_n12464, new_n12465, new_n12466, new_n12467, new_n12468, new_n12469,
    new_n12470, new_n12472, new_n12473, new_n12474, new_n12476, new_n12477,
    new_n12478, new_n12479, new_n12480, new_n12481, new_n12482_1,
    new_n12483, new_n12484, new_n12485, new_n12486, new_n12487, new_n12488,
    new_n12489, new_n12490, new_n12491, new_n12492, new_n12493, new_n12494,
    new_n12495, new_n12496, new_n12497, new_n12498, new_n12499, new_n12500,
    new_n12501, new_n12502, new_n12503_1, new_n12504, new_n12505,
    new_n12506, new_n12507, new_n12508, new_n12509, new_n12510, new_n12511,
    new_n12512, new_n12513, new_n12514, new_n12515_1, new_n12516,
    new_n12517, new_n12518, new_n12519, new_n12520, new_n12521, new_n12522,
    new_n12523, new_n12524, new_n12525, new_n12526, new_n12527, new_n12528,
    new_n12529, new_n12530, new_n12531, new_n12532, new_n12533, new_n12534,
    new_n12535, new_n12536, new_n12537, new_n12538, new_n12539, new_n12540,
    new_n12541, new_n12542, new_n12543, new_n12544, new_n12545, new_n12546,
    new_n12547, new_n12548, new_n12549, new_n12550, new_n12551, new_n12552,
    new_n12553, new_n12554, new_n12555, new_n12556, new_n12557, new_n12558,
    new_n12559, new_n12560, new_n12561, new_n12562, new_n12563, new_n12564,
    new_n12565, new_n12566, new_n12567, new_n12568, new_n12569, new_n12570,
    new_n12571, new_n12572, new_n12573, new_n12574, new_n12575, new_n12576,
    new_n12577, new_n12578, new_n12579_1, new_n12580, new_n12581,
    new_n12582, new_n12583, new_n12584, new_n12585, new_n12586, new_n12587,
    new_n12588, new_n12589, new_n12590, new_n12591, new_n12592_1,
    new_n12593, new_n12594, new_n12595, new_n12596, new_n12597, new_n12598,
    new_n12599, new_n12600, new_n12601, new_n12602, new_n12603, new_n12604,
    new_n12605_1, new_n12606, new_n12607, new_n12608, new_n12609,
    new_n12610, new_n12611, new_n12612, new_n12613, new_n12614, new_n12615,
    new_n12616_1, new_n12617, new_n12618, new_n12619, new_n12620,
    new_n12621, new_n12622, new_n12623, new_n12624, new_n12625, new_n12626,
    new_n12627, new_n12628, new_n12629, new_n12630, new_n12631, new_n12632,
    new_n12633, new_n12634, new_n12635, new_n12636, new_n12637, new_n12638,
    new_n12639, new_n12640, new_n12641, new_n12642, new_n12643, new_n12644,
    new_n12645, new_n12646, new_n12647, new_n12648, new_n12649, new_n12650,
    new_n12651_1, new_n12652, new_n12653, new_n12654, new_n12655,
    new_n12656, new_n12657, new_n12658, new_n12659, new_n12660, new_n12661,
    new_n12662, new_n12663, new_n12664, new_n12665, new_n12666, new_n12667,
    new_n12668, new_n12669, new_n12670, new_n12671, new_n12672, new_n12673,
    new_n12674, new_n12675, new_n12676, new_n12677, new_n12678, new_n12679,
    new_n12680, new_n12681, new_n12682, new_n12683, new_n12684, new_n12685,
    new_n12686, new_n12687, new_n12688, new_n12689, new_n12690, new_n12691,
    new_n12692, new_n12693_1, new_n12694, new_n12695, new_n12696,
    new_n12697, new_n12698, new_n12699, new_n12700, new_n12701, new_n12702,
    new_n12703, new_n12704, new_n12705, new_n12706, new_n12707, new_n12708,
    new_n12709, new_n12710, new_n12711, new_n12712, new_n12713, new_n12714,
    new_n12715, new_n12716, new_n12717, new_n12718, new_n12719, new_n12720,
    new_n12721, new_n12722, new_n12723, new_n12724, new_n12725, new_n12726,
    new_n12727, new_n12728, new_n12729, new_n12730, new_n12731, new_n12732,
    new_n12733, new_n12734, new_n12735, new_n12736, new_n12737, new_n12738,
    new_n12739, new_n12740, new_n12741, new_n12742, new_n12743, new_n12744,
    new_n12745, new_n12746, new_n12747, new_n12748, new_n12749,
    new_n12750_1, new_n12751, new_n12752, new_n12753, new_n12754,
    new_n12755, new_n12756, new_n12757, new_n12758, new_n12759, new_n12760,
    new_n12761, new_n12762, new_n12763, new_n12764, new_n12765, new_n12766,
    new_n12767, new_n12768, new_n12769, new_n12770, new_n12771, new_n12772,
    new_n12773, new_n12774, new_n12775, new_n12776, new_n12777, new_n12778,
    new_n12779, new_n12780, new_n12781, new_n12782, new_n12783, new_n12784,
    new_n12785, new_n12786, new_n12787, new_n12788, new_n12789, new_n12790,
    new_n12791, new_n12792, new_n12793, new_n12794, new_n12795, new_n12796,
    new_n12797, new_n12798, new_n12799, new_n12800, new_n12801, new_n12802,
    new_n12803, new_n12804, new_n12805, new_n12806, new_n12807, new_n12808,
    new_n12809, new_n12810, new_n12811, new_n12812, new_n12813, new_n12814,
    new_n12815, new_n12816, new_n12817, new_n12818, new_n12819, new_n12821,
    new_n12822, new_n12823, new_n12825, new_n12826, new_n12827, new_n12829,
    new_n12831, new_n12832, new_n12833, new_n12835, new_n12836, new_n12837,
    new_n12839_1, new_n12840, new_n12841, new_n12843, new_n12844,
    new_n12845, new_n12847, new_n12848, new_n12849, new_n12851,
    new_n12853_1, new_n12854, new_n12855, new_n12857, new_n12858,
    new_n12859, new_n12861, new_n12862, new_n12863, new_n12865, new_n12866,
    new_n12867, new_n12869, new_n12870, new_n12871, new_n12873, new_n12874,
    new_n12875, new_n12877, new_n12879, new_n12880, new_n12881, new_n12883,
    new_n12884, new_n12885, new_n12887, new_n12888, new_n12889, new_n12890,
    new_n12891, new_n12892, new_n12893, new_n12894, new_n12895, new_n12896,
    new_n12897, new_n12898, new_n12899, new_n12900, new_n12901, new_n12902,
    new_n12903, new_n12904, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912_1, new_n12913,
    new_n12914, new_n12915, new_n12916, new_n12917, new_n12918, new_n12919,
    new_n12920, new_n12921, new_n12922, new_n12923, new_n12924, new_n12925,
    new_n12926, new_n12927, new_n12928, new_n12929, new_n12930, new_n12931,
    new_n12932, new_n12933, new_n12934, new_n12935, new_n12936, new_n12937,
    new_n12938, new_n12939, new_n12940, new_n12941, new_n12942, new_n12943,
    new_n12944, new_n12945, new_n12946, new_n12947, new_n12948, new_n12949,
    new_n12950, new_n12951, new_n12952, new_n12953, new_n12954, new_n12955,
    new_n12956, new_n12957, new_n12958, new_n12959, new_n12960, new_n12961,
    new_n12962, new_n12963, new_n12964, new_n12965_1, new_n12966,
    new_n12967, new_n12968_1, new_n12969, new_n12970, new_n12971,
    new_n12972, new_n12973, new_n12974, new_n12975, new_n12976, new_n12977,
    new_n12978, new_n12979, new_n12980, new_n12981, new_n12982, new_n12983,
    new_n12984, new_n12985, new_n12986, new_n12987, new_n12988, new_n12989,
    new_n12990, new_n12991, new_n12992, new_n12993, new_n12994, new_n12995,
    new_n12996, new_n12997, new_n12998, new_n12999, new_n13000, new_n13001,
    new_n13002_1, new_n13003, new_n13004, new_n13005, new_n13006,
    new_n13007, new_n13008, new_n13009, new_n13010, new_n13011, new_n13012,
    new_n13013, new_n13014, new_n13015, new_n13016, new_n13017, new_n13018,
    new_n13019, new_n13020, new_n13021, new_n13022, new_n13023, new_n13024,
    new_n13025, new_n13026, new_n13027, new_n13028, new_n13029, new_n13030,
    new_n13031, new_n13032, new_n13033, new_n13034, new_n13035_1,
    new_n13036, new_n13037, new_n13038, new_n13039, new_n13040, new_n13041,
    new_n13042, new_n13043, new_n13044, new_n13045, new_n13046, new_n13047,
    new_n13048, new_n13049, new_n13050, new_n13051, new_n13052, new_n13053,
    new_n13054, new_n13055, new_n13056, new_n13057, new_n13058_1,
    new_n13059, new_n13060_1, new_n13061, new_n13062, new_n13063,
    new_n13064, new_n13065, new_n13066, new_n13067, new_n13068, new_n13069,
    new_n13070, new_n13071, new_n13072, new_n13073, new_n13074, new_n13075,
    new_n13076, new_n13077, new_n13078, new_n13079, new_n13080, new_n13081,
    new_n13082, new_n13083, new_n13084, new_n13085, new_n13086, new_n13087,
    new_n13088, new_n13089, new_n13090, new_n13091, new_n13092, new_n13093,
    new_n13094, new_n13095, new_n13096, new_n13097, new_n13098, new_n13099,
    new_n13100, new_n13101, new_n13102, new_n13103, new_n13104, new_n13105,
    new_n13106, new_n13107, new_n13108, new_n13109, new_n13110, new_n13111,
    new_n13112, new_n13113, new_n13114, new_n13115, new_n13116, new_n13117,
    new_n13118, new_n13119, new_n13120, new_n13121, new_n13122, new_n13123,
    new_n13124, new_n13125, new_n13126, new_n13127, new_n13128, new_n13129,
    new_n13130, new_n13131, new_n13132, new_n13133, new_n13134, new_n13135,
    new_n13136, new_n13137, new_n13138, new_n13139, new_n13140, new_n13141,
    new_n13142, new_n13143, new_n13144, new_n13145, new_n13146, new_n13147,
    new_n13148, new_n13149, new_n13150, new_n13151, new_n13152, new_n13153,
    new_n13154, new_n13155, new_n13156, new_n13157, new_n13158, new_n13159,
    new_n13160, new_n13161, new_n13162, new_n13163, new_n13164, new_n13165,
    new_n13166, new_n13167, new_n13168, new_n13169, new_n13170, new_n13171,
    new_n13172, new_n13173, new_n13174, new_n13175, new_n13176, new_n13177,
    new_n13178, new_n13179, new_n13180, new_n13181, new_n13182, new_n13183,
    new_n13184, new_n13185, new_n13186, new_n13187, new_n13188, new_n13189,
    new_n13190, new_n13191, new_n13192, new_n13193, new_n13194, new_n13195,
    new_n13196, new_n13197, new_n13198, new_n13199, new_n13200,
    new_n13201_1, new_n13202, new_n13203, new_n13204, new_n13205,
    new_n13206, new_n13207, new_n13208, new_n13209, new_n13210, new_n13211,
    new_n13212, new_n13213, new_n13214, new_n13215, new_n13216, new_n13217,
    new_n13218, new_n13219, new_n13220, new_n13221, new_n13222, new_n13223,
    new_n13224, new_n13225, new_n13226, new_n13227, new_n13228, new_n13229,
    new_n13230, new_n13231, new_n13232, new_n13233, new_n13234, new_n13235,
    new_n13236, new_n13237, new_n13238, new_n13239, new_n13240, new_n13241,
    new_n13242, new_n13243, new_n13244, new_n13245, new_n13246, new_n13247,
    new_n13248, new_n13249, new_n13250, new_n13251, new_n13252, new_n13253,
    new_n13254, new_n13255, new_n13256, new_n13257, new_n13258, new_n13259,
    new_n13260, new_n13261, new_n13262, new_n13263, new_n13264, new_n13265,
    new_n13266, new_n13267, new_n13268, new_n13269, new_n13270, new_n13271,
    new_n13272, new_n13273, new_n13274, new_n13275, new_n13276, new_n13277,
    new_n13278, new_n13280, new_n13282, new_n13283, new_n13284, new_n13286,
    new_n13287, new_n13288, new_n13290, new_n13291, new_n13292, new_n13293,
    new_n13294, new_n13295, new_n13296, new_n13297, new_n13298, new_n13299,
    new_n13300, new_n13301, new_n13302, new_n13303, new_n13304, new_n13305,
    new_n13306, new_n13307, new_n13308, new_n13309, new_n13310, new_n13311,
    new_n13312, new_n13313, new_n13314, new_n13315, new_n13316, new_n13317,
    new_n13318, new_n13319, new_n13320, new_n13321, new_n13322, new_n13323,
    new_n13324, new_n13325, new_n13326, new_n13327, new_n13328, new_n13329,
    new_n13330, new_n13331, new_n13332, new_n13333, new_n13334, new_n13335,
    new_n13336, new_n13337, new_n13338, new_n13339, new_n13340, new_n13341,
    new_n13342, new_n13343, new_n13344, new_n13345, new_n13346, new_n13347,
    new_n13348, new_n13349, new_n13350, new_n13351, new_n13352, new_n13353,
    new_n13354, new_n13355, new_n13356, new_n13357, new_n13358, new_n13359,
    new_n13360, new_n13361, new_n13362, new_n13363, new_n13364, new_n13365,
    new_n13366, new_n13367, new_n13368, new_n13369, new_n13370, new_n13371,
    new_n13372, new_n13373, new_n13374, new_n13375, new_n13376, new_n13377,
    new_n13378, new_n13379, new_n13380, new_n13381, new_n13382, new_n13383,
    new_n13384, new_n13385, new_n13386, new_n13387, new_n13388, new_n13389,
    new_n13390, new_n13391, new_n13392, new_n13393, new_n13394, new_n13395,
    new_n13396, new_n13397, new_n13398, new_n13399, new_n13400, new_n13401,
    new_n13402, new_n13403, new_n13404, new_n13405, new_n13406, new_n13407,
    new_n13408, new_n13409, new_n13410, new_n13411, new_n13412, new_n13413,
    new_n13414, new_n13415, new_n13416, new_n13417, new_n13418, new_n13419,
    new_n13420, new_n13421, new_n13422, new_n13423, new_n13424, new_n13425,
    new_n13426, new_n13427, new_n13428, new_n13429, new_n13430, new_n13431,
    new_n13432, new_n13433, new_n13434, new_n13435, new_n13436, new_n13437,
    new_n13438, new_n13439, new_n13440, new_n13441, new_n13442, new_n13443,
    new_n13444, new_n13445, new_n13446, new_n13447, new_n13448, new_n13449,
    new_n13450, new_n13451, new_n13452, new_n13453, new_n13454, new_n13455,
    new_n13456, new_n13457, new_n13458, new_n13459, new_n13460, new_n13461,
    new_n13462, new_n13463, new_n13464, new_n13465, new_n13466, new_n13467,
    new_n13468, new_n13469, new_n13470, new_n13471, new_n13472, new_n13473,
    new_n13474, new_n13475, new_n13476, new_n13477, new_n13478, new_n13479,
    new_n13480, new_n13481, new_n13482, new_n13483, new_n13484, new_n13485,
    new_n13486, new_n13487, new_n13488, new_n13489, new_n13490, new_n13491,
    new_n13492, new_n13493, new_n13494, new_n13495, new_n13496, new_n13497,
    new_n13498, new_n13499, new_n13500, new_n13501, new_n13502, new_n13503,
    new_n13504, new_n13505, new_n13506, new_n13507, new_n13508, new_n13509,
    new_n13510, new_n13511, new_n13512, new_n13513, new_n13514, new_n13515,
    new_n13516, new_n13517, new_n13518, new_n13519, new_n13520, new_n13521,
    new_n13522, new_n13523, new_n13524, new_n13525, new_n13526, new_n13527,
    new_n13529, new_n13530, new_n13531, new_n13533, new_n13534, new_n13535,
    new_n13536, new_n13537, new_n13538, new_n13539, new_n13540, new_n13541,
    new_n13542, new_n13543, new_n13544, new_n13545, new_n13546, new_n13547,
    new_n13548, new_n13549, new_n13550, new_n13551, new_n13552, new_n13553,
    new_n13554, new_n13555, new_n13556, new_n13557, new_n13558, new_n13559,
    new_n13560, new_n13561, new_n13562, new_n13563, new_n13564, new_n13565,
    new_n13566, new_n13567, new_n13568, new_n13569, new_n13570, new_n13571,
    new_n13572, new_n13573, new_n13574, new_n13575, new_n13576, new_n13577,
    new_n13578, new_n13579, new_n13580, new_n13581, new_n13582, new_n13583,
    new_n13584, new_n13585, new_n13586, new_n13587, new_n13588, new_n13589,
    new_n13590, new_n13591, new_n13592, new_n13593, new_n13594, new_n13595,
    new_n13596, new_n13597, new_n13598, new_n13599, new_n13600, new_n13601,
    new_n13602, new_n13603, new_n13604, new_n13605, new_n13606, new_n13607,
    new_n13608, new_n13609, new_n13610, new_n13611, new_n13612, new_n13613,
    new_n13614, new_n13615, new_n13616, new_n13617, new_n13618, new_n13619,
    new_n13620, new_n13621, new_n13622, new_n13623, new_n13624, new_n13625,
    new_n13626, new_n13627, new_n13628, new_n13629, new_n13630, new_n13631,
    new_n13632, new_n13633, new_n13634, new_n13635, new_n13636, new_n13637,
    new_n13638, new_n13639, new_n13640, new_n13641, new_n13642, new_n13643,
    new_n13644, new_n13645, new_n13646, new_n13647, new_n13648, new_n13649,
    new_n13650, new_n13651, new_n13652, new_n13653, new_n13654, new_n13655,
    new_n13656, new_n13657, new_n13658, new_n13659, new_n13660, new_n13661,
    new_n13662, new_n13663, new_n13664, new_n13665, new_n13666, new_n13667,
    new_n13668, new_n13669, new_n13670, new_n13671, new_n13672, new_n13673,
    new_n13674, new_n13675, new_n13676, new_n13677, new_n13678, new_n13679,
    new_n13680, new_n13681, new_n13682, new_n13683, new_n13684, new_n13685,
    new_n13686, new_n13687, new_n13688, new_n13689, new_n13690, new_n13691,
    new_n13692, new_n13693, new_n13694, new_n13695, new_n13696, new_n13697,
    new_n13698, new_n13699, new_n13700, new_n13701, new_n13702, new_n13703,
    new_n13704, new_n13705, new_n13706, new_n13707, new_n13708, new_n13709,
    new_n13710, new_n13711, new_n13712, new_n13713, new_n13714, new_n13715,
    new_n13716, new_n13717, new_n13718, new_n13719, new_n13720, new_n13721,
    new_n13722, new_n13723, new_n13724, new_n13725, new_n13726, new_n13727,
    new_n13728, new_n13729, new_n13730, new_n13731, new_n13732, new_n13733,
    new_n13734, new_n13735, new_n13736, new_n13737, new_n13738, new_n13739,
    new_n13740, new_n13741, new_n13742, new_n13743, new_n13744, new_n13745,
    new_n13746, new_n13747, new_n13748, new_n13749, new_n13750, new_n13751,
    new_n13752, new_n13753, new_n13754, new_n13755, new_n13756, new_n13757,
    new_n13758, new_n13759, new_n13760, new_n13761, new_n13762, new_n13763,
    new_n13764, new_n13765, new_n13766, new_n13767, new_n13768, new_n13769,
    new_n13770, new_n13771, new_n13772, new_n13773, new_n13774, new_n13775,
    new_n13776, new_n13777, new_n13778, new_n13779, new_n13780, new_n13781,
    new_n13782, new_n13783, new_n13784, new_n13785, new_n13786, new_n13787,
    new_n13788, new_n13789, new_n13790, new_n13791, new_n13792, new_n13793,
    new_n13794, new_n13795, new_n13796, new_n13797, new_n13798, new_n13799,
    new_n13800, new_n13801, new_n13802, new_n13803, new_n13804, new_n13805,
    new_n13806, new_n13807, new_n13808, new_n13809, new_n13810, new_n13811,
    new_n13812, new_n13813, new_n13814, new_n13815, new_n13816, new_n13817,
    new_n13818, new_n13819, new_n13820, new_n13821, new_n13822, new_n13823,
    new_n13824, new_n13825, new_n13826, new_n13827, new_n13828, new_n13829,
    new_n13830, new_n13831, new_n13832, new_n13833, new_n13834, new_n13835,
    new_n13836, new_n13837, new_n13838, new_n13839, new_n13840, new_n13841,
    new_n13842, new_n13843, new_n13844, new_n13845, new_n13846, new_n13847,
    new_n13848, new_n13849, new_n13850, new_n13851, new_n13852, new_n13853,
    new_n13854, new_n13855, new_n13856, new_n13857, new_n13858, new_n13859,
    new_n13860, new_n13861, new_n13862, new_n13863, new_n13864, new_n13865,
    new_n13866, new_n13867, new_n13868, new_n13869, new_n13870, new_n13871,
    new_n13872, new_n13873, new_n13874, new_n13875, new_n13876, new_n13877,
    new_n13878, new_n13879, new_n13880, new_n13881, new_n13882, new_n13883,
    new_n13884, new_n13885, new_n13886, new_n13887, new_n13888, new_n13889,
    new_n13890, new_n13891, new_n13892, new_n13893, new_n13894, new_n13895,
    new_n13896, new_n13897, new_n13898, new_n13899, new_n13900, new_n13901,
    new_n13902, new_n13903, new_n13904, new_n13905, new_n13906, new_n13907,
    new_n13908, new_n13909, new_n13910, new_n13911, new_n13912, new_n13913,
    new_n13914, new_n13915, new_n13916, new_n13917, new_n13918, new_n13919,
    new_n13920, new_n13921, new_n13922, new_n13923, new_n13924, new_n13925,
    new_n13926, new_n13927, new_n13928, new_n13929, new_n13930, new_n13931,
    new_n13932, new_n13933, new_n13934, new_n13935, new_n13936, new_n13937,
    new_n13938, new_n13939, new_n13940, new_n13941, new_n13942, new_n13943,
    new_n13944, new_n13945, new_n13946, new_n13947, new_n13948, new_n13949,
    new_n13950, new_n13951, new_n13952, new_n13953, new_n13954, new_n13955,
    new_n13956, new_n13957, new_n13958, new_n13959, new_n13960, new_n13961,
    new_n13962, new_n13963, new_n13964, new_n13965, new_n13966, new_n13967,
    new_n13968, new_n13969, new_n13970, new_n13971, new_n13972, new_n13973,
    new_n13974, new_n13975, new_n13976, new_n13977, new_n13978, new_n13979,
    new_n13980, new_n13981, new_n13982, new_n13983, new_n13984, new_n13985,
    new_n13986, new_n13987, new_n13988, new_n13989, new_n13990, new_n13991,
    new_n13992, new_n13993, new_n13994, new_n13995, new_n13996, new_n13997,
    new_n13998, new_n13999, new_n14000, new_n14001, new_n14002, new_n14003,
    new_n14004, new_n14005, new_n14006, new_n14007, new_n14008, new_n14009,
    new_n14010, new_n14011, new_n14012, new_n14013, new_n14014, new_n14015,
    new_n14016, new_n14017, new_n14018, new_n14019, new_n14020, new_n14021,
    new_n14022, new_n14023, new_n14024, new_n14025, new_n14026, new_n14027,
    new_n14028, new_n14029, new_n14030, new_n14031, new_n14032, new_n14033,
    new_n14034, new_n14035, new_n14036, new_n14037, new_n14038, new_n14039,
    new_n14040, new_n14041, new_n14042, new_n14043, new_n14044, new_n14045,
    new_n14046, new_n14047, new_n14048, new_n14049, new_n14050, new_n14051,
    new_n14052, new_n14053, new_n14054, new_n14055, new_n14056, new_n14057,
    new_n14058, new_n14059, new_n14060, new_n14061, new_n14063, new_n14065,
    new_n14066, new_n14067, new_n14069, new_n14070, new_n14071, new_n14073,
    new_n14074, new_n14075, new_n14077, new_n14078, new_n14079, new_n14081,
    new_n14082, new_n14083, new_n14084, new_n14085, new_n14086, new_n14087,
    new_n14088, new_n14089, new_n14090, new_n14091, new_n14092, new_n14093,
    new_n14094, new_n14095, new_n14096, new_n14097, new_n14098, new_n14099,
    new_n14100, new_n14101, new_n14102, new_n14103, new_n14104, new_n14105,
    new_n14106, new_n14107, new_n14108, new_n14109, new_n14110, new_n14111,
    new_n14112, new_n14113, new_n14114, new_n14115, new_n14116, new_n14117,
    new_n14118, new_n14119, new_n14120, new_n14121, new_n14122, new_n14123,
    new_n14124, new_n14125, new_n14126, new_n14127, new_n14128, new_n14129,
    new_n14130, new_n14131, new_n14132, new_n14133, new_n14134, new_n14135,
    new_n14136, new_n14137, new_n14138, new_n14139, new_n14140, new_n14141,
    new_n14142, new_n14143, new_n14144, new_n14145, new_n14146, new_n14147,
    new_n14148, new_n14149, new_n14150, new_n14151, new_n14152, new_n14153,
    new_n14154, new_n14155, new_n14156, new_n14157, new_n14158, new_n14159,
    new_n14160, new_n14161, new_n14162, new_n14163, new_n14164, new_n14165,
    new_n14166, new_n14167, new_n14168, new_n14169, new_n14170, new_n14171,
    new_n14172, new_n14173, new_n14174, new_n14175, new_n14176, new_n14177,
    new_n14178, new_n14179, new_n14180, new_n14181, new_n14182, new_n14183,
    new_n14184, new_n14185, new_n14186, new_n14187, new_n14188, new_n14189,
    new_n14190, new_n14191, new_n14192, new_n14193, new_n14194, new_n14195,
    new_n14196, new_n14197, new_n14198, new_n14199, new_n14200, new_n14201,
    new_n14202, new_n14203, new_n14204, new_n14205, new_n14206, new_n14207,
    new_n14208, new_n14209, new_n14210, new_n14211, new_n14212, new_n14213,
    new_n14214, new_n14215, new_n14216, new_n14217, new_n14218, new_n14219,
    new_n14220, new_n14221, new_n14222, new_n14223, new_n14224, new_n14225,
    new_n14226, new_n14227, new_n14228, new_n14229, new_n14230, new_n14231,
    new_n14232, new_n14233, new_n14234, new_n14235, new_n14236, new_n14237,
    new_n14238, new_n14239, new_n14240, new_n14241, new_n14242, new_n14243,
    new_n14244, new_n14245, new_n14246, new_n14247, new_n14248, new_n14249,
    new_n14250, new_n14251, new_n14252, new_n14253, new_n14254, new_n14255,
    new_n14256, new_n14257, new_n14258, new_n14259, new_n14260, new_n14261,
    new_n14262, new_n14263, new_n14264, new_n14265, new_n14266, new_n14267,
    new_n14268, new_n14269, new_n14270, new_n14271, new_n14272, new_n14273,
    new_n14274, new_n14275, new_n14276, new_n14277, new_n14278, new_n14279,
    new_n14280, new_n14281, new_n14282, new_n14283, new_n14284, new_n14285,
    new_n14286, new_n14287, new_n14288, new_n14289, new_n14290, new_n14291,
    new_n14292, new_n14293, new_n14294, new_n14295, new_n14296, new_n14297,
    new_n14298, new_n14299, new_n14300, new_n14301, new_n14302, new_n14303,
    new_n14304, new_n14305, new_n14306, new_n14307, new_n14308, new_n14309,
    new_n14310, new_n14311, new_n14312, new_n14313, new_n14314, new_n14316,
    new_n14317, new_n14318, new_n14320, new_n14321, new_n14322, new_n14324,
    new_n14325, new_n14326, new_n14327, new_n14328, new_n14329, new_n14330,
    new_n14331, new_n14332, new_n14333, new_n14334, new_n14335, new_n14336,
    new_n14337, new_n14338, new_n14339, new_n14340, new_n14341, new_n14342,
    new_n14343, new_n14344, new_n14345, new_n14346, new_n14347, new_n14348,
    new_n14349, new_n14350, new_n14351, new_n14352, new_n14353, new_n14354,
    new_n14355, new_n14356, new_n14357, new_n14358, new_n14359, new_n14360,
    new_n14361, new_n14362, new_n14363, new_n14364, new_n14365, new_n14366,
    new_n14367, new_n14368, new_n14369, new_n14370, new_n14371, new_n14372,
    new_n14373, new_n14374, new_n14375, new_n14376, new_n14377, new_n14378,
    new_n14379, new_n14380, new_n14381, new_n14382, new_n14383, new_n14384,
    new_n14385, new_n14386, new_n14387, new_n14388, new_n14389, new_n14390,
    new_n14391, new_n14392, new_n14393, new_n14394, new_n14395, new_n14396,
    new_n14397, new_n14398, new_n14399, new_n14400, new_n14401, new_n14402,
    new_n14403, new_n14404, new_n14405, new_n14406, new_n14407, new_n14408,
    new_n14409, new_n14410, new_n14411, new_n14412, new_n14413, new_n14414,
    new_n14415, new_n14416, new_n14417, new_n14418, new_n14419, new_n14420,
    new_n14421, new_n14422, new_n14423, new_n14424, new_n14425, new_n14426,
    new_n14427, new_n14428, new_n14429, new_n14430, new_n14431, new_n14432,
    new_n14433, new_n14434, new_n14435, new_n14436, new_n14437, new_n14438,
    new_n14439, new_n14440, new_n14441, new_n14442, new_n14443, new_n14444,
    new_n14445, new_n14446, new_n14447, new_n14448, new_n14449, new_n14450,
    new_n14451, new_n14452, new_n14453, new_n14454, new_n14455, new_n14456,
    new_n14457, new_n14458, new_n14459, new_n14460, new_n14461, new_n14462,
    new_n14463, new_n14464, new_n14465, new_n14466, new_n14467, new_n14468,
    new_n14469, new_n14470, new_n14471, new_n14472, new_n14473, new_n14474,
    new_n14475, new_n14476, new_n14477, new_n14478, new_n14479, new_n14480,
    new_n14481, new_n14482, new_n14483, new_n14484, new_n14485, new_n14486,
    new_n14487, new_n14488, new_n14489, new_n14490, new_n14491, new_n14492,
    new_n14493, new_n14494, new_n14495, new_n14496, new_n14497, new_n14498,
    new_n14499, new_n14500, new_n14501, new_n14502, new_n14503, new_n14504,
    new_n14505, new_n14506, new_n14507, new_n14508, new_n14509, new_n14510,
    new_n14511, new_n14512, new_n14513, new_n14514, new_n14515, new_n14516,
    new_n14517, new_n14518, new_n14519, new_n14520, new_n14521, new_n14522,
    new_n14523, new_n14524, new_n14525, new_n14526, new_n14527, new_n14528,
    new_n14529, new_n14530, new_n14531, new_n14532, new_n14533, new_n14534,
    new_n14535, new_n14536, new_n14538, new_n14539, new_n14540, new_n14542,
    new_n14543, new_n14544, new_n14546, new_n14548, new_n14549, new_n14550,
    new_n14552, new_n14553, new_n14554, new_n14556, new_n14557, new_n14558,
    new_n14560, new_n14561, new_n14562, new_n14564, new_n14565, new_n14566,
    new_n14568, new_n14569, new_n14570, new_n14572, new_n14573, new_n14574,
    new_n14576, new_n14577, new_n14578, new_n14579, new_n14580, new_n14581,
    new_n14582, new_n14583, new_n14584, new_n14585, new_n14586, new_n14587,
    new_n14588, new_n14589, new_n14590, new_n14591, new_n14592, new_n14593,
    new_n14594, new_n14595, new_n14596, new_n14597, new_n14598, new_n14599,
    new_n14600, new_n14601, new_n14602, new_n14603, new_n14604, new_n14605,
    new_n14606, new_n14607, new_n14608, new_n14609, new_n14610, new_n14611,
    new_n14612, new_n14613, new_n14614, new_n14615, new_n14616, new_n14617,
    new_n14618, new_n14619, new_n14620, new_n14621, new_n14622, new_n14623,
    new_n14624, new_n14625, new_n14626, new_n14627, new_n14628, new_n14629,
    new_n14630, new_n14631, new_n14632, new_n14633, new_n14634, new_n14635,
    new_n14636, new_n14637, new_n14638, new_n14639, new_n14640, new_n14641,
    new_n14642, new_n14643, new_n14644, new_n14645, new_n14646, new_n14647,
    new_n14648, new_n14649, new_n14650, new_n14651, new_n14652, new_n14653,
    new_n14654, new_n14655, new_n14656, new_n14657, new_n14658, new_n14659,
    new_n14660, new_n14661, new_n14662, new_n14663, new_n14664, new_n14665,
    new_n14666, new_n14667, new_n14668, new_n14669, new_n14670, new_n14671,
    new_n14672, new_n14673, new_n14674, new_n14675, new_n14676, new_n14677,
    new_n14678, new_n14679, new_n14680, new_n14681, new_n14682, new_n14683,
    new_n14684, new_n14685, new_n14686, new_n14687, new_n14688, new_n14689,
    new_n14690, new_n14691, new_n14692, new_n14693, new_n14694, new_n14695,
    new_n14696, new_n14697, new_n14698, new_n14699, new_n14700, new_n14701,
    new_n14702, new_n14703, new_n14704, new_n14705, new_n14706, new_n14707,
    new_n14708, new_n14709, new_n14710, new_n14711, new_n14712, new_n14713,
    new_n14714, new_n14715, new_n14716, new_n14717, new_n14718, new_n14719,
    new_n14720, new_n14721, new_n14722, new_n14723, new_n14724, new_n14725,
    new_n14726, new_n14727, new_n14728, new_n14729, new_n14730, new_n14731,
    new_n14732, new_n14733, new_n14734, new_n14735, new_n14736, new_n14737,
    new_n14738, new_n14739, new_n14740, new_n14741, new_n14742, new_n14743,
    new_n14744, new_n14745, new_n14746, new_n14747, new_n14748, new_n14749,
    new_n14750, new_n14751, new_n14752, new_n14753, new_n14754, new_n14755,
    new_n14756, new_n14757, new_n14758, new_n14759, new_n14760, new_n14761,
    new_n14762, new_n14763, new_n14764, new_n14765, new_n14766, new_n14767,
    new_n14768, new_n14769, new_n14770, new_n14771, new_n14772, new_n14773,
    new_n14774, new_n14775, new_n14776, new_n14777, new_n14778, new_n14779,
    new_n14780, new_n14781, new_n14782, new_n14783, new_n14784, new_n14785,
    new_n14786, new_n14787, new_n14788, new_n14789, new_n14790, new_n14791,
    new_n14792, new_n14793, new_n14794, new_n14795, new_n14796, new_n14797,
    new_n14798, new_n14799, new_n14800, new_n14801, new_n14802, new_n14803,
    new_n14804, new_n14805, new_n14806, new_n14807, new_n14808, new_n14809,
    new_n14810, new_n14811, new_n14812, new_n14813, new_n14814, new_n14815,
    new_n14816, new_n14817, new_n14818, new_n14819, new_n14820, new_n14821,
    new_n14822, new_n14823, new_n14824, new_n14825, new_n14826, new_n14827,
    new_n14828, new_n14829, new_n14830, new_n14831, new_n14832, new_n14833,
    new_n14834, new_n14835, new_n14836, new_n14837, new_n14838, new_n14839,
    new_n14840, new_n14841, new_n14842, new_n14843, new_n14844, new_n14845,
    new_n14846, new_n14847, new_n14848, new_n14849, new_n14850, new_n14851,
    new_n14852, new_n14853, new_n14854, new_n14855, new_n14856, new_n14857,
    new_n14858, new_n14859, new_n14860, new_n14861, new_n14862, new_n14863,
    new_n14864, new_n14865, new_n14866, new_n14867, new_n14868, new_n14869,
    new_n14870, new_n14871, new_n14872, new_n14873, new_n14874, new_n14875,
    new_n14876, new_n14877, new_n14878, new_n14879, new_n14880, new_n14881,
    new_n14882, new_n14883, new_n14884, new_n14885, new_n14886, new_n14887,
    new_n14888, new_n14889, new_n14890, new_n14891, new_n14892, new_n14893,
    new_n14894, new_n14895, new_n14896, new_n14897, new_n14898, new_n14899,
    new_n14900, new_n14901, new_n14902, new_n14903, new_n14904, new_n14905,
    new_n14906, new_n14907, new_n14908, new_n14909, new_n14910, new_n14911,
    new_n14912, new_n14913, new_n14914, new_n14915, new_n14916, new_n14917,
    new_n14918, new_n14919, new_n14920, new_n14921, new_n14922, new_n14923,
    new_n14924, new_n14925, new_n14926, new_n14927, new_n14928, new_n14929,
    new_n14930, new_n14931, new_n14932, new_n14933, new_n14934, new_n14935,
    new_n14936, new_n14937, new_n14938, new_n14939, new_n14940, new_n14941,
    new_n14942, new_n14943, new_n14944, new_n14945, new_n14946, new_n14947,
    new_n14948, new_n14949, new_n14950, new_n14951, new_n14952, new_n14953,
    new_n14954, new_n14955, new_n14956, new_n14957, new_n14958, new_n14959,
    new_n14960, new_n14961, new_n14962, new_n14963, new_n14964, new_n14965,
    new_n14966, new_n14967, new_n14969, new_n14970, new_n14971, new_n14973,
    new_n14974, new_n14975, new_n14977, new_n14978, new_n14979, new_n14981,
    new_n14982, new_n14983, new_n14985, new_n14986, new_n14987, new_n14989,
    new_n14990, new_n14991, new_n14993, new_n14995, new_n14996, new_n14997,
    new_n14998, new_n14999, new_n15000, new_n15001, new_n15002, new_n15003,
    new_n15004, new_n15005, new_n15006, new_n15007, new_n15008, new_n15009,
    new_n15010, new_n15011, new_n15012, new_n15013, new_n15014, new_n15015,
    new_n15016, new_n15017, new_n15018, new_n15019, new_n15020, new_n15021,
    new_n15022, new_n15023, new_n15024, new_n15025, new_n15026, new_n15027,
    new_n15028, new_n15029, new_n15030, new_n15031, new_n15032, new_n15033,
    new_n15034, new_n15035, new_n15036, new_n15037, new_n15038, new_n15039,
    new_n15040, new_n15041, new_n15042, new_n15043, new_n15044, new_n15045,
    new_n15046, new_n15047, new_n15048, new_n15049, new_n15050, new_n15051,
    new_n15052, new_n15053, new_n15054, new_n15055, new_n15056, new_n15057,
    new_n15058, new_n15059, new_n15060, new_n15061, new_n15062, new_n15063,
    new_n15064, new_n15065, new_n15066, new_n15067, new_n15068, new_n15069,
    new_n15070, new_n15071, new_n15072, new_n15073, new_n15074, new_n15075,
    new_n15076, new_n15077, new_n15078, new_n15079, new_n15080, new_n15081,
    new_n15082, new_n15083, new_n15084, new_n15085, new_n15086, new_n15087,
    new_n15088, new_n15089, new_n15090, new_n15091, new_n15092, new_n15093,
    new_n15094, new_n15095, new_n15096, new_n15097, new_n15098, new_n15099,
    new_n15100, new_n15101, new_n15102, new_n15103, new_n15104, new_n15105,
    new_n15106, new_n15107, new_n15108, new_n15109, new_n15110, new_n15111,
    new_n15112, new_n15113, new_n15114, new_n15115, new_n15116, new_n15117,
    new_n15118, new_n15119, new_n15120, new_n15121, new_n15122, new_n15123,
    new_n15124, new_n15125, new_n15126, new_n15127, new_n15128, new_n15129,
    new_n15130, new_n15131, new_n15132, new_n15133, new_n15134, new_n15135,
    new_n15136, new_n15137, new_n15138, new_n15139, new_n15140, new_n15141,
    new_n15142, new_n15143, new_n15144, new_n15145, new_n15146, new_n15147,
    new_n15148, new_n15149, new_n15150, new_n15151, new_n15152, new_n15153,
    new_n15154, new_n15155, new_n15156, new_n15157, new_n15158, new_n15159,
    new_n15160, new_n15161, new_n15162, new_n15163, new_n15164, new_n15165,
    new_n15166, new_n15167, new_n15168, new_n15169, new_n15170, new_n15171,
    new_n15172, new_n15173, new_n15174, new_n15175, new_n15176, new_n15177,
    new_n15178, new_n15179, new_n15180, new_n15181, new_n15182, new_n15183,
    new_n15184, new_n15185, new_n15186, new_n15187, new_n15188, new_n15189,
    new_n15190, new_n15191, new_n15192, new_n15193, new_n15194, new_n15195,
    new_n15196, new_n15197, new_n15198, new_n15199, new_n15200, new_n15201,
    new_n15202, new_n15203, new_n15204, new_n15205, new_n15206, new_n15207,
    new_n15208, new_n15209, new_n15210, new_n15211, new_n15212, new_n15213,
    new_n15214, new_n15215, new_n15216, new_n15217, new_n15218, new_n15219,
    new_n15220, new_n15221, new_n15222, new_n15223, new_n15224, new_n15225,
    new_n15226, new_n15227, new_n15228, new_n15229, new_n15230, new_n15231,
    new_n15232, new_n15233, new_n15234, new_n15235, new_n15236;
  assign new_n362 = n7772 & n9531;
  assign new_n363 = n7529 & n12853;
  assign new_n364 = new_n362 & new_n363;
  assign new_n365 = n7715 & n12853;
  assign new_n366 = n7529 & n9531;
  assign new_n367 = n7772 & n11891;
  assign new_n368 = ~new_n366 & ~new_n367;
  assign new_n369 = new_n366 & new_n367;
  assign new_n370_1 = ~new_n368 & ~new_n369;
  assign new_n371 = new_n365 & ~new_n370_1;
  assign new_n372 = ~new_n365 & new_n370_1;
  assign new_n373 = ~new_n371 & ~new_n372;
  assign new_n374 = ~new_n364 & new_n373;
  assign new_n375 = new_n364 & ~new_n373;
  assign new_n376 = ~new_n374 & ~new_n375;
  assign new_n377 = ~new_n362 & ~new_n363;
  assign new_n378 = ~new_n364 & ~new_n377;
  assign new_n379 = n510 & n8466;
  assign new_n380 = n834 & n3178;
  assign new_n381 = new_n379 & new_n380;
  assign new_n382 = ~new_n379 & ~new_n380;
  assign new_n383 = ~new_n381 & ~new_n382;
  assign new_n384 = n854 & n9216;
  assign new_n385 = new_n383 & new_n384;
  assign new_n386 = n12348 & new_n384;
  assign new_n387 = n854 & n12348;
  assign new_n388 = ~new_n384 & ~new_n387;
  assign new_n389_1 = ~new_n386 & ~new_n388;
  assign new_n390 = ~new_n385 & ~new_n389_1;
  assign new_n391 = ~n12348 & new_n385;
  assign new_n392 = ~new_n390 & ~new_n391;
  assign new_n393 = n3178 & n8716;
  assign new_n394 = n834 & n12592;
  assign new_n395 = ~new_n393 & ~new_n394;
  assign new_n396_1 = new_n393 & new_n394;
  assign new_n397 = ~new_n395 & ~new_n396_1;
  assign new_n398 = n8290 & n8466;
  assign new_n399 = n510 & n5031;
  assign new_n400 = ~new_n398 & ~new_n399;
  assign new_n401_1 = new_n398 & new_n399;
  assign new_n402 = ~new_n400 & ~new_n401_1;
  assign new_n403 = ~new_n381 & ~new_n402;
  assign new_n404 = new_n381 & new_n402;
  assign new_n405 = ~new_n403 & ~new_n404;
  assign new_n406 = ~new_n397 & new_n405;
  assign new_n407 = new_n397 & ~new_n405;
  assign new_n408 = ~new_n406 & ~new_n407;
  assign new_n409 = ~new_n392 & new_n408;
  assign new_n410 = new_n392 & ~new_n408;
  assign new_n411_1 = ~new_n409 & ~new_n410;
  assign new_n412 = ~new_n378 & ~new_n411_1;
  assign new_n413 = new_n378 & new_n411_1;
  assign new_n414 = n7772 & n12853;
  assign new_n415 = ~new_n383 & ~new_n384;
  assign new_n416 = ~new_n385 & ~new_n415;
  assign new_n417 = new_n414 & new_n416;
  assign new_n418 = ~new_n413 & ~new_n417;
  assign new_n419 = ~new_n412 & ~new_n418;
  assign new_n420 = ~new_n376 & ~new_n419;
  assign new_n421 = new_n376 & new_n419;
  assign new_n422 = ~new_n420 & ~new_n421;
  assign new_n423 = n2068 & ~new_n388;
  assign new_n424 = n854 & n2068;
  assign new_n425 = new_n388 & ~new_n424;
  assign new_n426 = ~new_n423 & ~new_n425;
  assign new_n427 = ~new_n391 & new_n408;
  assign new_n428 = ~new_n390 & ~new_n427;
  assign new_n429 = ~new_n426 & ~new_n428;
  assign new_n430 = new_n426 & new_n428;
  assign new_n431 = ~new_n429 & ~new_n430;
  assign new_n432 = n9 & n510;
  assign new_n433 = n5031 & n8290;
  assign new_n434 = n8466 & n9591;
  assign new_n435 = ~new_n433 & ~new_n434;
  assign new_n436 = new_n433 & new_n434;
  assign new_n437 = ~new_n435 & ~new_n436;
  assign new_n438 = new_n432 & ~new_n437;
  assign new_n439 = ~new_n432 & new_n437;
  assign new_n440 = ~new_n438 & ~new_n439;
  assign new_n441 = ~new_n401_1 & new_n440;
  assign new_n442 = new_n401_1 & ~new_n440;
  assign new_n443_1 = ~new_n441 & ~new_n442;
  assign new_n444 = n834 & n10168;
  assign new_n445 = n8716 & n12592;
  assign new_n446 = n3178 & n5189;
  assign new_n447 = ~new_n445 & ~new_n446;
  assign new_n448 = new_n445 & new_n446;
  assign new_n449 = ~new_n447 & ~new_n448;
  assign new_n450 = new_n444 & ~new_n449;
  assign new_n451 = ~new_n444 & new_n449;
  assign new_n452 = ~new_n450 & ~new_n451;
  assign new_n453 = ~new_n396_1 & new_n452;
  assign new_n454 = new_n396_1 & ~new_n452;
  assign new_n455 = ~new_n453 & ~new_n454;
  assign new_n456 = ~new_n443_1 & ~new_n455;
  assign new_n457 = new_n443_1 & new_n455;
  assign new_n458 = ~new_n456 & ~new_n457;
  assign new_n459 = ~new_n397 & ~new_n404;
  assign new_n460_1 = ~new_n403 & ~new_n459;
  assign new_n461 = ~new_n458 & ~new_n460_1;
  assign new_n462 = new_n458 & new_n460_1;
  assign new_n463 = ~new_n461 & ~new_n462;
  assign new_n464 = ~new_n431 & new_n463;
  assign new_n465 = new_n431 & ~new_n463;
  assign new_n466 = ~new_n464 & ~new_n465;
  assign new_n467 = ~new_n422 & new_n466;
  assign new_n468 = new_n422 & ~new_n466;
  assign n134 = ~new_n467 & ~new_n468;
  assign new_n470 = n3677 & n8228;
  assign new_n471 = n6937 & n8228;
  assign new_n472 = n1724 & n11236;
  assign new_n473 = n4382 & n10606;
  assign new_n474 = n11236 & n12965;
  assign new_n475 = new_n473 & new_n474;
  assign new_n476 = ~new_n473 & ~new_n474;
  assign new_n477 = n3130 & n10408;
  assign new_n478 = ~new_n476 & new_n477;
  assign new_n479 = ~new_n475 & ~new_n478;
  assign new_n480 = ~new_n472 & new_n479;
  assign new_n481 = new_n472 & ~new_n479;
  assign new_n482 = ~new_n480 & ~new_n481;
  assign new_n483 = n9732 & n10408;
  assign new_n484 = n4382 & n12965;
  assign new_n485 = n3130 & n10606;
  assign new_n486 = ~new_n484 & ~new_n485;
  assign new_n487 = new_n484 & new_n485;
  assign new_n488 = ~new_n486 & ~new_n487;
  assign new_n489 = new_n483 & ~new_n488;
  assign new_n490 = ~new_n483 & new_n488;
  assign new_n491 = ~new_n489 & ~new_n490;
  assign new_n492 = ~new_n482 & new_n491;
  assign new_n493 = new_n482 & ~new_n491;
  assign new_n494 = ~new_n492 & ~new_n493;
  assign new_n495 = new_n471 & new_n494;
  assign new_n496 = ~new_n471 & ~new_n494;
  assign new_n497_1 = n1724 & n8228;
  assign new_n498 = n10606 & n11236;
  assign new_n499_1 = n8228 & n12965;
  assign new_n500 = new_n498 & new_n499_1;
  assign new_n501 = ~new_n498 & ~new_n499_1;
  assign new_n502 = n4382 & n10408;
  assign new_n503 = ~new_n501 & new_n502;
  assign new_n504 = ~new_n500 & ~new_n503;
  assign new_n505 = ~new_n497_1 & new_n504;
  assign new_n506 = new_n497_1 & ~new_n504;
  assign new_n507 = ~new_n475 & ~new_n476;
  assign new_n508 = ~new_n477 & ~new_n507;
  assign new_n509 = new_n477 & new_n507;
  assign new_n510_1 = ~new_n508 & ~new_n509;
  assign new_n511 = ~new_n506 & ~new_n510_1;
  assign new_n512 = ~new_n505 & ~new_n511;
  assign new_n513 = ~new_n496 & new_n512;
  assign new_n514 = ~new_n495 & ~new_n513;
  assign new_n515 = n1724 & n4382;
  assign new_n516 = n6937 & n11236;
  assign new_n517 = ~new_n515 & ~new_n516;
  assign new_n518 = new_n515 & new_n516;
  assign new_n519 = ~new_n517 & ~new_n518;
  assign new_n520 = n3130 & n12965;
  assign new_n521 = n9732 & n10606;
  assign new_n522 = n103 & n10408;
  assign new_n523 = new_n521 & new_n522;
  assign new_n524 = ~new_n521 & ~new_n522;
  assign new_n525 = ~new_n523 & ~new_n524;
  assign new_n526 = ~new_n520 & ~new_n525;
  assign new_n527 = new_n520 & new_n525;
  assign new_n528 = ~new_n526 & ~new_n527;
  assign new_n529 = new_n483 & ~new_n486;
  assign new_n530 = ~new_n487 & ~new_n529;
  assign new_n531 = ~new_n528 & ~new_n530;
  assign new_n532 = new_n528 & new_n530;
  assign new_n533 = ~new_n531 & ~new_n532;
  assign new_n534 = ~new_n519 & new_n533;
  assign new_n535 = new_n519 & ~new_n533;
  assign new_n536 = ~new_n534 & ~new_n535;
  assign new_n537_1 = ~new_n481 & new_n491;
  assign new_n538 = ~new_n480 & ~new_n537_1;
  assign new_n539 = ~new_n536 & ~new_n538;
  assign new_n540 = new_n536 & new_n538;
  assign new_n541 = ~new_n539 & ~new_n540;
  assign new_n542 = ~new_n514 & new_n541;
  assign new_n543 = new_n514 & ~new_n541;
  assign new_n544 = ~new_n542 & ~new_n543;
  assign new_n545 = new_n470 & new_n544;
  assign new_n546 = n8228 & n10606;
  assign new_n547 = n10408 & n11236;
  assign new_n548 = new_n546 & new_n547;
  assign new_n549 = ~new_n500 & ~new_n501;
  assign new_n550 = ~new_n502 & ~new_n549;
  assign new_n551 = new_n502 & new_n549;
  assign new_n552 = ~new_n550 & ~new_n551;
  assign new_n553 = new_n548 & new_n552;
  assign new_n554 = ~new_n505 & ~new_n506;
  assign new_n555 = ~new_n510_1 & ~new_n554;
  assign new_n556 = new_n510_1 & new_n554;
  assign new_n557 = ~new_n555 & ~new_n556;
  assign new_n558 = new_n553 & new_n557;
  assign new_n559 = ~new_n495 & ~new_n496;
  assign new_n560 = new_n512 & new_n559;
  assign new_n561 = ~new_n512 & ~new_n559;
  assign new_n562 = ~new_n560 & ~new_n561;
  assign new_n563 = new_n558 & new_n562;
  assign new_n564 = ~new_n470 & ~new_n544;
  assign new_n565 = ~new_n545 & ~new_n564;
  assign new_n566 = new_n563 & new_n565;
  assign new_n567 = ~new_n545 & ~new_n566;
  assign new_n568 = n4382 & n6937;
  assign new_n569 = n7729 & n8228;
  assign new_n570 = n3677 & n11236;
  assign new_n571 = ~new_n569 & ~new_n570;
  assign new_n572 = new_n569 & new_n570;
  assign new_n573_1 = ~new_n571 & ~new_n572;
  assign new_n574 = ~new_n568 & ~new_n573_1;
  assign new_n575 = new_n568 & new_n573_1;
  assign new_n576 = ~new_n574 & ~new_n575;
  assign new_n577 = ~new_n527 & new_n530;
  assign new_n578 = ~new_n526 & ~new_n577;
  assign new_n579 = new_n576 & new_n578;
  assign new_n580 = ~new_n576 & ~new_n578;
  assign new_n581 = ~new_n579 & ~new_n580;
  assign new_n582 = n1724 & n3130;
  assign new_n583 = ~new_n523 & ~new_n582;
  assign new_n584 = new_n523 & new_n582;
  assign new_n585 = ~new_n583 & ~new_n584;
  assign new_n586 = n5320 & n10408;
  assign new_n587 = n103 & n10606;
  assign new_n588 = n9732 & n12965;
  assign new_n589 = ~new_n587 & ~new_n588;
  assign new_n590 = new_n587 & new_n588;
  assign new_n591 = ~new_n589 & ~new_n590;
  assign new_n592 = new_n586 & ~new_n591;
  assign new_n593 = ~new_n586 & new_n591;
  assign new_n594 = ~new_n592 & ~new_n593;
  assign new_n595 = ~new_n585 & new_n594;
  assign new_n596 = new_n585 & ~new_n594;
  assign new_n597 = ~new_n595 & ~new_n596;
  assign new_n598 = new_n581 & new_n597;
  assign new_n599 = ~new_n581 & ~new_n597;
  assign new_n600 = ~new_n598 & ~new_n599;
  assign new_n601 = new_n518 & new_n600;
  assign new_n602 = ~new_n518 & ~new_n600;
  assign new_n603_1 = ~new_n601 & ~new_n602;
  assign new_n604 = ~new_n534 & new_n538;
  assign new_n605 = ~new_n535 & ~new_n604;
  assign new_n606 = new_n603_1 & new_n605;
  assign new_n607 = ~new_n603_1 & ~new_n605;
  assign new_n608 = ~new_n606 & ~new_n607;
  assign new_n609 = new_n542 & ~new_n608;
  assign new_n610 = ~new_n542 & new_n608;
  assign new_n611 = ~new_n609 & ~new_n610;
  assign new_n612 = ~new_n567 & new_n611;
  assign new_n613 = new_n567 & ~new_n611;
  assign new_n614 = ~new_n612 & ~new_n613;
  assign new_n615 = n3112 & n8940;
  assign new_n616 = n2174 & n8940;
  assign new_n617 = n8233 & n10770;
  assign new_n618 = n4335 & n10522;
  assign new_n619 = n5684 & n9887;
  assign new_n620 = ~new_n618 & ~new_n619;
  assign new_n621 = new_n618 & new_n619;
  assign new_n622 = ~new_n620 & ~new_n621;
  assign new_n623 = ~new_n617 & ~new_n622;
  assign new_n624 = new_n617 & new_n622;
  assign new_n625 = ~new_n623 & ~new_n624;
  assign new_n626 = n497 & n4964;
  assign new_n627 = n4335 & n5684;
  assign new_n628 = n4964 & n9887;
  assign new_n629 = new_n627 & new_n628;
  assign new_n630 = ~new_n627 & ~new_n628;
  assign new_n631 = n8233 & n10522;
  assign new_n632 = ~new_n630 & new_n631;
  assign new_n633 = ~new_n629 & ~new_n632;
  assign new_n634 = new_n626 & ~new_n633;
  assign new_n635 = ~new_n626 & new_n633;
  assign new_n636 = ~new_n634 & ~new_n635;
  assign new_n637 = new_n625 & ~new_n636;
  assign new_n638 = ~new_n625 & new_n636;
  assign new_n639 = ~new_n637 & ~new_n638;
  assign new_n640 = new_n616 & ~new_n639;
  assign new_n641 = ~new_n616 & new_n639;
  assign new_n642 = n497 & n8940;
  assign new_n643 = n4335 & n4964;
  assign new_n644 = n8940 & n9887;
  assign new_n645 = new_n643 & new_n644;
  assign new_n646 = ~new_n643 & ~new_n644;
  assign new_n647 = n5684 & n8233;
  assign new_n648 = ~new_n646 & new_n647;
  assign new_n649 = ~new_n645 & ~new_n648;
  assign new_n650 = ~new_n642 & new_n649;
  assign new_n651 = new_n642 & ~new_n649;
  assign new_n652 = ~new_n629 & ~new_n630;
  assign new_n653 = ~new_n631 & ~new_n652;
  assign new_n654 = new_n631 & new_n652;
  assign new_n655 = ~new_n653 & ~new_n654;
  assign new_n656 = ~new_n651 & ~new_n655;
  assign new_n657 = ~new_n650 & ~new_n656;
  assign new_n658 = ~new_n641 & new_n657;
  assign new_n659 = ~new_n640 & ~new_n658;
  assign new_n660 = n497 & n5684;
  assign new_n661 = n2174 & n4964;
  assign new_n662 = new_n660 & new_n661;
  assign new_n663 = ~new_n660 & ~new_n661;
  assign new_n664 = ~new_n662 & ~new_n663;
  assign new_n665 = n9887 & n10522;
  assign new_n666 = n4335 & n10770;
  assign new_n667 = n8233 & new_n666;
  assign new_n668 = ~new_n617 & ~new_n666;
  assign new_n669 = ~new_n667 & ~new_n668;
  assign new_n670 = ~new_n665 & ~new_n669;
  assign new_n671 = new_n665 & new_n669;
  assign new_n672 = ~new_n670 & ~new_n671;
  assign new_n673 = new_n617 & ~new_n620;
  assign new_n674 = ~new_n621 & ~new_n673;
  assign new_n675 = ~new_n672 & new_n674;
  assign new_n676 = new_n672 & ~new_n674;
  assign new_n677 = ~new_n675 & ~new_n676;
  assign new_n678 = ~new_n664 & ~new_n677;
  assign new_n679 = new_n664 & new_n677;
  assign new_n680 = ~new_n678 & ~new_n679;
  assign new_n681 = ~new_n625 & ~new_n634;
  assign new_n682 = ~new_n635 & ~new_n681;
  assign new_n683 = ~new_n680 & ~new_n682;
  assign new_n684 = new_n680 & new_n682;
  assign new_n685 = ~new_n683 & ~new_n684;
  assign new_n686 = ~new_n659 & new_n685;
  assign new_n687 = new_n659 & ~new_n685;
  assign new_n688 = ~new_n686 & ~new_n687;
  assign new_n689 = new_n615 & new_n688;
  assign new_n690 = n4335 & n8940;
  assign new_n691 = n4964 & n8233;
  assign new_n692 = new_n690 & new_n691;
  assign new_n693 = ~new_n645 & ~new_n646;
  assign new_n694 = ~new_n647 & ~new_n693;
  assign new_n695 = new_n647 & new_n693;
  assign new_n696 = ~new_n694 & ~new_n695;
  assign new_n697 = new_n692 & new_n696;
  assign new_n698 = ~new_n650 & ~new_n651;
  assign new_n699 = ~new_n655 & ~new_n698;
  assign new_n700 = new_n655 & new_n698;
  assign new_n701 = ~new_n699 & ~new_n700;
  assign new_n702 = new_n697 & new_n701;
  assign new_n703 = ~new_n640 & ~new_n641;
  assign new_n704 = ~new_n657 & ~new_n703;
  assign new_n705 = new_n657 & new_n703;
  assign new_n706 = ~new_n704 & ~new_n705;
  assign new_n707 = new_n702 & new_n706;
  assign new_n708 = ~new_n615 & ~new_n688;
  assign new_n709 = ~new_n689 & ~new_n708;
  assign new_n710 = new_n707 & new_n709;
  assign new_n711 = ~new_n689 & ~new_n710;
  assign new_n712 = ~new_n678 & new_n682;
  assign new_n713 = new_n662 & new_n712;
  assign new_n714 = ~new_n662 & ~new_n712;
  assign new_n715 = ~new_n679 & new_n714;
  assign new_n716 = ~new_n713 & ~new_n715;
  assign new_n717 = ~new_n670 & ~new_n674;
  assign new_n718 = ~new_n671 & ~new_n717;
  assign new_n719 = n2174 & n5684;
  assign new_n720 = n4964 & new_n615;
  assign new_n721 = n3112 & n4964;
  assign new_n722 = ~new_n615 & ~new_n721;
  assign new_n723 = ~new_n720 & ~new_n722;
  assign new_n724 = ~new_n719 & new_n723;
  assign new_n725 = new_n719 & ~new_n723;
  assign new_n726 = ~new_n724 & ~new_n725;
  assign new_n727 = ~new_n718 & ~new_n726;
  assign new_n728_1 = new_n718 & new_n726;
  assign new_n729 = ~new_n727 & ~new_n728_1;
  assign new_n730 = ~n9887 & new_n669;
  assign new_n731 = n9887 & n10770;
  assign new_n732 = ~new_n669 & new_n731;
  assign new_n733 = ~new_n730 & ~new_n732;
  assign new_n734 = n497 & n10522;
  assign new_n735 = new_n667 & new_n734;
  assign new_n736 = ~new_n667 & ~new_n734;
  assign new_n737 = ~new_n735 & ~new_n736;
  assign new_n738 = new_n733 & ~new_n737;
  assign new_n739 = ~new_n733 & new_n737;
  assign new_n740 = ~new_n738 & ~new_n739;
  assign new_n741 = new_n729 & new_n740;
  assign new_n742 = ~new_n729 & ~new_n740;
  assign new_n743 = ~new_n741 & ~new_n742;
  assign new_n744 = new_n716 & ~new_n743;
  assign new_n745 = ~new_n716 & new_n743;
  assign new_n746 = ~new_n744 & ~new_n745;
  assign new_n747 = new_n686 & ~new_n746;
  assign new_n748 = ~new_n686 & new_n746;
  assign new_n749 = ~new_n747 & ~new_n748;
  assign new_n750 = ~new_n711 & new_n749;
  assign new_n751 = new_n711 & ~new_n749;
  assign new_n752 = ~new_n750 & ~new_n751;
  assign new_n753 = n4357 & n9353;
  assign new_n754 = n2882 & n9353;
  assign new_n755 = n3832 & n6333;
  assign new_n756 = n1912 & n9915;
  assign new_n757 = n6333 & n8332;
  assign new_n758_1 = new_n756 & new_n757;
  assign new_n759 = ~new_n756 & ~new_n757;
  assign new_n760 = n10063 & n12750;
  assign new_n761_1 = ~new_n759 & new_n760;
  assign new_n762_1 = ~new_n758_1 & ~new_n761_1;
  assign new_n763 = ~new_n755 & new_n762_1;
  assign new_n764 = new_n755 & ~new_n762_1;
  assign new_n765 = ~new_n763 & ~new_n764;
  assign new_n766 = n9620 & n10063;
  assign new_n767_1 = n1912 & n8332;
  assign new_n768 = n9915 & n12750;
  assign new_n769 = ~new_n767_1 & ~new_n768;
  assign new_n770 = new_n767_1 & new_n768;
  assign new_n771 = ~new_n769 & ~new_n770;
  assign new_n772_1 = new_n766 & ~new_n771;
  assign new_n773 = ~new_n766 & new_n771;
  assign new_n774 = ~new_n772_1 & ~new_n773;
  assign new_n775 = ~new_n765 & new_n774;
  assign new_n776 = new_n765 & ~new_n774;
  assign new_n777_1 = ~new_n775 & ~new_n776;
  assign new_n778 = new_n754 & new_n777_1;
  assign new_n779 = ~new_n754 & ~new_n777_1;
  assign new_n780 = n3832 & n9353;
  assign new_n781 = n6333 & n9915;
  assign new_n782 = n8332 & n9353;
  assign new_n783 = new_n781 & new_n782;
  assign new_n784 = ~new_n781 & ~new_n782;
  assign new_n785 = n1912 & n10063;
  assign new_n786 = ~new_n784 & new_n785;
  assign new_n787 = ~new_n783 & ~new_n786;
  assign new_n788 = ~new_n780 & new_n787;
  assign new_n789 = new_n780 & ~new_n787;
  assign new_n790 = ~new_n758_1 & ~new_n759;
  assign new_n791 = ~new_n760 & ~new_n790;
  assign new_n792 = new_n760 & new_n790;
  assign new_n793 = ~new_n791 & ~new_n792;
  assign new_n794 = ~new_n789 & ~new_n793;
  assign new_n795 = ~new_n788 & ~new_n794;
  assign new_n796 = ~new_n779 & new_n795;
  assign new_n797 = ~new_n778 & ~new_n796;
  assign new_n798 = n1912 & n3832;
  assign new_n799 = n2882 & n6333;
  assign new_n800_1 = ~new_n798 & ~new_n799;
  assign new_n801 = new_n798 & new_n799;
  assign new_n802 = ~new_n800_1 & ~new_n801;
  assign new_n803 = n8332 & n12750;
  assign new_n804 = n761 & n10063;
  assign new_n805 = n9620 & n9915;
  assign new_n806 = ~new_n804 & ~new_n805;
  assign new_n807 = new_n804 & new_n805;
  assign new_n808 = ~new_n806 & ~new_n807;
  assign new_n809 = ~new_n803 & ~new_n808;
  assign new_n810 = new_n803 & new_n808;
  assign new_n811 = ~new_n809 & ~new_n810;
  assign new_n812 = new_n766 & ~new_n769;
  assign new_n813 = ~new_n770 & ~new_n812;
  assign new_n814 = ~new_n811 & new_n813;
  assign new_n815 = new_n811 & ~new_n813;
  assign new_n816 = ~new_n814 & ~new_n815;
  assign new_n817_1 = ~new_n802 & ~new_n816;
  assign new_n818 = new_n802 & new_n816;
  assign new_n819 = ~new_n817_1 & ~new_n818;
  assign new_n820 = ~new_n764 & new_n774;
  assign new_n821 = ~new_n763 & ~new_n820;
  assign new_n822 = ~new_n819 & ~new_n821;
  assign new_n823 = new_n819 & new_n821;
  assign new_n824 = ~new_n822 & ~new_n823;
  assign new_n825 = ~new_n797 & new_n824;
  assign new_n826 = new_n797 & ~new_n824;
  assign new_n827 = ~new_n825 & ~new_n826;
  assign new_n828 = new_n753 & new_n827;
  assign new_n829 = n9353 & n9915;
  assign new_n830 = n6333 & n10063;
  assign new_n831_1 = new_n829 & new_n830;
  assign new_n832 = ~new_n783 & ~new_n784;
  assign new_n833 = ~new_n785 & ~new_n832;
  assign new_n834_1 = new_n785 & new_n832;
  assign new_n835 = ~new_n833 & ~new_n834_1;
  assign new_n836 = new_n831_1 & new_n835;
  assign new_n837 = ~new_n788 & ~new_n789;
  assign new_n838 = ~new_n793 & ~new_n837;
  assign new_n839 = new_n793 & new_n837;
  assign new_n840 = ~new_n838 & ~new_n839;
  assign new_n841 = new_n836 & new_n840;
  assign new_n842 = ~new_n778 & ~new_n779;
  assign new_n843 = new_n795 & new_n842;
  assign new_n844 = ~new_n795 & ~new_n842;
  assign new_n845 = ~new_n843 & ~new_n844;
  assign new_n846_1 = new_n841 & new_n845;
  assign new_n847 = ~new_n753 & ~new_n827;
  assign new_n848 = ~new_n828 & ~new_n847;
  assign new_n849 = new_n846_1 & new_n848;
  assign new_n850 = ~new_n828 & ~new_n849;
  assign new_n851 = ~new_n817_1 & new_n821;
  assign new_n852 = ~new_n801 & ~new_n851;
  assign new_n853 = ~new_n818 & new_n852;
  assign new_n854_1 = new_n801 & new_n851;
  assign new_n855 = ~new_n853 & ~new_n854_1;
  assign new_n856 = n1912 & n2882;
  assign new_n857 = n1165 & n9353;
  assign new_n858 = n4357 & n6333;
  assign new_n859 = ~new_n857 & ~new_n858;
  assign new_n860 = new_n857 & new_n858;
  assign new_n861 = ~new_n859 & ~new_n860;
  assign new_n862 = new_n856 & ~new_n861;
  assign new_n863 = ~new_n856 & new_n861;
  assign new_n864 = ~new_n862 & ~new_n863;
  assign new_n865 = ~new_n810 & new_n813;
  assign new_n866 = ~new_n809 & ~new_n865;
  assign new_n867 = new_n864 & ~new_n866;
  assign new_n868 = n3832 & n12750;
  assign new_n869 = new_n807 & new_n868;
  assign new_n870 = ~new_n807 & ~new_n868;
  assign new_n871 = ~new_n869 & ~new_n870;
  assign new_n872 = n5758 & n10063;
  assign new_n873 = n761 & n9915;
  assign new_n874 = n8332 & n9620;
  assign new_n875 = ~new_n873 & ~new_n874;
  assign new_n876 = new_n873 & new_n874;
  assign new_n877 = ~new_n875 & ~new_n876;
  assign new_n878 = new_n872 & ~new_n877;
  assign new_n879 = ~new_n872 & new_n877;
  assign new_n880 = ~new_n878 & ~new_n879;
  assign new_n881 = new_n871 & new_n880;
  assign new_n882 = ~new_n871 & ~new_n880;
  assign new_n883 = ~new_n881 & ~new_n882;
  assign new_n884 = new_n867 & new_n883;
  assign new_n885 = ~new_n864 & new_n866;
  assign new_n886 = ~new_n883 & new_n885;
  assign new_n887 = ~new_n867 & ~new_n883;
  assign new_n888 = ~new_n885 & ~new_n887;
  assign new_n889 = ~new_n886 & ~new_n888;
  assign new_n890 = ~new_n884 & ~new_n889;
  assign new_n891 = new_n855 & ~new_n890;
  assign new_n892 = ~new_n855 & new_n890;
  assign new_n893 = ~new_n891 & ~new_n892;
  assign new_n894 = new_n825 & ~new_n893;
  assign new_n895 = ~new_n825 & new_n893;
  assign new_n896 = ~new_n894 & ~new_n895;
  assign new_n897 = ~new_n850 & new_n896;
  assign new_n898 = new_n850 & ~new_n896;
  assign new_n899 = ~new_n897 & ~new_n898;
  assign new_n900 = new_n752 & new_n899;
  assign new_n901 = ~new_n752 & ~new_n899;
  assign new_n902 = ~new_n900 & ~new_n901;
  assign new_n903 = ~new_n707 & ~new_n709;
  assign new_n904 = ~new_n710 & ~new_n903;
  assign new_n905 = ~new_n846_1 & ~new_n848;
  assign new_n906 = ~new_n849 & ~new_n905;
  assign new_n907 = new_n904 & new_n906;
  assign new_n908 = ~new_n904 & ~new_n906;
  assign new_n909 = ~new_n841 & ~new_n845;
  assign new_n910 = ~new_n846_1 & ~new_n909;
  assign new_n911 = ~new_n702 & ~new_n706;
  assign new_n912 = ~new_n707 & ~new_n911;
  assign new_n913 = new_n910 & new_n912;
  assign new_n914 = ~new_n910 & ~new_n912;
  assign new_n915 = ~new_n836 & ~new_n840;
  assign new_n916 = ~new_n841 & ~new_n915;
  assign new_n917 = ~new_n697 & ~new_n701;
  assign new_n918 = ~new_n702 & ~new_n917;
  assign new_n919 = new_n916 & new_n918;
  assign new_n920 = ~new_n916 & ~new_n918;
  assign new_n921 = ~new_n831_1 & ~new_n835;
  assign new_n922_1 = ~new_n836 & ~new_n921;
  assign new_n923 = ~new_n692 & ~new_n696;
  assign new_n924 = ~new_n697 & ~new_n923;
  assign new_n925 = new_n922_1 & new_n924;
  assign new_n926 = ~new_n922_1 & ~new_n924;
  assign new_n927_1 = n9353 & n10063;
  assign new_n928 = n8233 & n8940;
  assign new_n929 = new_n927_1 & new_n928;
  assign new_n930 = ~new_n690 & ~new_n691;
  assign new_n931 = ~new_n692 & ~new_n930;
  assign new_n932 = new_n929 & new_n931;
  assign new_n933 = ~new_n929 & ~new_n931;
  assign new_n934 = ~new_n829 & ~new_n830;
  assign new_n935 = ~new_n831_1 & ~new_n934;
  assign new_n936 = ~new_n933 & new_n935;
  assign new_n937_1 = ~new_n932 & ~new_n936;
  assign new_n938 = ~new_n926 & ~new_n937_1;
  assign new_n939 = ~new_n925 & ~new_n938;
  assign new_n940 = ~new_n920 & ~new_n939;
  assign new_n941 = ~new_n919 & ~new_n940;
  assign new_n942 = ~new_n914 & ~new_n941;
  assign new_n943 = ~new_n913 & ~new_n942;
  assign new_n944 = ~new_n908 & ~new_n943;
  assign new_n945 = ~new_n907 & ~new_n944;
  assign new_n946 = ~new_n902 & ~new_n945;
  assign new_n947 = new_n902 & new_n945;
  assign new_n948 = ~new_n946 & ~new_n947;
  assign new_n949 = new_n614 & ~new_n948;
  assign new_n950 = ~new_n614 & new_n948;
  assign new_n951_1 = ~new_n563 & ~new_n565;
  assign new_n952 = ~new_n566 & ~new_n951_1;
  assign new_n953 = ~new_n558 & ~new_n562;
  assign new_n954 = ~new_n563 & ~new_n953;
  assign new_n955 = ~new_n913 & ~new_n914;
  assign new_n956 = new_n941 & ~new_n955;
  assign new_n957 = ~new_n941 & new_n955;
  assign new_n958 = ~new_n956 & ~new_n957;
  assign new_n959 = new_n954 & new_n958;
  assign new_n960 = ~new_n954 & ~new_n958;
  assign new_n961 = ~new_n553 & ~new_n557;
  assign new_n962 = ~new_n558 & ~new_n961;
  assign new_n963 = ~new_n919 & ~new_n920;
  assign new_n964 = new_n939 & ~new_n963;
  assign new_n965 = ~new_n939 & new_n963;
  assign new_n966 = ~new_n964 & ~new_n965;
  assign new_n967 = new_n962 & new_n966;
  assign new_n968 = ~new_n962 & ~new_n966;
  assign new_n969 = ~new_n548 & ~new_n552;
  assign new_n970 = ~new_n553 & ~new_n969;
  assign new_n971 = ~new_n925 & ~new_n926;
  assign new_n972 = new_n937_1 & ~new_n971;
  assign new_n973 = ~new_n937_1 & new_n971;
  assign new_n974 = ~new_n972 & ~new_n973;
  assign new_n975 = new_n970 & new_n974;
  assign new_n976 = ~new_n970 & ~new_n974;
  assign new_n977 = ~new_n546 & ~new_n547;
  assign new_n978 = ~new_n548 & ~new_n977;
  assign new_n979 = ~new_n932 & ~new_n933;
  assign new_n980 = new_n935 & ~new_n979;
  assign new_n981 = ~new_n935 & new_n979;
  assign new_n982 = ~new_n980 & ~new_n981;
  assign new_n983 = new_n978 & ~new_n982;
  assign new_n984 = ~new_n978 & new_n982;
  assign new_n985_1 = n8228 & n10408;
  assign new_n986 = ~new_n927_1 & ~new_n928;
  assign new_n987 = ~new_n929 & ~new_n986;
  assign new_n988 = new_n985_1 & new_n987;
  assign new_n989 = ~new_n984 & new_n988;
  assign new_n990 = ~new_n983 & ~new_n989;
  assign new_n991 = ~new_n976 & ~new_n990;
  assign new_n992 = ~new_n975 & ~new_n991;
  assign new_n993 = ~new_n968 & ~new_n992;
  assign new_n994 = ~new_n967 & ~new_n993;
  assign new_n995 = ~new_n960 & ~new_n994;
  assign new_n996 = ~new_n959 & ~new_n995;
  assign new_n997 = new_n952 & ~new_n996;
  assign new_n998 = ~new_n952 & new_n996;
  assign new_n999 = ~new_n907 & ~new_n908;
  assign new_n1000 = new_n943 & ~new_n999;
  assign new_n1001 = ~new_n943 & new_n999;
  assign new_n1002 = ~new_n1000 & ~new_n1001;
  assign new_n1003 = ~new_n998 & new_n1002;
  assign new_n1004 = ~new_n997 & ~new_n1003;
  assign new_n1005 = ~new_n950 & ~new_n1004;
  assign new_n1006 = ~new_n949 & ~new_n1005;
  assign new_n1007_1 = ~new_n609 & ~new_n612;
  assign new_n1008 = new_n733 & ~new_n735;
  assign new_n1009 = ~new_n736 & ~new_n1008;
  assign new_n1010 = new_n1007_1 & new_n1009;
  assign new_n1011 = ~new_n1007_1 & ~new_n1009;
  assign new_n1012 = ~new_n1010 & ~new_n1011;
  assign new_n1013 = new_n1006 & ~new_n1012;
  assign new_n1014 = ~new_n1006 & new_n1012;
  assign new_n1015 = ~new_n1013 & ~new_n1014;
  assign new_n1016 = ~new_n747 & ~new_n750;
  assign new_n1017 = n1757 & n12306;
  assign new_n1018 = n4748 & n10113;
  assign new_n1019 = new_n1017 & new_n1018;
  assign new_n1020 = ~new_n1017 & ~new_n1018;
  assign new_n1021 = ~new_n1019 & ~new_n1020;
  assign new_n1022 = n4006 & n10416;
  assign new_n1023 = n4470 & n11488;
  assign new_n1024 = n2758 & n11030;
  assign new_n1025 = ~new_n1023 & ~new_n1024;
  assign new_n1026 = new_n1023 & new_n1024;
  assign new_n1027 = ~new_n1025 & ~new_n1026;
  assign new_n1028 = ~new_n1022 & ~new_n1027;
  assign new_n1029 = new_n1022 & new_n1027;
  assign new_n1030 = ~new_n1028 & ~new_n1029;
  assign new_n1031 = n2758 & n10416;
  assign new_n1032 = n1757 & n4006;
  assign new_n1033 = new_n1031 & new_n1032;
  assign new_n1034 = n4470 & n11030;
  assign new_n1035 = ~new_n1031 & ~new_n1032;
  assign new_n1036 = new_n1034 & ~new_n1035;
  assign new_n1037 = ~new_n1033 & ~new_n1036;
  assign new_n1038 = ~new_n1030 & new_n1037;
  assign new_n1039 = new_n1030 & ~new_n1037;
  assign new_n1040 = ~new_n1038 & ~new_n1039;
  assign new_n1041 = ~new_n1021 & ~new_n1040;
  assign new_n1042 = n10113 & n12306;
  assign new_n1043 = n1757 & n2758;
  assign new_n1044 = n4006 & n10113;
  assign new_n1045 = new_n1043 & new_n1044;
  assign new_n1046 = ~new_n1043 & ~new_n1044;
  assign new_n1047 = n4470 & n10416;
  assign new_n1048 = ~new_n1046 & new_n1047;
  assign new_n1049 = ~new_n1045 & ~new_n1048;
  assign new_n1050 = ~new_n1042 & new_n1049;
  assign new_n1051 = new_n1042 & ~new_n1049;
  assign new_n1052 = ~new_n1033 & ~new_n1035;
  assign new_n1053 = ~new_n1034 & ~new_n1052;
  assign new_n1054 = new_n1034 & new_n1052;
  assign new_n1055 = ~new_n1053 & ~new_n1054;
  assign new_n1056 = ~new_n1051 & ~new_n1055;
  assign new_n1057 = ~new_n1050 & ~new_n1056;
  assign new_n1058 = ~new_n1041 & new_n1057;
  assign new_n1059 = new_n1019 & new_n1058;
  assign new_n1060 = new_n1021 & new_n1040;
  assign new_n1061 = ~new_n1019 & ~new_n1058;
  assign new_n1062 = ~new_n1060 & new_n1061;
  assign new_n1063 = n1757 & n4748;
  assign new_n1064 = n1231 & n2482;
  assign new_n1065 = n9187 & n10113;
  assign new_n1066 = ~new_n1064 & ~new_n1065;
  assign new_n1067 = new_n1064 & new_n1065;
  assign new_n1068 = ~new_n1066 & ~new_n1067;
  assign new_n1069 = new_n1063 & ~new_n1068;
  assign new_n1070 = ~new_n1063 & new_n1068;
  assign new_n1071 = ~new_n1069 & ~new_n1070;
  assign new_n1072 = ~new_n1029 & new_n1037;
  assign new_n1073 = ~new_n1028 & ~new_n1072;
  assign new_n1074 = new_n1071 & ~new_n1073;
  assign new_n1075 = n10416 & n12306;
  assign new_n1076 = ~new_n1026 & ~new_n1075;
  assign new_n1077 = new_n1026 & new_n1075;
  assign new_n1078 = ~new_n1076 & ~new_n1077;
  assign new_n1079 = n1982 & n4470;
  assign new_n1080 = n2758 & n11488;
  assign new_n1081 = n4006 & n11030;
  assign new_n1082 = ~new_n1080 & ~new_n1081;
  assign new_n1083 = new_n1080 & new_n1081;
  assign new_n1084_1 = ~new_n1082 & ~new_n1083;
  assign new_n1085 = new_n1079 & ~new_n1084_1;
  assign new_n1086 = ~new_n1079 & new_n1084_1;
  assign new_n1087 = ~new_n1085 & ~new_n1086;
  assign new_n1088 = new_n1078 & new_n1087;
  assign new_n1089 = ~new_n1078 & ~new_n1087;
  assign new_n1090 = ~new_n1088 & ~new_n1089;
  assign new_n1091 = new_n1074 & new_n1090;
  assign new_n1092 = ~new_n1071 & new_n1073;
  assign new_n1093 = new_n1090 & ~new_n1092;
  assign new_n1094 = ~new_n1074 & ~new_n1093;
  assign new_n1095 = ~new_n1091 & ~new_n1094;
  assign new_n1096 = ~new_n1090 & new_n1092;
  assign new_n1097_1 = ~new_n1095 & ~new_n1096;
  assign new_n1098 = ~new_n1062 & ~new_n1097_1;
  assign new_n1099 = ~new_n1059 & ~new_n1098;
  assign new_n1100 = ~new_n580 & new_n597;
  assign new_n1101 = ~new_n579 & ~new_n1100;
  assign new_n1102 = ~new_n872 & ~new_n876;
  assign new_n1103 = ~new_n875 & ~new_n1102;
  assign new_n1104 = n9887 & ~new_n668;
  assign new_n1105 = ~new_n667 & ~new_n1104;
  assign new_n1106 = ~new_n1103 & new_n1105;
  assign new_n1107 = new_n1103 & ~new_n1105;
  assign new_n1108 = ~new_n1106 & ~new_n1107;
  assign new_n1109 = new_n1101 & ~new_n1108;
  assign new_n1110 = ~new_n1101 & new_n1108;
  assign new_n1111 = ~new_n1109 & ~new_n1110;
  assign new_n1112_1 = new_n1099 & ~new_n1111;
  assign new_n1113 = ~new_n1099 & new_n1111;
  assign new_n1114 = ~new_n1112_1 & ~new_n1113;
  assign new_n1115 = ~new_n1016 & ~new_n1114;
  assign new_n1116 = new_n1016 & new_n1114;
  assign new_n1117 = ~new_n1115 & ~new_n1116;
  assign new_n1118 = ~new_n901 & ~new_n945;
  assign new_n1119 = ~new_n900 & ~new_n1118;
  assign new_n1120 = n2482 & n3641;
  assign new_n1121 = n4006 & n11488;
  assign new_n1122 = n1982 & n2758;
  assign new_n1123 = ~new_n1121 & ~new_n1122;
  assign new_n1124 = new_n1121 & new_n1122;
  assign new_n1125 = ~new_n1123 & ~new_n1124;
  assign new_n1126 = n11030 & n12306;
  assign new_n1127 = n4748 & n10416;
  assign new_n1128 = new_n1126 & ~new_n1127;
  assign new_n1129 = ~new_n1126 & new_n1127;
  assign new_n1130 = ~new_n1128 & ~new_n1129;
  assign new_n1131 = ~new_n1125 & ~new_n1130;
  assign new_n1132 = new_n1125 & new_n1130;
  assign new_n1133 = ~new_n1131 & ~new_n1132;
  assign new_n1134 = ~new_n1120 & ~new_n1133;
  assign new_n1135 = new_n1120 & new_n1133;
  assign new_n1136 = ~new_n1134 & ~new_n1135;
  assign new_n1137 = n7729 & n11236;
  assign new_n1138 = n4470 & n8820;
  assign new_n1139 = new_n1137 & ~new_n1138;
  assign new_n1140 = ~new_n1137 & new_n1138;
  assign new_n1141 = ~new_n1139 & ~new_n1140;
  assign new_n1142 = n497 & n10770;
  assign new_n1143 = n2174 & n10522;
  assign new_n1144 = ~new_n1142 & ~new_n1143;
  assign new_n1145 = new_n1142 & new_n1143;
  assign new_n1146 = ~new_n1144 & ~new_n1145;
  assign new_n1147 = ~new_n1141 & new_n1146;
  assign new_n1148 = new_n1141 & ~new_n1146;
  assign new_n1149 = ~new_n1147 & ~new_n1148;
  assign new_n1150 = new_n1136 & new_n1149;
  assign new_n1151 = ~new_n1136 & ~new_n1149;
  assign new_n1152 = ~new_n1150 & ~new_n1151;
  assign new_n1153 = n3130 & n6937;
  assign new_n1154 = n10063 & n12352;
  assign new_n1155 = ~new_n1153 & new_n1154;
  assign new_n1156 = new_n1153 & ~new_n1154;
  assign new_n1157 = ~new_n1155 & ~new_n1156;
  assign new_n1158 = n3677 & n4382;
  assign new_n1159 = n5758 & n9915;
  assign new_n1160 = new_n1158 & ~new_n1159;
  assign new_n1161 = ~new_n1158 & new_n1159;
  assign new_n1162 = ~new_n1160 & ~new_n1161;
  assign new_n1163 = ~new_n1157 & ~new_n1162;
  assign new_n1164 = new_n1157 & new_n1162;
  assign new_n1165_1 = ~new_n1163 & ~new_n1164;
  assign new_n1166 = new_n586 & ~new_n589;
  assign new_n1167 = ~new_n590 & ~new_n1166;
  assign new_n1168 = ~new_n1165_1 & ~new_n1167;
  assign new_n1169 = new_n1165_1 & new_n1167;
  assign new_n1170 = ~new_n1168 & ~new_n1169;
  assign new_n1171 = n1231 & n10113;
  assign new_n1172 = n1757 & n9187;
  assign new_n1173 = new_n1171 & ~new_n1172;
  assign new_n1174 = ~new_n1171 & new_n1172;
  assign new_n1175 = ~new_n1173 & ~new_n1174;
  assign new_n1176 = n9353 & n10874;
  assign new_n1177 = n4964 & n5684;
  assign new_n1178 = ~n4964 & ~n5684;
  assign new_n1179 = ~new_n1177 & ~new_n1178;
  assign new_n1180 = n3112 & new_n1179;
  assign new_n1181_1 = new_n1176 & new_n1180;
  assign new_n1182 = ~new_n1176 & ~new_n1180;
  assign new_n1183 = ~new_n1181_1 & ~new_n1182;
  assign new_n1184 = new_n1175 & ~new_n1183;
  assign new_n1185 = ~new_n1175 & new_n1183;
  assign new_n1186 = ~new_n1184 & ~new_n1185;
  assign new_n1187 = ~new_n1170 & new_n1186;
  assign new_n1188 = new_n1170 & ~new_n1186;
  assign new_n1189 = ~new_n1187 & ~new_n1188;
  assign new_n1190 = new_n1152 & new_n1189;
  assign new_n1191 = ~new_n1152 & ~new_n1189;
  assign new_n1192 = ~new_n1190 & ~new_n1191;
  assign new_n1193 = n761 & n8332;
  assign new_n1194 = n3591 & n8940;
  assign new_n1195 = ~new_n1193 & ~new_n1194;
  assign new_n1196 = new_n1193 & new_n1194;
  assign new_n1197 = ~new_n1195 & ~new_n1196;
  assign new_n1198_1 = n3832 & n9620;
  assign new_n1199 = n2882 & n12750;
  assign new_n1200 = ~new_n1198_1 & ~new_n1199;
  assign new_n1201 = new_n1198_1 & new_n1199;
  assign new_n1202 = ~new_n1200 & ~new_n1201;
  assign new_n1203 = n1165 & n6333;
  assign new_n1204 = n1912 & n4357;
  assign new_n1205 = new_n1203 & ~new_n1204;
  assign new_n1206 = ~new_n1203 & new_n1204;
  assign new_n1207 = ~new_n1205 & ~new_n1206;
  assign new_n1208 = ~new_n1202 & new_n1207;
  assign new_n1209 = new_n1202 & ~new_n1207;
  assign new_n1210 = ~new_n1208 & ~new_n1209;
  assign new_n1211 = ~new_n1197 & new_n1210;
  assign new_n1212 = new_n1197 & ~new_n1210;
  assign new_n1213 = ~new_n1211 & ~new_n1212;
  assign new_n1214 = ~new_n1192 & new_n1213;
  assign new_n1215 = new_n1192 & ~new_n1213;
  assign new_n1216 = ~new_n1214 & ~new_n1215;
  assign new_n1217 = n5320 & n10606;
  assign new_n1218 = n603 & n8228;
  assign new_n1219 = new_n1217 & ~new_n1218;
  assign new_n1220 = ~new_n1217 & new_n1218;
  assign new_n1221 = ~new_n1219 & ~new_n1220;
  assign new_n1222 = n103 & n12965;
  assign new_n1223 = n1724 & n9732;
  assign new_n1224 = ~new_n1222 & ~new_n1223;
  assign new_n1225 = new_n1222 & new_n1223;
  assign new_n1226 = ~new_n1224 & ~new_n1225;
  assign new_n1227 = ~new_n1221 & new_n1226;
  assign new_n1228 = new_n1221 & ~new_n1226;
  assign new_n1229 = ~new_n1227 & ~new_n1228;
  assign new_n1230 = n4743 & n10408;
  assign new_n1231_1 = new_n733 & new_n1230;
  assign new_n1232 = ~new_n733 & ~new_n1230;
  assign new_n1233 = ~new_n1231_1 & ~new_n1232;
  assign new_n1234 = new_n1229 & new_n1233;
  assign new_n1235 = ~new_n1229 & ~new_n1233;
  assign new_n1236 = ~new_n1234 & ~new_n1235;
  assign new_n1237 = ~new_n1216 & new_n1236;
  assign new_n1238 = new_n1216 & ~new_n1236;
  assign new_n1239 = ~new_n1237 & ~new_n1238;
  assign new_n1240 = ~new_n1077 & new_n1087;
  assign new_n1241 = ~new_n1076 & ~new_n1240;
  assign new_n1242 = ~new_n602 & ~new_n605;
  assign new_n1243 = ~new_n601 & ~new_n1242;
  assign new_n1244 = new_n1241 & new_n1243;
  assign new_n1245 = ~new_n1241 & ~new_n1243;
  assign new_n1246 = ~new_n1244 & ~new_n1245;
  assign new_n1247 = new_n1239 & new_n1246;
  assign new_n1248 = ~new_n1239 & ~new_n1246;
  assign new_n1249 = ~new_n1247 & ~new_n1248;
  assign new_n1250 = ~new_n869 & new_n880;
  assign new_n1251 = ~new_n870 & ~new_n1250;
  assign new_n1252 = ~new_n1249 & new_n1251;
  assign new_n1253 = new_n1249 & ~new_n1251;
  assign new_n1254 = ~new_n1252 & ~new_n1253;
  assign new_n1255 = ~new_n1119 & new_n1254;
  assign new_n1256 = new_n1119 & ~new_n1254;
  assign new_n1257 = ~new_n1255 & ~new_n1256;
  assign new_n1258 = new_n888 & ~new_n1257;
  assign new_n1259 = ~new_n888 & new_n1257;
  assign new_n1260 = ~new_n1258 & ~new_n1259;
  assign new_n1261 = new_n1063 & ~new_n1066;
  assign new_n1262 = ~new_n1067 & ~new_n1261;
  assign new_n1263 = ~new_n1260 & new_n1262;
  assign new_n1264 = new_n1260 & ~new_n1262;
  assign new_n1265 = ~new_n1263 & ~new_n1264;
  assign new_n1266 = ~new_n1117 & new_n1265;
  assign new_n1267 = new_n1117 & ~new_n1265;
  assign new_n1268 = ~new_n1266 & ~new_n1267;
  assign new_n1269 = ~new_n1015 & new_n1268;
  assign new_n1270 = new_n1015 & ~new_n1268;
  assign new_n1271 = ~new_n1269 & ~new_n1270;
  assign new_n1272 = n2482 & n9187;
  assign new_n1273 = ~new_n1041 & ~new_n1060;
  assign new_n1274 = ~new_n1057 & ~new_n1273;
  assign new_n1275 = new_n1057 & new_n1273;
  assign new_n1276 = ~new_n1274 & ~new_n1275;
  assign new_n1277 = n2482 & n4748;
  assign new_n1278 = ~new_n1050 & ~new_n1051;
  assign new_n1279 = ~new_n1055 & new_n1278;
  assign new_n1280 = new_n1055 & ~new_n1278;
  assign new_n1281 = ~new_n1279 & ~new_n1280;
  assign new_n1282 = new_n1277 & ~new_n1281;
  assign new_n1283 = ~new_n1277 & new_n1281;
  assign new_n1284 = n2482 & n12306;
  assign new_n1285 = n2758 & n10113;
  assign new_n1286 = n2482 & n4006;
  assign new_n1287 = new_n1285 & new_n1286;
  assign new_n1288 = ~new_n1285 & ~new_n1286;
  assign new_n1289 = n1757 & n4470;
  assign new_n1290 = ~new_n1288 & new_n1289;
  assign new_n1291 = ~new_n1287 & ~new_n1290;
  assign new_n1292 = ~new_n1284 & new_n1291;
  assign new_n1293 = new_n1284 & ~new_n1291;
  assign new_n1294 = ~new_n1045 & ~new_n1046;
  assign new_n1295 = ~new_n1047 & ~new_n1294;
  assign new_n1296 = new_n1047 & new_n1294;
  assign new_n1297 = ~new_n1295 & ~new_n1296;
  assign new_n1298 = ~new_n1293 & ~new_n1297;
  assign new_n1299 = ~new_n1292 & ~new_n1298;
  assign new_n1300 = ~new_n1283 & new_n1299;
  assign new_n1301 = ~new_n1282 & ~new_n1300;
  assign new_n1302_1 = new_n1276 & ~new_n1301;
  assign new_n1303 = ~new_n1276 & new_n1301;
  assign new_n1304 = ~new_n1302_1 & ~new_n1303;
  assign new_n1305 = new_n1272 & new_n1304;
  assign new_n1306 = n2482 & n2758;
  assign new_n1307_1 = n4470 & n10113;
  assign new_n1308 = new_n1306 & new_n1307_1;
  assign new_n1309 = ~new_n1287 & ~new_n1288;
  assign new_n1310 = ~new_n1289 & ~new_n1309;
  assign new_n1311 = new_n1289 & new_n1309;
  assign new_n1312 = ~new_n1310 & ~new_n1311;
  assign new_n1313 = new_n1308 & new_n1312;
  assign new_n1314 = ~new_n1292 & ~new_n1293;
  assign new_n1315 = ~new_n1297 & ~new_n1314;
  assign new_n1316 = new_n1297 & new_n1314;
  assign new_n1317 = ~new_n1315 & ~new_n1316;
  assign new_n1318 = new_n1313 & new_n1317;
  assign new_n1319 = ~new_n1282 & ~new_n1283;
  assign new_n1320 = ~new_n1299 & ~new_n1319;
  assign new_n1321 = new_n1299 & new_n1319;
  assign new_n1322 = ~new_n1320 & ~new_n1321;
  assign new_n1323 = new_n1318 & new_n1322;
  assign new_n1324 = ~new_n1272 & ~new_n1304;
  assign new_n1325 = ~new_n1305 & ~new_n1324;
  assign new_n1326 = new_n1323 & new_n1325;
  assign new_n1327 = ~new_n1305 & ~new_n1326;
  assign new_n1328 = ~new_n1059 & ~new_n1062;
  assign new_n1329 = new_n1097_1 & new_n1328;
  assign new_n1330 = ~new_n1097_1 & ~new_n1328;
  assign new_n1331 = ~new_n1329 & ~new_n1330;
  assign new_n1332 = new_n1302_1 & ~new_n1331;
  assign new_n1333 = ~new_n1302_1 & new_n1331;
  assign new_n1334 = ~new_n1332 & ~new_n1333;
  assign new_n1335 = ~new_n1327 & new_n1334;
  assign new_n1336 = new_n1327 & ~new_n1334;
  assign new_n1337 = ~new_n1335 & ~new_n1336;
  assign new_n1338 = ~new_n949 & ~new_n950;
  assign new_n1339 = new_n1004 & new_n1338;
  assign new_n1340 = ~new_n1004 & ~new_n1338;
  assign new_n1341 = ~new_n1339 & ~new_n1340;
  assign new_n1342 = ~new_n1337 & new_n1341;
  assign new_n1343 = new_n1337 & ~new_n1341;
  assign new_n1344 = ~new_n1323 & ~new_n1325;
  assign new_n1345 = ~new_n1326 & ~new_n1344;
  assign new_n1346 = ~new_n997 & ~new_n998;
  assign new_n1347 = ~new_n1002 & ~new_n1346;
  assign new_n1348 = new_n1002 & new_n1346;
  assign new_n1349 = ~new_n1347 & ~new_n1348;
  assign new_n1350 = new_n1345 & new_n1349;
  assign new_n1351 = ~new_n1345 & ~new_n1349;
  assign new_n1352 = ~new_n1318 & ~new_n1322;
  assign new_n1353 = ~new_n1323 & ~new_n1352;
  assign new_n1354 = ~new_n959 & ~new_n960;
  assign new_n1355 = new_n994 & ~new_n1354;
  assign new_n1356 = ~new_n994 & new_n1354;
  assign new_n1357 = ~new_n1355 & ~new_n1356;
  assign new_n1358 = ~new_n1353 & ~new_n1357;
  assign new_n1359 = new_n1353 & new_n1357;
  assign new_n1360 = ~new_n1313 & ~new_n1317;
  assign new_n1361 = ~new_n1318 & ~new_n1360;
  assign new_n1362 = ~new_n967 & ~new_n968;
  assign new_n1363 = new_n992 & ~new_n1362;
  assign new_n1364_1 = ~new_n992 & new_n1362;
  assign new_n1365 = ~new_n1363 & ~new_n1364_1;
  assign new_n1366 = ~new_n1361 & ~new_n1365;
  assign new_n1367 = new_n1361 & new_n1365;
  assign new_n1368 = ~new_n1308 & ~new_n1312;
  assign new_n1369 = ~new_n1313 & ~new_n1368;
  assign new_n1370 = ~new_n975 & ~new_n976;
  assign new_n1371 = new_n990 & ~new_n1370;
  assign new_n1372 = ~new_n990 & new_n1370;
  assign new_n1373 = ~new_n1371 & ~new_n1372;
  assign new_n1374 = ~new_n1369 & ~new_n1373;
  assign new_n1375 = new_n1369 & new_n1373;
  assign new_n1376 = ~new_n1306 & ~new_n1307_1;
  assign new_n1377 = ~new_n1308 & ~new_n1376;
  assign new_n1378 = n2482 & n4470;
  assign new_n1379 = ~new_n985_1 & ~new_n987;
  assign new_n1380 = ~new_n988 & ~new_n1379;
  assign new_n1381 = new_n1378 & new_n1380;
  assign new_n1382 = ~new_n1377 & ~new_n1381;
  assign new_n1383 = new_n1377 & new_n1381;
  assign new_n1384 = ~new_n983 & ~new_n984;
  assign new_n1385 = ~new_n988 & ~new_n1384;
  assign new_n1386 = new_n988 & new_n1384;
  assign new_n1387 = ~new_n1385 & ~new_n1386;
  assign new_n1388 = ~new_n1383 & ~new_n1387;
  assign new_n1389 = ~new_n1382 & ~new_n1388;
  assign new_n1390 = ~new_n1375 & ~new_n1389;
  assign new_n1391 = ~new_n1374 & ~new_n1390;
  assign new_n1392_1 = ~new_n1367 & ~new_n1391;
  assign new_n1393 = ~new_n1366 & ~new_n1392_1;
  assign new_n1394 = ~new_n1359 & ~new_n1393;
  assign new_n1395 = ~new_n1358 & ~new_n1394;
  assign new_n1396 = ~new_n1351 & new_n1395;
  assign new_n1397 = ~new_n1350 & ~new_n1396;
  assign new_n1398 = ~new_n1343 & new_n1397;
  assign new_n1399 = ~new_n1342 & ~new_n1398;
  assign new_n1400 = ~new_n1332 & ~new_n1335;
  assign new_n1401_1 = ~new_n584 & new_n594;
  assign new_n1402 = ~new_n583 & ~new_n1401_1;
  assign new_n1403 = ~new_n1400 & new_n1402;
  assign new_n1404 = new_n1400 & ~new_n1402;
  assign new_n1405 = ~new_n1403 & ~new_n1404;
  assign new_n1406 = ~new_n894 & ~new_n897;
  assign new_n1407 = ~new_n853 & new_n890;
  assign new_n1408 = ~new_n854_1 & ~new_n1407;
  assign new_n1409 = new_n856 & ~new_n859;
  assign new_n1410 = ~new_n860 & ~new_n1409;
  assign new_n1411 = ~new_n1408 & new_n1410;
  assign new_n1412 = new_n1408 & ~new_n1410;
  assign new_n1413 = ~new_n1411 & ~new_n1412;
  assign new_n1414 = new_n1406 & ~new_n1413;
  assign new_n1415 = ~new_n1406 & new_n1413;
  assign new_n1416 = ~new_n1414 & ~new_n1415;
  assign new_n1417 = ~new_n1405 & new_n1416;
  assign new_n1418 = new_n1405 & ~new_n1416;
  assign new_n1419 = ~new_n1417 & ~new_n1418;
  assign new_n1420 = ~new_n715 & new_n743;
  assign new_n1421 = ~new_n713 & ~new_n1420;
  assign new_n1422 = ~new_n719 & ~new_n720;
  assign new_n1423 = ~new_n722 & ~new_n1422;
  assign new_n1424 = ~new_n728_1 & new_n740;
  assign new_n1425 = ~new_n727 & ~new_n1424;
  assign new_n1426 = new_n1079 & ~new_n1082;
  assign new_n1427 = ~new_n1083 & ~new_n1426;
  assign new_n1428 = new_n568 & ~new_n571;
  assign new_n1429 = ~new_n572 & ~new_n1428;
  assign new_n1430 = ~new_n1427 & new_n1429;
  assign new_n1431 = new_n1427 & ~new_n1429;
  assign new_n1432 = ~new_n1430 & ~new_n1431;
  assign new_n1433 = new_n1425 & ~new_n1432;
  assign new_n1434 = ~new_n1425 & new_n1432;
  assign new_n1435 = ~new_n1433 & ~new_n1434;
  assign new_n1436 = ~new_n1423 & new_n1435;
  assign new_n1437 = new_n1423 & ~new_n1435;
  assign new_n1438 = ~new_n1436 & ~new_n1437;
  assign new_n1439 = ~new_n1421 & new_n1438;
  assign new_n1440 = new_n1421 & ~new_n1438;
  assign new_n1441 = ~new_n1439 & ~new_n1440;
  assign new_n1442 = new_n1094 & ~new_n1441;
  assign new_n1443 = ~new_n1094 & new_n1441;
  assign new_n1444 = ~new_n1442 & ~new_n1443;
  assign new_n1445 = ~new_n1419 & new_n1444;
  assign new_n1446 = new_n1419 & ~new_n1444;
  assign new_n1447 = ~new_n1445 & ~new_n1446;
  assign new_n1448 = new_n1399 & new_n1447;
  assign new_n1449 = ~new_n1399 & ~new_n1447;
  assign new_n1450 = ~new_n1448 & ~new_n1449;
  assign new_n1451 = new_n1271 & new_n1450;
  assign new_n1452 = ~new_n1271 & ~new_n1450;
  assign n201 = new_n1451 | new_n1452;
  assign new_n1454 = n3006 & n12853;
  assign new_n1455 = n854 & n5801;
  assign new_n1456 = n510 & n5671;
  assign new_n1457 = n834 & n13201;
  assign new_n1458 = new_n1456 & new_n1457;
  assign new_n1459 = ~new_n1456 & ~new_n1457;
  assign new_n1460 = ~new_n1458 & ~new_n1459;
  assign new_n1461 = new_n1455 & new_n1460;
  assign new_n1462 = ~new_n1455 & ~new_n1460;
  assign new_n1463 = ~new_n1461 & ~new_n1462;
  assign new_n1464 = new_n1454 & new_n1463;
  assign new_n1465 = ~new_n1454 & ~new_n1463;
  assign n211 = ~new_n1464 & ~new_n1465;
  assign new_n1467 = n2758 & n3006;
  assign new_n1468 = n4470 & n5568;
  assign new_n1469 = new_n1467 & new_n1468;
  assign new_n1470 = n4470 & n8308;
  assign new_n1471 = n2758 & n5568;
  assign new_n1472 = n3006 & n4006;
  assign new_n1473 = ~new_n1471 & ~new_n1472;
  assign new_n1474 = new_n1471 & new_n1472;
  assign new_n1475 = ~new_n1473 & ~new_n1474;
  assign new_n1476 = new_n1470 & ~new_n1475;
  assign new_n1477 = ~new_n1470 & new_n1475;
  assign new_n1478 = ~new_n1476 & ~new_n1477;
  assign new_n1479 = new_n1469 & ~new_n1478;
  assign new_n1480 = n3006 & n12306;
  assign new_n1481 = new_n1470 & ~new_n1473;
  assign new_n1482 = ~new_n1474 & ~new_n1481;
  assign new_n1483 = ~new_n1480 & new_n1482;
  assign new_n1484 = new_n1480 & ~new_n1482;
  assign new_n1485 = ~new_n1483 & ~new_n1484;
  assign new_n1486 = n4470 & n5214;
  assign new_n1487_1 = n4006 & n5568;
  assign new_n1488 = n2758 & n8308;
  assign new_n1489 = ~new_n1487_1 & ~new_n1488;
  assign new_n1490 = new_n1487_1 & new_n1488;
  assign new_n1491 = ~new_n1489 & ~new_n1490;
  assign new_n1492 = new_n1486 & ~new_n1491;
  assign new_n1493 = ~new_n1486 & new_n1491;
  assign new_n1494 = ~new_n1492 & ~new_n1493;
  assign new_n1495 = ~new_n1485 & new_n1494;
  assign new_n1496 = new_n1485 & ~new_n1494;
  assign new_n1497 = ~new_n1495 & ~new_n1496;
  assign new_n1498 = new_n1479 & new_n1497;
  assign new_n1499 = n3006 & n4748;
  assign new_n1500 = n5568 & n12306;
  assign new_n1501 = new_n1486 & ~new_n1489;
  assign new_n1502 = ~new_n1490 & ~new_n1501;
  assign new_n1503 = ~new_n1500 & new_n1502;
  assign new_n1504 = new_n1500 & ~new_n1502;
  assign new_n1505 = ~new_n1503 & ~new_n1504;
  assign new_n1506 = n2771 & n4470;
  assign new_n1507 = n4006 & n8308;
  assign new_n1508 = n2758 & n5214;
  assign new_n1509 = ~new_n1507 & ~new_n1508;
  assign new_n1510 = new_n1507 & new_n1508;
  assign new_n1511 = ~new_n1509 & ~new_n1510;
  assign new_n1512 = new_n1506 & ~new_n1511;
  assign new_n1513 = ~new_n1506 & new_n1511;
  assign new_n1514 = ~new_n1512 & ~new_n1513;
  assign new_n1515 = ~new_n1505 & new_n1514;
  assign new_n1516 = new_n1505 & ~new_n1514;
  assign new_n1517 = ~new_n1515 & ~new_n1516;
  assign new_n1518 = ~new_n1499 & ~new_n1517;
  assign new_n1519 = new_n1499 & new_n1517;
  assign new_n1520 = ~new_n1518 & ~new_n1519;
  assign new_n1521 = ~new_n1484 & new_n1494;
  assign new_n1522 = ~new_n1483 & ~new_n1521;
  assign new_n1523 = ~new_n1520 & ~new_n1522;
  assign new_n1524 = new_n1520 & new_n1522;
  assign new_n1525 = ~new_n1523 & ~new_n1524;
  assign new_n1526 = new_n1498 & new_n1525;
  assign new_n1527 = n3006 & n9187;
  assign new_n1528 = n8308 & n12306;
  assign new_n1529 = n4748 & n5568;
  assign new_n1530 = ~new_n1528 & ~new_n1529;
  assign new_n1531 = new_n1528 & new_n1529;
  assign new_n1532 = ~new_n1530 & ~new_n1531;
  assign new_n1533 = n4006 & n5214;
  assign new_n1534 = n2758 & n2771;
  assign new_n1535 = n4470 & n6168;
  assign new_n1536 = ~new_n1534 & ~new_n1535;
  assign new_n1537 = new_n1534 & new_n1535;
  assign new_n1538 = ~new_n1536 & ~new_n1537;
  assign new_n1539 = ~new_n1533 & ~new_n1538;
  assign new_n1540 = new_n1533 & new_n1538;
  assign new_n1541 = ~new_n1539 & ~new_n1540;
  assign new_n1542 = ~new_n1506 & ~new_n1510;
  assign new_n1543 = ~new_n1509 & ~new_n1542;
  assign new_n1544 = ~new_n1541 & ~new_n1543;
  assign new_n1545 = new_n1541 & new_n1543;
  assign new_n1546 = ~new_n1544 & ~new_n1545;
  assign new_n1547 = ~new_n1532 & ~new_n1546;
  assign new_n1548 = new_n1532 & new_n1546;
  assign new_n1549 = ~new_n1547 & ~new_n1548;
  assign new_n1550 = ~new_n1504 & new_n1514;
  assign new_n1551 = ~new_n1503 & ~new_n1550;
  assign new_n1552 = ~new_n1549 & ~new_n1551;
  assign new_n1553 = new_n1549 & new_n1551;
  assign new_n1554 = ~new_n1552 & ~new_n1553;
  assign new_n1555 = ~new_n1518 & new_n1522;
  assign new_n1556 = ~new_n1519 & ~new_n1555;
  assign new_n1557 = new_n1554 & ~new_n1556;
  assign new_n1558 = ~new_n1554 & new_n1556;
  assign new_n1559 = ~new_n1557 & ~new_n1558;
  assign new_n1560 = new_n1527 & new_n1559;
  assign new_n1561_1 = ~new_n1527 & ~new_n1559;
  assign new_n1562 = ~new_n1560 & ~new_n1561_1;
  assign new_n1563 = new_n1526 & new_n1562;
  assign new_n1564 = ~new_n1526 & ~new_n1562;
  assign new_n1565 = ~new_n1563 & ~new_n1564;
  assign new_n1566 = n5801 & n10606;
  assign new_n1567 = n10408 & n10908;
  assign new_n1568 = new_n1566 & new_n1567;
  assign new_n1569 = n10408 & n10560;
  assign new_n1570 = n10606 & n10908;
  assign new_n1571 = n5801 & n12965;
  assign new_n1572 = ~new_n1570 & ~new_n1571;
  assign new_n1573 = new_n1570 & new_n1571;
  assign new_n1574 = ~new_n1572 & ~new_n1573;
  assign new_n1575 = new_n1569 & ~new_n1574;
  assign new_n1576 = ~new_n1569 & new_n1574;
  assign new_n1577 = ~new_n1575 & ~new_n1576;
  assign new_n1578 = new_n1568 & ~new_n1577;
  assign new_n1579 = n1724 & n5801;
  assign new_n1580 = new_n1569 & ~new_n1572;
  assign new_n1581 = ~new_n1573 & ~new_n1580;
  assign new_n1582 = ~new_n1579 & new_n1581;
  assign new_n1583 = new_n1579 & ~new_n1581;
  assign new_n1584 = ~new_n1582 & ~new_n1583;
  assign new_n1585 = n10408 & n12003;
  assign new_n1586 = n10908 & n12965;
  assign new_n1587 = n10560 & n10606;
  assign new_n1588 = ~new_n1586 & ~new_n1587;
  assign new_n1589 = new_n1586 & new_n1587;
  assign new_n1590 = ~new_n1588 & ~new_n1589;
  assign new_n1591 = new_n1585 & ~new_n1590;
  assign new_n1592 = ~new_n1585 & new_n1590;
  assign new_n1593 = ~new_n1591 & ~new_n1592;
  assign new_n1594 = ~new_n1584 & new_n1593;
  assign new_n1595 = new_n1584 & ~new_n1593;
  assign new_n1596 = ~new_n1594 & ~new_n1595;
  assign new_n1597 = new_n1578 & new_n1596;
  assign new_n1598 = n5801 & n6937;
  assign new_n1599 = n1724 & n10908;
  assign new_n1600 = new_n1585 & ~new_n1588;
  assign new_n1601 = ~new_n1589 & ~new_n1600;
  assign new_n1602 = ~new_n1599 & new_n1601;
  assign new_n1603 = new_n1599 & ~new_n1601;
  assign new_n1604 = ~new_n1602 & ~new_n1603;
  assign new_n1605 = n8139 & n10408;
  assign new_n1606 = n10560 & n12965;
  assign new_n1607 = n10606 & n12003;
  assign new_n1608 = ~new_n1606 & ~new_n1607;
  assign new_n1609 = new_n1606 & new_n1607;
  assign new_n1610 = ~new_n1608 & ~new_n1609;
  assign new_n1611 = new_n1605 & ~new_n1610;
  assign new_n1612 = ~new_n1605 & new_n1610;
  assign new_n1613 = ~new_n1611 & ~new_n1612;
  assign new_n1614 = ~new_n1604 & new_n1613;
  assign new_n1615 = new_n1604 & ~new_n1613;
  assign new_n1616 = ~new_n1614 & ~new_n1615;
  assign new_n1617 = ~new_n1598 & ~new_n1616;
  assign new_n1618 = new_n1598 & new_n1616;
  assign new_n1619 = ~new_n1617 & ~new_n1618;
  assign new_n1620 = ~new_n1582 & ~new_n1593;
  assign new_n1621 = ~new_n1583 & ~new_n1620;
  assign new_n1622 = ~new_n1619 & new_n1621;
  assign new_n1623 = new_n1619 & ~new_n1621;
  assign new_n1624 = ~new_n1622 & ~new_n1623;
  assign new_n1625 = new_n1597 & new_n1624;
  assign new_n1626 = n3677 & n5801;
  assign new_n1627 = ~new_n1618 & new_n1621;
  assign new_n1628 = ~new_n1617 & ~new_n1627;
  assign new_n1629 = n6937 & n10908;
  assign new_n1630 = n1724 & n10560;
  assign new_n1631 = ~new_n1629 & ~new_n1630;
  assign new_n1632 = new_n1629 & new_n1630;
  assign new_n1633 = ~new_n1631 & ~new_n1632;
  assign new_n1634 = n12003 & n12965;
  assign new_n1635 = n8139 & n10606;
  assign new_n1636_1 = n3311 & n10408;
  assign new_n1637 = ~new_n1635 & ~new_n1636_1;
  assign new_n1638 = new_n1635 & new_n1636_1;
  assign new_n1639 = ~new_n1637 & ~new_n1638;
  assign new_n1640 = ~new_n1634 & ~new_n1639;
  assign new_n1641 = new_n1634 & new_n1639;
  assign new_n1642 = ~new_n1640 & ~new_n1641;
  assign new_n1643 = new_n1605 & ~new_n1608;
  assign new_n1644 = ~new_n1609 & ~new_n1643;
  assign new_n1645 = ~new_n1642 & ~new_n1644;
  assign new_n1646 = new_n1642 & new_n1644;
  assign new_n1647 = ~new_n1645 & ~new_n1646;
  assign new_n1648 = ~new_n1633 & new_n1647;
  assign new_n1649 = new_n1633 & ~new_n1647;
  assign new_n1650_1 = ~new_n1648 & ~new_n1649;
  assign new_n1651 = ~new_n1603 & new_n1613;
  assign new_n1652 = ~new_n1602 & ~new_n1651;
  assign new_n1653 = ~new_n1650_1 & ~new_n1652;
  assign new_n1654 = new_n1650_1 & new_n1652;
  assign new_n1655 = ~new_n1653 & ~new_n1654;
  assign new_n1656 = new_n1628 & new_n1655;
  assign new_n1657 = ~new_n1628 & ~new_n1655;
  assign new_n1658 = ~new_n1656 & ~new_n1657;
  assign new_n1659 = new_n1626 & new_n1658;
  assign new_n1660 = ~new_n1626 & ~new_n1658;
  assign new_n1661 = ~new_n1659 & ~new_n1660;
  assign new_n1662 = ~new_n1625 & ~new_n1661;
  assign new_n1663 = new_n1625 & new_n1661;
  assign new_n1664 = ~new_n1662 & ~new_n1663;
  assign new_n1665 = ~new_n1597 & ~new_n1624;
  assign new_n1666 = ~new_n1625 & ~new_n1665;
  assign new_n1667 = n4335 & n5671;
  assign new_n1668 = n4114 & n8233;
  assign new_n1669 = new_n1667 & new_n1668;
  assign new_n1670 = n8233 & n11665;
  assign new_n1671 = n4114 & n4335;
  assign new_n1672 = n5671 & n9887;
  assign new_n1673 = ~new_n1671 & ~new_n1672;
  assign new_n1674 = new_n1671 & new_n1672;
  assign new_n1675 = ~new_n1673 & ~new_n1674;
  assign new_n1676 = new_n1670 & ~new_n1675;
  assign new_n1677 = ~new_n1670 & new_n1675;
  assign new_n1678 = ~new_n1676 & ~new_n1677;
  assign new_n1679 = new_n1669 & ~new_n1678;
  assign new_n1680 = n497 & n5671;
  assign new_n1681 = new_n1670 & ~new_n1673;
  assign new_n1682 = ~new_n1674 & ~new_n1681;
  assign new_n1683 = ~new_n1680 & new_n1682;
  assign new_n1684 = new_n1680 & ~new_n1682;
  assign new_n1685 = ~new_n1683 & ~new_n1684;
  assign new_n1686 = n2777 & n8233;
  assign new_n1687 = n4114 & n9887;
  assign new_n1688 = n4335 & n11665;
  assign new_n1689 = ~new_n1687 & ~new_n1688;
  assign new_n1690 = new_n1687 & new_n1688;
  assign new_n1691 = ~new_n1689 & ~new_n1690;
  assign new_n1692 = new_n1686 & ~new_n1691;
  assign new_n1693 = ~new_n1686 & new_n1691;
  assign new_n1694 = ~new_n1692 & ~new_n1693;
  assign new_n1695 = ~new_n1685 & new_n1694;
  assign new_n1696 = new_n1685 & ~new_n1694;
  assign new_n1697 = ~new_n1695 & ~new_n1696;
  assign new_n1698 = new_n1679 & new_n1697;
  assign new_n1699 = n2174 & n5671;
  assign new_n1700 = n497 & n4114;
  assign new_n1701 = new_n1686 & ~new_n1689;
  assign new_n1702 = ~new_n1690 & ~new_n1701;
  assign new_n1703 = ~new_n1700 & new_n1702;
  assign new_n1704 = new_n1700 & ~new_n1702;
  assign new_n1705 = ~new_n1703 & ~new_n1704;
  assign new_n1706 = n8233 & n10642;
  assign new_n1707 = n9887 & n11665;
  assign new_n1708 = n2777 & n4335;
  assign new_n1709_1 = ~new_n1707 & ~new_n1708;
  assign new_n1710 = new_n1707 & new_n1708;
  assign new_n1711 = ~new_n1709_1 & ~new_n1710;
  assign new_n1712 = new_n1706 & ~new_n1711;
  assign new_n1713 = ~new_n1706 & new_n1711;
  assign new_n1714 = ~new_n1712 & ~new_n1713;
  assign new_n1715 = ~new_n1705 & new_n1714;
  assign new_n1716 = new_n1705 & ~new_n1714;
  assign new_n1717 = ~new_n1715 & ~new_n1716;
  assign new_n1718 = ~new_n1699 & ~new_n1717;
  assign new_n1719 = new_n1699 & new_n1717;
  assign new_n1720 = ~new_n1718 & ~new_n1719;
  assign new_n1721 = ~new_n1683 & ~new_n1694;
  assign new_n1722 = ~new_n1684 & ~new_n1721;
  assign new_n1723 = ~new_n1720 & new_n1722;
  assign new_n1724_1 = new_n1720 & ~new_n1722;
  assign new_n1725 = ~new_n1723 & ~new_n1724_1;
  assign new_n1726 = ~new_n1698 & ~new_n1725;
  assign new_n1727 = new_n1698 & new_n1725;
  assign new_n1728 = ~new_n1726 & ~new_n1727;
  assign new_n1729 = n9915 & n13201;
  assign new_n1730 = n2057 & n10063;
  assign new_n1731 = new_n1729 & new_n1730;
  assign new_n1732 = n5586 & n10063;
  assign new_n1733 = n2057 & n9915;
  assign new_n1734 = n8332 & n13201;
  assign new_n1735 = ~new_n1733 & ~new_n1734;
  assign new_n1736 = new_n1733 & new_n1734;
  assign new_n1737 = ~new_n1735 & ~new_n1736;
  assign new_n1738 = new_n1732 & ~new_n1737;
  assign new_n1739 = ~new_n1732 & new_n1737;
  assign new_n1740 = ~new_n1738 & ~new_n1739;
  assign new_n1741 = new_n1731 & ~new_n1740;
  assign new_n1742 = n3832 & n13201;
  assign new_n1743 = new_n1732 & ~new_n1735;
  assign new_n1744 = ~new_n1736 & ~new_n1743;
  assign new_n1745 = ~new_n1742 & new_n1744;
  assign new_n1746 = new_n1742 & ~new_n1744;
  assign new_n1747 = ~new_n1745 & ~new_n1746;
  assign new_n1748 = n4141 & n10063;
  assign new_n1749 = n2057 & n8332;
  assign new_n1750 = n5586 & n9915;
  assign new_n1751 = ~new_n1749 & ~new_n1750;
  assign new_n1752 = new_n1749 & new_n1750;
  assign new_n1753 = ~new_n1751 & ~new_n1752;
  assign new_n1754 = new_n1748 & ~new_n1753;
  assign new_n1755 = ~new_n1748 & new_n1753;
  assign new_n1756 = ~new_n1754 & ~new_n1755;
  assign new_n1757_1 = ~new_n1747 & new_n1756;
  assign new_n1758 = new_n1747 & ~new_n1756;
  assign new_n1759 = ~new_n1757_1 & ~new_n1758;
  assign new_n1760 = new_n1741 & new_n1759;
  assign new_n1761 = n2882 & n13201;
  assign new_n1762 = n2057 & n3832;
  assign new_n1763 = new_n1748 & ~new_n1751;
  assign new_n1764 = ~new_n1752 & ~new_n1763;
  assign new_n1765 = ~new_n1762 & new_n1764;
  assign new_n1766 = new_n1762 & ~new_n1764;
  assign new_n1767 = ~new_n1765 & ~new_n1766;
  assign new_n1768 = n1364 & n10063;
  assign new_n1769 = n5586 & n8332;
  assign new_n1770 = n4141 & n9915;
  assign new_n1771 = ~new_n1769 & ~new_n1770;
  assign new_n1772 = new_n1769 & new_n1770;
  assign new_n1773 = ~new_n1771 & ~new_n1772;
  assign new_n1774 = new_n1768 & ~new_n1773;
  assign new_n1775 = ~new_n1768 & new_n1773;
  assign new_n1776 = ~new_n1774 & ~new_n1775;
  assign new_n1777 = ~new_n1767 & new_n1776;
  assign new_n1778 = new_n1767 & ~new_n1776;
  assign new_n1779 = ~new_n1777 & ~new_n1778;
  assign new_n1780 = ~new_n1761 & ~new_n1779;
  assign new_n1781 = new_n1761 & new_n1779;
  assign new_n1782 = ~new_n1780 & ~new_n1781;
  assign new_n1783 = ~new_n1745 & ~new_n1756;
  assign new_n1784 = ~new_n1746 & ~new_n1783;
  assign new_n1785 = ~new_n1782 & new_n1784;
  assign new_n1786 = new_n1782 & ~new_n1784;
  assign new_n1787 = ~new_n1785 & ~new_n1786;
  assign new_n1788 = ~new_n1760 & ~new_n1787;
  assign new_n1789 = new_n1760 & new_n1787;
  assign new_n1790 = ~new_n1788 & ~new_n1789;
  assign new_n1791 = ~new_n1679 & ~new_n1697;
  assign new_n1792 = ~new_n1698 & ~new_n1791;
  assign new_n1793 = ~new_n1741 & ~new_n1759;
  assign new_n1794 = ~new_n1760 & ~new_n1793;
  assign new_n1795 = new_n1792 & new_n1794;
  assign new_n1796 = ~new_n1792 & ~new_n1794;
  assign new_n1797 = ~new_n1669 & new_n1678;
  assign new_n1798 = ~new_n1679 & ~new_n1797;
  assign new_n1799 = ~new_n1731 & new_n1740;
  assign new_n1800 = ~new_n1741 & ~new_n1799;
  assign new_n1801 = new_n1798 & new_n1800;
  assign new_n1802 = ~new_n1798 & ~new_n1800;
  assign new_n1803 = n5671 & n8233;
  assign new_n1804 = n10063 & n13201;
  assign new_n1805 = new_n1803 & new_n1804;
  assign new_n1806_1 = ~new_n1729 & ~new_n1730;
  assign new_n1807 = ~new_n1731 & ~new_n1806_1;
  assign new_n1808 = new_n1805 & new_n1807;
  assign new_n1809 = ~new_n1805 & ~new_n1807;
  assign new_n1810 = ~new_n1667 & ~new_n1668;
  assign new_n1811 = ~new_n1669 & ~new_n1810;
  assign new_n1812 = ~new_n1809 & new_n1811;
  assign new_n1813 = ~new_n1808 & ~new_n1812;
  assign new_n1814 = ~new_n1802 & ~new_n1813;
  assign new_n1815 = ~new_n1801 & ~new_n1814;
  assign new_n1816 = ~new_n1796 & ~new_n1815;
  assign new_n1817 = ~new_n1795 & ~new_n1816;
  assign new_n1818 = new_n1790 & ~new_n1817;
  assign new_n1819 = ~new_n1790 & new_n1817;
  assign new_n1820 = ~new_n1818 & ~new_n1819;
  assign new_n1821 = ~new_n1728 & new_n1820;
  assign new_n1822 = new_n1728 & ~new_n1820;
  assign new_n1823 = ~new_n1821 & ~new_n1822;
  assign new_n1824 = ~new_n1666 & new_n1823;
  assign new_n1825 = new_n1666 & ~new_n1823;
  assign new_n1826 = ~new_n1578 & ~new_n1596;
  assign new_n1827 = ~new_n1597 & ~new_n1826;
  assign new_n1828 = ~new_n1795 & ~new_n1796;
  assign new_n1829 = new_n1815 & ~new_n1828;
  assign new_n1830 = ~new_n1815 & new_n1828;
  assign new_n1831 = ~new_n1829 & ~new_n1830;
  assign new_n1832 = ~new_n1827 & ~new_n1831;
  assign new_n1833 = new_n1827 & new_n1831;
  assign new_n1834 = ~new_n1568 & new_n1577;
  assign new_n1835 = ~new_n1578 & ~new_n1834;
  assign new_n1836 = ~new_n1801 & ~new_n1802;
  assign new_n1837 = new_n1813 & ~new_n1836;
  assign new_n1838 = ~new_n1813 & new_n1836;
  assign new_n1839 = ~new_n1837 & ~new_n1838;
  assign new_n1840 = ~new_n1835 & ~new_n1839;
  assign new_n1841 = new_n1835 & new_n1839;
  assign new_n1842 = ~new_n1566 & ~new_n1567;
  assign new_n1843 = ~new_n1568 & ~new_n1842;
  assign new_n1844 = ~new_n1808 & ~new_n1809;
  assign new_n1845 = new_n1811 & ~new_n1844;
  assign new_n1846 = ~new_n1811 & new_n1844;
  assign new_n1847 = ~new_n1845 & ~new_n1846;
  assign new_n1848 = ~new_n1843 & new_n1847;
  assign new_n1849 = new_n1843 & ~new_n1847;
  assign new_n1850 = n5801 & n10408;
  assign new_n1851 = ~new_n1803 & ~new_n1804;
  assign new_n1852 = ~new_n1805 & ~new_n1851;
  assign new_n1853 = new_n1850 & new_n1852;
  assign new_n1854 = ~new_n1849 & ~new_n1853;
  assign new_n1855 = ~new_n1848 & ~new_n1854;
  assign new_n1856 = ~new_n1841 & ~new_n1855;
  assign new_n1857 = ~new_n1840 & ~new_n1856;
  assign new_n1858 = ~new_n1833 & ~new_n1857;
  assign new_n1859 = ~new_n1832 & ~new_n1858;
  assign new_n1860_1 = ~new_n1825 & ~new_n1859;
  assign new_n1861 = ~new_n1824 & ~new_n1860_1;
  assign new_n1862 = ~new_n1664 & ~new_n1861;
  assign new_n1863 = n4357 & n13201;
  assign new_n1864 = n2057 & n2882;
  assign new_n1865 = n3832 & n5586;
  assign new_n1866 = ~new_n1864 & ~new_n1865;
  assign new_n1867 = new_n1864 & new_n1865;
  assign new_n1868 = ~new_n1866 & ~new_n1867;
  assign new_n1869 = n4141 & n8332;
  assign new_n1870 = n3669 & n10063;
  assign new_n1871 = n1364 & n9915;
  assign new_n1872 = ~new_n1870 & ~new_n1871;
  assign new_n1873 = new_n1870 & new_n1871;
  assign new_n1874 = ~new_n1872 & ~new_n1873;
  assign new_n1875 = new_n1869 & new_n1874;
  assign new_n1876 = ~new_n1869 & ~new_n1874;
  assign new_n1877 = ~new_n1875 & ~new_n1876;
  assign new_n1878 = new_n1768 & ~new_n1771;
  assign new_n1879 = ~new_n1772 & ~new_n1878;
  assign new_n1880 = ~new_n1877 & new_n1879;
  assign new_n1881 = new_n1877 & ~new_n1879;
  assign new_n1882 = ~new_n1880 & ~new_n1881;
  assign new_n1883 = ~new_n1868 & ~new_n1882;
  assign new_n1884 = new_n1868 & new_n1882;
  assign new_n1885 = ~new_n1883 & ~new_n1884;
  assign new_n1886 = ~new_n1765 & ~new_n1776;
  assign new_n1887 = ~new_n1766 & ~new_n1886;
  assign new_n1888 = ~new_n1885 & ~new_n1887;
  assign new_n1889 = new_n1885 & new_n1887;
  assign new_n1890 = ~new_n1888 & ~new_n1889;
  assign new_n1891 = ~new_n1780 & ~new_n1784;
  assign new_n1892 = ~new_n1781 & ~new_n1891;
  assign new_n1893 = ~new_n1890 & ~new_n1892;
  assign new_n1894 = new_n1890 & new_n1892;
  assign new_n1895 = ~new_n1893 & ~new_n1894;
  assign new_n1896 = new_n1863 & new_n1895;
  assign new_n1897 = ~new_n1863 & ~new_n1895;
  assign new_n1898 = ~new_n1896 & ~new_n1897;
  assign new_n1899 = ~new_n1789 & ~new_n1898;
  assign new_n1900 = new_n1789 & new_n1898;
  assign new_n1901 = ~new_n1899 & ~new_n1900;
  assign new_n1902 = n3112 & n5671;
  assign new_n1903 = ~new_n1719 & new_n1722;
  assign new_n1904 = ~new_n1718 & ~new_n1903;
  assign new_n1905 = n2174 & n4114;
  assign new_n1906 = n497 & n11665;
  assign new_n1907 = ~new_n1905 & ~new_n1906;
  assign new_n1908 = new_n1905 & new_n1906;
  assign new_n1909 = ~new_n1907 & ~new_n1908;
  assign new_n1910 = n2777 & n9887;
  assign new_n1911 = n4335 & n10642;
  assign new_n1912_1 = n937 & n8233;
  assign new_n1913 = ~new_n1911 & ~new_n1912_1;
  assign new_n1914 = new_n1911 & new_n1912_1;
  assign new_n1915 = ~new_n1913 & ~new_n1914;
  assign new_n1916_1 = new_n1910 & new_n1915;
  assign new_n1917 = ~new_n1910 & ~new_n1915;
  assign new_n1918 = ~new_n1916_1 & ~new_n1917;
  assign new_n1919 = new_n1706 & ~new_n1709_1;
  assign new_n1920 = ~new_n1710 & ~new_n1919;
  assign new_n1921 = ~new_n1918 & new_n1920;
  assign new_n1922 = new_n1918 & ~new_n1920;
  assign new_n1923 = ~new_n1921 & ~new_n1922;
  assign new_n1924 = ~new_n1909 & ~new_n1923;
  assign new_n1925 = new_n1909 & new_n1923;
  assign new_n1926 = ~new_n1924 & ~new_n1925;
  assign new_n1927 = ~new_n1703 & ~new_n1714;
  assign new_n1928 = ~new_n1704 & ~new_n1927;
  assign new_n1929 = ~new_n1926 & ~new_n1928;
  assign new_n1930 = new_n1926 & new_n1928;
  assign new_n1931 = ~new_n1929 & ~new_n1930;
  assign new_n1932 = new_n1904 & ~new_n1931;
  assign new_n1933 = ~new_n1904 & new_n1931;
  assign new_n1934 = ~new_n1932 & ~new_n1933;
  assign new_n1935 = new_n1902 & new_n1934;
  assign new_n1936 = ~new_n1902 & ~new_n1934;
  assign new_n1937_1 = ~new_n1935 & ~new_n1936;
  assign new_n1938 = ~new_n1727 & ~new_n1937_1;
  assign new_n1939 = new_n1727 & new_n1937_1;
  assign new_n1940 = ~new_n1938 & ~new_n1939;
  assign new_n1941 = new_n1901 & new_n1940;
  assign new_n1942 = ~new_n1901 & ~new_n1940;
  assign new_n1943 = ~new_n1941 & ~new_n1942;
  assign new_n1944 = new_n1728 & ~new_n1819;
  assign new_n1945 = ~new_n1818 & ~new_n1944;
  assign new_n1946 = ~new_n1943 & ~new_n1945;
  assign new_n1947 = new_n1943 & new_n1945;
  assign new_n1948 = ~new_n1946 & ~new_n1947;
  assign new_n1949 = new_n1862 & new_n1948;
  assign new_n1950 = new_n1664 & new_n1861;
  assign new_n1951 = ~new_n1948 & new_n1950;
  assign new_n1952 = ~new_n1862 & ~new_n1948;
  assign new_n1953 = ~new_n1950 & ~new_n1952;
  assign new_n1954 = ~new_n1951 & ~new_n1953;
  assign new_n1955 = ~new_n1949 & ~new_n1954;
  assign new_n1956 = ~new_n1565 & ~new_n1955;
  assign new_n1957 = new_n1565 & new_n1955;
  assign new_n1958 = ~new_n1956 & ~new_n1957;
  assign new_n1959 = ~new_n1498 & ~new_n1525;
  assign new_n1960 = ~new_n1526 & ~new_n1959;
  assign new_n1961 = ~new_n1824 & ~new_n1825;
  assign new_n1962 = ~new_n1859 & ~new_n1961;
  assign new_n1963 = new_n1859 & new_n1961;
  assign new_n1964 = ~new_n1962 & ~new_n1963;
  assign new_n1965 = new_n1960 & new_n1964;
  assign new_n1966 = ~new_n1960 & ~new_n1964;
  assign new_n1967 = ~new_n1479 & ~new_n1497;
  assign new_n1968 = ~new_n1498 & ~new_n1967;
  assign new_n1969 = ~new_n1832 & ~new_n1833;
  assign new_n1970 = ~new_n1857 & ~new_n1969;
  assign new_n1971 = new_n1857 & new_n1969;
  assign new_n1972 = ~new_n1970 & ~new_n1971;
  assign new_n1973 = new_n1968 & new_n1972;
  assign new_n1974 = ~new_n1968 & ~new_n1972;
  assign new_n1975 = ~new_n1469 & new_n1478;
  assign new_n1976 = ~new_n1479 & ~new_n1975;
  assign new_n1977 = ~new_n1840 & ~new_n1841;
  assign new_n1978 = new_n1855 & ~new_n1977;
  assign new_n1979 = ~new_n1855 & new_n1977;
  assign new_n1980 = ~new_n1978 & ~new_n1979;
  assign new_n1981 = new_n1976 & ~new_n1980;
  assign new_n1982_1 = ~new_n1976 & new_n1980;
  assign new_n1983 = ~new_n1467 & ~new_n1468;
  assign new_n1984 = ~new_n1469 & ~new_n1983;
  assign new_n1985 = n3006 & n4470;
  assign new_n1986 = ~new_n1850 & ~new_n1852;
  assign new_n1987 = ~new_n1853 & ~new_n1986;
  assign new_n1988 = new_n1985 & new_n1987;
  assign new_n1989 = ~new_n1984 & ~new_n1988;
  assign new_n1990 = new_n1984 & new_n1988;
  assign new_n1991 = ~new_n1848 & ~new_n1849;
  assign new_n1992 = ~new_n1853 & new_n1991;
  assign new_n1993 = new_n1853 & ~new_n1991;
  assign new_n1994 = ~new_n1992 & ~new_n1993;
  assign new_n1995 = ~new_n1990 & new_n1994;
  assign new_n1996 = ~new_n1989 & ~new_n1995;
  assign new_n1997 = ~new_n1982_1 & new_n1996;
  assign new_n1998 = ~new_n1981 & ~new_n1997;
  assign new_n1999 = ~new_n1974 & ~new_n1998;
  assign new_n2000 = ~new_n1973 & ~new_n1999;
  assign new_n2001 = ~new_n1966 & ~new_n2000;
  assign new_n2002 = ~new_n1965 & ~new_n2001;
  assign new_n2003 = ~new_n1958 & new_n2002;
  assign new_n2004 = new_n1958 & ~new_n2002;
  assign n358 = ~new_n2003 & ~new_n2004;
  assign new_n2006 = n2482 & n6655;
  assign new_n2007 = n1757 & n9669;
  assign new_n2008 = n9528 & n10113;
  assign new_n2009 = ~new_n2007 & ~new_n2008;
  assign new_n2010 = new_n2007 & new_n2008;
  assign new_n2011 = ~new_n2009 & ~new_n2010;
  assign new_n2012 = n10416 & n11891;
  assign new_n2013 = n11488 & n12853;
  assign new_n2014 = n9531 & n11030;
  assign new_n2015 = ~new_n2013 & ~new_n2014;
  assign new_n2016 = new_n2013 & new_n2014;
  assign new_n2017 = ~new_n2015 & ~new_n2016;
  assign new_n2018 = ~new_n2012 & ~new_n2017;
  assign new_n2019 = new_n2012 & new_n2017;
  assign new_n2020 = ~new_n2018 & ~new_n2019;
  assign new_n2021 = n9531 & n10416;
  assign new_n2022 = n1757 & n11891;
  assign new_n2023 = new_n2021 & new_n2022;
  assign new_n2024 = ~new_n2021 & ~new_n2022;
  assign new_n2025 = n11030 & n12853;
  assign new_n2026 = ~new_n2024 & new_n2025;
  assign new_n2027 = ~new_n2023 & ~new_n2026;
  assign new_n2028 = ~new_n2020 & ~new_n2027;
  assign new_n2029 = new_n2020 & new_n2027;
  assign new_n2030 = ~new_n2028 & ~new_n2029;
  assign new_n2031 = new_n2011 & ~new_n2030;
  assign new_n2032 = ~new_n2011 & new_n2030;
  assign new_n2033 = ~new_n2031 & ~new_n2032;
  assign new_n2034 = n9669 & n10113;
  assign new_n2035 = n1757 & n9531;
  assign new_n2036 = n10113 & n11891;
  assign new_n2037 = new_n2035 & new_n2036;
  assign new_n2038 = ~new_n2035 & ~new_n2036;
  assign new_n2039 = n10416 & n12853;
  assign new_n2040 = ~new_n2038 & new_n2039;
  assign new_n2041 = ~new_n2037 & ~new_n2040;
  assign new_n2042 = ~new_n2034 & new_n2041;
  assign new_n2043 = new_n2034 & ~new_n2041;
  assign new_n2044 = ~new_n2023 & ~new_n2024;
  assign new_n2045 = ~new_n2025 & ~new_n2044;
  assign new_n2046 = new_n2025 & new_n2044;
  assign new_n2047 = ~new_n2045 & ~new_n2046;
  assign new_n2048 = ~new_n2043 & ~new_n2047;
  assign new_n2049 = ~new_n2042 & ~new_n2048;
  assign new_n2050 = ~new_n2033 & new_n2049;
  assign new_n2051 = new_n2033 & ~new_n2049;
  assign new_n2052 = ~new_n2050 & ~new_n2051;
  assign new_n2053 = n2482 & n9528;
  assign new_n2054 = ~new_n2042 & ~new_n2043;
  assign new_n2055 = new_n2047 & ~new_n2054;
  assign new_n2056 = ~new_n2047 & new_n2054;
  assign new_n2057_1 = ~new_n2055 & ~new_n2056;
  assign new_n2058 = new_n2053 & ~new_n2057_1;
  assign new_n2059 = ~new_n2053 & new_n2057_1;
  assign new_n2060 = n2482 & n9669;
  assign new_n2061_1 = n9531 & n10113;
  assign new_n2062 = n2482 & n11891;
  assign new_n2063 = new_n2061_1 & new_n2062;
  assign new_n2064 = ~new_n2061_1 & ~new_n2062;
  assign new_n2065 = n1757 & n12853;
  assign new_n2066 = ~new_n2064 & new_n2065;
  assign new_n2067 = ~new_n2063 & ~new_n2066;
  assign new_n2068_1 = ~new_n2060 & new_n2067;
  assign new_n2069 = new_n2060 & ~new_n2067;
  assign new_n2070 = ~new_n2037 & ~new_n2038;
  assign new_n2071 = ~new_n2039 & ~new_n2070;
  assign new_n2072 = new_n2039 & new_n2070;
  assign new_n2073 = ~new_n2071 & ~new_n2072;
  assign new_n2074 = ~new_n2069 & ~new_n2073;
  assign new_n2075 = ~new_n2068_1 & ~new_n2074;
  assign new_n2076 = ~new_n2059 & new_n2075;
  assign new_n2077 = ~new_n2058 & ~new_n2076;
  assign new_n2078 = ~new_n2052 & ~new_n2077;
  assign new_n2079 = new_n2052 & new_n2077;
  assign new_n2080 = ~new_n2078 & ~new_n2079;
  assign new_n2081 = new_n2006 & new_n2080;
  assign new_n2082 = n2482 & n9531;
  assign new_n2083 = n10113 & n12853;
  assign new_n2084 = new_n2082 & new_n2083;
  assign new_n2085 = ~new_n2063 & ~new_n2064;
  assign new_n2086 = ~new_n2065 & ~new_n2085;
  assign new_n2087 = new_n2065 & new_n2085;
  assign new_n2088 = ~new_n2086 & ~new_n2087;
  assign new_n2089 = new_n2084 & new_n2088;
  assign new_n2090 = ~new_n2068_1 & ~new_n2069;
  assign new_n2091 = ~new_n2073 & ~new_n2090;
  assign new_n2092 = new_n2073 & new_n2090;
  assign new_n2093 = ~new_n2091 & ~new_n2092;
  assign new_n2094 = new_n2089 & new_n2093;
  assign new_n2095 = ~new_n2058 & ~new_n2059;
  assign new_n2096 = ~new_n2075 & ~new_n2095;
  assign new_n2097 = new_n2075 & new_n2095;
  assign new_n2098 = ~new_n2096 & ~new_n2097;
  assign new_n2099 = new_n2094 & new_n2098;
  assign new_n2100 = ~new_n2006 & ~new_n2080;
  assign new_n2101 = ~new_n2081 & ~new_n2100;
  assign new_n2102 = new_n2099 & new_n2101;
  assign new_n2103 = ~new_n2081 & ~new_n2102;
  assign new_n2104 = ~new_n2032 & new_n2049;
  assign new_n2105 = ~new_n2010 & ~new_n2104;
  assign new_n2106 = ~new_n2031 & new_n2105;
  assign new_n2107 = new_n2010 & new_n2104;
  assign new_n2108 = ~new_n2106 & ~new_n2107;
  assign new_n2109 = n1757 & n9528;
  assign new_n2110 = n6655 & n10113;
  assign new_n2111 = n2482 & n8522;
  assign new_n2112 = ~new_n2110 & ~new_n2111;
  assign new_n2113 = new_n2110 & new_n2111;
  assign new_n2114 = ~new_n2112 & ~new_n2113;
  assign new_n2115 = new_n2109 & ~new_n2114;
  assign new_n2116 = ~new_n2109 & new_n2114;
  assign new_n2117 = ~new_n2115 & ~new_n2116;
  assign new_n2118 = ~new_n2019 & new_n2027;
  assign new_n2119 = ~new_n2018 & ~new_n2118;
  assign new_n2120 = ~new_n2117 & new_n2119;
  assign new_n2121 = new_n2117 & ~new_n2119;
  assign new_n2122 = ~new_n2120 & ~new_n2121;
  assign new_n2123 = n9669 & n10416;
  assign new_n2124 = new_n2016 & new_n2123;
  assign new_n2125 = ~new_n2016 & ~new_n2123;
  assign new_n2126 = ~new_n2124 & ~new_n2125;
  assign new_n2127 = n1982 & n12853;
  assign new_n2128 = n9531 & n11488;
  assign new_n2129 = n11030 & n11891;
  assign new_n2130 = ~new_n2128 & ~new_n2129;
  assign new_n2131 = new_n2128 & new_n2129;
  assign new_n2132 = ~new_n2130 & ~new_n2131;
  assign new_n2133 = new_n2127 & ~new_n2132;
  assign new_n2134 = ~new_n2127 & new_n2132;
  assign new_n2135 = ~new_n2133 & ~new_n2134;
  assign new_n2136 = new_n2126 & new_n2135;
  assign new_n2137 = ~new_n2126 & ~new_n2135;
  assign new_n2138 = ~new_n2136 & ~new_n2137;
  assign new_n2139 = ~new_n2122 & ~new_n2138;
  assign new_n2140 = new_n2122 & new_n2138;
  assign new_n2141 = ~new_n2139 & ~new_n2140;
  assign new_n2142 = ~new_n2108 & new_n2141;
  assign new_n2143 = new_n2108 & ~new_n2141;
  assign new_n2144 = ~new_n2142 & ~new_n2143;
  assign new_n2145 = new_n2078 & new_n2144;
  assign new_n2146 = ~new_n2078 & ~new_n2144;
  assign new_n2147 = ~new_n2145 & ~new_n2146;
  assign new_n2148 = ~new_n2103 & new_n2147;
  assign new_n2149 = new_n2103 & ~new_n2147;
  assign new_n2150 = ~new_n2148 & ~new_n2149;
  assign new_n2151 = n854 & n8228;
  assign new_n2152 = n854 & n11236;
  assign new_n2153 = n854 & n3130;
  assign new_n2154 = n854 & n4382;
  assign new_n2155 = ~new_n2153 & ~new_n2154;
  assign new_n2156 = ~new_n2152 & new_n2155;
  assign new_n2157 = n4382 & new_n2153;
  assign new_n2158 = n11236 & new_n2157;
  assign new_n2159 = ~new_n2151 & ~new_n2158;
  assign new_n2160 = ~new_n2156 & ~new_n2159;
  assign new_n2161 = n854 & n9732;
  assign new_n2162 = ~new_n2156 & ~new_n2158;
  assign new_n2163 = ~new_n2161 & ~new_n2162;
  assign new_n2164 = new_n2161 & new_n2162;
  assign new_n2165 = ~new_n2163 & ~new_n2164;
  assign new_n2166 = new_n2160 & new_n2165;
  assign new_n2167 = new_n2155 & ~new_n2161;
  assign new_n2168 = n11236 & ~new_n2167;
  assign new_n2169 = n9732 & new_n2157;
  assign new_n2170 = ~new_n2168 & ~new_n2169;
  assign new_n2171 = new_n2154 & ~new_n2170;
  assign new_n2172 = ~new_n2154 & new_n2170;
  assign new_n2173 = ~new_n2171 & ~new_n2172;
  assign new_n2174_1 = ~new_n2157 & ~new_n2161;
  assign new_n2175 = ~new_n2155 & ~new_n2174_1;
  assign new_n2176 = n103 & n854;
  assign new_n2177 = n9732 & new_n2176;
  assign new_n2178 = ~new_n2161 & ~new_n2176;
  assign new_n2179 = ~new_n2177 & ~new_n2178;
  assign new_n2180 = ~new_n2153 & ~new_n2179;
  assign new_n2181 = n3130 & new_n2179;
  assign new_n2182 = ~new_n2180 & ~new_n2181;
  assign new_n2183 = ~new_n2175 & ~new_n2182;
  assign new_n2184 = new_n2175 & new_n2182;
  assign new_n2185 = ~new_n2183 & ~new_n2184;
  assign new_n2186 = ~new_n2173 & new_n2185;
  assign new_n2187 = new_n2173 & ~new_n2185;
  assign new_n2188 = ~new_n2186 & ~new_n2187;
  assign new_n2189 = new_n2166 & ~new_n2188;
  assign new_n2190_1 = ~new_n2166 & new_n2188;
  assign new_n2191 = ~new_n2189 & ~new_n2190_1;
  assign new_n2192 = new_n2151 & new_n2191;
  assign new_n2193 = ~new_n2160 & ~new_n2165;
  assign new_n2194 = ~new_n2166 & ~new_n2193;
  assign new_n2195 = n8228 & new_n2158;
  assign new_n2196 = new_n2194 & new_n2195;
  assign new_n2197 = ~new_n2151 & ~new_n2191;
  assign new_n2198 = ~new_n2192 & ~new_n2197;
  assign new_n2199 = new_n2196 & new_n2198;
  assign new_n2200 = ~new_n2192 & ~new_n2199;
  assign new_n2201 = ~new_n2171 & ~new_n2185;
  assign new_n2202 = ~new_n2172 & ~new_n2201;
  assign new_n2203 = n11236 & new_n2151;
  assign new_n2204 = ~new_n2151 & ~new_n2152;
  assign new_n2205 = ~new_n2203 & ~new_n2204;
  assign new_n2206 = ~new_n2175 & ~new_n2181;
  assign new_n2207 = ~new_n2180 & ~new_n2206;
  assign new_n2208 = new_n2205 & new_n2207;
  assign new_n2209 = ~new_n2205 & ~new_n2207;
  assign new_n2210 = ~new_n2208 & ~new_n2209;
  assign new_n2211 = ~new_n2153 & ~new_n2177;
  assign new_n2212 = n3130 & new_n2177;
  assign new_n2213 = ~new_n2211 & ~new_n2212;
  assign new_n2214 = ~n5320 & new_n2179;
  assign new_n2215 = n854 & n5320;
  assign new_n2216 = ~new_n2179 & new_n2215;
  assign new_n2217 = ~new_n2214 & ~new_n2216;
  assign new_n2218 = ~new_n2213 & new_n2217;
  assign new_n2219 = new_n2213 & ~new_n2217;
  assign new_n2220 = ~new_n2218 & ~new_n2219;
  assign new_n2221 = new_n2210 & ~new_n2220;
  assign new_n2222 = ~new_n2210 & new_n2220;
  assign new_n2223 = ~new_n2221 & ~new_n2222;
  assign new_n2224 = new_n2202 & ~new_n2223;
  assign new_n2225 = ~new_n2202 & new_n2223;
  assign new_n2226 = ~new_n2224 & ~new_n2225;
  assign new_n2227 = new_n2189 & new_n2226;
  assign new_n2228 = ~new_n2189 & ~new_n2226;
  assign new_n2229 = ~new_n2227 & ~new_n2228;
  assign new_n2230 = ~new_n2200 & new_n2229;
  assign new_n2231 = new_n2200 & ~new_n2229;
  assign new_n2232 = ~new_n2230 & ~new_n2231;
  assign new_n2233 = n1912 & n13060;
  assign new_n2234 = n2295 & n6333;
  assign new_n2235_1 = ~new_n2233 & ~new_n2234;
  assign new_n2236 = new_n2233 & new_n2234;
  assign new_n2237 = ~new_n2235_1 & ~new_n2236;
  assign new_n2238 = n5189 & n12750;
  assign new_n2239 = n761 & n834;
  assign new_n2240 = n8716 & n9620;
  assign new_n2241 = ~new_n2239 & ~new_n2240;
  assign new_n2242 = new_n2239 & new_n2240;
  assign new_n2243 = ~new_n2241 & ~new_n2242;
  assign new_n2244 = ~new_n2238 & ~new_n2243;
  assign new_n2245 = new_n2238 & new_n2243;
  assign new_n2246 = ~new_n2244 & ~new_n2245;
  assign new_n2247 = n1912 & n5189;
  assign new_n2248 = n8716 & n12750;
  assign new_n2249 = new_n2247 & new_n2248;
  assign new_n2250 = n834 & n9620;
  assign new_n2251 = ~new_n2247 & ~new_n2248;
  assign new_n2252_1 = new_n2250 & ~new_n2251;
  assign new_n2253 = ~new_n2249 & ~new_n2252_1;
  assign new_n2254 = ~new_n2246 & new_n2253;
  assign new_n2255 = new_n2246 & ~new_n2253;
  assign new_n2256 = ~new_n2254 & ~new_n2255;
  assign new_n2257 = ~new_n2237 & ~new_n2256;
  assign new_n2258 = new_n2237 & new_n2256;
  assign new_n2259 = ~new_n2257 & ~new_n2258;
  assign new_n2260 = n6333 & n13060;
  assign new_n2261 = n1912 & n8716;
  assign new_n2262 = n5189 & n6333;
  assign new_n2263 = new_n2261 & new_n2262;
  assign new_n2264 = ~new_n2261 & ~new_n2262;
  assign new_n2265 = n834 & n12750;
  assign new_n2266 = ~new_n2264 & new_n2265;
  assign new_n2267 = ~new_n2263 & ~new_n2266;
  assign new_n2268 = ~new_n2260 & new_n2267;
  assign new_n2269 = new_n2260 & ~new_n2267;
  assign new_n2270 = ~new_n2249 & ~new_n2251;
  assign new_n2271 = new_n2250 & ~new_n2270;
  assign new_n2272 = ~new_n2250 & new_n2270;
  assign new_n2273 = ~new_n2271 & ~new_n2272;
  assign new_n2274 = ~new_n2269 & new_n2273;
  assign new_n2275 = ~new_n2268 & ~new_n2274;
  assign new_n2276 = ~new_n2259 & ~new_n2275;
  assign new_n2277 = new_n2259 & new_n2275;
  assign new_n2278 = ~new_n2276 & ~new_n2277;
  assign new_n2279 = n2295 & n9353;
  assign new_n2280 = ~new_n2268 & ~new_n2269;
  assign new_n2281 = new_n2273 & ~new_n2280;
  assign new_n2282 = ~new_n2273 & new_n2280;
  assign new_n2283 = ~new_n2281 & ~new_n2282;
  assign new_n2284 = new_n2279 & new_n2283;
  assign new_n2285 = ~new_n2279 & ~new_n2283;
  assign new_n2286 = n9353 & n13060;
  assign new_n2287 = n6333 & n8716;
  assign new_n2288 = n5189 & n9353;
  assign new_n2289 = new_n2287 & new_n2288;
  assign new_n2290 = ~new_n2287 & ~new_n2288;
  assign new_n2291 = n834 & n1912;
  assign new_n2292 = ~new_n2290 & new_n2291;
  assign new_n2293 = ~new_n2289 & ~new_n2292;
  assign new_n2294 = ~new_n2286 & new_n2293;
  assign new_n2295_1 = new_n2286 & ~new_n2293;
  assign new_n2296 = ~new_n2263 & ~new_n2264;
  assign new_n2297 = ~new_n2265 & ~new_n2296;
  assign new_n2298 = new_n2265 & new_n2296;
  assign new_n2299 = ~new_n2297 & ~new_n2298;
  assign new_n2300 = ~new_n2295_1 & ~new_n2299;
  assign new_n2301 = ~new_n2294 & ~new_n2300;
  assign new_n2302 = ~new_n2285 & new_n2301;
  assign new_n2303 = ~new_n2284 & ~new_n2302;
  assign new_n2304 = new_n2278 & ~new_n2303;
  assign new_n2305 = ~new_n2257 & new_n2275;
  assign new_n2306 = ~new_n2236 & ~new_n2305;
  assign new_n2307 = ~new_n2258 & new_n2306;
  assign new_n2308 = new_n2236 & new_n2305;
  assign new_n2309 = ~new_n2307 & ~new_n2308;
  assign new_n2310 = n1912 & n2295;
  assign new_n2311 = n1650 & n6333;
  assign new_n2312 = n2341 & n9353;
  assign new_n2313 = ~new_n2311 & ~new_n2312;
  assign new_n2314 = new_n2311 & new_n2312;
  assign new_n2315 = ~new_n2313 & ~new_n2314;
  assign new_n2316 = new_n2310 & ~new_n2315;
  assign new_n2317 = ~new_n2310 & new_n2315;
  assign new_n2318 = ~new_n2316 & ~new_n2317;
  assign new_n2319 = ~new_n2245 & new_n2253;
  assign new_n2320 = ~new_n2244 & ~new_n2319;
  assign new_n2321 = new_n2318 & ~new_n2320;
  assign new_n2322 = n12750 & n13060;
  assign new_n2323 = new_n2242 & new_n2322;
  assign new_n2324 = ~new_n2242 & ~new_n2322;
  assign new_n2325 = ~new_n2323 & ~new_n2324;
  assign new_n2326 = n834 & n5758;
  assign new_n2327 = n761 & n8716;
  assign new_n2328 = n5189 & n9620;
  assign new_n2329 = ~new_n2327 & ~new_n2328;
  assign new_n2330 = new_n2327 & new_n2328;
  assign new_n2331 = ~new_n2329 & ~new_n2330;
  assign new_n2332 = new_n2326 & ~new_n2331;
  assign new_n2333 = ~new_n2326 & new_n2331;
  assign new_n2334 = ~new_n2332 & ~new_n2333;
  assign new_n2335 = new_n2325 & new_n2334;
  assign new_n2336 = ~new_n2325 & ~new_n2334;
  assign new_n2337 = ~new_n2335 & ~new_n2336;
  assign new_n2338 = new_n2321 & new_n2337;
  assign new_n2339_1 = ~new_n2318 & new_n2320;
  assign new_n2340 = new_n2337 & ~new_n2339_1;
  assign new_n2341_1 = ~new_n2321 & ~new_n2340;
  assign new_n2342 = ~new_n2338 & ~new_n2341_1;
  assign new_n2343 = ~new_n2337 & new_n2339_1;
  assign new_n2344 = ~new_n2342 & ~new_n2343;
  assign new_n2345 = ~new_n2309 & new_n2344;
  assign new_n2346 = new_n2309 & ~new_n2344;
  assign new_n2347 = ~new_n2345 & ~new_n2346;
  assign new_n2348 = new_n2304 & new_n2347;
  assign new_n2349 = ~new_n2304 & ~new_n2347;
  assign new_n2350 = ~new_n2348 & ~new_n2349;
  assign new_n2351 = n1650 & n9353;
  assign new_n2352 = ~new_n2278 & new_n2303;
  assign new_n2353 = ~new_n2304 & ~new_n2352;
  assign new_n2354 = new_n2351 & new_n2353;
  assign new_n2355 = n8716 & n9353;
  assign new_n2356 = n834 & n6333;
  assign new_n2357 = new_n2355 & new_n2356;
  assign new_n2358 = ~new_n2289 & ~new_n2290;
  assign new_n2359 = ~new_n2291 & ~new_n2358;
  assign new_n2360 = new_n2291 & new_n2358;
  assign new_n2361 = ~new_n2359 & ~new_n2360;
  assign new_n2362 = new_n2357 & new_n2361;
  assign new_n2363 = ~new_n2294 & ~new_n2295_1;
  assign new_n2364 = ~new_n2299 & new_n2363;
  assign new_n2365 = new_n2299 & ~new_n2363;
  assign new_n2366 = ~new_n2364 & ~new_n2365;
  assign new_n2367 = new_n2362 & ~new_n2366;
  assign new_n2368 = ~new_n2284 & ~new_n2285;
  assign new_n2369 = new_n2301 & new_n2368;
  assign new_n2370 = ~new_n2301 & ~new_n2368;
  assign new_n2371 = ~new_n2369 & ~new_n2370;
  assign new_n2372 = new_n2367 & new_n2371;
  assign new_n2373 = ~new_n2351 & ~new_n2353;
  assign new_n2374 = ~new_n2354 & ~new_n2373;
  assign new_n2375 = new_n2372 & new_n2374;
  assign new_n2376 = ~new_n2354 & ~new_n2375;
  assign new_n2377 = new_n2350 & ~new_n2376;
  assign new_n2378 = ~new_n2350 & new_n2376;
  assign new_n2379 = ~new_n2377 & ~new_n2378;
  assign new_n2380 = n8940 & n12579;
  assign new_n2381 = n4964 & n9591;
  assign new_n2382 = n5684 & n8290;
  assign new_n2383 = new_n2381 & new_n2382;
  assign new_n2384 = ~new_n2381 & ~new_n2382;
  assign new_n2385 = n510 & n10522;
  assign new_n2386 = ~new_n2384 & new_n2385;
  assign new_n2387 = ~new_n2383 & ~new_n2386;
  assign new_n2388 = n510 & n10770;
  assign new_n2389 = n5684 & n9591;
  assign new_n2390 = n8290 & n10522;
  assign new_n2391 = ~new_n2389 & ~new_n2390;
  assign new_n2392 = new_n2389 & new_n2390;
  assign new_n2393 = ~new_n2391 & ~new_n2392;
  assign new_n2394 = new_n2388 & ~new_n2393;
  assign new_n2395 = ~new_n2388 & new_n2393;
  assign new_n2396 = ~new_n2394 & ~new_n2395;
  assign new_n2397 = ~new_n2387 & ~new_n2396;
  assign new_n2398 = n4964 & n11222;
  assign new_n2399 = ~new_n2397 & ~new_n2398;
  assign new_n2400 = new_n2397 & new_n2398;
  assign new_n2401 = ~new_n2399 & ~new_n2400;
  assign new_n2402 = ~new_n2388 & ~new_n2392;
  assign new_n2403 = ~new_n2391 & ~new_n2402;
  assign new_n2404 = n9591 & n10522;
  assign new_n2405 = ~n510 & ~n8290;
  assign new_n2406 = n10770 & ~new_n2405;
  assign new_n2407 = n510 & n8290;
  assign new_n2408 = new_n2406 & ~new_n2407;
  assign new_n2409 = ~new_n2404 & ~new_n2408;
  assign new_n2410 = new_n2404 & new_n2408;
  assign new_n2411 = ~new_n2409 & ~new_n2410;
  assign new_n2412 = new_n2403 & ~new_n2411;
  assign new_n2413 = ~new_n2403 & new_n2411;
  assign new_n2414 = ~new_n2412 & ~new_n2413;
  assign new_n2415 = new_n2401 & new_n2414;
  assign new_n2416 = ~new_n2401 & ~new_n2414;
  assign new_n2417 = ~new_n2415 & ~new_n2416;
  assign new_n2418 = n8940 & n11222;
  assign new_n2419 = ~new_n2383 & ~new_n2384;
  assign new_n2420 = ~new_n2385 & ~new_n2419;
  assign new_n2421 = new_n2385 & new_n2419;
  assign new_n2422 = ~new_n2420 & ~new_n2421;
  assign new_n2423 = n4964 & n8290;
  assign new_n2424 = n8940 & n9591;
  assign new_n2425 = new_n2423 & new_n2424;
  assign new_n2426 = ~new_n2423 & ~new_n2424;
  assign new_n2427 = n510 & n5684;
  assign new_n2428 = ~new_n2426 & new_n2427;
  assign new_n2429 = ~new_n2425 & ~new_n2428;
  assign new_n2430 = new_n2422 & ~new_n2429;
  assign new_n2431 = ~new_n2418 & ~new_n2430;
  assign new_n2432 = new_n2418 & new_n2430;
  assign new_n2433 = new_n2387 & new_n2396;
  assign new_n2434 = ~new_n2397 & ~new_n2433;
  assign new_n2435 = ~new_n2432 & ~new_n2434;
  assign new_n2436 = ~new_n2431 & ~new_n2435;
  assign new_n2437 = ~new_n2417 & new_n2436;
  assign new_n2438 = new_n2417 & ~new_n2436;
  assign new_n2439 = ~new_n2437 & ~new_n2438;
  assign new_n2440 = new_n2380 & new_n2439;
  assign new_n2441 = n8290 & n8940;
  assign new_n2442 = n510 & n4964;
  assign new_n2443 = new_n2441 & new_n2442;
  assign new_n2444 = ~new_n2425 & ~new_n2426;
  assign new_n2445 = ~new_n2427 & ~new_n2444;
  assign new_n2446 = new_n2427 & new_n2444;
  assign new_n2447 = ~new_n2445 & ~new_n2446;
  assign new_n2448 = new_n2443 & new_n2447;
  assign new_n2449 = ~new_n2422 & new_n2429;
  assign new_n2450 = ~new_n2430 & ~new_n2449;
  assign new_n2451 = new_n2448 & new_n2450;
  assign new_n2452 = ~new_n2431 & ~new_n2432;
  assign new_n2453 = new_n2434 & ~new_n2452;
  assign new_n2454 = ~new_n2434 & new_n2452;
  assign new_n2455 = ~new_n2453 & ~new_n2454;
  assign new_n2456 = new_n2451 & ~new_n2455;
  assign new_n2457 = ~new_n2380 & ~new_n2439;
  assign new_n2458_1 = ~new_n2440 & ~new_n2457;
  assign new_n2459 = new_n2456 & new_n2458_1;
  assign new_n2460 = ~new_n2440 & ~new_n2459;
  assign new_n2461 = ~new_n2399 & ~new_n2414;
  assign new_n2462 = ~new_n2400 & ~new_n2461;
  assign new_n2463 = ~new_n2403 & ~new_n2410;
  assign new_n2464 = ~new_n2409 & ~new_n2463;
  assign new_n2465 = n9591 & n10770;
  assign new_n2466 = ~new_n2406 & new_n2465;
  assign new_n2467 = ~n9591 & new_n2406;
  assign new_n2468 = ~new_n2466 & ~new_n2467;
  assign new_n2469 = ~new_n2464 & new_n2468;
  assign new_n2470 = new_n2464 & ~new_n2468;
  assign new_n2471 = ~new_n2469 & ~new_n2470;
  assign new_n2472 = n5684 & n11222;
  assign new_n2473 = n6023 & n8940;
  assign new_n2474 = n4964 & n12579;
  assign new_n2475 = ~new_n2473 & ~new_n2474;
  assign new_n2476 = new_n2473 & new_n2474;
  assign new_n2477 = ~new_n2475 & ~new_n2476;
  assign new_n2478 = new_n2472 & ~new_n2477;
  assign new_n2479 = ~new_n2472 & new_n2477;
  assign new_n2480 = ~new_n2478 & ~new_n2479;
  assign new_n2481 = new_n2471 & ~new_n2480;
  assign new_n2482_1 = ~new_n2471 & new_n2480;
  assign new_n2483 = ~new_n2481 & ~new_n2482_1;
  assign new_n2484 = ~new_n2462 & new_n2483;
  assign new_n2485 = new_n2462 & ~new_n2483;
  assign new_n2486 = ~new_n2484 & ~new_n2485;
  assign new_n2487 = new_n2437 & new_n2486;
  assign new_n2488 = ~new_n2437 & ~new_n2486;
  assign new_n2489 = ~new_n2487 & ~new_n2488;
  assign new_n2490 = ~new_n2460 & new_n2489;
  assign new_n2491 = new_n2460 & ~new_n2489;
  assign new_n2492 = ~new_n2490 & ~new_n2491;
  assign new_n2493 = new_n2379 & new_n2492;
  assign new_n2494 = ~new_n2379 & ~new_n2492;
  assign new_n2495 = ~new_n2493 & ~new_n2494;
  assign new_n2496 = ~new_n2456 & ~new_n2458_1;
  assign new_n2497 = ~new_n2459 & ~new_n2496;
  assign new_n2498_1 = ~new_n2372 & ~new_n2374;
  assign new_n2499 = ~new_n2375 & ~new_n2498_1;
  assign new_n2500 = new_n2497 & new_n2499;
  assign new_n2501 = ~new_n2497 & ~new_n2499;
  assign new_n2502 = ~new_n2367 & ~new_n2371;
  assign new_n2503 = ~new_n2372 & ~new_n2502;
  assign new_n2504 = ~new_n2451 & new_n2455;
  assign new_n2505 = ~new_n2456 & ~new_n2504;
  assign new_n2506 = new_n2503 & new_n2505;
  assign new_n2507 = ~new_n2503 & ~new_n2505;
  assign new_n2508 = ~new_n2448 & ~new_n2450;
  assign new_n2509 = ~new_n2451 & ~new_n2508;
  assign new_n2510 = ~new_n2362 & new_n2366;
  assign new_n2511 = ~new_n2367 & ~new_n2510;
  assign new_n2512 = new_n2509 & new_n2511;
  assign new_n2513 = ~new_n2509 & ~new_n2511;
  assign new_n2514 = ~new_n2357 & ~new_n2361;
  assign new_n2515 = ~new_n2362 & ~new_n2514;
  assign new_n2516 = ~new_n2443 & ~new_n2447;
  assign new_n2517 = ~new_n2448 & ~new_n2516;
  assign new_n2518 = new_n2515 & new_n2517;
  assign new_n2519 = ~new_n2515 & ~new_n2517;
  assign new_n2520 = n834 & n9353;
  assign new_n2521 = n510 & n8940;
  assign new_n2522 = new_n2520 & new_n2521;
  assign new_n2523 = ~new_n2441 & ~new_n2442;
  assign new_n2524 = ~new_n2443 & ~new_n2523;
  assign new_n2525 = new_n2522 & new_n2524;
  assign new_n2526 = ~new_n2522 & ~new_n2524;
  assign new_n2527 = ~new_n2355 & ~new_n2356;
  assign new_n2528 = ~new_n2357 & ~new_n2527;
  assign new_n2529 = ~new_n2526 & new_n2528;
  assign new_n2530 = ~new_n2525 & ~new_n2529;
  assign new_n2531 = ~new_n2519 & ~new_n2530;
  assign new_n2532 = ~new_n2518 & ~new_n2531;
  assign new_n2533 = ~new_n2513 & ~new_n2532;
  assign new_n2534 = ~new_n2512 & ~new_n2533;
  assign new_n2535 = ~new_n2507 & ~new_n2534;
  assign new_n2536 = ~new_n2506 & ~new_n2535;
  assign new_n2537 = ~new_n2501 & ~new_n2536;
  assign new_n2538 = ~new_n2500 & ~new_n2537;
  assign new_n2539 = ~new_n2495 & ~new_n2538;
  assign new_n2540 = new_n2495 & new_n2538;
  assign new_n2541 = ~new_n2539 & ~new_n2540;
  assign new_n2542 = ~new_n2232 & new_n2541;
  assign new_n2543 = new_n2232 & ~new_n2541;
  assign new_n2544 = ~new_n2542 & ~new_n2543;
  assign new_n2545 = ~new_n2196 & ~new_n2198;
  assign new_n2546 = ~new_n2199 & ~new_n2545;
  assign new_n2547 = ~new_n2500 & ~new_n2501;
  assign new_n2548 = new_n2536 & ~new_n2547;
  assign new_n2549_1 = ~new_n2536 & new_n2547;
  assign new_n2550 = ~new_n2548 & ~new_n2549_1;
  assign new_n2551 = ~new_n2546 & ~new_n2550;
  assign new_n2552 = new_n2546 & new_n2550;
  assign new_n2553 = ~new_n2194 & ~new_n2195;
  assign new_n2554 = ~new_n2196 & ~new_n2553;
  assign new_n2555 = ~new_n2506 & ~new_n2507;
  assign new_n2556 = new_n2534 & ~new_n2555;
  assign new_n2557 = ~new_n2534 & new_n2555;
  assign new_n2558 = ~new_n2556 & ~new_n2557;
  assign new_n2559 = ~new_n2554 & ~new_n2558;
  assign new_n2560 = new_n2554 & new_n2558;
  assign new_n2561 = ~new_n2512 & ~new_n2513;
  assign new_n2562 = new_n2532 & ~new_n2561;
  assign new_n2563 = ~new_n2532 & new_n2561;
  assign new_n2564 = ~new_n2562 & ~new_n2563;
  assign new_n2565 = ~new_n2154 & new_n2204;
  assign new_n2566 = ~new_n2153 & ~new_n2565;
  assign new_n2567 = new_n2153 & new_n2565;
  assign new_n2568 = ~new_n2566 & ~new_n2567;
  assign new_n2569 = ~new_n2564 & new_n2568;
  assign new_n2570 = new_n2564 & ~new_n2568;
  assign new_n2571 = n4382 & ~new_n2204;
  assign new_n2572 = ~new_n2565 & ~new_n2571;
  assign new_n2573 = ~new_n2518 & ~new_n2519;
  assign new_n2574 = new_n2530 & ~new_n2573;
  assign new_n2575 = ~new_n2530 & new_n2573;
  assign new_n2576 = ~new_n2574 & ~new_n2575;
  assign new_n2577 = ~new_n2572 & ~new_n2576;
  assign new_n2578 = new_n2572 & new_n2576;
  assign new_n2579 = ~new_n2525 & ~new_n2526;
  assign new_n2580 = new_n2528 & ~new_n2579;
  assign new_n2581 = ~new_n2528 & new_n2579;
  assign new_n2582 = ~new_n2580 & ~new_n2581;
  assign new_n2583 = ~new_n2205 & new_n2582;
  assign new_n2584 = new_n2205 & ~new_n2582;
  assign new_n2585 = ~new_n2520 & ~new_n2521;
  assign new_n2586 = ~new_n2522 & ~new_n2585;
  assign new_n2587 = new_n2151 & new_n2586;
  assign new_n2588 = ~new_n2584 & ~new_n2587;
  assign new_n2589 = ~new_n2583 & ~new_n2588;
  assign new_n2590_1 = ~new_n2578 & ~new_n2589;
  assign new_n2591 = ~new_n2577 & ~new_n2590_1;
  assign new_n2592_1 = ~new_n2570 & ~new_n2591;
  assign new_n2593 = ~new_n2569 & ~new_n2592_1;
  assign new_n2594 = ~new_n2560 & ~new_n2593;
  assign new_n2595 = ~new_n2559 & ~new_n2594;
  assign new_n2596 = ~new_n2552 & ~new_n2595;
  assign new_n2597 = ~new_n2551 & ~new_n2596;
  assign new_n2598 = new_n2544 & new_n2597;
  assign new_n2599 = ~new_n2544 & ~new_n2597;
  assign new_n2600 = ~new_n2598 & ~new_n2599;
  assign new_n2601 = ~new_n2150 & ~new_n2600;
  assign new_n2602 = new_n2150 & new_n2600;
  assign new_n2603 = ~new_n2099 & ~new_n2101;
  assign new_n2604 = ~new_n2102 & ~new_n2603;
  assign new_n2605 = ~new_n2551 & ~new_n2552;
  assign new_n2606 = new_n2595 & ~new_n2605;
  assign new_n2607 = ~new_n2595 & new_n2605;
  assign new_n2608 = ~new_n2606 & ~new_n2607;
  assign new_n2609 = ~new_n2604 & new_n2608;
  assign new_n2610 = new_n2604 & ~new_n2608;
  assign new_n2611 = ~new_n2094 & ~new_n2098;
  assign new_n2612 = ~new_n2099 & ~new_n2611;
  assign new_n2613 = ~new_n2559 & ~new_n2560;
  assign new_n2614 = ~new_n2593 & ~new_n2613;
  assign new_n2615 = new_n2593 & new_n2613;
  assign new_n2616 = ~new_n2614 & ~new_n2615;
  assign new_n2617 = ~new_n2612 & ~new_n2616;
  assign new_n2618 = new_n2612 & new_n2616;
  assign new_n2619 = ~new_n2089 & ~new_n2093;
  assign new_n2620 = ~new_n2094 & ~new_n2619;
  assign new_n2621 = ~new_n2569 & ~new_n2570;
  assign new_n2622 = ~new_n2591 & ~new_n2621;
  assign new_n2623 = new_n2591 & new_n2621;
  assign new_n2624 = ~new_n2622 & ~new_n2623;
  assign new_n2625 = new_n2620 & new_n2624;
  assign new_n2626 = ~new_n2620 & ~new_n2624;
  assign new_n2627 = ~new_n2084 & ~new_n2088;
  assign new_n2628 = ~new_n2089 & ~new_n2627;
  assign new_n2629 = ~new_n2577 & ~new_n2578;
  assign new_n2630 = new_n2589 & ~new_n2629;
  assign new_n2631 = ~new_n2589 & new_n2629;
  assign new_n2632 = ~new_n2630 & ~new_n2631;
  assign new_n2633 = new_n2628 & ~new_n2632;
  assign new_n2634 = ~new_n2628 & new_n2632;
  assign new_n2635 = ~new_n2082 & ~new_n2083;
  assign new_n2636 = ~new_n2084 & ~new_n2635;
  assign new_n2637 = n2482 & n12853;
  assign new_n2638 = ~new_n2151 & ~new_n2586;
  assign new_n2639 = ~new_n2587 & ~new_n2638;
  assign new_n2640 = new_n2637 & new_n2639;
  assign new_n2641 = ~new_n2636 & ~new_n2640;
  assign new_n2642 = new_n2636 & new_n2640;
  assign new_n2643 = ~new_n2583 & ~new_n2584;
  assign new_n2644 = new_n2587 & ~new_n2643;
  assign new_n2645 = ~new_n2587 & new_n2643;
  assign new_n2646 = ~new_n2644 & ~new_n2645;
  assign new_n2647 = ~new_n2642 & new_n2646;
  assign new_n2648 = ~new_n2641 & ~new_n2647;
  assign new_n2649 = ~new_n2634 & new_n2648;
  assign new_n2650 = ~new_n2633 & ~new_n2649;
  assign new_n2651 = ~new_n2626 & ~new_n2650;
  assign new_n2652 = ~new_n2625 & ~new_n2651;
  assign new_n2653 = ~new_n2618 & new_n2652;
  assign new_n2654 = ~new_n2617 & ~new_n2653;
  assign new_n2655 = ~new_n2610 & ~new_n2654;
  assign new_n2656 = ~new_n2609 & ~new_n2655;
  assign new_n2657 = ~new_n2602 & ~new_n2656;
  assign new_n2658 = ~new_n2601 & ~new_n2657;
  assign new_n2659 = ~new_n2145 & ~new_n2148;
  assign new_n2660 = ~new_n2106 & ~new_n2141;
  assign new_n2661 = ~new_n2107 & ~new_n2660;
  assign new_n2662 = n1982 & n9531;
  assign new_n2663 = n9669 & n11030;
  assign new_n2664 = n9528 & n10416;
  assign new_n2665 = ~new_n2663 & ~new_n2664;
  assign new_n2666_1 = new_n2663 & new_n2664;
  assign new_n2667 = ~new_n2665 & ~new_n2666_1;
  assign new_n2668 = n8522 & n10113;
  assign new_n2669 = n1757 & n6655;
  assign new_n2670 = new_n2668 & ~new_n2669;
  assign new_n2671 = ~new_n2668 & new_n2669;
  assign new_n2672 = ~new_n2670 & ~new_n2671;
  assign new_n2673 = ~new_n2667 & ~new_n2672;
  assign new_n2674 = new_n2667 & new_n2672;
  assign new_n2675 = ~new_n2673 & ~new_n2674;
  assign new_n2676 = ~new_n2662 & new_n2675;
  assign new_n2677 = new_n2662 & ~new_n2675;
  assign new_n2678 = ~new_n2676 & ~new_n2677;
  assign new_n2679 = ~new_n2408 & new_n2465;
  assign new_n2680 = ~n9591 & new_n2408;
  assign new_n2681 = ~new_n2679 & ~new_n2680;
  assign new_n2682 = n10522 & n11222;
  assign new_n2683 = n2666 & n8940;
  assign new_n2684 = new_n2682 & ~new_n2683;
  assign new_n2685 = ~new_n2682 & new_n2683;
  assign new_n2686 = ~new_n2684 & ~new_n2685;
  assign new_n2687 = new_n2681 & ~new_n2686;
  assign new_n2688 = ~new_n2681 & new_n2686;
  assign new_n2689 = ~new_n2687 & ~new_n2688;
  assign new_n2690 = n4964 & n6023;
  assign new_n2691 = n5684 & n12579;
  assign new_n2692 = ~new_n2690 & new_n2691;
  assign new_n2693 = new_n2690 & ~new_n2691;
  assign new_n2694 = ~new_n2692 & ~new_n2693;
  assign new_n2695 = n8820 & n12853;
  assign new_n2696 = n11488 & n11891;
  assign new_n2697 = n2482 & n5427;
  assign new_n2698 = new_n2696 & new_n2697;
  assign new_n2699 = ~new_n2696 & ~new_n2697;
  assign new_n2700 = ~new_n2698 & ~new_n2699;
  assign new_n2701 = new_n2695 & ~new_n2700;
  assign new_n2702 = ~new_n2695 & new_n2700;
  assign new_n2703 = ~new_n2701 & ~new_n2702;
  assign new_n2704 = ~new_n2694 & new_n2703;
  assign new_n2705 = new_n2694 & ~new_n2703;
  assign new_n2706 = ~new_n2704 & ~new_n2705;
  assign new_n2707 = new_n2689 & ~new_n2706;
  assign new_n2708 = ~new_n2689 & new_n2706;
  assign new_n2709_1 = ~new_n2707 & ~new_n2708;
  assign new_n2710 = new_n2406 & new_n2681;
  assign new_n2711 = new_n2472 & ~new_n2475;
  assign new_n2712 = ~new_n2476 & ~new_n2711;
  assign new_n2713 = ~new_n2710 & ~new_n2712;
  assign new_n2714 = new_n2710 & new_n2712;
  assign new_n2715 = ~new_n2713 & ~new_n2714;
  assign new_n2716 = new_n2709_1 & new_n2715;
  assign new_n2717 = ~new_n2709_1 & ~new_n2715;
  assign new_n2718 = ~new_n2716 & ~new_n2717;
  assign new_n2719 = ~new_n2678 & new_n2718;
  assign new_n2720 = new_n2678 & ~new_n2718;
  assign new_n2721 = ~new_n2719 & ~new_n2720;
  assign new_n2722 = ~new_n2661 & new_n2721;
  assign new_n2723 = new_n2661 & ~new_n2721;
  assign new_n2724 = ~new_n2722 & ~new_n2723;
  assign new_n2725 = new_n2659 & ~new_n2724;
  assign new_n2726 = ~new_n2659 & new_n2724;
  assign new_n2727 = ~new_n2725 & ~new_n2726;
  assign new_n2728 = new_n2658 & new_n2727;
  assign new_n2729 = ~new_n2658 & ~new_n2727;
  assign new_n2730 = ~new_n2728 & ~new_n2729;
  assign new_n2731 = ~new_n2542 & new_n2597;
  assign new_n2732 = ~new_n2543 & ~new_n2731;
  assign new_n2733 = ~new_n2125 & ~new_n2135;
  assign new_n2734 = ~new_n2124 & ~new_n2733;
  assign new_n2735 = n9353 & n12693;
  assign new_n2736 = ~new_n2348 & ~new_n2377;
  assign new_n2737_1 = ~new_n2735 & new_n2736;
  assign new_n2738 = new_n2735 & ~new_n2736;
  assign new_n2739 = ~new_n2737_1 & ~new_n2738;
  assign new_n2740 = new_n2734 & new_n2739;
  assign new_n2741 = ~new_n2734 & ~new_n2739;
  assign new_n2742 = ~new_n2740 & ~new_n2741;
  assign new_n2743 = ~new_n2494 & ~new_n2538;
  assign new_n2744 = ~new_n2493 & ~new_n2743;
  assign new_n2745 = ~new_n2227 & ~new_n2230;
  assign new_n2746 = ~new_n2224 & new_n2745;
  assign new_n2747 = new_n2224 & ~new_n2745;
  assign new_n2748 = ~new_n2746 & ~new_n2747;
  assign new_n2749 = ~new_n2208 & ~new_n2220;
  assign new_n2750 = ~new_n2209 & ~new_n2749;
  assign new_n2751 = ~new_n2212 & new_n2217;
  assign new_n2752 = ~new_n2211 & ~new_n2751;
  assign new_n2753 = new_n2203 & new_n2752;
  assign new_n2754 = ~new_n2203 & ~new_n2752;
  assign new_n2755 = ~new_n2753 & ~new_n2754;
  assign new_n2756 = new_n2750 & ~new_n2755;
  assign new_n2757 = ~new_n2750 & new_n2755;
  assign new_n2758_1 = ~new_n2756 & ~new_n2757;
  assign new_n2759 = n389 & n8228;
  assign new_n2760 = new_n2217 & ~new_n2759;
  assign new_n2761 = ~new_n2217 & new_n2759;
  assign new_n2762 = ~new_n2760 & ~new_n2761;
  assign new_n2763 = ~new_n2152 & ~new_n2154;
  assign new_n2764 = n11236 & new_n2154;
  assign new_n2765 = ~new_n2763 & ~new_n2764;
  assign new_n2766 = n5320 & ~new_n2178;
  assign new_n2767 = ~new_n2177 & ~new_n2766;
  assign new_n2768 = new_n2765 & new_n2767;
  assign new_n2769 = ~new_n2765 & ~new_n2767;
  assign new_n2770 = ~new_n2768 & ~new_n2769;
  assign new_n2771_1 = new_n2762 & ~new_n2770;
  assign new_n2772 = ~new_n2762 & new_n2770;
  assign new_n2773 = ~new_n2771_1 & ~new_n2772;
  assign new_n2774 = ~new_n2758_1 & new_n2773;
  assign new_n2775 = new_n2758_1 & ~new_n2773;
  assign new_n2776 = ~new_n2774 & ~new_n2775;
  assign new_n2777_1 = ~new_n2748 & new_n2776;
  assign new_n2778 = new_n2748 & ~new_n2776;
  assign new_n2779 = ~new_n2777_1 & ~new_n2778;
  assign new_n2780 = new_n2744 & new_n2779;
  assign new_n2781 = ~new_n2744 & ~new_n2779;
  assign new_n2782 = ~new_n2780 & ~new_n2781;
  assign new_n2783 = new_n2742 & ~new_n2782;
  assign new_n2784 = ~new_n2742 & new_n2782;
  assign new_n2785 = ~new_n2783 & ~new_n2784;
  assign new_n2786 = ~new_n2469 & ~new_n2480;
  assign new_n2787 = n854 & n4743;
  assign new_n2788 = new_n2109 & ~new_n2112;
  assign new_n2789 = ~new_n2113 & ~new_n2788;
  assign new_n2790 = new_n2127 & ~new_n2130;
  assign new_n2791 = ~new_n2131 & ~new_n2790;
  assign new_n2792 = ~new_n2789 & new_n2791;
  assign new_n2793 = new_n2789 & ~new_n2791;
  assign new_n2794 = ~new_n2792 & ~new_n2793;
  assign new_n2795 = new_n2787 & new_n2794;
  assign new_n2796 = ~new_n2787 & ~new_n2794;
  assign new_n2797 = ~new_n2795 & ~new_n2796;
  assign new_n2798 = ~new_n2484 & ~new_n2487;
  assign new_n2799 = ~new_n2490 & new_n2798;
  assign new_n2800 = n761 & n5189;
  assign new_n2801 = n5758 & n8716;
  assign new_n2802 = ~new_n2800 & ~new_n2801;
  assign new_n2803 = new_n2800 & new_n2801;
  assign new_n2804 = ~new_n2802 & ~new_n2803;
  assign new_n2805_1 = n9620 & n13060;
  assign new_n2806 = n2295 & n12750;
  assign new_n2807 = new_n2805_1 & ~new_n2806;
  assign new_n2808 = ~new_n2805_1 & new_n2806;
  assign new_n2809 = ~new_n2807 & ~new_n2808;
  assign new_n2810 = ~new_n2804 & new_n2809;
  assign new_n2811 = new_n2804 & ~new_n2809;
  assign new_n2812 = ~new_n2810 & ~new_n2811;
  assign new_n2813 = ~new_n2307 & ~new_n2344;
  assign new_n2814 = ~new_n2308 & ~new_n2813;
  assign new_n2815 = new_n2310 & ~new_n2313;
  assign new_n2816 = ~new_n2314 & ~new_n2815;
  assign new_n2817 = ~new_n2323 & new_n2334;
  assign new_n2818 = ~new_n2324 & ~new_n2817;
  assign new_n2819 = ~new_n2816 & ~new_n2818;
  assign new_n2820 = new_n2816 & new_n2818;
  assign new_n2821 = ~new_n2819 & ~new_n2820;
  assign new_n2822 = new_n2326 & ~new_n2329;
  assign new_n2823 = ~new_n2330 & ~new_n2822;
  assign new_n2824 = ~new_n2821 & new_n2823;
  assign new_n2825 = new_n2821 & ~new_n2823;
  assign new_n2826 = ~new_n2824 & ~new_n2825;
  assign new_n2827 = n834 & n12352;
  assign new_n2828 = n2341 & n6333;
  assign new_n2829 = n1650 & n1912;
  assign new_n2830 = ~new_n2828 & new_n2829;
  assign new_n2831 = new_n2828 & ~new_n2829;
  assign new_n2832 = ~new_n2830 & ~new_n2831;
  assign new_n2833 = new_n2827 & new_n2832;
  assign new_n2834 = ~new_n2827 & ~new_n2832;
  assign new_n2835 = ~new_n2833 & ~new_n2834;
  assign new_n2836 = new_n2341_1 & new_n2835;
  assign new_n2837 = ~new_n2341_1 & ~new_n2835;
  assign new_n2838 = ~new_n2836 & ~new_n2837;
  assign new_n2839 = new_n2826 & new_n2838;
  assign new_n2840 = ~new_n2826 & ~new_n2838;
  assign new_n2841 = ~new_n2839 & ~new_n2840;
  assign new_n2842 = new_n2814 & new_n2841;
  assign new_n2843 = ~new_n2814 & ~new_n2841;
  assign new_n2844 = ~new_n2842 & ~new_n2843;
  assign new_n2845 = new_n2812 & new_n2844;
  assign new_n2846 = ~new_n2812 & ~new_n2844;
  assign new_n2847 = ~new_n2845 & ~new_n2846;
  assign new_n2848 = ~new_n2799 & new_n2847;
  assign new_n2849 = new_n2799 & ~new_n2847;
  assign new_n2850 = ~new_n2848 & ~new_n2849;
  assign new_n2851 = ~new_n2120 & new_n2138;
  assign new_n2852 = ~new_n2121 & ~new_n2851;
  assign new_n2853 = ~new_n2850 & new_n2852;
  assign new_n2854 = new_n2850 & ~new_n2852;
  assign new_n2855 = ~new_n2853 & ~new_n2854;
  assign new_n2856 = ~new_n2797 & new_n2855;
  assign new_n2857 = new_n2797 & ~new_n2855;
  assign new_n2858 = ~new_n2856 & ~new_n2857;
  assign new_n2859 = new_n2786 & new_n2858;
  assign new_n2860 = ~new_n2786 & ~new_n2858;
  assign new_n2861 = ~new_n2859 & ~new_n2860;
  assign new_n2862 = new_n2785 & ~new_n2861;
  assign new_n2863 = ~new_n2785 & new_n2861;
  assign new_n2864 = ~new_n2862 & ~new_n2863;
  assign new_n2865 = ~new_n2732 & new_n2864;
  assign new_n2866 = new_n2732 & ~new_n2864;
  assign new_n2867 = ~new_n2865 & ~new_n2866;
  assign new_n2868 = new_n2730 & new_n2867;
  assign new_n2869 = ~new_n2730 & ~new_n2867;
  assign n370 = ~new_n2868 & ~new_n2869;
  assign new_n2871 = n5568 & n9528;
  assign new_n2872 = n8308 & n9669;
  assign new_n2873 = ~new_n2871 & ~new_n2872;
  assign new_n2874 = new_n2871 & new_n2872;
  assign new_n2875 = ~new_n2873 & ~new_n2874;
  assign new_n2876 = n5214 & n11891;
  assign new_n2877 = n2771 & n9531;
  assign new_n2878 = n6168 & n12853;
  assign new_n2879 = ~new_n2877 & ~new_n2878;
  assign new_n2880 = new_n2877 & new_n2878;
  assign new_n2881 = ~new_n2879 & ~new_n2880;
  assign new_n2882_1 = ~new_n2876 & ~new_n2881;
  assign new_n2883 = new_n2876 & new_n2881;
  assign new_n2884 = ~new_n2882_1 & ~new_n2883;
  assign new_n2885 = n8308 & n11891;
  assign new_n2886 = n5214 & n9531;
  assign new_n2887 = new_n2885 & new_n2886;
  assign new_n2888 = n2771 & n12853;
  assign new_n2889 = ~new_n2885 & ~new_n2886;
  assign new_n2890 = new_n2888 & ~new_n2889;
  assign new_n2891 = ~new_n2887 & ~new_n2890;
  assign new_n2892 = ~new_n2884 & new_n2891;
  assign new_n2893 = new_n2884 & ~new_n2891;
  assign new_n2894 = ~new_n2892 & ~new_n2893;
  assign new_n2895 = ~new_n2875 & ~new_n2894;
  assign new_n2896 = new_n2875 & new_n2894;
  assign new_n2897 = ~new_n2895 & ~new_n2896;
  assign new_n2898 = n5568 & n9669;
  assign new_n2899 = n8308 & n9531;
  assign new_n2900 = n5568 & n11891;
  assign new_n2901 = new_n2899 & new_n2900;
  assign new_n2902 = ~new_n2899 & ~new_n2900;
  assign new_n2903 = n5214 & n12853;
  assign new_n2904_1 = ~new_n2902 & new_n2903;
  assign new_n2905 = ~new_n2901 & ~new_n2904_1;
  assign new_n2906 = ~new_n2898 & new_n2905;
  assign new_n2907 = new_n2898 & ~new_n2905;
  assign new_n2908 = ~new_n2887 & ~new_n2889;
  assign new_n2909 = new_n2888 & ~new_n2908;
  assign new_n2910 = ~new_n2888 & new_n2908;
  assign new_n2911 = ~new_n2909 & ~new_n2910;
  assign new_n2912 = ~new_n2907 & new_n2911;
  assign new_n2913 = ~new_n2906 & ~new_n2912;
  assign new_n2914 = ~new_n2897 & ~new_n2913;
  assign new_n2915 = new_n2897 & new_n2913;
  assign new_n2916 = ~new_n2914 & ~new_n2915;
  assign new_n2917 = n3006 & n9528;
  assign new_n2918 = ~new_n2906 & ~new_n2907;
  assign new_n2919 = new_n2911 & ~new_n2918;
  assign new_n2920 = ~new_n2911 & new_n2918;
  assign new_n2921 = ~new_n2919 & ~new_n2920;
  assign new_n2922 = new_n2917 & new_n2921;
  assign new_n2923 = ~new_n2917 & ~new_n2921;
  assign new_n2924 = n3006 & n9669;
  assign new_n2925 = n5568 & n9531;
  assign new_n2926 = n3006 & n11891;
  assign new_n2927 = new_n2925 & new_n2926;
  assign new_n2928 = ~new_n2925 & ~new_n2926;
  assign new_n2929 = n8308 & n12853;
  assign new_n2930 = ~new_n2928 & new_n2929;
  assign new_n2931 = ~new_n2927 & ~new_n2930;
  assign new_n2932 = ~new_n2924 & new_n2931;
  assign new_n2933 = new_n2924 & ~new_n2931;
  assign new_n2934_1 = ~new_n2901 & ~new_n2902;
  assign new_n2935 = ~new_n2903 & ~new_n2934_1;
  assign new_n2936 = new_n2903 & new_n2934_1;
  assign new_n2937 = ~new_n2935 & ~new_n2936;
  assign new_n2938 = ~new_n2933 & ~new_n2937;
  assign new_n2939 = ~new_n2932 & ~new_n2938;
  assign new_n2940 = ~new_n2923 & new_n2939;
  assign new_n2941 = ~new_n2922 & ~new_n2940;
  assign new_n2942 = new_n2916 & ~new_n2941;
  assign new_n2943 = ~new_n2895 & new_n2913;
  assign new_n2944 = ~new_n2874 & ~new_n2943;
  assign new_n2945 = ~new_n2896 & new_n2944;
  assign new_n2946 = new_n2874 & new_n2943;
  assign new_n2947 = ~new_n2945 & ~new_n2946;
  assign new_n2948 = n8308 & n9528;
  assign new_n2949 = n3006 & n8522;
  assign new_n2950 = n5568 & n6655;
  assign new_n2951 = ~new_n2949 & ~new_n2950;
  assign new_n2952 = new_n2949 & new_n2950;
  assign new_n2953 = ~new_n2951 & ~new_n2952;
  assign new_n2954 = new_n2948 & ~new_n2953;
  assign new_n2955 = ~new_n2948 & new_n2953;
  assign new_n2956 = ~new_n2954 & ~new_n2955;
  assign new_n2957 = ~new_n2883 & new_n2891;
  assign new_n2958 = ~new_n2882_1 & ~new_n2957;
  assign new_n2959 = new_n2956 & ~new_n2958;
  assign new_n2960 = n5214 & n9669;
  assign new_n2961 = ~new_n2880 & ~new_n2960;
  assign new_n2962 = new_n2880 & new_n2960;
  assign new_n2963 = ~new_n2961 & ~new_n2962;
  assign new_n2964 = n11411 & n12853;
  assign new_n2965 = n6168 & n9531;
  assign new_n2966 = n2771 & n11891;
  assign new_n2967 = ~new_n2965 & ~new_n2966;
  assign new_n2968 = new_n2965 & new_n2966;
  assign new_n2969 = ~new_n2967 & ~new_n2968;
  assign new_n2970 = new_n2964 & ~new_n2969;
  assign new_n2971 = ~new_n2964 & new_n2969;
  assign new_n2972 = ~new_n2970 & ~new_n2971;
  assign new_n2973 = new_n2963 & new_n2972;
  assign new_n2974 = ~new_n2963 & ~new_n2972;
  assign new_n2975 = ~new_n2973 & ~new_n2974;
  assign new_n2976 = new_n2959 & new_n2975;
  assign new_n2977 = ~new_n2956 & new_n2958;
  assign new_n2978 = ~new_n2975 & new_n2977;
  assign new_n2979 = ~new_n2959 & ~new_n2975;
  assign new_n2980 = ~new_n2977 & ~new_n2979;
  assign new_n2981 = ~new_n2978 & ~new_n2980;
  assign new_n2982 = ~new_n2976 & ~new_n2981;
  assign new_n2983 = ~new_n2947 & ~new_n2982;
  assign new_n2984 = new_n2947 & new_n2982;
  assign new_n2985 = ~new_n2983 & ~new_n2984;
  assign new_n2986 = ~new_n2942 & ~new_n2985;
  assign new_n2987 = new_n2942 & new_n2985;
  assign new_n2988 = ~new_n2986 & ~new_n2987;
  assign new_n2989 = n3006 & n6655;
  assign new_n2990 = ~new_n2916 & new_n2941;
  assign new_n2991 = ~new_n2942 & ~new_n2990;
  assign new_n2992 = new_n2989 & new_n2991;
  assign new_n2993 = n3006 & n9531;
  assign new_n2994 = n5568 & n12853;
  assign new_n2995 = new_n2993 & new_n2994;
  assign new_n2996 = ~new_n2927 & ~new_n2928;
  assign new_n2997 = ~new_n2929 & ~new_n2996;
  assign new_n2998 = new_n2929 & new_n2996;
  assign new_n2999 = ~new_n2997 & ~new_n2998;
  assign new_n3000 = new_n2995 & new_n2999;
  assign new_n3001 = ~new_n2932 & ~new_n2933;
  assign new_n3002 = new_n2937 & ~new_n3001;
  assign new_n3003 = ~new_n2937 & new_n3001;
  assign new_n3004 = ~new_n3002 & ~new_n3003;
  assign new_n3005 = new_n3000 & ~new_n3004;
  assign new_n3006_1 = ~new_n2922 & ~new_n2923;
  assign new_n3007 = ~new_n2939 & ~new_n3006_1;
  assign new_n3008 = new_n2939 & new_n3006_1;
  assign new_n3009 = ~new_n3007 & ~new_n3008;
  assign new_n3010 = new_n3005 & new_n3009;
  assign new_n3011 = ~new_n2989 & ~new_n2991;
  assign new_n3012 = ~new_n2992 & ~new_n3011;
  assign new_n3013 = new_n3010 & new_n3012;
  assign new_n3014 = ~new_n2992 & ~new_n3013;
  assign new_n3015 = ~new_n2988 & new_n3014;
  assign new_n3016 = new_n2988 & ~new_n3014;
  assign new_n3017 = ~new_n3015 & ~new_n3016;
  assign new_n3018 = n854 & n10560;
  assign new_n3019 = n12003 & new_n3018;
  assign new_n3020 = ~n5801 & ~new_n3019;
  assign new_n3021 = n854 & n12003;
  assign new_n3022 = ~new_n3018 & ~new_n3021;
  assign new_n3023 = n5801 & ~new_n3022;
  assign new_n3024 = n854 & n10908;
  assign new_n3025 = ~new_n3023 & ~new_n3024;
  assign new_n3026 = ~new_n3020 & ~new_n3025;
  assign new_n3027 = ~new_n3018 & ~new_n3024;
  assign new_n3028 = n10908 & new_n3018;
  assign new_n3029 = ~new_n3027 & ~new_n3028;
  assign new_n3030 = n854 & n8139;
  assign new_n3031 = ~new_n3019 & ~new_n3022;
  assign new_n3032 = ~new_n3030 & ~new_n3031;
  assign new_n3033 = new_n3030 & new_n3031;
  assign new_n3034 = ~new_n3032 & ~new_n3033;
  assign new_n3035 = ~new_n3029 & ~new_n3034;
  assign new_n3036 = new_n3029 & new_n3030;
  assign new_n3037 = ~new_n3035 & ~new_n3036;
  assign new_n3038 = new_n3026 & new_n3037;
  assign new_n3039 = new_n3018 & new_n3021;
  assign new_n3040 = new_n3034 & new_n3039;
  assign new_n3041 = ~new_n3028 & ~new_n3040;
  assign new_n3042 = ~n12003 & ~new_n3030;
  assign new_n3043 = new_n3024 & ~new_n3042;
  assign new_n3044 = ~new_n3018 & ~new_n3043;
  assign new_n3045 = new_n3041 & ~new_n3044;
  assign new_n3046 = n854 & n3311;
  assign new_n3047 = ~n8139 & n10560;
  assign new_n3048 = ~n10560 & new_n3030;
  assign new_n3049 = ~new_n3021 & ~new_n3048;
  assign new_n3050 = ~new_n3047 & ~new_n3049;
  assign new_n3051 = new_n3046 & new_n3050;
  assign new_n3052 = ~new_n3046 & ~new_n3050;
  assign new_n3053 = ~new_n3051 & ~new_n3052;
  assign new_n3054 = ~new_n3045 & new_n3053;
  assign new_n3055 = new_n3045 & ~new_n3053;
  assign new_n3056 = ~new_n3054 & ~new_n3055;
  assign new_n3057 = new_n3038 & ~new_n3056;
  assign new_n3058 = ~new_n3038 & new_n3056;
  assign new_n3059 = ~new_n3057 & ~new_n3058;
  assign new_n3060 = new_n1455 & new_n3059;
  assign new_n3061 = ~new_n3026 & ~new_n3037;
  assign new_n3062 = ~new_n3038 & ~new_n3061;
  assign new_n3063 = n10908 & new_n1455;
  assign new_n3064 = n12003 & ~new_n3029;
  assign new_n3065 = new_n3063 & new_n3064;
  assign new_n3066 = new_n3062 & new_n3065;
  assign new_n3067 = ~new_n1455 & ~new_n3059;
  assign new_n3068 = ~new_n3060 & ~new_n3067;
  assign new_n3069 = new_n3066 & new_n3068;
  assign new_n3070 = ~new_n3060 & ~new_n3069;
  assign new_n3071 = new_n3041 & ~new_n3053;
  assign new_n3072 = ~new_n3044 & ~new_n3071;
  assign new_n3073 = ~new_n1455 & ~new_n3024;
  assign new_n3074 = ~new_n3063 & ~new_n3073;
  assign new_n3075 = ~new_n3030 & ~new_n3046;
  assign new_n3076_1 = ~new_n3019 & new_n3075;
  assign new_n3077 = n3311 & ~new_n3021;
  assign new_n3078 = ~new_n3022 & ~new_n3077;
  assign new_n3079 = ~new_n3076_1 & new_n3078;
  assign new_n3080 = ~new_n3074 & ~new_n3079;
  assign new_n3081 = new_n3074 & new_n3079;
  assign new_n3082 = ~new_n3080 & ~new_n3081;
  assign new_n3083 = n8139 & new_n3046;
  assign new_n3084 = ~new_n3075 & ~new_n3083;
  assign new_n3085_1 = n854 & ~n10866;
  assign new_n3086 = ~new_n3084 & ~new_n3085_1;
  assign new_n3087 = new_n3084 & new_n3085_1;
  assign new_n3088 = ~new_n3086 & ~new_n3087;
  assign new_n3089 = n12003 & new_n3083;
  assign new_n3090 = ~new_n3021 & ~new_n3083;
  assign new_n3091 = ~new_n3089 & ~new_n3090;
  assign new_n3092 = new_n3088 & new_n3091;
  assign new_n3093 = ~new_n3088 & ~new_n3091;
  assign new_n3094 = ~new_n3092 & ~new_n3093;
  assign new_n3095 = new_n3082 & ~new_n3094;
  assign new_n3096 = ~new_n3082 & new_n3094;
  assign new_n3097 = ~new_n3095 & ~new_n3096;
  assign new_n3098 = new_n3072 & ~new_n3097;
  assign new_n3099 = ~new_n3072 & new_n3097;
  assign new_n3100 = ~new_n3098 & ~new_n3099;
  assign new_n3101 = new_n3057 & new_n3100;
  assign new_n3102 = ~new_n3057 & ~new_n3100;
  assign new_n3103 = ~new_n3101 & ~new_n3102;
  assign new_n3104 = ~new_n3070 & new_n3103;
  assign new_n3105 = new_n3070 & ~new_n3103;
  assign new_n3106 = ~new_n3104 & ~new_n3105;
  assign new_n3107 = n8290 & n11665;
  assign new_n3108 = n4114 & n9591;
  assign new_n3109 = new_n3107 & new_n3108;
  assign new_n3110 = ~new_n3107 & ~new_n3108;
  assign new_n3111 = n510 & n2777;
  assign new_n3112_1 = ~new_n3110 & new_n3111;
  assign new_n3113 = ~new_n3109 & ~new_n3112_1;
  assign new_n3114 = n510 & n10642;
  assign new_n3115 = n9591 & n11665;
  assign new_n3116 = n2777 & n8290;
  assign new_n3117 = ~new_n3115 & ~new_n3116;
  assign new_n3118 = new_n3115 & new_n3116;
  assign new_n3119 = ~new_n3117 & ~new_n3118;
  assign new_n3120 = new_n3114 & ~new_n3119;
  assign new_n3121 = ~new_n3114 & new_n3119;
  assign new_n3122 = ~new_n3120 & ~new_n3121;
  assign new_n3123 = ~new_n3113 & ~new_n3122;
  assign new_n3124 = n4114 & n11222;
  assign new_n3125 = ~new_n3123 & ~new_n3124;
  assign new_n3126 = new_n3123 & new_n3124;
  assign new_n3127 = ~new_n3125 & ~new_n3126;
  assign new_n3128 = n2777 & n9591;
  assign new_n3129 = n8290 & n10642;
  assign new_n3130_1 = n510 & n937;
  assign new_n3131 = ~new_n3129 & ~new_n3130_1;
  assign new_n3132 = new_n3129 & new_n3130_1;
  assign new_n3133 = ~new_n3131 & ~new_n3132;
  assign new_n3134 = ~new_n3128 & ~new_n3133;
  assign new_n3135 = new_n3128 & new_n3133;
  assign new_n3136 = ~new_n3134 & ~new_n3135;
  assign new_n3137 = new_n3114 & ~new_n3117;
  assign new_n3138 = ~new_n3118 & ~new_n3137;
  assign new_n3139 = ~new_n3136 & new_n3138;
  assign new_n3140 = new_n3136 & ~new_n3138;
  assign new_n3141 = ~new_n3139 & ~new_n3140;
  assign new_n3142 = new_n3127 & new_n3141;
  assign new_n3143 = ~new_n3127 & ~new_n3141;
  assign new_n3144 = ~new_n3142 & ~new_n3143;
  assign new_n3145 = ~new_n3109 & ~new_n3110;
  assign new_n3146 = ~new_n3111 & ~new_n3145;
  assign new_n3147 = new_n3111 & new_n3145;
  assign new_n3148 = ~new_n3146 & ~new_n3147;
  assign new_n3149 = n4114 & n8290;
  assign new_n3150 = n5671 & n9591;
  assign new_n3151 = new_n3149 & new_n3150;
  assign new_n3152 = ~new_n3149 & ~new_n3150;
  assign new_n3153 = n510 & n11665;
  assign new_n3154 = ~new_n3152 & new_n3153;
  assign new_n3155 = ~new_n3151 & ~new_n3154;
  assign new_n3156 = new_n3148 & ~new_n3155;
  assign new_n3157 = n5671 & n11222;
  assign new_n3158 = ~new_n3156 & ~new_n3157;
  assign new_n3159 = new_n3156 & new_n3157;
  assign new_n3160 = new_n3113 & new_n3122;
  assign new_n3161 = ~new_n3123 & ~new_n3160;
  assign new_n3162 = ~new_n3159 & ~new_n3161;
  assign new_n3163 = ~new_n3158 & ~new_n3162;
  assign new_n3164 = new_n3144 & new_n3163;
  assign new_n3165 = n510 & n12605;
  assign new_n3166 = n937 & n8290;
  assign new_n3167 = n9591 & n10642;
  assign new_n3168 = ~new_n3166 & ~new_n3167;
  assign new_n3169 = new_n3166 & new_n3167;
  assign new_n3170 = ~new_n3168 & ~new_n3169;
  assign new_n3171 = new_n3165 & ~new_n3170;
  assign new_n3172 = ~new_n3165 & new_n3170;
  assign new_n3173 = ~new_n3171 & ~new_n3172;
  assign new_n3174 = ~new_n3132 & new_n3173;
  assign new_n3175 = new_n3132 & ~new_n3173;
  assign new_n3176 = ~new_n3174 & ~new_n3175;
  assign new_n3177 = n11222 & n11665;
  assign new_n3178_1 = n5671 & n6023;
  assign new_n3179 = n4114 & n12579;
  assign new_n3180 = ~new_n3178_1 & ~new_n3179;
  assign new_n3181 = new_n3178_1 & new_n3179;
  assign new_n3182 = ~new_n3180 & ~new_n3181;
  assign new_n3183 = new_n3177 & ~new_n3182;
  assign new_n3184 = ~new_n3177 & new_n3182;
  assign new_n3185 = ~new_n3183 & ~new_n3184;
  assign new_n3186 = ~new_n3135 & new_n3138;
  assign new_n3187 = ~new_n3134 & ~new_n3186;
  assign new_n3188 = ~new_n3185 & new_n3187;
  assign new_n3189 = new_n3185 & ~new_n3187;
  assign new_n3190 = ~new_n3188 & ~new_n3189;
  assign new_n3191 = ~new_n3176 & new_n3190;
  assign new_n3192 = new_n3176 & ~new_n3190;
  assign new_n3193 = ~new_n3191 & ~new_n3192;
  assign new_n3194 = ~new_n3126 & ~new_n3141;
  assign new_n3195 = ~new_n3125 & ~new_n3194;
  assign new_n3196 = new_n3193 & ~new_n3195;
  assign new_n3197 = ~new_n3193 & new_n3195;
  assign new_n3198 = ~new_n3196 & ~new_n3197;
  assign new_n3199 = ~new_n3164 & ~new_n3198;
  assign new_n3200 = new_n3164 & new_n3198;
  assign new_n3201 = ~new_n3199 & ~new_n3200;
  assign new_n3202 = n5671 & n12579;
  assign new_n3203 = ~new_n3144 & ~new_n3163;
  assign new_n3204 = ~new_n3164 & ~new_n3203;
  assign new_n3205 = new_n3202 & new_n3204;
  assign new_n3206 = n5671 & n8290;
  assign new_n3207 = n510 & n4114;
  assign new_n3208 = new_n3206 & new_n3207;
  assign new_n3209 = ~new_n3151 & ~new_n3152;
  assign new_n3210 = ~new_n3153 & ~new_n3209;
  assign new_n3211 = new_n3153 & new_n3209;
  assign new_n3212 = ~new_n3210 & ~new_n3211;
  assign new_n3213 = new_n3208 & new_n3212;
  assign new_n3214 = ~new_n3148 & new_n3155;
  assign new_n3215 = ~new_n3156 & ~new_n3214;
  assign new_n3216 = new_n3213 & new_n3215;
  assign new_n3217 = ~new_n3158 & ~new_n3159;
  assign new_n3218 = new_n3161 & ~new_n3217;
  assign new_n3219 = ~new_n3161 & new_n3217;
  assign new_n3220 = ~new_n3218 & ~new_n3219;
  assign new_n3221 = new_n3216 & ~new_n3220;
  assign new_n3222 = ~new_n3202 & ~new_n3204;
  assign new_n3223 = ~new_n3205 & ~new_n3222;
  assign new_n3224 = new_n3221 & new_n3223;
  assign new_n3225 = ~new_n3205 & ~new_n3224;
  assign new_n3226 = ~new_n3201 & new_n3225;
  assign new_n3227 = new_n3201 & ~new_n3225;
  assign new_n3228 = ~new_n3226 & ~new_n3227;
  assign new_n3229 = n5586 & n13060;
  assign new_n3230 = n2057 & n2295;
  assign new_n3231 = ~new_n3229 & ~new_n3230;
  assign new_n3232 = new_n3229 & new_n3230;
  assign new_n3233 = ~new_n3231 & ~new_n3232;
  assign new_n3234 = n4141 & n5189;
  assign new_n3235 = n1364 & n8716;
  assign new_n3236 = n834 & n3669;
  assign new_n3237 = ~new_n3235 & ~new_n3236;
  assign new_n3238 = new_n3235 & new_n3236;
  assign new_n3239 = ~new_n3237 & ~new_n3238;
  assign new_n3240 = new_n3234 & new_n3239;
  assign new_n3241 = ~new_n3234 & ~new_n3239;
  assign new_n3242 = ~new_n3240 & ~new_n3241;
  assign new_n3243 = n5189 & n5586;
  assign new_n3244 = n4141 & n8716;
  assign new_n3245 = new_n3243 & new_n3244;
  assign new_n3246 = ~new_n3243 & ~new_n3244;
  assign new_n3247 = n834 & n1364;
  assign new_n3248 = ~new_n3246 & new_n3247;
  assign new_n3249 = ~new_n3245 & ~new_n3248;
  assign new_n3250 = ~new_n3242 & new_n3249;
  assign new_n3251 = new_n3242 & ~new_n3249;
  assign new_n3252 = ~new_n3250 & ~new_n3251;
  assign new_n3253 = ~new_n3233 & ~new_n3252;
  assign new_n3254 = new_n3233 & new_n3252;
  assign new_n3255 = ~new_n3253 & ~new_n3254;
  assign new_n3256 = n2057 & n13060;
  assign new_n3257 = n5586 & n8716;
  assign new_n3258 = n2057 & n5189;
  assign new_n3259 = new_n3257 & new_n3258;
  assign new_n3260 = ~new_n3257 & ~new_n3258;
  assign new_n3261 = n834 & n4141;
  assign new_n3262_1 = ~new_n3260 & new_n3261;
  assign new_n3263 = ~new_n3259 & ~new_n3262_1;
  assign new_n3264 = ~new_n3256 & new_n3263;
  assign new_n3265 = new_n3256 & ~new_n3263;
  assign new_n3266 = ~new_n3245 & ~new_n3246;
  assign new_n3267 = ~new_n3247 & ~new_n3266;
  assign new_n3268 = new_n3247 & new_n3266;
  assign new_n3269 = ~new_n3267 & ~new_n3268;
  assign new_n3270 = ~new_n3265 & ~new_n3269;
  assign new_n3271 = ~new_n3264 & ~new_n3270;
  assign new_n3272 = ~new_n3255 & new_n3271;
  assign new_n3273 = new_n3255 & ~new_n3271;
  assign new_n3274 = ~new_n3272 & ~new_n3273;
  assign new_n3275 = n2295 & n13201;
  assign new_n3276 = ~new_n3264 & ~new_n3265;
  assign new_n3277 = ~new_n3269 & ~new_n3276;
  assign new_n3278 = new_n3269 & new_n3276;
  assign new_n3279 = ~new_n3277 & ~new_n3278;
  assign new_n3280 = new_n3275 & new_n3279;
  assign new_n3281 = ~new_n3275 & ~new_n3279;
  assign new_n3282 = n13060 & n13201;
  assign new_n3283 = n2057 & n8716;
  assign new_n3284 = n5189 & n13201;
  assign new_n3285 = new_n3283 & new_n3284;
  assign new_n3286 = ~new_n3283 & ~new_n3284;
  assign new_n3287 = n834 & n5586;
  assign new_n3288 = ~new_n3286 & new_n3287;
  assign new_n3289 = ~new_n3285 & ~new_n3288;
  assign new_n3290 = ~new_n3282 & new_n3289;
  assign new_n3291 = new_n3282 & ~new_n3289;
  assign new_n3292 = ~new_n3259 & ~new_n3260;
  assign new_n3293 = ~new_n3261 & ~new_n3292;
  assign new_n3294 = new_n3261 & new_n3292;
  assign new_n3295 = ~new_n3293 & ~new_n3294;
  assign new_n3296 = ~new_n3291 & ~new_n3295;
  assign new_n3297 = ~new_n3290 & ~new_n3296;
  assign new_n3298 = ~new_n3281 & new_n3297;
  assign new_n3299 = ~new_n3280 & ~new_n3298;
  assign new_n3300 = ~new_n3274 & ~new_n3299;
  assign new_n3301 = ~new_n3253 & new_n3271;
  assign new_n3302 = ~new_n3232 & ~new_n3301;
  assign new_n3303 = ~new_n3254 & new_n3302;
  assign new_n3304 = new_n3232 & new_n3301;
  assign new_n3305 = ~new_n3303 & ~new_n3304;
  assign new_n3306 = n2295 & n5586;
  assign new_n3307 = n2341 & n13201;
  assign new_n3308 = n1650 & n2057;
  assign new_n3309 = ~new_n3307 & ~new_n3308;
  assign new_n3310 = new_n3307 & new_n3308;
  assign new_n3311_1 = ~new_n3309 & ~new_n3310;
  assign new_n3312 = new_n3306 & ~new_n3311_1;
  assign new_n3313 = ~new_n3306 & new_n3311_1;
  assign new_n3314 = ~new_n3312 & ~new_n3313;
  assign new_n3315 = ~new_n3240 & new_n3249;
  assign new_n3316 = ~new_n3241 & ~new_n3315;
  assign new_n3317 = new_n3314 & ~new_n3316;
  assign new_n3318 = n4141 & n13060;
  assign new_n3319 = new_n3238 & new_n3318;
  assign new_n3320 = ~new_n3238 & ~new_n3318;
  assign new_n3321 = ~new_n3319 & ~new_n3320;
  assign new_n3322 = n834 & n5470;
  assign new_n3323_1 = n3669 & n8716;
  assign new_n3324 = n1364 & n5189;
  assign new_n3325 = ~new_n3323_1 & ~new_n3324;
  assign new_n3326 = new_n3323_1 & new_n3324;
  assign new_n3327 = ~new_n3325 & ~new_n3326;
  assign new_n3328 = new_n3322 & ~new_n3327;
  assign new_n3329 = ~new_n3322 & new_n3327;
  assign new_n3330 = ~new_n3328 & ~new_n3329;
  assign new_n3331 = new_n3321 & new_n3330;
  assign new_n3332 = ~new_n3321 & ~new_n3330;
  assign new_n3333 = ~new_n3331 & ~new_n3332;
  assign new_n3334 = new_n3317 & new_n3333;
  assign new_n3335 = ~new_n3314 & new_n3316;
  assign new_n3336 = new_n3333 & ~new_n3335;
  assign new_n3337 = ~new_n3317 & ~new_n3336;
  assign new_n3338 = ~new_n3334 & ~new_n3337;
  assign new_n3339 = ~new_n3333 & new_n3335;
  assign new_n3340 = ~new_n3338 & ~new_n3339;
  assign new_n3341 = ~new_n3305 & new_n3340;
  assign new_n3342 = new_n3305 & ~new_n3340;
  assign new_n3343 = ~new_n3341 & ~new_n3342;
  assign new_n3344 = ~new_n3300 & ~new_n3343;
  assign new_n3345 = new_n3300 & new_n3343;
  assign new_n3346 = ~new_n3344 & ~new_n3345;
  assign new_n3347 = n1650 & n13201;
  assign new_n3348 = new_n3274 & new_n3299;
  assign new_n3349 = ~new_n3300 & ~new_n3348;
  assign new_n3350 = new_n3347 & new_n3349;
  assign new_n3351 = n8716 & n13201;
  assign new_n3352 = n834 & n2057;
  assign new_n3353 = new_n3351 & new_n3352;
  assign new_n3354 = ~new_n3285 & ~new_n3286;
  assign new_n3355 = ~new_n3287 & ~new_n3354;
  assign new_n3356 = new_n3287 & new_n3354;
  assign new_n3357 = ~new_n3355 & ~new_n3356;
  assign new_n3358 = new_n3353 & new_n3357;
  assign new_n3359 = ~new_n3290 & ~new_n3291;
  assign new_n3360 = new_n3295 & ~new_n3359;
  assign new_n3361 = ~new_n3295 & new_n3359;
  assign new_n3362_1 = ~new_n3360 & ~new_n3361;
  assign new_n3363 = new_n3358 & ~new_n3362_1;
  assign new_n3364 = ~new_n3280 & ~new_n3281;
  assign new_n3365 = new_n3297 & new_n3364;
  assign new_n3366 = ~new_n3297 & ~new_n3364;
  assign new_n3367 = ~new_n3365 & ~new_n3366;
  assign new_n3368 = new_n3363 & new_n3367;
  assign new_n3369 = ~new_n3347 & ~new_n3349;
  assign new_n3370 = ~new_n3350 & ~new_n3369;
  assign new_n3371 = new_n3368 & new_n3370;
  assign new_n3372 = ~new_n3350 & ~new_n3371;
  assign new_n3373 = ~new_n3346 & new_n3372;
  assign new_n3374 = new_n3346 & ~new_n3372;
  assign new_n3375 = ~new_n3373 & ~new_n3374;
  assign new_n3376 = new_n3228 & new_n3375;
  assign new_n3377 = ~new_n3228 & ~new_n3375;
  assign new_n3378 = ~new_n3376 & ~new_n3377;
  assign new_n3379 = ~new_n3221 & ~new_n3223;
  assign new_n3380 = ~new_n3224 & ~new_n3379;
  assign new_n3381 = ~new_n3368 & ~new_n3370;
  assign new_n3382 = ~new_n3371 & ~new_n3381;
  assign new_n3383 = ~new_n3380 & ~new_n3382;
  assign new_n3384 = new_n3380 & new_n3382;
  assign new_n3385 = ~new_n3363 & ~new_n3367;
  assign new_n3386 = ~new_n3368 & ~new_n3385;
  assign new_n3387 = ~new_n3216 & new_n3220;
  assign new_n3388 = ~new_n3221 & ~new_n3387;
  assign new_n3389 = new_n3386 & new_n3388;
  assign new_n3390 = ~new_n3386 & ~new_n3388;
  assign new_n3391 = ~new_n3213 & ~new_n3215;
  assign new_n3392 = ~new_n3216 & ~new_n3391;
  assign new_n3393 = ~new_n3358 & new_n3362_1;
  assign new_n3394 = ~new_n3363 & ~new_n3393;
  assign new_n3395 = new_n3392 & new_n3394;
  assign new_n3396 = ~new_n3392 & ~new_n3394;
  assign new_n3397 = ~new_n3353 & ~new_n3357;
  assign new_n3398 = ~new_n3358 & ~new_n3397;
  assign new_n3399 = ~new_n3351 & ~new_n3352;
  assign new_n3400 = ~new_n3353 & ~new_n3399;
  assign new_n3401 = ~new_n1458 & ~new_n3400;
  assign new_n3402 = new_n1458 & new_n3400;
  assign new_n3403 = ~new_n3206 & ~new_n3207;
  assign new_n3404 = ~new_n3208 & ~new_n3403;
  assign new_n3405 = ~new_n3402 & ~new_n3404;
  assign new_n3406 = ~new_n3401 & ~new_n3405;
  assign new_n3407 = new_n3398 & new_n3406;
  assign new_n3408 = ~new_n3398 & ~new_n3406;
  assign new_n3409_1 = ~new_n3208 & ~new_n3212;
  assign new_n3410 = ~new_n3213 & ~new_n3409_1;
  assign new_n3411 = ~new_n3408 & new_n3410;
  assign new_n3412 = ~new_n3407 & ~new_n3411;
  assign new_n3413 = ~new_n3396 & ~new_n3412;
  assign new_n3414 = ~new_n3395 & ~new_n3413;
  assign new_n3415 = ~new_n3390 & ~new_n3414;
  assign new_n3416 = ~new_n3389 & ~new_n3415;
  assign new_n3417 = ~new_n3384 & new_n3416;
  assign new_n3418 = ~new_n3383 & ~new_n3417;
  assign new_n3419 = ~new_n3378 & new_n3418;
  assign new_n3420 = new_n3378 & ~new_n3418;
  assign new_n3421 = ~new_n3419 & ~new_n3420;
  assign new_n3422 = ~new_n3106 & new_n3421;
  assign new_n3423 = new_n3106 & ~new_n3421;
  assign new_n3424 = ~new_n3422 & ~new_n3423;
  assign new_n3425 = ~new_n3066 & ~new_n3068;
  assign new_n3426 = ~new_n3069 & ~new_n3425;
  assign new_n3427 = ~new_n3062 & ~new_n3065;
  assign new_n3428 = ~new_n3066 & ~new_n3427;
  assign new_n3429 = ~new_n3389 & ~new_n3390;
  assign new_n3430 = new_n3414 & ~new_n3429;
  assign new_n3431 = ~new_n3414 & new_n3429;
  assign new_n3432 = ~new_n3430 & ~new_n3431;
  assign new_n3433 = ~new_n3428 & ~new_n3432;
  assign new_n3434 = new_n3428 & new_n3432;
  assign new_n3435 = ~new_n3395 & ~new_n3396;
  assign new_n3436 = new_n3412 & ~new_n3435;
  assign new_n3437 = ~new_n3412 & new_n3435;
  assign new_n3438 = ~new_n3436 & ~new_n3437;
  assign new_n3439 = new_n3031 & new_n3073;
  assign new_n3440 = ~n12003 & ~new_n3073;
  assign new_n3441 = ~new_n3439 & ~new_n3440;
  assign new_n3442 = ~new_n3438 & new_n3441;
  assign new_n3443 = new_n3438 & ~new_n3441;
  assign new_n3444 = new_n3018 & new_n3073;
  assign new_n3445 = ~n10560 & ~new_n3073;
  assign new_n3446 = ~new_n3444 & ~new_n3445;
  assign new_n3447 = ~new_n3407 & ~new_n3408;
  assign new_n3448 = ~new_n3410 & ~new_n3447;
  assign new_n3449 = new_n3410 & new_n3447;
  assign new_n3450 = ~new_n3448 & ~new_n3449;
  assign new_n3451 = new_n3446 & ~new_n3450;
  assign new_n3452 = ~new_n3446 & new_n3450;
  assign new_n3453 = ~new_n1461 & ~new_n3074;
  assign new_n3454 = ~n10908 & new_n1461;
  assign new_n3455 = ~new_n3401 & ~new_n3402;
  assign new_n3456 = new_n3404 & ~new_n3455;
  assign new_n3457 = ~new_n3404 & new_n3455;
  assign new_n3458 = ~new_n3456 & ~new_n3457;
  assign new_n3459 = ~new_n3454 & new_n3458;
  assign new_n3460 = ~new_n3453 & ~new_n3459;
  assign new_n3461 = ~new_n3452 & ~new_n3460;
  assign new_n3462 = ~new_n3451 & ~new_n3461;
  assign new_n3463 = ~new_n3443 & ~new_n3462;
  assign new_n3464 = ~new_n3442 & ~new_n3463;
  assign new_n3465 = ~new_n3434 & ~new_n3464;
  assign new_n3466 = ~new_n3433 & ~new_n3465;
  assign new_n3467 = new_n3426 & new_n3466;
  assign new_n3468 = ~new_n3426 & ~new_n3466;
  assign new_n3469 = ~new_n3383 & ~new_n3384;
  assign new_n3470 = ~new_n3416 & ~new_n3469;
  assign new_n3471 = ~new_n3383 & new_n3417;
  assign new_n3472 = ~new_n3470 & ~new_n3471;
  assign new_n3473 = ~new_n3468 & ~new_n3472;
  assign new_n3474 = ~new_n3467 & ~new_n3473;
  assign new_n3475 = ~new_n3424 & new_n3474;
  assign new_n3476 = new_n3424 & ~new_n3474;
  assign new_n3477 = ~new_n3475 & ~new_n3476;
  assign new_n3478 = new_n3017 & new_n3477;
  assign new_n3479 = ~new_n3017 & ~new_n3477;
  assign new_n3480 = ~new_n3478 & ~new_n3479;
  assign new_n3481 = ~new_n3010 & ~new_n3012;
  assign new_n3482 = ~new_n3013 & ~new_n3481;
  assign new_n3483 = ~new_n3005 & ~new_n3009;
  assign new_n3484 = ~new_n3010 & ~new_n3483;
  assign new_n3485 = ~new_n3433 & ~new_n3434;
  assign new_n3486 = new_n3464 & ~new_n3485;
  assign new_n3487 = ~new_n3464 & new_n3485;
  assign new_n3488 = ~new_n3486 & ~new_n3487;
  assign new_n3489 = new_n3484 & ~new_n3488;
  assign new_n3490 = ~new_n3484 & new_n3488;
  assign new_n3491 = ~new_n3000 & new_n3004;
  assign new_n3492 = ~new_n3005 & ~new_n3491;
  assign new_n3493 = ~new_n3442 & ~new_n3443;
  assign new_n3494 = new_n3462 & ~new_n3493;
  assign new_n3495 = ~new_n3462 & new_n3493;
  assign new_n3496 = ~new_n3494 & ~new_n3495;
  assign new_n3497 = new_n3492 & ~new_n3496;
  assign new_n3498 = ~new_n3492 & new_n3496;
  assign new_n3499 = ~new_n2995 & ~new_n2999;
  assign new_n3500 = ~new_n3000 & ~new_n3499;
  assign new_n3501 = ~new_n3451 & ~new_n3452;
  assign new_n3502 = new_n3460 & ~new_n3501;
  assign new_n3503 = ~new_n3460 & new_n3501;
  assign new_n3504 = ~new_n3502 & ~new_n3503;
  assign new_n3505 = new_n3500 & ~new_n3504;
  assign new_n3506 = ~new_n3500 & new_n3504;
  assign new_n3507 = ~new_n3453 & ~new_n3454;
  assign new_n3508 = ~new_n3458 & ~new_n3507;
  assign new_n3509 = new_n3458 & new_n3507;
  assign new_n3510 = ~new_n3508 & ~new_n3509;
  assign new_n3511 = ~new_n1464 & new_n3510;
  assign new_n3512 = new_n1464 & ~new_n3510;
  assign new_n3513 = ~new_n2993 & ~new_n2994;
  assign new_n3514 = ~new_n2995 & ~new_n3513;
  assign new_n3515 = ~new_n3512 & ~new_n3514;
  assign new_n3516 = ~new_n3511 & ~new_n3515;
  assign new_n3517 = ~new_n3506 & new_n3516;
  assign new_n3518 = ~new_n3505 & ~new_n3517;
  assign new_n3519 = ~new_n3498 & ~new_n3518;
  assign new_n3520 = ~new_n3497 & ~new_n3519;
  assign new_n3521 = ~new_n3490 & ~new_n3520;
  assign new_n3522 = ~new_n3489 & ~new_n3521;
  assign new_n3523 = ~new_n3482 & new_n3522;
  assign new_n3524 = new_n3482 & ~new_n3522;
  assign new_n3525 = ~new_n3467 & ~new_n3468;
  assign new_n3526 = new_n3472 & ~new_n3525;
  assign new_n3527 = ~new_n3472 & new_n3525;
  assign new_n3528 = ~new_n3526 & ~new_n3527;
  assign new_n3529 = ~new_n3524 & ~new_n3528;
  assign new_n3530 = ~new_n3523 & ~new_n3529;
  assign new_n3531 = ~new_n3480 & new_n3530;
  assign new_n3532 = new_n3480 & ~new_n3530;
  assign n396 = new_n3531 | new_n3532;
  assign new_n3534 = ~new_n2987 & ~new_n3016;
  assign new_n3535 = n8290 & n12605;
  assign new_n3536 = new_n3197 & ~new_n3535;
  assign new_n3537 = ~new_n3197 & new_n3535;
  assign new_n3538 = ~new_n3536 & ~new_n3537;
  assign new_n3539 = n937 & n9591;
  assign new_n3540 = n4114 & n6023;
  assign new_n3541 = new_n3539 & ~new_n3540;
  assign new_n3542 = ~new_n3539 & new_n3540;
  assign new_n3543 = ~new_n3541 & ~new_n3542;
  assign new_n3544 = n510 & n5167;
  assign new_n3545 = n11665 & n12579;
  assign new_n3546 = new_n3544 & new_n3545;
  assign new_n3547 = ~new_n3544 & ~new_n3545;
  assign new_n3548 = ~new_n3546 & ~new_n3547;
  assign new_n3549 = new_n3543 & ~new_n3548;
  assign new_n3550 = ~new_n3543 & new_n3548;
  assign new_n3551 = ~new_n3549 & ~new_n3550;
  assign new_n3552 = new_n3165 & ~new_n3168;
  assign new_n3553 = ~new_n3169 & ~new_n3552;
  assign new_n3554 = ~new_n3551 & new_n3553;
  assign new_n3555 = new_n3551 & ~new_n3553;
  assign new_n3556 = ~new_n3554 & ~new_n3555;
  assign new_n3557 = n2666 & n5671;
  assign new_n3558 = n2777 & n11222;
  assign new_n3559 = ~new_n3557 & new_n3558;
  assign new_n3560 = new_n3557 & ~new_n3558;
  assign new_n3561 = ~new_n3559 & ~new_n3560;
  assign new_n3562 = new_n3175 & new_n3561;
  assign new_n3563 = ~new_n3175 & ~new_n3561;
  assign new_n3564 = ~new_n3562 & ~new_n3563;
  assign new_n3565 = new_n3556 & ~new_n3564;
  assign new_n3566 = ~new_n3556 & new_n3564;
  assign new_n3567 = ~new_n3565 & ~new_n3566;
  assign new_n3568 = ~new_n3538 & ~new_n3567;
  assign new_n3569 = new_n3538 & new_n3567;
  assign new_n3570 = ~new_n3568 & ~new_n3569;
  assign new_n3571 = ~new_n2945 & new_n2982;
  assign new_n3572 = ~new_n2946 & ~new_n3571;
  assign new_n3573 = n6168 & n11891;
  assign new_n3574 = n5214 & n9528;
  assign new_n3575 = ~new_n3573 & ~new_n3574;
  assign new_n3576 = new_n3573 & new_n3574;
  assign new_n3577 = ~new_n3575 & ~new_n3576;
  assign new_n3578 = n9531 & n11411;
  assign new_n3579 = n3006 & n5427;
  assign new_n3580 = ~new_n3578 & new_n3579;
  assign new_n3581 = new_n3578 & ~new_n3579;
  assign new_n3582 = ~new_n3580 & ~new_n3581;
  assign new_n3583 = ~new_n3577 & new_n3582;
  assign new_n3584 = new_n3577 & ~new_n3582;
  assign new_n3585 = ~new_n3583 & ~new_n3584;
  assign new_n3586 = n7061 & n12853;
  assign new_n3587 = n2771 & n9669;
  assign new_n3588 = n6655 & n8308;
  assign new_n3589 = new_n3587 & ~new_n3588;
  assign new_n3590 = ~new_n3587 & new_n3588;
  assign new_n3591_1 = ~new_n3589 & ~new_n3590;
  assign new_n3592 = new_n3586 & new_n3591_1;
  assign new_n3593 = ~new_n3586 & ~new_n3591_1;
  assign new_n3594 = ~new_n3592 & ~new_n3593;
  assign new_n3595 = new_n3585 & new_n3594;
  assign new_n3596 = ~new_n3585 & ~new_n3594;
  assign new_n3597 = ~new_n3595 & ~new_n3596;
  assign new_n3598 = new_n3572 & ~new_n3597;
  assign new_n3599 = ~new_n3572 & new_n3597;
  assign new_n3600 = ~new_n3598 & ~new_n3599;
  assign new_n3601 = new_n3176 & ~new_n3189;
  assign new_n3602 = ~new_n3188 & ~new_n3601;
  assign new_n3603 = ~new_n3600 & new_n3602;
  assign new_n3604 = new_n3600 & ~new_n3602;
  assign new_n3605 = ~new_n3603 & ~new_n3604;
  assign new_n3606 = ~new_n3570 & new_n3605;
  assign new_n3607 = new_n3570 & ~new_n3605;
  assign new_n3608 = ~new_n3606 & ~new_n3607;
  assign new_n3609 = new_n3534 & ~new_n3608;
  assign new_n3610 = ~new_n3534 & new_n3608;
  assign new_n3611 = ~new_n3609 & ~new_n3610;
  assign new_n3612 = new_n3177 & ~new_n3180;
  assign new_n3613 = ~new_n3181 & ~new_n3612;
  assign new_n3614 = ~new_n3422 & ~new_n3474;
  assign new_n3615 = ~new_n3423 & ~new_n3614;
  assign new_n3616 = ~new_n3613 & new_n3615;
  assign new_n3617 = new_n3613 & ~new_n3615;
  assign new_n3618 = ~new_n3616 & ~new_n3617;
  assign new_n3619 = ~new_n3098 & ~new_n3104;
  assign new_n3620 = ~new_n3101 & new_n3619;
  assign new_n3621 = ~new_n3080 & new_n3094;
  assign new_n3622 = ~new_n3081 & ~new_n3621;
  assign new_n3623 = new_n2948 & ~new_n2951;
  assign new_n3624 = ~new_n2952 & ~new_n3623;
  assign new_n3625 = ~new_n3622 & ~new_n3624;
  assign new_n3626 = new_n3622 & new_n3624;
  assign new_n3627 = ~new_n3625 & ~new_n3626;
  assign new_n3628 = n854 & n9041;
  assign new_n3629 = new_n3029 & ~new_n3628;
  assign new_n3630 = ~new_n3029 & new_n3628;
  assign new_n3631 = ~new_n3629 & ~new_n3630;
  assign new_n3632 = ~new_n3088 & ~new_n3089;
  assign new_n3633 = ~new_n3090 & ~new_n3632;
  assign new_n3634 = new_n3631 & new_n3633;
  assign new_n3635 = ~new_n3631 & ~new_n3633;
  assign new_n3636 = ~new_n3634 & ~new_n3635;
  assign new_n3637 = ~new_n3083 & ~new_n3085_1;
  assign new_n3638 = ~new_n3075 & ~new_n3637;
  assign new_n3639 = ~new_n3063 & ~new_n3638;
  assign new_n3640 = new_n3063 & new_n3638;
  assign new_n3641_1 = ~new_n3639 & ~new_n3640;
  assign new_n3642 = n389 & n5801;
  assign new_n3643 = new_n3088 & new_n3642;
  assign new_n3644 = ~new_n3088 & ~new_n3642;
  assign new_n3645 = ~new_n3643 & ~new_n3644;
  assign new_n3646 = new_n3641_1 & ~new_n3645;
  assign new_n3647 = ~new_n3641_1 & new_n3645;
  assign new_n3648 = ~new_n3646 & ~new_n3647;
  assign new_n3649 = ~new_n3636 & new_n3648;
  assign new_n3650 = new_n3636 & ~new_n3648;
  assign new_n3651 = ~new_n3649 & ~new_n3650;
  assign new_n3652 = ~new_n3627 & ~new_n3651;
  assign new_n3653 = new_n3627 & new_n3651;
  assign new_n3654 = ~new_n3652 & ~new_n3653;
  assign new_n3655 = ~new_n2962 & new_n2972;
  assign new_n3656 = ~new_n2961 & ~new_n3655;
  assign new_n3657 = n5568 & n8522;
  assign new_n3658 = new_n2964 & ~new_n2967;
  assign new_n3659 = ~new_n2968 & ~new_n3658;
  assign new_n3660 = ~new_n3657 & new_n3659;
  assign new_n3661 = new_n3657 & ~new_n3659;
  assign new_n3662 = ~new_n3660 & ~new_n3661;
  assign new_n3663 = new_n3656 & ~new_n3662;
  assign new_n3664 = ~new_n3656 & new_n3662;
  assign new_n3665 = ~new_n3663 & ~new_n3664;
  assign new_n3666 = new_n2980 & ~new_n3665;
  assign new_n3667 = ~new_n2980 & new_n3665;
  assign new_n3668 = ~new_n3666 & ~new_n3667;
  assign new_n3669_1 = ~new_n3654 & new_n3668;
  assign new_n3670 = new_n3654 & ~new_n3668;
  assign new_n3671 = ~new_n3669_1 & ~new_n3670;
  assign new_n3672 = new_n3620 & ~new_n3671;
  assign new_n3673 = ~new_n3620 & new_n3671;
  assign new_n3674 = ~new_n3672 & ~new_n3673;
  assign new_n3675 = ~new_n3377 & new_n3418;
  assign new_n3676 = ~new_n3376 & ~new_n3675;
  assign new_n3677_1 = ~new_n3674 & new_n3676;
  assign new_n3678 = new_n3674 & ~new_n3676;
  assign new_n3679 = ~new_n3677_1 & ~new_n3678;
  assign new_n3680 = ~new_n3200 & ~new_n3227;
  assign new_n3681 = n2057 & n2341;
  assign new_n3682 = n1650 & n5586;
  assign new_n3683 = ~new_n3319 & new_n3330;
  assign new_n3684 = ~new_n3320 & ~new_n3683;
  assign new_n3685 = new_n3682 & ~new_n3684;
  assign new_n3686 = ~new_n3682 & new_n3684;
  assign new_n3687 = ~new_n3685 & ~new_n3686;
  assign new_n3688 = n2295 & n4141;
  assign new_n3689 = ~new_n3322 & ~new_n3326;
  assign new_n3690 = ~new_n3325 & ~new_n3689;
  assign new_n3691 = new_n3306 & ~new_n3309;
  assign new_n3692 = ~new_n3310 & ~new_n3691;
  assign new_n3693 = ~new_n3690 & new_n3692;
  assign new_n3694 = new_n3690 & ~new_n3692;
  assign new_n3695 = ~new_n3693 & ~new_n3694;
  assign new_n3696 = new_n3688 & new_n3695;
  assign new_n3697 = ~new_n3688 & ~new_n3695;
  assign new_n3698 = ~new_n3696 & ~new_n3697;
  assign new_n3699 = new_n3337 & ~new_n3698;
  assign new_n3700 = ~new_n3337 & new_n3698;
  assign new_n3701 = ~new_n3699 & ~new_n3700;
  assign new_n3702 = ~new_n3687 & ~new_n3701;
  assign new_n3703 = new_n3687 & new_n3701;
  assign new_n3704 = ~new_n3702 & ~new_n3703;
  assign new_n3705 = ~new_n3681 & new_n3704;
  assign new_n3706 = new_n3681 & ~new_n3704;
  assign new_n3707 = ~new_n3705 & ~new_n3706;
  assign new_n3708 = ~new_n3680 & new_n3707;
  assign new_n3709 = new_n3680 & ~new_n3707;
  assign new_n3710 = ~new_n3708 & ~new_n3709;
  assign new_n3711 = ~new_n3345 & ~new_n3374;
  assign new_n3712 = ~new_n3303 & ~new_n3340;
  assign new_n3713 = ~new_n3304 & ~new_n3712;
  assign new_n3714 = n834 & n6409;
  assign new_n3715 = n5470 & n8716;
  assign new_n3716 = n12693 & n13201;
  assign new_n3717 = ~new_n3715 & ~new_n3716;
  assign new_n3718 = new_n3715 & new_n3716;
  assign new_n3719 = ~new_n3717 & ~new_n3718;
  assign new_n3720 = n3669 & n5189;
  assign new_n3721 = n1364 & n13060;
  assign new_n3722 = new_n3720 & ~new_n3721;
  assign new_n3723 = ~new_n3720 & new_n3721;
  assign new_n3724 = ~new_n3722 & ~new_n3723;
  assign new_n3725 = ~new_n3719 & ~new_n3724;
  assign new_n3726 = new_n3719 & new_n3724;
  assign new_n3727 = ~new_n3725 & ~new_n3726;
  assign new_n3728 = ~new_n3714 & new_n3727;
  assign new_n3729 = new_n3714 & ~new_n3727;
  assign new_n3730 = ~new_n3728 & ~new_n3729;
  assign new_n3731 = new_n3713 & new_n3730;
  assign new_n3732 = ~new_n3713 & ~new_n3730;
  assign new_n3733 = ~new_n3731 & ~new_n3732;
  assign new_n3734 = new_n3711 & new_n3733;
  assign new_n3735 = ~new_n3711 & ~new_n3733;
  assign new_n3736 = ~new_n3734 & ~new_n3735;
  assign new_n3737 = new_n3710 & new_n3736;
  assign new_n3738 = ~new_n3710 & ~new_n3736;
  assign new_n3739 = ~new_n3737 & ~new_n3738;
  assign new_n3740 = new_n3679 & ~new_n3739;
  assign new_n3741 = ~new_n3679 & new_n3739;
  assign new_n3742 = ~new_n3740 & ~new_n3741;
  assign new_n3743 = ~new_n3618 & ~new_n3742;
  assign new_n3744 = new_n3618 & new_n3742;
  assign new_n3745 = ~new_n3743 & ~new_n3744;
  assign new_n3746 = ~new_n3478 & ~new_n3530;
  assign new_n3747 = ~new_n3479 & ~new_n3746;
  assign new_n3748_1 = new_n3745 & new_n3747;
  assign new_n3749 = ~new_n3745 & ~new_n3747;
  assign new_n3750 = ~new_n3748_1 & ~new_n3749;
  assign new_n3751 = ~new_n3611 & new_n3750;
  assign new_n3752 = new_n3611 & ~new_n3750;
  assign n460 = ~new_n3751 & ~new_n3752;
  assign new_n3754 = ~new_n2633 & ~new_n2634;
  assign new_n3755 = new_n2648 & new_n3754;
  assign new_n3756 = ~new_n2648 & ~new_n3754;
  assign n537 = ~new_n3755 & ~new_n3756;
  assign new_n3758 = n2482 & n10451;
  assign new_n3759 = n9353 & n11058;
  assign new_n3760 = n287 & n8940;
  assign new_n3761 = new_n3759 & new_n3760;
  assign new_n3762 = ~new_n3759 & ~new_n3760;
  assign new_n3763 = ~new_n3761 & ~new_n3762;
  assign new_n3764 = n5962 & n8228;
  assign new_n3765 = new_n3763 & new_n3764;
  assign new_n3766 = ~new_n3763 & ~new_n3764;
  assign new_n3767 = ~new_n3765 & ~new_n3766;
  assign new_n3768 = new_n3758 & new_n3767;
  assign new_n3769_1 = ~new_n3758 & ~new_n3767;
  assign n573 = ~new_n3768 & ~new_n3769_1;
  assign new_n3771 = ~new_n1956 & ~new_n2002;
  assign new_n3772 = ~new_n1957 & ~new_n3771;
  assign new_n3773 = ~new_n1547 & new_n1551;
  assign new_n3774 = ~new_n1531 & ~new_n3773;
  assign new_n3775 = ~new_n1548 & new_n3774;
  assign new_n3776 = new_n1531 & new_n3773;
  assign new_n3777 = ~new_n3775 & ~new_n3776;
  assign new_n3778 = n4748 & n8308;
  assign new_n3779 = n1231 & n3006;
  assign new_n3780 = n5568 & n9187;
  assign new_n3781 = ~new_n3779 & ~new_n3780;
  assign new_n3782 = new_n3779 & new_n3780;
  assign new_n3783 = ~new_n3781 & ~new_n3782;
  assign new_n3784 = new_n3778 & ~new_n3783;
  assign new_n3785 = ~new_n3778 & new_n3783;
  assign new_n3786 = ~new_n3784 & ~new_n3785;
  assign new_n3787 = ~new_n1540 & ~new_n1543;
  assign new_n3788 = ~new_n1539 & ~new_n3787;
  assign new_n3789 = new_n3786 & ~new_n3788;
  assign new_n3790_1 = n5214 & n12306;
  assign new_n3791 = new_n1537 & new_n3790_1;
  assign new_n3792 = ~new_n1537 & ~new_n3790_1;
  assign new_n3793 = ~new_n3791 & ~new_n3792;
  assign new_n3794 = n4470 & n11411;
  assign new_n3795 = n2758 & n6168;
  assign new_n3796 = n2771 & n4006;
  assign new_n3797 = ~new_n3795 & ~new_n3796;
  assign new_n3798 = new_n3795 & new_n3796;
  assign new_n3799 = ~new_n3797 & ~new_n3798;
  assign new_n3800 = new_n3794 & ~new_n3799;
  assign new_n3801 = ~new_n3794 & new_n3799;
  assign new_n3802 = ~new_n3800 & ~new_n3801;
  assign new_n3803 = new_n3793 & new_n3802;
  assign new_n3804 = ~new_n3793 & ~new_n3802;
  assign new_n3805 = ~new_n3803 & ~new_n3804;
  assign new_n3806 = new_n3789 & new_n3805;
  assign new_n3807 = ~new_n3786 & new_n3788;
  assign new_n3808 = new_n3805 & ~new_n3807;
  assign new_n3809 = ~new_n3789 & ~new_n3808;
  assign new_n3810 = ~new_n3806 & ~new_n3809;
  assign new_n3811 = ~new_n3805 & new_n3807;
  assign new_n3812 = ~new_n3810 & ~new_n3811;
  assign new_n3813 = ~new_n3777 & new_n3812;
  assign new_n3814 = new_n3777 & ~new_n3812;
  assign new_n3815_1 = ~new_n3813 & ~new_n3814;
  assign new_n3816 = ~new_n1557 & ~new_n3815_1;
  assign new_n3817 = new_n1557 & new_n3815_1;
  assign new_n3818 = ~new_n3816 & ~new_n3817;
  assign new_n3819 = ~new_n1560 & ~new_n1563;
  assign new_n3820 = ~new_n3818 & new_n3819;
  assign new_n3821 = new_n3818 & ~new_n3819;
  assign new_n3822 = ~new_n3820 & ~new_n3821;
  assign new_n3823 = ~new_n1659 & ~new_n1663;
  assign new_n3824 = n6937 & n10560;
  assign new_n3825 = n5801 & n7729;
  assign new_n3826 = n3677 & n10908;
  assign new_n3827 = ~new_n3825 & ~new_n3826;
  assign new_n3828 = new_n3825 & new_n3826;
  assign new_n3829 = ~new_n3827 & ~new_n3828;
  assign new_n3830 = new_n3824 & ~new_n3829;
  assign new_n3831 = ~new_n3824 & new_n3829;
  assign new_n3832_1 = ~new_n3830 & ~new_n3831;
  assign new_n3833 = ~new_n1641 & new_n1644;
  assign new_n3834 = ~new_n1640 & ~new_n3833;
  assign new_n3835 = new_n3832_1 & ~new_n3834;
  assign new_n3836 = n1724 & n12003;
  assign new_n3837 = new_n1638 & new_n3836;
  assign new_n3838 = ~new_n1638 & ~new_n3836;
  assign new_n3839 = ~new_n3837 & ~new_n3838;
  assign new_n3840 = n10408 & ~n10866;
  assign new_n3841 = n3311 & n10606;
  assign new_n3842 = n8139 & n12965;
  assign new_n3843 = ~new_n3841 & ~new_n3842;
  assign new_n3844 = new_n3841 & new_n3842;
  assign new_n3845 = ~new_n3843 & ~new_n3844;
  assign new_n3846 = new_n3840 & ~new_n3845;
  assign new_n3847 = ~new_n3840 & new_n3845;
  assign new_n3848 = ~new_n3846 & ~new_n3847;
  assign new_n3849 = new_n3839 & new_n3848;
  assign new_n3850 = ~new_n3839 & ~new_n3848;
  assign new_n3851 = ~new_n3849 & ~new_n3850;
  assign new_n3852 = new_n3835 & new_n3851;
  assign new_n3853 = ~new_n3832_1 & new_n3834;
  assign new_n3854 = new_n3851 & ~new_n3853;
  assign new_n3855 = ~new_n3835 & ~new_n3854;
  assign new_n3856 = ~new_n3852 & ~new_n3855;
  assign new_n3857 = ~new_n3851 & new_n3853;
  assign new_n3858 = ~new_n3856 & ~new_n3857;
  assign new_n3859 = new_n1632 & ~new_n3858;
  assign new_n3860 = ~new_n1632 & new_n3858;
  assign new_n3861 = ~new_n3859 & ~new_n3860;
  assign new_n3862 = ~new_n1648 & new_n1652;
  assign new_n3863 = ~new_n1649 & ~new_n3862;
  assign new_n3864 = ~new_n3861 & new_n3863;
  assign new_n3865 = new_n3861 & ~new_n3863;
  assign new_n3866 = ~new_n3864 & ~new_n3865;
  assign new_n3867 = new_n1656 & new_n3866;
  assign new_n3868 = ~new_n1656 & ~new_n3866;
  assign new_n3869 = ~new_n3867 & ~new_n3868;
  assign new_n3870 = ~new_n3823 & new_n3869;
  assign new_n3871 = new_n3823 & ~new_n3869;
  assign new_n3872 = ~new_n3870 & ~new_n3871;
  assign new_n3873 = ~new_n1924 & ~new_n1928;
  assign new_n3874 = ~new_n1908 & ~new_n3873;
  assign new_n3875 = ~new_n1925 & new_n3874;
  assign new_n3876 = new_n1908 & new_n3873;
  assign new_n3877 = ~new_n3875 & ~new_n3876;
  assign new_n3878 = n2174 & n11665;
  assign new_n3879 = n4114 & new_n1902;
  assign new_n3880 = n3112 & n4114;
  assign new_n3881 = ~new_n1902 & ~new_n3880;
  assign new_n3882 = ~new_n3879 & ~new_n3881;
  assign new_n3883 = ~new_n3878 & new_n3882;
  assign new_n3884 = new_n3878 & ~new_n3882;
  assign new_n3885 = ~new_n3883 & ~new_n3884;
  assign new_n3886 = ~new_n1916_1 & new_n1920;
  assign new_n3887 = ~new_n1917 & ~new_n3886;
  assign new_n3888 = new_n3885 & ~new_n3887;
  assign new_n3889 = n497 & n2777;
  assign new_n3890 = new_n1914 & new_n3889;
  assign new_n3891 = ~new_n1914 & ~new_n3889;
  assign new_n3892 = ~new_n3890 & ~new_n3891;
  assign new_n3893 = n8233 & n12605;
  assign new_n3894 = n937 & n4335;
  assign new_n3895 = n9887 & n10642;
  assign new_n3896 = ~new_n3894 & ~new_n3895;
  assign new_n3897 = new_n3894 & new_n3895;
  assign new_n3898 = ~new_n3896 & ~new_n3897;
  assign new_n3899 = new_n3893 & ~new_n3898;
  assign new_n3900 = ~new_n3893 & new_n3898;
  assign new_n3901 = ~new_n3899 & ~new_n3900;
  assign new_n3902 = new_n3892 & new_n3901;
  assign new_n3903 = ~new_n3892 & ~new_n3901;
  assign new_n3904 = ~new_n3902 & ~new_n3903;
  assign new_n3905 = new_n3888 & new_n3904;
  assign new_n3906 = ~new_n3885 & new_n3887;
  assign new_n3907 = new_n3904 & ~new_n3906;
  assign new_n3908 = ~new_n3888 & ~new_n3907;
  assign new_n3909 = ~new_n3905 & ~new_n3908;
  assign new_n3910 = ~new_n3904 & new_n3906;
  assign new_n3911 = ~new_n3909 & ~new_n3910;
  assign new_n3912 = ~new_n3877 & new_n3911;
  assign new_n3913 = new_n3877 & ~new_n3911;
  assign new_n3914 = ~new_n3912 & ~new_n3913;
  assign new_n3915 = ~new_n1932 & ~new_n3914;
  assign new_n3916 = new_n1932 & new_n3914;
  assign new_n3917 = ~new_n3915 & ~new_n3916;
  assign new_n3918 = ~new_n1935 & ~new_n1939;
  assign new_n3919 = ~new_n3917 & new_n3918;
  assign new_n3920 = new_n3917 & ~new_n3918;
  assign new_n3921 = ~new_n3919 & ~new_n3920;
  assign new_n3922 = ~new_n1883 & ~new_n1887;
  assign new_n3923 = ~new_n1867 & ~new_n3922;
  assign new_n3924 = ~new_n1884 & new_n3923;
  assign new_n3925 = new_n1867 & new_n3922;
  assign new_n3926 = ~new_n3924 & ~new_n3925;
  assign new_n3927 = n2882 & n5586;
  assign new_n3928 = n1165 & n13201;
  assign new_n3929 = n2057 & n4357;
  assign new_n3930 = ~new_n3928 & ~new_n3929;
  assign new_n3931 = new_n3928 & new_n3929;
  assign new_n3932 = ~new_n3930 & ~new_n3931;
  assign new_n3933 = new_n3927 & ~new_n3932;
  assign new_n3934 = ~new_n3927 & new_n3932;
  assign new_n3935 = ~new_n3933 & ~new_n3934;
  assign new_n3936 = ~new_n1875 & new_n1879;
  assign new_n3937 = ~new_n1876 & ~new_n3936;
  assign new_n3938 = new_n3935 & ~new_n3937;
  assign new_n3939 = n3832 & n4141;
  assign new_n3940 = new_n1873 & new_n3939;
  assign new_n3941 = ~new_n1873 & ~new_n3939;
  assign new_n3942 = ~new_n3940 & ~new_n3941;
  assign new_n3943 = n5470 & n10063;
  assign new_n3944 = n3669 & n9915;
  assign new_n3945 = n1364 & n8332;
  assign new_n3946_1 = ~new_n3944 & ~new_n3945;
  assign new_n3947 = new_n3944 & new_n3945;
  assign new_n3948 = ~new_n3946_1 & ~new_n3947;
  assign new_n3949 = new_n3943 & ~new_n3948;
  assign new_n3950 = ~new_n3943 & new_n3948;
  assign new_n3951 = ~new_n3949 & ~new_n3950;
  assign new_n3952 = new_n3942 & new_n3951;
  assign new_n3953 = ~new_n3942 & ~new_n3951;
  assign new_n3954 = ~new_n3952 & ~new_n3953;
  assign new_n3955 = new_n3938 & new_n3954;
  assign new_n3956 = ~new_n3935 & new_n3937;
  assign new_n3957 = new_n3954 & ~new_n3956;
  assign new_n3958 = ~new_n3938 & ~new_n3957;
  assign new_n3959 = ~new_n3955 & ~new_n3958;
  assign new_n3960 = ~new_n3954 & new_n3956;
  assign new_n3961 = ~new_n3959 & ~new_n3960;
  assign new_n3962 = ~new_n3926 & new_n3961;
  assign new_n3963 = new_n3926 & ~new_n3961;
  assign new_n3964 = ~new_n3962 & ~new_n3963;
  assign new_n3965 = ~new_n1893 & ~new_n3964;
  assign new_n3966 = new_n1893 & new_n3964;
  assign new_n3967 = ~new_n3965 & ~new_n3966;
  assign new_n3968 = ~new_n1896 & ~new_n1900;
  assign new_n3969 = ~new_n3967 & new_n3968;
  assign new_n3970 = new_n3967 & ~new_n3968;
  assign new_n3971 = ~new_n3969 & ~new_n3970;
  assign new_n3972 = ~new_n3921 & ~new_n3971;
  assign new_n3973 = ~new_n1942 & ~new_n1945;
  assign new_n3974 = ~new_n1941 & ~new_n3973;
  assign new_n3975 = new_n3972 & new_n3974;
  assign new_n3976 = new_n3921 & new_n3971;
  assign new_n3977 = ~new_n3974 & new_n3976;
  assign new_n3978 = ~new_n3972 & ~new_n3974;
  assign new_n3979 = ~new_n3976 & ~new_n3978;
  assign new_n3980 = ~new_n3977 & ~new_n3979;
  assign new_n3981 = ~new_n3975 & ~new_n3980;
  assign new_n3982 = new_n3872 & new_n3981;
  assign new_n3983 = ~new_n3872 & ~new_n3981;
  assign new_n3984 = ~new_n3982 & ~new_n3983;
  assign new_n3985 = ~new_n1953 & new_n3984;
  assign new_n3986 = new_n1953 & ~new_n3984;
  assign new_n3987 = ~new_n3985 & ~new_n3986;
  assign new_n3988 = ~new_n3822 & ~new_n3987;
  assign new_n3989 = new_n3822 & new_n3987;
  assign new_n3990 = ~new_n3988 & ~new_n3989;
  assign new_n3991 = new_n3772 & new_n3990;
  assign new_n3992 = ~new_n3772 & ~new_n3990;
  assign n728 = new_n3991 | new_n3992;
  assign new_n3994 = n2482 & n12289;
  assign new_n3995 = n5729 & n10113;
  assign new_n3996 = new_n3994 & new_n3995;
  assign new_n3997 = n1757 & n5729;
  assign new_n3998 = n10113 & n12289;
  assign new_n3999 = n2482 & n7659;
  assign new_n4000 = ~new_n3998 & ~new_n3999;
  assign new_n4001 = new_n3998 & new_n3999;
  assign new_n4002 = ~new_n4000 & ~new_n4001;
  assign new_n4003 = new_n3997 & ~new_n4002;
  assign new_n4004 = ~new_n3997 & new_n4002;
  assign new_n4005 = ~new_n4003 & ~new_n4004;
  assign new_n4006_1 = ~new_n3996 & new_n4005;
  assign new_n4007 = new_n3996 & ~new_n4005;
  assign new_n4008 = ~new_n4006_1 & ~new_n4007;
  assign new_n4009 = ~new_n3994 & ~new_n3995;
  assign new_n4010 = ~new_n3996 & ~new_n4009;
  assign new_n4011 = n2482 & n5729;
  assign new_n4012 = n8228 & n13058;
  assign new_n4013 = n3769 & n8940;
  assign new_n4014 = n5548 & n9353;
  assign new_n4015 = new_n4013 & new_n4014;
  assign new_n4016 = ~new_n4013 & ~new_n4014;
  assign new_n4017 = ~new_n4015 & ~new_n4016;
  assign new_n4018 = new_n4012 & new_n4017;
  assign new_n4019 = ~new_n4012 & ~new_n4017;
  assign new_n4020 = ~new_n4018 & ~new_n4019;
  assign new_n4021 = new_n4011 & new_n4020;
  assign new_n4022 = ~new_n4010 & ~new_n4021;
  assign new_n4023 = new_n4010 & new_n4021;
  assign new_n4024 = n11236 & n13058;
  assign new_n4025 = n5920 & n8228;
  assign new_n4026 = ~new_n4024 & ~new_n4025;
  assign new_n4027 = new_n4024 & new_n4025;
  assign new_n4028 = ~new_n4026 & ~new_n4027;
  assign new_n4029 = n5548 & n6333;
  assign new_n4030 = n3815 & n9353;
  assign new_n4031 = ~new_n4029 & ~new_n4030;
  assign new_n4032 = new_n4029 & new_n4030;
  assign new_n4033 = ~new_n4031 & ~new_n4032;
  assign new_n4034 = n3769 & n4964;
  assign new_n4035 = n6392 & n8940;
  assign new_n4036 = ~new_n4034 & ~new_n4035;
  assign new_n4037 = new_n4034 & new_n4035;
  assign new_n4038 = ~new_n4036 & ~new_n4037;
  assign new_n4039 = ~new_n4015 & ~new_n4038;
  assign new_n4040 = new_n4015 & new_n4038;
  assign new_n4041 = ~new_n4039 & ~new_n4040;
  assign new_n4042 = ~new_n4033 & new_n4041;
  assign new_n4043 = new_n4033 & ~new_n4041;
  assign new_n4044 = ~new_n4042 & ~new_n4043;
  assign new_n4045 = ~new_n4028 & new_n4044;
  assign new_n4046 = new_n4028 & ~new_n4044;
  assign new_n4047 = ~new_n4045 & ~new_n4046;
  assign new_n4048 = ~new_n4018 & ~new_n4047;
  assign new_n4049 = new_n4018 & new_n4047;
  assign new_n4050 = ~new_n4048 & ~new_n4049;
  assign new_n4051 = ~new_n4023 & ~new_n4050;
  assign new_n4052 = ~new_n4022 & ~new_n4051;
  assign new_n4053 = new_n4008 & new_n4052;
  assign new_n4054 = n4382 & n13058;
  assign new_n4055 = n5920 & n11236;
  assign new_n4056 = n4862 & n8228;
  assign new_n4057 = ~new_n4055 & ~new_n4056;
  assign new_n4058 = new_n4055 & new_n4056;
  assign new_n4059_1 = ~new_n4057 & ~new_n4058;
  assign new_n4060 = new_n4054 & ~new_n4059_1;
  assign new_n4061 = ~new_n4054 & new_n4059_1;
  assign new_n4062 = ~new_n4060 & ~new_n4061;
  assign new_n4063 = ~new_n4027 & new_n4062;
  assign new_n4064 = new_n4027 & ~new_n4062;
  assign new_n4065 = ~new_n4063 & ~new_n4064;
  assign new_n4066 = n3769 & n5684;
  assign new_n4067 = n4964 & n6392;
  assign new_n4068 = n8940 & n10162;
  assign new_n4069 = ~new_n4067 & ~new_n4068;
  assign new_n4070 = new_n4067 & new_n4068;
  assign new_n4071 = ~new_n4069 & ~new_n4070;
  assign new_n4072 = new_n4066 & ~new_n4071;
  assign new_n4073 = ~new_n4066 & new_n4071;
  assign new_n4074 = ~new_n4072 & ~new_n4073;
  assign new_n4075_1 = ~new_n4037 & new_n4074;
  assign new_n4076 = new_n4037 & ~new_n4074;
  assign new_n4077 = ~new_n4075_1 & ~new_n4076;
  assign new_n4078 = n1912 & n5548;
  assign new_n4079 = n3815 & n6333;
  assign new_n4080 = n817 & n9353;
  assign new_n4081 = ~new_n4079 & ~new_n4080;
  assign new_n4082 = new_n4079 & new_n4080;
  assign new_n4083 = ~new_n4081 & ~new_n4082;
  assign new_n4084 = new_n4078 & ~new_n4083;
  assign new_n4085 = ~new_n4078 & new_n4083;
  assign new_n4086 = ~new_n4084 & ~new_n4085;
  assign new_n4087 = ~new_n4032 & new_n4086;
  assign new_n4088 = new_n4032 & ~new_n4086;
  assign new_n4089 = ~new_n4087 & ~new_n4088;
  assign new_n4090 = new_n4077 & new_n4089;
  assign new_n4091 = ~new_n4077 & ~new_n4089;
  assign new_n4092 = ~new_n4090 & ~new_n4091;
  assign new_n4093 = ~new_n4033 & ~new_n4040;
  assign new_n4094 = ~new_n4039 & ~new_n4093;
  assign new_n4095 = ~new_n4092 & new_n4094;
  assign new_n4096 = new_n4092 & ~new_n4094;
  assign new_n4097 = ~new_n4095 & ~new_n4096;
  assign new_n4098 = ~new_n4065 & new_n4097;
  assign new_n4099 = new_n4065 & ~new_n4097;
  assign new_n4100 = ~new_n4098 & ~new_n4099;
  assign new_n4101 = ~new_n4018 & ~new_n4046;
  assign new_n4102 = ~new_n4045 & ~new_n4101;
  assign new_n4103 = new_n4100 & new_n4102;
  assign new_n4104 = ~new_n4100 & ~new_n4102;
  assign new_n4105 = ~new_n4103 & ~new_n4104;
  assign new_n4106 = new_n4053 & new_n4105;
  assign new_n4107 = ~new_n4008 & ~new_n4052;
  assign new_n4108 = new_n4105 & ~new_n4107;
  assign new_n4109 = ~new_n4053 & ~new_n4108;
  assign new_n4110 = ~new_n4106 & ~new_n4109;
  assign new_n4111 = ~new_n4105 & new_n4107;
  assign n758 = ~new_n4110 & ~new_n4111;
  assign new_n4113 = n3769 & n8466;
  assign new_n4114_1 = n3178 & n5548;
  assign new_n4115 = new_n4113 & new_n4114_1;
  assign new_n4116 = ~new_n4113 & ~new_n4114_1;
  assign new_n4117 = ~new_n4115 & ~new_n4116;
  assign new_n4118 = n9216 & n13058;
  assign new_n4119 = new_n4117 & new_n4118;
  assign new_n4120 = ~new_n4117 & ~new_n4118;
  assign new_n4121 = ~new_n4119 & ~new_n4120;
  assign new_n4122_1 = n5729 & n7772;
  assign new_n4123 = new_n4121 & new_n4122_1;
  assign new_n4124 = n7772 & n12289;
  assign new_n4125 = n5729 & n7529;
  assign new_n4126 = ~new_n4124 & ~new_n4125;
  assign new_n4127 = new_n4124 & new_n4125;
  assign new_n4128 = ~new_n4126 & ~new_n4127;
  assign new_n4129 = ~new_n4123 & ~new_n4128;
  assign new_n4130 = new_n4123 & new_n4128;
  assign new_n4131 = ~new_n4129 & ~new_n4130;
  assign new_n4132 = n12348 & n13058;
  assign new_n4133 = n5920 & n9216;
  assign new_n4134 = ~new_n4132 & ~new_n4133;
  assign new_n4135 = new_n4132 & new_n4133;
  assign new_n4136 = ~new_n4134 & ~new_n4135;
  assign new_n4137 = n6392 & n8466;
  assign new_n4138 = n3769 & n5031;
  assign new_n4139 = ~new_n4137 & ~new_n4138;
  assign new_n4140 = new_n4137 & new_n4138;
  assign new_n4141_1 = ~new_n4139 & ~new_n4140;
  assign new_n4142 = ~new_n4115 & ~new_n4141_1;
  assign new_n4143 = new_n4115 & new_n4141_1;
  assign new_n4144 = ~new_n4142 & ~new_n4143;
  assign new_n4145 = n3178 & n3815;
  assign new_n4146 = n5548 & n12592;
  assign new_n4147 = ~new_n4145 & ~new_n4146;
  assign new_n4148 = new_n4145 & new_n4146;
  assign new_n4149 = ~new_n4147 & ~new_n4148;
  assign new_n4150 = ~new_n4144 & new_n4149;
  assign new_n4151 = ~new_n4143 & ~new_n4149;
  assign new_n4152 = ~new_n4142 & new_n4151;
  assign new_n4153 = ~new_n4150 & ~new_n4152;
  assign new_n4154 = new_n4136 & ~new_n4153;
  assign new_n4155 = ~new_n4136 & new_n4153;
  assign new_n4156 = ~new_n4154 & ~new_n4155;
  assign new_n4157 = ~new_n4119 & new_n4156;
  assign new_n4158 = new_n4119 & ~new_n4156;
  assign new_n4159 = ~new_n4157 & ~new_n4158;
  assign new_n4160 = new_n4131 & ~new_n4159;
  assign new_n4161 = ~new_n4131 & new_n4159;
  assign n762 = ~new_n4160 & ~new_n4161;
  assign new_n4163 = ~new_n4121 & ~new_n4122_1;
  assign n777 = ~new_n4123 & ~new_n4163;
  assign new_n4165 = ~new_n3523 & ~new_n3524;
  assign new_n4166 = ~new_n3528 & new_n4165;
  assign new_n4167 = new_n3528 & ~new_n4165;
  assign n800 = new_n4166 | new_n4167;
  assign new_n4169 = n4330 & n8308;
  assign new_n4170 = n2252 & n5568;
  assign new_n4171 = ~new_n4169 & ~new_n4170;
  assign new_n4172 = new_n4169 & new_n4170;
  assign new_n4173 = ~new_n4171 & ~new_n4172;
  assign new_n4174 = n5214 & n7659;
  assign new_n4175 = n2771 & n12289;
  assign new_n4176 = n5729 & n6168;
  assign new_n4177 = new_n4175 & new_n4176;
  assign new_n4178 = ~new_n4175 & ~new_n4176;
  assign new_n4179 = ~new_n4177 & ~new_n4178;
  assign new_n4180 = new_n4174 & new_n4179;
  assign new_n4181 = ~new_n4174 & ~new_n4179;
  assign new_n4182 = ~new_n4180 & ~new_n4181;
  assign new_n4183 = n5214 & n12289;
  assign new_n4184 = n7659 & n8308;
  assign new_n4185 = new_n4183 & new_n4184;
  assign new_n4186 = n2771 & n5729;
  assign new_n4187 = ~new_n4183 & ~new_n4184;
  assign new_n4188 = new_n4186 & ~new_n4187;
  assign new_n4189 = ~new_n4185 & ~new_n4188;
  assign new_n4190 = ~new_n4182 & ~new_n4189;
  assign new_n4191 = new_n4182 & new_n4189;
  assign new_n4192 = ~new_n4190 & ~new_n4191;
  assign new_n4193 = ~new_n4173 & new_n4192;
  assign new_n4194 = new_n4173 & ~new_n4192;
  assign new_n4195 = ~new_n4193 & ~new_n4194;
  assign new_n4196 = n4330 & n5568;
  assign new_n4197 = n8308 & n12289;
  assign new_n4198 = n5568 & n7659;
  assign new_n4199 = new_n4197 & new_n4198;
  assign new_n4200 = ~new_n4197 & ~new_n4198;
  assign new_n4201 = n5214 & n5729;
  assign new_n4202_1 = ~new_n4200 & new_n4201;
  assign new_n4203 = ~new_n4199 & ~new_n4202_1;
  assign new_n4204 = ~new_n4196 & new_n4203;
  assign new_n4205 = new_n4196 & ~new_n4203;
  assign new_n4206 = ~new_n4185 & ~new_n4187;
  assign new_n4207 = ~new_n4186 & ~new_n4206;
  assign new_n4208 = new_n4186 & new_n4206;
  assign new_n4209 = ~new_n4207 & ~new_n4208;
  assign new_n4210 = ~new_n4205 & ~new_n4209;
  assign new_n4211 = ~new_n4204 & ~new_n4210;
  assign new_n4212 = ~new_n4195 & new_n4211;
  assign new_n4213 = new_n4195 & ~new_n4211;
  assign new_n4214 = ~new_n4212 & ~new_n4213;
  assign new_n4215 = n2252 & n3006;
  assign new_n4216 = ~new_n4204 & ~new_n4205;
  assign new_n4217 = new_n4209 & ~new_n4216;
  assign new_n4218 = ~new_n4209 & new_n4216;
  assign new_n4219 = ~new_n4217 & ~new_n4218;
  assign new_n4220 = new_n4215 & ~new_n4219;
  assign new_n4221 = ~new_n4215 & new_n4219;
  assign new_n4222 = n3006 & n4330;
  assign new_n4223 = n5568 & n12289;
  assign new_n4224 = n3006 & n7659;
  assign new_n4225 = new_n4223 & new_n4224;
  assign new_n4226 = ~new_n4223 & ~new_n4224;
  assign new_n4227 = n5729 & n8308;
  assign new_n4228 = ~new_n4226 & new_n4227;
  assign new_n4229 = ~new_n4225 & ~new_n4228;
  assign new_n4230 = ~new_n4222 & new_n4229;
  assign new_n4231 = new_n4222 & ~new_n4229;
  assign new_n4232 = ~new_n4199 & ~new_n4200;
  assign new_n4233 = ~new_n4201 & ~new_n4232;
  assign new_n4234 = new_n4201 & new_n4232;
  assign new_n4235 = ~new_n4233 & ~new_n4234;
  assign new_n4236 = ~new_n4231 & ~new_n4235;
  assign new_n4237 = ~new_n4230 & ~new_n4236;
  assign new_n4238 = ~new_n4221 & new_n4237;
  assign new_n4239 = ~new_n4220 & ~new_n4238;
  assign new_n4240 = ~new_n4214 & ~new_n4239;
  assign new_n4241 = ~new_n4193 & new_n4211;
  assign new_n4242 = ~new_n4172 & ~new_n4241;
  assign new_n4243 = ~new_n4194 & new_n4242;
  assign new_n4244 = new_n4172 & new_n4241;
  assign new_n4245 = ~new_n4243 & ~new_n4244;
  assign new_n4246 = ~new_n4180 & new_n4189;
  assign new_n4247 = ~new_n4181 & ~new_n4246;
  assign new_n4248 = n2252 & n8308;
  assign new_n4249 = n5568 & n9747;
  assign new_n4250 = n3006 & n5884;
  assign new_n4251 = ~new_n4249 & ~new_n4250;
  assign new_n4252 = new_n4249 & new_n4250;
  assign new_n4253 = ~new_n4251 & ~new_n4252;
  assign new_n4254 = new_n4248 & ~new_n4253;
  assign new_n4255 = ~new_n4248 & new_n4253;
  assign new_n4256 = ~new_n4254 & ~new_n4255;
  assign new_n4257 = new_n4247 & ~new_n4256;
  assign new_n4258 = ~new_n4247 & new_n4256;
  assign new_n4259 = ~new_n4257 & ~new_n4258;
  assign new_n4260 = n4330 & n5214;
  assign new_n4261 = new_n4177 & new_n4260;
  assign new_n4262 = ~new_n4177 & ~new_n4260;
  assign new_n4263 = ~new_n4261 & ~new_n4262;
  assign new_n4264 = n5729 & n11411;
  assign new_n4265 = n6168 & n12289;
  assign new_n4266 = n2771 & n7659;
  assign new_n4267 = ~new_n4265 & ~new_n4266;
  assign new_n4268 = new_n4265 & new_n4266;
  assign new_n4269 = ~new_n4267 & ~new_n4268;
  assign new_n4270 = new_n4264 & ~new_n4269;
  assign new_n4271 = ~new_n4264 & new_n4269;
  assign new_n4272 = ~new_n4270 & ~new_n4271;
  assign new_n4273 = ~new_n4263 & ~new_n4272;
  assign new_n4274 = new_n4263 & new_n4272;
  assign new_n4275 = ~new_n4273 & ~new_n4274;
  assign new_n4276 = ~new_n4259 & new_n4275;
  assign new_n4277 = new_n4259 & ~new_n4275;
  assign new_n4278 = ~new_n4276 & ~new_n4277;
  assign new_n4279 = new_n4245 & new_n4278;
  assign new_n4280 = ~new_n4245 & ~new_n4278;
  assign new_n4281 = ~new_n4279 & ~new_n4280;
  assign new_n4282 = new_n4240 & new_n4281;
  assign new_n4283 = ~new_n4240 & ~new_n4281;
  assign new_n4284 = ~new_n4282 & ~new_n4283;
  assign new_n4285 = n3006 & n9747;
  assign new_n4286 = new_n4214 & new_n4239;
  assign new_n4287 = ~new_n4240 & ~new_n4286;
  assign new_n4288 = new_n4285 & new_n4287;
  assign new_n4289 = n3006 & n12289;
  assign new_n4290 = n5568 & n5729;
  assign new_n4291 = new_n4289 & new_n4290;
  assign new_n4292 = ~new_n4225 & ~new_n4226;
  assign new_n4293 = ~new_n4227 & ~new_n4292;
  assign new_n4294 = new_n4227 & new_n4292;
  assign new_n4295 = ~new_n4293 & ~new_n4294;
  assign new_n4296 = new_n4291 & new_n4295;
  assign new_n4297 = ~new_n4230 & ~new_n4231;
  assign new_n4298 = ~new_n4235 & ~new_n4297;
  assign new_n4299 = new_n4235 & new_n4297;
  assign new_n4300 = ~new_n4298 & ~new_n4299;
  assign new_n4301 = new_n4296 & new_n4300;
  assign new_n4302 = ~new_n4220 & ~new_n4221;
  assign new_n4303 = ~new_n4237 & ~new_n4302;
  assign new_n4304 = new_n4237 & new_n4302;
  assign new_n4305 = ~new_n4303 & ~new_n4304;
  assign new_n4306 = new_n4301 & new_n4305;
  assign new_n4307 = ~new_n4285 & ~new_n4287;
  assign new_n4308 = ~new_n4288 & ~new_n4307;
  assign new_n4309 = new_n4306 & new_n4308;
  assign new_n4310 = ~new_n4288 & ~new_n4309;
  assign new_n4311 = new_n4284 & ~new_n4310;
  assign new_n4312 = ~new_n4284 & new_n4310;
  assign new_n4313 = ~new_n4311 & ~new_n4312;
  assign new_n4314 = n443 & n5801;
  assign new_n4315 = n5065 & n5801;
  assign new_n4316 = n8139 & n13058;
  assign new_n4317 = n5920 & n12003;
  assign new_n4318 = n4862 & n10560;
  assign new_n4319 = ~new_n4317 & ~new_n4318;
  assign new_n4320 = new_n4317 & new_n4318;
  assign new_n4321 = ~new_n4319 & ~new_n4320;
  assign new_n4322 = ~new_n4316 & ~new_n4321;
  assign new_n4323 = new_n4316 & new_n4321;
  assign new_n4324 = ~new_n4322 & ~new_n4323;
  assign new_n4325 = n1636 & n10908;
  assign new_n4326 = n5920 & n10560;
  assign new_n4327 = n4862 & n10908;
  assign new_n4328 = new_n4326 & new_n4327;
  assign new_n4329 = ~new_n4326 & ~new_n4327;
  assign new_n4330_1 = n12003 & n13058;
  assign new_n4331 = ~new_n4329 & new_n4330_1;
  assign new_n4332 = ~new_n4328 & ~new_n4331;
  assign new_n4333 = new_n4325 & ~new_n4332;
  assign new_n4334 = ~new_n4325 & new_n4332;
  assign new_n4335_1 = ~new_n4333 & ~new_n4334;
  assign new_n4336 = ~new_n4324 & new_n4335_1;
  assign new_n4337 = new_n4324 & ~new_n4335_1;
  assign new_n4338 = ~new_n4336 & ~new_n4337;
  assign new_n4339 = new_n4315 & ~new_n4338;
  assign new_n4340 = ~new_n4315 & new_n4338;
  assign new_n4341 = n1636 & n5801;
  assign new_n4342 = n5920 & n10908;
  assign new_n4343 = n4862 & n5801;
  assign new_n4344 = new_n4342 & new_n4343;
  assign new_n4345 = ~new_n4342 & ~new_n4343;
  assign new_n4346 = n10560 & n13058;
  assign new_n4347 = ~new_n4345 & new_n4346;
  assign new_n4348 = ~new_n4344 & ~new_n4347;
  assign new_n4349 = ~new_n4341 & new_n4348;
  assign new_n4350 = new_n4341 & ~new_n4348;
  assign new_n4351 = ~new_n4328 & ~new_n4329;
  assign new_n4352 = ~new_n4330_1 & ~new_n4351;
  assign new_n4353 = new_n4330_1 & new_n4351;
  assign new_n4354 = ~new_n4352 & ~new_n4353;
  assign new_n4355 = ~new_n4350 & ~new_n4354;
  assign new_n4356 = ~new_n4349 & ~new_n4355;
  assign new_n4357_1 = ~new_n4340 & new_n4356;
  assign new_n4358 = ~new_n4339 & ~new_n4357_1;
  assign new_n4359 = new_n4324 & ~new_n4334;
  assign new_n4360 = ~new_n4333 & ~new_n4359;
  assign new_n4361 = n1636 & n10560;
  assign new_n4362 = n5065 & n10908;
  assign new_n4363 = new_n4361 & new_n4362;
  assign new_n4364 = ~new_n4361 & ~new_n4362;
  assign new_n4365 = ~new_n4363 & ~new_n4364;
  assign new_n4366 = n4862 & n12003;
  assign new_n4367 = n5920 & n8139;
  assign new_n4368 = n3311 & n13058;
  assign new_n4369 = new_n4367 & new_n4368;
  assign new_n4370 = ~new_n4367 & ~new_n4368;
  assign new_n4371 = ~new_n4369 & ~new_n4370;
  assign new_n4372 = ~new_n4366 & ~new_n4371;
  assign new_n4373 = new_n4366 & new_n4371;
  assign new_n4374 = ~new_n4372 & ~new_n4373;
  assign new_n4375 = new_n4316 & ~new_n4319;
  assign new_n4376 = ~new_n4320 & ~new_n4375;
  assign new_n4377 = ~new_n4374 & new_n4376;
  assign new_n4378 = new_n4374 & ~new_n4376;
  assign new_n4379 = ~new_n4377 & ~new_n4378;
  assign new_n4380 = ~new_n4365 & ~new_n4379;
  assign new_n4381 = new_n4365 & new_n4379;
  assign new_n4382_1 = ~new_n4380 & ~new_n4381;
  assign new_n4383 = ~new_n4360 & new_n4382_1;
  assign new_n4384 = new_n4360 & ~new_n4382_1;
  assign new_n4385 = ~new_n4383 & ~new_n4384;
  assign new_n4386 = ~new_n4358 & new_n4385;
  assign new_n4387 = new_n4358 & ~new_n4385;
  assign new_n4388 = ~new_n4386 & ~new_n4387;
  assign new_n4389 = new_n4314 & new_n4388;
  assign new_n4390 = n5801 & n5920;
  assign new_n4391 = n10908 & n13058;
  assign new_n4392 = new_n4390 & new_n4391;
  assign new_n4393 = ~new_n4344 & ~new_n4345;
  assign new_n4394 = ~new_n4346 & ~new_n4393;
  assign new_n4395 = new_n4346 & new_n4393;
  assign new_n4396 = ~new_n4394 & ~new_n4395;
  assign new_n4397 = new_n4392 & new_n4396;
  assign new_n4398 = ~new_n4349 & ~new_n4350;
  assign new_n4399 = ~new_n4354 & new_n4398;
  assign new_n4400 = new_n4354 & ~new_n4398;
  assign new_n4401 = ~new_n4399 & ~new_n4400;
  assign new_n4402 = new_n4397 & ~new_n4401;
  assign new_n4403 = ~new_n4339 & ~new_n4340;
  assign new_n4404 = ~new_n4356 & ~new_n4403;
  assign new_n4405 = new_n4356 & new_n4403;
  assign new_n4406 = ~new_n4404 & ~new_n4405;
  assign new_n4407 = new_n4402 & new_n4406;
  assign new_n4408 = ~new_n4314 & ~new_n4388;
  assign new_n4409 = ~new_n4389 & ~new_n4408;
  assign new_n4410 = new_n4407 & new_n4409;
  assign new_n4411 = ~new_n4389 & ~new_n4410;
  assign new_n4412 = ~n10866 & n13058;
  assign new_n4413 = n3311 & n5920;
  assign new_n4414 = n4862 & n8139;
  assign new_n4415 = ~new_n4413 & ~new_n4414;
  assign new_n4416 = new_n4413 & new_n4414;
  assign new_n4417 = ~new_n4415 & ~new_n4416;
  assign new_n4418 = ~new_n4412 & ~new_n4417;
  assign new_n4419_1 = new_n4412 & new_n4417;
  assign new_n4420 = ~new_n4418 & ~new_n4419_1;
  assign new_n4421 = n1636 & n12003;
  assign new_n4422 = new_n4369 & new_n4421;
  assign new_n4423 = ~new_n4369 & ~new_n4421;
  assign new_n4424 = ~new_n4422 & ~new_n4423;
  assign new_n4425 = ~new_n4420 & ~new_n4424;
  assign new_n4426 = new_n4420 & new_n4424;
  assign new_n4427 = ~new_n4425 & ~new_n4426;
  assign new_n4428 = ~new_n4372 & ~new_n4376;
  assign new_n4429 = ~new_n4373 & ~new_n4428;
  assign new_n4430 = n5065 & n10560;
  assign new_n4431 = n5801 & n11835;
  assign new_n4432 = n443 & n10908;
  assign new_n4433 = ~new_n4431 & ~new_n4432;
  assign new_n4434 = new_n4431 & new_n4432;
  assign new_n4435 = ~new_n4433 & ~new_n4434;
  assign new_n4436 = new_n4430 & ~new_n4435;
  assign new_n4437 = ~new_n4430 & new_n4435;
  assign new_n4438 = ~new_n4436 & ~new_n4437;
  assign new_n4439 = ~new_n4429 & ~new_n4438;
  assign new_n4440 = new_n4429 & new_n4438;
  assign new_n4441 = ~new_n4439 & ~new_n4440;
  assign new_n4442 = new_n4427 & ~new_n4441;
  assign new_n4443 = ~new_n4427 & ~new_n4439;
  assign new_n4444 = ~new_n4440 & new_n4443;
  assign new_n4445 = ~new_n4442 & ~new_n4444;
  assign new_n4446 = ~new_n4360 & ~new_n4380;
  assign new_n4447 = new_n4363 & new_n4446;
  assign new_n4448 = ~new_n4363 & ~new_n4446;
  assign new_n4449 = ~new_n4381 & new_n4448;
  assign new_n4450 = ~new_n4447 & ~new_n4449;
  assign new_n4451 = ~new_n4445 & new_n4450;
  assign new_n4452_1 = new_n4445 & ~new_n4450;
  assign new_n4453 = ~new_n4451 & ~new_n4452_1;
  assign new_n4454 = new_n4386 & new_n4453;
  assign new_n4455 = ~new_n4386 & ~new_n4453;
  assign new_n4456 = ~new_n4454 & ~new_n4455;
  assign new_n4457 = ~new_n4411 & new_n4456;
  assign new_n4458 = new_n4411 & ~new_n4456;
  assign new_n4459 = ~new_n4457 & ~new_n4458;
  assign new_n4460 = n8163 & n13201;
  assign new_n4461 = n5586 & n11634;
  assign new_n4462 = n2057 & n3076;
  assign new_n4463 = ~new_n4461 & ~new_n4462;
  assign new_n4464 = new_n4461 & new_n4462;
  assign new_n4465 = ~new_n4463 & ~new_n4464;
  assign new_n4466 = n1364 & n3815;
  assign new_n4467 = n3669 & n5548;
  assign new_n4468 = ~new_n4466 & ~new_n4467;
  assign new_n4469 = new_n4466 & new_n4467;
  assign new_n4470_1 = ~new_n4468 & ~new_n4469;
  assign new_n4471 = n817 & n4141;
  assign new_n4472 = ~new_n4470_1 & ~new_n4471;
  assign new_n4473 = new_n4470_1 & new_n4471;
  assign new_n4474 = ~new_n4472 & ~new_n4473;
  assign new_n4475 = n3815 & n4141;
  assign new_n4476 = n817 & n5586;
  assign new_n4477 = new_n4475 & new_n4476;
  assign new_n4478 = n1364 & n5548;
  assign new_n4479 = ~new_n4475 & ~new_n4476;
  assign new_n4480 = new_n4478 & ~new_n4479;
  assign new_n4481 = ~new_n4477 & ~new_n4480;
  assign new_n4482 = ~new_n4474 & ~new_n4481;
  assign new_n4483 = new_n4474 & new_n4481;
  assign new_n4484 = ~new_n4482 & ~new_n4483;
  assign new_n4485 = ~new_n4465 & new_n4484;
  assign new_n4486 = new_n4465 & ~new_n4484;
  assign new_n4487 = ~new_n4485 & ~new_n4486;
  assign new_n4488 = n2057 & n11634;
  assign new_n4489 = n3815 & n5586;
  assign new_n4490 = n817 & n2057;
  assign new_n4491 = new_n4489 & new_n4490;
  assign new_n4492 = ~new_n4489 & ~new_n4490;
  assign new_n4493 = n4141 & n5548;
  assign new_n4494 = ~new_n4492 & new_n4493;
  assign new_n4495 = ~new_n4491 & ~new_n4494;
  assign new_n4496 = ~new_n4488 & new_n4495;
  assign new_n4497 = new_n4488 & ~new_n4495;
  assign new_n4498 = ~new_n4477 & ~new_n4479;
  assign new_n4499 = ~new_n4478 & ~new_n4498;
  assign new_n4500 = new_n4478 & new_n4498;
  assign new_n4501 = ~new_n4499 & ~new_n4500;
  assign new_n4502 = ~new_n4497 & ~new_n4501;
  assign new_n4503 = ~new_n4496 & ~new_n4502;
  assign new_n4504 = ~new_n4487 & ~new_n4503;
  assign new_n4505 = new_n4487 & new_n4503;
  assign new_n4506 = ~new_n4504 & ~new_n4505;
  assign new_n4507 = n3076 & n13201;
  assign new_n4508 = ~new_n4496 & new_n4502;
  assign new_n4509 = ~new_n4496 & ~new_n4497;
  assign new_n4510 = new_n4501 & ~new_n4509;
  assign new_n4511 = ~new_n4508 & ~new_n4510;
  assign new_n4512 = new_n4507 & ~new_n4511;
  assign new_n4513 = ~new_n4507 & new_n4511;
  assign new_n4514 = n11634 & n13201;
  assign new_n4515 = n2057 & n3815;
  assign new_n4516 = n817 & n13201;
  assign new_n4517 = new_n4515 & new_n4516;
  assign new_n4518 = ~new_n4515 & ~new_n4516;
  assign new_n4519 = n5548 & n5586;
  assign new_n4520 = ~new_n4518 & new_n4519;
  assign new_n4521 = ~new_n4517 & ~new_n4520;
  assign new_n4522 = ~new_n4514 & new_n4521;
  assign new_n4523 = new_n4514 & ~new_n4521;
  assign new_n4524 = ~new_n4491 & ~new_n4492;
  assign new_n4525 = ~new_n4493 & ~new_n4524;
  assign new_n4526 = new_n4493 & new_n4524;
  assign new_n4527 = ~new_n4525 & ~new_n4526;
  assign new_n4528 = ~new_n4523 & ~new_n4527;
  assign new_n4529 = ~new_n4522 & ~new_n4528;
  assign new_n4530 = ~new_n4513 & new_n4529;
  assign new_n4531 = ~new_n4512 & ~new_n4530;
  assign new_n4532 = new_n4506 & ~new_n4531;
  assign new_n4533 = ~new_n4506 & new_n4531;
  assign new_n4534 = ~new_n4532 & ~new_n4533;
  assign new_n4535 = new_n4460 & new_n4534;
  assign new_n4536 = n3815 & n13201;
  assign new_n4537 = n2057 & n5548;
  assign new_n4538 = new_n4536 & new_n4537;
  assign new_n4539 = ~new_n4517 & ~new_n4518;
  assign new_n4540 = ~new_n4519 & ~new_n4539;
  assign new_n4541 = new_n4519 & new_n4539;
  assign new_n4542 = ~new_n4540 & ~new_n4541;
  assign new_n4543 = new_n4538 & new_n4542;
  assign new_n4544 = ~new_n4522 & ~new_n4523;
  assign new_n4545 = ~new_n4527 & new_n4544;
  assign new_n4546 = new_n4527 & ~new_n4544;
  assign new_n4547 = ~new_n4545 & ~new_n4546;
  assign new_n4548 = new_n4543 & ~new_n4547;
  assign new_n4549 = ~new_n4512 & ~new_n4513;
  assign new_n4550 = ~new_n4529 & ~new_n4549;
  assign new_n4551 = new_n4529 & new_n4549;
  assign new_n4552 = ~new_n4550 & ~new_n4551;
  assign new_n4553_1 = new_n4548 & new_n4552;
  assign new_n4554 = ~new_n4460 & ~new_n4534;
  assign new_n4555 = ~new_n4535 & ~new_n4554;
  assign new_n4556 = new_n4553_1 & new_n4555;
  assign new_n4557 = ~new_n4535 & ~new_n4556;
  assign new_n4558 = ~new_n4485 & new_n4503;
  assign new_n4559 = ~new_n4464 & ~new_n4558;
  assign new_n4560 = ~new_n4486 & new_n4559;
  assign new_n4561 = new_n4464 & new_n4558;
  assign new_n4562 = ~new_n4560 & ~new_n4561;
  assign new_n4563 = n3076 & n5586;
  assign new_n4564 = n7974 & n13201;
  assign new_n4565 = n2057 & n8163;
  assign new_n4566 = ~new_n4564 & ~new_n4565;
  assign new_n4567 = new_n4564 & new_n4565;
  assign new_n4568 = ~new_n4566 & ~new_n4567;
  assign new_n4569 = new_n4563 & ~new_n4568;
  assign new_n4570 = ~new_n4563 & new_n4568;
  assign new_n4571 = ~new_n4569 & ~new_n4570;
  assign new_n4572 = ~new_n4473 & new_n4481;
  assign new_n4573 = ~new_n4472 & ~new_n4572;
  assign new_n4574 = new_n4571 & ~new_n4573;
  assign new_n4575 = ~new_n4571 & new_n4573;
  assign new_n4576 = ~new_n4574 & ~new_n4575;
  assign new_n4577 = n4141 & n11634;
  assign new_n4578 = ~new_n4469 & ~new_n4577;
  assign new_n4579 = new_n4469 & new_n4577;
  assign new_n4580 = ~new_n4578 & ~new_n4579;
  assign new_n4581 = n5470 & n5548;
  assign new_n4582 = n3669 & n3815;
  assign new_n4583 = n817 & n1364;
  assign new_n4584 = ~new_n4582 & ~new_n4583;
  assign new_n4585 = new_n4582 & new_n4583;
  assign new_n4586 = ~new_n4584 & ~new_n4585;
  assign new_n4587 = new_n4581 & ~new_n4586;
  assign new_n4588 = ~new_n4581 & new_n4586;
  assign new_n4589 = ~new_n4587 & ~new_n4588;
  assign new_n4590 = ~new_n4580 & new_n4589;
  assign new_n4591 = new_n4580 & ~new_n4589;
  assign new_n4592 = ~new_n4590 & ~new_n4591;
  assign new_n4593 = ~new_n4576 & ~new_n4592;
  assign new_n4594 = new_n4576 & new_n4592;
  assign new_n4595 = ~new_n4593 & ~new_n4594;
  assign new_n4596 = new_n4562 & ~new_n4595;
  assign new_n4597 = ~new_n4562 & new_n4595;
  assign new_n4598 = ~new_n4596 & ~new_n4597;
  assign new_n4599 = new_n4532 & ~new_n4598;
  assign new_n4600 = ~new_n4532 & new_n4598;
  assign new_n4601 = ~new_n4599 & ~new_n4600;
  assign new_n4602 = ~new_n4557 & new_n4601;
  assign new_n4603 = new_n4557 & ~new_n4601;
  assign new_n4604 = ~new_n4602 & ~new_n4603;
  assign new_n4605 = n1916 & n4114;
  assign new_n4606 = n8860 & n11665;
  assign new_n4607 = ~new_n4605 & ~new_n4606;
  assign new_n4608 = new_n4605 & new_n4606;
  assign new_n4609 = ~new_n4607 & ~new_n4608;
  assign new_n4610 = n2777 & n10162;
  assign new_n4611 = n6392 & n10642;
  assign new_n4612 = n937 & n3769;
  assign new_n4613 = ~new_n4611 & ~new_n4612;
  assign new_n4614 = new_n4611 & new_n4612;
  assign new_n4615 = ~new_n4613 & ~new_n4614;
  assign new_n4616 = new_n4610 & new_n4615;
  assign new_n4617 = ~new_n4610 & ~new_n4615;
  assign new_n4618 = ~new_n4616 & ~new_n4617;
  assign new_n4619 = n10162 & n11665;
  assign new_n4620 = n2777 & n6392;
  assign new_n4621 = new_n4619 & new_n4620;
  assign new_n4622 = ~new_n4619 & ~new_n4620;
  assign new_n4623 = n3769 & n10642;
  assign new_n4624 = ~new_n4622 & new_n4623;
  assign new_n4625 = ~new_n4621 & ~new_n4624;
  assign new_n4626 = ~new_n4618 & ~new_n4625;
  assign new_n4627 = new_n4618 & new_n4625;
  assign new_n4628 = ~new_n4626 & ~new_n4627;
  assign new_n4629 = ~new_n4609 & new_n4628;
  assign new_n4630 = new_n4609 & ~new_n4628;
  assign new_n4631 = ~new_n4629 & ~new_n4630;
  assign new_n4632 = n4114 & n8860;
  assign new_n4633 = n6392 & n11665;
  assign new_n4634 = n4114 & n10162;
  assign new_n4635 = new_n4633 & new_n4634;
  assign new_n4636 = ~new_n4633 & ~new_n4634;
  assign new_n4637 = n2777 & n3769;
  assign new_n4638 = ~new_n4636 & new_n4637;
  assign new_n4639 = ~new_n4635 & ~new_n4638;
  assign new_n4640 = ~new_n4632 & new_n4639;
  assign new_n4641 = new_n4632 & ~new_n4639;
  assign new_n4642 = ~new_n4621 & ~new_n4622;
  assign new_n4643 = ~new_n4623 & ~new_n4642;
  assign new_n4644 = new_n4623 & new_n4642;
  assign new_n4645 = ~new_n4643 & ~new_n4644;
  assign new_n4646 = ~new_n4641 & ~new_n4645;
  assign new_n4647 = ~new_n4640 & ~new_n4646;
  assign new_n4648 = ~new_n4631 & new_n4647;
  assign new_n4649 = new_n4631 & ~new_n4647;
  assign new_n4650 = ~new_n4648 & ~new_n4649;
  assign new_n4651 = n1916 & n5671;
  assign new_n4652 = ~new_n4640 & ~new_n4641;
  assign new_n4653 = ~new_n4645 & ~new_n4652;
  assign new_n4654 = new_n4645 & new_n4652;
  assign new_n4655 = ~new_n4653 & ~new_n4654;
  assign new_n4656 = new_n4651 & new_n4655;
  assign new_n4657 = ~new_n4651 & ~new_n4655;
  assign new_n4658 = n5671 & n8860;
  assign new_n4659 = n4114 & n6392;
  assign new_n4660 = n5671 & n10162;
  assign new_n4661 = new_n4659 & new_n4660;
  assign new_n4662 = ~new_n4659 & ~new_n4660;
  assign new_n4663 = n3769 & n11665;
  assign new_n4664 = ~new_n4662 & new_n4663;
  assign new_n4665 = ~new_n4661 & ~new_n4664;
  assign new_n4666 = ~new_n4658 & new_n4665;
  assign new_n4667 = new_n4658 & ~new_n4665;
  assign new_n4668 = ~new_n4635 & ~new_n4636;
  assign new_n4669 = ~new_n4637 & ~new_n4668;
  assign new_n4670 = new_n4637 & new_n4668;
  assign new_n4671 = ~new_n4669 & ~new_n4670;
  assign new_n4672 = ~new_n4667 & ~new_n4671;
  assign new_n4673 = ~new_n4666 & ~new_n4672;
  assign new_n4674 = ~new_n4657 & new_n4673;
  assign new_n4675 = ~new_n4656 & ~new_n4674;
  assign new_n4676 = ~new_n4650 & ~new_n4675;
  assign new_n4677 = ~new_n4629 & new_n4647;
  assign new_n4678 = ~new_n4608 & ~new_n4677;
  assign new_n4679 = ~new_n4630 & new_n4678;
  assign new_n4680 = new_n4608 & new_n4677;
  assign new_n4681 = ~new_n4679 & ~new_n4680;
  assign new_n4682 = n1916 & n11665;
  assign new_n4683 = n5671 & n11429;
  assign new_n4684 = n4114 & n7374;
  assign new_n4685 = ~new_n4683 & ~new_n4684;
  assign new_n4686 = new_n4683 & new_n4684;
  assign new_n4687 = ~new_n4685 & ~new_n4686;
  assign new_n4688 = new_n4682 & ~new_n4687;
  assign new_n4689 = ~new_n4682 & new_n4687;
  assign new_n4690 = ~new_n4688 & ~new_n4689;
  assign new_n4691 = ~new_n4616 & new_n4625;
  assign new_n4692 = ~new_n4617 & ~new_n4691;
  assign new_n4693 = new_n4690 & ~new_n4692;
  assign new_n4694 = n2777 & n8860;
  assign new_n4695 = ~new_n4614 & ~new_n4694;
  assign new_n4696 = new_n4614 & new_n4694;
  assign new_n4697 = ~new_n4695 & ~new_n4696;
  assign new_n4698 = n3769 & n12605;
  assign new_n4699 = n937 & n6392;
  assign new_n4700 = n10162 & n10642;
  assign new_n4701 = ~new_n4699 & ~new_n4700;
  assign new_n4702 = new_n4699 & new_n4700;
  assign new_n4703 = ~new_n4701 & ~new_n4702;
  assign new_n4704 = new_n4698 & ~new_n4703;
  assign new_n4705 = ~new_n4698 & new_n4703;
  assign new_n4706 = ~new_n4704 & ~new_n4705;
  assign new_n4707 = new_n4697 & new_n4706;
  assign new_n4708 = ~new_n4697 & ~new_n4706;
  assign new_n4709 = ~new_n4707 & ~new_n4708;
  assign new_n4710 = new_n4693 & new_n4709;
  assign new_n4711 = ~new_n4690 & new_n4692;
  assign new_n4712 = new_n4709 & ~new_n4711;
  assign new_n4713 = ~new_n4693 & ~new_n4712;
  assign new_n4714 = ~new_n4710 & ~new_n4713;
  assign new_n4715 = ~new_n4709 & new_n4711;
  assign new_n4716 = ~new_n4714 & ~new_n4715;
  assign new_n4717 = new_n4681 & ~new_n4716;
  assign new_n4718 = ~new_n4681 & new_n4716;
  assign new_n4719 = ~new_n4717 & ~new_n4718;
  assign new_n4720 = new_n4676 & new_n4719;
  assign new_n4721 = ~new_n4676 & ~new_n4719;
  assign new_n4722 = ~new_n4720 & ~new_n4721;
  assign new_n4723 = n5671 & n7374;
  assign new_n4724 = new_n4650 & new_n4675;
  assign new_n4725 = ~new_n4676 & ~new_n4724;
  assign new_n4726 = new_n4723 & new_n4725;
  assign new_n4727 = n5671 & n6392;
  assign new_n4728 = n3769 & n4114;
  assign new_n4729 = new_n4727 & new_n4728;
  assign new_n4730 = ~new_n4661 & ~new_n4662;
  assign new_n4731 = ~new_n4663 & ~new_n4730;
  assign new_n4732 = new_n4663 & new_n4730;
  assign new_n4733 = ~new_n4731 & ~new_n4732;
  assign new_n4734 = new_n4729 & new_n4733;
  assign new_n4735 = ~new_n4666 & new_n4672;
  assign new_n4736 = ~new_n4666 & ~new_n4667;
  assign new_n4737 = new_n4671 & ~new_n4736;
  assign new_n4738 = ~new_n4735 & ~new_n4737;
  assign new_n4739 = new_n4734 & ~new_n4738;
  assign new_n4740 = ~new_n4656 & ~new_n4657;
  assign new_n4741 = ~new_n4673 & ~new_n4740;
  assign new_n4742 = new_n4673 & new_n4740;
  assign new_n4743_1 = ~new_n4741 & ~new_n4742;
  assign new_n4744 = new_n4739 & new_n4743_1;
  assign new_n4745 = ~new_n4723 & ~new_n4725;
  assign new_n4746 = ~new_n4726 & ~new_n4745;
  assign new_n4747 = new_n4744 & new_n4746;
  assign new_n4748_1 = ~new_n4726 & ~new_n4747;
  assign new_n4749 = new_n4722 & ~new_n4748_1;
  assign new_n4750 = ~new_n4722 & new_n4748_1;
  assign new_n4751 = ~new_n4749 & ~new_n4750;
  assign new_n4752 = ~new_n4604 & ~new_n4751;
  assign new_n4753 = new_n4604 & new_n4751;
  assign new_n4754 = ~new_n4752 & ~new_n4753;
  assign new_n4755 = ~new_n4744 & ~new_n4746;
  assign new_n4756 = ~new_n4747 & ~new_n4755;
  assign new_n4757 = ~new_n4553_1 & ~new_n4555;
  assign new_n4758 = ~new_n4556 & ~new_n4757;
  assign new_n4759 = new_n4756 & new_n4758;
  assign new_n4760 = ~new_n4756 & ~new_n4758;
  assign new_n4761 = ~new_n4548 & ~new_n4552;
  assign new_n4762 = ~new_n4553_1 & ~new_n4761;
  assign new_n4763 = ~new_n4739 & ~new_n4743_1;
  assign new_n4764 = ~new_n4744 & ~new_n4763;
  assign new_n4765 = new_n4762 & new_n4764;
  assign new_n4766 = ~new_n4762 & ~new_n4764;
  assign new_n4767 = ~new_n4543 & new_n4547;
  assign new_n4768 = ~new_n4548 & ~new_n4767;
  assign new_n4769 = ~new_n4734 & new_n4738;
  assign new_n4770 = ~new_n4739 & ~new_n4769;
  assign new_n4771 = new_n4768 & new_n4770;
  assign new_n4772 = ~new_n4768 & ~new_n4770;
  assign new_n4773 = ~new_n4729 & ~new_n4733;
  assign new_n4774 = ~new_n4734 & ~new_n4773;
  assign new_n4775 = n5548 & n13201;
  assign new_n4776 = n3769 & n5671;
  assign new_n4777_1 = new_n4775 & new_n4776;
  assign new_n4778 = ~new_n4536 & ~new_n4537;
  assign new_n4779 = ~new_n4538 & ~new_n4778;
  assign new_n4780 = ~new_n4777_1 & ~new_n4779;
  assign new_n4781 = new_n4777_1 & new_n4779;
  assign new_n4782 = ~new_n4727 & ~new_n4728;
  assign new_n4783 = ~new_n4729 & ~new_n4782;
  assign new_n4784 = ~new_n4781 & ~new_n4783;
  assign new_n4785 = ~new_n4780 & ~new_n4784;
  assign new_n4786 = new_n4774 & new_n4785;
  assign new_n4787 = ~new_n4774 & ~new_n4785;
  assign new_n4788 = ~new_n4538 & ~new_n4542;
  assign new_n4789 = ~new_n4543 & ~new_n4788;
  assign new_n4790 = ~new_n4787 & new_n4789;
  assign new_n4791 = ~new_n4786 & ~new_n4790;
  assign new_n4792 = ~new_n4772 & ~new_n4791;
  assign new_n4793 = ~new_n4771 & ~new_n4792;
  assign new_n4794 = ~new_n4766 & ~new_n4793;
  assign new_n4795 = ~new_n4765 & ~new_n4794;
  assign new_n4796 = ~new_n4760 & ~new_n4795;
  assign new_n4797 = ~new_n4759 & ~new_n4796;
  assign new_n4798 = ~new_n4754 & new_n4797;
  assign new_n4799 = new_n4754 & ~new_n4797;
  assign new_n4800 = ~new_n4798 & ~new_n4799;
  assign new_n4801 = new_n4459 & new_n4800;
  assign new_n4802 = ~new_n4459 & ~new_n4800;
  assign new_n4803 = ~new_n4801 & ~new_n4802;
  assign new_n4804 = ~new_n4407 & ~new_n4409;
  assign new_n4805 = ~new_n4410 & ~new_n4804;
  assign new_n4806 = ~new_n4759 & ~new_n4760;
  assign new_n4807 = new_n4795 & ~new_n4806;
  assign new_n4808 = ~new_n4795 & new_n4806;
  assign new_n4809 = ~new_n4807 & ~new_n4808;
  assign new_n4810 = ~new_n4805 & ~new_n4809;
  assign new_n4811 = new_n4805 & new_n4809;
  assign new_n4812 = ~new_n4402 & ~new_n4406;
  assign new_n4813 = ~new_n4407 & ~new_n4812;
  assign new_n4814 = ~new_n4765 & ~new_n4766;
  assign new_n4815 = new_n4793 & ~new_n4814;
  assign new_n4816 = ~new_n4793 & new_n4814;
  assign new_n4817 = ~new_n4815 & ~new_n4816;
  assign new_n4818 = ~new_n4813 & ~new_n4817;
  assign new_n4819 = new_n4813 & new_n4817;
  assign new_n4820 = ~new_n4397 & new_n4401;
  assign new_n4821 = ~new_n4402 & ~new_n4820;
  assign new_n4822 = ~new_n4771 & ~new_n4772;
  assign new_n4823 = new_n4791 & ~new_n4822;
  assign new_n4824_1 = ~new_n4791 & new_n4822;
  assign new_n4825 = ~new_n4823 & ~new_n4824_1;
  assign new_n4826 = ~new_n4821 & ~new_n4825;
  assign new_n4827 = new_n4821 & new_n4825;
  assign new_n4828 = ~new_n4392 & ~new_n4396;
  assign new_n4829 = ~new_n4397 & ~new_n4828;
  assign new_n4830 = ~new_n4786 & ~new_n4787;
  assign new_n4831 = ~new_n4789 & new_n4830;
  assign new_n4832 = new_n4789 & ~new_n4830;
  assign new_n4833 = ~new_n4831 & ~new_n4832;
  assign new_n4834 = ~new_n4829 & new_n4833;
  assign new_n4835 = new_n4829 & ~new_n4833;
  assign new_n4836 = ~new_n4390 & ~new_n4391;
  assign new_n4837 = ~new_n4392 & ~new_n4836;
  assign new_n4838 = ~new_n4780 & ~new_n4781;
  assign new_n4839 = new_n4783 & ~new_n4838;
  assign new_n4840 = ~new_n4783 & new_n4838;
  assign new_n4841 = ~new_n4839 & ~new_n4840;
  assign new_n4842 = ~new_n4837 & new_n4841;
  assign new_n4843 = new_n4837 & ~new_n4841;
  assign new_n4844 = n5801 & n13058;
  assign new_n4845 = ~new_n4775 & ~new_n4776;
  assign new_n4846 = ~new_n4777_1 & ~new_n4845;
  assign new_n4847 = new_n4844 & new_n4846;
  assign new_n4848 = ~new_n4843 & ~new_n4847;
  assign new_n4849 = ~new_n4842 & ~new_n4848;
  assign new_n4850 = ~new_n4835 & ~new_n4849;
  assign new_n4851 = ~new_n4834 & ~new_n4850;
  assign new_n4852 = ~new_n4827 & ~new_n4851;
  assign new_n4853 = ~new_n4826 & ~new_n4852;
  assign new_n4854 = ~new_n4819 & ~new_n4853;
  assign new_n4855 = ~new_n4818 & ~new_n4854;
  assign new_n4856 = ~new_n4811 & ~new_n4855;
  assign new_n4857 = ~new_n4810 & ~new_n4856;
  assign new_n4858 = ~new_n4803 & ~new_n4857;
  assign new_n4859 = new_n4803 & new_n4857;
  assign new_n4860 = ~new_n4858 & ~new_n4859;
  assign new_n4861 = new_n4313 & new_n4860;
  assign new_n4862_1 = ~new_n4313 & ~new_n4860;
  assign new_n4863 = ~new_n4306 & ~new_n4308;
  assign new_n4864_1 = ~new_n4309 & ~new_n4863;
  assign new_n4865 = ~new_n4301 & ~new_n4305;
  assign new_n4866 = ~new_n4306 & ~new_n4865;
  assign new_n4867 = ~new_n4818 & ~new_n4819;
  assign new_n4868 = new_n4853 & ~new_n4867;
  assign new_n4869 = ~new_n4853 & new_n4867;
  assign new_n4870 = ~new_n4868 & ~new_n4869;
  assign new_n4871 = new_n4866 & ~new_n4870;
  assign new_n4872 = ~new_n4866 & new_n4870;
  assign new_n4873 = ~new_n4296 & ~new_n4300;
  assign new_n4874 = ~new_n4301 & ~new_n4873;
  assign new_n4875 = ~new_n4826 & ~new_n4827;
  assign new_n4876 = ~new_n4851 & new_n4875;
  assign new_n4877 = new_n4851 & ~new_n4875;
  assign new_n4878 = ~new_n4876 & ~new_n4877;
  assign new_n4879 = new_n4874 & ~new_n4878;
  assign new_n4880 = ~new_n4874 & new_n4878;
  assign new_n4881 = ~new_n4291 & ~new_n4295;
  assign new_n4882 = ~new_n4296 & ~new_n4881;
  assign new_n4883 = ~new_n4834 & ~new_n4835;
  assign new_n4884 = new_n4849 & ~new_n4883;
  assign new_n4885 = ~new_n4849 & new_n4883;
  assign new_n4886 = ~new_n4884 & ~new_n4885;
  assign new_n4887 = new_n4882 & ~new_n4886;
  assign new_n4888 = ~new_n4882 & new_n4886;
  assign new_n4889 = n3006 & n5729;
  assign new_n4890 = ~new_n4844 & ~new_n4846;
  assign new_n4891 = ~new_n4847 & ~new_n4890;
  assign new_n4892 = new_n4889 & new_n4891;
  assign new_n4893 = ~new_n4289 & ~new_n4290;
  assign new_n4894 = ~new_n4291 & ~new_n4893;
  assign new_n4895 = new_n4892 & new_n4894;
  assign new_n4896 = ~new_n4892 & ~new_n4894;
  assign new_n4897 = ~new_n4842 & ~new_n4843;
  assign new_n4898 = ~new_n4847 & new_n4897;
  assign new_n4899 = new_n4847 & ~new_n4897;
  assign new_n4900 = ~new_n4898 & ~new_n4899;
  assign new_n4901 = ~new_n4896 & ~new_n4900;
  assign new_n4902 = ~new_n4895 & ~new_n4901;
  assign new_n4903 = ~new_n4888 & ~new_n4902;
  assign new_n4904 = ~new_n4887 & ~new_n4903;
  assign new_n4905 = ~new_n4880 & ~new_n4904;
  assign new_n4906 = ~new_n4879 & ~new_n4905;
  assign new_n4907 = ~new_n4872 & ~new_n4906;
  assign new_n4908 = ~new_n4871 & ~new_n4907;
  assign new_n4909 = new_n4864_1 & ~new_n4908;
  assign new_n4910 = ~new_n4864_1 & new_n4908;
  assign new_n4911 = ~new_n4810 & ~new_n4811;
  assign new_n4912 = new_n4855 & ~new_n4911;
  assign new_n4913 = ~new_n4855 & new_n4911;
  assign new_n4914 = ~new_n4912 & ~new_n4913;
  assign new_n4915 = ~new_n4910 & ~new_n4914;
  assign new_n4916 = ~new_n4909 & ~new_n4915;
  assign new_n4917 = ~new_n4862_1 & ~new_n4916;
  assign new_n4918 = ~new_n4861 & ~new_n4917;
  assign new_n4919 = ~new_n4599 & ~new_n4602;
  assign new_n4920 = n10908 & n11835;
  assign new_n4921 = new_n4412 & ~new_n4415;
  assign new_n4922 = ~new_n4416 & ~new_n4921;
  assign new_n4923 = ~new_n4920 & new_n4922;
  assign new_n4924 = new_n4920 & ~new_n4922;
  assign new_n4925 = ~new_n4923 & ~new_n4924;
  assign new_n4926 = ~new_n4420 & ~new_n4422;
  assign new_n4927 = ~new_n4423 & ~new_n4926;
  assign new_n4928 = new_n4925 & new_n4927;
  assign new_n4929 = ~new_n4925 & ~new_n4927;
  assign new_n4930 = ~new_n4928 & ~new_n4929;
  assign new_n4931 = n1636 & n8139;
  assign new_n4932 = n443 & n10560;
  assign new_n4933 = ~new_n4931 & new_n4932;
  assign new_n4934 = new_n4931 & ~new_n4932;
  assign new_n4935 = ~new_n4933 & ~new_n4934;
  assign new_n4936 = n3311 & n4862;
  assign new_n4937 = n5065 & n12003;
  assign new_n4938 = ~new_n4936 & ~new_n4937;
  assign new_n4939 = new_n4936 & new_n4937;
  assign new_n4940 = ~new_n4938 & ~new_n4939;
  assign new_n4941 = ~new_n4935 & new_n4940;
  assign new_n4942 = new_n4935 & ~new_n4940;
  assign new_n4943 = ~new_n4941 & ~new_n4942;
  assign new_n4944 = new_n4930 & new_n4943;
  assign new_n4945 = ~new_n4930 & ~new_n4943;
  assign new_n4946 = ~new_n4944 & ~new_n4945;
  assign new_n4947 = n5356 & n5801;
  assign new_n4948 = ~new_n4445 & ~new_n4449;
  assign new_n4949 = ~new_n4447 & ~new_n4948;
  assign new_n4950 = ~new_n4947 & new_n4949;
  assign new_n4951 = new_n4947 & ~new_n4949;
  assign new_n4952 = ~new_n4950 & ~new_n4951;
  assign new_n4953 = ~new_n4946 & new_n4952;
  assign new_n4954 = new_n4946 & ~new_n4952;
  assign new_n4955 = ~new_n4953 & ~new_n4954;
  assign new_n4956 = ~new_n4440 & ~new_n4443;
  assign new_n4957 = ~new_n4560 & new_n4595;
  assign new_n4958 = ~new_n4561 & ~new_n4957;
  assign new_n4959 = new_n4430 & ~new_n4433;
  assign new_n4960 = ~new_n4434 & ~new_n4959;
  assign new_n4961 = n5548 & n6409;
  assign new_n4962 = n1709 & n13201;
  assign new_n4963 = ~new_n4961 & ~new_n4962;
  assign new_n4964_1 = new_n4961 & new_n4962;
  assign new_n4965 = ~new_n4963 & ~new_n4964_1;
  assign new_n4966 = n817 & n3669;
  assign new_n4967 = n3815 & n5470;
  assign new_n4968 = new_n4966 & ~new_n4967;
  assign new_n4969 = ~new_n4966 & new_n4967;
  assign new_n4970 = ~new_n4968 & ~new_n4969;
  assign new_n4971 = ~new_n4965 & ~new_n4970;
  assign new_n4972 = new_n4965 & new_n4970;
  assign new_n4973 = ~new_n4971 & ~new_n4972;
  assign new_n4974 = ~new_n4960 & new_n4973;
  assign new_n4975 = new_n4960 & ~new_n4973;
  assign new_n4976 = ~new_n4974 & ~new_n4975;
  assign new_n4977 = new_n4958 & ~new_n4976;
  assign new_n4978 = ~new_n4958 & new_n4976;
  assign new_n4979 = ~new_n4977 & ~new_n4978;
  assign new_n4980 = new_n4956 & new_n4979;
  assign new_n4981 = ~new_n4956 & ~new_n4979;
  assign new_n4982 = ~new_n4980 & ~new_n4981;
  assign new_n4983 = new_n4955 & new_n4982;
  assign new_n4984 = ~new_n4955 & ~new_n4982;
  assign new_n4985 = ~new_n4983 & ~new_n4984;
  assign new_n4986 = ~new_n4919 & new_n4985;
  assign new_n4987 = new_n4919 & ~new_n4985;
  assign new_n4988 = ~new_n4986 & ~new_n4987;
  assign new_n4989 = ~new_n4802 & new_n4857;
  assign new_n4990 = ~new_n4801 & ~new_n4989;
  assign new_n4991 = new_n4988 & new_n4990;
  assign new_n4992 = ~new_n4988 & ~new_n4990;
  assign new_n4993 = ~new_n4991 & ~new_n4992;
  assign new_n4994 = ~new_n4282 & ~new_n4311;
  assign new_n4995 = ~new_n4243 & new_n4278;
  assign new_n4996 = ~new_n4244 & ~new_n4995;
  assign new_n4997 = n5729 & n7061;
  assign new_n4998_1 = n3006 & n10122;
  assign new_n4999 = ~new_n4997 & new_n4998_1;
  assign new_n5000 = new_n4997 & ~new_n4998_1;
  assign new_n5001 = ~new_n4999 & ~new_n5000;
  assign new_n5002 = new_n4996 & ~new_n5001;
  assign new_n5003_1 = ~new_n4996 & new_n5001;
  assign new_n5004 = ~new_n5002 & ~new_n5003_1;
  assign new_n5005 = ~new_n4994 & new_n5004;
  assign new_n5006 = new_n4994 & ~new_n5004;
  assign new_n5007 = ~new_n5005 & ~new_n5006;
  assign new_n5008 = n2057 & n7974;
  assign new_n5009 = n5586 & n8163;
  assign new_n5010 = new_n5008 & ~new_n5009;
  assign new_n5011 = ~new_n5008 & new_n5009;
  assign new_n5012 = ~new_n5010 & ~new_n5011;
  assign new_n5013 = n1364 & n11634;
  assign new_n5014 = n3076 & n4141;
  assign new_n5015 = ~new_n5013 & ~new_n5014;
  assign new_n5016 = new_n5013 & new_n5014;
  assign new_n5017 = ~new_n5015 & ~new_n5016;
  assign new_n5018 = n3769 & n5167;
  assign new_n5019 = n4075 & n5671;
  assign new_n5020 = new_n5018 & new_n5019;
  assign new_n5021 = ~new_n5018 & ~new_n5019;
  assign new_n5022 = ~new_n5020 & ~new_n5021;
  assign new_n5023 = new_n5017 & ~new_n5022;
  assign new_n5024 = ~new_n5017 & new_n5022;
  assign new_n5025 = ~new_n5023 & ~new_n5024;
  assign new_n5026 = ~new_n5012 & new_n5025;
  assign new_n5027 = new_n5012 & ~new_n5025;
  assign new_n5028 = ~new_n5026 & ~new_n5027;
  assign new_n5029 = ~new_n4579 & new_n4589;
  assign new_n5030 = ~new_n4578 & ~new_n5029;
  assign new_n5031_1 = new_n4581 & ~new_n4584;
  assign new_n5032 = ~new_n4585 & ~new_n5031_1;
  assign new_n5033 = new_n4563 & ~new_n4566;
  assign new_n5034 = ~new_n4567 & ~new_n5033;
  assign new_n5035 = ~new_n5032 & new_n5034;
  assign new_n5036 = new_n5032 & ~new_n5034;
  assign new_n5037 = ~new_n5035 & ~new_n5036;
  assign new_n5038 = new_n5030 & new_n5037;
  assign new_n5039 = ~new_n5030 & ~new_n5037;
  assign new_n5040 = ~new_n5038 & ~new_n5039;
  assign new_n5041 = new_n5028 & new_n5040;
  assign new_n5042 = ~new_n5028 & ~new_n5040;
  assign new_n5043 = ~new_n5041 & ~new_n5042;
  assign new_n5044 = n937 & n10162;
  assign new_n5045 = n6392 & n12605;
  assign new_n5046 = ~new_n5044 & ~new_n5045;
  assign new_n5047 = new_n5044 & new_n5045;
  assign new_n5048 = ~new_n5046 & ~new_n5047;
  assign new_n5049 = n8860 & n10642;
  assign new_n5050 = n1916 & n2777;
  assign new_n5051 = new_n5049 & ~new_n5050;
  assign new_n5052 = ~new_n5049 & new_n5050;
  assign new_n5053 = ~new_n5051 & ~new_n5052;
  assign new_n5054 = ~new_n5048 & ~new_n5053;
  assign new_n5055 = new_n5048 & new_n5053;
  assign new_n5056 = ~new_n5054 & ~new_n5055;
  assign new_n5057 = ~new_n5043 & new_n5056;
  assign new_n5058 = new_n5043 & ~new_n5056;
  assign new_n5059 = ~new_n5057 & ~new_n5058;
  assign new_n5060_1 = new_n4682 & ~new_n4685;
  assign new_n5061 = ~new_n4686 & ~new_n5060_1;
  assign new_n5062 = ~new_n4696 & new_n4706;
  assign new_n5063 = ~new_n4695 & ~new_n5062;
  assign new_n5064 = ~new_n5061 & ~new_n5063;
  assign new_n5065_1 = new_n5061 & new_n5063;
  assign new_n5066 = ~new_n5064 & ~new_n5065_1;
  assign new_n5067 = ~new_n4713 & new_n5066;
  assign new_n5068 = new_n4713 & ~new_n5066;
  assign new_n5069 = ~new_n5067 & ~new_n5068;
  assign new_n5070 = ~new_n5059 & new_n5069;
  assign new_n5071 = new_n5059 & ~new_n5069;
  assign new_n5072 = ~new_n5070 & ~new_n5071;
  assign new_n5073 = ~new_n4679 & ~new_n4716;
  assign new_n5074 = ~new_n4680 & ~new_n5073;
  assign new_n5075 = ~new_n4698 & ~new_n4702;
  assign new_n5076 = ~new_n4701 & ~new_n5075;
  assign new_n5077 = n4114 & n11429;
  assign new_n5078 = n7374 & n11665;
  assign new_n5079 = ~new_n5077 & new_n5078;
  assign new_n5080 = new_n5077 & ~new_n5078;
  assign new_n5081 = ~new_n5079 & ~new_n5080;
  assign new_n5082 = new_n5076 & ~new_n5081;
  assign new_n5083 = ~new_n5076 & new_n5081;
  assign new_n5084 = ~new_n5082 & ~new_n5083;
  assign new_n5085 = new_n5074 & new_n5084;
  assign new_n5086 = ~new_n5074 & ~new_n5084;
  assign new_n5087 = ~new_n5085 & ~new_n5086;
  assign new_n5088 = new_n5072 & new_n5087;
  assign new_n5089 = ~new_n5072 & ~new_n5087;
  assign new_n5090 = ~new_n5088 & ~new_n5089;
  assign new_n5091 = ~new_n4720 & ~new_n4749;
  assign new_n5092 = ~new_n4574 & new_n4592;
  assign new_n5093 = ~new_n4575 & ~new_n5092;
  assign new_n5094 = ~new_n5091 & ~new_n5093;
  assign new_n5095 = new_n5091 & new_n5093;
  assign new_n5096 = ~new_n5094 & ~new_n5095;
  assign new_n5097 = ~new_n5090 & new_n5096;
  assign new_n5098 = new_n5090 & ~new_n5096;
  assign new_n5099 = ~new_n5097 & ~new_n5098;
  assign new_n5100 = ~new_n5007 & ~new_n5099;
  assign new_n5101 = new_n5007 & new_n5099;
  assign new_n5102 = ~new_n5100 & ~new_n5101;
  assign new_n5103 = ~new_n4454 & ~new_n4457;
  assign new_n5104 = n6168 & n7659;
  assign new_n5105 = n11411 & n12289;
  assign new_n5106 = ~new_n5104 & ~new_n5105;
  assign new_n5107 = new_n5104 & new_n5105;
  assign new_n5108 = ~new_n5106 & ~new_n5107;
  assign new_n5109 = n2771 & n4330;
  assign new_n5110 = n2252 & n5214;
  assign new_n5111 = new_n5109 & ~new_n5110;
  assign new_n5112 = ~new_n5109 & new_n5110;
  assign new_n5113 = ~new_n5111 & ~new_n5112;
  assign new_n5114 = ~new_n5108 & ~new_n5113;
  assign new_n5115 = new_n5108 & new_n5113;
  assign new_n5116 = ~new_n5114 & ~new_n5115;
  assign new_n5117 = new_n4264 & ~new_n4267;
  assign new_n5118 = ~new_n4268 & ~new_n5117;
  assign new_n5119 = n5568 & n5884;
  assign new_n5120 = n8308 & n9747;
  assign new_n5121 = ~new_n5119 & new_n5120;
  assign new_n5122 = new_n5119 & ~new_n5120;
  assign new_n5123 = ~new_n5121 & ~new_n5122;
  assign new_n5124 = new_n5118 & ~new_n5123;
  assign new_n5125 = ~new_n5118 & new_n5123;
  assign new_n5126 = ~new_n5124 & ~new_n5125;
  assign new_n5127 = new_n5116 & new_n5126;
  assign new_n5128 = ~new_n5116 & ~new_n5126;
  assign new_n5129 = ~new_n5127 & ~new_n5128;
  assign new_n5130 = new_n4248 & ~new_n4251;
  assign new_n5131 = ~new_n4252 & ~new_n5130;
  assign new_n5132 = ~new_n4261 & new_n4272;
  assign new_n5133 = ~new_n4262 & ~new_n5132;
  assign new_n5134 = ~new_n5131 & new_n5133;
  assign new_n5135 = new_n5131 & ~new_n5133;
  assign new_n5136 = ~new_n5134 & ~new_n5135;
  assign new_n5137 = new_n5129 & new_n5136;
  assign new_n5138 = ~new_n5129 & ~new_n5136;
  assign new_n5139 = ~new_n5137 & ~new_n5138;
  assign new_n5140 = ~new_n4258 & ~new_n4275;
  assign new_n5141 = ~new_n4257 & ~new_n5140;
  assign new_n5142 = new_n5139 & ~new_n5141;
  assign new_n5143 = ~new_n5139 & new_n5141;
  assign new_n5144 = ~new_n5142 & ~new_n5143;
  assign new_n5145 = n5920 & ~n10866;
  assign new_n5146 = n9041 & n13058;
  assign new_n5147 = ~new_n5145 & new_n5146;
  assign new_n5148 = new_n5145 & ~new_n5146;
  assign new_n5149 = ~new_n5147 & ~new_n5148;
  assign new_n5150 = ~new_n5144 & new_n5149;
  assign new_n5151 = new_n5144 & ~new_n5149;
  assign new_n5152 = ~new_n5150 & ~new_n5151;
  assign new_n5153 = new_n5103 & new_n5152;
  assign new_n5154 = ~new_n5103 & ~new_n5152;
  assign new_n5155 = ~new_n5153 & ~new_n5154;
  assign new_n5156 = ~new_n4752 & ~new_n4797;
  assign new_n5157 = ~new_n4753 & ~new_n5156;
  assign new_n5158 = new_n5155 & new_n5157;
  assign new_n5159 = ~new_n5155 & ~new_n5157;
  assign new_n5160 = ~new_n5158 & ~new_n5159;
  assign new_n5161 = new_n5102 & new_n5160;
  assign new_n5162 = ~new_n5102 & ~new_n5160;
  assign new_n5163 = ~new_n5161 & ~new_n5162;
  assign new_n5164 = new_n4993 & ~new_n5163;
  assign new_n5165 = ~new_n4993 & new_n5163;
  assign new_n5166 = ~new_n5164 & ~new_n5165;
  assign new_n5167_1 = ~new_n4918 & ~new_n5166;
  assign new_n5168 = new_n4918 & new_n5166;
  assign n831 = new_n5167_1 | new_n5168;
  assign new_n5170 = n8506 & n8940;
  assign new_n5171 = n3085 & n9353;
  assign new_n5172 = new_n5170 & new_n5171;
  assign new_n5173 = ~new_n5170 & ~new_n5171;
  assign new_n5174 = ~new_n5172 & ~new_n5173;
  assign new_n5175 = n411 & n8228;
  assign new_n5176 = new_n5174 & new_n5175;
  assign new_n5177 = ~new_n5174 & ~new_n5175;
  assign new_n5178 = ~new_n5176 & ~new_n5177;
  assign new_n5179 = n2482 & new_n5178;
  assign new_n5180 = ~n2482 & ~new_n5178;
  assign n846 = ~new_n5179 & ~new_n5180;
  assign new_n5182 = n3006 & n9093;
  assign new_n5183 = n5568 & n10451;
  assign new_n5184 = new_n5182 & new_n5183;
  assign new_n5185 = n8308 & n10451;
  assign new_n5186 = n5568 & n9093;
  assign new_n5187 = n3006 & n10594;
  assign new_n5188 = ~new_n5186 & ~new_n5187;
  assign new_n5189_1 = new_n5186 & new_n5187;
  assign new_n5190 = ~new_n5188 & ~new_n5189_1;
  assign new_n5191 = new_n5185 & ~new_n5190;
  assign new_n5192 = ~new_n5185 & new_n5190;
  assign new_n5193 = ~new_n5191 & ~new_n5192;
  assign new_n5194 = new_n5184 & ~new_n5193;
  assign new_n5195 = ~new_n5184 & new_n5193;
  assign new_n5196 = ~new_n5194 & ~new_n5195;
  assign new_n5197 = n5671 & n7720;
  assign new_n5198 = n287 & n4114;
  assign new_n5199 = new_n5197 & new_n5198;
  assign new_n5200 = n287 & n11665;
  assign new_n5201 = n4114 & n7720;
  assign new_n5202 = n5671 & n12482;
  assign new_n5203 = ~new_n5201 & ~new_n5202;
  assign new_n5204 = new_n5201 & new_n5202;
  assign new_n5205 = ~new_n5203 & ~new_n5204;
  assign new_n5206 = new_n5200 & ~new_n5205;
  assign new_n5207 = ~new_n5200 & new_n5205;
  assign new_n5208 = ~new_n5206 & ~new_n5207;
  assign new_n5209 = new_n5199 & ~new_n5208;
  assign new_n5210 = ~new_n5199 & new_n5208;
  assign new_n5211 = ~new_n5209 & ~new_n5210;
  assign new_n5212 = n1007 & n13201;
  assign new_n5213 = n2057 & n11058;
  assign new_n5214_1 = new_n5212 & new_n5213;
  assign new_n5215 = n5586 & n11058;
  assign new_n5216 = n1007 & n2057;
  assign new_n5217 = n5969 & n13201;
  assign new_n5218 = ~new_n5216 & ~new_n5217;
  assign new_n5219 = new_n5216 & new_n5217;
  assign new_n5220 = ~new_n5218 & ~new_n5219;
  assign new_n5221 = new_n5215 & ~new_n5220;
  assign new_n5222 = ~new_n5215 & new_n5220;
  assign new_n5223 = ~new_n5221 & ~new_n5222;
  assign new_n5224 = new_n5214_1 & ~new_n5223;
  assign new_n5225 = ~new_n5214_1 & new_n5223;
  assign new_n5226 = ~new_n5224 & ~new_n5225;
  assign new_n5227 = ~new_n5211 & ~new_n5226;
  assign new_n5228 = new_n5211 & new_n5226;
  assign new_n5229 = ~new_n5227 & ~new_n5228;
  assign new_n5230 = n287 & n5671;
  assign new_n5231 = n11058 & n13201;
  assign new_n5232 = new_n5230 & new_n5231;
  assign new_n5233 = ~new_n5197 & ~new_n5198;
  assign new_n5234 = ~new_n5199 & ~new_n5233;
  assign new_n5235 = new_n5232 & new_n5234;
  assign new_n5236 = ~new_n5232 & ~new_n5234;
  assign new_n5237 = ~new_n5212 & ~new_n5213;
  assign new_n5238 = ~new_n5214_1 & ~new_n5237;
  assign new_n5239 = ~new_n5236 & new_n5238;
  assign new_n5240 = ~new_n5235 & ~new_n5239;
  assign new_n5241 = ~new_n5229 & ~new_n5240;
  assign new_n5242 = new_n5229 & new_n5240;
  assign new_n5243 = ~new_n5241 & ~new_n5242;
  assign new_n5244 = n5801 & n6085;
  assign new_n5245 = n5962 & n10908;
  assign new_n5246 = new_n5244 & new_n5245;
  assign new_n5247 = n5962 & n10560;
  assign new_n5248 = n6085 & n10908;
  assign new_n5249 = n5801 & n9906;
  assign new_n5250 = ~new_n5248 & ~new_n5249;
  assign new_n5251 = new_n5248 & new_n5249;
  assign new_n5252 = ~new_n5250 & ~new_n5251;
  assign new_n5253 = new_n5247 & ~new_n5252;
  assign new_n5254 = ~new_n5247 & new_n5252;
  assign new_n5255 = ~new_n5253 & ~new_n5254;
  assign new_n5256 = new_n5246 & ~new_n5255;
  assign new_n5257 = ~new_n5246 & new_n5255;
  assign new_n5258 = ~new_n5256 & ~new_n5257;
  assign new_n5259 = ~new_n5244 & ~new_n5245;
  assign new_n5260 = ~new_n5246 & ~new_n5259;
  assign new_n5261 = ~new_n5235 & ~new_n5236;
  assign new_n5262 = new_n5238 & ~new_n5261;
  assign new_n5263 = ~new_n5238 & new_n5261;
  assign new_n5264 = ~new_n5262 & ~new_n5263;
  assign new_n5265 = new_n5260 & ~new_n5264;
  assign new_n5266 = ~new_n5260 & new_n5264;
  assign new_n5267 = n5801 & n5962;
  assign new_n5268 = ~new_n5230 & ~new_n5231;
  assign new_n5269 = ~new_n5232 & ~new_n5268;
  assign new_n5270 = new_n5267 & new_n5269;
  assign new_n5271 = ~new_n5266 & new_n5270;
  assign new_n5272 = ~new_n5265 & ~new_n5271;
  assign new_n5273 = ~new_n5258 & new_n5272;
  assign new_n5274 = new_n5258 & ~new_n5272;
  assign new_n5275 = ~new_n5273 & ~new_n5274;
  assign new_n5276 = ~new_n5243 & new_n5275;
  assign new_n5277 = new_n5243 & ~new_n5275;
  assign new_n5278 = ~new_n5276 & ~new_n5277;
  assign new_n5279 = ~new_n5196 & ~new_n5278;
  assign new_n5280 = new_n5196 & new_n5278;
  assign new_n5281 = ~new_n5182 & ~new_n5183;
  assign new_n5282 = ~new_n5184 & ~new_n5281;
  assign new_n5283 = n3006 & n10451;
  assign new_n5284 = ~new_n5267 & ~new_n5269;
  assign new_n5285 = ~new_n5270 & ~new_n5284;
  assign new_n5286 = new_n5283 & new_n5285;
  assign new_n5287 = ~new_n5282 & ~new_n5286;
  assign new_n5288 = new_n5282 & new_n5286;
  assign new_n5289 = ~new_n5265 & ~new_n5266;
  assign new_n5290 = ~new_n5270 & ~new_n5289;
  assign new_n5291 = new_n5270 & new_n5289;
  assign new_n5292 = ~new_n5290 & ~new_n5291;
  assign new_n5293 = ~new_n5288 & ~new_n5292;
  assign new_n5294 = ~new_n5287 & ~new_n5293;
  assign new_n5295 = ~new_n5280 & ~new_n5294;
  assign new_n5296 = ~new_n5279 & ~new_n5295;
  assign new_n5297 = n3006 & n3409;
  assign new_n5298 = new_n5185 & ~new_n5188;
  assign new_n5299 = ~new_n5189_1 & ~new_n5298;
  assign new_n5300 = ~new_n5297 & new_n5299;
  assign new_n5301 = new_n5297 & ~new_n5299;
  assign new_n5302 = ~new_n5300 & ~new_n5301;
  assign new_n5303 = n5214 & n10451;
  assign new_n5304 = n5568 & n10594;
  assign new_n5305 = n8308 & n9093;
  assign new_n5306 = ~new_n5304 & ~new_n5305;
  assign new_n5307 = new_n5304 & new_n5305;
  assign new_n5308 = ~new_n5306 & ~new_n5307;
  assign new_n5309 = new_n5303 & ~new_n5308;
  assign new_n5310 = ~new_n5303 & new_n5308;
  assign new_n5311 = ~new_n5309 & ~new_n5310;
  assign new_n5312 = ~new_n5302 & new_n5311;
  assign new_n5313 = new_n5302 & ~new_n5311;
  assign new_n5314 = ~new_n5312 & ~new_n5313;
  assign new_n5315 = ~new_n5194 & ~new_n5314;
  assign new_n5316 = new_n5194 & new_n5314;
  assign new_n5317 = ~new_n5315 & ~new_n5316;
  assign new_n5318 = n5801 & n11109;
  assign new_n5319 = new_n5247 & ~new_n5250;
  assign new_n5320_1 = ~new_n5251 & ~new_n5319;
  assign new_n5321 = ~new_n5318 & new_n5320_1;
  assign new_n5322 = new_n5318 & ~new_n5320_1;
  assign new_n5323 = ~new_n5321 & ~new_n5322;
  assign new_n5324 = n5962 & n12003;
  assign new_n5325 = n9906 & n10908;
  assign new_n5326 = n6085 & n10560;
  assign new_n5327 = ~new_n5325 & ~new_n5326;
  assign new_n5328 = new_n5325 & new_n5326;
  assign new_n5329 = ~new_n5327 & ~new_n5328;
  assign new_n5330 = new_n5324 & ~new_n5329;
  assign new_n5331 = ~new_n5324 & new_n5329;
  assign new_n5332 = ~new_n5330 & ~new_n5331;
  assign new_n5333 = ~new_n5323 & new_n5332;
  assign new_n5334 = new_n5323 & ~new_n5332;
  assign new_n5335 = ~new_n5333 & ~new_n5334;
  assign new_n5336 = ~new_n5256 & ~new_n5335;
  assign new_n5337 = new_n5256 & new_n5335;
  assign new_n5338 = ~new_n5336 & ~new_n5337;
  assign new_n5339 = n5671 & n9570;
  assign new_n5340 = new_n5200 & ~new_n5203;
  assign new_n5341 = ~new_n5204 & ~new_n5340;
  assign new_n5342 = ~new_n5339 & new_n5341;
  assign new_n5343 = new_n5339 & ~new_n5341;
  assign new_n5344 = ~new_n5342 & ~new_n5343;
  assign new_n5345 = n287 & n2777;
  assign new_n5346 = n4114 & n12482;
  assign new_n5347 = n7720 & n11665;
  assign new_n5348 = ~new_n5346 & ~new_n5347;
  assign new_n5349 = new_n5346 & new_n5347;
  assign new_n5350 = ~new_n5348 & ~new_n5349;
  assign new_n5351 = new_n5345 & ~new_n5350;
  assign new_n5352 = ~new_n5345 & new_n5350;
  assign new_n5353 = ~new_n5351 & ~new_n5352;
  assign new_n5354 = ~new_n5344 & new_n5353;
  assign new_n5355 = new_n5344 & ~new_n5353;
  assign new_n5356_1 = ~new_n5354 & ~new_n5355;
  assign new_n5357 = ~new_n5209 & ~new_n5356_1;
  assign new_n5358 = new_n5209 & new_n5356_1;
  assign new_n5359 = ~new_n5357 & ~new_n5358;
  assign new_n5360 = n2498 & n13201;
  assign new_n5361 = new_n5215 & ~new_n5218;
  assign new_n5362 = ~new_n5219 & ~new_n5361;
  assign new_n5363 = ~new_n5360 & new_n5362;
  assign new_n5364_1 = new_n5360 & ~new_n5362;
  assign new_n5365 = ~new_n5363 & ~new_n5364_1;
  assign new_n5366 = n4141 & n11058;
  assign new_n5367 = n2057 & n5969;
  assign new_n5368 = n1007 & n5586;
  assign new_n5369 = ~new_n5367 & ~new_n5368;
  assign new_n5370 = new_n5367 & new_n5368;
  assign new_n5371 = ~new_n5369 & ~new_n5370;
  assign new_n5372 = new_n5366 & ~new_n5371;
  assign new_n5373 = ~new_n5366 & new_n5371;
  assign new_n5374 = ~new_n5372 & ~new_n5373;
  assign new_n5375 = ~new_n5365 & new_n5374;
  assign new_n5376 = new_n5365 & ~new_n5374;
  assign new_n5377 = ~new_n5375 & ~new_n5376;
  assign new_n5378 = new_n5224 & new_n5377;
  assign new_n5379 = ~new_n5224 & ~new_n5377;
  assign new_n5380 = ~new_n5378 & ~new_n5379;
  assign new_n5381 = new_n5359 & new_n5380;
  assign new_n5382 = ~new_n5359 & ~new_n5380;
  assign new_n5383 = ~new_n5381 & ~new_n5382;
  assign new_n5384 = ~new_n5227 & ~new_n5240;
  assign new_n5385 = ~new_n5228 & ~new_n5384;
  assign new_n5386 = new_n5383 & new_n5385;
  assign new_n5387 = ~new_n5383 & ~new_n5385;
  assign new_n5388 = ~new_n5386 & ~new_n5387;
  assign new_n5389 = new_n5338 & ~new_n5388;
  assign new_n5390 = ~new_n5338 & new_n5388;
  assign new_n5391 = ~new_n5389 & ~new_n5390;
  assign new_n5392 = ~new_n5243 & ~new_n5273;
  assign new_n5393 = ~new_n5274 & ~new_n5392;
  assign new_n5394 = new_n5391 & new_n5393;
  assign new_n5395 = ~new_n5391 & ~new_n5393;
  assign new_n5396 = ~new_n5394 & ~new_n5395;
  assign new_n5397 = new_n5317 & ~new_n5396;
  assign new_n5398 = ~new_n5317 & new_n5396;
  assign new_n5399 = ~new_n5397 & ~new_n5398;
  assign new_n5400 = new_n5296 & new_n5399;
  assign new_n5401 = ~new_n5296 & ~new_n5399;
  assign n922 = ~new_n5400 & ~new_n5401;
  assign new_n5403 = n2482 & n4330;
  assign new_n5404 = new_n3997 & ~new_n4000;
  assign new_n5405 = ~new_n4001 & ~new_n5404;
  assign new_n5406 = ~new_n5403 & new_n5405;
  assign new_n5407 = new_n5403 & ~new_n5405;
  assign new_n5408 = ~new_n5406 & ~new_n5407;
  assign new_n5409 = n5729 & n10416;
  assign new_n5410 = n7659 & n10113;
  assign new_n5411 = n1757 & n12289;
  assign new_n5412 = ~new_n5410 & ~new_n5411;
  assign new_n5413 = new_n5410 & new_n5411;
  assign new_n5414 = ~new_n5412 & ~new_n5413;
  assign new_n5415 = new_n5409 & ~new_n5414;
  assign new_n5416 = ~new_n5409 & new_n5414;
  assign new_n5417 = ~new_n5415 & ~new_n5416;
  assign new_n5418 = ~new_n5408 & new_n5417;
  assign new_n5419 = new_n5408 & ~new_n5417;
  assign new_n5420 = ~new_n5418 & ~new_n5419;
  assign new_n5421 = new_n4007 & new_n5420;
  assign new_n5422 = n2252 & n2482;
  assign new_n5423 = n4330 & n10113;
  assign new_n5424 = new_n5409 & ~new_n5412;
  assign new_n5425 = ~new_n5413 & ~new_n5424;
  assign new_n5426 = ~new_n5423 & new_n5425;
  assign new_n5427_1 = new_n5423 & ~new_n5425;
  assign new_n5428 = ~new_n5426 & ~new_n5427_1;
  assign new_n5429 = n5729 & n11030;
  assign new_n5430 = n1757 & n7659;
  assign new_n5431 = n10416 & n12289;
  assign new_n5432 = ~new_n5430 & ~new_n5431;
  assign new_n5433 = new_n5430 & new_n5431;
  assign new_n5434 = ~new_n5432 & ~new_n5433;
  assign new_n5435 = new_n5429 & ~new_n5434;
  assign new_n5436 = ~new_n5429 & new_n5434;
  assign new_n5437 = ~new_n5435 & ~new_n5436;
  assign new_n5438 = ~new_n5428 & new_n5437;
  assign new_n5439 = new_n5428 & ~new_n5437;
  assign new_n5440 = ~new_n5438 & ~new_n5439;
  assign new_n5441 = ~new_n5422 & ~new_n5440;
  assign new_n5442 = new_n5422 & new_n5440;
  assign new_n5443 = ~new_n5441 & ~new_n5442;
  assign new_n5444 = ~new_n5407 & new_n5417;
  assign new_n5445 = ~new_n5406 & ~new_n5444;
  assign new_n5446 = ~new_n5443 & ~new_n5445;
  assign new_n5447 = new_n5443 & new_n5445;
  assign new_n5448 = ~new_n5446 & ~new_n5447;
  assign new_n5449 = ~new_n5421 & ~new_n5448;
  assign new_n5450 = new_n5421 & new_n5448;
  assign new_n5451 = ~new_n5449 & ~new_n5450;
  assign new_n5452 = ~new_n4007 & ~new_n5420;
  assign new_n5453 = ~new_n5421 & ~new_n5452;
  assign new_n5454 = ~new_n4098 & new_n4102;
  assign new_n5455 = ~new_n4099 & ~new_n5454;
  assign new_n5456 = n1636 & n8228;
  assign new_n5457 = new_n4054 & ~new_n4057;
  assign new_n5458 = ~new_n4058 & ~new_n5457;
  assign new_n5459 = ~new_n5456 & new_n5458;
  assign new_n5460 = new_n5456 & ~new_n5458;
  assign new_n5461 = ~new_n5459 & ~new_n5460;
  assign new_n5462 = n3130 & n13058;
  assign new_n5463 = n4862 & n11236;
  assign new_n5464 = n4382 & n5920;
  assign new_n5465 = ~new_n5463 & ~new_n5464;
  assign new_n5466 = new_n5463 & new_n5464;
  assign new_n5467 = ~new_n5465 & ~new_n5466;
  assign new_n5468 = new_n5462 & ~new_n5467;
  assign new_n5469 = ~new_n5462 & new_n5467;
  assign new_n5470_1 = ~new_n5468 & ~new_n5469;
  assign new_n5471 = ~new_n5461 & new_n5470_1;
  assign new_n5472 = new_n5461 & ~new_n5470_1;
  assign new_n5473 = ~new_n5471 & ~new_n5472;
  assign new_n5474 = ~new_n4064 & ~new_n5473;
  assign new_n5475 = new_n4064 & new_n5473;
  assign new_n5476 = ~new_n5474 & ~new_n5475;
  assign new_n5477 = ~new_n4090 & ~new_n4094;
  assign new_n5478 = ~new_n4091 & ~new_n5477;
  assign new_n5479 = n8860 & n8940;
  assign new_n5480 = new_n4066 & ~new_n4069;
  assign new_n5481 = ~new_n4070 & ~new_n5480;
  assign new_n5482 = ~new_n5479 & new_n5481;
  assign new_n5483 = new_n5479 & ~new_n5481;
  assign new_n5484 = ~new_n5482 & ~new_n5483;
  assign new_n5485 = n3769 & n10522;
  assign new_n5486 = n4964 & n10162;
  assign new_n5487 = n5684 & n6392;
  assign new_n5488 = ~new_n5486 & ~new_n5487;
  assign new_n5489 = new_n5486 & new_n5487;
  assign new_n5490 = ~new_n5488 & ~new_n5489;
  assign new_n5491 = new_n5485 & ~new_n5490;
  assign new_n5492 = ~new_n5485 & new_n5490;
  assign new_n5493 = ~new_n5491 & ~new_n5492;
  assign new_n5494 = ~new_n5484 & new_n5493;
  assign new_n5495 = new_n5484 & ~new_n5493;
  assign new_n5496 = ~new_n5494 & ~new_n5495;
  assign new_n5497 = ~new_n4076 & ~new_n5496;
  assign new_n5498 = new_n4076 & new_n5496;
  assign new_n5499 = ~new_n5497 & ~new_n5498;
  assign new_n5500 = n9353 & n11634;
  assign new_n5501 = new_n4078 & ~new_n4081;
  assign new_n5502 = ~new_n4082 & ~new_n5501;
  assign new_n5503 = ~new_n5500 & new_n5502;
  assign new_n5504 = new_n5500 & ~new_n5502;
  assign new_n5505 = ~new_n5503 & ~new_n5504;
  assign new_n5506 = n5548 & n12750;
  assign new_n5507 = n817 & n6333;
  assign new_n5508 = n1912 & n3815;
  assign new_n5509 = ~new_n5507 & ~new_n5508;
  assign new_n5510 = new_n5507 & new_n5508;
  assign new_n5511 = ~new_n5509 & ~new_n5510;
  assign new_n5512 = new_n5506 & ~new_n5511;
  assign new_n5513 = ~new_n5506 & new_n5511;
  assign new_n5514 = ~new_n5512 & ~new_n5513;
  assign new_n5515 = ~new_n5505 & new_n5514;
  assign new_n5516 = new_n5505 & ~new_n5514;
  assign new_n5517 = ~new_n5515 & ~new_n5516;
  assign new_n5518 = new_n4088 & new_n5517;
  assign new_n5519 = ~new_n4088 & ~new_n5517;
  assign new_n5520 = ~new_n5518 & ~new_n5519;
  assign new_n5521 = new_n5499 & new_n5520;
  assign new_n5522 = ~new_n5499 & ~new_n5520;
  assign new_n5523 = ~new_n5521 & ~new_n5522;
  assign new_n5524 = new_n5478 & ~new_n5523;
  assign new_n5525 = ~new_n5478 & new_n5523;
  assign new_n5526 = ~new_n5524 & ~new_n5525;
  assign new_n5527 = ~new_n5476 & new_n5526;
  assign new_n5528 = new_n5476 & ~new_n5526;
  assign new_n5529 = ~new_n5527 & ~new_n5528;
  assign new_n5530 = new_n5455 & new_n5529;
  assign new_n5531 = ~new_n5455 & ~new_n5529;
  assign new_n5532 = ~new_n5530 & ~new_n5531;
  assign new_n5533 = new_n5453 & ~new_n5532;
  assign new_n5534 = ~new_n5453 & new_n5532;
  assign new_n5535 = ~new_n4109 & ~new_n5534;
  assign new_n5536_1 = ~new_n5533 & ~new_n5535;
  assign new_n5537 = ~new_n5451 & new_n5536_1;
  assign new_n5538 = new_n5451 & ~new_n5536_1;
  assign new_n5539 = ~new_n5537 & ~new_n5538;
  assign new_n5540 = n5065 & n8228;
  assign new_n5541 = n1636 & n11236;
  assign new_n5542 = new_n5462 & ~new_n5465;
  assign new_n5543 = ~new_n5466 & ~new_n5542;
  assign new_n5544 = ~new_n5541 & new_n5543;
  assign new_n5545 = new_n5541 & ~new_n5543;
  assign new_n5546 = ~new_n5544 & ~new_n5545;
  assign new_n5547 = n9732 & n13058;
  assign new_n5548_1 = n4382 & n4862;
  assign new_n5549_1 = n3130 & n5920;
  assign new_n5550 = ~new_n5548_1 & ~new_n5549_1;
  assign new_n5551 = new_n5548_1 & new_n5549_1;
  assign new_n5552 = ~new_n5550 & ~new_n5551;
  assign new_n5553 = new_n5547 & ~new_n5552;
  assign new_n5554 = ~new_n5547 & new_n5552;
  assign new_n5555 = ~new_n5553 & ~new_n5554;
  assign new_n5556 = ~new_n5546 & new_n5555;
  assign new_n5557_1 = new_n5546 & ~new_n5555;
  assign new_n5558 = ~new_n5556 & ~new_n5557_1;
  assign new_n5559 = ~new_n5540 & ~new_n5558;
  assign new_n5560 = new_n5540 & new_n5558;
  assign new_n5561 = ~new_n5559 & ~new_n5560;
  assign new_n5562 = ~new_n5459 & ~new_n5470_1;
  assign new_n5563 = ~new_n5460 & ~new_n5562;
  assign new_n5564 = ~new_n5561 & new_n5563;
  assign new_n5565 = new_n5561 & ~new_n5563;
  assign new_n5566 = ~new_n5564 & ~new_n5565;
  assign new_n5567 = ~new_n5475 & ~new_n5566;
  assign new_n5568_1 = new_n5475 & new_n5566;
  assign new_n5569 = ~new_n5567 & ~new_n5568_1;
  assign new_n5570 = n1916 & n8940;
  assign new_n5571 = n4964 & n8860;
  assign new_n5572 = new_n5485 & ~new_n5488;
  assign new_n5573 = ~new_n5489 & ~new_n5572;
  assign new_n5574 = ~new_n5571 & new_n5573;
  assign new_n5575 = new_n5571 & ~new_n5573;
  assign new_n5576 = ~new_n5574 & ~new_n5575;
  assign new_n5577 = n3769 & n10770;
  assign new_n5578 = n5684 & n10162;
  assign new_n5579 = n6392 & n10522;
  assign new_n5580 = ~new_n5578 & ~new_n5579;
  assign new_n5581 = new_n5578 & new_n5579;
  assign new_n5582 = ~new_n5580 & ~new_n5581;
  assign new_n5583 = new_n5577 & ~new_n5582;
  assign new_n5584 = ~new_n5577 & new_n5582;
  assign new_n5585 = ~new_n5583 & ~new_n5584;
  assign new_n5586_1 = ~new_n5576 & new_n5585;
  assign new_n5587 = new_n5576 & ~new_n5585;
  assign new_n5588 = ~new_n5586_1 & ~new_n5587;
  assign new_n5589 = ~new_n5570 & ~new_n5588;
  assign new_n5590 = new_n5570 & new_n5588;
  assign new_n5591 = ~new_n5589 & ~new_n5590;
  assign new_n5592 = ~new_n5482 & ~new_n5493;
  assign new_n5593 = ~new_n5483 & ~new_n5592;
  assign new_n5594 = ~new_n5591 & ~new_n5593;
  assign new_n5595 = ~new_n5590 & new_n5593;
  assign new_n5596 = ~new_n5589 & new_n5595;
  assign new_n5597 = ~new_n5594 & ~new_n5596;
  assign new_n5598 = ~new_n5498 & new_n5597;
  assign new_n5599 = new_n5498 & ~new_n5597;
  assign new_n5600 = ~new_n5598 & ~new_n5599;
  assign new_n5601 = n3076 & n9353;
  assign new_n5602 = n6333 & n11634;
  assign new_n5603 = new_n5506 & ~new_n5509;
  assign new_n5604 = ~new_n5510 & ~new_n5603;
  assign new_n5605 = ~new_n5602 & new_n5604;
  assign new_n5606 = new_n5602 & ~new_n5604;
  assign new_n5607 = ~new_n5605 & ~new_n5606;
  assign new_n5608 = n5548 & n9620;
  assign new_n5609_1 = n817 & n1912;
  assign new_n5610 = n3815 & n12750;
  assign new_n5611 = ~new_n5609_1 & ~new_n5610;
  assign new_n5612 = new_n5609_1 & new_n5610;
  assign new_n5613 = ~new_n5611 & ~new_n5612;
  assign new_n5614 = new_n5608 & ~new_n5613;
  assign new_n5615 = ~new_n5608 & new_n5613;
  assign new_n5616 = ~new_n5614 & ~new_n5615;
  assign new_n5617 = ~new_n5607 & new_n5616;
  assign new_n5618 = new_n5607 & ~new_n5616;
  assign new_n5619 = ~new_n5617 & ~new_n5618;
  assign new_n5620 = ~new_n5601 & ~new_n5619;
  assign new_n5621 = new_n5601 & new_n5619;
  assign new_n5622 = ~new_n5620 & ~new_n5621;
  assign new_n5623 = ~new_n5504 & new_n5514;
  assign new_n5624 = ~new_n5503 & ~new_n5623;
  assign new_n5625 = ~new_n5622 & ~new_n5624;
  assign new_n5626 = new_n5622 & new_n5624;
  assign new_n5627 = ~new_n5625 & ~new_n5626;
  assign new_n5628 = ~new_n5518 & ~new_n5627;
  assign new_n5629 = new_n5518 & new_n5627;
  assign new_n5630 = ~new_n5628 & ~new_n5629;
  assign new_n5631 = new_n5600 & new_n5630;
  assign new_n5632 = ~new_n5600 & ~new_n5630;
  assign new_n5633 = ~new_n5631 & ~new_n5632;
  assign new_n5634 = ~new_n5478 & ~new_n5521;
  assign new_n5635 = ~new_n5522 & ~new_n5634;
  assign new_n5636 = new_n5633 & new_n5635;
  assign new_n5637 = ~new_n5633 & ~new_n5635;
  assign new_n5638 = ~new_n5636 & ~new_n5637;
  assign new_n5639 = ~new_n5569 & ~new_n5638;
  assign new_n5640 = new_n5569 & new_n5638;
  assign new_n5641 = ~new_n5639 & ~new_n5640;
  assign new_n5642 = ~new_n5455 & ~new_n5527;
  assign new_n5643 = ~new_n5528 & ~new_n5642;
  assign new_n5644 = new_n5641 & new_n5643;
  assign new_n5645 = ~new_n5641 & ~new_n5643;
  assign new_n5646 = ~new_n5644 & ~new_n5645;
  assign new_n5647 = ~new_n5539 & new_n5646;
  assign new_n5648 = new_n5539 & ~new_n5646;
  assign n927 = ~new_n5647 & ~new_n5648;
  assign new_n5650 = n3085 & n3178;
  assign new_n5651 = n8466 & n8506;
  assign new_n5652 = new_n5650 & new_n5651;
  assign new_n5653 = ~new_n5650 & ~new_n5651;
  assign new_n5654 = ~new_n5652 & ~new_n5653;
  assign new_n5655 = n411 & n9216;
  assign new_n5656 = new_n5654 & new_n5655;
  assign new_n5657 = ~new_n5654 & ~new_n5655;
  assign new_n5658 = ~new_n5656 & ~new_n5657;
  assign new_n5659 = n7772 & new_n5658;
  assign new_n5660 = ~n7772 & ~new_n5658;
  assign n985 = ~new_n5659 & ~new_n5660;
  assign new_n5662 = n2758 & n7772;
  assign new_n5663 = n4470 & n7529;
  assign new_n5664 = new_n5662 & new_n5663;
  assign new_n5665 = n4470 & n7715;
  assign new_n5666 = n2758 & n7529;
  assign new_n5667 = n4006 & n7772;
  assign new_n5668 = ~new_n5666 & ~new_n5667;
  assign new_n5669 = new_n5666 & new_n5667;
  assign new_n5670 = ~new_n5668 & ~new_n5669;
  assign new_n5671_1 = new_n5665 & ~new_n5670;
  assign new_n5672 = ~new_n5665 & new_n5670;
  assign new_n5673 = ~new_n5671_1 & ~new_n5672;
  assign new_n5674 = new_n5664 & ~new_n5673;
  assign new_n5675 = n7772 & n12306;
  assign new_n5676 = new_n5665 & ~new_n5668;
  assign new_n5677 = ~new_n5669 & ~new_n5676;
  assign new_n5678 = ~new_n5675 & new_n5677;
  assign new_n5679 = new_n5675 & ~new_n5677;
  assign new_n5680 = ~new_n5678 & ~new_n5679;
  assign new_n5681 = n4006 & n7529;
  assign new_n5682 = n2458 & n4470;
  assign new_n5683 = n2758 & n7715;
  assign new_n5684_1 = ~new_n5682 & ~new_n5683;
  assign new_n5685 = n2458 & n2758;
  assign new_n5686 = new_n5665 & new_n5685;
  assign new_n5687 = ~new_n5684_1 & ~new_n5686;
  assign new_n5688 = ~new_n5681 & new_n5687;
  assign new_n5689 = new_n5681 & ~new_n5687;
  assign new_n5690 = ~new_n5688 & ~new_n5689;
  assign new_n5691 = new_n5680 & ~new_n5690;
  assign new_n5692 = ~new_n5680 & new_n5690;
  assign new_n5693 = ~new_n5691 & ~new_n5692;
  assign new_n5694 = new_n5674 & new_n5693;
  assign new_n5695 = n4748 & n7772;
  assign new_n5696 = n7529 & n12306;
  assign new_n5697 = ~new_n5681 & ~new_n5686;
  assign new_n5698 = ~new_n5684_1 & ~new_n5697;
  assign new_n5699 = ~new_n5696 & ~new_n5698;
  assign new_n5700 = new_n5696 & new_n5698;
  assign new_n5701 = ~new_n5699 & ~new_n5700;
  assign new_n5702 = n4006 & n7715;
  assign new_n5703 = n4470 & n8230;
  assign new_n5704 = ~new_n5685 & ~new_n5703;
  assign new_n5705 = new_n5685 & new_n5703;
  assign new_n5706 = ~new_n5704 & ~new_n5705;
  assign new_n5707 = new_n5702 & ~new_n5706;
  assign new_n5708 = ~new_n5702 & new_n5706;
  assign new_n5709 = ~new_n5707 & ~new_n5708;
  assign new_n5710 = ~new_n5701 & new_n5709;
  assign new_n5711 = new_n5701 & ~new_n5709;
  assign new_n5712 = ~new_n5710 & ~new_n5711;
  assign new_n5713 = ~new_n5695 & ~new_n5712;
  assign new_n5714 = new_n5695 & new_n5712;
  assign new_n5715_1 = ~new_n5713 & ~new_n5714;
  assign new_n5716 = ~new_n5678 & ~new_n5690;
  assign new_n5717 = ~new_n5679 & ~new_n5716;
  assign new_n5718 = ~new_n5715_1 & new_n5717;
  assign new_n5719 = new_n5715_1 & ~new_n5717;
  assign new_n5720 = ~new_n5718 & ~new_n5719;
  assign new_n5721 = new_n5694 & new_n5720;
  assign new_n5722 = n7772 & n9187;
  assign new_n5723 = n4748 & n7529;
  assign new_n5724 = n7715 & n12306;
  assign new_n5725 = ~new_n5723 & ~new_n5724;
  assign new_n5726 = new_n5723 & new_n5724;
  assign new_n5727 = ~new_n5725 & ~new_n5726;
  assign new_n5728 = n2458 & n4006;
  assign new_n5729_1 = n2758 & n8230;
  assign new_n5730 = n4470 & n6668;
  assign new_n5731 = ~new_n5729_1 & ~new_n5730;
  assign new_n5732 = new_n5729_1 & new_n5730;
  assign new_n5733 = ~new_n5731 & ~new_n5732;
  assign new_n5734 = new_n5728 & new_n5733;
  assign new_n5735 = ~new_n5728 & ~new_n5733;
  assign new_n5736 = ~new_n5734 & ~new_n5735;
  assign new_n5737 = new_n5702 & ~new_n5704;
  assign new_n5738 = ~new_n5705 & ~new_n5737;
  assign new_n5739 = ~new_n5736 & new_n5738;
  assign new_n5740 = new_n5736 & ~new_n5738;
  assign new_n5741 = ~new_n5739 & ~new_n5740;
  assign new_n5742 = ~new_n5727 & ~new_n5741;
  assign new_n5743 = new_n5727 & new_n5741;
  assign new_n5744 = ~new_n5742 & ~new_n5743;
  assign new_n5745 = ~new_n5700 & new_n5709;
  assign new_n5746 = ~new_n5699 & ~new_n5745;
  assign new_n5747 = ~new_n5744 & new_n5746;
  assign new_n5748 = new_n5744 & ~new_n5746;
  assign new_n5749 = ~new_n5747 & ~new_n5748;
  assign new_n5750 = ~new_n5713 & ~new_n5717;
  assign new_n5751 = ~new_n5714 & ~new_n5750;
  assign new_n5752 = ~new_n5749 & ~new_n5751;
  assign new_n5753 = new_n5749 & new_n5751;
  assign new_n5754 = ~new_n5752 & ~new_n5753;
  assign new_n5755 = new_n5722 & new_n5754;
  assign new_n5756 = ~new_n5722 & ~new_n5754;
  assign new_n5757 = ~new_n5755 & ~new_n5756;
  assign new_n5758_1 = ~new_n5721 & ~new_n5757;
  assign new_n5759 = new_n5721 & new_n5757;
  assign new_n5760 = ~new_n5758_1 & ~new_n5759;
  assign new_n5761 = ~new_n5694 & ~new_n5720;
  assign new_n5762 = ~new_n5721 & ~new_n5761;
  assign new_n5763 = n10408 & n12348;
  assign new_n5764 = n9216 & n10606;
  assign new_n5765 = new_n5763 & new_n5764;
  assign new_n5766 = n9216 & n12965;
  assign new_n5767 = n10606 & n12348;
  assign new_n5768 = n2068 & n10408;
  assign new_n5769 = ~new_n5767 & ~new_n5768;
  assign new_n5770 = new_n5767 & new_n5768;
  assign new_n5771 = ~new_n5769 & ~new_n5770;
  assign new_n5772 = new_n5766 & ~new_n5771;
  assign new_n5773 = ~new_n5766 & new_n5771;
  assign new_n5774 = ~new_n5772 & ~new_n5773;
  assign new_n5775 = new_n5765 & ~new_n5774;
  assign new_n5776 = n1724 & n9216;
  assign new_n5777 = new_n5766 & ~new_n5769;
  assign new_n5778 = ~new_n5770 & ~new_n5777;
  assign new_n5779 = ~new_n5776 & new_n5778;
  assign new_n5780 = new_n5776 & ~new_n5778;
  assign new_n5781 = ~new_n5779 & ~new_n5780;
  assign new_n5782 = n12348 & n12965;
  assign new_n5783 = n2068 & n10606;
  assign new_n5784 = n10408 & n11324;
  assign new_n5785 = ~new_n5783 & ~new_n5784;
  assign new_n5786 = new_n5783 & new_n5784;
  assign new_n5787 = ~new_n5785 & ~new_n5786;
  assign new_n5788 = new_n5782 & ~new_n5787;
  assign new_n5789 = ~new_n5782 & new_n5787;
  assign new_n5790 = ~new_n5788 & ~new_n5789;
  assign new_n5791 = ~new_n5781 & new_n5790;
  assign new_n5792 = new_n5781 & ~new_n5790;
  assign new_n5793 = ~new_n5791 & ~new_n5792;
  assign new_n5794 = new_n5775 & new_n5793;
  assign new_n5795 = n6937 & n9216;
  assign new_n5796 = n1724 & n12348;
  assign new_n5797 = new_n5782 & ~new_n5785;
  assign new_n5798 = ~new_n5786 & ~new_n5797;
  assign new_n5799 = ~new_n5796 & new_n5798;
  assign new_n5800 = new_n5796 & ~new_n5798;
  assign new_n5801_1 = ~new_n5799 & ~new_n5800;
  assign new_n5802 = n2068 & n12965;
  assign new_n5803 = n10606 & n11324;
  assign new_n5804 = n8183 & n10408;
  assign new_n5805 = ~new_n5803 & ~new_n5804;
  assign new_n5806 = new_n5803 & new_n5804;
  assign new_n5807 = ~new_n5805 & ~new_n5806;
  assign new_n5808 = new_n5802 & ~new_n5807;
  assign new_n5809 = ~new_n5802 & new_n5807;
  assign new_n5810 = ~new_n5808 & ~new_n5809;
  assign new_n5811 = ~new_n5801_1 & new_n5810;
  assign new_n5812 = new_n5801_1 & ~new_n5810;
  assign new_n5813 = ~new_n5811 & ~new_n5812;
  assign new_n5814 = ~new_n5795 & ~new_n5813;
  assign new_n5815 = new_n5795 & new_n5813;
  assign new_n5816 = ~new_n5814 & ~new_n5815;
  assign new_n5817 = ~new_n5779 & ~new_n5790;
  assign new_n5818 = ~new_n5780 & ~new_n5817;
  assign new_n5819 = ~new_n5816 & new_n5818;
  assign new_n5820 = new_n5816 & ~new_n5818;
  assign new_n5821 = ~new_n5819 & ~new_n5820;
  assign new_n5822 = ~new_n5794 & ~new_n5821;
  assign new_n5823 = new_n5794 & new_n5821;
  assign new_n5824 = ~new_n5822 & ~new_n5823;
  assign new_n5825 = n5031 & n8233;
  assign new_n5826 = n4335 & n8466;
  assign new_n5827 = new_n5825 & new_n5826;
  assign new_n5828 = n8466 & n9887;
  assign new_n5829 = n4335 & n5031;
  assign new_n5830 = n9 & n8233;
  assign new_n5831 = ~new_n5829 & ~new_n5830;
  assign new_n5832 = new_n5829 & new_n5830;
  assign new_n5833 = ~new_n5831 & ~new_n5832;
  assign new_n5834 = new_n5828 & ~new_n5833;
  assign new_n5835 = ~new_n5828 & new_n5833;
  assign new_n5836 = ~new_n5834 & ~new_n5835;
  assign new_n5837 = new_n5827 & ~new_n5836;
  assign new_n5838 = n497 & n8466;
  assign new_n5839 = new_n5828 & ~new_n5831;
  assign new_n5840 = ~new_n5832 & ~new_n5839;
  assign new_n5841 = ~new_n5838 & new_n5840;
  assign new_n5842 = new_n5838 & ~new_n5840;
  assign new_n5843 = ~new_n5841 & ~new_n5842;
  assign new_n5844 = n5031 & n9887;
  assign new_n5845 = n9 & n4335;
  assign new_n5846 = n2592 & n8233;
  assign new_n5847 = ~new_n5845 & ~new_n5846;
  assign new_n5848 = new_n5845 & new_n5846;
  assign new_n5849 = ~new_n5847 & ~new_n5848;
  assign new_n5850 = new_n5844 & ~new_n5849;
  assign new_n5851 = ~new_n5844 & new_n5849;
  assign new_n5852 = ~new_n5850 & ~new_n5851;
  assign new_n5853 = ~new_n5843 & new_n5852;
  assign new_n5854 = new_n5843 & ~new_n5852;
  assign new_n5855 = ~new_n5853 & ~new_n5854;
  assign new_n5856 = new_n5837 & new_n5855;
  assign new_n5857 = n2174 & n8466;
  assign new_n5858 = n497 & n5031;
  assign new_n5859 = new_n5844 & ~new_n5847;
  assign new_n5860 = ~new_n5848 & ~new_n5859;
  assign new_n5861 = ~new_n5858 & new_n5860;
  assign new_n5862 = new_n5858 & ~new_n5860;
  assign new_n5863 = ~new_n5861 & ~new_n5862;
  assign new_n5864 = n9 & n9887;
  assign new_n5865 = n2592 & n4335;
  assign new_n5866 = n2590 & n8233;
  assign new_n5867 = ~new_n5865 & ~new_n5866;
  assign new_n5868 = new_n5865 & new_n5866;
  assign new_n5869 = ~new_n5867 & ~new_n5868;
  assign new_n5870 = new_n5864 & ~new_n5869;
  assign new_n5871 = ~new_n5864 & new_n5869;
  assign new_n5872 = ~new_n5870 & ~new_n5871;
  assign new_n5873 = ~new_n5863 & new_n5872;
  assign new_n5874 = new_n5863 & ~new_n5872;
  assign new_n5875 = ~new_n5873 & ~new_n5874;
  assign new_n5876 = ~new_n5857 & ~new_n5875;
  assign new_n5877 = new_n5857 & new_n5875;
  assign new_n5878 = ~new_n5876 & ~new_n5877;
  assign new_n5879 = ~new_n5841 & ~new_n5852;
  assign new_n5880 = ~new_n5842 & ~new_n5879;
  assign new_n5881 = ~new_n5878 & new_n5880;
  assign new_n5882_1 = new_n5878 & ~new_n5880;
  assign new_n5883 = ~new_n5881 & ~new_n5882_1;
  assign new_n5884_1 = ~new_n5856 & ~new_n5883;
  assign new_n5885 = new_n5856 & new_n5883;
  assign new_n5886 = ~new_n5884_1 & ~new_n5885;
  assign new_n5887 = n10063 & n12592;
  assign new_n5888 = n3178 & n9915;
  assign new_n5889 = new_n5887 & new_n5888;
  assign new_n5890 = n3178 & n8332;
  assign new_n5891 = n9915 & n12592;
  assign new_n5892 = n10063 & n10168;
  assign new_n5893 = ~new_n5891 & ~new_n5892;
  assign new_n5894 = new_n5891 & new_n5892;
  assign new_n5895 = ~new_n5893 & ~new_n5894;
  assign new_n5896 = new_n5890 & ~new_n5895;
  assign new_n5897 = ~new_n5890 & new_n5895;
  assign new_n5898 = ~new_n5896 & ~new_n5897;
  assign new_n5899 = new_n5889 & ~new_n5898;
  assign new_n5900 = n3178 & n3832;
  assign new_n5901 = new_n5890 & ~new_n5893;
  assign new_n5902 = ~new_n5894 & ~new_n5901;
  assign new_n5903 = ~new_n5900 & new_n5902;
  assign new_n5904 = new_n5900 & ~new_n5902;
  assign new_n5905 = ~new_n5903 & ~new_n5904;
  assign new_n5906 = n8332 & n12592;
  assign new_n5907 = n9915 & n10168;
  assign new_n5908 = n767 & n10063;
  assign new_n5909 = ~new_n5907 & ~new_n5908;
  assign new_n5910 = new_n5907 & new_n5908;
  assign new_n5911 = ~new_n5909 & ~new_n5910;
  assign new_n5912 = new_n5906 & ~new_n5911;
  assign new_n5913 = ~new_n5906 & new_n5911;
  assign new_n5914 = ~new_n5912 & ~new_n5913;
  assign new_n5915 = ~new_n5905 & new_n5914;
  assign new_n5916 = new_n5905 & ~new_n5914;
  assign new_n5917 = ~new_n5915 & ~new_n5916;
  assign new_n5918 = new_n5899 & new_n5917;
  assign new_n5919 = n2882 & n3178;
  assign new_n5920_1 = n3832 & n12592;
  assign new_n5921 = new_n5906 & ~new_n5909;
  assign new_n5922 = ~new_n5910 & ~new_n5921;
  assign new_n5923 = ~new_n5920_1 & new_n5922;
  assign new_n5924 = new_n5920_1 & ~new_n5922;
  assign new_n5925 = ~new_n5923 & ~new_n5924;
  assign new_n5926 = n8332 & n10168;
  assign new_n5927 = n767 & n9915;
  assign new_n5928 = n10063 & n11537;
  assign new_n5929 = ~new_n5927 & ~new_n5928;
  assign new_n5930 = new_n5927 & new_n5928;
  assign new_n5931 = ~new_n5929 & ~new_n5930;
  assign new_n5932 = new_n5926 & ~new_n5931;
  assign new_n5933 = ~new_n5926 & new_n5931;
  assign new_n5934 = ~new_n5932 & ~new_n5933;
  assign new_n5935 = ~new_n5925 & new_n5934;
  assign new_n5936 = new_n5925 & ~new_n5934;
  assign new_n5937 = ~new_n5935 & ~new_n5936;
  assign new_n5938 = ~new_n5919 & ~new_n5937;
  assign new_n5939 = new_n5919 & new_n5937;
  assign new_n5940 = ~new_n5938 & ~new_n5939;
  assign new_n5941 = ~new_n5903 & ~new_n5914;
  assign new_n5942 = ~new_n5904 & ~new_n5941;
  assign new_n5943 = ~new_n5940 & new_n5942;
  assign new_n5944 = new_n5940 & ~new_n5942;
  assign new_n5945 = ~new_n5943 & ~new_n5944;
  assign new_n5946 = ~new_n5918 & ~new_n5945;
  assign new_n5947 = new_n5918 & new_n5945;
  assign new_n5948 = ~new_n5946 & ~new_n5947;
  assign new_n5949 = ~new_n5837 & ~new_n5855;
  assign new_n5950 = ~new_n5856 & ~new_n5949;
  assign new_n5951 = ~new_n5899 & ~new_n5917;
  assign new_n5952 = ~new_n5918 & ~new_n5951;
  assign new_n5953 = new_n5950 & new_n5952;
  assign new_n5954 = ~new_n5950 & ~new_n5952;
  assign new_n5955 = ~new_n5889 & new_n5898;
  assign new_n5956 = ~new_n5899 & ~new_n5955;
  assign new_n5957 = n8233 & n8466;
  assign new_n5958 = n3178 & n10063;
  assign new_n5959 = new_n5957 & new_n5958;
  assign new_n5960 = ~new_n5887 & ~new_n5888;
  assign new_n5961 = ~new_n5889 & ~new_n5960;
  assign new_n5962_1 = new_n5959 & new_n5961;
  assign new_n5963 = ~new_n5959 & ~new_n5961;
  assign new_n5964 = ~new_n5825 & ~new_n5826;
  assign new_n5965 = ~new_n5827 & ~new_n5964;
  assign new_n5966 = ~new_n5963 & new_n5965;
  assign new_n5967 = ~new_n5962_1 & ~new_n5966;
  assign new_n5968 = new_n5956 & ~new_n5967;
  assign new_n5969_1 = ~new_n5956 & new_n5967;
  assign new_n5970 = ~new_n5827 & new_n5836;
  assign new_n5971 = ~new_n5837 & ~new_n5970;
  assign new_n5972 = ~new_n5969_1 & new_n5971;
  assign new_n5973 = ~new_n5968 & ~new_n5972;
  assign new_n5974 = ~new_n5954 & ~new_n5973;
  assign new_n5975 = ~new_n5953 & ~new_n5974;
  assign new_n5976 = new_n5948 & ~new_n5975;
  assign new_n5977 = ~new_n5948 & new_n5975;
  assign new_n5978 = ~new_n5976 & ~new_n5977;
  assign new_n5979 = new_n5886 & new_n5978;
  assign new_n5980 = ~new_n5886 & ~new_n5978;
  assign new_n5981 = ~new_n5979 & ~new_n5980;
  assign new_n5982 = ~new_n5824 & ~new_n5981;
  assign new_n5983 = new_n5824 & new_n5981;
  assign new_n5984 = ~new_n5982 & ~new_n5983;
  assign new_n5985 = ~new_n5775 & ~new_n5793;
  assign new_n5986 = ~new_n5794 & ~new_n5985;
  assign new_n5987 = ~new_n5953 & ~new_n5954;
  assign new_n5988 = new_n5973 & ~new_n5987;
  assign new_n5989 = ~new_n5973 & new_n5987;
  assign new_n5990 = ~new_n5988 & ~new_n5989;
  assign new_n5991 = ~new_n5986 & ~new_n5990;
  assign new_n5992 = new_n5986 & new_n5990;
  assign new_n5993 = ~new_n5765 & new_n5774;
  assign new_n5994 = ~new_n5775 & ~new_n5993;
  assign new_n5995 = ~new_n5968 & ~new_n5969_1;
  assign new_n5996 = new_n5971 & new_n5995;
  assign new_n5997 = ~new_n5971 & ~new_n5995;
  assign new_n5998 = ~new_n5996 & ~new_n5997;
  assign new_n5999 = ~new_n5994 & ~new_n5998;
  assign new_n6000 = new_n5994 & new_n5998;
  assign new_n6001 = ~new_n5763 & ~new_n5764;
  assign new_n6002 = ~new_n5765 & ~new_n6001;
  assign new_n6003 = ~new_n5962_1 & ~new_n5963;
  assign new_n6004 = new_n5965 & ~new_n6003;
  assign new_n6005 = ~new_n5965 & new_n6003;
  assign new_n6006 = ~new_n6004 & ~new_n6005;
  assign new_n6007 = ~new_n6002 & new_n6006;
  assign new_n6008 = new_n6002 & ~new_n6006;
  assign new_n6009 = n9216 & n10408;
  assign new_n6010 = ~new_n5957 & ~new_n5958;
  assign new_n6011 = ~new_n5959 & ~new_n6010;
  assign new_n6012 = new_n6009 & new_n6011;
  assign new_n6013 = ~new_n6008 & ~new_n6012;
  assign new_n6014 = ~new_n6007 & ~new_n6013;
  assign new_n6015 = ~new_n6000 & ~new_n6014;
  assign new_n6016 = ~new_n5999 & ~new_n6015;
  assign new_n6017 = ~new_n5992 & ~new_n6016;
  assign new_n6018 = ~new_n5991 & ~new_n6017;
  assign new_n6019_1 = ~new_n5984 & ~new_n6018;
  assign new_n6020 = new_n5984 & new_n6018;
  assign new_n6021 = ~new_n6019_1 & ~new_n6020;
  assign new_n6022 = new_n5762 & new_n6021;
  assign new_n6023_1 = ~new_n5762 & ~new_n6021;
  assign new_n6024 = ~new_n5674 & ~new_n5693;
  assign new_n6025 = ~new_n5694 & ~new_n6024;
  assign new_n6026 = ~new_n5991 & ~new_n5992;
  assign new_n6027 = new_n6016 & ~new_n6026;
  assign new_n6028 = ~new_n6016 & new_n6026;
  assign new_n6029 = ~new_n6027 & ~new_n6028;
  assign new_n6030 = new_n6025 & ~new_n6029;
  assign new_n6031 = ~new_n6025 & new_n6029;
  assign new_n6032 = ~new_n5664 & new_n5673;
  assign new_n6033 = ~new_n5674 & ~new_n6032;
  assign new_n6034 = ~new_n5999 & ~new_n6000;
  assign new_n6035 = new_n6014 & ~new_n6034;
  assign new_n6036 = ~new_n6014 & new_n6034;
  assign new_n6037 = ~new_n6035 & ~new_n6036;
  assign new_n6038 = new_n6033 & ~new_n6037;
  assign new_n6039 = ~new_n6033 & new_n6037;
  assign new_n6040 = n4470 & n7772;
  assign new_n6041 = ~new_n6009 & ~new_n6011;
  assign new_n6042 = ~new_n6012 & ~new_n6041;
  assign new_n6043 = new_n6040 & new_n6042;
  assign new_n6044 = ~new_n5662 & ~new_n5663;
  assign new_n6045 = ~new_n5664 & ~new_n6044;
  assign new_n6046 = new_n6043 & new_n6045;
  assign new_n6047 = ~new_n6043 & ~new_n6045;
  assign new_n6048 = ~new_n6007 & ~new_n6008;
  assign new_n6049 = ~new_n6012 & new_n6048;
  assign new_n6050 = new_n6012 & ~new_n6048;
  assign new_n6051 = ~new_n6049 & ~new_n6050;
  assign new_n6052 = ~new_n6047 & ~new_n6051;
  assign new_n6053 = ~new_n6046 & ~new_n6052;
  assign new_n6054 = ~new_n6039 & ~new_n6053;
  assign new_n6055 = ~new_n6038 & ~new_n6054;
  assign new_n6056 = ~new_n6031 & ~new_n6055;
  assign new_n6057 = ~new_n6030 & ~new_n6056;
  assign new_n6058 = ~new_n6023_1 & ~new_n6057;
  assign new_n6059 = ~new_n6022 & ~new_n6058;
  assign new_n6060 = ~new_n5760 & new_n6059;
  assign new_n6061 = new_n5760 & ~new_n6059;
  assign new_n6062 = ~new_n6060 & ~new_n6061;
  assign new_n6063 = n3677 & n9216;
  assign new_n6064 = n1724 & n2068;
  assign new_n6065 = n6937 & n12348;
  assign new_n6066 = ~new_n6064 & ~new_n6065;
  assign new_n6067 = new_n6064 & new_n6065;
  assign new_n6068 = ~new_n6066 & ~new_n6067;
  assign new_n6069 = n11324 & n12965;
  assign new_n6070 = n8183 & n10606;
  assign new_n6071 = n10142 & n10408;
  assign new_n6072 = ~new_n6070 & ~new_n6071;
  assign new_n6073 = new_n6070 & new_n6071;
  assign new_n6074 = ~new_n6072 & ~new_n6073;
  assign new_n6075 = new_n6069 & new_n6074;
  assign new_n6076 = ~new_n6069 & ~new_n6074;
  assign new_n6077 = ~new_n6075 & ~new_n6076;
  assign new_n6078 = new_n5802 & ~new_n5805;
  assign new_n6079 = ~new_n5806 & ~new_n6078;
  assign new_n6080 = ~new_n6077 & new_n6079;
  assign new_n6081 = new_n6077 & ~new_n6079;
  assign new_n6082 = ~new_n6080 & ~new_n6081;
  assign new_n6083 = new_n6068 & new_n6082;
  assign new_n6084 = ~new_n6068 & ~new_n6082;
  assign new_n6085_1 = ~new_n6083 & ~new_n6084;
  assign new_n6086 = ~new_n5799 & ~new_n5810;
  assign new_n6087 = ~new_n5800 & ~new_n6086;
  assign new_n6088 = new_n6085_1 & new_n6087;
  assign new_n6089 = ~new_n6085_1 & ~new_n6087;
  assign new_n6090 = ~new_n6088 & ~new_n6089;
  assign new_n6091 = ~new_n5814 & ~new_n5818;
  assign new_n6092 = ~new_n5815 & ~new_n6091;
  assign new_n6093 = ~new_n6090 & ~new_n6092;
  assign new_n6094 = new_n6090 & new_n6092;
  assign new_n6095 = ~new_n6093 & ~new_n6094;
  assign new_n6096 = new_n6063 & new_n6095;
  assign new_n6097 = ~new_n6063 & ~new_n6095;
  assign new_n6098 = ~new_n6096 & ~new_n6097;
  assign new_n6099 = ~new_n5823 & ~new_n6098;
  assign new_n6100 = new_n5823 & new_n6098;
  assign new_n6101 = ~new_n6099 & ~new_n6100;
  assign new_n6102 = ~new_n5983 & ~new_n6018;
  assign new_n6103_1 = ~new_n5982 & ~new_n6102;
  assign new_n6104 = ~new_n6101 & ~new_n6103_1;
  assign new_n6105 = n3178 & n4357;
  assign new_n6106 = n2882 & n12592;
  assign new_n6107 = n3832 & n10168;
  assign new_n6108 = ~new_n6106 & ~new_n6107;
  assign new_n6109_1 = new_n6106 & new_n6107;
  assign new_n6110 = ~new_n6108 & ~new_n6109_1;
  assign new_n6111 = n767 & n8332;
  assign new_n6112 = n9915 & n11537;
  assign new_n6113 = n951 & n10063;
  assign new_n6114 = ~new_n6112 & ~new_n6113;
  assign new_n6115 = new_n6112 & new_n6113;
  assign new_n6116 = ~new_n6114 & ~new_n6115;
  assign new_n6117 = ~new_n6111 & ~new_n6116;
  assign new_n6118 = new_n6111 & new_n6116;
  assign new_n6119 = ~new_n6117 & ~new_n6118;
  assign new_n6120 = new_n5926 & ~new_n5929;
  assign new_n6121 = ~new_n5930 & ~new_n6120;
  assign new_n6122 = ~new_n6119 & ~new_n6121;
  assign new_n6123 = new_n6119 & new_n6121;
  assign new_n6124 = ~new_n6122 & ~new_n6123;
  assign new_n6125 = ~new_n6110 & new_n6124;
  assign new_n6126 = new_n6110 & ~new_n6124;
  assign new_n6127 = ~new_n6125 & ~new_n6126;
  assign new_n6128 = ~new_n5923 & ~new_n5934;
  assign new_n6129 = ~new_n5924 & ~new_n6128;
  assign new_n6130 = ~new_n6127 & new_n6129;
  assign new_n6131 = new_n6127 & ~new_n6129;
  assign new_n6132 = ~new_n6130 & ~new_n6131;
  assign new_n6133 = ~new_n5938 & ~new_n5942;
  assign new_n6134 = ~new_n5939 & ~new_n6133;
  assign new_n6135 = new_n6132 & ~new_n6134;
  assign new_n6136 = ~new_n6132 & new_n6134;
  assign new_n6137 = ~new_n6135 & ~new_n6136;
  assign new_n6138 = new_n6105 & new_n6137;
  assign new_n6139 = ~new_n6105 & ~new_n6137;
  assign new_n6140 = ~new_n6138 & ~new_n6139;
  assign new_n6141 = ~new_n5947 & ~new_n6140;
  assign new_n6142 = new_n5947 & new_n6140;
  assign new_n6143 = ~new_n6141 & ~new_n6142;
  assign new_n6144 = n3112 & n8466;
  assign new_n6145 = ~new_n5876 & ~new_n5880;
  assign new_n6146 = ~new_n5877 & ~new_n6145;
  assign new_n6147 = n2174 & n5031;
  assign new_n6148 = n9 & n497;
  assign new_n6149_1 = ~new_n6147 & ~new_n6148;
  assign new_n6150 = new_n6147 & new_n6148;
  assign new_n6151 = ~new_n6149_1 & ~new_n6150;
  assign new_n6152 = n2592 & n9887;
  assign new_n6153 = n2590 & n4335;
  assign new_n6154 = n8233 & n11061;
  assign new_n6155 = ~new_n6153 & ~new_n6154;
  assign new_n6156 = new_n6153 & new_n6154;
  assign new_n6157 = ~new_n6155 & ~new_n6156;
  assign new_n6158 = ~new_n6152 & ~new_n6157;
  assign new_n6159 = new_n6152 & new_n6157;
  assign new_n6160 = ~new_n6158 & ~new_n6159;
  assign new_n6161 = new_n5864 & ~new_n5867;
  assign new_n6162 = ~new_n5868 & ~new_n6161;
  assign new_n6163 = ~new_n6160 & new_n6162;
  assign new_n6164 = new_n6160 & ~new_n6162;
  assign new_n6165 = ~new_n6163 & ~new_n6164;
  assign new_n6166 = ~new_n6151 & ~new_n6165;
  assign new_n6167 = new_n6151 & new_n6165;
  assign new_n6168_1 = ~new_n6166 & ~new_n6167;
  assign new_n6169 = ~new_n5861 & ~new_n5872;
  assign new_n6170 = ~new_n5862 & ~new_n6169;
  assign new_n6171 = ~new_n6168_1 & ~new_n6170;
  assign new_n6172 = new_n6168_1 & new_n6170;
  assign new_n6173 = ~new_n6171 & ~new_n6172;
  assign new_n6174 = ~new_n6146 & ~new_n6173;
  assign new_n6175 = new_n6146 & new_n6173;
  assign new_n6176 = ~new_n6174 & ~new_n6175;
  assign new_n6177 = new_n6144 & new_n6176;
  assign new_n6178 = ~new_n6144 & ~new_n6176;
  assign new_n6179 = ~new_n6177 & ~new_n6178;
  assign new_n6180 = ~new_n5885 & ~new_n6179;
  assign new_n6181 = new_n5885 & new_n6179;
  assign new_n6182 = ~new_n6180 & ~new_n6181;
  assign new_n6183 = new_n6143 & new_n6182;
  assign new_n6184 = ~new_n6143 & ~new_n6182;
  assign new_n6185 = ~new_n6183 & ~new_n6184;
  assign new_n6186 = new_n5886 & ~new_n5977;
  assign new_n6187 = ~new_n5976 & ~new_n6186;
  assign new_n6188 = ~new_n6185 & ~new_n6187;
  assign new_n6189 = new_n6185 & new_n6187;
  assign new_n6190 = ~new_n6188 & ~new_n6189;
  assign new_n6191 = new_n6104 & new_n6190;
  assign new_n6192 = new_n6101 & new_n6103_1;
  assign new_n6193 = ~new_n6190 & new_n6192;
  assign new_n6194 = ~new_n6104 & ~new_n6190;
  assign new_n6195 = ~new_n6192 & ~new_n6194;
  assign new_n6196 = ~new_n6193 & ~new_n6195;
  assign new_n6197 = ~new_n6191 & ~new_n6196;
  assign new_n6198 = ~new_n6062 & ~new_n6197;
  assign new_n6199 = new_n6062 & new_n6197;
  assign n1097 = new_n6198 | new_n6199;
  assign new_n6201 = ~new_n5755 & ~new_n5759;
  assign new_n6202 = ~new_n5742 & new_n5746;
  assign new_n6203 = new_n5726 & new_n6202;
  assign new_n6204 = ~new_n5726 & ~new_n6202;
  assign new_n6205 = ~new_n5743 & new_n6204;
  assign new_n6206 = ~new_n6203 & ~new_n6205;
  assign new_n6207 = n1231 & n7772;
  assign new_n6208 = n4748 & n7715;
  assign new_n6209 = n7529 & n9187;
  assign new_n6210 = ~new_n6208 & ~new_n6209;
  assign new_n6211 = new_n6208 & new_n6209;
  assign new_n6212 = ~new_n6210 & ~new_n6211;
  assign new_n6213 = new_n6207 & ~new_n6212;
  assign new_n6214 = ~new_n6207 & new_n6212;
  assign new_n6215 = ~new_n6213 & ~new_n6214;
  assign new_n6216 = ~new_n5734 & new_n5738;
  assign new_n6217 = ~new_n5735 & ~new_n6216;
  assign new_n6218 = new_n6215 & ~new_n6217;
  assign new_n6219 = ~new_n6215 & new_n6217;
  assign new_n6220 = ~new_n6218 & ~new_n6219;
  assign new_n6221 = n2458 & n12306;
  assign new_n6222 = new_n5732 & new_n6221;
  assign new_n6223 = ~new_n5732 & ~new_n6221;
  assign new_n6224 = ~new_n6222 & ~new_n6223;
  assign new_n6225 = n4006 & n8230;
  assign new_n6226 = n2758 & n6668;
  assign new_n6227 = n4470 & n7812;
  assign new_n6228 = ~new_n6226 & ~new_n6227;
  assign new_n6229 = new_n6226 & new_n6227;
  assign new_n6230 = ~new_n6228 & ~new_n6229;
  assign new_n6231 = new_n6225 & ~new_n6230;
  assign new_n6232 = ~new_n6225 & new_n6230;
  assign new_n6233 = ~new_n6231 & ~new_n6232;
  assign new_n6234 = new_n6224 & new_n6233;
  assign new_n6235 = ~new_n6224 & ~new_n6233;
  assign new_n6236 = ~new_n6234 & ~new_n6235;
  assign new_n6237 = new_n6220 & new_n6236;
  assign new_n6238 = ~new_n6220 & ~new_n6236;
  assign new_n6239 = ~new_n6237 & ~new_n6238;
  assign new_n6240 = ~new_n6206 & new_n6239;
  assign new_n6241 = new_n6206 & ~new_n6239;
  assign new_n6242 = ~new_n6240 & ~new_n6241;
  assign new_n6243 = new_n5752 & new_n6242;
  assign new_n6244 = ~new_n5752 & ~new_n6242;
  assign new_n6245 = ~new_n6243 & ~new_n6244;
  assign new_n6246 = ~new_n6201 & new_n6245;
  assign new_n6247 = new_n6201 & ~new_n6245;
  assign new_n6248 = ~new_n6246 & ~new_n6247;
  assign new_n6249 = ~new_n6096 & ~new_n6100;
  assign new_n6250 = ~new_n6084 & ~new_n6087;
  assign new_n6251 = new_n6067 & new_n6250;
  assign new_n6252 = ~new_n6067 & ~new_n6250;
  assign new_n6253 = ~new_n6083 & new_n6252;
  assign new_n6254 = n7729 & n9216;
  assign new_n6255 = n2068 & n6937;
  assign new_n6256 = n3677 & n12348;
  assign new_n6257 = ~new_n6255 & ~new_n6256;
  assign new_n6258 = new_n6255 & new_n6256;
  assign new_n6259 = ~new_n6257 & ~new_n6258;
  assign new_n6260 = new_n6254 & ~new_n6259;
  assign new_n6261 = ~new_n6254 & new_n6259;
  assign new_n6262 = ~new_n6260 & ~new_n6261;
  assign new_n6263 = ~new_n6075 & new_n6079;
  assign new_n6264 = ~new_n6076 & ~new_n6263;
  assign new_n6265 = ~new_n6262 & new_n6264;
  assign new_n6266 = new_n6262 & ~new_n6264;
  assign new_n6267 = ~new_n6265 & ~new_n6266;
  assign new_n6268 = n1724 & n11324;
  assign new_n6269 = new_n6073 & new_n6268;
  assign new_n6270 = ~new_n6073 & ~new_n6268;
  assign new_n6271 = ~new_n6269 & ~new_n6270;
  assign new_n6272 = n8183 & n12965;
  assign new_n6273 = n10142 & n10606;
  assign new_n6274 = n10408 & n10657;
  assign new_n6275 = ~new_n6273 & ~new_n6274;
  assign new_n6276 = new_n6273 & new_n6274;
  assign new_n6277 = ~new_n6275 & ~new_n6276;
  assign new_n6278 = new_n6272 & ~new_n6277;
  assign new_n6279 = ~new_n6272 & new_n6277;
  assign new_n6280 = ~new_n6278 & ~new_n6279;
  assign new_n6281 = new_n6271 & new_n6280;
  assign new_n6282 = ~new_n6271 & ~new_n6280;
  assign new_n6283 = ~new_n6281 & ~new_n6282;
  assign new_n6284 = ~new_n6267 & ~new_n6283;
  assign new_n6285 = new_n6267 & new_n6283;
  assign new_n6286 = ~new_n6284 & ~new_n6285;
  assign new_n6287 = ~new_n6253 & ~new_n6286;
  assign new_n6288 = ~new_n6251 & ~new_n6287;
  assign new_n6289 = new_n6253 & new_n6286;
  assign new_n6290 = new_n6288 & ~new_n6289;
  assign new_n6291 = new_n6251 & ~new_n6286;
  assign new_n6292 = ~new_n6290 & ~new_n6291;
  assign new_n6293 = new_n6093 & ~new_n6292;
  assign new_n6294 = ~new_n6093 & new_n6292;
  assign new_n6295 = ~new_n6293 & ~new_n6294;
  assign new_n6296 = ~new_n6249 & new_n6295;
  assign new_n6297_1 = new_n6249 & ~new_n6295;
  assign new_n6298 = ~new_n6296 & ~new_n6297_1;
  assign new_n6299 = ~new_n6125 & ~new_n6129;
  assign new_n6300 = ~new_n6109_1 & ~new_n6299;
  assign new_n6301_1 = ~new_n6126 & new_n6300;
  assign new_n6302 = new_n6109_1 & new_n6299;
  assign new_n6303 = ~new_n6301_1 & ~new_n6302;
  assign new_n6304 = n8332 & n11537;
  assign new_n6305 = n951 & n9915;
  assign new_n6306 = n401 & n10063;
  assign new_n6307 = ~new_n6305 & ~new_n6306;
  assign new_n6308 = n401 & n9915;
  assign new_n6309 = new_n6113 & new_n6308;
  assign new_n6310 = ~new_n6307 & ~new_n6309;
  assign new_n6311 = ~new_n6304 & ~new_n6310;
  assign new_n6312 = new_n6304 & new_n6310;
  assign new_n6313 = ~new_n6311 & ~new_n6312;
  assign new_n6314 = n767 & n3832;
  assign new_n6315 = ~new_n6115 & ~new_n6314;
  assign new_n6316 = new_n6115 & new_n6314;
  assign new_n6317 = ~new_n6315 & ~new_n6316;
  assign new_n6318 = ~new_n6313 & new_n6317;
  assign new_n6319 = new_n6313 & ~new_n6317;
  assign new_n6320 = ~new_n6318 & ~new_n6319;
  assign new_n6321 = n1165 & n3178;
  assign new_n6322 = n2882 & n10168;
  assign new_n6323 = n4357 & n12592;
  assign new_n6324 = ~new_n6322 & ~new_n6323;
  assign new_n6325 = new_n6322 & new_n6323;
  assign new_n6326 = ~new_n6324 & ~new_n6325;
  assign new_n6327 = ~new_n6321 & ~new_n6326;
  assign new_n6328 = new_n6321 & new_n6326;
  assign new_n6329 = ~new_n6327 & ~new_n6328;
  assign new_n6330 = ~new_n6118 & new_n6121;
  assign new_n6331 = ~new_n6117 & ~new_n6330;
  assign new_n6332 = ~new_n6329 & ~new_n6331;
  assign new_n6333_1 = new_n6329 & new_n6331;
  assign new_n6334 = ~new_n6332 & ~new_n6333_1;
  assign new_n6335 = new_n6320 & new_n6334;
  assign new_n6336 = ~new_n6320 & ~new_n6334;
  assign new_n6337 = ~new_n6335 & ~new_n6336;
  assign new_n6338 = ~new_n6303 & new_n6337;
  assign new_n6339 = new_n6303 & ~new_n6337;
  assign new_n6340 = ~new_n6338 & ~new_n6339;
  assign new_n6341 = new_n6135 & new_n6340;
  assign new_n6342 = ~new_n6135 & ~new_n6340;
  assign new_n6343 = ~new_n6341 & ~new_n6342;
  assign new_n6344 = ~new_n6138 & ~new_n6142;
  assign new_n6345 = new_n6343 & ~new_n6344;
  assign new_n6346 = ~new_n6343 & new_n6344;
  assign new_n6347 = ~new_n6345 & ~new_n6346;
  assign new_n6348 = ~new_n6166 & ~new_n6170;
  assign new_n6349 = new_n6150 & new_n6348;
  assign new_n6350 = ~new_n6150 & ~new_n6348;
  assign new_n6351 = ~new_n6167 & new_n6350;
  assign new_n6352 = ~new_n6349 & ~new_n6351;
  assign new_n6353 = ~new_n6158 & ~new_n6162;
  assign new_n6354 = ~new_n6159 & ~new_n6353;
  assign new_n6355 = n9 & n2174;
  assign new_n6356 = n3112 & n5031;
  assign new_n6357 = ~new_n6144 & ~new_n6356;
  assign new_n6358 = n5031 & new_n6144;
  assign new_n6359 = ~new_n6357 & ~new_n6358;
  assign new_n6360 = ~new_n6355 & new_n6359;
  assign new_n6361 = new_n6355 & ~new_n6359;
  assign new_n6362 = ~new_n6360 & ~new_n6361;
  assign new_n6363 = new_n6354 & new_n6362;
  assign new_n6364 = n2590 & n9887;
  assign new_n6365 = n4335 & n11061;
  assign new_n6366 = n8233 & n8768;
  assign new_n6367 = ~new_n6365 & ~new_n6366;
  assign new_n6368 = new_n6365 & new_n6366;
  assign new_n6369 = ~new_n6367 & ~new_n6368;
  assign new_n6370 = ~new_n6364 & ~new_n6369;
  assign new_n6371 = new_n6364 & new_n6369;
  assign new_n6372 = ~new_n6370 & ~new_n6371;
  assign new_n6373 = n497 & n2592;
  assign new_n6374 = new_n6156 & new_n6373;
  assign new_n6375 = ~new_n6156 & ~new_n6373;
  assign new_n6376 = ~new_n6374 & ~new_n6375;
  assign new_n6377 = ~new_n6372 & ~new_n6376;
  assign new_n6378 = new_n6372 & ~new_n6375;
  assign new_n6379 = ~new_n6374 & new_n6378;
  assign new_n6380 = ~new_n6377 & ~new_n6379;
  assign new_n6381 = new_n6363 & ~new_n6380;
  assign new_n6382 = ~new_n6354 & ~new_n6362;
  assign new_n6383 = ~new_n6380 & ~new_n6382;
  assign new_n6384 = ~new_n6363 & ~new_n6383;
  assign new_n6385 = new_n6380 & new_n6382;
  assign new_n6386 = new_n6384 & ~new_n6385;
  assign new_n6387 = ~new_n6381 & ~new_n6386;
  assign new_n6388 = new_n6352 & ~new_n6387;
  assign new_n6389 = ~new_n6352 & new_n6387;
  assign new_n6390 = ~new_n6388 & ~new_n6389;
  assign new_n6391 = new_n6174 & ~new_n6390;
  assign new_n6392_1 = ~new_n6174 & new_n6390;
  assign new_n6393 = ~new_n6391 & ~new_n6392_1;
  assign new_n6394 = ~new_n6177 & ~new_n6181;
  assign new_n6395 = new_n6393 & ~new_n6394;
  assign new_n6396 = ~new_n6393 & new_n6394;
  assign new_n6397 = ~new_n6395 & ~new_n6396;
  assign new_n6398 = new_n6347 & new_n6397;
  assign new_n6399 = ~new_n6347 & ~new_n6397;
  assign new_n6400 = ~new_n6398 & ~new_n6399;
  assign new_n6401 = ~new_n6184 & ~new_n6187;
  assign new_n6402 = ~new_n6183 & ~new_n6401;
  assign new_n6403 = ~new_n6400 & ~new_n6402;
  assign new_n6404 = new_n6400 & new_n6402;
  assign new_n6405 = ~new_n6403 & ~new_n6404;
  assign new_n6406 = new_n6298 & ~new_n6405;
  assign new_n6407 = ~new_n6298 & new_n6405;
  assign new_n6408 = ~new_n6406 & ~new_n6407;
  assign new_n6409_1 = new_n6195 & new_n6408;
  assign new_n6410 = ~new_n6195 & ~new_n6408;
  assign new_n6411 = ~new_n6409_1 & ~new_n6410;
  assign new_n6412 = new_n6248 & ~new_n6411;
  assign new_n6413 = ~new_n6248 & new_n6411;
  assign new_n6414 = ~new_n6060 & new_n6197;
  assign new_n6415 = ~new_n6061 & ~new_n6414;
  assign new_n6416 = ~new_n6413 & ~new_n6415;
  assign new_n6417 = ~new_n6412 & ~new_n6416;
  assign new_n6418 = ~new_n6243 & ~new_n6246;
  assign new_n6419 = ~new_n6391 & ~new_n6395;
  assign new_n6420 = new_n6418 & new_n6419;
  assign new_n6421 = ~new_n6418 & ~new_n6419;
  assign new_n6422 = ~new_n6420 & ~new_n6421;
  assign new_n6423 = ~new_n6205 & ~new_n6239;
  assign new_n6424 = ~new_n6203 & ~new_n6423;
  assign new_n6425 = ~new_n6374 & ~new_n6378;
  assign new_n6426 = new_n6364 & ~new_n6367;
  assign new_n6427 = ~new_n6368 & ~new_n6426;
  assign new_n6428 = n4006 & n6668;
  assign new_n6429 = n2758 & n7812;
  assign new_n6430 = n3641 & n7772;
  assign new_n6431 = new_n6429 & ~new_n6430;
  assign new_n6432 = ~new_n6429 & new_n6430;
  assign new_n6433 = ~new_n6431 & ~new_n6432;
  assign new_n6434_1 = new_n6428 & ~new_n6433;
  assign new_n6435 = ~new_n6428 & new_n6433;
  assign new_n6436 = ~new_n6434_1 & ~new_n6435;
  assign new_n6437 = ~new_n6427 & new_n6436;
  assign new_n6438 = new_n6427 & ~new_n6436;
  assign new_n6439 = ~new_n6437 & ~new_n6438;
  assign new_n6440 = new_n6425 & new_n6439;
  assign new_n6441 = ~new_n6425 & ~new_n6439;
  assign new_n6442 = ~new_n6440 & ~new_n6441;
  assign new_n6443 = new_n6424 & new_n6442;
  assign new_n6444 = ~new_n6424 & ~new_n6442;
  assign new_n6445 = ~new_n6443 & ~new_n6444;
  assign new_n6446 = ~new_n6320 & ~new_n6332;
  assign new_n6447 = ~new_n6333_1 & ~new_n6446;
  assign new_n6448 = new_n6313 & ~new_n6315;
  assign new_n6449 = ~new_n6316 & ~new_n6448;
  assign new_n6450 = new_n6304 & ~new_n6307;
  assign new_n6451 = ~new_n6309 & ~new_n6450;
  assign new_n6452 = n4357 & n10168;
  assign new_n6453 = n1165 & n12592;
  assign new_n6454 = ~new_n6452 & new_n6453;
  assign new_n6455 = new_n6452 & ~new_n6453;
  assign new_n6456 = ~new_n6454 & ~new_n6455;
  assign new_n6457 = new_n6451 & ~new_n6456;
  assign new_n6458 = ~new_n6451 & new_n6456;
  assign new_n6459 = ~new_n6457 & ~new_n6458;
  assign new_n6460 = ~new_n6449 & new_n6459;
  assign new_n6461 = new_n6449 & ~new_n6459;
  assign new_n6462 = ~new_n6460 & ~new_n6461;
  assign new_n6463 = new_n6447 & new_n6462;
  assign new_n6464 = ~new_n6447 & ~new_n6462;
  assign new_n6465 = ~new_n6463 & ~new_n6464;
  assign new_n6466 = n2174 & n2592;
  assign new_n6467 = n3591 & n8466;
  assign new_n6468 = ~new_n6466 & new_n6467;
  assign new_n6469 = new_n6466 & ~new_n6467;
  assign new_n6470 = ~new_n6468 & ~new_n6469;
  assign new_n6471 = n497 & n2590;
  assign new_n6472 = new_n6356 & ~new_n6471;
  assign new_n6473 = ~new_n6356 & new_n6471;
  assign new_n6474 = ~new_n6472 & ~new_n6473;
  assign new_n6475 = ~new_n6470 & ~new_n6474;
  assign new_n6476 = new_n6470 & new_n6474;
  assign new_n6477 = ~new_n6475 & ~new_n6476;
  assign new_n6478 = n9 & n3112;
  assign new_n6479 = n4998 & n8233;
  assign new_n6480 = ~new_n6478 & new_n6479;
  assign new_n6481 = new_n6478 & ~new_n6479;
  assign new_n6482 = ~new_n6480 & ~new_n6481;
  assign new_n6483 = n4335 & n8768;
  assign new_n6484 = n9887 & n11061;
  assign new_n6485 = ~new_n6483 & ~new_n6484;
  assign new_n6486 = new_n6483 & new_n6484;
  assign new_n6487 = ~new_n6485 & ~new_n6486;
  assign new_n6488 = ~new_n6482 & new_n6487;
  assign new_n6489 = new_n6482 & ~new_n6487;
  assign new_n6490 = ~new_n6488 & ~new_n6489;
  assign new_n6491 = new_n6477 & new_n6490;
  assign new_n6492 = ~new_n6477 & ~new_n6490;
  assign new_n6493 = ~new_n6491 & ~new_n6492;
  assign new_n6494 = new_n6321 & ~new_n6324;
  assign new_n6495 = ~new_n6325 & ~new_n6494;
  assign new_n6496 = ~new_n6493 & new_n6495;
  assign new_n6497 = new_n6493 & ~new_n6495;
  assign new_n6498 = ~new_n6496 & ~new_n6497;
  assign new_n6499 = ~new_n6465 & ~new_n6498;
  assign new_n6500 = new_n6465 & new_n6498;
  assign new_n6501 = ~new_n6499 & ~new_n6500;
  assign new_n6502 = ~new_n6351 & new_n6387;
  assign new_n6503 = ~new_n6349 & ~new_n6502;
  assign new_n6504 = new_n6384 & ~new_n6503;
  assign new_n6505 = ~new_n6384 & new_n6503;
  assign new_n6506 = ~new_n6504 & ~new_n6505;
  assign new_n6507 = ~new_n6501 & new_n6506;
  assign new_n6508 = new_n6501 & ~new_n6506;
  assign new_n6509 = ~new_n6507 & ~new_n6508;
  assign new_n6510 = ~new_n6445 & new_n6509;
  assign new_n6511 = new_n6445 & ~new_n6509;
  assign new_n6512 = ~new_n6510 & ~new_n6511;
  assign new_n6513 = ~new_n6422 & ~new_n6512;
  assign new_n6514 = new_n6422 & new_n6512;
  assign new_n6515 = ~new_n6513 & ~new_n6514;
  assign new_n6516 = new_n6195 & ~new_n6406;
  assign new_n6517 = ~new_n6407 & ~new_n6516;
  assign new_n6518 = ~new_n6341 & ~new_n6345;
  assign new_n6519 = ~new_n6301_1 & ~new_n6337;
  assign new_n6520 = ~new_n6302 & ~new_n6519;
  assign new_n6521 = n951 & n8332;
  assign new_n6522 = n767 & n2882;
  assign new_n6523 = new_n6521 & ~new_n6522;
  assign new_n6524 = ~new_n6521 & new_n6522;
  assign new_n6525 = ~new_n6523 & ~new_n6524;
  assign new_n6526 = n3832 & n11537;
  assign new_n6527 = ~new_n6308 & ~new_n6526;
  assign new_n6528 = new_n6308 & new_n6526;
  assign new_n6529 = ~new_n6527 & ~new_n6528;
  assign new_n6530 = ~new_n6525 & new_n6529;
  assign new_n6531 = new_n6525 & ~new_n6529;
  assign new_n6532 = ~new_n6530 & ~new_n6531;
  assign new_n6533 = n4419 & n10063;
  assign new_n6534 = n3178 & n10874;
  assign new_n6535 = ~new_n6533 & new_n6534;
  assign new_n6536 = new_n6533 & ~new_n6534;
  assign new_n6537 = ~new_n6535 & ~new_n6536;
  assign new_n6538 = ~new_n6532 & new_n6537;
  assign new_n6539 = new_n6532 & ~new_n6537;
  assign new_n6540 = ~new_n6538 & ~new_n6539;
  assign new_n6541 = ~new_n6270 & ~new_n6280;
  assign new_n6542 = ~new_n6269 & ~new_n6541;
  assign new_n6543 = ~new_n6266 & ~new_n6283;
  assign new_n6544 = ~new_n6265 & ~new_n6543;
  assign new_n6545 = new_n6542 & new_n6544;
  assign new_n6546 = ~new_n6542 & ~new_n6544;
  assign new_n6547 = ~new_n6545 & ~new_n6546;
  assign new_n6548 = ~new_n6540 & new_n6547;
  assign new_n6549 = new_n6540 & ~new_n6547;
  assign new_n6550 = ~new_n6548 & ~new_n6549;
  assign new_n6551 = new_n6520 & ~new_n6550;
  assign new_n6552 = ~new_n6520 & new_n6550;
  assign new_n6553 = ~new_n6551 & ~new_n6552;
  assign new_n6554 = n2068 & n3677;
  assign new_n6555 = n7729 & n12348;
  assign new_n6556 = ~new_n6554 & new_n6555;
  assign new_n6557 = new_n6554 & ~new_n6555;
  assign new_n6558 = ~new_n6556 & ~new_n6557;
  assign new_n6559 = new_n6272 & ~new_n6275;
  assign new_n6560 = ~new_n6276 & ~new_n6559;
  assign new_n6561 = ~new_n6558 & new_n6560;
  assign new_n6562 = new_n6558 & ~new_n6560;
  assign new_n6563 = ~new_n6561 & ~new_n6562;
  assign new_n6564 = n6937 & n11324;
  assign new_n6565 = new_n6254 & ~new_n6257;
  assign new_n6566 = ~new_n6258 & ~new_n6565;
  assign new_n6567 = new_n6564 & new_n6566;
  assign new_n6568 = ~new_n6564 & ~new_n6566;
  assign new_n6569 = ~new_n6567 & ~new_n6568;
  assign new_n6570 = new_n6563 & new_n6569;
  assign new_n6571 = ~new_n6563 & ~new_n6569;
  assign new_n6572 = ~new_n6570 & ~new_n6571;
  assign new_n6573 = ~new_n6553 & new_n6572;
  assign new_n6574 = new_n6553 & ~new_n6572;
  assign new_n6575 = ~new_n6573 & ~new_n6574;
  assign new_n6576 = new_n6518 & new_n6575;
  assign new_n6577 = ~new_n6518 & ~new_n6575;
  assign new_n6578 = ~new_n6576 & ~new_n6577;
  assign new_n6579 = ~new_n6293 & ~new_n6296;
  assign new_n6580 = n4452 & n10408;
  assign new_n6581 = ~new_n6219 & new_n6236;
  assign new_n6582 = ~new_n6218 & ~new_n6581;
  assign new_n6583 = ~new_n6223 & ~new_n6233;
  assign new_n6584 = ~new_n6222 & ~new_n6583;
  assign new_n6585 = n8230 & n12306;
  assign new_n6586_1 = n2458 & n4748;
  assign new_n6587 = ~new_n6585 & ~new_n6586_1;
  assign new_n6588 = new_n6585 & new_n6586_1;
  assign new_n6589 = ~new_n6587 & ~new_n6588;
  assign new_n6590 = n7715 & n9187;
  assign new_n6591 = n1231 & n7529;
  assign new_n6592 = new_n6590 & ~new_n6591;
  assign new_n6593 = ~new_n6590 & new_n6591;
  assign new_n6594 = ~new_n6592 & ~new_n6593;
  assign new_n6595 = ~new_n6589 & ~new_n6594;
  assign new_n6596 = new_n6589 & new_n6594;
  assign new_n6597 = ~new_n6595 & ~new_n6596;
  assign new_n6598 = new_n6225 & ~new_n6228;
  assign new_n6599 = ~new_n6229 & ~new_n6598;
  assign new_n6600 = new_n6207 & ~new_n6210;
  assign new_n6601 = ~new_n6211 & ~new_n6600;
  assign new_n6602 = ~new_n6599 & new_n6601;
  assign new_n6603 = new_n6599 & ~new_n6601;
  assign new_n6604 = ~new_n6602 & ~new_n6603;
  assign new_n6605 = new_n6597 & new_n6604;
  assign new_n6606 = ~new_n6597 & ~new_n6604;
  assign new_n6607 = ~new_n6605 & ~new_n6606;
  assign new_n6608 = ~new_n6584 & new_n6607;
  assign new_n6609 = new_n6584 & ~new_n6607;
  assign new_n6610 = ~new_n6608 & ~new_n6609;
  assign new_n6611 = ~new_n6582 & ~new_n6610;
  assign new_n6612 = new_n6582 & new_n6610;
  assign new_n6613 = ~new_n6611 & ~new_n6612;
  assign new_n6614 = ~new_n6580 & new_n6613;
  assign new_n6615 = new_n6580 & ~new_n6613;
  assign new_n6616 = ~new_n6614 & ~new_n6615;
  assign new_n6617 = n603 & n9216;
  assign new_n6618 = n1724 & n8183;
  assign new_n6619 = new_n6617 & ~new_n6618;
  assign new_n6620 = ~new_n6617 & new_n6618;
  assign new_n6621 = ~new_n6619 & ~new_n6620;
  assign new_n6622 = n10606 & n10657;
  assign new_n6623 = n10142 & n12965;
  assign new_n6624 = ~new_n6622 & ~new_n6623;
  assign new_n6625 = new_n6622 & new_n6623;
  assign new_n6626 = ~new_n6624 & ~new_n6625;
  assign new_n6627 = ~new_n6621 & new_n6626;
  assign new_n6628 = new_n6621 & ~new_n6626;
  assign new_n6629 = ~new_n6627 & ~new_n6628;
  assign new_n6630 = ~new_n6288 & new_n6629;
  assign new_n6631 = new_n6288 & ~new_n6629;
  assign new_n6632 = ~new_n6630 & ~new_n6631;
  assign new_n6633 = ~new_n6616 & ~new_n6632;
  assign new_n6634 = new_n6616 & new_n6632;
  assign new_n6635 = ~new_n6633 & ~new_n6634;
  assign new_n6636 = ~new_n6579 & ~new_n6635;
  assign new_n6637 = new_n6579 & new_n6635;
  assign new_n6638 = ~new_n6636 & ~new_n6637;
  assign new_n6639 = ~new_n6578 & new_n6638;
  assign new_n6640 = new_n6578 & ~new_n6638;
  assign new_n6641 = ~new_n6639 & ~new_n6640;
  assign new_n6642 = ~new_n6355 & ~new_n6358;
  assign new_n6643 = ~new_n6357 & ~new_n6642;
  assign new_n6644 = ~new_n6399 & ~new_n6402;
  assign new_n6645 = ~new_n6398 & ~new_n6644;
  assign new_n6646 = new_n6643 & new_n6645;
  assign new_n6647 = ~new_n6643 & ~new_n6645;
  assign new_n6648 = ~new_n6646 & ~new_n6647;
  assign new_n6649 = new_n6641 & ~new_n6648;
  assign new_n6650 = ~new_n6641 & new_n6648;
  assign new_n6651 = ~new_n6649 & ~new_n6650;
  assign new_n6652 = ~new_n6517 & ~new_n6651;
  assign new_n6653 = new_n6517 & new_n6651;
  assign new_n6654 = ~new_n6652 & ~new_n6653;
  assign new_n6655_1 = ~new_n6515 & new_n6654;
  assign new_n6656 = new_n6515 & ~new_n6654;
  assign new_n6657 = ~new_n6655_1 & ~new_n6656;
  assign new_n6658 = ~new_n6417 & ~new_n6657;
  assign new_n6659 = new_n6417 & new_n6657;
  assign n1112 = ~new_n6658 & ~new_n6659;
  assign new_n6661 = n2339 & n4114;
  assign new_n6662 = n9570 & n11665;
  assign new_n6663 = ~new_n6661 & ~new_n6662;
  assign new_n6664 = new_n6661 & new_n6662;
  assign new_n6665 = ~new_n6663 & ~new_n6664;
  assign new_n6666 = n2777 & n12482;
  assign new_n6667 = n7720 & n10642;
  assign new_n6668_1 = n287 & n937;
  assign new_n6669 = ~new_n6667 & ~new_n6668_1;
  assign new_n6670 = new_n6667 & new_n6668_1;
  assign new_n6671 = ~new_n6669 & ~new_n6670;
  assign new_n6672 = ~new_n6666 & ~new_n6671;
  assign new_n6673 = new_n6666 & new_n6671;
  assign new_n6674 = ~new_n6672 & ~new_n6673;
  assign new_n6675 = n11665 & n12482;
  assign new_n6676 = n2777 & n7720;
  assign new_n6677 = new_n6675 & new_n6676;
  assign new_n6678 = n287 & n10642;
  assign new_n6679 = ~new_n6675 & ~new_n6676;
  assign new_n6680 = new_n6678 & ~new_n6679;
  assign new_n6681 = ~new_n6677 & ~new_n6680;
  assign new_n6682 = ~new_n6674 & ~new_n6681;
  assign new_n6683_1 = new_n6674 & new_n6681;
  assign new_n6684 = ~new_n6682 & ~new_n6683_1;
  assign new_n6685 = ~new_n6665 & new_n6684;
  assign new_n6686 = new_n6665 & ~new_n6684;
  assign new_n6687 = ~new_n6685 & ~new_n6686;
  assign new_n6688 = n4114 & n9570;
  assign new_n6689 = new_n5345 & ~new_n5348;
  assign new_n6690 = ~new_n5349 & ~new_n6689;
  assign new_n6691 = ~new_n6688 & new_n6690;
  assign new_n6692 = new_n6688 & ~new_n6690;
  assign new_n6693 = ~new_n6677 & ~new_n6679;
  assign new_n6694 = ~new_n6678 & ~new_n6693;
  assign new_n6695 = new_n6678 & new_n6693;
  assign new_n6696 = ~new_n6694 & ~new_n6695;
  assign new_n6697 = ~new_n6692 & ~new_n6696;
  assign new_n6698 = ~new_n6691 & ~new_n6697;
  assign new_n6699 = new_n6687 & ~new_n6698;
  assign new_n6700 = ~new_n6687 & new_n6698;
  assign new_n6701 = ~new_n6699 & ~new_n6700;
  assign new_n6702 = n2339 & n5671;
  assign new_n6703 = ~new_n6691 & ~new_n6692;
  assign new_n6704 = ~new_n6696 & ~new_n6703;
  assign new_n6705 = new_n6696 & new_n6703;
  assign new_n6706 = ~new_n6704 & ~new_n6705;
  assign new_n6707 = ~new_n6702 & ~new_n6706;
  assign new_n6708 = new_n6702 & new_n6706;
  assign new_n6709 = ~new_n5342 & ~new_n5353;
  assign new_n6710 = ~new_n5343 & ~new_n6709;
  assign new_n6711 = ~new_n6708 & new_n6710;
  assign new_n6712 = ~new_n6707 & ~new_n6711;
  assign new_n6713 = ~new_n6701 & new_n6712;
  assign new_n6714 = ~new_n6685 & new_n6698;
  assign new_n6715 = ~new_n6664 & ~new_n6714;
  assign new_n6716 = ~new_n6686 & new_n6715;
  assign new_n6717 = new_n6664 & new_n6714;
  assign new_n6718 = ~new_n6716 & ~new_n6717;
  assign new_n6719 = n2339 & n11665;
  assign new_n6720 = n1307 & n4114;
  assign new_n6721 = ~new_n6719 & ~new_n6720;
  assign new_n6722 = new_n6719 & new_n6720;
  assign new_n6723 = ~new_n6721 & ~new_n6722;
  assign new_n6724 = ~new_n6673 & new_n6681;
  assign new_n6725 = ~new_n6672 & ~new_n6724;
  assign new_n6726 = new_n6723 & new_n6725;
  assign new_n6727 = ~new_n6723 & ~new_n6725;
  assign new_n6728 = ~new_n6726 & ~new_n6727;
  assign new_n6729 = n2777 & n9570;
  assign new_n6730 = ~new_n6670 & ~new_n6729;
  assign new_n6731 = new_n6670 & new_n6729;
  assign new_n6732 = ~new_n6730 & ~new_n6731;
  assign new_n6733 = n287 & n12605;
  assign new_n6734 = n937 & n7720;
  assign new_n6735 = n10642 & n12482;
  assign new_n6736 = ~new_n6734 & ~new_n6735;
  assign new_n6737 = new_n6734 & new_n6735;
  assign new_n6738 = ~new_n6736 & ~new_n6737;
  assign new_n6739 = new_n6733 & ~new_n6738;
  assign new_n6740 = ~new_n6733 & new_n6738;
  assign new_n6741 = ~new_n6739 & ~new_n6740;
  assign new_n6742 = new_n6732 & ~new_n6741;
  assign new_n6743 = ~new_n6732 & new_n6741;
  assign new_n6744 = ~new_n6742 & ~new_n6743;
  assign new_n6745 = new_n6728 & ~new_n6744;
  assign new_n6746 = ~new_n6728 & new_n6744;
  assign new_n6747 = ~new_n6745 & ~new_n6746;
  assign new_n6748 = new_n6718 & ~new_n6747;
  assign new_n6749 = ~new_n6718 & new_n6747;
  assign new_n6750 = ~new_n6748 & ~new_n6749;
  assign new_n6751 = new_n6713 & new_n6750;
  assign new_n6752 = ~new_n6713 & ~new_n6750;
  assign new_n6753 = ~new_n6751 & ~new_n6752;
  assign new_n6754 = n1307 & n5671;
  assign new_n6755 = new_n6701 & ~new_n6712;
  assign new_n6756 = ~new_n6713 & ~new_n6755;
  assign new_n6757 = new_n6754 & new_n6756;
  assign new_n6758 = ~new_n6707 & ~new_n6708;
  assign new_n6759 = ~new_n6710 & ~new_n6758;
  assign new_n6760 = new_n6710 & new_n6758;
  assign new_n6761 = ~new_n6759 & ~new_n6760;
  assign new_n6762 = new_n5358 & ~new_n6761;
  assign new_n6763 = ~new_n6754 & ~new_n6756;
  assign new_n6764 = ~new_n6757 & ~new_n6763;
  assign new_n6765 = new_n6762 & new_n6764;
  assign new_n6766 = ~new_n6757 & ~new_n6765;
  assign new_n6767 = new_n6753 & ~new_n6766;
  assign new_n6768 = ~new_n6751 & ~new_n6767;
  assign new_n6769 = n3409 & n8308;
  assign new_n6770 = n5568 & n7113;
  assign new_n6771 = ~new_n6769 & ~new_n6770;
  assign new_n6772 = new_n6769 & new_n6770;
  assign new_n6773 = ~new_n6771 & ~new_n6772;
  assign new_n6774 = n5214 & n10594;
  assign new_n6775 = n6168 & n10451;
  assign new_n6776 = n2771 & n9093;
  assign new_n6777 = new_n6775 & new_n6776;
  assign new_n6778 = ~new_n6775 & ~new_n6776;
  assign new_n6779 = ~new_n6777 & ~new_n6778;
  assign new_n6780 = new_n6774 & new_n6779;
  assign new_n6781 = ~new_n6774 & ~new_n6779;
  assign new_n6782 = ~new_n6780 & ~new_n6781;
  assign new_n6783 = n8308 & n10594;
  assign new_n6784 = n5214 & n9093;
  assign new_n6785 = new_n6783 & new_n6784;
  assign new_n6786 = ~new_n6783 & ~new_n6784;
  assign new_n6787 = n2771 & n10451;
  assign new_n6788 = ~new_n6786 & new_n6787;
  assign new_n6789 = ~new_n6785 & ~new_n6788;
  assign new_n6790 = ~new_n6782 & ~new_n6789;
  assign new_n6791 = new_n6782 & new_n6789;
  assign new_n6792 = ~new_n6790 & ~new_n6791;
  assign new_n6793 = new_n6773 & ~new_n6792;
  assign new_n6794 = ~new_n6773 & new_n6792;
  assign new_n6795 = ~new_n6793 & ~new_n6794;
  assign new_n6796 = n3409 & n5568;
  assign new_n6797 = new_n5303 & ~new_n5306;
  assign new_n6798 = ~new_n5307 & ~new_n6797;
  assign new_n6799 = ~new_n6796 & new_n6798;
  assign new_n6800 = new_n6796 & ~new_n6798;
  assign new_n6801 = ~new_n6785 & ~new_n6786;
  assign new_n6802 = ~new_n6787 & ~new_n6801;
  assign new_n6803 = new_n6787 & new_n6801;
  assign new_n6804 = ~new_n6802 & ~new_n6803;
  assign new_n6805 = ~new_n6800 & ~new_n6804;
  assign new_n6806 = ~new_n6799 & ~new_n6805;
  assign new_n6807 = new_n6795 & ~new_n6806;
  assign new_n6808 = ~new_n6795 & new_n6806;
  assign new_n6809 = ~new_n6807 & ~new_n6808;
  assign new_n6810 = n3006 & n7113;
  assign new_n6811 = ~new_n6799 & ~new_n6800;
  assign new_n6812 = ~new_n6804 & ~new_n6811;
  assign new_n6813 = new_n6804 & new_n6811;
  assign new_n6814 = ~new_n6812 & ~new_n6813;
  assign new_n6815 = ~new_n6810 & ~new_n6814;
  assign new_n6816 = new_n6810 & new_n6814;
  assign new_n6817 = ~new_n5300 & ~new_n5311;
  assign new_n6818_1 = ~new_n5301 & ~new_n6817;
  assign new_n6819 = ~new_n6816 & new_n6818_1;
  assign new_n6820 = ~new_n6815 & ~new_n6819;
  assign new_n6821 = ~new_n6809 & new_n6820;
  assign new_n6822 = ~new_n6794 & new_n6806;
  assign new_n6823 = new_n6772 & new_n6822;
  assign new_n6824 = ~new_n6772 & ~new_n6822;
  assign new_n6825 = ~new_n6793 & new_n6824;
  assign new_n6826_1 = ~new_n6823 & ~new_n6825;
  assign new_n6827 = n7113 & n8308;
  assign new_n6828 = n499 & n3006;
  assign new_n6829 = n1302 & n5568;
  assign new_n6830 = ~new_n6828 & ~new_n6829;
  assign new_n6831 = new_n6828 & new_n6829;
  assign new_n6832 = ~new_n6830 & ~new_n6831;
  assign new_n6833 = new_n6827 & ~new_n6832;
  assign new_n6834 = ~new_n6827 & new_n6832;
  assign new_n6835 = ~new_n6833 & ~new_n6834;
  assign new_n6836 = ~new_n6780 & new_n6789;
  assign new_n6837 = ~new_n6781 & ~new_n6836;
  assign new_n6838 = ~new_n6835 & new_n6837;
  assign new_n6839 = new_n6835 & ~new_n6837;
  assign new_n6840 = ~new_n6838 & ~new_n6839;
  assign new_n6841 = n10451 & n11411;
  assign new_n6842 = n6168 & n9093;
  assign new_n6843_1 = n2771 & n10594;
  assign new_n6844 = ~new_n6842 & ~new_n6843_1;
  assign new_n6845 = new_n6842 & new_n6843_1;
  assign new_n6846 = ~new_n6844 & ~new_n6845;
  assign new_n6847 = new_n6841 & ~new_n6846;
  assign new_n6848 = ~new_n6841 & new_n6846;
  assign new_n6849 = ~new_n6847 & ~new_n6848;
  assign new_n6850 = n3409 & n5214;
  assign new_n6851 = new_n6777 & new_n6850;
  assign new_n6852 = ~new_n6777 & ~new_n6850;
  assign new_n6853 = ~new_n6851 & ~new_n6852;
  assign new_n6854 = ~new_n6849 & new_n6853;
  assign new_n6855 = new_n6849 & ~new_n6853;
  assign new_n6856 = ~new_n6854 & ~new_n6855;
  assign new_n6857 = ~new_n6840 & new_n6856;
  assign new_n6858 = new_n6840 & ~new_n6856;
  assign new_n6859 = ~new_n6857 & ~new_n6858;
  assign new_n6860 = ~new_n6826_1 & ~new_n6859;
  assign new_n6861 = new_n6826_1 & new_n6859;
  assign new_n6862_1 = ~new_n6860 & ~new_n6861;
  assign new_n6863 = new_n6821 & ~new_n6862_1;
  assign new_n6864 = n1302 & n3006;
  assign new_n6865 = new_n6809 & ~new_n6820;
  assign new_n6866 = ~new_n6821 & ~new_n6865;
  assign new_n6867 = new_n6864 & new_n6866;
  assign new_n6868 = ~new_n6815 & ~new_n6816;
  assign new_n6869 = new_n6818_1 & new_n6868;
  assign new_n6870 = ~new_n6818_1 & ~new_n6868;
  assign new_n6871 = ~new_n6869 & ~new_n6870;
  assign new_n6872 = new_n5316 & ~new_n6871;
  assign new_n6873 = ~new_n6864 & ~new_n6866;
  assign new_n6874 = ~new_n6867 & ~new_n6873;
  assign new_n6875 = new_n6872 & new_n6874;
  assign new_n6876 = ~new_n6867 & ~new_n6875;
  assign new_n6877 = ~new_n6821 & new_n6862_1;
  assign new_n6878 = ~new_n6863 & ~new_n6877;
  assign new_n6879 = ~new_n6876 & new_n6878;
  assign new_n6880 = ~new_n6863 & ~new_n6879;
  assign new_n6881 = new_n6768 & new_n6880;
  assign new_n6882 = ~new_n6768 & ~new_n6880;
  assign new_n6883 = ~new_n6881 & ~new_n6882;
  assign new_n6884 = n9300 & n13201;
  assign new_n6885 = n1198 & n13201;
  assign new_n6886 = n2057 & n2498;
  assign new_n6887 = new_n5366 & ~new_n5369;
  assign new_n6888 = ~new_n5370 & ~new_n6887;
  assign new_n6889 = new_n6886 & ~new_n6888;
  assign new_n6890 = ~new_n6886 & new_n6888;
  assign new_n6891 = ~new_n6889 & ~new_n6890;
  assign new_n6892 = n1364 & n11058;
  assign new_n6893 = n5586 & n5969;
  assign new_n6894 = n1007 & n4141;
  assign new_n6895 = ~new_n6893 & ~new_n6894;
  assign new_n6896 = new_n6893 & new_n6894;
  assign new_n6897 = ~new_n6895 & ~new_n6896;
  assign new_n6898 = new_n6892 & ~new_n6897;
  assign new_n6899 = ~new_n6892 & new_n6897;
  assign new_n6900 = ~new_n6898 & ~new_n6899;
  assign new_n6901 = ~new_n6891 & ~new_n6900;
  assign new_n6902 = new_n6891 & new_n6900;
  assign new_n6903 = ~new_n6901 & ~new_n6902;
  assign new_n6904 = ~new_n6885 & new_n6903;
  assign new_n6905 = new_n6885 & ~new_n6903;
  assign new_n6906 = ~new_n5364_1 & new_n5374;
  assign new_n6907 = ~new_n5363 & ~new_n6906;
  assign new_n6908 = ~new_n6905 & ~new_n6907;
  assign new_n6909 = ~new_n6904 & ~new_n6908;
  assign new_n6910 = n2498 & n5586;
  assign new_n6911 = n1198 & n2057;
  assign new_n6912 = new_n6910 & new_n6911;
  assign new_n6913 = ~new_n6910 & ~new_n6911;
  assign new_n6914 = ~new_n6912 & ~new_n6913;
  assign new_n6915 = n4141 & n5969;
  assign new_n6916 = n1007 & n1364;
  assign new_n6917 = n3669 & n11058;
  assign new_n6918 = ~new_n6916 & ~new_n6917;
  assign new_n6919 = new_n6916 & new_n6917;
  assign new_n6920 = ~new_n6918 & ~new_n6919;
  assign new_n6921 = ~new_n6915 & ~new_n6920;
  assign new_n6922 = new_n6915 & new_n6920;
  assign new_n6923 = ~new_n6921 & ~new_n6922;
  assign new_n6924 = new_n6892 & ~new_n6895;
  assign new_n6925 = ~new_n6896 & ~new_n6924;
  assign new_n6926 = ~new_n6923 & new_n6925;
  assign new_n6927 = new_n6923 & ~new_n6925;
  assign new_n6928 = ~new_n6926 & ~new_n6927;
  assign new_n6929 = ~new_n6914 & ~new_n6928;
  assign new_n6930 = new_n6914 & new_n6928;
  assign new_n6931 = ~new_n6929 & ~new_n6930;
  assign new_n6932 = ~new_n6890 & ~new_n6900;
  assign new_n6933 = ~new_n6889 & ~new_n6932;
  assign new_n6934 = ~new_n6931 & ~new_n6933;
  assign new_n6935 = new_n6931 & new_n6933;
  assign new_n6936 = ~new_n6934 & ~new_n6935;
  assign new_n6937_1 = new_n6909 & ~new_n6936;
  assign new_n6938 = ~new_n6909 & new_n6936;
  assign new_n6939 = ~new_n6937_1 & ~new_n6938;
  assign new_n6940 = new_n6884 & new_n6939;
  assign new_n6941 = ~new_n6904 & ~new_n6905;
  assign new_n6942 = ~new_n6907 & ~new_n6941;
  assign new_n6943 = new_n6907 & new_n6941;
  assign new_n6944 = ~new_n6942 & ~new_n6943;
  assign new_n6945 = new_n5378 & new_n6944;
  assign new_n6946 = ~new_n6884 & ~new_n6939;
  assign new_n6947 = ~new_n6940 & ~new_n6946;
  assign new_n6948 = new_n6945 & new_n6947;
  assign new_n6949 = ~new_n6940 & ~new_n6948;
  assign new_n6950 = ~new_n6929 & ~new_n6933;
  assign new_n6951 = new_n6912 & new_n6950;
  assign new_n6952 = ~new_n6912 & ~new_n6950;
  assign new_n6953 = ~new_n6930 & new_n6952;
  assign new_n6954 = ~new_n6951 & ~new_n6953;
  assign new_n6955 = ~new_n6921 & ~new_n6925;
  assign new_n6956 = ~new_n6922 & ~new_n6955;
  assign new_n6957 = n1198 & n5586;
  assign new_n6958 = n11574 & n13201;
  assign new_n6959 = n2057 & n9300;
  assign new_n6960 = ~new_n6958 & ~new_n6959;
  assign new_n6961 = new_n6958 & new_n6959;
  assign new_n6962 = ~new_n6960 & ~new_n6961;
  assign new_n6963 = new_n6957 & ~new_n6962;
  assign new_n6964 = ~new_n6957 & new_n6962;
  assign new_n6965 = ~new_n6963 & ~new_n6964;
  assign new_n6966 = new_n6956 & new_n6965;
  assign new_n6967 = ~new_n6956 & ~new_n6965;
  assign new_n6968 = ~new_n6966 & ~new_n6967;
  assign new_n6969 = n2498 & n4141;
  assign new_n6970 = ~new_n6919 & ~new_n6969;
  assign new_n6971 = new_n6919 & new_n6969;
  assign new_n6972 = ~new_n6970 & ~new_n6971;
  assign new_n6973 = n5470 & n11058;
  assign new_n6974 = n1007 & n3669;
  assign new_n6975 = n1364 & n5969;
  assign new_n6976 = ~new_n6974 & ~new_n6975;
  assign new_n6977 = new_n6974 & new_n6975;
  assign new_n6978 = ~new_n6976 & ~new_n6977;
  assign new_n6979 = new_n6973 & ~new_n6978;
  assign new_n6980 = ~new_n6973 & new_n6978;
  assign new_n6981 = ~new_n6979 & ~new_n6980;
  assign new_n6982 = ~new_n6972 & new_n6981;
  assign new_n6983 = new_n6972 & ~new_n6981;
  assign new_n6984 = ~new_n6982 & ~new_n6983;
  assign new_n6985 = new_n6968 & new_n6984;
  assign new_n6986 = ~new_n6968 & ~new_n6984;
  assign new_n6987 = ~new_n6985 & ~new_n6986;
  assign new_n6988 = new_n6954 & ~new_n6987;
  assign new_n6989 = ~new_n6954 & new_n6987;
  assign new_n6990 = ~new_n6988 & ~new_n6989;
  assign new_n6991 = new_n6937_1 & ~new_n6990;
  assign new_n6992 = ~new_n6937_1 & new_n6990;
  assign new_n6993 = ~new_n6991 & ~new_n6992;
  assign new_n6994 = ~new_n6949 & new_n6993;
  assign new_n6995 = new_n6949 & ~new_n6993;
  assign new_n6996 = ~new_n6994 & ~new_n6995;
  assign new_n6997 = ~new_n6753 & new_n6766;
  assign new_n6998 = ~new_n6767 & ~new_n6997;
  assign new_n6999 = new_n6996 & new_n6998;
  assign new_n7000 = ~new_n6996 & ~new_n6998;
  assign new_n7001 = ~new_n6945 & ~new_n6947;
  assign new_n7002 = ~new_n6948 & ~new_n7001;
  assign new_n7003 = ~new_n6762 & ~new_n6764;
  assign new_n7004 = ~new_n6765 & ~new_n7003;
  assign new_n7005 = new_n7002 & new_n7004;
  assign new_n7006 = ~new_n7002 & ~new_n7004;
  assign new_n7007 = ~new_n5378 & ~new_n6944;
  assign new_n7008 = ~new_n6945 & ~new_n7007;
  assign new_n7009 = ~new_n5358 & new_n6761;
  assign new_n7010 = ~new_n6762 & ~new_n7009;
  assign new_n7011 = new_n7008 & new_n7010;
  assign new_n7012 = ~new_n7008 & ~new_n7010;
  assign new_n7013 = ~new_n5382 & ~new_n5385;
  assign new_n7014 = ~new_n5381 & ~new_n7013;
  assign new_n7015 = ~new_n7012 & ~new_n7014;
  assign new_n7016 = ~new_n7011 & ~new_n7015;
  assign new_n7017 = ~new_n7006 & ~new_n7016;
  assign new_n7018 = ~new_n7005 & ~new_n7017;
  assign new_n7019 = ~new_n7000 & ~new_n7018;
  assign new_n7020 = ~new_n6999 & ~new_n7019;
  assign new_n7021 = ~new_n6991 & ~new_n6994;
  assign new_n7022 = n3311 & n9906;
  assign new_n7023 = n5962 & n9041;
  assign new_n7024 = n1392 & n5801;
  assign new_n7025 = ~new_n7023 & new_n7024;
  assign new_n7026 = new_n7023 & ~new_n7024;
  assign new_n7027 = ~new_n7025 & ~new_n7026;
  assign new_n7028 = new_n7022 & new_n7027;
  assign new_n7029 = ~new_n7022 & ~new_n7027;
  assign new_n7030 = ~new_n7028 & ~new_n7029;
  assign new_n7031 = n6409 & n11058;
  assign new_n7032 = n1007 & n5470;
  assign new_n7033 = n8859 & n13201;
  assign new_n7034_1 = ~new_n7032 & ~new_n7033;
  assign new_n7035 = new_n7032 & new_n7033;
  assign new_n7036 = ~new_n7034_1 & ~new_n7035;
  assign new_n7037 = n3669 & n5969;
  assign new_n7038 = n1364 & n2498;
  assign new_n7039 = new_n7037 & ~new_n7038;
  assign new_n7040 = ~new_n7037 & new_n7038;
  assign new_n7041 = ~new_n7039 & ~new_n7040;
  assign new_n7042 = ~new_n7036 & ~new_n7041;
  assign new_n7043 = new_n7036 & new_n7041;
  assign new_n7044 = ~new_n7042 & ~new_n7043;
  assign new_n7045 = ~new_n7031 & new_n7044;
  assign new_n7046 = new_n7031 & ~new_n7044;
  assign new_n7047 = ~new_n7045 & ~new_n7046;
  assign new_n7048 = ~new_n7030 & new_n7047;
  assign new_n7049 = new_n7030 & ~new_n7047;
  assign new_n7050 = ~new_n7048 & ~new_n7049;
  assign new_n7051 = new_n7021 & new_n7050;
  assign new_n7052 = ~new_n7021 & ~new_n7050;
  assign new_n7053 = ~new_n7051 & ~new_n7052;
  assign new_n7054 = ~new_n6727 & new_n6744;
  assign new_n7055 = new_n6722 & ~new_n7054;
  assign new_n7056 = ~new_n6722 & new_n7054;
  assign new_n7057 = ~new_n7055 & ~new_n7056;
  assign new_n7058 = ~new_n6726 & new_n7057;
  assign new_n7059 = ~new_n6953 & new_n6987;
  assign new_n7060 = ~new_n6951 & ~new_n7059;
  assign new_n7061_1 = n8468 & n10560;
  assign new_n7062 = n6818 & n10908;
  assign new_n7063 = n1084 & n5801;
  assign new_n7064 = ~new_n7062 & ~new_n7063;
  assign new_n7065 = new_n7062 & new_n7063;
  assign new_n7066 = ~new_n7064 & ~new_n7065;
  assign new_n7067 = new_n7061_1 & ~new_n7066;
  assign new_n7068 = ~new_n7061_1 & new_n7066;
  assign new_n7069 = ~new_n7067 & ~new_n7068;
  assign new_n7070 = n9906 & n12003;
  assign new_n7071 = n3311 & n5962;
  assign new_n7072 = n6085 & n8139;
  assign new_n7073 = ~new_n7071 & ~new_n7072;
  assign new_n7074 = new_n7071 & new_n7072;
  assign new_n7075 = ~new_n7073 & ~new_n7074;
  assign new_n7076 = ~new_n7070 & ~new_n7075;
  assign new_n7077 = n9906 & n10560;
  assign new_n7078 = n6085 & n12003;
  assign new_n7079 = ~new_n7077 & ~new_n7078;
  assign new_n7080 = n5962 & n8139;
  assign new_n7081 = new_n7077 & new_n7078;
  assign new_n7082 = ~new_n7080 & ~new_n7081;
  assign new_n7083 = ~new_n7079 & ~new_n7082;
  assign new_n7084 = new_n7070 & new_n7075;
  assign new_n7085 = ~new_n7083 & ~new_n7084;
  assign new_n7086 = ~new_n7076 & ~new_n7085;
  assign new_n7087 = new_n7069 & ~new_n7086;
  assign new_n7088 = ~new_n7069 & new_n7086;
  assign new_n7089 = n11109 & n12003;
  assign new_n7090 = new_n7074 & new_n7089;
  assign new_n7091 = ~new_n7074 & ~new_n7089;
  assign new_n7092 = ~new_n7090 & ~new_n7091;
  assign new_n7093 = n5962 & ~n10866;
  assign new_n7094 = n3311 & n6085;
  assign new_n7095 = n8139 & n9906;
  assign new_n7096 = ~new_n7094 & ~new_n7095;
  assign new_n7097 = new_n7094 & new_n7095;
  assign new_n7098 = ~new_n7096 & ~new_n7097;
  assign new_n7099 = new_n7093 & ~new_n7098;
  assign new_n7100 = ~new_n7093 & new_n7098;
  assign new_n7101 = ~new_n7099 & ~new_n7100;
  assign new_n7102 = new_n7092 & new_n7101;
  assign new_n7103 = ~new_n7092 & ~new_n7101;
  assign new_n7104 = ~new_n7102 & ~new_n7103;
  assign new_n7105 = ~new_n7088 & new_n7104;
  assign new_n7106 = ~new_n7087 & ~new_n7105;
  assign new_n7107 = ~new_n7091 & ~new_n7101;
  assign new_n7108 = ~new_n7090 & ~new_n7107;
  assign new_n7109 = n8139 & n11109;
  assign new_n7110 = n8468 & n12003;
  assign new_n7111_1 = ~new_n7109 & ~new_n7110;
  assign new_n7112 = new_n7109 & new_n7110;
  assign new_n7113_1 = ~new_n7111_1 & ~new_n7112;
  assign new_n7114 = n1084 & n10908;
  assign new_n7115 = n6818 & n10560;
  assign new_n7116 = new_n7114 & ~new_n7115;
  assign new_n7117 = ~new_n7114 & new_n7115;
  assign new_n7118 = ~new_n7116 & ~new_n7117;
  assign new_n7119 = ~new_n7113_1 & ~new_n7118;
  assign new_n7120 = new_n7113_1 & new_n7118;
  assign new_n7121 = ~new_n7119 & ~new_n7120;
  assign new_n7122 = new_n7093 & ~new_n7096;
  assign new_n7123 = ~new_n7097 & ~new_n7122;
  assign new_n7124 = new_n7061_1 & ~new_n7064;
  assign new_n7125 = ~new_n7065 & ~new_n7124;
  assign new_n7126 = ~new_n7123 & new_n7125;
  assign new_n7127 = new_n7123 & ~new_n7125;
  assign new_n7128 = ~new_n7126 & ~new_n7127;
  assign new_n7129 = new_n7121 & new_n7128;
  assign new_n7130 = ~new_n7121 & ~new_n7128;
  assign new_n7131 = ~new_n7129 & ~new_n7130;
  assign new_n7132_1 = new_n7108 & ~new_n7131;
  assign new_n7133 = ~new_n7108 & new_n7131;
  assign new_n7134 = ~new_n7132_1 & ~new_n7133;
  assign new_n7135 = ~new_n7106 & ~new_n7134;
  assign new_n7136 = new_n7106 & new_n7134;
  assign new_n7137 = ~new_n7135 & ~new_n7136;
  assign new_n7138 = new_n7060 & new_n7137;
  assign new_n7139 = ~new_n7060 & ~new_n7137;
  assign new_n7140 = ~new_n7138 & ~new_n7139;
  assign new_n7141 = ~new_n7058 & new_n7140;
  assign new_n7142 = new_n7058 & ~new_n7140;
  assign new_n7143 = ~new_n7141 & ~new_n7142;
  assign new_n7144 = ~new_n7053 & new_n7143;
  assign new_n7145 = new_n7053 & ~new_n7143;
  assign new_n7146 = ~new_n7144 & ~new_n7145;
  assign new_n7147 = ~new_n7020 & ~new_n7146;
  assign new_n7148 = new_n7020 & new_n7146;
  assign new_n7149 = ~new_n7147 & ~new_n7148;
  assign new_n7150 = n6085 & ~n10866;
  assign new_n7151 = n5801 & n8468;
  assign new_n7152 = n10908 & n11109;
  assign new_n7153 = new_n5324 & ~new_n5327;
  assign new_n7154 = ~new_n5328 & ~new_n7153;
  assign new_n7155 = ~new_n7152 & new_n7154;
  assign new_n7156 = new_n7152 & ~new_n7154;
  assign new_n7157 = ~new_n7155 & ~new_n7156;
  assign new_n7158 = ~new_n7079 & ~new_n7081;
  assign new_n7159 = new_n7080 & ~new_n7158;
  assign new_n7160 = ~new_n7080 & new_n7158;
  assign new_n7161_1 = ~new_n7159 & ~new_n7160;
  assign new_n7162 = ~new_n7157 & new_n7161_1;
  assign new_n7163 = new_n7157 & ~new_n7161_1;
  assign new_n7164 = ~new_n7162 & ~new_n7163;
  assign new_n7165 = ~new_n7151 & ~new_n7164;
  assign new_n7166 = new_n7151 & new_n7164;
  assign new_n7167 = ~new_n5322 & new_n5332;
  assign new_n7168 = ~new_n5321 & ~new_n7167;
  assign new_n7169 = ~new_n7166 & ~new_n7168;
  assign new_n7170 = ~new_n7165 & ~new_n7169;
  assign new_n7171 = n10560 & n11109;
  assign new_n7172 = n8468 & n10908;
  assign new_n7173 = ~new_n7171 & ~new_n7172;
  assign new_n7174 = new_n7171 & new_n7172;
  assign new_n7175 = ~new_n7173 & ~new_n7174;
  assign new_n7176 = ~new_n7076 & ~new_n7084;
  assign new_n7177 = ~new_n7083 & ~new_n7176;
  assign new_n7178 = new_n7083 & new_n7176;
  assign new_n7179 = ~new_n7177 & ~new_n7178;
  assign new_n7180 = ~new_n7175 & ~new_n7179;
  assign new_n7181 = new_n7175 & new_n7179;
  assign new_n7182 = ~new_n7180 & ~new_n7181;
  assign new_n7183 = ~new_n7156 & new_n7161_1;
  assign new_n7184 = ~new_n7155 & ~new_n7183;
  assign new_n7185 = ~new_n7182 & ~new_n7184;
  assign new_n7186 = new_n7182 & new_n7184;
  assign new_n7187 = ~new_n7185 & ~new_n7186;
  assign new_n7188 = new_n7170 & new_n7187;
  assign new_n7189 = ~new_n7180 & new_n7184;
  assign new_n7190 = ~new_n7174 & ~new_n7189;
  assign new_n7191 = ~new_n7181 & new_n7190;
  assign new_n7192 = new_n7174 & new_n7189;
  assign new_n7193 = ~new_n7191 & ~new_n7192;
  assign new_n7194 = ~new_n7087 & ~new_n7088;
  assign new_n7195 = new_n7104 & new_n7194;
  assign new_n7196 = ~new_n7104 & ~new_n7194;
  assign new_n7197 = ~new_n7195 & ~new_n7196;
  assign new_n7198 = new_n7193 & ~new_n7197;
  assign new_n7199 = ~new_n7193 & new_n7197;
  assign new_n7200 = ~new_n7198 & ~new_n7199;
  assign new_n7201 = new_n7188 & new_n7200;
  assign new_n7202 = n5801 & n6818;
  assign new_n7203 = ~new_n7170 & ~new_n7187;
  assign new_n7204 = ~new_n7188 & ~new_n7203;
  assign new_n7205 = new_n7202 & new_n7204;
  assign new_n7206 = ~new_n7165 & ~new_n7166;
  assign new_n7207 = new_n7168 & ~new_n7206;
  assign new_n7208 = ~new_n7168 & new_n7206;
  assign new_n7209 = ~new_n7207 & ~new_n7208;
  assign new_n7210 = new_n5337 & ~new_n7209;
  assign new_n7211 = ~new_n7202 & ~new_n7204;
  assign new_n7212 = ~new_n7205 & ~new_n7211;
  assign new_n7213 = new_n7210 & new_n7212;
  assign new_n7214 = ~new_n7205 & ~new_n7213;
  assign new_n7215 = ~new_n7188 & ~new_n7200;
  assign new_n7216 = ~new_n7201 & ~new_n7215;
  assign new_n7217 = ~new_n7214 & new_n7216;
  assign new_n7218 = ~new_n7201 & ~new_n7217;
  assign new_n7219 = ~new_n6839 & new_n6856;
  assign new_n7220 = ~new_n6838 & ~new_n7219;
  assign new_n7221 = new_n6841 & ~new_n6844;
  assign new_n7222 = ~new_n6845 & ~new_n7221;
  assign new_n7223 = n2771 & n3409;
  assign new_n7224 = n1302 & n8308;
  assign new_n7225 = new_n7223 & new_n7224;
  assign new_n7226 = ~new_n7223 & ~new_n7224;
  assign new_n7227 = ~new_n7225 & ~new_n7226;
  assign new_n7228 = new_n7222 & ~new_n7227;
  assign new_n7229 = ~new_n7222 & new_n7227;
  assign new_n7230 = ~new_n7228 & ~new_n7229;
  assign new_n7231 = n499 & n5568;
  assign new_n7232 = n6168 & n10594;
  assign new_n7233 = n5214 & n7113;
  assign new_n7234 = ~new_n7232 & new_n7233;
  assign new_n7235 = new_n7232 & ~new_n7233;
  assign new_n7236 = ~new_n7234 & ~new_n7235;
  assign new_n7237 = new_n7231 & new_n7236;
  assign new_n7238 = ~new_n7231 & ~new_n7236;
  assign new_n7239 = ~new_n7237 & ~new_n7238;
  assign new_n7240 = new_n6849 & ~new_n6851;
  assign new_n7241_1 = ~new_n6852 & ~new_n7240;
  assign new_n7242 = new_n7239 & new_n7241_1;
  assign new_n7243 = ~new_n7239 & ~new_n7241_1;
  assign new_n7244 = ~new_n7242 & ~new_n7243;
  assign new_n7245 = new_n7230 & ~new_n7244;
  assign new_n7246 = ~new_n7230 & new_n7244;
  assign new_n7247 = ~new_n7245 & ~new_n7246;
  assign new_n7248 = ~new_n7220 & new_n7247;
  assign new_n7249 = new_n7220 & ~new_n7247;
  assign new_n7250 = ~new_n7248 & ~new_n7249;
  assign new_n7251 = ~new_n7191 & ~new_n7197;
  assign new_n7252 = ~new_n7192 & ~new_n7251;
  assign new_n7253 = new_n6827 & ~new_n6830;
  assign new_n7254 = ~new_n6831 & ~new_n7253;
  assign new_n7255 = new_n7252 & new_n7254;
  assign new_n7256 = ~new_n7252 & ~new_n7254;
  assign new_n7257 = ~new_n7255 & ~new_n7256;
  assign new_n7258 = new_n7250 & new_n7257;
  assign new_n7259 = ~new_n7250 & ~new_n7257;
  assign new_n7260 = ~new_n7258 & ~new_n7259;
  assign new_n7261 = ~new_n7218 & ~new_n7260;
  assign new_n7262 = new_n7218 & new_n7260;
  assign new_n7263 = ~new_n7261 & ~new_n7262;
  assign new_n7264 = new_n7150 & ~new_n7263;
  assign new_n7265 = ~new_n7150 & new_n7263;
  assign new_n7266 = ~new_n7264 & ~new_n7265;
  assign new_n7267 = ~new_n7149 & new_n7266;
  assign new_n7268 = new_n7149 & ~new_n7266;
  assign new_n7269 = ~new_n7267 & ~new_n7268;
  assign new_n7270 = new_n7214 & ~new_n7216;
  assign new_n7271 = ~new_n7217 & ~new_n7270;
  assign new_n7272 = ~new_n6999 & ~new_n7000;
  assign new_n7273 = ~new_n7018 & ~new_n7272;
  assign new_n7274 = new_n7018 & new_n7272;
  assign new_n7275 = ~new_n7273 & ~new_n7274;
  assign new_n7276 = ~new_n7271 & new_n7275;
  assign new_n7277 = new_n7271 & ~new_n7275;
  assign new_n7278 = ~new_n7210 & ~new_n7212;
  assign new_n7279 = ~new_n7213 & ~new_n7278;
  assign new_n7280 = ~new_n7005 & ~new_n7006;
  assign new_n7281 = new_n7016 & ~new_n7280;
  assign new_n7282 = ~new_n7016 & new_n7280;
  assign new_n7283 = ~new_n7281 & ~new_n7282;
  assign new_n7284 = ~new_n7279 & ~new_n7283;
  assign new_n7285 = new_n7279 & new_n7283;
  assign new_n7286 = ~new_n5337 & new_n7209;
  assign new_n7287 = ~new_n7210 & ~new_n7286;
  assign new_n7288 = ~new_n7011 & ~new_n7012;
  assign new_n7289 = new_n7014 & ~new_n7288;
  assign new_n7290 = ~new_n7014 & new_n7288;
  assign new_n7291 = ~new_n7289 & ~new_n7290;
  assign new_n7292 = new_n7287 & new_n7291;
  assign new_n7293 = ~new_n7287 & ~new_n7291;
  assign new_n7294 = ~new_n5390 & ~new_n5393;
  assign new_n7295 = ~new_n5389 & ~new_n7294;
  assign new_n7296 = ~new_n7293 & ~new_n7295;
  assign new_n7297 = ~new_n7292 & ~new_n7296;
  assign new_n7298 = ~new_n7285 & new_n7297;
  assign new_n7299 = ~new_n7284 & ~new_n7298;
  assign new_n7300 = ~new_n7277 & ~new_n7299;
  assign new_n7301 = ~new_n7276 & ~new_n7300;
  assign new_n7302 = ~new_n6825 & ~new_n6859;
  assign new_n7303 = ~new_n6823 & ~new_n7302;
  assign new_n7304 = ~new_n6733 & ~new_n6737;
  assign new_n7305 = ~new_n6736 & ~new_n7304;
  assign new_n7306 = n3006 & n11111;
  assign new_n7307 = n7061 & n10451;
  assign new_n7308 = n9093 & n11411;
  assign new_n7309 = ~new_n7307 & new_n7308;
  assign new_n7310 = new_n7307 & ~new_n7308;
  assign new_n7311 = ~new_n7309 & ~new_n7310;
  assign new_n7312 = new_n7306 & ~new_n7311;
  assign new_n7313 = ~new_n7306 & new_n7311;
  assign new_n7314 = ~new_n7312 & ~new_n7313;
  assign new_n7315 = ~new_n7305 & new_n7314;
  assign new_n7316 = new_n7305 & ~new_n7314;
  assign new_n7317 = ~new_n7315 & ~new_n7316;
  assign new_n7318 = new_n7303 & new_n7317;
  assign new_n7319 = ~new_n7303 & ~new_n7317;
  assign new_n7320 = ~new_n7318 & ~new_n7319;
  assign new_n7321 = new_n7301 & ~new_n7320;
  assign new_n7322 = ~new_n7301 & new_n7320;
  assign new_n7323 = ~new_n7321 & ~new_n7322;
  assign new_n7324 = ~new_n7269 & ~new_n7323;
  assign new_n7325 = new_n7269 & new_n7323;
  assign new_n7326 = ~new_n7324 & ~new_n7325;
  assign new_n7327 = ~new_n6883 & new_n7326;
  assign new_n7328 = new_n6883 & ~new_n7326;
  assign new_n7329 = ~new_n7327 & ~new_n7328;
  assign new_n7330 = new_n6876 & ~new_n6878;
  assign new_n7331 = ~new_n6879 & ~new_n7330;
  assign new_n7332 = ~new_n7276 & ~new_n7277;
  assign new_n7333 = ~new_n7299 & ~new_n7332;
  assign new_n7334 = new_n7299 & new_n7332;
  assign new_n7335 = ~new_n7333 & ~new_n7334;
  assign new_n7336 = new_n7331 & new_n7335;
  assign new_n7337 = ~new_n7331 & ~new_n7335;
  assign new_n7338 = ~new_n6872 & ~new_n6874;
  assign new_n7339 = ~new_n6875 & ~new_n7338;
  assign new_n7340 = ~new_n7284 & ~new_n7285;
  assign new_n7341 = ~new_n7297 & new_n7340;
  assign new_n7342 = new_n7297 & ~new_n7340;
  assign new_n7343 = ~new_n7341 & ~new_n7342;
  assign new_n7344 = new_n7339 & new_n7343;
  assign new_n7345 = ~new_n7339 & ~new_n7343;
  assign new_n7346 = ~new_n5316 & new_n6871;
  assign new_n7347 = ~new_n6872 & ~new_n7346;
  assign new_n7348 = ~new_n7292 & ~new_n7293;
  assign new_n7349 = new_n7295 & ~new_n7348;
  assign new_n7350 = ~new_n7295 & new_n7348;
  assign new_n7351 = ~new_n7349 & ~new_n7350;
  assign new_n7352 = ~new_n7347 & ~new_n7351;
  assign new_n7353 = new_n7347 & new_n7351;
  assign new_n7354 = ~new_n5296 & ~new_n5397;
  assign new_n7355 = ~new_n5398 & ~new_n7354;
  assign new_n7356 = ~new_n7353 & ~new_n7355;
  assign new_n7357 = ~new_n7352 & ~new_n7356;
  assign new_n7358 = ~new_n7345 & new_n7357;
  assign new_n7359 = ~new_n7344 & ~new_n7358;
  assign new_n7360 = ~new_n7337 & ~new_n7359;
  assign new_n7361 = ~new_n7336 & ~new_n7360;
  assign new_n7362 = ~new_n6731 & new_n6741;
  assign new_n7363 = ~new_n6730 & ~new_n7362;
  assign new_n7364 = ~new_n6966 & new_n6984;
  assign new_n7365 = ~new_n6967 & ~new_n7364;
  assign new_n7366 = n1198 & n4141;
  assign new_n7367 = new_n6957 & ~new_n6960;
  assign new_n7368 = ~new_n6961 & ~new_n7367;
  assign new_n7369 = ~new_n7366 & ~new_n7368;
  assign new_n7370 = new_n7366 & new_n7368;
  assign new_n7371 = ~new_n7369 & ~new_n7370;
  assign new_n7372 = new_n6973 & ~new_n6976;
  assign new_n7373 = ~new_n6977 & ~new_n7372;
  assign new_n7374_1 = n2057 & n11574;
  assign new_n7375 = n5586 & n9300;
  assign new_n7376 = new_n7374_1 & new_n7375;
  assign new_n7377 = ~new_n7374_1 & ~new_n7375;
  assign new_n7378 = ~new_n7376 & ~new_n7377;
  assign new_n7379 = new_n7373 & ~new_n7378;
  assign new_n7380 = ~new_n7373 & new_n7378;
  assign new_n7381 = ~new_n7379 & ~new_n7380;
  assign new_n7382 = ~new_n7371 & new_n7381;
  assign new_n7383 = new_n7371 & ~new_n7381;
  assign new_n7384 = ~new_n7382 & ~new_n7383;
  assign new_n7385 = new_n7365 & ~new_n7384;
  assign new_n7386 = ~new_n7365 & new_n7384;
  assign new_n7387 = ~new_n7385 & ~new_n7386;
  assign new_n7388 = ~new_n6716 & ~new_n6747;
  assign new_n7389 = ~new_n6717 & ~new_n7388;
  assign new_n7390 = ~new_n6971 & new_n6981;
  assign new_n7391 = ~new_n6970 & ~new_n7390;
  assign new_n7392 = n287 & n5167;
  assign new_n7393 = n7720 & n12605;
  assign new_n7394 = n5671 & n6843;
  assign new_n7395 = ~new_n7393 & new_n7394;
  assign new_n7396 = new_n7393 & ~new_n7394;
  assign new_n7397 = ~new_n7395 & ~new_n7396;
  assign new_n7398 = new_n7392 & new_n7397;
  assign new_n7399 = ~new_n7392 & ~new_n7397;
  assign new_n7400 = ~new_n7398 & ~new_n7399;
  assign new_n7401 = n937 & n12482;
  assign new_n7402 = n9570 & n10642;
  assign new_n7403 = ~new_n7401 & ~new_n7402;
  assign new_n7404 = new_n7401 & new_n7402;
  assign new_n7405 = ~new_n7403 & ~new_n7404;
  assign new_n7406 = n1307 & n11665;
  assign new_n7407 = n2339 & n2777;
  assign new_n7408 = new_n7406 & ~new_n7407;
  assign new_n7409 = ~new_n7406 & new_n7407;
  assign new_n7410 = ~new_n7408 & ~new_n7409;
  assign new_n7411_1 = ~new_n7405 & new_n7410;
  assign new_n7412 = new_n7405 & ~new_n7410;
  assign new_n7413 = ~new_n7411_1 & ~new_n7412;
  assign new_n7414 = new_n7400 & ~new_n7413;
  assign new_n7415 = ~new_n7400 & new_n7413;
  assign new_n7416 = ~new_n7414 & ~new_n7415;
  assign new_n7417 = new_n7391 & ~new_n7416;
  assign new_n7418 = ~new_n7391 & new_n7416;
  assign new_n7419 = ~new_n7417 & ~new_n7418;
  assign new_n7420 = new_n7389 & new_n7419;
  assign new_n7421 = ~new_n7389 & ~new_n7419;
  assign new_n7422 = ~new_n7420 & ~new_n7421;
  assign new_n7423 = ~new_n7387 & new_n7422;
  assign new_n7424 = new_n7387 & ~new_n7422;
  assign new_n7425 = ~new_n7423 & ~new_n7424;
  assign new_n7426 = ~new_n7363 & new_n7425;
  assign new_n7427 = new_n7363 & ~new_n7425;
  assign new_n7428 = ~new_n7426 & ~new_n7427;
  assign new_n7429 = new_n7361 & new_n7428;
  assign new_n7430 = ~new_n7361 & ~new_n7428;
  assign new_n7431 = ~new_n7429 & ~new_n7430;
  assign new_n7432 = new_n7329 & new_n7431;
  assign new_n7433 = ~new_n7329 & ~new_n7431;
  assign n1181 = ~new_n7432 & ~new_n7433;
  assign new_n7435 = ~new_n414 & ~new_n416;
  assign n1401 = ~new_n417 & ~new_n7435;
  assign new_n7437 = ~new_n6046 & ~new_n6047;
  assign new_n7438 = ~new_n6051 & new_n7437;
  assign new_n7439 = new_n6051 & ~new_n7437;
  assign n1487 = new_n7438 | new_n7439;
  assign new_n7441 = n2482 & n9093;
  assign new_n7442 = n10113 & n10451;
  assign new_n7443 = new_n7441 & new_n7442;
  assign new_n7444 = n1757 & n10451;
  assign new_n7445 = n9093 & n10113;
  assign new_n7446 = n2482 & n10594;
  assign new_n7447 = ~new_n7445 & ~new_n7446;
  assign new_n7448 = new_n7445 & new_n7446;
  assign new_n7449 = ~new_n7447 & ~new_n7448;
  assign new_n7450 = new_n7444 & ~new_n7449;
  assign new_n7451 = ~new_n7444 & new_n7449;
  assign new_n7452 = ~new_n7450 & ~new_n7451;
  assign new_n7453 = new_n7443 & ~new_n7452;
  assign new_n7454 = n2482 & n3409;
  assign new_n7455 = new_n7444 & ~new_n7447;
  assign new_n7456 = ~new_n7448 & ~new_n7455;
  assign new_n7457 = ~new_n7454 & new_n7456;
  assign new_n7458 = new_n7454 & ~new_n7456;
  assign new_n7459 = ~new_n7457 & ~new_n7458;
  assign new_n7460 = n10416 & n10451;
  assign new_n7461 = n10113 & n10594;
  assign new_n7462 = n1757 & n9093;
  assign new_n7463 = ~new_n7461 & ~new_n7462;
  assign new_n7464 = new_n7461 & new_n7462;
  assign new_n7465 = ~new_n7463 & ~new_n7464;
  assign new_n7466 = new_n7460 & ~new_n7465;
  assign new_n7467 = ~new_n7460 & new_n7465;
  assign new_n7468 = ~new_n7466 & ~new_n7467;
  assign new_n7469 = ~new_n7459 & new_n7468;
  assign new_n7470 = new_n7459 & ~new_n7468;
  assign new_n7471 = ~new_n7469 & ~new_n7470;
  assign new_n7472 = new_n7453 & new_n7471;
  assign new_n7473 = n2482 & n7113;
  assign new_n7474 = n3409 & n10113;
  assign new_n7475 = new_n7460 & ~new_n7463;
  assign new_n7476 = ~new_n7464 & ~new_n7475;
  assign new_n7477 = ~new_n7474 & new_n7476;
  assign new_n7478 = new_n7474 & ~new_n7476;
  assign new_n7479 = ~new_n7477 & ~new_n7478;
  assign new_n7480 = n10451 & n11030;
  assign new_n7481 = n1757 & n10594;
  assign new_n7482 = n9093 & n10416;
  assign new_n7483 = ~new_n7481 & ~new_n7482;
  assign new_n7484 = new_n7481 & new_n7482;
  assign new_n7485 = ~new_n7483 & ~new_n7484;
  assign new_n7486 = new_n7480 & ~new_n7485;
  assign new_n7487 = ~new_n7480 & new_n7485;
  assign new_n7488 = ~new_n7486 & ~new_n7487;
  assign new_n7489 = ~new_n7479 & new_n7488;
  assign new_n7490 = new_n7479 & ~new_n7488;
  assign new_n7491 = ~new_n7489 & ~new_n7490;
  assign new_n7492 = ~new_n7473 & ~new_n7491;
  assign new_n7493 = new_n7473 & new_n7491;
  assign new_n7494 = ~new_n7492 & ~new_n7493;
  assign new_n7495 = ~new_n7457 & ~new_n7468;
  assign new_n7496 = ~new_n7458 & ~new_n7495;
  assign new_n7497 = ~new_n7494 & new_n7496;
  assign new_n7498 = new_n7494 & ~new_n7496;
  assign new_n7499 = ~new_n7497 & ~new_n7498;
  assign new_n7500 = new_n7472 & new_n7499;
  assign new_n7501 = n1302 & n2482;
  assign new_n7502 = ~new_n7493 & new_n7496;
  assign new_n7503 = ~new_n7492 & ~new_n7502;
  assign new_n7504 = n7113 & n10113;
  assign new_n7505 = n1757 & n3409;
  assign new_n7506 = ~new_n7504 & ~new_n7505;
  assign new_n7507 = new_n7504 & new_n7505;
  assign new_n7508 = ~new_n7506 & ~new_n7507;
  assign new_n7509 = n10416 & n10594;
  assign new_n7510 = n9093 & n11030;
  assign new_n7511 = n10451 & n11488;
  assign new_n7512 = ~new_n7510 & ~new_n7511;
  assign new_n7513 = new_n7510 & new_n7511;
  assign new_n7514 = ~new_n7512 & ~new_n7513;
  assign new_n7515 = ~new_n7509 & ~new_n7514;
  assign new_n7516 = new_n7509 & new_n7514;
  assign new_n7517 = ~new_n7515 & ~new_n7516;
  assign new_n7518 = new_n7480 & ~new_n7483;
  assign new_n7519 = ~new_n7484 & ~new_n7518;
  assign new_n7520 = ~new_n7517 & ~new_n7519;
  assign new_n7521 = new_n7517 & new_n7519;
  assign new_n7522 = ~new_n7520 & ~new_n7521;
  assign new_n7523 = ~new_n7508 & new_n7522;
  assign new_n7524 = new_n7508 & ~new_n7522;
  assign new_n7525 = ~new_n7523 & ~new_n7524;
  assign new_n7526 = ~new_n7478 & new_n7488;
  assign new_n7527 = ~new_n7477 & ~new_n7526;
  assign new_n7528 = ~new_n7525 & ~new_n7527;
  assign new_n7529_1 = new_n7525 & new_n7527;
  assign new_n7530 = ~new_n7528 & ~new_n7529_1;
  assign new_n7531 = new_n7503 & new_n7530;
  assign new_n7532 = ~new_n7503 & ~new_n7530;
  assign new_n7533 = ~new_n7531 & ~new_n7532;
  assign new_n7534 = new_n7501 & new_n7533;
  assign new_n7535 = ~new_n7501 & ~new_n7533;
  assign new_n7536 = ~new_n7534 & ~new_n7535;
  assign new_n7537 = new_n7500 & new_n7536;
  assign new_n7538 = ~new_n7500 & ~new_n7536;
  assign new_n7539 = ~new_n7537 & ~new_n7538;
  assign new_n7540 = ~new_n7472 & ~new_n7499;
  assign new_n7541 = ~new_n7500 & ~new_n7540;
  assign new_n7542 = n6085 & n8228;
  assign new_n7543 = n5962 & n11236;
  assign new_n7544 = new_n7542 & new_n7543;
  assign new_n7545 = n4382 & n5962;
  assign new_n7546 = n6085 & n11236;
  assign new_n7547 = n8228 & n9906;
  assign new_n7548 = ~new_n7546 & ~new_n7547;
  assign new_n7549 = new_n7546 & new_n7547;
  assign new_n7550 = ~new_n7548 & ~new_n7549;
  assign new_n7551 = new_n7545 & ~new_n7550;
  assign new_n7552 = ~new_n7545 & new_n7550;
  assign new_n7553_1 = ~new_n7551 & ~new_n7552;
  assign new_n7554 = new_n7544 & ~new_n7553_1;
  assign new_n7555 = n8228 & n11109;
  assign new_n7556 = new_n7545 & ~new_n7548;
  assign new_n7557 = ~new_n7549 & ~new_n7556;
  assign new_n7558 = ~new_n7555 & new_n7557;
  assign new_n7559 = new_n7555 & ~new_n7557;
  assign new_n7560 = ~new_n7558 & ~new_n7559;
  assign new_n7561 = n3130 & n5962;
  assign new_n7562 = n9906 & n11236;
  assign new_n7563 = n4382 & n6085;
  assign new_n7564 = ~new_n7562 & ~new_n7563;
  assign new_n7565 = new_n7562 & new_n7563;
  assign new_n7566 = ~new_n7564 & ~new_n7565;
  assign new_n7567 = new_n7561 & ~new_n7566;
  assign new_n7568 = ~new_n7561 & new_n7566;
  assign new_n7569 = ~new_n7567 & ~new_n7568;
  assign new_n7570 = ~new_n7560 & new_n7569;
  assign new_n7571 = new_n7560 & ~new_n7569;
  assign new_n7572 = ~new_n7570 & ~new_n7571;
  assign new_n7573 = new_n7554 & new_n7572;
  assign new_n7574 = n8228 & n8468;
  assign new_n7575 = n11109 & n11236;
  assign new_n7576 = new_n7561 & ~new_n7564;
  assign new_n7577 = ~new_n7565 & ~new_n7576;
  assign new_n7578 = ~new_n7575 & new_n7577;
  assign new_n7579 = new_n7575 & ~new_n7577;
  assign new_n7580 = ~new_n7578 & ~new_n7579;
  assign new_n7581 = n5962 & n9732;
  assign new_n7582_1 = n4382 & n9906;
  assign new_n7583 = n3130 & n6085;
  assign new_n7584 = ~new_n7582_1 & ~new_n7583;
  assign new_n7585 = new_n7582_1 & new_n7583;
  assign new_n7586 = ~new_n7584 & ~new_n7585;
  assign new_n7587 = new_n7581 & ~new_n7586;
  assign new_n7588 = ~new_n7581 & new_n7586;
  assign new_n7589 = ~new_n7587 & ~new_n7588;
  assign new_n7590 = ~new_n7580 & new_n7589;
  assign new_n7591 = new_n7580 & ~new_n7589;
  assign new_n7592 = ~new_n7590 & ~new_n7591;
  assign new_n7593 = ~new_n7574 & ~new_n7592;
  assign new_n7594 = new_n7574 & new_n7592;
  assign new_n7595 = ~new_n7593 & ~new_n7594;
  assign new_n7596 = ~new_n7559 & new_n7569;
  assign new_n7597 = ~new_n7558 & ~new_n7596;
  assign new_n7598 = ~new_n7595 & ~new_n7597;
  assign new_n7599 = new_n7595 & new_n7597;
  assign new_n7600 = ~new_n7598 & ~new_n7599;
  assign new_n7601 = ~new_n7573 & ~new_n7600;
  assign new_n7602 = new_n7573 & new_n7600;
  assign new_n7603 = ~new_n7601 & ~new_n7602;
  assign new_n7604 = n7720 & n8940;
  assign new_n7605 = n287 & n4964;
  assign new_n7606 = new_n7604 & new_n7605;
  assign new_n7607 = n287 & n5684;
  assign new_n7608 = n4964 & n7720;
  assign new_n7609 = n8940 & n12482;
  assign new_n7610 = ~new_n7608 & ~new_n7609;
  assign new_n7611 = new_n7608 & new_n7609;
  assign new_n7612 = ~new_n7610 & ~new_n7611;
  assign new_n7613 = new_n7607 & ~new_n7612;
  assign new_n7614 = ~new_n7607 & new_n7612;
  assign new_n7615 = ~new_n7613 & ~new_n7614;
  assign new_n7616 = new_n7606 & ~new_n7615;
  assign new_n7617 = n8940 & n9570;
  assign new_n7618 = new_n7607 & ~new_n7610;
  assign new_n7619 = ~new_n7611 & ~new_n7618;
  assign new_n7620 = ~new_n7617 & new_n7619;
  assign new_n7621 = new_n7617 & ~new_n7619;
  assign new_n7622 = ~new_n7620 & ~new_n7621;
  assign new_n7623 = n287 & n10522;
  assign new_n7624 = n4964 & n12482;
  assign new_n7625 = n5684 & n7720;
  assign new_n7626 = ~new_n7624 & ~new_n7625;
  assign new_n7627 = new_n7624 & new_n7625;
  assign new_n7628 = ~new_n7626 & ~new_n7627;
  assign new_n7629 = new_n7623 & ~new_n7628;
  assign new_n7630 = ~new_n7623 & new_n7628;
  assign new_n7631 = ~new_n7629 & ~new_n7630;
  assign new_n7632 = ~new_n7622 & new_n7631;
  assign new_n7633 = new_n7622 & ~new_n7631;
  assign new_n7634 = ~new_n7632 & ~new_n7633;
  assign new_n7635 = new_n7616 & new_n7634;
  assign new_n7636 = n2339 & n8940;
  assign new_n7637 = n4964 & n9570;
  assign new_n7638 = new_n7623 & ~new_n7626;
  assign new_n7639 = ~new_n7627 & ~new_n7638;
  assign new_n7640 = ~new_n7637 & new_n7639;
  assign new_n7641 = new_n7637 & ~new_n7639;
  assign new_n7642 = ~new_n7640 & ~new_n7641;
  assign new_n7643 = n287 & n10770;
  assign new_n7644 = n5684 & n12482;
  assign new_n7645 = n7720 & n10522;
  assign new_n7646 = ~new_n7644 & ~new_n7645;
  assign new_n7647 = new_n7644 & new_n7645;
  assign new_n7648 = ~new_n7646 & ~new_n7647;
  assign new_n7649 = new_n7643 & ~new_n7648;
  assign new_n7650 = ~new_n7643 & new_n7648;
  assign new_n7651 = ~new_n7649 & ~new_n7650;
  assign new_n7652 = ~new_n7642 & new_n7651;
  assign new_n7653 = new_n7642 & ~new_n7651;
  assign new_n7654 = ~new_n7652 & ~new_n7653;
  assign new_n7655 = ~new_n7636 & ~new_n7654;
  assign new_n7656 = new_n7636 & new_n7654;
  assign new_n7657 = ~new_n7655 & ~new_n7656;
  assign new_n7658 = ~new_n7620 & ~new_n7631;
  assign new_n7659_1 = ~new_n7621 & ~new_n7658;
  assign new_n7660 = ~new_n7657 & ~new_n7659_1;
  assign new_n7661 = new_n7657 & new_n7659_1;
  assign new_n7662 = ~new_n7660 & ~new_n7661;
  assign new_n7663 = ~new_n7635 & new_n7662;
  assign new_n7664 = new_n7635 & ~new_n7662;
  assign new_n7665 = ~new_n7663 & ~new_n7664;
  assign new_n7666 = n1007 & n9353;
  assign new_n7667 = n6333 & n11058;
  assign new_n7668 = new_n7666 & new_n7667;
  assign new_n7669 = n1912 & n11058;
  assign new_n7670 = n1007 & n6333;
  assign new_n7671 = n5969 & n9353;
  assign new_n7672 = ~new_n7670 & ~new_n7671;
  assign new_n7673 = new_n7670 & new_n7671;
  assign new_n7674 = ~new_n7672 & ~new_n7673;
  assign new_n7675 = new_n7669 & ~new_n7674;
  assign new_n7676 = ~new_n7669 & new_n7674;
  assign new_n7677 = ~new_n7675 & ~new_n7676;
  assign new_n7678 = new_n7668 & ~new_n7677;
  assign new_n7679 = n2498 & n9353;
  assign new_n7680 = new_n7669 & ~new_n7672;
  assign new_n7681 = ~new_n7673 & ~new_n7680;
  assign new_n7682 = ~new_n7679 & new_n7681;
  assign new_n7683 = new_n7679 & ~new_n7681;
  assign new_n7684 = ~new_n7682 & ~new_n7683;
  assign new_n7685 = n11058 & n12750;
  assign new_n7686 = n5969 & n6333;
  assign new_n7687_1 = n1007 & n1912;
  assign new_n7688 = ~new_n7686 & ~new_n7687_1;
  assign new_n7689 = new_n7686 & new_n7687_1;
  assign new_n7690 = ~new_n7688 & ~new_n7689;
  assign new_n7691 = new_n7685 & ~new_n7690;
  assign new_n7692 = ~new_n7685 & new_n7690;
  assign new_n7693 = ~new_n7691 & ~new_n7692;
  assign new_n7694 = ~new_n7684 & new_n7693;
  assign new_n7695 = new_n7684 & ~new_n7693;
  assign new_n7696 = ~new_n7694 & ~new_n7695;
  assign new_n7697 = new_n7678 & new_n7696;
  assign new_n7698 = n1198 & n9353;
  assign new_n7699 = n2498 & n6333;
  assign new_n7700 = new_n7685 & ~new_n7688;
  assign new_n7701 = ~new_n7689 & ~new_n7700;
  assign new_n7702 = ~new_n7699 & new_n7701;
  assign new_n7703 = new_n7699 & ~new_n7701;
  assign new_n7704 = ~new_n7702 & ~new_n7703;
  assign new_n7705 = n9620 & n11058;
  assign new_n7706 = n1912 & n5969;
  assign new_n7707 = n1007 & n12750;
  assign new_n7708 = ~new_n7706 & ~new_n7707;
  assign new_n7709 = new_n7706 & new_n7707;
  assign new_n7710 = ~new_n7708 & ~new_n7709;
  assign new_n7711 = new_n7705 & ~new_n7710;
  assign new_n7712 = ~new_n7705 & new_n7710;
  assign new_n7713 = ~new_n7711 & ~new_n7712;
  assign new_n7714 = ~new_n7704 & new_n7713;
  assign new_n7715_1 = new_n7704 & ~new_n7713;
  assign new_n7716 = ~new_n7714 & ~new_n7715_1;
  assign new_n7717 = ~new_n7698 & ~new_n7716;
  assign new_n7718 = new_n7698 & new_n7716;
  assign new_n7719 = ~new_n7717 & ~new_n7718;
  assign new_n7720_1 = ~new_n7683 & new_n7693;
  assign new_n7721 = ~new_n7682 & ~new_n7720_1;
  assign new_n7722 = ~new_n7719 & ~new_n7721;
  assign new_n7723 = new_n7719 & new_n7721;
  assign new_n7724 = ~new_n7722 & ~new_n7723;
  assign new_n7725 = ~new_n7697 & ~new_n7724;
  assign new_n7726 = new_n7697 & new_n7724;
  assign new_n7727 = ~new_n7725 & ~new_n7726;
  assign new_n7728 = ~new_n7665 & ~new_n7727;
  assign new_n7729_1 = new_n7665 & new_n7727;
  assign new_n7730 = ~new_n7728 & ~new_n7729_1;
  assign new_n7731 = ~new_n7616 & ~new_n7634;
  assign new_n7732 = ~new_n7635 & ~new_n7731;
  assign new_n7733 = ~new_n7678 & ~new_n7696;
  assign new_n7734 = ~new_n7697 & ~new_n7733;
  assign new_n7735 = new_n7732 & new_n7734;
  assign new_n7736 = ~new_n7732 & ~new_n7734;
  assign new_n7737 = ~new_n7606 & new_n7615;
  assign new_n7738 = ~new_n7616 & ~new_n7737;
  assign new_n7739 = ~new_n7668 & new_n7677;
  assign new_n7740 = ~new_n7678 & ~new_n7739;
  assign new_n7741 = new_n7738 & new_n7740;
  assign new_n7742 = ~new_n7738 & ~new_n7740;
  assign new_n7743 = ~new_n7666 & ~new_n7667;
  assign new_n7744 = ~new_n7668 & ~new_n7743;
  assign new_n7745 = new_n3761 & new_n7744;
  assign new_n7746 = ~new_n3761 & ~new_n7744;
  assign new_n7747 = ~new_n7604 & ~new_n7605;
  assign new_n7748 = ~new_n7606 & ~new_n7747;
  assign new_n7749 = ~new_n7746 & new_n7748;
  assign new_n7750 = ~new_n7745 & ~new_n7749;
  assign new_n7751 = ~new_n7742 & ~new_n7750;
  assign new_n7752 = ~new_n7741 & ~new_n7751;
  assign new_n7753 = ~new_n7736 & ~new_n7752;
  assign new_n7754 = ~new_n7735 & ~new_n7753;
  assign new_n7755_1 = ~new_n7730 & new_n7754;
  assign new_n7756 = new_n7730 & ~new_n7754;
  assign new_n7757 = ~new_n7755_1 & ~new_n7756;
  assign new_n7758 = new_n7603 & new_n7757;
  assign new_n7759 = ~new_n7603 & ~new_n7757;
  assign new_n7760 = ~new_n7758 & ~new_n7759;
  assign new_n7761 = ~new_n7554 & ~new_n7572;
  assign new_n7762 = ~new_n7573 & ~new_n7761;
  assign new_n7763 = ~new_n7735 & ~new_n7736;
  assign new_n7764 = new_n7752 & ~new_n7763;
  assign new_n7765 = ~new_n7752 & new_n7763;
  assign new_n7766 = ~new_n7764 & ~new_n7765;
  assign new_n7767 = ~new_n7762 & ~new_n7766;
  assign new_n7768 = new_n7762 & new_n7766;
  assign new_n7769 = ~new_n7544 & new_n7553_1;
  assign new_n7770 = ~new_n7554 & ~new_n7769;
  assign new_n7771 = ~new_n7741 & ~new_n7742;
  assign new_n7772_1 = new_n7750 & ~new_n7771;
  assign new_n7773 = ~new_n7750 & new_n7771;
  assign new_n7774 = ~new_n7772_1 & ~new_n7773;
  assign new_n7775 = ~new_n7770 & ~new_n7774;
  assign new_n7776 = new_n7770 & new_n7774;
  assign new_n7777 = ~new_n7542 & ~new_n7543;
  assign new_n7778 = ~new_n7544 & ~new_n7777;
  assign new_n7779 = ~new_n7745 & ~new_n7746;
  assign new_n7780 = new_n7748 & ~new_n7779;
  assign new_n7781 = ~new_n7748 & new_n7779;
  assign new_n7782 = ~new_n7780 & ~new_n7781;
  assign new_n7783 = ~new_n7778 & new_n7782;
  assign new_n7784 = new_n7778 & ~new_n7782;
  assign new_n7785 = ~new_n3765 & ~new_n7784;
  assign new_n7786 = ~new_n7783 & ~new_n7785;
  assign new_n7787 = ~new_n7776 & ~new_n7786;
  assign new_n7788 = ~new_n7775 & ~new_n7787;
  assign new_n7789 = ~new_n7768 & ~new_n7788;
  assign new_n7790_1 = ~new_n7767 & ~new_n7789;
  assign new_n7791 = ~new_n7760 & new_n7790_1;
  assign new_n7792 = new_n7760 & ~new_n7790_1;
  assign new_n7793 = ~new_n7791 & ~new_n7792;
  assign new_n7794 = ~new_n7541 & new_n7793;
  assign new_n7795 = new_n7541 & ~new_n7793;
  assign new_n7796 = ~new_n7453 & ~new_n7471;
  assign new_n7797 = ~new_n7472 & ~new_n7796;
  assign new_n7798 = ~new_n7767 & ~new_n7768;
  assign new_n7799 = new_n7788 & ~new_n7798;
  assign new_n7800 = ~new_n7788 & new_n7798;
  assign new_n7801 = ~new_n7799 & ~new_n7800;
  assign new_n7802 = new_n7797 & ~new_n7801;
  assign new_n7803 = ~new_n7797 & new_n7801;
  assign new_n7804 = ~new_n7443 & new_n7452;
  assign new_n7805 = ~new_n7453 & ~new_n7804;
  assign new_n7806 = ~new_n7775 & ~new_n7776;
  assign new_n7807 = new_n7786 & ~new_n7806;
  assign new_n7808 = ~new_n7786 & new_n7806;
  assign new_n7809 = ~new_n7807 & ~new_n7808;
  assign new_n7810 = new_n7805 & ~new_n7809;
  assign new_n7811 = ~new_n7805 & new_n7809;
  assign new_n7812_1 = ~new_n7441 & ~new_n7442;
  assign new_n7813 = ~new_n7443 & ~new_n7812_1;
  assign new_n7814 = ~new_n3768 & ~new_n7813;
  assign new_n7815 = new_n3768 & new_n7813;
  assign new_n7816 = ~new_n7783 & ~new_n7784;
  assign new_n7817 = new_n3765 & ~new_n7816;
  assign new_n7818 = ~new_n3765 & new_n7816;
  assign new_n7819 = ~new_n7817 & ~new_n7818;
  assign new_n7820 = ~new_n7815 & new_n7819;
  assign new_n7821 = ~new_n7814 & ~new_n7820;
  assign new_n7822 = ~new_n7811 & new_n7821;
  assign new_n7823 = ~new_n7810 & ~new_n7822;
  assign new_n7824 = ~new_n7803 & ~new_n7823;
  assign new_n7825 = ~new_n7802 & ~new_n7824;
  assign new_n7826 = ~new_n7795 & new_n7825;
  assign new_n7827 = ~new_n7794 & ~new_n7826;
  assign new_n7828 = ~new_n7539 & ~new_n7827;
  assign new_n7829 = new_n7539 & new_n7827;
  assign new_n7830 = ~new_n7828 & ~new_n7829;
  assign new_n7831 = n6818 & n8228;
  assign new_n7832 = n8468 & n11236;
  assign new_n7833 = n4382 & n11109;
  assign new_n7834 = ~new_n7832 & ~new_n7833;
  assign new_n7835 = new_n7832 & new_n7833;
  assign new_n7836 = ~new_n7834 & ~new_n7835;
  assign new_n7837 = n3130 & n9906;
  assign new_n7838 = n6085 & n9732;
  assign new_n7839 = n103 & n5962;
  assign new_n7840 = ~new_n7838 & ~new_n7839;
  assign new_n7841 = new_n7838 & new_n7839;
  assign new_n7842 = ~new_n7840 & ~new_n7841;
  assign new_n7843 = ~new_n7837 & ~new_n7842;
  assign new_n7844 = new_n7837 & new_n7842;
  assign new_n7845 = ~new_n7843 & ~new_n7844;
  assign new_n7846 = new_n7581 & ~new_n7584;
  assign new_n7847 = ~new_n7585 & ~new_n7846;
  assign new_n7848 = ~new_n7845 & ~new_n7847;
  assign new_n7849 = new_n7845 & new_n7847;
  assign new_n7850 = ~new_n7848 & ~new_n7849;
  assign new_n7851 = ~new_n7836 & new_n7850;
  assign new_n7852 = new_n7836 & ~new_n7850;
  assign new_n7853 = ~new_n7851 & ~new_n7852;
  assign new_n7854 = ~new_n7578 & ~new_n7589;
  assign new_n7855 = ~new_n7579 & ~new_n7854;
  assign new_n7856 = ~new_n7853 & new_n7855;
  assign new_n7857 = new_n7853 & ~new_n7855;
  assign new_n7858_1 = ~new_n7856 & ~new_n7857;
  assign new_n7859 = ~new_n7593 & new_n7597;
  assign new_n7860_1 = ~new_n7594 & ~new_n7859;
  assign new_n7861 = new_n7858_1 & ~new_n7860_1;
  assign new_n7862 = ~new_n7858_1 & new_n7860_1;
  assign new_n7863 = ~new_n7861 & ~new_n7862;
  assign new_n7864 = new_n7831 & new_n7863;
  assign new_n7865 = ~new_n7831 & ~new_n7863;
  assign new_n7866 = ~new_n7864 & ~new_n7865;
  assign new_n7867 = ~new_n7602 & ~new_n7866;
  assign new_n7868 = new_n7602 & new_n7866;
  assign new_n7869 = ~new_n7867 & ~new_n7868;
  assign new_n7870 = ~new_n7758 & ~new_n7790_1;
  assign new_n7871 = ~new_n7759 & ~new_n7870;
  assign new_n7872 = ~new_n7869 & ~new_n7871;
  assign new_n7873 = new_n7869 & new_n7871;
  assign new_n7874 = ~new_n7872 & ~new_n7873;
  assign new_n7875 = n1307 & n8940;
  assign new_n7876 = n5684 & n9570;
  assign new_n7877 = n2339 & n4964;
  assign new_n7878 = ~new_n7876 & ~new_n7877;
  assign new_n7879 = new_n7876 & new_n7877;
  assign new_n7880 = ~new_n7878 & ~new_n7879;
  assign new_n7881 = n10522 & n12482;
  assign new_n7882 = n7720 & n10770;
  assign new_n7883 = n287 & new_n7882;
  assign new_n7884 = ~new_n7643 & ~new_n7882;
  assign new_n7885 = ~new_n7883 & ~new_n7884;
  assign new_n7886 = ~new_n7881 & ~new_n7885;
  assign new_n7887 = new_n7881 & new_n7885;
  assign new_n7888 = ~new_n7886 & ~new_n7887;
  assign new_n7889 = new_n7643 & ~new_n7646;
  assign new_n7890 = ~new_n7647 & ~new_n7889;
  assign new_n7891 = ~new_n7888 & new_n7890;
  assign new_n7892 = new_n7888 & ~new_n7890;
  assign new_n7893 = ~new_n7891 & ~new_n7892;
  assign new_n7894 = ~new_n7880 & ~new_n7893;
  assign new_n7895 = new_n7880 & new_n7893;
  assign new_n7896 = ~new_n7894 & ~new_n7895;
  assign new_n7897 = ~new_n7641 & new_n7651;
  assign new_n7898 = ~new_n7640 & ~new_n7897;
  assign new_n7899 = ~new_n7896 & ~new_n7898;
  assign new_n7900 = new_n7896 & new_n7898;
  assign new_n7901 = ~new_n7899 & ~new_n7900;
  assign new_n7902 = ~new_n7655 & ~new_n7659_1;
  assign new_n7903 = ~new_n7656 & ~new_n7902;
  assign new_n7904 = new_n7901 & ~new_n7903;
  assign new_n7905 = ~new_n7901 & new_n7903;
  assign new_n7906 = ~new_n7904 & ~new_n7905;
  assign new_n7907 = new_n7875 & new_n7906;
  assign new_n7908 = ~new_n7875 & ~new_n7906;
  assign new_n7909 = ~new_n7907 & ~new_n7908;
  assign new_n7910 = new_n7664 & new_n7909;
  assign new_n7911 = ~new_n7664 & ~new_n7909;
  assign new_n7912 = ~new_n7910 & ~new_n7911;
  assign new_n7913 = n9300 & n9353;
  assign new_n7914 = n1198 & n6333;
  assign new_n7915 = n1912 & n2498;
  assign new_n7916 = ~new_n7914 & ~new_n7915;
  assign new_n7917 = new_n7914 & new_n7915;
  assign new_n7918 = ~new_n7916 & ~new_n7917;
  assign new_n7919 = n5969 & n12750;
  assign new_n7920 = n1007 & n9620;
  assign new_n7921 = n761 & n11058;
  assign new_n7922 = ~new_n7920 & ~new_n7921;
  assign new_n7923 = new_n7920 & new_n7921;
  assign new_n7924 = ~new_n7922 & ~new_n7923;
  assign new_n7925 = new_n7919 & new_n7924;
  assign new_n7926 = ~new_n7919 & ~new_n7924;
  assign new_n7927 = ~new_n7925 & ~new_n7926;
  assign new_n7928 = new_n7705 & ~new_n7708;
  assign new_n7929 = ~new_n7709 & ~new_n7928;
  assign new_n7930 = ~new_n7927 & new_n7929;
  assign new_n7931 = new_n7927 & ~new_n7929;
  assign new_n7932 = ~new_n7930 & ~new_n7931;
  assign new_n7933 = ~new_n7918 & ~new_n7932;
  assign new_n7934 = new_n7918 & new_n7932;
  assign new_n7935 = ~new_n7933 & ~new_n7934;
  assign new_n7936 = ~new_n7702 & ~new_n7713;
  assign new_n7937 = ~new_n7703 & ~new_n7936;
  assign new_n7938 = ~new_n7935 & ~new_n7937;
  assign new_n7939 = new_n7935 & new_n7937;
  assign new_n7940 = ~new_n7938 & ~new_n7939;
  assign new_n7941 = ~new_n7717 & new_n7721;
  assign new_n7942 = ~new_n7718 & ~new_n7941;
  assign new_n7943 = ~new_n7940 & ~new_n7942;
  assign new_n7944 = new_n7940 & new_n7942;
  assign new_n7945 = ~new_n7943 & ~new_n7944;
  assign new_n7946 = new_n7913 & new_n7945;
  assign new_n7947 = ~new_n7913 & ~new_n7945;
  assign new_n7948 = ~new_n7946 & ~new_n7947;
  assign new_n7949 = new_n7726 & new_n7948;
  assign new_n7950 = ~new_n7726 & ~new_n7948;
  assign new_n7951 = ~new_n7949 & ~new_n7950;
  assign new_n7952 = new_n7912 & new_n7951;
  assign new_n7953 = ~new_n7912 & ~new_n7951;
  assign new_n7954 = ~new_n7952 & ~new_n7953;
  assign new_n7955 = ~new_n7728 & ~new_n7754;
  assign new_n7956 = ~new_n7729_1 & ~new_n7955;
  assign new_n7957 = ~new_n7954 & ~new_n7956;
  assign new_n7958 = ~new_n7952 & new_n7956;
  assign new_n7959 = ~new_n7953 & new_n7958;
  assign new_n7960 = ~new_n7957 & ~new_n7959;
  assign new_n7961 = ~new_n7874 & new_n7960;
  assign new_n7962 = new_n7874 & ~new_n7960;
  assign new_n7963 = ~new_n7961 & ~new_n7962;
  assign new_n7964 = ~new_n7830 & new_n7963;
  assign new_n7965 = ~new_n7829 & ~new_n7963;
  assign new_n7966 = ~new_n7828 & new_n7965;
  assign n1561 = new_n7964 | new_n7966;
  assign new_n7968_1 = ~new_n7814 & ~new_n7815;
  assign new_n7969 = ~new_n7819 & new_n7968_1;
  assign new_n7970 = new_n7819 & ~new_n7968_1;
  assign n1806 = ~new_n7969 & ~new_n7970;
  assign new_n7972 = ~new_n2641 & ~new_n2642;
  assign new_n7973 = ~new_n2646 & ~new_n7972;
  assign new_n7974_1 = new_n2646 & new_n7972;
  assign n1860 = new_n7973 | new_n7974_1;
  assign new_n7976 = ~new_n6412 & ~new_n6413;
  assign new_n7977 = new_n6415 & ~new_n7976;
  assign new_n7978 = ~new_n6415 & new_n7976;
  assign n1937 = new_n7977 | new_n7978;
  assign new_n7980 = n7772 & n9747;
  assign new_n7981 = n4330 & n7715;
  assign new_n7982 = n2252 & n7529;
  assign new_n7983 = ~new_n7981 & ~new_n7982;
  assign new_n7984 = new_n7981 & new_n7982;
  assign new_n7985 = ~new_n7983 & ~new_n7984;
  assign new_n7986 = n2458 & n7659;
  assign new_n7987 = n8230 & n12289;
  assign new_n7988 = n5729 & n6668;
  assign new_n7989 = ~new_n7987 & ~new_n7988;
  assign new_n7990 = new_n7987 & new_n7988;
  assign new_n7991 = ~new_n7989 & ~new_n7990;
  assign new_n7992 = ~new_n7986 & ~new_n7991;
  assign new_n7993 = new_n7986 & new_n7991;
  assign new_n7994 = ~new_n7992 & ~new_n7993;
  assign new_n7995 = n2458 & n12289;
  assign new_n7996 = n5729 & n8230;
  assign new_n7997 = new_n7995 & new_n7996;
  assign new_n7998 = ~new_n7995 & ~new_n7996;
  assign new_n7999 = n7659 & n7715;
  assign new_n8000 = ~new_n7998 & new_n7999;
  assign new_n8001 = ~new_n7997 & ~new_n8000;
  assign new_n8002 = ~new_n7994 & ~new_n8001;
  assign new_n8003 = new_n7994 & new_n8001;
  assign new_n8004 = ~new_n8002 & ~new_n8003;
  assign new_n8005 = ~new_n7985 & new_n8004;
  assign new_n8006 = new_n7985 & ~new_n8004;
  assign new_n8007 = ~new_n8005 & ~new_n8006;
  assign new_n8008 = n4330 & n7529;
  assign new_n8009 = new_n4125 & new_n7986;
  assign new_n8010 = n2458 & n5729;
  assign new_n8011 = n7529 & n7659;
  assign new_n8012 = ~new_n8010 & ~new_n8011;
  assign new_n8013 = n7715 & n12289;
  assign new_n8014 = ~new_n8012 & new_n8013;
  assign new_n8015 = ~new_n8009 & ~new_n8014;
  assign new_n8016 = ~new_n8008 & new_n8015;
  assign new_n8017 = new_n8008 & ~new_n8015;
  assign new_n8018 = ~new_n7997 & ~new_n7998;
  assign new_n8019 = ~new_n7999 & ~new_n8018;
  assign new_n8020 = new_n7999 & new_n8018;
  assign new_n8021 = ~new_n8019 & ~new_n8020;
  assign new_n8022 = ~new_n8017 & ~new_n8021;
  assign new_n8023 = ~new_n8016 & ~new_n8022;
  assign new_n8024 = ~new_n8007 & new_n8023;
  assign new_n8025 = new_n8007 & ~new_n8023;
  assign new_n8026 = ~new_n8024 & ~new_n8025;
  assign new_n8027 = n2252 & n7772;
  assign new_n8028 = ~new_n8016 & ~new_n8017;
  assign new_n8029 = new_n8021 & ~new_n8028;
  assign new_n8030 = ~new_n8021 & new_n8028;
  assign new_n8031 = ~new_n8029 & ~new_n8030;
  assign new_n8032 = new_n8027 & ~new_n8031;
  assign new_n8033 = ~new_n8027 & new_n8031;
  assign new_n8034 = n4330 & n7772;
  assign new_n8035 = new_n4122_1 & new_n7999;
  assign new_n8036 = n7529 & n12289;
  assign new_n8037 = n5729 & n7715;
  assign new_n8038 = n7659 & n7772;
  assign new_n8039 = ~new_n8037 & ~new_n8038;
  assign new_n8040 = new_n8036 & ~new_n8039;
  assign new_n8041 = ~new_n8035 & ~new_n8040;
  assign new_n8042 = ~new_n8034 & new_n8041;
  assign new_n8043 = new_n8034 & ~new_n8041;
  assign new_n8044 = ~new_n8009 & ~new_n8012;
  assign new_n8045 = ~new_n8013 & ~new_n8044;
  assign new_n8046 = new_n8013 & new_n8044;
  assign new_n8047 = ~new_n8045 & ~new_n8046;
  assign new_n8048 = ~new_n8043 & ~new_n8047;
  assign new_n8049 = ~new_n8042 & ~new_n8048;
  assign new_n8050 = ~new_n8033 & new_n8049;
  assign new_n8051 = ~new_n8032 & ~new_n8050;
  assign new_n8052 = ~new_n8026 & ~new_n8051;
  assign new_n8053 = new_n8026 & new_n8051;
  assign new_n8054 = ~new_n8052 & ~new_n8053;
  assign new_n8055 = new_n7980 & new_n8054;
  assign new_n8056 = ~new_n8035 & ~new_n8039;
  assign new_n8057 = new_n4127 & ~new_n8056;
  assign new_n8058 = ~new_n8042 & ~new_n8043;
  assign new_n8059 = ~new_n8047 & ~new_n8058;
  assign new_n8060 = new_n8047 & new_n8058;
  assign new_n8061 = ~new_n8059 & ~new_n8060;
  assign new_n8062 = new_n8057 & new_n8061;
  assign new_n8063 = ~new_n8032 & ~new_n8033;
  assign new_n8064 = ~new_n8049 & ~new_n8063;
  assign new_n8065 = new_n8049 & new_n8063;
  assign new_n8066 = ~new_n8064 & ~new_n8065;
  assign new_n8067 = new_n8062 & new_n8066;
  assign new_n8068 = ~new_n7980 & ~new_n8054;
  assign new_n8069 = ~new_n8055 & ~new_n8068;
  assign new_n8070 = new_n8067 & new_n8069;
  assign new_n8071 = ~new_n8055 & ~new_n8070;
  assign new_n8072 = n5884 & n7772;
  assign new_n8073 = n2252 & n7715;
  assign new_n8074 = n7529 & n9747;
  assign new_n8075 = ~new_n8073 & ~new_n8074;
  assign new_n8076 = new_n8073 & new_n8074;
  assign new_n8077 = ~new_n8075 & ~new_n8076;
  assign new_n8078 = new_n8072 & ~new_n8077;
  assign new_n8079 = ~new_n8072 & new_n8077;
  assign new_n8080 = ~new_n8078 & ~new_n8079;
  assign new_n8081 = ~new_n7993 & new_n8001;
  assign new_n8082 = ~new_n7992 & ~new_n8081;
  assign new_n8083 = new_n8080 & ~new_n8082;
  assign new_n8084 = ~new_n8080 & new_n8082;
  assign new_n8085 = ~new_n8083 & ~new_n8084;
  assign new_n8086 = n2458 & n4330;
  assign new_n8087 = new_n7990 & new_n8086;
  assign new_n8088 = ~new_n7990 & ~new_n8086;
  assign new_n8089 = ~new_n8087 & ~new_n8088;
  assign new_n8090 = n7659 & n8230;
  assign new_n8091 = n6668 & n12289;
  assign new_n8092 = n5729 & n7812;
  assign new_n8093 = ~new_n8091 & ~new_n8092;
  assign new_n8094 = new_n8091 & new_n8092;
  assign new_n8095 = ~new_n8093 & ~new_n8094;
  assign new_n8096 = new_n8090 & ~new_n8095;
  assign new_n8097 = ~new_n8090 & new_n8095;
  assign new_n8098 = ~new_n8096 & ~new_n8097;
  assign new_n8099 = new_n8089 & new_n8098;
  assign new_n8100 = ~new_n8089 & ~new_n8098;
  assign new_n8101 = ~new_n8099 & ~new_n8100;
  assign new_n8102 = new_n8085 & new_n8101;
  assign new_n8103 = ~new_n8085 & ~new_n8101;
  assign new_n8104 = ~new_n8102 & ~new_n8103;
  assign new_n8105 = ~new_n8005 & new_n8023;
  assign new_n8106 = ~new_n7984 & ~new_n8105;
  assign new_n8107 = ~new_n8006 & new_n8106;
  assign new_n8108 = new_n7984 & new_n8105;
  assign new_n8109 = ~new_n8107 & ~new_n8108;
  assign new_n8110 = ~new_n8104 & new_n8109;
  assign new_n8111 = new_n8104 & ~new_n8109;
  assign new_n8112 = ~new_n8110 & ~new_n8111;
  assign new_n8113 = new_n8052 & new_n8112;
  assign new_n8114 = ~new_n8052 & ~new_n8112;
  assign new_n8115 = ~new_n8113 & ~new_n8114;
  assign new_n8116 = ~new_n8071 & new_n8115;
  assign new_n8117 = new_n8071 & ~new_n8115;
  assign new_n8118 = ~new_n8116 & ~new_n8117;
  assign new_n8119 = n1636 & n2068;
  assign new_n8120 = n5065 & n12348;
  assign new_n8121 = ~new_n8119 & ~new_n8120;
  assign new_n8122 = new_n8119 & new_n8120;
  assign new_n8123 = ~new_n8121 & ~new_n8122;
  assign new_n8124 = n4862 & n11324;
  assign new_n8125 = n5920 & n8183;
  assign new_n8126 = n10142 & n13058;
  assign new_n8127 = ~new_n8125 & ~new_n8126;
  assign new_n8128 = new_n8125 & new_n8126;
  assign new_n8129 = ~new_n8127 & ~new_n8128;
  assign new_n8130 = ~new_n8124 & ~new_n8129;
  assign new_n8131 = new_n8124 & new_n8129;
  assign new_n8132 = ~new_n8130 & ~new_n8131;
  assign new_n8133 = n5920 & n11324;
  assign new_n8134 = n8183 & n13058;
  assign new_n8135 = new_n8133 & new_n8134;
  assign new_n8136 = ~new_n8133 & ~new_n8134;
  assign new_n8137 = n2068 & n4862;
  assign new_n8138 = ~new_n8136 & new_n8137;
  assign new_n8139_1 = ~new_n8135 & ~new_n8138;
  assign new_n8140 = ~new_n8132 & ~new_n8139_1;
  assign new_n8141 = new_n8132 & new_n8139_1;
  assign new_n8142 = ~new_n8140 & ~new_n8141;
  assign new_n8143 = ~new_n8123 & new_n8142;
  assign new_n8144 = new_n8123 & ~new_n8142;
  assign new_n8145 = ~new_n8143 & ~new_n8144;
  assign new_n8146 = n1636 & n12348;
  assign new_n8147 = new_n4132 & new_n8124;
  assign new_n8148 = n11324 & n13058;
  assign new_n8149 = n4862 & n12348;
  assign new_n8150 = ~new_n8148 & ~new_n8149;
  assign new_n8151 = n2068 & n5920;
  assign new_n8152 = ~new_n8150 & new_n8151;
  assign new_n8153 = ~new_n8147 & ~new_n8152;
  assign new_n8154 = ~new_n8146 & new_n8153;
  assign new_n8155 = new_n8146 & ~new_n8153;
  assign new_n8156 = ~new_n8135 & ~new_n8136;
  assign new_n8157 = ~new_n8137 & ~new_n8156;
  assign new_n8158 = new_n8137 & new_n8156;
  assign new_n8159 = ~new_n8157 & ~new_n8158;
  assign new_n8160 = ~new_n8155 & ~new_n8159;
  assign new_n8161 = ~new_n8154 & ~new_n8160;
  assign new_n8162 = ~new_n8145 & new_n8161;
  assign new_n8163_1 = new_n8145 & ~new_n8161;
  assign new_n8164 = ~new_n8162 & ~new_n8163_1;
  assign new_n8165 = n5065 & n9216;
  assign new_n8166 = ~new_n8154 & ~new_n8155;
  assign new_n8167 = new_n8159 & ~new_n8166;
  assign new_n8168 = ~new_n8159 & new_n8166;
  assign new_n8169 = ~new_n8167 & ~new_n8168;
  assign new_n8170 = new_n8165 & ~new_n8169;
  assign new_n8171 = ~new_n8165 & new_n8169;
  assign new_n8172_1 = n1636 & n9216;
  assign new_n8173 = new_n4118 & new_n8137;
  assign new_n8174 = n5920 & n12348;
  assign new_n8175 = n2068 & n13058;
  assign new_n8176 = n4862 & n9216;
  assign new_n8177 = ~new_n8175 & ~new_n8176;
  assign new_n8178 = new_n8174 & ~new_n8177;
  assign new_n8179 = ~new_n8173 & ~new_n8178;
  assign new_n8180 = ~new_n8172_1 & new_n8179;
  assign new_n8181 = new_n8172_1 & ~new_n8179;
  assign new_n8182 = ~new_n8147 & ~new_n8150;
  assign new_n8183_1 = ~new_n8151 & ~new_n8182;
  assign new_n8184 = new_n8151 & new_n8182;
  assign new_n8185 = ~new_n8183_1 & ~new_n8184;
  assign new_n8186 = ~new_n8181 & ~new_n8185;
  assign new_n8187 = ~new_n8180 & ~new_n8186;
  assign new_n8188 = ~new_n8171 & new_n8187;
  assign new_n8189 = ~new_n8170 & ~new_n8188;
  assign new_n8190 = ~new_n8164 & ~new_n8189;
  assign new_n8191 = ~new_n8143 & new_n8161;
  assign new_n8192 = new_n8122 & new_n8191;
  assign new_n8193 = ~new_n8122 & ~new_n8191;
  assign new_n8194 = ~new_n8144 & new_n8193;
  assign new_n8195 = ~new_n8192 & ~new_n8194;
  assign new_n8196 = n9216 & n11835;
  assign new_n8197 = n2068 & n5065;
  assign new_n8198 = n443 & n12348;
  assign new_n8199 = ~new_n8197 & ~new_n8198;
  assign new_n8200 = new_n8197 & new_n8198;
  assign new_n8201 = ~new_n8199 & ~new_n8200;
  assign new_n8202 = new_n8196 & ~new_n8201;
  assign new_n8203 = ~new_n8196 & new_n8201;
  assign new_n8204 = ~new_n8202 & ~new_n8203;
  assign new_n8205 = ~new_n8131 & new_n8139_1;
  assign new_n8206 = ~new_n8130 & ~new_n8205;
  assign new_n8207 = ~new_n8204 & new_n8206;
  assign new_n8208 = new_n8204 & ~new_n8206;
  assign new_n8209 = ~new_n8207 & ~new_n8208;
  assign new_n8210 = n1636 & n11324;
  assign new_n8211 = new_n8128 & new_n8210;
  assign new_n8212 = ~new_n8128 & ~new_n8210;
  assign new_n8213 = ~new_n8211 & ~new_n8212;
  assign new_n8214 = n4862 & n8183;
  assign new_n8215 = n5920 & n10142;
  assign new_n8216 = n10657 & n13058;
  assign new_n8217 = ~new_n8215 & ~new_n8216;
  assign new_n8218 = new_n8215 & new_n8216;
  assign new_n8219_1 = ~new_n8217 & ~new_n8218;
  assign new_n8220 = new_n8214 & ~new_n8219_1;
  assign new_n8221 = ~new_n8214 & new_n8219_1;
  assign new_n8222 = ~new_n8220 & ~new_n8221;
  assign new_n8223 = new_n8213 & new_n8222;
  assign new_n8224 = ~new_n8213 & ~new_n8222;
  assign new_n8225 = ~new_n8223 & ~new_n8224;
  assign new_n8226 = ~new_n8209 & ~new_n8225;
  assign new_n8227 = new_n8209 & new_n8225;
  assign new_n8228_1 = ~new_n8226 & ~new_n8227;
  assign new_n8229 = new_n8195 & new_n8228_1;
  assign new_n8230_1 = ~new_n8195 & ~new_n8228_1;
  assign new_n8231 = ~new_n8229 & ~new_n8230_1;
  assign new_n8232 = ~new_n8190 & new_n8231;
  assign new_n8233_1 = new_n8190 & ~new_n8231;
  assign new_n8234 = ~new_n8232 & ~new_n8233_1;
  assign new_n8235 = n443 & n9216;
  assign new_n8236 = new_n8164 & new_n8189;
  assign new_n8237 = ~new_n8190 & ~new_n8236;
  assign new_n8238 = new_n8235 & new_n8237;
  assign new_n8239 = ~new_n8173 & ~new_n8177;
  assign new_n8240 = new_n4135 & ~new_n8239;
  assign new_n8241 = ~new_n8180 & ~new_n8181;
  assign new_n8242 = ~new_n8185 & ~new_n8241;
  assign new_n8243 = new_n8185 & new_n8241;
  assign new_n8244 = ~new_n8242 & ~new_n8243;
  assign new_n8245 = new_n8240 & new_n8244;
  assign new_n8246 = ~new_n8170 & ~new_n8171;
  assign new_n8247 = ~new_n8187 & ~new_n8246;
  assign new_n8248 = new_n8187 & new_n8246;
  assign new_n8249 = ~new_n8247 & ~new_n8248;
  assign new_n8250 = new_n8245 & new_n8249;
  assign new_n8251 = ~new_n8235 & ~new_n8237;
  assign new_n8252 = ~new_n8238 & ~new_n8251;
  assign new_n8253 = new_n8250 & new_n8252;
  assign new_n8254 = ~new_n8238 & ~new_n8253;
  assign new_n8255 = ~new_n8234 & new_n8254;
  assign new_n8256 = new_n8234 & ~new_n8254;
  assign new_n8257 = ~new_n8255 & ~new_n8256;
  assign new_n8258 = n3076 & n12592;
  assign new_n8259 = n10168 & n11634;
  assign new_n8260 = ~new_n8258 & ~new_n8259;
  assign new_n8261 = new_n8258 & new_n8259;
  assign new_n8262 = ~new_n8260 & ~new_n8261;
  assign new_n8263 = n767 & n817;
  assign new_n8264 = n951 & n5548;
  assign new_n8265_1 = n3815 & n11537;
  assign new_n8266 = ~new_n8264 & ~new_n8265_1;
  assign new_n8267 = new_n8264 & new_n8265_1;
  assign new_n8268 = ~new_n8266 & ~new_n8267;
  assign new_n8269 = ~new_n8263 & ~new_n8268;
  assign new_n8270 = new_n8263 & new_n8268;
  assign new_n8271 = ~new_n8269 & ~new_n8270;
  assign new_n8272 = n5548 & n10168;
  assign new_n8273 = n817 & n11537;
  assign new_n8274 = new_n8272 & new_n8273;
  assign new_n8275 = n767 & n3815;
  assign new_n8276 = n5548 & n11537;
  assign new_n8277 = n817 & n10168;
  assign new_n8278 = ~new_n8276 & ~new_n8277;
  assign new_n8279 = new_n8275 & ~new_n8278;
  assign new_n8280 = ~new_n8274 & ~new_n8279;
  assign new_n8281 = ~new_n8271 & new_n8280;
  assign new_n8282 = new_n8271 & ~new_n8280;
  assign new_n8283 = ~new_n8281 & ~new_n8282;
  assign new_n8284 = ~new_n8262 & ~new_n8283;
  assign new_n8285 = new_n8262 & new_n8283;
  assign new_n8286 = ~new_n8284 & ~new_n8285;
  assign new_n8287 = n11634 & n12592;
  assign new_n8288 = new_n4146 & new_n8263;
  assign new_n8289 = n767 & n5548;
  assign new_n8290_1 = n817 & n12592;
  assign new_n8291 = ~new_n8289 & ~new_n8290_1;
  assign new_n8292 = n3815 & n10168;
  assign new_n8293 = ~new_n8291 & new_n8292;
  assign new_n8294 = ~new_n8288 & ~new_n8293;
  assign new_n8295 = ~new_n8287 & new_n8294;
  assign new_n8296 = new_n8287 & ~new_n8294;
  assign new_n8297 = ~new_n8274 & ~new_n8278;
  assign new_n8298 = ~new_n8275 & ~new_n8297;
  assign new_n8299 = new_n8275 & new_n8297;
  assign new_n8300 = ~new_n8298 & ~new_n8299;
  assign new_n8301 = ~new_n8296 & ~new_n8300;
  assign new_n8302 = ~new_n8295 & ~new_n8301;
  assign new_n8303 = ~new_n8286 & ~new_n8302;
  assign new_n8304 = new_n8286 & new_n8302;
  assign new_n8305 = ~new_n8303 & ~new_n8304;
  assign new_n8306 = n3076 & n3178;
  assign new_n8307 = ~new_n8295 & ~new_n8296;
  assign new_n8308_1 = ~new_n8300 & ~new_n8307;
  assign new_n8309 = new_n8300 & new_n8307;
  assign new_n8310 = ~new_n8308_1 & ~new_n8309;
  assign new_n8311 = new_n8306 & new_n8310;
  assign new_n8312 = ~new_n8306 & ~new_n8310;
  assign new_n8313 = n3178 & n11634;
  assign new_n8314 = new_n4114_1 & new_n8277;
  assign new_n8315 = n3815 & n12592;
  assign new_n8316 = n817 & n3178;
  assign new_n8317 = ~new_n8272 & ~new_n8316;
  assign new_n8318 = new_n8315 & ~new_n8317;
  assign new_n8319 = ~new_n8314 & ~new_n8318;
  assign new_n8320 = ~new_n8313 & new_n8319;
  assign new_n8321 = new_n8313 & ~new_n8319;
  assign new_n8322 = ~new_n8288 & ~new_n8291;
  assign new_n8323 = ~new_n8292 & ~new_n8322;
  assign new_n8324 = new_n8292 & new_n8322;
  assign new_n8325 = ~new_n8323 & ~new_n8324;
  assign new_n8326 = ~new_n8321 & ~new_n8325;
  assign new_n8327 = ~new_n8320 & ~new_n8326;
  assign new_n8328 = ~new_n8312 & new_n8327;
  assign new_n8329 = ~new_n8311 & ~new_n8328;
  assign new_n8330 = new_n8305 & ~new_n8329;
  assign new_n8331 = ~new_n8284 & new_n8302;
  assign new_n8332_1 = ~new_n8261 & ~new_n8331;
  assign new_n8333 = ~new_n8285 & new_n8332_1;
  assign new_n8334 = new_n8261 & new_n8331;
  assign new_n8335 = ~new_n8333 & ~new_n8334;
  assign new_n8336_1 = n3178 & n7974;
  assign new_n8337 = n3076 & n10168;
  assign new_n8338 = n8163 & n12592;
  assign new_n8339 = ~new_n8337 & ~new_n8338;
  assign new_n8340 = n8163 & n10168;
  assign new_n8341 = new_n8258 & new_n8340;
  assign new_n8342 = ~new_n8339 & ~new_n8341;
  assign new_n8343 = ~new_n8336_1 & ~new_n8342;
  assign new_n8344 = new_n8336_1 & new_n8342;
  assign new_n8345 = ~new_n8343 & ~new_n8344;
  assign new_n8346 = ~new_n8270 & new_n8280;
  assign new_n8347 = ~new_n8269 & ~new_n8346;
  assign new_n8348 = ~new_n8345 & ~new_n8347;
  assign new_n8349 = new_n8345 & new_n8347;
  assign new_n8350 = ~new_n8348 & ~new_n8349;
  assign new_n8351 = n951 & n3815;
  assign new_n8352 = n401 & n5548;
  assign new_n8353 = ~new_n8351 & ~new_n8352;
  assign new_n8354 = n401 & n3815;
  assign new_n8355 = new_n8264 & new_n8354;
  assign new_n8356 = ~new_n8353 & ~new_n8355;
  assign new_n8357 = ~new_n8273 & ~new_n8356;
  assign new_n8358 = new_n8273 & new_n8356;
  assign new_n8359 = ~new_n8357 & ~new_n8358;
  assign new_n8360 = n767 & n11634;
  assign new_n8361 = ~new_n8267 & ~new_n8360;
  assign new_n8362 = new_n8267 & new_n8360;
  assign new_n8363 = ~new_n8361 & ~new_n8362;
  assign new_n8364 = ~new_n8359 & new_n8363;
  assign new_n8365 = new_n8359 & ~new_n8363;
  assign new_n8366 = ~new_n8364 & ~new_n8365;
  assign new_n8367 = ~new_n8350 & new_n8366;
  assign new_n8368 = new_n8350 & ~new_n8366;
  assign new_n8369 = ~new_n8367 & ~new_n8368;
  assign new_n8370 = new_n8335 & ~new_n8369;
  assign new_n8371 = ~new_n8335 & new_n8369;
  assign new_n8372 = ~new_n8370 & ~new_n8371;
  assign new_n8373 = new_n8330 & ~new_n8372;
  assign new_n8374 = ~new_n8330 & new_n8372;
  assign new_n8375 = ~new_n8373 & ~new_n8374;
  assign new_n8376 = n3178 & n8163;
  assign new_n8377 = ~new_n8305 & new_n8329;
  assign new_n8378 = ~new_n8330 & ~new_n8377;
  assign new_n8379 = new_n8376 & new_n8378;
  assign new_n8380 = ~new_n8314 & ~new_n8317;
  assign new_n8381 = new_n4148 & ~new_n8380;
  assign new_n8382 = ~new_n8320 & ~new_n8321;
  assign new_n8383 = ~new_n8325 & ~new_n8382;
  assign new_n8384 = new_n8325 & new_n8382;
  assign new_n8385 = ~new_n8383 & ~new_n8384;
  assign new_n8386 = new_n8381 & new_n8385;
  assign new_n8387 = ~new_n8311 & ~new_n8312;
  assign new_n8388 = ~new_n8327 & ~new_n8387;
  assign new_n8389 = new_n8327 & new_n8387;
  assign new_n8390 = ~new_n8388 & ~new_n8389;
  assign new_n8391 = new_n8386 & new_n8390;
  assign new_n8392 = ~new_n8376 & ~new_n8378;
  assign new_n8393 = ~new_n8379 & ~new_n8392;
  assign new_n8394 = new_n8391 & new_n8393;
  assign new_n8395 = ~new_n8379 & ~new_n8394;
  assign new_n8396 = new_n8375 & ~new_n8395;
  assign new_n8397 = ~new_n8375 & new_n8395;
  assign new_n8398 = ~new_n8396 & ~new_n8397;
  assign new_n8399 = n9 & n8860;
  assign new_n8400 = n1916 & n5031;
  assign new_n8401 = ~new_n8399 & ~new_n8400;
  assign new_n8402 = new_n8399 & new_n8400;
  assign new_n8403 = ~new_n8401 & ~new_n8402;
  assign new_n8404 = n2592 & n10162;
  assign new_n8405 = n2590 & n6392;
  assign new_n8406 = n3769 & n11061;
  assign new_n8407 = ~new_n8405 & ~new_n8406;
  assign new_n8408 = new_n8405 & new_n8406;
  assign new_n8409 = ~new_n8407 & ~new_n8408;
  assign new_n8410 = ~new_n8404 & ~new_n8409;
  assign new_n8411 = new_n8404 & new_n8409;
  assign new_n8412 = ~new_n8410 & ~new_n8411;
  assign new_n8413 = n2592 & n3769;
  assign new_n8414 = new_n8405 & new_n8413;
  assign new_n8415 = n9 & n10162;
  assign new_n8416 = n2590 & n3769;
  assign new_n8417 = n2592 & n6392;
  assign new_n8418 = ~new_n8416 & ~new_n8417;
  assign new_n8419 = new_n8415 & ~new_n8418;
  assign new_n8420 = ~new_n8414 & ~new_n8419;
  assign new_n8421 = ~new_n8412 & new_n8420;
  assign new_n8422 = new_n8412 & ~new_n8420;
  assign new_n8423 = ~new_n8421 & ~new_n8422;
  assign new_n8424 = ~new_n8403 & ~new_n8423;
  assign new_n8425 = new_n8403 & new_n8423;
  assign new_n8426 = ~new_n8424 & ~new_n8425;
  assign new_n8427 = n5031 & n8860;
  assign new_n8428 = new_n4138 & new_n8404;
  assign new_n8429 = n5031 & n10162;
  assign new_n8430 = ~new_n8413 & ~new_n8429;
  assign new_n8431 = n9 & n6392;
  assign new_n8432 = ~new_n8430 & new_n8431;
  assign new_n8433 = ~new_n8428 & ~new_n8432;
  assign new_n8434 = ~new_n8427 & new_n8433;
  assign new_n8435 = new_n8427 & ~new_n8433;
  assign new_n8436 = ~new_n8414 & ~new_n8418;
  assign new_n8437 = ~new_n8415 & ~new_n8436;
  assign new_n8438 = new_n8415 & new_n8436;
  assign new_n8439 = ~new_n8437 & ~new_n8438;
  assign new_n8440 = ~new_n8435 & ~new_n8439;
  assign new_n8441 = ~new_n8434 & ~new_n8440;
  assign new_n8442 = ~new_n8426 & new_n8441;
  assign new_n8443 = new_n8426 & ~new_n8441;
  assign new_n8444 = ~new_n8442 & ~new_n8443;
  assign new_n8445 = n1916 & n8466;
  assign new_n8446 = ~new_n8434 & ~new_n8435;
  assign new_n8447 = ~new_n8439 & ~new_n8446;
  assign new_n8448 = new_n8439 & new_n8446;
  assign new_n8449 = ~new_n8447 & ~new_n8448;
  assign new_n8450 = new_n8445 & new_n8449;
  assign new_n8451 = ~new_n8445 & ~new_n8449;
  assign new_n8452 = n8466 & n8860;
  assign new_n8453 = new_n4113 & new_n8415;
  assign new_n8454 = n5031 & n6392;
  assign new_n8455 = n9 & n3769;
  assign new_n8456 = n8466 & n10162;
  assign new_n8457 = ~new_n8455 & ~new_n8456;
  assign new_n8458 = new_n8454 & ~new_n8457;
  assign new_n8459 = ~new_n8453 & ~new_n8458;
  assign new_n8460 = ~new_n8452 & new_n8459;
  assign new_n8461 = new_n8452 & ~new_n8459;
  assign new_n8462 = ~new_n8428 & ~new_n8430;
  assign new_n8463 = ~new_n8431 & ~new_n8462;
  assign new_n8464 = new_n8431 & new_n8462;
  assign new_n8465 = ~new_n8463 & ~new_n8464;
  assign new_n8466_1 = ~new_n8461 & ~new_n8465;
  assign new_n8467 = ~new_n8460 & ~new_n8466_1;
  assign new_n8468_1 = ~new_n8451 & new_n8467;
  assign new_n8469 = ~new_n8450 & ~new_n8468_1;
  assign new_n8470 = ~new_n8444 & ~new_n8469;
  assign new_n8471 = ~new_n8424 & new_n8441;
  assign new_n8472 = ~new_n8402 & ~new_n8471;
  assign new_n8473 = ~new_n8425 & new_n8472;
  assign new_n8474 = new_n8402 & new_n8471;
  assign new_n8475 = ~new_n8473 & ~new_n8474;
  assign new_n8476 = n8466 & n11429;
  assign new_n8477 = n9 & n1916;
  assign new_n8478 = n5031 & n7374;
  assign new_n8479 = ~new_n8477 & ~new_n8478;
  assign new_n8480 = new_n8477 & new_n8478;
  assign new_n8481 = ~new_n8479 & ~new_n8480;
  assign new_n8482 = new_n8476 & ~new_n8481;
  assign new_n8483 = ~new_n8476 & new_n8481;
  assign new_n8484 = ~new_n8482 & ~new_n8483;
  assign new_n8485 = ~new_n8411 & new_n8420;
  assign new_n8486 = ~new_n8410 & ~new_n8485;
  assign new_n8487 = new_n8484 & ~new_n8486;
  assign new_n8488 = n2592 & n8860;
  assign new_n8489 = ~new_n8408 & ~new_n8488;
  assign new_n8490 = new_n8408 & new_n8488;
  assign new_n8491 = ~new_n8489 & ~new_n8490;
  assign new_n8492 = n2590 & n10162;
  assign new_n8493 = n6392 & n11061;
  assign new_n8494 = n3769 & n8768;
  assign new_n8495 = ~new_n8493 & ~new_n8494;
  assign new_n8496 = new_n8493 & new_n8494;
  assign new_n8497 = ~new_n8495 & ~new_n8496;
  assign new_n8498 = new_n8492 & ~new_n8497;
  assign new_n8499 = ~new_n8492 & new_n8497;
  assign new_n8500 = ~new_n8498 & ~new_n8499;
  assign new_n8501 = new_n8491 & new_n8500;
  assign new_n8502 = ~new_n8491 & ~new_n8500;
  assign new_n8503 = ~new_n8501 & ~new_n8502;
  assign new_n8504 = new_n8487 & new_n8503;
  assign new_n8505 = ~new_n8484 & new_n8486;
  assign new_n8506_1 = new_n8503 & ~new_n8505;
  assign new_n8507 = ~new_n8487 & ~new_n8506_1;
  assign new_n8508 = ~new_n8504 & ~new_n8507;
  assign new_n8509 = ~new_n8503 & new_n8505;
  assign new_n8510 = ~new_n8508 & ~new_n8509;
  assign new_n8511 = ~new_n8475 & new_n8510;
  assign new_n8512 = new_n8475 & ~new_n8510;
  assign new_n8513 = ~new_n8511 & ~new_n8512;
  assign new_n8514 = new_n8470 & new_n8513;
  assign new_n8515 = ~new_n8470 & ~new_n8513;
  assign new_n8516_1 = ~new_n8514 & ~new_n8515;
  assign new_n8517 = n7374 & n8466;
  assign new_n8518 = new_n8444 & new_n8469;
  assign new_n8519 = ~new_n8470 & ~new_n8518;
  assign new_n8520 = new_n8517 & new_n8519;
  assign new_n8521 = ~new_n8453 & ~new_n8457;
  assign new_n8522_1 = new_n4140 & ~new_n8521;
  assign new_n8523 = ~new_n8460 & ~new_n8461;
  assign new_n8524 = ~new_n8465 & ~new_n8523;
  assign new_n8525 = new_n8465 & new_n8523;
  assign new_n8526 = ~new_n8524 & ~new_n8525;
  assign new_n8527 = new_n8522_1 & new_n8526;
  assign new_n8528 = ~new_n8450 & ~new_n8451;
  assign new_n8529 = ~new_n8467 & ~new_n8528;
  assign new_n8530 = new_n8467 & new_n8528;
  assign new_n8531 = ~new_n8529 & ~new_n8530;
  assign new_n8532 = new_n8527 & new_n8531;
  assign new_n8533 = ~new_n8517 & ~new_n8519;
  assign new_n8534 = ~new_n8520 & ~new_n8533;
  assign new_n8535 = new_n8532 & new_n8534;
  assign new_n8536 = ~new_n8520 & ~new_n8535;
  assign new_n8537 = new_n8516_1 & ~new_n8536;
  assign new_n8538 = ~new_n8516_1 & new_n8536;
  assign new_n8539 = ~new_n8537 & ~new_n8538;
  assign new_n8540 = new_n8398 & new_n8539;
  assign new_n8541 = ~new_n8398 & ~new_n8539;
  assign new_n8542 = ~new_n8540 & ~new_n8541;
  assign new_n8543 = ~new_n8532 & ~new_n8534;
  assign new_n8544 = ~new_n8535 & ~new_n8543;
  assign new_n8545 = ~new_n8391 & ~new_n8393;
  assign new_n8546 = ~new_n8394 & ~new_n8545;
  assign new_n8547 = new_n8544 & new_n8546;
  assign new_n8548 = ~new_n8544 & ~new_n8546;
  assign new_n8549 = ~new_n8386 & ~new_n8390;
  assign new_n8550 = ~new_n8391 & ~new_n8549;
  assign new_n8551 = ~new_n8527 & ~new_n8531;
  assign new_n8552 = ~new_n8532 & ~new_n8551;
  assign new_n8553 = new_n8550 & new_n8552;
  assign new_n8554 = ~new_n8550 & ~new_n8552;
  assign new_n8555 = ~new_n8381 & ~new_n8385;
  assign new_n8556 = ~new_n8386 & ~new_n8555;
  assign new_n8557 = ~new_n8522_1 & ~new_n8526;
  assign new_n8558 = ~new_n8527 & ~new_n8557;
  assign new_n8559 = new_n8556 & new_n8558;
  assign new_n8560 = ~new_n8556 & ~new_n8558;
  assign new_n8561 = ~new_n4114_1 & new_n8315;
  assign new_n8562 = ~new_n8380 & ~new_n8561;
  assign new_n8563 = ~new_n4114_1 & new_n8318;
  assign new_n8564 = ~new_n8562 & ~new_n8563;
  assign new_n8565 = ~new_n4113 & new_n8454;
  assign new_n8566 = ~new_n8521 & ~new_n8565;
  assign new_n8567 = ~new_n4113 & new_n8458;
  assign new_n8568 = ~new_n8566 & ~new_n8567;
  assign new_n8569 = ~new_n8564 & ~new_n8568;
  assign new_n8570 = new_n8564 & new_n8568;
  assign new_n8571 = ~new_n4142 & ~new_n4151;
  assign new_n8572 = ~new_n8570 & ~new_n8571;
  assign new_n8573 = ~new_n8569 & ~new_n8572;
  assign new_n8574 = ~new_n8560 & new_n8573;
  assign new_n8575 = ~new_n8559 & ~new_n8574;
  assign new_n8576 = ~new_n8554 & ~new_n8575;
  assign new_n8577 = ~new_n8553 & ~new_n8576;
  assign new_n8578 = ~new_n8548 & ~new_n8577;
  assign new_n8579 = ~new_n8547 & ~new_n8578;
  assign new_n8580 = ~new_n8542 & ~new_n8579;
  assign new_n8581 = new_n8542 & new_n8579;
  assign new_n8582 = ~new_n8580 & ~new_n8581;
  assign new_n8583 = ~new_n8257 & new_n8582;
  assign new_n8584 = ~new_n8250 & ~new_n8252;
  assign new_n8585 = ~new_n8253 & ~new_n8584;
  assign new_n8586 = ~new_n8547 & ~new_n8548;
  assign new_n8587 = new_n8577 & ~new_n8586;
  assign new_n8588 = ~new_n8577 & new_n8586;
  assign new_n8589 = ~new_n8587 & ~new_n8588;
  assign new_n8590 = new_n8585 & new_n8589;
  assign new_n8591 = ~new_n8585 & ~new_n8589;
  assign new_n8592 = ~new_n8245 & ~new_n8249;
  assign new_n8593 = ~new_n8250 & ~new_n8592;
  assign new_n8594 = ~new_n8553 & ~new_n8554;
  assign new_n8595 = new_n8575 & ~new_n8594;
  assign new_n8596 = ~new_n8575 & new_n8594;
  assign new_n8597 = ~new_n8595 & ~new_n8596;
  assign new_n8598 = new_n8593 & new_n8597;
  assign new_n8599 = ~new_n8593 & ~new_n8597;
  assign new_n8600 = ~new_n8240 & ~new_n8244;
  assign new_n8601 = ~new_n8245 & ~new_n8600;
  assign new_n8602 = ~new_n8559 & ~new_n8560;
  assign new_n8603 = ~new_n8573 & ~new_n8602;
  assign new_n8604 = new_n8573 & new_n8602;
  assign new_n8605 = ~new_n8603 & ~new_n8604;
  assign new_n8606 = new_n8601 & new_n8605;
  assign new_n8607 = ~new_n8601 & ~new_n8605;
  assign new_n8608 = ~new_n8569 & ~new_n8570;
  assign new_n8609 = new_n8571 & ~new_n8608;
  assign new_n8610 = ~new_n8571 & new_n8608;
  assign new_n8611 = ~new_n8609 & ~new_n8610;
  assign new_n8612 = ~new_n4118 & new_n8174;
  assign new_n8613 = ~new_n8239 & ~new_n8612;
  assign new_n8614 = ~new_n4118 & new_n8178;
  assign new_n8615 = ~new_n8613 & ~new_n8614;
  assign new_n8616 = ~new_n8611 & new_n8615;
  assign new_n8617 = new_n8611 & ~new_n8615;
  assign new_n8618 = new_n4119 & ~new_n4155;
  assign new_n8619 = ~new_n4154 & ~new_n8618;
  assign new_n8620 = ~new_n8617 & ~new_n8619;
  assign new_n8621 = ~new_n8616 & ~new_n8620;
  assign new_n8622 = ~new_n8607 & ~new_n8621;
  assign new_n8623 = ~new_n8606 & ~new_n8622;
  assign new_n8624 = ~new_n8599 & ~new_n8623;
  assign new_n8625 = ~new_n8598 & ~new_n8624;
  assign new_n8626 = ~new_n8591 & ~new_n8625;
  assign new_n8627 = ~new_n8590 & ~new_n8626;
  assign new_n8628 = new_n8583 & new_n8627;
  assign new_n8629 = new_n8257 & ~new_n8582;
  assign new_n8630 = ~new_n8627 & new_n8629;
  assign new_n8631 = ~new_n8583 & ~new_n8627;
  assign new_n8632 = ~new_n8629 & ~new_n8631;
  assign new_n8633 = ~new_n8630 & ~new_n8632;
  assign new_n8634 = ~new_n8628 & ~new_n8633;
  assign new_n8635 = new_n8118 & new_n8634;
  assign new_n8636 = ~new_n8118 & ~new_n8634;
  assign new_n8637 = ~new_n8067 & ~new_n8069;
  assign new_n8638 = ~new_n8070 & ~new_n8637;
  assign new_n8639 = ~new_n8062 & ~new_n8066;
  assign new_n8640 = ~new_n8067 & ~new_n8639;
  assign new_n8641 = ~new_n8598 & ~new_n8599;
  assign new_n8642 = new_n8623 & ~new_n8641;
  assign new_n8643 = ~new_n8623 & new_n8641;
  assign new_n8644 = ~new_n8642 & ~new_n8643;
  assign new_n8645 = new_n8640 & new_n8644;
  assign new_n8646 = ~new_n8640 & ~new_n8644;
  assign new_n8647 = ~new_n8057 & ~new_n8061;
  assign new_n8648 = ~new_n8062 & ~new_n8647;
  assign new_n8649 = ~new_n8606 & ~new_n8607;
  assign new_n8650 = ~new_n8621 & new_n8649;
  assign new_n8651 = new_n8621 & ~new_n8649;
  assign new_n8652 = ~new_n8650 & ~new_n8651;
  assign new_n8653 = new_n8648 & new_n8652;
  assign new_n8654 = ~new_n8648 & ~new_n8652;
  assign new_n8655 = ~new_n4122_1 & new_n8036;
  assign new_n8656 = ~new_n8056 & ~new_n8655;
  assign new_n8657 = ~new_n4122_1 & new_n8040;
  assign new_n8658 = ~new_n8656 & ~new_n8657;
  assign new_n8659 = ~new_n8616 & ~new_n8617;
  assign new_n8660 = ~new_n8619 & ~new_n8659;
  assign new_n8661 = new_n8619 & new_n8659;
  assign new_n8662 = ~new_n8660 & ~new_n8661;
  assign new_n8663 = new_n8658 & ~new_n8662;
  assign new_n8664 = ~new_n8658 & new_n8662;
  assign new_n8665 = ~new_n4129 & ~new_n4159;
  assign new_n8666 = ~new_n4130 & ~new_n8665;
  assign new_n8667 = ~new_n8664 & ~new_n8666;
  assign new_n8668 = ~new_n8663 & ~new_n8667;
  assign new_n8669 = ~new_n8654 & ~new_n8668;
  assign new_n8670 = ~new_n8653 & ~new_n8669;
  assign new_n8671 = ~new_n8646 & ~new_n8670;
  assign new_n8672 = ~new_n8645 & ~new_n8671;
  assign new_n8673 = new_n8638 & ~new_n8672;
  assign new_n8674 = ~new_n8638 & new_n8672;
  assign new_n8675 = ~new_n8590 & ~new_n8591;
  assign new_n8676 = new_n8625 & ~new_n8675;
  assign new_n8677 = ~new_n8625 & new_n8675;
  assign new_n8678 = ~new_n8676 & ~new_n8677;
  assign new_n8679 = ~new_n8674 & new_n8678;
  assign new_n8680 = ~new_n8673 & ~new_n8679;
  assign new_n8681 = ~new_n8636 & ~new_n8680;
  assign new_n8682 = ~new_n8635 & ~new_n8681;
  assign new_n8683 = ~new_n8514 & ~new_n8537;
  assign new_n8684 = ~new_n8113 & ~new_n8116;
  assign new_n8685 = ~new_n8683 & new_n8684;
  assign new_n8686 = new_n8683 & ~new_n8684;
  assign new_n8687 = ~new_n8685 & ~new_n8686;
  assign new_n8688 = new_n8492 & ~new_n8495;
  assign new_n8689 = ~new_n8496 & ~new_n8688;
  assign new_n8690 = new_n8476 & ~new_n8479;
  assign new_n8691 = ~new_n8480 & ~new_n8690;
  assign new_n8692 = ~new_n8689 & new_n8691;
  assign new_n8693 = new_n8689 & ~new_n8691;
  assign new_n8694 = ~new_n8692 & ~new_n8693;
  assign new_n8695 = ~new_n8104 & ~new_n8107;
  assign new_n8696 = ~new_n8108 & ~new_n8695;
  assign new_n8697 = n6668 & n7659;
  assign new_n8698 = n7812 & n12289;
  assign new_n8699 = n7772 & n10122;
  assign new_n8700 = new_n8698 & ~new_n8699;
  assign new_n8701_1 = ~new_n8698 & new_n8699;
  assign new_n8702 = ~new_n8700 & ~new_n8701_1;
  assign new_n8703 = new_n8697 & ~new_n8702;
  assign new_n8704 = ~new_n8697 & new_n8702;
  assign new_n8705 = ~new_n8703 & ~new_n8704;
  assign new_n8706 = ~new_n8490 & new_n8500;
  assign new_n8707 = ~new_n8489 & ~new_n8706;
  assign new_n8708 = ~new_n8705 & ~new_n8707;
  assign new_n8709 = new_n8705 & new_n8707;
  assign new_n8710 = ~new_n8708 & ~new_n8709;
  assign new_n8711 = new_n8696 & ~new_n8710;
  assign new_n8712 = ~new_n8696 & new_n8710;
  assign new_n8713 = ~new_n8711 & ~new_n8712;
  assign new_n8714 = ~new_n8348 & ~new_n8366;
  assign new_n8715 = ~new_n8349 & ~new_n8714;
  assign new_n8716_1 = n4075 & n8466;
  assign new_n8717 = n2590 & n8860;
  assign new_n8718 = ~new_n8716_1 & new_n8717;
  assign new_n8719 = new_n8716_1 & ~new_n8717;
  assign new_n8720 = ~new_n8718 & ~new_n8719;
  assign new_n8721 = n9 & n7374;
  assign new_n8722 = n5031 & n11429;
  assign new_n8723 = ~new_n8721 & ~new_n8722;
  assign new_n8724 = new_n8721 & new_n8722;
  assign new_n8725 = ~new_n8723 & ~new_n8724;
  assign new_n8726 = ~new_n8720 & new_n8725;
  assign new_n8727 = new_n8720 & ~new_n8725;
  assign new_n8728 = ~new_n8726 & ~new_n8727;
  assign new_n8729 = new_n8336_1 & ~new_n8339;
  assign new_n8730 = ~new_n8341 & ~new_n8729;
  assign new_n8731 = n3769 & n4998;
  assign new_n8732 = n1916 & n2592;
  assign new_n8733 = new_n8731 & ~new_n8732;
  assign new_n8734 = ~new_n8731 & new_n8732;
  assign new_n8735 = ~new_n8733 & ~new_n8734;
  assign new_n8736 = n6392 & n8768;
  assign new_n8737 = n10162 & n11061;
  assign new_n8738 = new_n8736 & ~new_n8737;
  assign new_n8739 = ~new_n8736 & new_n8737;
  assign new_n8740 = ~new_n8738 & ~new_n8739;
  assign new_n8741 = ~new_n8735 & ~new_n8740;
  assign new_n8742 = new_n8735 & new_n8740;
  assign new_n8743 = ~new_n8741 & ~new_n8742;
  assign new_n8744 = new_n8730 & new_n8743;
  assign new_n8745 = ~new_n8730 & ~new_n8743;
  assign new_n8746 = ~new_n8744 & ~new_n8745;
  assign new_n8747 = new_n8728 & ~new_n8746;
  assign new_n8748 = ~new_n8728 & new_n8746;
  assign new_n8749 = ~new_n8747 & ~new_n8748;
  assign new_n8750 = ~new_n8715 & ~new_n8749;
  assign new_n8751 = new_n8715 & new_n8749;
  assign new_n8752 = ~new_n8750 & ~new_n8751;
  assign new_n8753 = new_n8359 & ~new_n8361;
  assign new_n8754 = ~new_n8362 & ~new_n8753;
  assign new_n8755 = new_n8273 & ~new_n8353;
  assign new_n8756 = ~new_n8355 & ~new_n8755;
  assign new_n8757 = n7974 & n12592;
  assign new_n8758 = ~new_n8340 & new_n8757;
  assign new_n8759 = new_n8340 & ~new_n8757;
  assign new_n8760 = ~new_n8758 & ~new_n8759;
  assign new_n8761 = new_n8756 & ~new_n8760;
  assign new_n8762 = ~new_n8756 & new_n8760;
  assign new_n8763 = ~new_n8761 & ~new_n8762;
  assign new_n8764 = ~new_n8754 & new_n8763;
  assign new_n8765 = new_n8754 & ~new_n8763;
  assign new_n8766 = ~new_n8764 & ~new_n8765;
  assign new_n8767 = ~new_n8752 & new_n8766;
  assign new_n8768_1 = new_n8752 & ~new_n8766;
  assign new_n8769 = ~new_n8767 & ~new_n8768_1;
  assign new_n8770 = ~new_n8473 & ~new_n8510;
  assign new_n8771 = ~new_n8474 & ~new_n8770;
  assign new_n8772 = new_n8507 & new_n8771;
  assign new_n8773 = ~new_n8507 & ~new_n8771;
  assign new_n8774 = ~new_n8772 & ~new_n8773;
  assign new_n8775 = new_n8769 & ~new_n8774;
  assign new_n8776 = ~new_n8769 & new_n8774;
  assign new_n8777 = ~new_n8775 & ~new_n8776;
  assign new_n8778 = ~new_n8713 & ~new_n8777;
  assign new_n8779 = new_n8713 & new_n8777;
  assign new_n8780 = ~new_n8778 & ~new_n8779;
  assign new_n8781 = ~new_n8694 & new_n8780;
  assign new_n8782 = new_n8694 & ~new_n8780;
  assign new_n8783 = ~new_n8781 & ~new_n8782;
  assign new_n8784 = ~new_n8541 & ~new_n8579;
  assign new_n8785 = ~new_n8540 & ~new_n8784;
  assign new_n8786 = n4452 & n13058;
  assign new_n8787 = ~new_n8087 & new_n8098;
  assign new_n8788 = ~new_n8088 & ~new_n8787;
  assign new_n8789 = n4330 & n8230;
  assign new_n8790 = n2252 & n2458;
  assign new_n8791 = ~new_n8789 & ~new_n8790;
  assign new_n8792 = new_n8789 & new_n8790;
  assign new_n8793 = ~new_n8791 & ~new_n8792;
  assign new_n8794 = n7715 & n9747;
  assign new_n8795 = n5884 & n7529;
  assign new_n8796 = new_n8794 & ~new_n8795;
  assign new_n8797 = ~new_n8794 & new_n8795;
  assign new_n8798 = ~new_n8796 & ~new_n8797;
  assign new_n8799 = ~new_n8793 & ~new_n8798;
  assign new_n8800 = new_n8793 & new_n8798;
  assign new_n8801 = ~new_n8799 & ~new_n8800;
  assign new_n8802 = new_n8090 & ~new_n8093;
  assign new_n8803 = ~new_n8094 & ~new_n8802;
  assign new_n8804 = new_n8072 & ~new_n8075;
  assign new_n8805 = ~new_n8076 & ~new_n8804;
  assign new_n8806 = ~new_n8803 & new_n8805;
  assign new_n8807 = new_n8803 & ~new_n8805;
  assign new_n8808 = ~new_n8806 & ~new_n8807;
  assign new_n8809 = ~new_n8801 & new_n8808;
  assign new_n8810 = new_n8801 & ~new_n8808;
  assign new_n8811 = ~new_n8809 & ~new_n8810;
  assign new_n8812 = new_n8788 & new_n8811;
  assign new_n8813 = ~new_n8788 & ~new_n8811;
  assign new_n8814 = ~new_n8812 & ~new_n8813;
  assign new_n8815 = ~new_n8084 & new_n8101;
  assign new_n8816 = ~new_n8083 & ~new_n8815;
  assign new_n8817 = ~new_n8814 & new_n8816;
  assign new_n8818 = new_n8814 & ~new_n8816;
  assign new_n8819 = ~new_n8817 & ~new_n8818;
  assign new_n8820_1 = ~new_n8786 & new_n8819;
  assign new_n8821 = new_n8786 & ~new_n8819;
  assign new_n8822 = ~new_n8820_1 & ~new_n8821;
  assign new_n8823 = ~new_n8194 & ~new_n8228_1;
  assign new_n8824 = ~new_n8192 & ~new_n8823;
  assign new_n8825 = n5356 & n9216;
  assign new_n8826 = n1636 & n8183;
  assign new_n8827 = new_n8825 & ~new_n8826;
  assign new_n8828 = ~new_n8825 & new_n8826;
  assign new_n8829 = ~new_n8827 & ~new_n8828;
  assign new_n8830 = n5920 & n10657;
  assign new_n8831 = n4862 & n10142;
  assign new_n8832 = ~new_n8830 & ~new_n8831;
  assign new_n8833 = new_n8830 & new_n8831;
  assign new_n8834 = ~new_n8832 & ~new_n8833;
  assign new_n8835 = ~new_n8829 & new_n8834;
  assign new_n8836 = new_n8829 & ~new_n8834;
  assign new_n8837 = ~new_n8835 & ~new_n8836;
  assign new_n8838 = ~new_n8824 & new_n8837;
  assign new_n8839 = new_n8824 & ~new_n8837;
  assign new_n8840 = ~new_n8838 & ~new_n8839;
  assign new_n8841 = ~new_n8822 & ~new_n8840;
  assign new_n8842 = new_n8822 & new_n8840;
  assign new_n8843 = ~new_n8841 & ~new_n8842;
  assign new_n8844 = ~new_n8785 & new_n8843;
  assign new_n8845 = new_n8785 & ~new_n8843;
  assign new_n8846 = ~new_n8844 & ~new_n8845;
  assign new_n8847 = ~new_n8373 & ~new_n8396;
  assign new_n8848 = ~new_n8333 & new_n8369;
  assign new_n8849 = ~new_n8334 & ~new_n8848;
  assign new_n8850 = n817 & n951;
  assign new_n8851 = n767 & n3076;
  assign new_n8852 = ~new_n8850 & new_n8851;
  assign new_n8853 = new_n8850 & ~new_n8851;
  assign new_n8854 = ~new_n8852 & ~new_n8853;
  assign new_n8855 = n11537 & n11634;
  assign new_n8856 = ~new_n8354 & ~new_n8855;
  assign new_n8857 = new_n8354 & new_n8855;
  assign new_n8858 = ~new_n8856 & ~new_n8857;
  assign new_n8859_1 = ~new_n8854 & new_n8858;
  assign new_n8860_1 = new_n8854 & ~new_n8858;
  assign new_n8861 = ~new_n8859_1 & ~new_n8860_1;
  assign new_n8862 = n4419 & n5548;
  assign new_n8863 = n1709 & n3178;
  assign new_n8864 = ~new_n8862 & new_n8863;
  assign new_n8865 = new_n8862 & ~new_n8863;
  assign new_n8866 = ~new_n8864 & ~new_n8865;
  assign new_n8867 = ~new_n8861 & new_n8866;
  assign new_n8868 = new_n8861 & ~new_n8866;
  assign new_n8869 = ~new_n8867 & ~new_n8868;
  assign new_n8870 = ~new_n8208 & ~new_n8225;
  assign new_n8871 = ~new_n8207 & ~new_n8870;
  assign new_n8872 = ~new_n8211 & new_n8222;
  assign new_n8873 = ~new_n8212 & ~new_n8872;
  assign new_n8874 = ~new_n8871 & new_n8873;
  assign new_n8875 = new_n8871 & ~new_n8873;
  assign new_n8876 = ~new_n8874 & ~new_n8875;
  assign new_n8877 = ~new_n8869 & new_n8876;
  assign new_n8878 = new_n8869 & ~new_n8876;
  assign new_n8879 = ~new_n8877 & ~new_n8878;
  assign new_n8880 = ~new_n8849 & new_n8879;
  assign new_n8881 = new_n8849 & ~new_n8879;
  assign new_n8882 = ~new_n8880 & ~new_n8881;
  assign new_n8883 = n11835 & n12348;
  assign new_n8884 = n443 & n2068;
  assign new_n8885 = n5065 & n11324;
  assign new_n8886 = new_n8884 & new_n8885;
  assign new_n8887 = ~new_n8884 & ~new_n8885;
  assign new_n8888 = ~new_n8886 & ~new_n8887;
  assign new_n8889 = new_n8883 & ~new_n8888;
  assign new_n8890 = ~new_n8883 & new_n8888;
  assign new_n8891 = ~new_n8889 & ~new_n8890;
  assign new_n8892 = new_n8196 & ~new_n8199;
  assign new_n8893 = ~new_n8200 & ~new_n8892;
  assign new_n8894 = new_n8214 & ~new_n8217;
  assign new_n8895 = ~new_n8218 & ~new_n8894;
  assign new_n8896 = ~new_n8893 & new_n8895;
  assign new_n8897 = new_n8893 & ~new_n8895;
  assign new_n8898 = ~new_n8896 & ~new_n8897;
  assign new_n8899 = ~new_n8891 & ~new_n8898;
  assign new_n8900 = new_n8891 & new_n8898;
  assign new_n8901 = ~new_n8899 & ~new_n8900;
  assign new_n8902 = ~new_n8882 & new_n8901;
  assign new_n8903 = new_n8882 & ~new_n8901;
  assign new_n8904 = ~new_n8902 & ~new_n8903;
  assign new_n8905 = new_n8847 & ~new_n8904;
  assign new_n8906 = ~new_n8847 & new_n8904;
  assign new_n8907 = ~new_n8905 & ~new_n8906;
  assign new_n8908 = ~new_n8233_1 & ~new_n8256;
  assign new_n8909 = new_n8907 & new_n8908;
  assign new_n8910 = ~new_n8907 & ~new_n8908;
  assign new_n8911 = ~new_n8909 & ~new_n8910;
  assign new_n8912 = new_n8846 & new_n8911;
  assign new_n8913 = ~new_n8846 & ~new_n8911;
  assign new_n8914 = ~new_n8912 & ~new_n8913;
  assign new_n8915 = new_n8632 & new_n8914;
  assign new_n8916 = ~new_n8632 & ~new_n8914;
  assign new_n8917 = ~new_n8915 & ~new_n8916;
  assign new_n8918 = new_n8783 & new_n8917;
  assign new_n8919 = ~new_n8783 & ~new_n8917;
  assign new_n8920 = ~new_n8918 & ~new_n8919;
  assign new_n8921 = ~new_n8687 & new_n8920;
  assign new_n8922 = new_n8687 & ~new_n8920;
  assign new_n8923 = ~new_n8921 & ~new_n8922;
  assign new_n8924 = new_n8682 & ~new_n8923;
  assign new_n8925 = ~new_n8682 & new_n8923;
  assign n2061 = new_n8924 | new_n8925;
  assign new_n8927 = ~new_n3489 & ~new_n3490;
  assign new_n8928 = new_n3520 & ~new_n8927;
  assign new_n8929 = ~new_n3520 & new_n8927;
  assign n2190 = ~new_n8928 & ~new_n8929;
  assign new_n8931 = n5962 & n9216;
  assign new_n8932 = n287 & n8466;
  assign new_n8933 = n3178 & n11058;
  assign new_n8934 = new_n8932 & new_n8933;
  assign new_n8935 = ~new_n8932 & ~new_n8933;
  assign new_n8936 = ~new_n8934 & ~new_n8935;
  assign new_n8937 = new_n8931 & new_n8936;
  assign new_n8938 = ~new_n8931 & ~new_n8936;
  assign new_n8939 = ~new_n8937 & ~new_n8938;
  assign new_n8940_1 = n7772 & n10451;
  assign new_n8941 = new_n8939 & new_n8940_1;
  assign new_n8942 = n7772 & n9093;
  assign new_n8943 = n7529 & n10451;
  assign new_n8944 = ~new_n8942 & ~new_n8943;
  assign new_n8945 = new_n8942 & new_n8943;
  assign new_n8946 = ~new_n8944 & ~new_n8945;
  assign new_n8947 = ~new_n8941 & ~new_n8946;
  assign new_n8948 = new_n8941 & new_n8946;
  assign new_n8949 = ~new_n8947 & ~new_n8948;
  assign new_n8950 = n6085 & n9216;
  assign new_n8951 = n5962 & n12348;
  assign new_n8952 = ~new_n8950 & ~new_n8951;
  assign new_n8953 = new_n8950 & new_n8951;
  assign new_n8954 = ~new_n8952 & ~new_n8953;
  assign new_n8955 = new_n8937 & new_n8954;
  assign new_n8956 = ~new_n8937 & ~new_n8954;
  assign new_n8957 = ~new_n8955 & ~new_n8956;
  assign new_n8958 = n7720 & n8466;
  assign new_n8959 = n287 & n5031;
  assign new_n8960 = ~new_n8958 & ~new_n8959;
  assign new_n8961 = new_n8958 & new_n8959;
  assign new_n8962 = ~new_n8960 & ~new_n8961;
  assign new_n8963 = ~new_n8934 & ~new_n8962;
  assign new_n8964 = new_n8934 & new_n8962;
  assign new_n8965 = ~new_n8963 & ~new_n8964;
  assign new_n8966 = n1007 & n3178;
  assign new_n8967 = n11058 & n12592;
  assign new_n8968 = ~new_n8966 & ~new_n8967;
  assign new_n8969 = new_n8966 & new_n8967;
  assign new_n8970 = ~new_n8968 & ~new_n8969;
  assign new_n8971 = ~new_n8965 & new_n8970;
  assign new_n8972 = new_n8965 & ~new_n8970;
  assign new_n8973 = ~new_n8971 & ~new_n8972;
  assign new_n8974 = new_n8957 & new_n8973;
  assign new_n8975 = ~new_n8957 & ~new_n8973;
  assign new_n8976 = ~new_n8974 & ~new_n8975;
  assign new_n8977 = new_n8949 & ~new_n8976;
  assign new_n8978 = ~new_n8949 & new_n8976;
  assign n2235 = ~new_n8977 & ~new_n8978;
  assign new_n8980 = ~new_n3511 & ~new_n3512;
  assign new_n8981 = new_n3514 & ~new_n8980;
  assign new_n8982 = ~new_n3514 & new_n8980;
  assign n2549 = new_n8981 | new_n8982;
  assign new_n8984 = ~new_n4887 & ~new_n4888;
  assign new_n8985 = new_n4902 & ~new_n8984;
  assign new_n8986 = ~new_n4902 & new_n8984;
  assign n2709 = ~new_n8985 & ~new_n8986;
  assign new_n8988 = ~new_n4889 & ~new_n4891;
  assign n2805 = ~new_n4892 & ~new_n8988;
  assign new_n8990 = ~new_n412 & ~new_n413;
  assign new_n8991 = ~new_n417 & new_n8990;
  assign new_n8992 = new_n417 & ~new_n8990;
  assign n2904 = new_n8991 | new_n8992;
  assign new_n8994 = ~new_n1973 & ~new_n1974;
  assign new_n8995 = new_n1998 & ~new_n8994;
  assign new_n8996 = ~new_n1998 & new_n8994;
  assign n2934 = ~new_n8995 & ~new_n8996;
  assign new_n8998 = ~new_n1366 & ~new_n1367;
  assign new_n8999 = ~new_n1391 & ~new_n8998;
  assign new_n9000 = new_n1391 & new_n8998;
  assign n3262 = ~new_n8999 & ~new_n9000;
  assign new_n9002 = n5801 & n9475;
  assign new_n9003 = n411 & n10908;
  assign new_n9004 = new_n9002 & new_n9003;
  assign new_n9005 = n411 & n10560;
  assign new_n9006 = n9475 & n10908;
  assign new_n9007 = n5801 & n6826;
  assign new_n9008 = ~new_n9006 & ~new_n9007;
  assign new_n9009 = new_n9006 & new_n9007;
  assign new_n9010 = ~new_n9008 & ~new_n9009;
  assign new_n9011 = new_n9005 & ~new_n9010;
  assign new_n9012 = ~new_n9005 & new_n9010;
  assign new_n9013 = ~new_n9011 & ~new_n9012;
  assign new_n9014 = new_n9004 & ~new_n9013;
  assign new_n9015 = n5801 & n12284;
  assign new_n9016 = new_n9005 & ~new_n9008;
  assign new_n9017 = ~new_n9009 & ~new_n9016;
  assign new_n9018 = ~new_n9015 & new_n9017;
  assign new_n9019 = new_n9015 & ~new_n9017;
  assign new_n9020 = ~new_n9018 & ~new_n9019;
  assign new_n9021 = n411 & n12003;
  assign new_n9022 = n6826 & n10908;
  assign new_n9023 = n9475 & n10560;
  assign new_n9024 = ~new_n9022 & ~new_n9023;
  assign new_n9025 = new_n9022 & new_n9023;
  assign new_n9026 = ~new_n9024 & ~new_n9025;
  assign new_n9027 = new_n9021 & ~new_n9026;
  assign new_n9028 = ~new_n9021 & new_n9026;
  assign new_n9029 = ~new_n9027 & ~new_n9028;
  assign new_n9030 = ~new_n9020 & new_n9029;
  assign new_n9031 = new_n9020 & ~new_n9029;
  assign new_n9032 = ~new_n9030 & ~new_n9031;
  assign new_n9033 = new_n9014 & new_n9032;
  assign new_n9034 = n469 & n5801;
  assign new_n9035 = n10908 & n12284;
  assign new_n9036 = new_n9021 & ~new_n9024;
  assign new_n9037 = ~new_n9025 & ~new_n9036;
  assign new_n9038 = ~new_n9035 & new_n9037;
  assign new_n9039 = new_n9035 & ~new_n9037;
  assign new_n9040 = ~new_n9038 & ~new_n9039;
  assign new_n9041_1 = n411 & n8139;
  assign new_n9042 = n6826 & n10560;
  assign new_n9043 = n9475 & n12003;
  assign new_n9044 = ~new_n9042 & ~new_n9043;
  assign new_n9045 = new_n9042 & new_n9043;
  assign new_n9046 = ~new_n9044 & ~new_n9045;
  assign new_n9047 = new_n9041_1 & ~new_n9046;
  assign new_n9048 = ~new_n9041_1 & new_n9046;
  assign new_n9049 = ~new_n9047 & ~new_n9048;
  assign new_n9050 = ~new_n9040 & new_n9049;
  assign new_n9051 = new_n9040 & ~new_n9049;
  assign new_n9052 = ~new_n9050 & ~new_n9051;
  assign new_n9053 = ~new_n9034 & ~new_n9052;
  assign new_n9054 = new_n9034 & new_n9052;
  assign new_n9055 = ~new_n9053 & ~new_n9054;
  assign new_n9056 = ~new_n9018 & ~new_n9029;
  assign new_n9057 = ~new_n9019 & ~new_n9056;
  assign new_n9058 = ~new_n9055 & new_n9057;
  assign new_n9059 = new_n9055 & ~new_n9057;
  assign new_n9060 = ~new_n9058 & ~new_n9059;
  assign new_n9061 = ~new_n9033 & ~new_n9060;
  assign new_n9062 = new_n9033 & new_n9060;
  assign new_n9063 = ~new_n9061 & ~new_n9062;
  assign new_n9064 = n5536 & n5671;
  assign new_n9065 = n4114 & n8506;
  assign new_n9066 = new_n9064 & new_n9065;
  assign new_n9067 = n8506 & n11665;
  assign new_n9068 = n4114 & n5536;
  assign new_n9069 = n772 & n5671;
  assign new_n9070 = ~new_n9068 & ~new_n9069;
  assign new_n9071 = new_n9068 & new_n9069;
  assign new_n9072 = ~new_n9070 & ~new_n9071;
  assign new_n9073 = new_n9067 & ~new_n9072;
  assign new_n9074 = ~new_n9067 & new_n9072;
  assign new_n9075 = ~new_n9073 & ~new_n9074;
  assign new_n9076 = new_n9066 & ~new_n9075;
  assign new_n9077 = n2737 & n5671;
  assign new_n9078 = new_n9067 & ~new_n9070;
  assign new_n9079 = ~new_n9071 & ~new_n9078;
  assign new_n9080 = ~new_n9077 & new_n9079;
  assign new_n9081 = new_n9077 & ~new_n9079;
  assign new_n9082 = ~new_n9080 & ~new_n9081;
  assign new_n9083 = n2777 & n8506;
  assign new_n9084 = n772 & n4114;
  assign new_n9085 = n5536 & n11665;
  assign new_n9086 = ~new_n9084 & ~new_n9085;
  assign new_n9087 = new_n9084 & new_n9085;
  assign new_n9088 = ~new_n9086 & ~new_n9087;
  assign new_n9089 = new_n9083 & ~new_n9088;
  assign new_n9090 = ~new_n9083 & new_n9088;
  assign new_n9091 = ~new_n9089 & ~new_n9090;
  assign new_n9092 = ~new_n9082 & new_n9091;
  assign new_n9093_1 = new_n9082 & ~new_n9091;
  assign new_n9094 = ~new_n9092 & ~new_n9093_1;
  assign new_n9095 = new_n9076 & new_n9094;
  assign new_n9096 = n5671 & n12408;
  assign new_n9097 = n2737 & n4114;
  assign new_n9098 = new_n9083 & ~new_n9086;
  assign new_n9099 = ~new_n9087 & ~new_n9098;
  assign new_n9100_1 = ~new_n9097 & new_n9099;
  assign new_n9101 = new_n9097 & ~new_n9099;
  assign new_n9102 = ~new_n9100_1 & ~new_n9101;
  assign new_n9103 = n8506 & n10642;
  assign new_n9104 = n772 & n11665;
  assign new_n9105 = n2777 & n5536;
  assign new_n9106 = ~new_n9104 & ~new_n9105;
  assign new_n9107 = new_n9104 & new_n9105;
  assign new_n9108 = ~new_n9106 & ~new_n9107;
  assign new_n9109 = new_n9103 & ~new_n9108;
  assign new_n9110 = ~new_n9103 & new_n9108;
  assign new_n9111 = ~new_n9109 & ~new_n9110;
  assign new_n9112 = ~new_n9102 & new_n9111;
  assign new_n9113 = new_n9102 & ~new_n9111;
  assign new_n9114 = ~new_n9112 & ~new_n9113;
  assign new_n9115 = ~new_n9096 & ~new_n9114;
  assign new_n9116 = new_n9096 & new_n9114;
  assign new_n9117 = ~new_n9115 & ~new_n9116;
  assign new_n9118 = ~new_n9080 & ~new_n9091;
  assign new_n9119 = ~new_n9081 & ~new_n9118;
  assign new_n9120 = ~new_n9117 & new_n9119;
  assign new_n9121 = new_n9117 & ~new_n9119;
  assign new_n9122 = ~new_n9120 & ~new_n9121;
  assign new_n9123 = ~new_n9095 & ~new_n9122;
  assign new_n9124 = new_n9095 & new_n9122;
  assign new_n9125 = ~new_n9123 & ~new_n9124;
  assign new_n9126 = n124 & n13201;
  assign new_n9127 = n2057 & n3085;
  assign new_n9128 = new_n9126 & new_n9127;
  assign new_n9129 = n3085 & n5586;
  assign new_n9130 = n124 & n2057;
  assign new_n9131 = n10805 & n13201;
  assign new_n9132 = ~new_n9130 & ~new_n9131;
  assign new_n9133 = new_n9130 & new_n9131;
  assign new_n9134 = ~new_n9132 & ~new_n9133;
  assign new_n9135 = new_n9129 & ~new_n9134;
  assign new_n9136 = ~new_n9129 & new_n9134;
  assign new_n9137 = ~new_n9135 & ~new_n9136;
  assign new_n9138 = new_n9128 & ~new_n9137;
  assign new_n9139 = n12263 & n13201;
  assign new_n9140 = new_n9129 & ~new_n9132;
  assign new_n9141 = ~new_n9133 & ~new_n9140;
  assign new_n9142 = ~new_n9139 & new_n9141;
  assign new_n9143 = new_n9139 & ~new_n9141;
  assign new_n9144 = ~new_n9142 & ~new_n9143;
  assign new_n9145 = n3085 & n4141;
  assign new_n9146 = n2057 & n10805;
  assign new_n9147 = n124 & n5586;
  assign new_n9148 = ~new_n9146 & ~new_n9147;
  assign new_n9149 = new_n9146 & new_n9147;
  assign new_n9150 = ~new_n9148 & ~new_n9149;
  assign new_n9151 = new_n9145 & ~new_n9150;
  assign new_n9152 = ~new_n9145 & new_n9150;
  assign new_n9153 = ~new_n9151 & ~new_n9152;
  assign new_n9154 = ~new_n9144 & new_n9153;
  assign new_n9155 = new_n9144 & ~new_n9153;
  assign new_n9156 = ~new_n9154 & ~new_n9155;
  assign new_n9157 = new_n9138 & new_n9156;
  assign new_n9158 = n353 & n13201;
  assign new_n9159 = n2057 & n12263;
  assign new_n9160 = new_n9145 & ~new_n9148;
  assign new_n9161 = ~new_n9149 & ~new_n9160;
  assign new_n9162 = ~new_n9159 & new_n9161;
  assign new_n9163 = new_n9159 & ~new_n9161;
  assign new_n9164 = ~new_n9162 & ~new_n9163;
  assign new_n9165 = n1364 & n3085;
  assign new_n9166 = n5586 & n10805;
  assign new_n9167 = n124 & n4141;
  assign new_n9168 = ~new_n9166 & ~new_n9167;
  assign new_n9169 = new_n9166 & new_n9167;
  assign new_n9170 = ~new_n9168 & ~new_n9169;
  assign new_n9171 = new_n9165 & ~new_n9170;
  assign new_n9172 = ~new_n9165 & new_n9170;
  assign new_n9173 = ~new_n9171 & ~new_n9172;
  assign new_n9174 = ~new_n9164 & new_n9173;
  assign new_n9175 = new_n9164 & ~new_n9173;
  assign new_n9176 = ~new_n9174 & ~new_n9175;
  assign new_n9177 = ~new_n9158 & ~new_n9176;
  assign new_n9178 = new_n9158 & new_n9176;
  assign new_n9179 = ~new_n9177 & ~new_n9178;
  assign new_n9180 = ~new_n9142 & ~new_n9153;
  assign new_n9181 = ~new_n9143 & ~new_n9180;
  assign new_n9182 = ~new_n9179 & new_n9181;
  assign new_n9183 = new_n9179 & ~new_n9181;
  assign new_n9184 = ~new_n9182 & ~new_n9183;
  assign new_n9185 = ~new_n9157 & ~new_n9184;
  assign new_n9186 = new_n9157 & new_n9184;
  assign new_n9187_1 = ~new_n9185 & ~new_n9186;
  assign new_n9188 = ~new_n9125 & ~new_n9187_1;
  assign new_n9189 = new_n9125 & new_n9187_1;
  assign new_n9190 = ~new_n9188 & ~new_n9189;
  assign new_n9191 = ~new_n9076 & ~new_n9094;
  assign new_n9192 = ~new_n9095 & ~new_n9191;
  assign new_n9193 = ~new_n9138 & ~new_n9156;
  assign new_n9194 = ~new_n9157 & ~new_n9193;
  assign new_n9195 = new_n9192 & new_n9194;
  assign new_n9196 = ~new_n9192 & ~new_n9194;
  assign new_n9197 = ~new_n9066 & new_n9075;
  assign new_n9198 = ~new_n9076 & ~new_n9197;
  assign new_n9199 = ~new_n9128 & new_n9137;
  assign new_n9200 = ~new_n9138 & ~new_n9199;
  assign new_n9201 = new_n9198 & new_n9200;
  assign new_n9202 = ~new_n9198 & ~new_n9200;
  assign new_n9203 = n5671 & n8506;
  assign new_n9204 = n3085 & n13201;
  assign new_n9205 = new_n9203 & new_n9204;
  assign new_n9206 = ~new_n9064 & ~new_n9065;
  assign new_n9207 = ~new_n9066 & ~new_n9206;
  assign new_n9208 = new_n9205 & new_n9207;
  assign new_n9209 = ~new_n9205 & ~new_n9207;
  assign new_n9210 = ~new_n9126 & ~new_n9127;
  assign new_n9211 = ~new_n9128 & ~new_n9210;
  assign new_n9212 = ~new_n9209 & new_n9211;
  assign new_n9213 = ~new_n9208 & ~new_n9212;
  assign new_n9214 = ~new_n9202 & ~new_n9213;
  assign new_n9215 = ~new_n9201 & ~new_n9214;
  assign new_n9216_1 = ~new_n9196 & ~new_n9215;
  assign new_n9217 = ~new_n9195 & ~new_n9216_1;
  assign new_n9218 = ~new_n9190 & new_n9217;
  assign new_n9219 = new_n9190 & ~new_n9217;
  assign new_n9220 = ~new_n9218 & ~new_n9219;
  assign new_n9221 = ~new_n9063 & ~new_n9220;
  assign new_n9222 = new_n9063 & new_n9220;
  assign new_n9223 = ~new_n9221 & ~new_n9222;
  assign new_n9224 = ~new_n9014 & ~new_n9032;
  assign new_n9225 = ~new_n9033 & ~new_n9224;
  assign new_n9226 = new_n9195 & ~new_n9215;
  assign new_n9227 = new_n9196 & new_n9215;
  assign new_n9228 = new_n9217 & ~new_n9227;
  assign new_n9229 = ~new_n9226 & ~new_n9228;
  assign new_n9230 = new_n9225 & ~new_n9229;
  assign new_n9231 = ~new_n9225 & new_n9229;
  assign new_n9232 = ~new_n9004 & new_n9013;
  assign new_n9233 = ~new_n9014 & ~new_n9232;
  assign new_n9234 = ~new_n9002 & ~new_n9003;
  assign new_n9235 = ~new_n9004 & ~new_n9234;
  assign new_n9236 = ~new_n9208 & ~new_n9209;
  assign new_n9237 = new_n9211 & ~new_n9236;
  assign new_n9238 = ~new_n9211 & new_n9236;
  assign new_n9239 = ~new_n9237 & ~new_n9238;
  assign new_n9240 = new_n9235 & ~new_n9239;
  assign new_n9241 = ~new_n9235 & new_n9239;
  assign new_n9242 = n411 & n5801;
  assign new_n9243 = ~new_n9203 & ~new_n9204;
  assign new_n9244 = ~new_n9205 & ~new_n9243;
  assign new_n9245 = new_n9242 & new_n9244;
  assign new_n9246 = ~new_n9241 & new_n9245;
  assign new_n9247 = ~new_n9240 & ~new_n9246;
  assign new_n9248 = ~new_n9233 & new_n9247;
  assign new_n9249 = new_n9233 & ~new_n9247;
  assign new_n9250 = ~new_n9201 & ~new_n9202;
  assign new_n9251 = new_n9213 & ~new_n9250;
  assign new_n9252 = ~new_n9213 & new_n9250;
  assign new_n9253 = ~new_n9251 & ~new_n9252;
  assign new_n9254 = ~new_n9249 & ~new_n9253;
  assign new_n9255 = ~new_n9248 & ~new_n9254;
  assign new_n9256 = ~new_n9231 & new_n9255;
  assign new_n9257 = ~new_n9230 & ~new_n9256;
  assign new_n9258 = ~new_n9223 & new_n9257;
  assign new_n9259 = new_n9223 & ~new_n9257;
  assign new_n9260 = ~new_n9258 & ~new_n9259;
  assign new_n9261 = n3006 & n5568;
  assign new_n9262 = n3006 & n11734;
  assign new_n9263 = n5568 & new_n9262;
  assign new_n9264 = ~n5568 & ~new_n9262;
  assign new_n9265 = ~new_n9263 & ~new_n9264;
  assign new_n9266 = n8308 & ~new_n9265;
  assign new_n9267 = ~n8308 & new_n9265;
  assign new_n9268 = ~new_n9266 & ~new_n9267;
  assign new_n9269 = new_n9261 & ~new_n9268;
  assign new_n9270 = n3006 & n12651;
  assign new_n9271 = n8308 & ~new_n9264;
  assign new_n9272 = ~new_n9263 & ~new_n9271;
  assign new_n9273 = ~new_n9270 & new_n9272;
  assign new_n9274 = new_n9270 & ~new_n9272;
  assign new_n9275 = ~new_n9273 & ~new_n9274;
  assign new_n9276 = n5568 & n11734;
  assign new_n9277 = n8308 & new_n9276;
  assign new_n9278 = ~n8308 & ~new_n9276;
  assign new_n9279 = ~new_n9277 & ~new_n9278;
  assign new_n9280 = n5214 & ~new_n9279;
  assign new_n9281 = n5214 & ~new_n9278;
  assign new_n9282 = new_n9279 & ~new_n9281;
  assign new_n9283 = ~new_n9280 & ~new_n9282;
  assign new_n9284 = ~new_n9275 & new_n9283;
  assign new_n9285 = new_n9275 & ~new_n9283;
  assign new_n9286 = ~new_n9284 & ~new_n9285;
  assign new_n9287 = new_n9269 & new_n9286;
  assign new_n9288 = n3006 & n7411;
  assign new_n9289 = n8308 & n11734;
  assign new_n9290 = n5214 & new_n9289;
  assign new_n9291 = ~n5214 & ~new_n9289;
  assign new_n9292 = n2771 & ~new_n9291;
  assign new_n9293 = ~new_n9290 & ~new_n9292;
  assign new_n9294 = ~n2771 & new_n9291;
  assign new_n9295 = new_n9293 & ~new_n9294;
  assign new_n9296 = n2771 & new_n9290;
  assign new_n9297 = ~new_n9295 & ~new_n9296;
  assign new_n9298 = n5568 & n12651;
  assign new_n9299 = ~new_n9277 & ~new_n9281;
  assign new_n9300_1 = ~new_n9298 & new_n9299;
  assign new_n9301 = new_n9298 & ~new_n9299;
  assign new_n9302 = ~new_n9300_1 & ~new_n9301;
  assign new_n9303 = new_n9297 & ~new_n9302;
  assign new_n9304 = ~new_n9297 & new_n9302;
  assign new_n9305 = ~new_n9303 & ~new_n9304;
  assign new_n9306 = ~new_n9288 & ~new_n9305;
  assign new_n9307 = new_n9288 & new_n9305;
  assign new_n9308 = ~new_n9306 & ~new_n9307;
  assign new_n9309 = ~new_n9273 & ~new_n9283;
  assign new_n9310 = ~new_n9274 & ~new_n9309;
  assign new_n9311 = ~new_n9308 & new_n9310;
  assign new_n9312 = new_n9308 & ~new_n9310;
  assign new_n9313 = ~new_n9311 & ~new_n9312;
  assign new_n9314 = new_n9287 & new_n9313;
  assign new_n9315 = ~new_n9287 & ~new_n9313;
  assign new_n9316 = ~new_n9314 & ~new_n9315;
  assign new_n9317 = ~new_n9269 & ~new_n9286;
  assign new_n9318 = ~new_n9287 & ~new_n9317;
  assign new_n9319 = ~new_n9230 & ~new_n9231;
  assign new_n9320 = ~new_n9255 & ~new_n9319;
  assign new_n9321 = new_n9255 & new_n9319;
  assign new_n9322 = ~new_n9320 & ~new_n9321;
  assign new_n9323 = new_n9318 & new_n9322;
  assign new_n9324 = ~new_n9318 & ~new_n9322;
  assign new_n9325 = ~new_n9261 & new_n9268;
  assign new_n9326 = ~new_n9269 & ~new_n9325;
  assign new_n9327 = ~new_n9248 & ~new_n9249;
  assign new_n9328 = new_n9253 & new_n9327;
  assign new_n9329_1 = ~new_n9253 & ~new_n9327;
  assign new_n9330 = ~new_n9328 & ~new_n9329_1;
  assign new_n9331 = new_n9326 & new_n9330;
  assign new_n9332 = ~new_n9326 & ~new_n9330;
  assign new_n9333 = ~n3006 & ~n5568;
  assign new_n9334 = ~new_n9242 & ~new_n9244;
  assign new_n9335 = ~new_n9245 & ~new_n9334;
  assign new_n9336 = new_n9261 & ~new_n9335;
  assign new_n9337 = ~new_n9333 & ~new_n9336;
  assign new_n9338 = ~new_n9240 & ~new_n9241;
  assign new_n9339 = ~new_n9245 & ~new_n9338;
  assign new_n9340 = new_n9245 & new_n9338;
  assign new_n9341 = ~new_n9339 & ~new_n9340;
  assign new_n9342 = new_n9337 & new_n9341;
  assign new_n9343 = n3006 & new_n9335;
  assign new_n9344 = ~n5568 & new_n9343;
  assign new_n9345 = ~new_n9342 & ~new_n9344;
  assign new_n9346 = ~new_n9332 & ~new_n9345;
  assign new_n9347 = ~new_n9331 & ~new_n9346;
  assign new_n9348 = ~new_n9324 & ~new_n9347;
  assign new_n9349 = ~new_n9323 & ~new_n9348;
  assign new_n9350 = ~new_n9316 & new_n9349;
  assign new_n9351 = new_n9316 & ~new_n9349;
  assign new_n9352 = ~new_n9350 & ~new_n9351;
  assign new_n9353_1 = ~new_n9260 & new_n9352;
  assign new_n9354 = new_n9260 & ~new_n9352;
  assign n3323 = new_n9353_1 | new_n9354;
  assign new_n9356 = ~new_n8673 & ~new_n8674;
  assign new_n9357 = ~new_n8678 & ~new_n9356;
  assign new_n9358 = new_n8678 & new_n9356;
  assign n3362 = new_n9357 | new_n9358;
  assign new_n9360 = ~new_n1358 & ~new_n1359;
  assign new_n9361 = new_n1393 & ~new_n9360;
  assign new_n9362 = ~new_n1393 & new_n9360;
  assign n3748 = new_n9361 | new_n9362;
  assign new_n9364 = ~new_n3497 & ~new_n3498;
  assign new_n9365 = new_n3518 & ~new_n9364;
  assign new_n9366 = ~new_n3518 & new_n9364;
  assign n3790 = ~new_n9365 & ~new_n9366;
  assign new_n9368 = ~new_n1374 & ~new_n1375;
  assign new_n9369 = new_n1389 & ~new_n9368;
  assign new_n9370 = ~new_n1389 & new_n9368;
  assign n3946 = new_n9369 | new_n9370;
  assign new_n9372 = ~new_n4871 & ~new_n4872;
  assign new_n9373 = new_n4906 & ~new_n9372;
  assign new_n9374 = ~new_n4906 & new_n9372;
  assign n4059 = ~new_n9373 & ~new_n9374;
  assign new_n9376 = ~new_n7810 & ~new_n7811;
  assign new_n9377 = new_n7821 & new_n9376;
  assign new_n9378 = ~new_n7821 & ~new_n9376;
  assign n4202 = ~new_n9377 & ~new_n9378;
  assign new_n9380 = ~new_n7534 & ~new_n7537;
  assign new_n9381 = n1757 & n7113;
  assign new_n9382 = n499 & n2482;
  assign new_n9383 = n1302 & n10113;
  assign new_n9384 = ~new_n9382 & ~new_n9383;
  assign new_n9385 = new_n9382 & new_n9383;
  assign new_n9386 = ~new_n9384 & ~new_n9385;
  assign new_n9387 = ~new_n9381 & ~new_n9386;
  assign new_n9388 = new_n9381 & new_n9386;
  assign new_n9389 = ~new_n9387 & ~new_n9388;
  assign new_n9390 = ~new_n7516 & new_n7519;
  assign new_n9391 = ~new_n7515 & ~new_n9390;
  assign new_n9392 = ~new_n9389 & ~new_n9391;
  assign new_n9393 = new_n9389 & new_n9391;
  assign new_n9394 = ~new_n9392 & ~new_n9393;
  assign new_n9395 = n1982 & n10451;
  assign new_n9396 = n9093 & n11488;
  assign new_n9397 = n10594 & n11030;
  assign new_n9398 = ~new_n9396 & ~new_n9397;
  assign new_n9399 = new_n9396 & new_n9397;
  assign new_n9400 = ~new_n9398 & ~new_n9399;
  assign new_n9401 = new_n9395 & ~new_n9400;
  assign new_n9402 = ~new_n9395 & new_n9400;
  assign new_n9403 = ~new_n9401 & ~new_n9402;
  assign new_n9404 = n3409 & n10416;
  assign new_n9405 = new_n7513 & new_n9404;
  assign new_n9406 = ~new_n7513 & ~new_n9404;
  assign new_n9407 = ~new_n9405 & ~new_n9406;
  assign new_n9408 = ~new_n9403 & new_n9407;
  assign new_n9409 = new_n9403 & ~new_n9407;
  assign new_n9410 = ~new_n9408 & ~new_n9409;
  assign new_n9411 = new_n9394 & new_n9410;
  assign new_n9412 = ~new_n9394 & ~new_n9410;
  assign new_n9413 = ~new_n9411 & ~new_n9412;
  assign new_n9414 = ~new_n7523 & new_n7527;
  assign new_n9415 = ~new_n7507 & ~new_n9414;
  assign new_n9416 = ~new_n7524 & new_n9415;
  assign new_n9417 = new_n7507 & new_n9414;
  assign new_n9418 = ~new_n9416 & ~new_n9417;
  assign new_n9419 = ~new_n9413 & new_n9418;
  assign new_n9420 = new_n9413 & ~new_n9418;
  assign new_n9421 = ~new_n9419 & ~new_n9420;
  assign new_n9422 = new_n7531 & ~new_n9421;
  assign new_n9423 = ~new_n7531 & new_n9421;
  assign new_n9424 = ~new_n9422 & ~new_n9423;
  assign new_n9425 = ~new_n9380 & new_n9424;
  assign new_n9426 = new_n9380 & ~new_n9424;
  assign new_n9427 = ~new_n9425 & ~new_n9426;
  assign new_n9428 = ~new_n7864 & ~new_n7868;
  assign new_n9429 = n4382 & n8468;
  assign new_n9430 = n6818 & n11236;
  assign new_n9431 = n1084 & n8228;
  assign new_n9432 = ~new_n9430 & ~new_n9431;
  assign new_n9433 = new_n9430 & new_n9431;
  assign new_n9434 = ~new_n9432 & ~new_n9433;
  assign new_n9435 = new_n9429 & ~new_n9434;
  assign new_n9436 = ~new_n9429 & new_n9434;
  assign new_n9437 = ~new_n9435 & ~new_n9436;
  assign new_n9438 = ~new_n7844 & new_n7847;
  assign new_n9439 = ~new_n7843 & ~new_n9438;
  assign new_n9440 = new_n9437 & ~new_n9439;
  assign new_n9441 = n3130 & n11109;
  assign new_n9442 = new_n7841 & new_n9441;
  assign new_n9443 = ~new_n7841 & ~new_n9441;
  assign new_n9444 = ~new_n9442 & ~new_n9443;
  assign new_n9445 = n5320 & n5962;
  assign new_n9446 = n103 & n6085;
  assign new_n9447 = n9732 & n9906;
  assign new_n9448 = ~new_n9446 & ~new_n9447;
  assign new_n9449 = new_n9446 & new_n9447;
  assign new_n9450 = ~new_n9448 & ~new_n9449;
  assign new_n9451 = new_n9445 & ~new_n9450;
  assign new_n9452 = ~new_n9445 & new_n9450;
  assign new_n9453 = ~new_n9451 & ~new_n9452;
  assign new_n9454 = new_n9444 & new_n9453;
  assign new_n9455 = ~new_n9444 & ~new_n9453;
  assign new_n9456 = ~new_n9454 & ~new_n9455;
  assign new_n9457 = new_n9440 & new_n9456;
  assign new_n9458 = ~new_n9437 & new_n9439;
  assign new_n9459 = new_n9456 & ~new_n9458;
  assign new_n9460 = ~new_n9440 & ~new_n9459;
  assign new_n9461 = ~new_n9456 & new_n9458;
  assign new_n9462 = new_n9460 & ~new_n9461;
  assign new_n9463 = ~new_n9457 & ~new_n9462;
  assign new_n9464 = ~new_n7851 & ~new_n7855;
  assign new_n9465 = new_n7835 & new_n9464;
  assign new_n9466 = ~new_n7835 & ~new_n9464;
  assign new_n9467 = ~new_n7852 & new_n9466;
  assign new_n9468 = ~new_n9465 & ~new_n9467;
  assign new_n9469 = ~new_n9463 & ~new_n9468;
  assign new_n9470 = new_n9463 & new_n9468;
  assign new_n9471 = ~new_n9469 & ~new_n9470;
  assign new_n9472 = new_n7861 & new_n9471;
  assign new_n9473 = ~new_n7861 & ~new_n9471;
  assign new_n9474 = ~new_n9472 & ~new_n9473;
  assign new_n9475_1 = ~new_n9428 & new_n9474;
  assign new_n9476 = new_n9428 & ~new_n9474;
  assign new_n9477 = ~new_n9475_1 & ~new_n9476;
  assign new_n9478 = ~new_n7953 & ~new_n7958;
  assign new_n9479 = ~new_n7946 & ~new_n7949;
  assign new_n9480 = ~new_n7933 & ~new_n7937;
  assign new_n9481 = new_n7917 & new_n9480;
  assign new_n9482 = ~new_n7917 & ~new_n9480;
  assign new_n9483 = ~new_n7934 & new_n9482;
  assign new_n9484 = ~new_n9481 & ~new_n9483;
  assign new_n9485 = n1198 & n1912;
  assign new_n9486 = n9353 & n11574;
  assign new_n9487 = n6333 & n9300;
  assign new_n9488 = ~new_n9486 & ~new_n9487;
  assign new_n9489 = new_n9486 & new_n9487;
  assign new_n9490 = ~new_n9488 & ~new_n9489;
  assign new_n9491 = new_n9485 & ~new_n9490;
  assign new_n9492 = ~new_n9485 & new_n9490;
  assign new_n9493 = ~new_n9491 & ~new_n9492;
  assign new_n9494 = ~new_n7925 & new_n7929;
  assign new_n9495 = ~new_n7926 & ~new_n9494;
  assign new_n9496 = new_n9493 & ~new_n9495;
  assign new_n9497 = n2498 & n12750;
  assign new_n9498 = new_n7923 & new_n9497;
  assign new_n9499 = ~new_n7923 & ~new_n9497;
  assign new_n9500 = ~new_n9498 & ~new_n9499;
  assign new_n9501 = n5758 & n11058;
  assign new_n9502 = n761 & n1007;
  assign new_n9503 = n5969 & n9620;
  assign new_n9504 = ~new_n9502 & ~new_n9503;
  assign new_n9505 = new_n9502 & new_n9503;
  assign new_n9506 = ~new_n9504 & ~new_n9505;
  assign new_n9507 = new_n9501 & ~new_n9506;
  assign new_n9508 = ~new_n9501 & new_n9506;
  assign new_n9509 = ~new_n9507 & ~new_n9508;
  assign new_n9510 = new_n9500 & new_n9509;
  assign new_n9511 = ~new_n9500 & ~new_n9509;
  assign new_n9512 = ~new_n9510 & ~new_n9511;
  assign new_n9513 = new_n9496 & new_n9512;
  assign new_n9514 = ~new_n9493 & new_n9495;
  assign new_n9515 = ~new_n9512 & new_n9514;
  assign new_n9516 = ~new_n9496 & ~new_n9512;
  assign new_n9517 = ~new_n9514 & ~new_n9516;
  assign new_n9518 = ~new_n9515 & ~new_n9517;
  assign new_n9519 = ~new_n9513 & ~new_n9518;
  assign new_n9520 = ~new_n9484 & new_n9519;
  assign new_n9521 = new_n9484 & ~new_n9519;
  assign new_n9522 = ~new_n9520 & ~new_n9521;
  assign new_n9523 = new_n7943 & ~new_n9522;
  assign new_n9524 = ~new_n7943 & new_n9522;
  assign new_n9525 = ~new_n9523 & ~new_n9524;
  assign new_n9526 = ~new_n9479 & new_n9525;
  assign new_n9527 = new_n9479 & ~new_n9525;
  assign new_n9528_1 = ~new_n9526 & ~new_n9527;
  assign new_n9529 = ~new_n7894 & new_n7898;
  assign new_n9530 = ~new_n7879 & ~new_n9529;
  assign new_n9531_1 = ~new_n7895 & new_n9530;
  assign new_n9532 = new_n7879 & new_n9529;
  assign new_n9533 = ~new_n9531_1 & ~new_n9532;
  assign new_n9534 = n2339 & n5684;
  assign new_n9535 = n1307 & n4964;
  assign new_n9536 = ~new_n9534 & ~new_n9535;
  assign new_n9537 = new_n9534 & new_n9535;
  assign new_n9538 = ~new_n9536 & ~new_n9537;
  assign new_n9539 = ~new_n7886 & ~new_n7890;
  assign new_n9540 = ~new_n7887 & ~new_n9539;
  assign new_n9541 = new_n9538 & ~new_n9540;
  assign new_n9542 = ~new_n9538 & new_n9540;
  assign new_n9543 = ~new_n9541 & ~new_n9542;
  assign new_n9544 = ~n12482 & new_n7885;
  assign new_n9545 = n10770 & n12482;
  assign new_n9546 = ~new_n7885 & new_n9545;
  assign new_n9547 = ~new_n9544 & ~new_n9546;
  assign new_n9548 = n9570 & n10522;
  assign new_n9549 = new_n7883 & new_n9548;
  assign new_n9550 = ~new_n7883 & ~new_n9548;
  assign new_n9551 = ~new_n9549 & ~new_n9550;
  assign new_n9552 = new_n9547 & ~new_n9551;
  assign new_n9553 = ~new_n9547 & new_n9551;
  assign new_n9554 = ~new_n9552 & ~new_n9553;
  assign new_n9555 = new_n9543 & new_n9554;
  assign new_n9556 = ~new_n9543 & ~new_n9554;
  assign new_n9557 = ~new_n9555 & ~new_n9556;
  assign new_n9558 = new_n9533 & new_n9557;
  assign new_n9559 = ~new_n9533 & ~new_n9557;
  assign new_n9560 = ~new_n9558 & ~new_n9559;
  assign new_n9561 = ~new_n7904 & ~new_n9560;
  assign new_n9562 = new_n7904 & new_n9560;
  assign new_n9563 = ~new_n9561 & ~new_n9562;
  assign new_n9564 = ~new_n7907 & ~new_n7910;
  assign new_n9565 = ~new_n9563 & new_n9564;
  assign new_n9566 = new_n9563 & ~new_n9564;
  assign new_n9567 = ~new_n9565 & ~new_n9566;
  assign new_n9568 = ~new_n9528_1 & ~new_n9567;
  assign new_n9569 = new_n9528_1 & new_n9567;
  assign new_n9570_1 = ~new_n9568 & ~new_n9569;
  assign new_n9571 = ~new_n9478 & ~new_n9570_1;
  assign new_n9572 = new_n9478 & new_n9570_1;
  assign new_n9573 = ~new_n9571 & ~new_n9572;
  assign new_n9574 = ~new_n9477 & ~new_n9573;
  assign new_n9575 = new_n9477 & new_n9573;
  assign new_n9576 = ~new_n9574 & ~new_n9575;
  assign new_n9577 = ~new_n7872 & ~new_n7960;
  assign new_n9578 = ~new_n7873 & ~new_n9577;
  assign new_n9579 = ~new_n9576 & new_n9578;
  assign new_n9580 = new_n9576 & ~new_n9578;
  assign new_n9581 = ~new_n9579 & ~new_n9580;
  assign new_n9582 = new_n9427 & new_n9581;
  assign new_n9583 = ~new_n9427 & ~new_n9581;
  assign new_n9584 = ~new_n7828 & ~new_n7965;
  assign new_n9585 = ~new_n9583 & new_n9584;
  assign new_n9586 = ~new_n9582 & ~new_n9585;
  assign new_n9587 = new_n9537 & new_n9547;
  assign new_n9588 = ~new_n9537 & ~new_n9547;
  assign new_n9589 = ~new_n9587 & ~new_n9588;
  assign new_n9590 = new_n9485 & ~new_n9488;
  assign new_n9591_1 = ~new_n9489 & ~new_n9590;
  assign new_n9592 = n8820 & n10451;
  assign new_n9593 = n9570 & n10770;
  assign new_n9594 = n6843 & n8940;
  assign new_n9595 = ~new_n9593 & new_n9594;
  assign new_n9596 = new_n9593 & ~new_n9594;
  assign new_n9597 = ~new_n9595 & ~new_n9596;
  assign new_n9598 = ~new_n9592 & new_n9597;
  assign new_n9599 = new_n9592 & ~new_n9597;
  assign new_n9600 = ~new_n9598 & ~new_n9599;
  assign new_n9601 = new_n9591_1 & ~new_n9600;
  assign new_n9602 = ~new_n9591_1 & new_n9600;
  assign new_n9603 = ~new_n9601 & ~new_n9602;
  assign new_n9604 = n6333 & n11574;
  assign new_n9605 = n1912 & n9300;
  assign new_n9606 = new_n9604 & ~new_n9605;
  assign new_n9607 = ~new_n9604 & new_n9605;
  assign new_n9608 = ~new_n9606 & ~new_n9607;
  assign new_n9609 = n1982 & n9093;
  assign new_n9610 = n2482 & n11111;
  assign new_n9611 = ~new_n9609 & new_n9610;
  assign new_n9612 = new_n9609 & ~new_n9610;
  assign new_n9613 = ~new_n9611 & ~new_n9612;
  assign new_n9614 = ~new_n9608 & new_n9613;
  assign new_n9615 = new_n9608 & ~new_n9613;
  assign new_n9616 = ~new_n9614 & ~new_n9615;
  assign new_n9617 = n1198 & n12750;
  assign new_n9618 = new_n9501 & ~new_n9504;
  assign new_n9619 = ~new_n9505 & ~new_n9618;
  assign new_n9620_1 = new_n9617 & new_n9619;
  assign new_n9621 = ~new_n9617 & ~new_n9619;
  assign new_n9622 = ~new_n9620_1 & ~new_n9621;
  assign new_n9623 = new_n9616 & new_n9622;
  assign new_n9624 = ~new_n9616 & ~new_n9622;
  assign new_n9625 = ~new_n9623 & ~new_n9624;
  assign new_n9626 = new_n9603 & ~new_n9625;
  assign new_n9627 = ~new_n9603 & new_n9625;
  assign new_n9628 = ~new_n9626 & ~new_n9627;
  assign new_n9629 = ~new_n9517 & new_n9628;
  assign new_n9630 = new_n9517 & ~new_n9628;
  assign new_n9631 = ~new_n9629 & ~new_n9630;
  assign new_n9632 = ~new_n9589 & new_n9631;
  assign new_n9633 = new_n9589 & ~new_n9631;
  assign new_n9634 = ~new_n9632 & ~new_n9633;
  assign new_n9635 = new_n9413 & ~new_n9416;
  assign new_n9636 = ~new_n9417 & ~new_n9635;
  assign new_n9637 = n1307 & n5684;
  assign new_n9638 = n2339 & n10522;
  assign new_n9639 = ~new_n9637 & new_n9638;
  assign new_n9640 = new_n9637 & ~new_n9638;
  assign new_n9641 = ~new_n9639 & ~new_n9640;
  assign new_n9642 = new_n9636 & ~new_n9641;
  assign new_n9643 = ~new_n9636 & new_n9641;
  assign new_n9644 = ~new_n9642 & ~new_n9643;
  assign new_n9645 = ~new_n9541 & ~new_n9554;
  assign new_n9646 = ~new_n9542 & ~new_n9645;
  assign new_n9647 = new_n9644 & new_n9646;
  assign new_n9648 = ~new_n9644 & ~new_n9646;
  assign new_n9649 = ~new_n9647 & ~new_n9648;
  assign new_n9650 = ~new_n9634 & new_n9649;
  assign new_n9651 = new_n9634 & ~new_n9649;
  assign new_n9652 = ~new_n9650 & ~new_n9651;
  assign new_n9653 = ~new_n9531_1 & new_n9557;
  assign new_n9654 = ~new_n9532 & ~new_n9653;
  assign new_n9655 = n12482 & ~new_n7884;
  assign new_n9656 = ~new_n7883 & ~new_n9655;
  assign new_n9657 = ~new_n9654 & new_n9656;
  assign new_n9658 = new_n9654 & ~new_n9656;
  assign new_n9659 = ~new_n9657 & ~new_n9658;
  assign new_n9660 = ~new_n9652 & new_n9659;
  assign new_n9661 = new_n9652 & ~new_n9659;
  assign new_n9662 = ~new_n9660 & ~new_n9661;
  assign new_n9663 = ~new_n9422 & ~new_n9425;
  assign new_n9664 = ~new_n9562 & ~new_n9566;
  assign new_n9665 = new_n9547 & ~new_n9549;
  assign new_n9666 = ~new_n9550 & ~new_n9665;
  assign new_n9667 = ~new_n9664 & ~new_n9666;
  assign new_n9668 = new_n9664 & new_n9666;
  assign new_n9669_1 = ~new_n9667 & ~new_n9668;
  assign new_n9670 = new_n9663 & new_n9669_1;
  assign new_n9671 = ~new_n9663 & ~new_n9669_1;
  assign new_n9672 = ~new_n9670 & ~new_n9671;
  assign new_n9673 = new_n9662 & new_n9672;
  assign new_n9674 = ~new_n9662 & ~new_n9672;
  assign new_n9675 = ~new_n9673 & ~new_n9674;
  assign new_n9676 = new_n9586 & new_n9675;
  assign new_n9677 = ~new_n9586 & ~new_n9675;
  assign new_n9678 = ~new_n9676 & ~new_n9677;
  assign new_n9679 = new_n9463 & ~new_n9467;
  assign new_n9680 = ~new_n9465 & ~new_n9679;
  assign new_n9681 = n1007 & n5758;
  assign new_n9682 = n8859 & n9353;
  assign new_n9683 = ~new_n9681 & ~new_n9682;
  assign new_n9684 = new_n9681 & new_n9682;
  assign new_n9685 = ~new_n9683 & ~new_n9684;
  assign new_n9686 = n761 & n5969;
  assign new_n9687 = n2498 & n9620;
  assign new_n9688 = new_n9686 & ~new_n9687;
  assign new_n9689 = ~new_n9686 & new_n9687;
  assign new_n9690 = ~new_n9688 & ~new_n9689;
  assign new_n9691 = ~new_n9685 & ~new_n9690;
  assign new_n9692 = new_n9685 & new_n9690;
  assign new_n9693 = ~new_n9691 & ~new_n9692;
  assign new_n9694 = ~new_n9680 & ~new_n9693;
  assign new_n9695 = new_n9680 & new_n9693;
  assign new_n9696 = ~new_n9694 & ~new_n9695;
  assign new_n9697 = ~new_n9574 & ~new_n9578;
  assign new_n9698 = ~new_n9575 & ~new_n9697;
  assign new_n9699 = ~new_n9696 & new_n9698;
  assign new_n9700 = new_n9696 & ~new_n9698;
  assign new_n9701 = ~new_n9699 & ~new_n9700;
  assign new_n9702 = ~new_n9483 & new_n9519;
  assign new_n9703 = ~new_n9481 & ~new_n9702;
  assign new_n9704 = ~new_n9442 & new_n9453;
  assign new_n9705 = ~new_n9443 & ~new_n9704;
  assign new_n9706 = n9732 & n11109;
  assign new_n9707 = n3130 & n8468;
  assign new_n9708 = ~new_n9706 & ~new_n9707;
  assign new_n9709 = new_n9706 & new_n9707;
  assign new_n9710 = ~new_n9708 & ~new_n9709;
  assign new_n9711 = n1084 & n11236;
  assign new_n9712 = n4382 & n6818;
  assign new_n9713 = new_n9711 & ~new_n9712;
  assign new_n9714 = ~new_n9711 & new_n9712;
  assign new_n9715 = ~new_n9713 & ~new_n9714;
  assign new_n9716 = ~new_n9710 & ~new_n9715;
  assign new_n9717 = new_n9710 & new_n9715;
  assign new_n9718 = ~new_n9716 & ~new_n9717;
  assign new_n9719 = new_n9429 & ~new_n9432;
  assign new_n9720 = ~new_n9433 & ~new_n9719;
  assign new_n9721 = new_n9445 & ~new_n9448;
  assign new_n9722 = ~new_n9449 & ~new_n9721;
  assign new_n9723 = ~new_n9720 & new_n9722;
  assign new_n9724 = new_n9720 & ~new_n9722;
  assign new_n9725 = ~new_n9723 & ~new_n9724;
  assign new_n9726 = new_n9718 & new_n9725;
  assign new_n9727 = ~new_n9718 & ~new_n9725;
  assign new_n9728 = ~new_n9726 & ~new_n9727;
  assign new_n9729 = ~new_n9705 & new_n9728;
  assign new_n9730 = new_n9705 & ~new_n9728;
  assign new_n9731 = ~new_n9729 & ~new_n9730;
  assign new_n9732_1 = new_n9460 & ~new_n9731;
  assign new_n9733 = ~new_n9460 & new_n9731;
  assign new_n9734 = ~new_n9732_1 & ~new_n9733;
  assign new_n9735 = new_n9703 & new_n9734;
  assign new_n9736 = ~new_n9703 & ~new_n9734;
  assign new_n9737 = ~new_n9735 & ~new_n9736;
  assign new_n9738 = n11058 & n12352;
  assign new_n9739 = ~new_n9523 & ~new_n9526;
  assign new_n9740 = new_n9738 & new_n9739;
  assign new_n9741 = ~new_n9738 & ~new_n9739;
  assign new_n9742 = ~new_n9740 & ~new_n9741;
  assign new_n9743 = new_n9737 & ~new_n9742;
  assign new_n9744 = ~new_n9737 & new_n9742;
  assign new_n9745 = ~new_n9743 & ~new_n9744;
  assign new_n9746 = ~new_n9499 & ~new_n9509;
  assign new_n9747_1 = ~new_n9498 & ~new_n9746;
  assign new_n9748 = new_n9478 & ~new_n9568;
  assign new_n9749 = ~new_n9569 & ~new_n9748;
  assign new_n9750 = new_n9747_1 & ~new_n9749;
  assign new_n9751 = ~new_n9747_1 & new_n9749;
  assign new_n9752 = ~new_n9750 & ~new_n9751;
  assign new_n9753 = ~new_n9745 & ~new_n9752;
  assign new_n9754 = new_n9745 & new_n9752;
  assign new_n9755 = ~new_n9753 & ~new_n9754;
  assign new_n9756 = ~new_n9472 & ~new_n9475_1;
  assign new_n9757 = new_n9381 & ~new_n9384;
  assign new_n9758 = ~new_n9385 & ~new_n9757;
  assign new_n9759 = new_n9403 & ~new_n9405;
  assign new_n9760 = ~new_n9406 & ~new_n9759;
  assign new_n9761 = new_n9395 & ~new_n9398;
  assign new_n9762 = ~new_n9399 & ~new_n9761;
  assign new_n9763 = n3409 & n11030;
  assign new_n9764 = n1302 & n1757;
  assign new_n9765 = new_n9763 & new_n9764;
  assign new_n9766 = ~new_n9763 & ~new_n9764;
  assign new_n9767 = ~new_n9765 & ~new_n9766;
  assign new_n9768 = new_n9762 & ~new_n9767;
  assign new_n9769 = ~new_n9762 & new_n9767;
  assign new_n9770 = ~new_n9768 & ~new_n9769;
  assign new_n9771 = ~new_n9760 & ~new_n9770;
  assign new_n9772 = new_n9760 & new_n9770;
  assign new_n9773 = ~new_n9771 & ~new_n9772;
  assign new_n9774 = ~new_n9393 & ~new_n9410;
  assign new_n9775 = ~new_n9392 & ~new_n9774;
  assign new_n9776 = n499 & n10113;
  assign new_n9777 = n10594 & n11488;
  assign new_n9778 = n7113 & n10416;
  assign new_n9779 = ~new_n9777 & new_n9778;
  assign new_n9780 = new_n9777 & ~new_n9778;
  assign new_n9781 = ~new_n9779 & ~new_n9780;
  assign new_n9782 = ~new_n9776 & new_n9781;
  assign new_n9783 = new_n9776 & ~new_n9781;
  assign new_n9784 = ~new_n9782 & ~new_n9783;
  assign new_n9785 = new_n9775 & ~new_n9784;
  assign new_n9786 = ~new_n9775 & new_n9784;
  assign new_n9787 = ~new_n9785 & ~new_n9786;
  assign new_n9788 = new_n9773 & ~new_n9787;
  assign new_n9789 = ~new_n9773 & new_n9787;
  assign new_n9790 = ~new_n9788 & ~new_n9789;
  assign new_n9791 = ~new_n9758 & new_n9790;
  assign new_n9792 = new_n9758 & ~new_n9790;
  assign new_n9793 = ~new_n9791 & ~new_n9792;
  assign new_n9794 = n4743 & n5962;
  assign new_n9795 = n1392 & n8228;
  assign new_n9796 = ~new_n9794 & ~new_n9795;
  assign new_n9797 = new_n9794 & new_n9795;
  assign new_n9798 = ~new_n9796 & ~new_n9797;
  assign new_n9799 = n103 & n9906;
  assign new_n9800 = n5320 & n6085;
  assign new_n9801 = new_n9799 & ~new_n9800;
  assign new_n9802 = ~new_n9799 & new_n9800;
  assign new_n9803 = ~new_n9801 & ~new_n9802;
  assign new_n9804 = ~new_n9798 & ~new_n9803;
  assign new_n9805 = new_n9798 & new_n9803;
  assign new_n9806 = ~new_n9804 & ~new_n9805;
  assign new_n9807 = ~new_n9793 & new_n9806;
  assign new_n9808 = new_n9793 & ~new_n9806;
  assign new_n9809 = ~new_n9807 & ~new_n9808;
  assign new_n9810 = new_n9756 & ~new_n9809;
  assign new_n9811 = ~new_n9756 & new_n9809;
  assign new_n9812 = ~new_n9810 & ~new_n9811;
  assign new_n9813 = new_n9755 & new_n9812;
  assign new_n9814 = ~new_n9755 & ~new_n9812;
  assign new_n9815 = ~new_n9813 & ~new_n9814;
  assign new_n9816 = ~new_n9701 & new_n9815;
  assign new_n9817 = new_n9701 & ~new_n9815;
  assign new_n9818 = ~new_n9816 & ~new_n9817;
  assign new_n9819 = new_n9678 & ~new_n9818;
  assign new_n9820 = ~new_n9678 & new_n9818;
  assign n4553 = ~new_n9819 & ~new_n9820;
  assign new_n9822 = ~new_n3772 & ~new_n3988;
  assign new_n9823 = ~new_n3989 & ~new_n9822;
  assign new_n9824 = ~new_n3775 & ~new_n3812;
  assign new_n9825 = ~new_n3776 & ~new_n9824;
  assign new_n9826 = ~new_n3878 & ~new_n3879;
  assign new_n9827 = ~new_n3881 & ~new_n9826;
  assign new_n9828 = n4470 & n7061;
  assign new_n9829 = n3006 & n3641;
  assign new_n9830 = ~new_n9828 & new_n9829;
  assign new_n9831 = new_n9828 & ~new_n9829;
  assign new_n9832 = ~new_n9830 & ~new_n9831;
  assign new_n9833 = ~new_n9827 & new_n9832;
  assign new_n9834 = new_n9827 & ~new_n9832;
  assign new_n9835 = ~new_n9833 & ~new_n9834;
  assign new_n9836 = new_n9825 & ~new_n9835;
  assign new_n9837 = ~new_n9825 & new_n9835;
  assign new_n9838 = ~new_n9836 & ~new_n9837;
  assign new_n9839 = ~new_n3890 & new_n3901;
  assign new_n9840 = ~new_n3891 & ~new_n9839;
  assign new_n9841 = n4114 & n11665;
  assign new_n9842 = ~n4114 & ~n11665;
  assign new_n9843 = n3112 & ~new_n9842;
  assign new_n9844 = ~new_n9841 & new_n9843;
  assign new_n9845 = new_n3893 & ~new_n3896;
  assign new_n9846_1 = ~new_n3897 & ~new_n9845;
  assign new_n9847 = new_n9844 & ~new_n9846_1;
  assign new_n9848 = ~new_n9844 & new_n9846_1;
  assign new_n9849 = ~new_n9847 & ~new_n9848;
  assign new_n9850 = ~new_n9840 & new_n9849;
  assign new_n9851 = new_n9840 & ~new_n9849;
  assign new_n9852 = ~new_n9850 & ~new_n9851;
  assign new_n9853 = new_n3908 & new_n9852;
  assign new_n9854 = ~new_n3908 & ~new_n9852;
  assign new_n9855 = ~new_n9853 & ~new_n9854;
  assign new_n9856 = ~new_n9838 & new_n9855;
  assign new_n9857 = new_n9838 & ~new_n9855;
  assign new_n9858 = ~new_n9856 & ~new_n9857;
  assign new_n9859 = ~new_n9823 & new_n9858;
  assign new_n9860 = new_n9823 & ~new_n9858;
  assign new_n9861 = ~new_n9859 & ~new_n9860;
  assign new_n9862 = ~new_n3817 & ~new_n3821;
  assign new_n9863 = ~new_n1953 & ~new_n3983;
  assign new_n9864 = ~new_n3982 & ~new_n9863;
  assign new_n9865 = ~new_n3867 & ~new_n3870;
  assign new_n9866_1 = new_n3778 & ~new_n3781;
  assign new_n9867 = ~new_n3782 & ~new_n9866_1;
  assign new_n9868 = ~new_n3792 & ~new_n3802;
  assign new_n9869 = ~new_n3791 & ~new_n9868;
  assign new_n9870 = n2771 & n12306;
  assign new_n9871 = n4748 & n5214;
  assign new_n9872_1 = new_n9870 & ~new_n9871;
  assign new_n9873 = ~new_n9870 & new_n9871;
  assign new_n9874 = ~new_n9872_1 & ~new_n9873;
  assign new_n9875 = n1231 & n5568;
  assign new_n9876 = n8308 & n9187;
  assign new_n9877 = ~new_n9875 & new_n9876;
  assign new_n9878 = new_n9875 & ~new_n9876;
  assign new_n9879 = ~new_n9877 & ~new_n9878;
  assign new_n9880 = ~new_n9874 & new_n9879;
  assign new_n9881 = new_n9874 & ~new_n9879;
  assign new_n9882 = ~new_n9880 & ~new_n9881;
  assign new_n9883 = ~new_n3794 & ~new_n3798;
  assign new_n9884 = ~new_n3797 & ~new_n9883;
  assign new_n9885 = n4006 & n6168;
  assign new_n9886 = n2758 & n11411;
  assign new_n9887_1 = ~new_n9885 & ~new_n9886;
  assign new_n9888 = new_n9885 & new_n9886;
  assign new_n9889 = ~new_n9887_1 & ~new_n9888;
  assign new_n9890 = new_n9884 & new_n9889;
  assign new_n9891 = ~new_n9884 & ~new_n9889;
  assign new_n9892 = ~new_n9890 & ~new_n9891;
  assign new_n9893 = new_n9882 & new_n9892;
  assign new_n9894 = ~new_n9882 & ~new_n9892;
  assign new_n9895 = ~new_n9893 & ~new_n9894;
  assign new_n9896 = ~new_n9869 & new_n9895;
  assign new_n9897 = new_n9869 & ~new_n9895;
  assign new_n9898 = ~new_n9896 & ~new_n9897;
  assign new_n9899 = ~new_n9867 & new_n9898;
  assign new_n9900 = new_n9867 & ~new_n9898;
  assign new_n9901 = ~new_n9899 & ~new_n9900;
  assign new_n9902 = ~new_n3809 & new_n9901;
  assign new_n9903 = new_n3809 & ~new_n9901;
  assign new_n9904 = ~new_n9902 & ~new_n9903;
  assign new_n9905 = new_n9865 & ~new_n9904;
  assign new_n9906_1 = ~new_n9865 & new_n9904;
  assign new_n9907 = ~new_n9905 & ~new_n9906_1;
  assign new_n9908 = new_n9864 & ~new_n9907;
  assign new_n9909 = ~new_n9864 & new_n9907;
  assign new_n9910 = ~new_n9908 & ~new_n9909;
  assign new_n9911 = ~new_n3966 & ~new_n3970;
  assign new_n9912 = ~new_n3924 & ~new_n3961;
  assign new_n9913 = ~new_n3925 & ~new_n9912;
  assign new_n9914 = new_n3824 & ~new_n3827;
  assign new_n9915_1 = ~new_n3828 & ~new_n9914;
  assign new_n9916 = n6409 & n10063;
  assign new_n9917 = n10874 & n13201;
  assign new_n9918 = ~new_n9916 & ~new_n9917;
  assign new_n9919 = new_n9916 & new_n9917;
  assign new_n9920 = ~new_n9918 & ~new_n9919;
  assign new_n9921 = n3669 & n8332;
  assign new_n9922 = n5470 & n9915;
  assign new_n9923 = new_n9921 & ~new_n9922;
  assign new_n9924 = ~new_n9921 & new_n9922;
  assign new_n9925 = ~new_n9923 & ~new_n9924;
  assign new_n9926 = ~new_n9920 & ~new_n9925;
  assign new_n9927 = new_n9920 & new_n9925;
  assign new_n9928 = ~new_n9926 & ~new_n9927;
  assign new_n9929 = ~new_n9915_1 & new_n9928;
  assign new_n9930 = new_n9915_1 & ~new_n9928;
  assign new_n9931 = ~new_n9929 & ~new_n9930;
  assign new_n9932 = new_n9913 & ~new_n9931;
  assign new_n9933 = ~new_n9913 & new_n9931;
  assign new_n9934 = ~new_n9932 & ~new_n9933;
  assign new_n9935 = n7729 & n10908;
  assign new_n9936 = new_n3840 & ~new_n3843;
  assign new_n9937 = ~new_n3844 & ~new_n9936;
  assign new_n9938 = ~new_n9935 & new_n9937;
  assign new_n9939 = new_n9935 & ~new_n9937;
  assign new_n9940 = ~new_n9938 & ~new_n9939;
  assign new_n9941 = ~new_n3838 & ~new_n3848;
  assign new_n9942 = ~new_n3837 & ~new_n9941;
  assign new_n9943 = n1724 & n8139;
  assign new_n9944 = n3677 & n10560;
  assign new_n9945 = ~new_n9943 & new_n9944;
  assign new_n9946 = new_n9943 & ~new_n9944;
  assign new_n9947 = ~new_n9945 & ~new_n9946;
  assign new_n9948 = n3311 & n12965;
  assign new_n9949 = n6937 & n12003;
  assign new_n9950 = ~new_n9948 & ~new_n9949;
  assign new_n9951 = new_n9948 & new_n9949;
  assign new_n9952 = ~new_n9950 & ~new_n9951;
  assign new_n9953 = ~new_n9947 & new_n9952;
  assign new_n9954 = new_n9947 & ~new_n9952;
  assign new_n9955 = ~new_n9953 & ~new_n9954;
  assign new_n9956 = new_n9942 & new_n9955;
  assign new_n9957 = ~new_n9942 & ~new_n9955;
  assign new_n9958 = ~new_n9956 & ~new_n9957;
  assign new_n9959 = new_n3855 & ~new_n9958;
  assign new_n9960 = ~new_n3855 & new_n9958;
  assign new_n9961 = ~new_n9959 & ~new_n9960;
  assign new_n9962 = ~new_n9940 & ~new_n9961;
  assign new_n9963 = new_n9940 & new_n9961;
  assign new_n9964 = ~new_n9962 & ~new_n9963;
  assign new_n9965 = ~new_n9934 & new_n9964;
  assign new_n9966 = new_n9934 & ~new_n9964;
  assign new_n9967 = ~new_n9965 & ~new_n9966;
  assign new_n9968 = new_n9911 & new_n9967;
  assign new_n9969 = ~new_n9911 & ~new_n9967;
  assign new_n9970 = ~new_n9968 & ~new_n9969;
  assign new_n9971 = ~new_n3860 & ~new_n3863;
  assign new_n9972 = ~new_n3859 & ~new_n9971;
  assign new_n9973 = n603 & n5801;
  assign new_n9974 = n10606 & ~n10866;
  assign new_n9975 = n9041 & n10408;
  assign new_n9976 = new_n9974 & ~new_n9975;
  assign new_n9977 = ~new_n9974 & new_n9975;
  assign new_n9978 = ~new_n9976 & ~new_n9977;
  assign new_n9979 = new_n9973 & ~new_n9978;
  assign new_n9980 = ~new_n9973 & new_n9978;
  assign new_n9981 = ~new_n9979 & ~new_n9980;
  assign new_n9982 = new_n9972 & ~new_n9981;
  assign new_n9983 = ~new_n9972 & new_n9981;
  assign new_n9984 = ~new_n9982 & ~new_n9983;
  assign new_n9985 = ~new_n9970 & new_n9984;
  assign new_n9986 = new_n9970 & ~new_n9984;
  assign new_n9987 = ~new_n9985 & ~new_n9986;
  assign new_n9988 = ~new_n3979 & new_n9987;
  assign new_n9989 = new_n3979 & ~new_n9987;
  assign new_n9990 = ~new_n9988 & ~new_n9989;
  assign new_n9991 = ~new_n3916 & ~new_n3920;
  assign new_n9992 = ~new_n3941 & ~new_n3951;
  assign new_n9993 = ~new_n3940 & ~new_n9992;
  assign new_n9994 = n1165 & n2057;
  assign new_n9995 = n4357 & n5586;
  assign new_n9996 = new_n9994 & ~new_n9995;
  assign new_n9997 = ~new_n9994 & new_n9995;
  assign new_n9998 = ~new_n9996 & ~new_n9997;
  assign new_n9999 = new_n3943 & ~new_n3946_1;
  assign new_n10000 = ~new_n3947 & ~new_n9999;
  assign new_n10001 = ~new_n9998 & new_n10000;
  assign new_n10002 = new_n9998 & ~new_n10000;
  assign new_n10003 = ~new_n10001 & ~new_n10002;
  assign new_n10004 = ~new_n3927 & ~new_n3931;
  assign new_n10005 = ~new_n3930 & ~new_n10004;
  assign new_n10006 = n1364 & n3832;
  assign new_n10007 = n2882 & n4141;
  assign new_n10008 = ~new_n10006 & ~new_n10007;
  assign new_n10009 = new_n10006 & new_n10007;
  assign new_n10010 = ~new_n10008 & ~new_n10009;
  assign new_n10011 = new_n10005 & new_n10010;
  assign new_n10012 = ~new_n10005 & ~new_n10010;
  assign new_n10013 = ~new_n10011 & ~new_n10012;
  assign new_n10014 = new_n10003 & new_n10013;
  assign new_n10015 = ~new_n10003 & ~new_n10013;
  assign new_n10016 = ~new_n10014 & ~new_n10015;
  assign new_n10017 = ~new_n9993 & new_n10016;
  assign new_n10018 = new_n9993 & ~new_n10016;
  assign new_n10019 = ~new_n10017 & ~new_n10018;
  assign new_n10020 = n5167 & n8233;
  assign new_n10021 = n937 & n9887;
  assign new_n10022 = n4335 & n12605;
  assign new_n10023 = ~new_n10021 & ~new_n10022;
  assign new_n10024 = new_n10021 & new_n10022;
  assign new_n10025 = ~new_n10023 & ~new_n10024;
  assign new_n10026 = new_n10020 & new_n10025;
  assign new_n10027 = ~new_n10020 & ~new_n10025;
  assign new_n10028 = ~new_n10026 & ~new_n10027;
  assign new_n10029 = n497 & n10642;
  assign new_n10030 = n2174 & n2777;
  assign new_n10031 = new_n10029 & ~new_n10030;
  assign new_n10032 = ~new_n10029 & new_n10030;
  assign new_n10033 = ~new_n10031 & ~new_n10032;
  assign new_n10034 = new_n3958 & new_n10033;
  assign new_n10035 = ~new_n3958 & ~new_n10033;
  assign new_n10036 = ~new_n10034 & ~new_n10035;
  assign new_n10037 = new_n10028 & ~new_n10036;
  assign new_n10038 = ~new_n10028 & new_n10036;
  assign new_n10039 = ~new_n10037 & ~new_n10038;
  assign new_n10040 = ~new_n10019 & new_n10039;
  assign new_n10041 = new_n10019 & ~new_n10039;
  assign new_n10042 = ~new_n10040 & ~new_n10041;
  assign new_n10043 = n3591 & n5671;
  assign new_n10044 = ~new_n3875 & ~new_n3911;
  assign new_n10045 = ~new_n3876 & ~new_n10044;
  assign new_n10046 = new_n10043 & new_n10045;
  assign new_n10047 = ~new_n10043 & ~new_n10045;
  assign new_n10048 = ~new_n10046 & ~new_n10047;
  assign new_n10049 = new_n10042 & new_n10048;
  assign new_n10050 = ~new_n10042 & ~new_n10048;
  assign new_n10051 = ~new_n10049 & ~new_n10050;
  assign new_n10052 = new_n9991 & ~new_n10051;
  assign new_n10053 = ~new_n9991 & new_n10051;
  assign new_n10054 = ~new_n10052 & ~new_n10053;
  assign new_n10055 = ~new_n9990 & new_n10054;
  assign new_n10056 = new_n9990 & ~new_n10054;
  assign new_n10057 = ~new_n10055 & ~new_n10056;
  assign new_n10058 = new_n9910 & ~new_n10057;
  assign new_n10059 = ~new_n9910 & new_n10057;
  assign new_n10060 = ~new_n10058 & ~new_n10059;
  assign new_n10061 = new_n9862 & new_n10060;
  assign new_n10062 = ~new_n9862 & ~new_n10060;
  assign new_n10063_1 = ~new_n10061 & ~new_n10062;
  assign new_n10064 = new_n9861 & new_n10063_1;
  assign new_n10065 = ~new_n9861 & ~new_n10063_1;
  assign n4777 = ~new_n10064 & ~new_n10065;
  assign new_n10067 = ~new_n8939 & ~new_n8940_1;
  assign n4824 = ~new_n8941 & ~new_n10067;
  assign new_n10069 = ~new_n2625 & ~new_n2626;
  assign new_n10070 = new_n2650 & ~new_n10069;
  assign new_n10071 = ~new_n2650 & new_n10069;
  assign n4864 = ~new_n10070 & ~new_n10071;
  assign new_n10073 = ~new_n2601 & ~new_n2602;
  assign new_n10074 = new_n2656 & ~new_n10073;
  assign new_n10075 = ~new_n2656 & new_n10073;
  assign n5003 = new_n10074 | new_n10075;
  assign new_n10077 = ~new_n7802 & ~new_n7803;
  assign new_n10078 = new_n7823 & new_n10077;
  assign new_n10079 = ~new_n7823 & ~new_n10077;
  assign n5060 = new_n10078 | new_n10079;
  assign new_n10081 = ~new_n4022 & ~new_n4023;
  assign new_n10082 = ~new_n4050 & new_n10081;
  assign new_n10083 = new_n4050 & ~new_n10081;
  assign n5364 = new_n10082 | new_n10083;
  assign new_n10085 = ~new_n9331 & ~new_n9332;
  assign new_n10086 = new_n9345 & ~new_n10085;
  assign new_n10087 = ~new_n9345 & new_n10085;
  assign n5549 = ~new_n10086 & ~new_n10087;
  assign new_n10089 = n7772 & n10594;
  assign new_n10090 = n7529 & n9093;
  assign new_n10091 = n7715 & n10451;
  assign new_n10092 = ~new_n10090 & ~new_n10091;
  assign new_n10093 = new_n10090 & new_n10091;
  assign new_n10094 = ~new_n10092 & ~new_n10093;
  assign new_n10095 = new_n10089 & ~new_n10094;
  assign new_n10096 = ~new_n10089 & new_n10094;
  assign new_n10097 = ~new_n10095 & ~new_n10096;
  assign new_n10098 = new_n8945 & ~new_n10097;
  assign new_n10099 = n3409 & n7772;
  assign new_n10100 = new_n10089 & ~new_n10092;
  assign new_n10101_1 = ~new_n10093 & ~new_n10100;
  assign new_n10102 = ~new_n10099 & new_n10101_1;
  assign new_n10103 = new_n10099 & ~new_n10101_1;
  assign new_n10104 = ~new_n10102 & ~new_n10103;
  assign new_n10105 = n7529 & n10594;
  assign new_n10106 = n7715 & n9093;
  assign new_n10107 = n2458 & n10451;
  assign new_n10108 = ~new_n10106 & ~new_n10107;
  assign new_n10109 = new_n10106 & new_n10107;
  assign new_n10110 = ~new_n10108 & ~new_n10109;
  assign new_n10111 = new_n10105 & ~new_n10110;
  assign new_n10112 = ~new_n10105 & new_n10110;
  assign new_n10113_1 = ~new_n10111 & ~new_n10112;
  assign new_n10114 = ~new_n10104 & new_n10113_1;
  assign new_n10115 = new_n10104 & ~new_n10113_1;
  assign new_n10116 = ~new_n10114 & ~new_n10115;
  assign new_n10117 = ~new_n10098 & ~new_n10116;
  assign new_n10118 = new_n10098 & new_n10116;
  assign new_n10119 = ~new_n10117 & ~new_n10118;
  assign new_n10120 = n9216 & n9906;
  assign new_n10121 = n6085 & n12348;
  assign new_n10122_1 = n2068 & n5962;
  assign new_n10123 = ~new_n10121 & ~new_n10122_1;
  assign new_n10124 = new_n10121 & new_n10122_1;
  assign new_n10125 = ~new_n10123 & ~new_n10124;
  assign new_n10126 = new_n10120 & ~new_n10125;
  assign new_n10127 = ~new_n10120 & new_n10125;
  assign new_n10128 = ~new_n10126 & ~new_n10127;
  assign new_n10129 = new_n8953 & ~new_n10128;
  assign new_n10130 = n9216 & n11109;
  assign new_n10131 = new_n10120 & ~new_n10123;
  assign new_n10132 = ~new_n10124 & ~new_n10131;
  assign new_n10133 = ~new_n10130 & new_n10132;
  assign new_n10134 = new_n10130 & ~new_n10132;
  assign new_n10135 = ~new_n10133 & ~new_n10134;
  assign new_n10136 = n9906 & n12348;
  assign new_n10137 = n2068 & n6085;
  assign new_n10138 = n5962 & n11324;
  assign new_n10139 = ~new_n10137 & ~new_n10138;
  assign new_n10140 = new_n10137 & new_n10138;
  assign new_n10141 = ~new_n10139 & ~new_n10140;
  assign new_n10142_1 = new_n10136 & ~new_n10141;
  assign new_n10143 = ~new_n10136 & new_n10141;
  assign new_n10144 = ~new_n10142_1 & ~new_n10143;
  assign new_n10145 = ~new_n10135 & new_n10144;
  assign new_n10146 = new_n10135 & ~new_n10144;
  assign new_n10147 = ~new_n10145 & ~new_n10146;
  assign new_n10148 = ~new_n10129 & ~new_n10147;
  assign new_n10149 = new_n10129 & new_n10147;
  assign new_n10150 = ~new_n10148 & ~new_n10149;
  assign new_n10151 = n8466 & n12482;
  assign new_n10152 = n5031 & n7720;
  assign new_n10153 = n9 & n287;
  assign new_n10154 = ~new_n10152 & ~new_n10153;
  assign new_n10155 = new_n10152 & new_n10153;
  assign new_n10156 = ~new_n10154 & ~new_n10155;
  assign new_n10157 = new_n10151 & ~new_n10156;
  assign new_n10158 = ~new_n10151 & new_n10156;
  assign new_n10159 = ~new_n10157 & ~new_n10158;
  assign new_n10160 = new_n8961 & ~new_n10159;
  assign new_n10161 = n8466 & n9570;
  assign new_n10162_1 = new_n10151 & ~new_n10154;
  assign new_n10163 = ~new_n10155 & ~new_n10162_1;
  assign new_n10164 = ~new_n10161 & new_n10163;
  assign new_n10165 = new_n10161 & ~new_n10163;
  assign new_n10166 = ~new_n10164 & ~new_n10165;
  assign new_n10167 = n5031 & n12482;
  assign new_n10168_1 = n9 & n7720;
  assign new_n10169 = n287 & n2592;
  assign new_n10170 = ~new_n10168_1 & ~new_n10169;
  assign new_n10171 = new_n10168_1 & new_n10169;
  assign new_n10172 = ~new_n10170 & ~new_n10171;
  assign new_n10173 = new_n10167 & ~new_n10172;
  assign new_n10174 = ~new_n10167 & new_n10172;
  assign new_n10175 = ~new_n10173 & ~new_n10174;
  assign new_n10176 = ~new_n10166 & new_n10175;
  assign new_n10177 = new_n10166 & ~new_n10175;
  assign new_n10178 = ~new_n10176 & ~new_n10177;
  assign new_n10179 = ~new_n10160 & ~new_n10178;
  assign new_n10180 = new_n10160 & new_n10178;
  assign new_n10181 = ~new_n10179 & ~new_n10180;
  assign new_n10182 = n3178 & n5969;
  assign new_n10183 = n1007 & n12592;
  assign new_n10184 = n10168 & n11058;
  assign new_n10185 = ~new_n10183 & ~new_n10184;
  assign new_n10186 = new_n10183 & new_n10184;
  assign new_n10187 = ~new_n10185 & ~new_n10186;
  assign new_n10188 = new_n10182 & ~new_n10187;
  assign new_n10189 = ~new_n10182 & new_n10187;
  assign new_n10190 = ~new_n10188 & ~new_n10189;
  assign new_n10191 = new_n8969 & ~new_n10190;
  assign new_n10192 = n2498 & n3178;
  assign new_n10193 = new_n10182 & ~new_n10185;
  assign new_n10194 = ~new_n10186 & ~new_n10193;
  assign new_n10195 = ~new_n10192 & new_n10194;
  assign new_n10196 = new_n10192 & ~new_n10194;
  assign new_n10197 = ~new_n10195 & ~new_n10196;
  assign new_n10198 = n5969 & n12592;
  assign new_n10199 = n1007 & n10168;
  assign new_n10200 = n767 & n11058;
  assign new_n10201 = ~new_n10199 & ~new_n10200;
  assign new_n10202 = new_n10199 & new_n10200;
  assign new_n10203 = ~new_n10201 & ~new_n10202;
  assign new_n10204 = new_n10198 & ~new_n10203;
  assign new_n10205 = ~new_n10198 & new_n10203;
  assign new_n10206 = ~new_n10204 & ~new_n10205;
  assign new_n10207 = ~new_n10197 & new_n10206;
  assign new_n10208 = new_n10197 & ~new_n10206;
  assign new_n10209 = ~new_n10207 & ~new_n10208;
  assign new_n10210 = new_n10191 & new_n10209;
  assign new_n10211 = ~new_n10191 & ~new_n10209;
  assign new_n10212 = ~new_n10210 & ~new_n10211;
  assign new_n10213 = new_n10181 & new_n10212;
  assign new_n10214 = ~new_n10181 & ~new_n10212;
  assign new_n10215 = ~new_n10213 & ~new_n10214;
  assign new_n10216 = ~new_n8961 & new_n10159;
  assign new_n10217 = ~new_n10160 & ~new_n10216;
  assign new_n10218 = ~new_n8969 & new_n10190;
  assign new_n10219 = ~new_n10191 & ~new_n10218;
  assign new_n10220 = new_n10217 & new_n10219;
  assign new_n10221 = ~new_n10217 & ~new_n10219;
  assign new_n10222 = ~new_n8963 & new_n8970;
  assign new_n10223 = ~new_n8964 & ~new_n10222;
  assign new_n10224 = ~new_n10221 & ~new_n10223;
  assign new_n10225 = ~new_n10220 & ~new_n10224;
  assign new_n10226 = new_n10215 & new_n10225;
  assign new_n10227 = ~new_n10215 & ~new_n10225;
  assign new_n10228 = ~new_n10226 & ~new_n10227;
  assign new_n10229 = new_n10150 & ~new_n10228;
  assign new_n10230 = ~new_n10150 & new_n10228;
  assign new_n10231 = ~new_n10229 & ~new_n10230;
  assign new_n10232 = ~new_n8953 & new_n10128;
  assign new_n10233 = ~new_n10129 & ~new_n10232;
  assign new_n10234 = ~new_n8956 & ~new_n8973;
  assign new_n10235 = ~new_n8955 & ~new_n10234;
  assign new_n10236 = new_n10233 & ~new_n10235;
  assign new_n10237 = ~new_n10233 & new_n10235;
  assign new_n10238 = ~new_n10220 & ~new_n10221;
  assign new_n10239 = ~new_n10223 & ~new_n10238;
  assign new_n10240 = new_n10223 & new_n10238;
  assign new_n10241 = ~new_n10239 & ~new_n10240;
  assign new_n10242 = ~new_n10237 & ~new_n10241;
  assign new_n10243_1 = ~new_n10236 & ~new_n10242;
  assign new_n10244 = ~new_n10231 & ~new_n10243_1;
  assign new_n10245 = new_n10231 & new_n10243_1;
  assign new_n10246 = ~new_n10244 & ~new_n10245;
  assign new_n10247 = new_n10119 & ~new_n10246;
  assign new_n10248 = ~new_n10119 & new_n10246;
  assign new_n10249 = ~new_n10247 & ~new_n10248;
  assign new_n10250 = ~new_n8945 & new_n10097;
  assign new_n10251 = ~new_n10098 & ~new_n10250;
  assign new_n10252 = ~new_n10236 & ~new_n10237;
  assign new_n10253 = new_n10241 & ~new_n10252;
  assign new_n10254 = ~new_n10241 & new_n10252;
  assign new_n10255 = ~new_n10253 & ~new_n10254;
  assign new_n10256 = new_n10251 & new_n10255;
  assign new_n10257 = ~new_n10251 & ~new_n10255;
  assign new_n10258 = ~new_n8947 & ~new_n8976;
  assign new_n10259 = ~new_n8948 & ~new_n10258;
  assign new_n10260 = ~new_n10257 & ~new_n10259;
  assign new_n10261 = ~new_n10256 & ~new_n10260;
  assign new_n10262 = new_n10249 & new_n10261;
  assign new_n10263 = ~new_n10249 & ~new_n10261;
  assign n5557 = new_n10262 | new_n10263;
  assign new_n10265 = n7772 & n9669;
  assign new_n10266 = new_n365 & ~new_n368;
  assign new_n10267 = ~new_n369 & ~new_n10266;
  assign new_n10268 = ~new_n10265 & new_n10267;
  assign new_n10269 = new_n10265 & ~new_n10267;
  assign new_n10270 = ~new_n10268 & ~new_n10269;
  assign new_n10271 = n2458 & n12853;
  assign new_n10272 = n7529 & n11891;
  assign new_n10273 = n7715 & n9531;
  assign new_n10274 = ~new_n10272 & ~new_n10273;
  assign new_n10275 = new_n10272 & new_n10273;
  assign new_n10276 = ~new_n10274 & ~new_n10275;
  assign new_n10277 = new_n10271 & ~new_n10276;
  assign new_n10278 = ~new_n10271 & new_n10276;
  assign new_n10279 = ~new_n10277 & ~new_n10278;
  assign new_n10280 = ~new_n10270 & new_n10279;
  assign new_n10281 = new_n10270 & ~new_n10279;
  assign new_n10282 = ~new_n10280 & ~new_n10281;
  assign new_n10283 = ~new_n375 & ~new_n10282;
  assign new_n10284 = new_n375 & new_n10282;
  assign new_n10285 = ~new_n10283 & ~new_n10284;
  assign new_n10286 = ~new_n457 & ~new_n460_1;
  assign new_n10287 = ~new_n456 & ~new_n10286;
  assign new_n10288 = new_n432 & ~new_n435;
  assign new_n10289 = ~new_n436 & ~new_n10288;
  assign new_n10290 = n510 & n2592;
  assign new_n10291 = n5031 & n9591;
  assign new_n10292 = n9 & n8290;
  assign new_n10293 = ~new_n10291 & ~new_n10292;
  assign new_n10294 = new_n10291 & new_n10292;
  assign new_n10295 = ~new_n10293 & ~new_n10294;
  assign new_n10296 = new_n10290 & ~new_n10295;
  assign new_n10297 = ~new_n10290 & new_n10295;
  assign new_n10298 = ~new_n10296 & ~new_n10297;
  assign new_n10299 = ~new_n10289 & ~new_n10298;
  assign new_n10300 = new_n10289 & new_n10298;
  assign new_n10301 = ~new_n10299 & ~new_n10300;
  assign new_n10302 = ~new_n442 & ~new_n10301;
  assign new_n10303 = new_n442 & new_n10301;
  assign new_n10304 = ~new_n10302 & ~new_n10303;
  assign new_n10305 = n3178 & n13060;
  assign new_n10306 = new_n444 & ~new_n447;
  assign new_n10307 = ~new_n448 & ~new_n10306;
  assign new_n10308 = ~new_n10305 & new_n10307;
  assign new_n10309 = new_n10305 & ~new_n10307;
  assign new_n10310 = ~new_n10308 & ~new_n10309;
  assign new_n10311 = n767 & n834;
  assign new_n10312 = n5189 & n12592;
  assign new_n10313 = n8716 & n10168;
  assign new_n10314 = ~new_n10312 & ~new_n10313;
  assign new_n10315 = new_n10312 & new_n10313;
  assign new_n10316 = ~new_n10314 & ~new_n10315;
  assign new_n10317 = new_n10311 & ~new_n10316;
  assign new_n10318 = ~new_n10311 & new_n10316;
  assign new_n10319 = ~new_n10317 & ~new_n10318;
  assign new_n10320 = ~new_n10310 & new_n10319;
  assign new_n10321 = new_n10310 & ~new_n10319;
  assign new_n10322 = ~new_n10320 & ~new_n10321;
  assign new_n10323 = new_n454 & new_n10322;
  assign new_n10324 = ~new_n454 & ~new_n10322;
  assign new_n10325 = ~new_n10323 & ~new_n10324;
  assign new_n10326 = new_n10304 & new_n10325;
  assign new_n10327 = ~new_n10304 & ~new_n10325;
  assign new_n10328 = ~new_n10326 & ~new_n10327;
  assign new_n10329 = new_n10287 & ~new_n10328;
  assign new_n10330 = ~new_n10287 & new_n10328;
  assign new_n10331 = ~new_n10329 & ~new_n10330;
  assign new_n10332 = n854 & n11324;
  assign new_n10333 = ~new_n424 & ~new_n10332;
  assign new_n10334 = new_n388 & new_n10333;
  assign new_n10335 = ~new_n425 & new_n10332;
  assign new_n10336 = ~new_n10334 & ~new_n10335;
  assign new_n10337 = new_n10331 & ~new_n10336;
  assign new_n10338 = ~new_n10331 & new_n10336;
  assign new_n10339 = ~new_n10337 & ~new_n10338;
  assign new_n10340 = ~new_n429 & new_n463;
  assign new_n10341 = ~new_n430 & ~new_n10340;
  assign new_n10342 = ~new_n10339 & new_n10341;
  assign new_n10343 = new_n10339 & ~new_n10341;
  assign new_n10344 = ~new_n10342 & ~new_n10343;
  assign new_n10345 = new_n10285 & new_n10344;
  assign new_n10346 = ~new_n10285 & ~new_n10344;
  assign new_n10347 = ~new_n10345 & ~new_n10346;
  assign new_n10348 = ~new_n420 & ~new_n466;
  assign new_n10349 = ~new_n421 & ~new_n10348;
  assign new_n10350 = new_n10347 & new_n10349;
  assign new_n10351 = ~new_n10347 & ~new_n10349;
  assign n5609 = new_n10350 | new_n10351;
  assign new_n10353 = ~new_n4879 & ~new_n4880;
  assign new_n10354 = new_n4904 & ~new_n10353;
  assign new_n10355 = ~new_n4904 & new_n10353;
  assign n5882 = ~new_n10354 & ~new_n10355;
  assign new_n10357 = ~new_n5279 & ~new_n5280;
  assign new_n10358 = new_n5294 & ~new_n10357;
  assign new_n10359 = ~new_n5294 & new_n10357;
  assign n6019 = new_n10358 | new_n10359;
  assign new_n10361 = ~new_n7352 & ~new_n7353;
  assign new_n10362 = new_n7355 & ~new_n10361;
  assign new_n10363 = ~new_n7355 & new_n10361;
  assign n6103 = new_n10362 | new_n10363;
  assign new_n10365 = ~new_n1342 & ~new_n1343;
  assign new_n10366 = ~new_n1397 & ~new_n10365;
  assign new_n10367 = new_n1397 & new_n10365;
  assign n6109 = new_n10366 | new_n10367;
  assign new_n10369 = n2482 & n10113;
  assign new_n10370 = n2482 & n11734;
  assign new_n10371 = n10113 & new_n10370;
  assign new_n10372 = ~n10113 & ~new_n10370;
  assign new_n10373 = ~new_n10371 & ~new_n10372;
  assign new_n10374 = ~n1757 & ~new_n10373;
  assign new_n10375 = n1757 & ~new_n10372;
  assign new_n10376 = ~new_n10371 & new_n10375;
  assign new_n10377 = ~new_n10374 & ~new_n10376;
  assign new_n10378 = new_n10369 & new_n10377;
  assign new_n10379 = ~new_n10369 & ~new_n10377;
  assign new_n10380 = ~new_n10378 & ~new_n10379;
  assign new_n10381 = n8228 & n9475;
  assign new_n10382 = n411 & n11236;
  assign new_n10383 = new_n10381 & new_n10382;
  assign new_n10384 = n411 & n4382;
  assign new_n10385 = n9475 & n11236;
  assign new_n10386 = n6826 & n8228;
  assign new_n10387 = ~new_n10385 & ~new_n10386;
  assign new_n10388 = new_n10385 & new_n10386;
  assign new_n10389 = ~new_n10387 & ~new_n10388;
  assign new_n10390 = new_n10384 & ~new_n10389;
  assign new_n10391 = ~new_n10384 & new_n10389;
  assign new_n10392 = ~new_n10390 & ~new_n10391;
  assign new_n10393 = new_n10383 & ~new_n10392;
  assign new_n10394 = ~new_n10383 & new_n10392;
  assign new_n10395 = ~new_n10393 & ~new_n10394;
  assign new_n10396 = n5536 & n8940;
  assign new_n10397 = n4964 & n8506;
  assign new_n10398 = new_n10396 & new_n10397;
  assign new_n10399 = n5684 & n8506;
  assign new_n10400 = n4964 & n5536;
  assign new_n10401 = n772 & n8940;
  assign new_n10402 = ~new_n10400 & ~new_n10401;
  assign new_n10403 = new_n10400 & new_n10401;
  assign new_n10404 = ~new_n10402 & ~new_n10403;
  assign new_n10405 = new_n10399 & ~new_n10404;
  assign new_n10406 = ~new_n10399 & new_n10404;
  assign new_n10407 = ~new_n10405 & ~new_n10406;
  assign new_n10408_1 = new_n10398 & ~new_n10407;
  assign new_n10409 = ~new_n10398 & new_n10407;
  assign new_n10410 = ~new_n10408_1 & ~new_n10409;
  assign new_n10411 = n124 & n9353;
  assign new_n10412 = n3085 & n6333;
  assign new_n10413 = new_n10411 & new_n10412;
  assign new_n10414 = n1912 & n3085;
  assign new_n10415 = n124 & n6333;
  assign new_n10416_1 = n9353 & n10805;
  assign new_n10417 = ~new_n10415 & ~new_n10416_1;
  assign new_n10418 = new_n10415 & new_n10416_1;
  assign new_n10419 = ~new_n10417 & ~new_n10418;
  assign new_n10420 = new_n10414 & ~new_n10419;
  assign new_n10421 = ~new_n10414 & new_n10419;
  assign new_n10422 = ~new_n10420 & ~new_n10421;
  assign new_n10423 = new_n10413 & ~new_n10422;
  assign new_n10424 = ~new_n10413 & new_n10422;
  assign new_n10425 = ~new_n10423 & ~new_n10424;
  assign new_n10426 = ~new_n10410 & ~new_n10425;
  assign new_n10427 = new_n10410 & new_n10425;
  assign new_n10428 = ~new_n10426 & ~new_n10427;
  assign new_n10429 = ~new_n10396 & ~new_n10397;
  assign new_n10430 = ~new_n10398 & ~new_n10429;
  assign new_n10431 = new_n5172 & new_n10430;
  assign new_n10432 = ~new_n10411 & ~new_n10412;
  assign new_n10433 = ~new_n10413 & ~new_n10432;
  assign new_n10434 = ~new_n5172 & ~new_n10430;
  assign new_n10435 = new_n10433 & ~new_n10434;
  assign new_n10436 = ~new_n10431 & ~new_n10435;
  assign new_n10437 = ~new_n10428 & ~new_n10436;
  assign new_n10438 = new_n10428 & new_n10436;
  assign new_n10439 = ~new_n10437 & ~new_n10438;
  assign new_n10440 = new_n10395 & ~new_n10439;
  assign new_n10441 = ~new_n10395 & new_n10439;
  assign new_n10442 = ~new_n10440 & ~new_n10441;
  assign new_n10443 = ~new_n10381 & ~new_n10382;
  assign new_n10444 = ~new_n10383 & ~new_n10443;
  assign new_n10445 = ~new_n10431 & ~new_n10434;
  assign new_n10446 = ~new_n10433 & new_n10445;
  assign new_n10447 = new_n10433 & ~new_n10445;
  assign new_n10448 = ~new_n10446 & ~new_n10447;
  assign new_n10449 = ~new_n10444 & new_n10448;
  assign new_n10450 = new_n10444 & ~new_n10448;
  assign new_n10451_1 = ~new_n5176 & ~new_n10450;
  assign new_n10452 = ~new_n10449 & ~new_n10451_1;
  assign new_n10453_1 = ~new_n10442 & ~new_n10452;
  assign new_n10454 = new_n10442 & new_n10452;
  assign new_n10455 = ~new_n10453_1 & ~new_n10454;
  assign new_n10456 = new_n10380 & new_n10455;
  assign new_n10457 = ~new_n10380 & ~new_n10455;
  assign new_n10458 = ~n10113 & new_n5179;
  assign new_n10459 = ~new_n10449 & ~new_n10450;
  assign new_n10460 = new_n5176 & ~new_n10459;
  assign new_n10461 = ~new_n5176 & new_n10459;
  assign new_n10462 = ~new_n10460 & ~new_n10461;
  assign new_n10463 = ~new_n10458 & new_n10462;
  assign new_n10464 = ~n2482 & ~n10113;
  assign new_n10465 = ~new_n5178 & new_n10369;
  assign new_n10466 = ~new_n10464 & ~new_n10465;
  assign new_n10467 = ~new_n10463 & new_n10466;
  assign new_n10468 = ~new_n10457 & new_n10467;
  assign new_n10469 = ~new_n10456 & ~new_n10468;
  assign new_n10470 = n10113 & n11734;
  assign new_n10471 = n1757 & new_n10470;
  assign new_n10472 = ~n1757 & ~new_n10470;
  assign new_n10473 = ~new_n10471 & ~new_n10472;
  assign new_n10474 = n10416 & ~new_n10473;
  assign new_n10475 = ~n10416 & new_n10473;
  assign new_n10476 = ~new_n10474 & ~new_n10475;
  assign new_n10477 = n2482 & n12651;
  assign new_n10478 = ~new_n10371 & ~new_n10375;
  assign new_n10479 = ~new_n10477 & new_n10478;
  assign new_n10480 = new_n10477 & ~new_n10478;
  assign new_n10481 = ~new_n10479 & ~new_n10480;
  assign new_n10482 = ~new_n10476 & new_n10481;
  assign new_n10483 = new_n10476 & ~new_n10481;
  assign new_n10484 = ~new_n10482 & ~new_n10483;
  assign new_n10485 = ~new_n10378 & ~new_n10484;
  assign new_n10486 = new_n10378 & new_n10484;
  assign new_n10487 = ~new_n10485 & ~new_n10486;
  assign new_n10488 = n8228 & n12284;
  assign new_n10489 = new_n10384 & ~new_n10387;
  assign new_n10490 = ~new_n10388 & ~new_n10489;
  assign new_n10491 = ~new_n10488 & new_n10490;
  assign new_n10492 = new_n10488 & ~new_n10490;
  assign new_n10493 = ~new_n10491 & ~new_n10492;
  assign new_n10494 = n411 & n3130;
  assign new_n10495 = n6826 & n11236;
  assign new_n10496 = n4382 & n9475;
  assign new_n10497 = ~new_n10495 & ~new_n10496;
  assign new_n10498 = new_n10495 & new_n10496;
  assign new_n10499 = ~new_n10497 & ~new_n10498;
  assign new_n10500 = new_n10494 & ~new_n10499;
  assign new_n10501 = ~new_n10494 & new_n10499;
  assign new_n10502 = ~new_n10500 & ~new_n10501;
  assign new_n10503 = ~new_n10493 & new_n10502;
  assign new_n10504 = new_n10493 & ~new_n10502;
  assign new_n10505 = ~new_n10503 & ~new_n10504;
  assign new_n10506 = ~new_n10393 & ~new_n10505;
  assign new_n10507 = new_n10393 & new_n10505;
  assign new_n10508 = ~new_n10506 & ~new_n10507;
  assign new_n10509 = n2737 & n8940;
  assign new_n10510 = new_n10399 & ~new_n10402;
  assign new_n10511 = ~new_n10403 & ~new_n10510;
  assign new_n10512 = ~new_n10509 & new_n10511;
  assign new_n10513 = new_n10509 & ~new_n10511;
  assign new_n10514 = ~new_n10512 & ~new_n10513;
  assign new_n10515 = n8506 & n10522;
  assign new_n10516 = n772 & n4964;
  assign new_n10517 = n5536 & n5684;
  assign new_n10518 = ~new_n10516 & ~new_n10517;
  assign new_n10519 = new_n10516 & new_n10517;
  assign new_n10520 = ~new_n10518 & ~new_n10519;
  assign new_n10521 = new_n10515 & ~new_n10520;
  assign new_n10522_1 = ~new_n10515 & new_n10520;
  assign new_n10523 = ~new_n10521 & ~new_n10522_1;
  assign new_n10524_1 = ~new_n10514 & new_n10523;
  assign new_n10525 = new_n10514 & ~new_n10523;
  assign new_n10526 = ~new_n10524_1 & ~new_n10525;
  assign new_n10527 = ~new_n10408_1 & ~new_n10526;
  assign new_n10528 = new_n10408_1 & new_n10526;
  assign new_n10529 = ~new_n10527 & ~new_n10528;
  assign new_n10530 = n9353 & n12263;
  assign new_n10531 = ~new_n10414 & ~new_n10418;
  assign new_n10532 = ~new_n10417 & ~new_n10531;
  assign new_n10533 = ~new_n10530 & ~new_n10532;
  assign new_n10534 = new_n10530 & new_n10532;
  assign new_n10535 = ~new_n10533 & ~new_n10534;
  assign new_n10536 = n124 & n1912;
  assign new_n10537 = n6333 & n10805;
  assign new_n10538 = n3085 & n12750;
  assign new_n10539 = ~new_n10537 & ~new_n10538;
  assign new_n10540 = new_n10537 & new_n10538;
  assign new_n10541 = ~new_n10539 & ~new_n10540;
  assign new_n10542 = new_n10536 & ~new_n10541;
  assign new_n10543 = ~new_n10536 & new_n10541;
  assign new_n10544 = ~new_n10542 & ~new_n10543;
  assign new_n10545 = ~new_n10535 & new_n10544;
  assign new_n10546 = new_n10535 & ~new_n10544;
  assign new_n10547 = ~new_n10545 & ~new_n10546;
  assign new_n10548 = new_n10423 & new_n10547;
  assign new_n10549 = ~new_n10423 & ~new_n10547;
  assign new_n10550 = ~new_n10548 & ~new_n10549;
  assign new_n10551 = new_n10529 & new_n10550;
  assign new_n10552 = ~new_n10529 & ~new_n10550;
  assign new_n10553 = ~new_n10551 & ~new_n10552;
  assign new_n10554 = ~new_n10426 & ~new_n10436;
  assign new_n10555 = ~new_n10427 & ~new_n10554;
  assign new_n10556 = new_n10553 & new_n10555;
  assign new_n10557 = ~new_n10553 & ~new_n10555;
  assign new_n10558 = ~new_n10556 & ~new_n10557;
  assign new_n10559 = new_n10508 & ~new_n10558;
  assign new_n10560_1 = ~new_n10508 & new_n10558;
  assign new_n10561 = ~new_n10559 & ~new_n10560_1;
  assign new_n10562 = ~new_n10440 & ~new_n10452;
  assign new_n10563 = ~new_n10441 & ~new_n10562;
  assign new_n10564 = ~new_n10561 & new_n10563;
  assign new_n10565 = new_n10561 & ~new_n10563;
  assign new_n10566 = ~new_n10564 & ~new_n10565;
  assign new_n10567 = ~new_n10487 & new_n10566;
  assign new_n10568 = new_n10487 & ~new_n10566;
  assign new_n10569 = ~new_n10567 & ~new_n10568;
  assign new_n10570 = new_n10469 & new_n10569;
  assign new_n10571 = ~new_n10469 & ~new_n10569;
  assign n6297 = new_n10570 | new_n10571;
  assign new_n10573 = new_n7344 & new_n7357;
  assign new_n10574 = new_n7345 & ~new_n7357;
  assign new_n10575 = new_n7359 & ~new_n10574;
  assign n6301 = new_n10573 | new_n10575;
  assign new_n10577 = ~new_n10256 & ~new_n10257;
  assign new_n10578 = new_n10259 & ~new_n10577;
  assign new_n10579 = ~new_n10259 & new_n10577;
  assign n6434 = ~new_n10578 & ~new_n10579;
  assign new_n10581 = ~new_n10456 & ~new_n10457;
  assign new_n10582 = ~new_n10467 & ~new_n10581;
  assign new_n10583 = new_n10467 & new_n10581;
  assign n6586 = ~new_n10582 & ~new_n10583;
  assign new_n10585 = n3006 & ~n7161;
  assign new_n10586 = ~new_n9306 & ~new_n9310;
  assign new_n10587 = ~new_n9307 & ~new_n10586;
  assign new_n10588 = n8308 & n12651;
  assign new_n10589 = n5568 & n7411;
  assign new_n10590 = new_n10588 & new_n10589;
  assign new_n10591 = ~new_n10588 & ~new_n10589;
  assign new_n10592 = ~new_n10590 & ~new_n10591;
  assign new_n10593 = n5214 & n11734;
  assign new_n10594_1 = n2771 & n6168;
  assign new_n10595 = ~n2771 & ~n6168;
  assign new_n10596 = ~new_n10594_1 & ~new_n10595;
  assign new_n10597 = ~new_n10593 & ~new_n10596;
  assign new_n10598 = new_n10593 & new_n10596;
  assign new_n10599 = ~new_n10597 & ~new_n10598;
  assign new_n10600 = new_n9293 & new_n10599;
  assign new_n10601 = ~new_n9293 & ~new_n10599;
  assign new_n10602 = ~new_n10600 & ~new_n10601;
  assign new_n10603 = ~new_n10592 & new_n10602;
  assign new_n10604 = new_n10592 & ~new_n10602;
  assign new_n10605 = ~new_n10603 & ~new_n10604;
  assign new_n10606_1 = ~new_n9297 & ~new_n9300_1;
  assign new_n10607 = ~new_n9301 & ~new_n10606_1;
  assign new_n10608 = ~new_n10605 & new_n10607;
  assign new_n10609 = new_n10605 & ~new_n10607;
  assign new_n10610 = ~new_n10608 & ~new_n10609;
  assign new_n10611 = ~new_n10587 & new_n10610;
  assign new_n10612 = new_n10587 & ~new_n10610;
  assign new_n10613 = ~new_n10611 & ~new_n10612;
  assign new_n10614 = new_n10585 & new_n10613;
  assign new_n10615 = ~new_n10585 & ~new_n10613;
  assign new_n10616 = ~new_n10614 & ~new_n10615;
  assign new_n10617 = new_n9314 & new_n10616;
  assign new_n10618 = ~new_n10614 & ~new_n10617;
  assign new_n10619 = ~new_n10603 & ~new_n10607;
  assign new_n10620 = new_n10590 & new_n10619;
  assign new_n10621 = ~new_n10590 & ~new_n10619;
  assign new_n10622 = ~new_n10604 & new_n10621;
  assign new_n10623 = ~new_n10620 & ~new_n10622;
  assign new_n10624 = new_n9293 & ~new_n10598;
  assign new_n10625 = ~new_n10597 & ~new_n10624;
  assign new_n10626 = n7411 & n8308;
  assign new_n10627 = n5568 & ~n7161;
  assign new_n10628_1 = n3006 & n6149;
  assign new_n10629 = ~new_n10627 & ~new_n10628_1;
  assign new_n10630 = new_n10627 & new_n10628_1;
  assign new_n10631 = ~new_n10629 & ~new_n10630;
  assign new_n10632 = new_n10626 & ~new_n10631;
  assign new_n10633 = ~new_n10626 & new_n10631;
  assign new_n10634 = ~new_n10632 & ~new_n10633;
  assign new_n10635 = new_n10625 & ~new_n10634;
  assign new_n10636 = ~new_n10625 & new_n10634;
  assign new_n10637 = ~new_n10635 & ~new_n10636;
  assign new_n10638 = n5214 & n12651;
  assign new_n10639 = ~new_n10594_1 & ~new_n10638;
  assign new_n10640 = new_n10594_1 & new_n10638;
  assign new_n10641 = ~new_n10639 & ~new_n10640;
  assign new_n10642_1 = n2771 & n11734;
  assign new_n10643 = n6168 & new_n10642_1;
  assign new_n10644 = ~n6168 & ~new_n10642_1;
  assign new_n10645 = ~new_n10643 & ~new_n10644;
  assign new_n10646 = n11411 & ~new_n10645;
  assign new_n10647 = ~n11411 & new_n10645;
  assign new_n10648 = ~new_n10646 & ~new_n10647;
  assign new_n10649 = new_n10641 & ~new_n10648;
  assign new_n10650 = ~new_n10641 & new_n10648;
  assign new_n10651 = ~new_n10649 & ~new_n10650;
  assign new_n10652 = new_n10637 & new_n10651;
  assign new_n10653 = ~new_n10637 & ~new_n10651;
  assign new_n10654 = ~new_n10652 & ~new_n10653;
  assign new_n10655 = new_n10623 & ~new_n10654;
  assign new_n10656 = ~new_n10623 & new_n10654;
  assign new_n10657_1 = ~new_n10655 & ~new_n10656;
  assign new_n10658 = new_n10611 & ~new_n10657_1;
  assign new_n10659 = ~new_n10611 & new_n10657_1;
  assign new_n10660 = ~new_n10658 & ~new_n10659;
  assign new_n10661 = ~new_n10618 & new_n10660;
  assign new_n10662 = new_n10618 & ~new_n10660;
  assign new_n10663 = ~new_n10661 & ~new_n10662;
  assign new_n10664 = n5801 & n12065;
  assign new_n10665 = ~new_n9054 & new_n9057;
  assign new_n10666 = ~new_n9053 & ~new_n10665;
  assign new_n10667 = n10560 & n12284;
  assign new_n10668 = n469 & n10908;
  assign new_n10669 = new_n10667 & new_n10668;
  assign new_n10670 = ~new_n10667 & ~new_n10668;
  assign new_n10671 = ~new_n10669 & ~new_n10670;
  assign new_n10672 = ~new_n9041_1 & ~new_n9045;
  assign new_n10673 = ~new_n9044 & ~new_n10672;
  assign new_n10674 = n6826 & n12003;
  assign new_n10675 = n8139 & n9475;
  assign new_n10676 = n411 & n3311;
  assign new_n10677 = new_n10675 & new_n10676;
  assign new_n10678 = ~new_n10675 & ~new_n10676;
  assign new_n10679 = ~new_n10677 & ~new_n10678;
  assign new_n10680 = new_n10674 & new_n10679;
  assign new_n10681 = ~new_n10674 & ~new_n10679;
  assign new_n10682 = ~new_n10680 & ~new_n10681;
  assign new_n10683 = new_n10673 & ~new_n10682;
  assign new_n10684 = ~new_n10673 & new_n10682;
  assign new_n10685 = ~new_n10683 & ~new_n10684;
  assign new_n10686 = ~new_n10671 & new_n10685;
  assign new_n10687 = new_n10671 & ~new_n10685;
  assign new_n10688 = ~new_n10686 & ~new_n10687;
  assign new_n10689 = ~new_n9039 & new_n9049;
  assign new_n10690 = ~new_n9038 & ~new_n10689;
  assign new_n10691 = ~new_n10688 & new_n10690;
  assign new_n10692 = new_n10688 & ~new_n10690;
  assign new_n10693 = ~new_n10691 & ~new_n10692;
  assign new_n10694 = new_n10666 & ~new_n10693;
  assign new_n10695 = ~new_n10666 & new_n10693;
  assign new_n10696 = ~new_n10694 & ~new_n10695;
  assign new_n10697 = new_n10664 & new_n10696;
  assign new_n10698 = ~new_n10664 & ~new_n10696;
  assign new_n10699 = ~new_n10697 & ~new_n10698;
  assign new_n10700 = new_n9062 & new_n10699;
  assign new_n10701 = ~new_n10697 & ~new_n10700;
  assign new_n10702 = ~new_n10686 & new_n10690;
  assign new_n10703 = new_n10669 & new_n10702;
  assign new_n10704 = ~new_n10669 & ~new_n10702;
  assign new_n10705 = ~new_n10687 & new_n10704;
  assign new_n10706 = ~new_n10703 & ~new_n10705;
  assign new_n10707 = n411 & ~n10866;
  assign new_n10708 = n3311 & n9475;
  assign new_n10709 = n6826 & n8139;
  assign new_n10710 = ~new_n10708 & ~new_n10709;
  assign new_n10711 = new_n10708 & new_n10709;
  assign new_n10712 = ~new_n10710 & ~new_n10711;
  assign new_n10713 = ~new_n10707 & ~new_n10712;
  assign new_n10714 = new_n10707 & new_n10712;
  assign new_n10715 = ~new_n10713 & ~new_n10714;
  assign new_n10716 = n12003 & n12284;
  assign new_n10717 = new_n10677 & new_n10716;
  assign new_n10718 = ~new_n10677 & ~new_n10716;
  assign new_n10719 = ~new_n10717 & ~new_n10718;
  assign new_n10720 = ~new_n10715 & ~new_n10719;
  assign new_n10721 = new_n10715 & new_n10719;
  assign new_n10722 = ~new_n10720 & ~new_n10721;
  assign new_n10723 = n469 & n10560;
  assign new_n10724 = n5801 & n11180;
  assign new_n10725 = n10908 & n12065;
  assign new_n10726 = ~new_n10724 & ~new_n10725;
  assign new_n10727 = new_n10724 & new_n10725;
  assign new_n10728 = ~new_n10726 & ~new_n10727;
  assign new_n10729 = new_n10723 & ~new_n10728;
  assign new_n10730 = ~new_n10723 & new_n10728;
  assign new_n10731 = ~new_n10729 & ~new_n10730;
  assign new_n10732 = ~new_n10673 & ~new_n10680;
  assign new_n10733 = ~new_n10681 & ~new_n10732;
  assign new_n10734 = ~new_n10731 & new_n10733;
  assign new_n10735 = new_n10731 & ~new_n10733;
  assign new_n10736_1 = ~new_n10734 & ~new_n10735;
  assign new_n10737 = ~new_n10722 & new_n10736_1;
  assign new_n10738 = new_n10722 & ~new_n10736_1;
  assign new_n10739 = ~new_n10737 & ~new_n10738;
  assign new_n10740 = new_n10706 & ~new_n10739;
  assign new_n10741 = ~new_n10706 & new_n10739;
  assign new_n10742 = ~new_n10740 & ~new_n10741;
  assign new_n10743 = new_n10694 & new_n10742;
  assign new_n10744 = ~new_n10694 & ~new_n10742;
  assign new_n10745 = ~new_n10743 & ~new_n10744;
  assign new_n10746 = ~new_n10701 & new_n10745;
  assign new_n10747 = new_n10701 & ~new_n10745;
  assign new_n10748 = ~new_n10746 & ~new_n10747;
  assign new_n10749 = n22 & n13201;
  assign new_n10750 = n5586 & n12263;
  assign new_n10751 = n353 & n2057;
  assign new_n10752 = new_n10750 & new_n10751;
  assign new_n10753 = ~new_n10750 & ~new_n10751;
  assign new_n10754 = ~new_n10752 & ~new_n10753;
  assign new_n10755 = n4141 & n10805;
  assign new_n10756 = n124 & n1364;
  assign new_n10757 = n3085 & n3669;
  assign new_n10758 = new_n10756 & new_n10757;
  assign new_n10759 = ~new_n10756 & ~new_n10757;
  assign new_n10760 = ~new_n10758 & ~new_n10759;
  assign new_n10761 = new_n10755 & new_n10760;
  assign new_n10762 = ~new_n10755 & ~new_n10760;
  assign new_n10763 = ~new_n10761 & ~new_n10762;
  assign new_n10764 = new_n9165 & ~new_n9168;
  assign new_n10765 = ~new_n9169 & ~new_n10764;
  assign new_n10766 = ~new_n10763 & ~new_n10765;
  assign new_n10767 = new_n10763 & new_n10765;
  assign new_n10768 = ~new_n10766 & ~new_n10767;
  assign new_n10769 = ~new_n10754 & new_n10768;
  assign new_n10770_1 = new_n10754 & ~new_n10768;
  assign new_n10771 = ~new_n10769 & ~new_n10770_1;
  assign new_n10772 = ~new_n9162 & ~new_n9173;
  assign new_n10773 = ~new_n9163 & ~new_n10772;
  assign new_n10774 = ~new_n10771 & new_n10773;
  assign new_n10775 = new_n10771 & ~new_n10773;
  assign new_n10776 = ~new_n10774 & ~new_n10775;
  assign new_n10777 = ~new_n9177 & ~new_n9181;
  assign new_n10778 = ~new_n9178 & ~new_n10777;
  assign new_n10779 = new_n10776 & ~new_n10778;
  assign new_n10780 = ~new_n10776 & new_n10778;
  assign new_n10781 = ~new_n10779 & ~new_n10780;
  assign new_n10782 = new_n10749 & new_n10781;
  assign new_n10783 = ~new_n10749 & ~new_n10781;
  assign new_n10784 = ~new_n10782 & ~new_n10783;
  assign new_n10785 = new_n9186 & new_n10784;
  assign new_n10786 = ~new_n10782 & ~new_n10785;
  assign new_n10787 = n353 & n5586;
  assign new_n10788 = n11396 & n13201;
  assign new_n10789 = n22 & n2057;
  assign new_n10790 = ~new_n10788 & ~new_n10789;
  assign new_n10791 = new_n10788 & new_n10789;
  assign new_n10792 = ~new_n10790 & ~new_n10791;
  assign new_n10793 = ~new_n10787 & ~new_n10792;
  assign new_n10794 = new_n10787 & new_n10792;
  assign new_n10795 = ~new_n10793 & ~new_n10794;
  assign new_n10796 = ~new_n10761 & new_n10765;
  assign new_n10797_1 = ~new_n10762 & ~new_n10796;
  assign new_n10798 = ~new_n10795 & ~new_n10797_1;
  assign new_n10799 = new_n10795 & new_n10797_1;
  assign new_n10800 = ~new_n10798 & ~new_n10799;
  assign new_n10801 = n4141 & n12263;
  assign new_n10802 = ~new_n10758 & ~new_n10801;
  assign new_n10803 = new_n10758 & new_n10801;
  assign new_n10804 = ~new_n10802 & ~new_n10803;
  assign new_n10805_1 = n3085 & n5470;
  assign new_n10806 = n124 & n3669;
  assign new_n10807 = n1364 & n10805;
  assign new_n10808 = ~new_n10806 & ~new_n10807;
  assign new_n10809 = new_n10806 & new_n10807;
  assign new_n10810 = ~new_n10808 & ~new_n10809;
  assign new_n10811 = new_n10805_1 & ~new_n10810;
  assign new_n10812 = ~new_n10805_1 & new_n10810;
  assign new_n10813 = ~new_n10811 & ~new_n10812;
  assign new_n10814 = ~new_n10804 & new_n10813;
  assign new_n10815 = new_n10804 & ~new_n10813;
  assign new_n10816 = ~new_n10814 & ~new_n10815;
  assign new_n10817 = ~new_n10800 & ~new_n10816;
  assign new_n10818 = new_n10800 & new_n10816;
  assign new_n10819 = ~new_n10817 & ~new_n10818;
  assign new_n10820 = ~new_n10769 & ~new_n10773;
  assign new_n10821 = new_n10752 & new_n10820;
  assign new_n10822 = ~new_n10752 & ~new_n10820;
  assign new_n10823 = ~new_n10770_1 & new_n10822;
  assign new_n10824 = ~new_n10821 & ~new_n10823;
  assign new_n10825 = ~new_n10819 & new_n10824;
  assign new_n10826 = new_n10819 & ~new_n10824;
  assign new_n10827 = ~new_n10825 & ~new_n10826;
  assign new_n10828 = new_n10779 & ~new_n10827;
  assign new_n10829 = ~new_n10779 & new_n10827;
  assign new_n10830 = ~new_n10828 & ~new_n10829;
  assign new_n10831 = ~new_n10786 & new_n10830;
  assign new_n10832 = new_n10786 & ~new_n10830;
  assign new_n10833 = ~new_n10831 & ~new_n10832;
  assign new_n10834 = n4114 & n12408;
  assign new_n10835 = n2737 & n11665;
  assign new_n10836 = new_n10834 & new_n10835;
  assign new_n10837 = ~new_n10834 & ~new_n10835;
  assign new_n10838 = ~new_n10836 & ~new_n10837;
  assign new_n10839 = n772 & n2777;
  assign new_n10840 = n5536 & n10642;
  assign new_n10841 = n937 & n8506;
  assign new_n10842 = new_n10840 & new_n10841;
  assign new_n10843 = ~new_n10840 & ~new_n10841;
  assign new_n10844 = ~new_n10842 & ~new_n10843;
  assign new_n10845 = new_n10839 & new_n10844;
  assign new_n10846 = ~new_n10839 & ~new_n10844;
  assign new_n10847 = ~new_n10845 & ~new_n10846;
  assign new_n10848 = new_n9103 & ~new_n9106;
  assign new_n10849 = ~new_n9107 & ~new_n10848;
  assign new_n10850 = ~new_n10847 & ~new_n10849;
  assign new_n10851 = new_n10847 & new_n10849;
  assign new_n10852 = ~new_n10850 & ~new_n10851;
  assign new_n10853 = ~new_n10838 & new_n10852;
  assign new_n10854 = new_n10838 & ~new_n10852;
  assign new_n10855 = ~new_n10853 & ~new_n10854;
  assign new_n10856 = ~new_n9100_1 & ~new_n9111;
  assign new_n10857 = ~new_n9101 & ~new_n10856;
  assign new_n10858 = ~new_n10855 & new_n10857;
  assign new_n10859 = new_n10855 & ~new_n10857;
  assign new_n10860 = ~new_n10858 & ~new_n10859;
  assign new_n10861 = ~new_n9115 & ~new_n9119;
  assign new_n10862 = ~new_n9116 & ~new_n10861;
  assign new_n10863 = new_n10860 & ~new_n10862;
  assign new_n10864 = n11665 & n12408;
  assign new_n10865 = n5671 & n11350;
  assign new_n10866_1 = n4114 & n9846;
  assign new_n10867 = ~new_n10865 & ~new_n10866_1;
  assign new_n10868 = new_n10865 & new_n10866_1;
  assign new_n10869 = ~new_n10867 & ~new_n10868;
  assign new_n10870 = ~new_n10864 & ~new_n10869;
  assign new_n10871 = new_n10864 & new_n10869;
  assign new_n10872 = ~new_n10870 & ~new_n10871;
  assign new_n10873 = ~new_n10845 & new_n10849;
  assign new_n10874_1 = ~new_n10846 & ~new_n10873;
  assign new_n10875 = ~new_n10872 & ~new_n10874_1;
  assign new_n10876 = n2737 & n2777;
  assign new_n10877 = new_n10842 & new_n10876;
  assign new_n10878 = ~new_n10842 & ~new_n10876;
  assign new_n10879 = ~new_n10877 & ~new_n10878;
  assign new_n10880 = n8506 & n12605;
  assign new_n10881 = n937 & n5536;
  assign new_n10882 = n772 & n10642;
  assign new_n10883 = ~new_n10881 & ~new_n10882;
  assign new_n10884 = new_n10881 & new_n10882;
  assign new_n10885 = ~new_n10883 & ~new_n10884;
  assign new_n10886 = new_n10880 & ~new_n10885;
  assign new_n10887 = ~new_n10880 & new_n10885;
  assign new_n10888 = ~new_n10886 & ~new_n10887;
  assign new_n10889 = new_n10879 & new_n10888;
  assign new_n10890 = ~new_n10879 & ~new_n10888;
  assign new_n10891 = ~new_n10889 & ~new_n10890;
  assign new_n10892 = new_n10875 & new_n10891;
  assign new_n10893 = new_n10872 & new_n10874_1;
  assign new_n10894 = new_n10891 & ~new_n10893;
  assign new_n10895 = ~new_n10875 & ~new_n10894;
  assign new_n10896 = ~new_n10891 & new_n10893;
  assign new_n10897 = new_n10895 & ~new_n10896;
  assign new_n10898 = ~new_n10892 & ~new_n10897;
  assign new_n10899 = ~new_n10853 & ~new_n10857;
  assign new_n10900 = new_n10836 & new_n10899;
  assign new_n10901 = ~new_n10836 & ~new_n10899;
  assign new_n10902 = ~new_n10854 & new_n10901;
  assign new_n10903 = ~new_n10900 & ~new_n10902;
  assign new_n10904 = new_n10898 & new_n10903;
  assign new_n10905 = ~new_n10898 & ~new_n10903;
  assign new_n10906 = ~new_n10904 & ~new_n10905;
  assign new_n10907 = new_n10863 & new_n10906;
  assign new_n10908_1 = ~new_n10863 & ~new_n10906;
  assign new_n10909 = ~new_n10907 & ~new_n10908_1;
  assign new_n10910 = n5671 & n9846;
  assign new_n10911 = ~new_n10860 & new_n10862;
  assign new_n10912 = ~new_n10863 & ~new_n10911;
  assign new_n10913 = new_n10910 & new_n10912;
  assign new_n10914 = ~new_n10910 & ~new_n10912;
  assign new_n10915 = ~new_n10913 & ~new_n10914;
  assign new_n10916 = new_n9124 & new_n10915;
  assign new_n10917 = ~new_n10913 & ~new_n10916;
  assign new_n10918 = new_n10909 & ~new_n10917;
  assign new_n10919 = ~new_n10909 & new_n10917;
  assign new_n10920 = ~new_n10918 & ~new_n10919;
  assign new_n10921 = ~new_n10833 & ~new_n10920;
  assign new_n10922 = new_n10833 & new_n10920;
  assign new_n10923 = ~new_n10921 & ~new_n10922;
  assign new_n10924 = ~new_n9124 & ~new_n10915;
  assign new_n10925 = ~new_n10916 & ~new_n10924;
  assign new_n10926 = ~new_n9186 & ~new_n10784;
  assign new_n10927 = ~new_n10785 & ~new_n10926;
  assign new_n10928 = new_n10925 & new_n10927;
  assign new_n10929 = ~new_n10925 & ~new_n10927;
  assign new_n10930 = ~new_n9188 & ~new_n9217;
  assign new_n10931 = ~new_n9189 & ~new_n10930;
  assign new_n10932 = ~new_n10929 & ~new_n10931;
  assign new_n10933 = ~new_n10928 & ~new_n10932;
  assign new_n10934 = ~new_n10923 & new_n10933;
  assign new_n10935 = new_n10923 & ~new_n10933;
  assign new_n10936 = ~new_n10934 & ~new_n10935;
  assign new_n10937 = ~new_n10748 & ~new_n10936;
  assign new_n10938 = new_n10748 & new_n10936;
  assign new_n10939 = ~new_n10937 & ~new_n10938;
  assign new_n10940 = ~new_n9062 & ~new_n10699;
  assign new_n10941 = ~new_n10700 & ~new_n10940;
  assign new_n10942 = ~new_n10928 & ~new_n10929;
  assign new_n10943 = new_n10931 & ~new_n10942;
  assign new_n10944 = ~new_n10931 & new_n10942;
  assign new_n10945 = ~new_n10943 & ~new_n10944;
  assign new_n10946 = new_n10941 & new_n10945;
  assign new_n10947 = ~new_n10941 & ~new_n10945;
  assign new_n10948 = ~new_n9221 & ~new_n9257;
  assign new_n10949 = ~new_n9222 & ~new_n10948;
  assign new_n10950 = ~new_n10947 & ~new_n10949;
  assign new_n10951 = ~new_n10946 & ~new_n10950;
  assign new_n10952 = ~new_n10939 & new_n10951;
  assign new_n10953 = new_n10939 & ~new_n10951;
  assign new_n10954 = ~new_n10952 & ~new_n10953;
  assign new_n10955 = ~new_n10663 & ~new_n10954;
  assign new_n10956 = new_n10663 & new_n10954;
  assign new_n10957 = ~new_n9314 & ~new_n10616;
  assign new_n10958 = ~new_n10617 & ~new_n10957;
  assign new_n10959 = new_n9260 & ~new_n9350;
  assign new_n10960 = ~new_n9351 & ~new_n10959;
  assign new_n10961 = new_n10958 & ~new_n10960;
  assign new_n10962 = ~new_n10958 & new_n10960;
  assign new_n10963 = ~new_n10946 & ~new_n10947;
  assign new_n10964 = new_n10949 & ~new_n10963;
  assign new_n10965 = ~new_n10949 & new_n10963;
  assign new_n10966 = ~new_n10964 & ~new_n10965;
  assign new_n10967 = ~new_n10962 & new_n10966;
  assign new_n10968 = ~new_n10961 & ~new_n10967;
  assign new_n10969 = ~new_n10956 & new_n10968;
  assign new_n10970 = ~new_n10955 & ~new_n10969;
  assign new_n10971 = ~new_n10907 & ~new_n10918;
  assign new_n10972 = ~new_n10798 & new_n10816;
  assign new_n10973 = ~new_n10799 & ~new_n10972;
  assign new_n10974 = new_n10971 & new_n10973;
  assign new_n10975 = ~new_n10971 & ~new_n10973;
  assign new_n10976 = ~new_n10974 & ~new_n10975;
  assign new_n10977 = ~new_n10658 & ~new_n10661;
  assign new_n10978 = n772 & n937;
  assign new_n10979 = n5536 & n12605;
  assign new_n10980 = ~new_n10978 & ~new_n10979;
  assign new_n10981 = new_n10978 & new_n10979;
  assign new_n10982 = ~new_n10980 & ~new_n10981;
  assign new_n10983 = n2737 & n10642;
  assign new_n10984 = n2777 & n12408;
  assign new_n10985 = new_n10983 & ~new_n10984;
  assign new_n10986 = ~new_n10983 & new_n10984;
  assign new_n10987 = ~new_n10985 & ~new_n10986;
  assign new_n10988 = ~new_n10982 & ~new_n10987;
  assign new_n10989 = new_n10982 & new_n10987;
  assign new_n10990 = ~new_n10988 & ~new_n10989;
  assign new_n10991 = ~new_n10895 & new_n10990;
  assign new_n10992 = new_n10895 & ~new_n10990;
  assign new_n10993 = ~new_n10991 & ~new_n10992;
  assign new_n10994 = ~new_n10877 & new_n10888;
  assign new_n10995 = ~new_n10878 & ~new_n10994;
  assign new_n10996 = n9846 & n11665;
  assign new_n10997 = n4114 & n11350;
  assign new_n10998 = new_n10996 & ~new_n10997;
  assign new_n10999 = ~new_n10996 & new_n10997;
  assign new_n11000 = ~new_n10998 & ~new_n10999;
  assign new_n11001 = new_n10880 & ~new_n10883;
  assign new_n11002 = ~new_n10884 & ~new_n11001;
  assign new_n11003 = new_n10864 & ~new_n10867;
  assign new_n11004 = ~new_n10868 & ~new_n11003;
  assign new_n11005 = ~new_n11002 & new_n11004;
  assign new_n11006 = new_n11002 & ~new_n11004;
  assign new_n11007 = ~new_n11005 & ~new_n11006;
  assign new_n11008 = ~new_n11000 & ~new_n11007;
  assign new_n11009 = new_n11000 & new_n11007;
  assign new_n11010 = ~new_n11008 & ~new_n11009;
  assign new_n11011 = new_n10995 & new_n11010;
  assign new_n11012 = ~new_n10995 & ~new_n11010;
  assign new_n11013 = ~new_n11011 & ~new_n11012;
  assign new_n11014 = new_n10993 & ~new_n11013;
  assign new_n11015 = ~new_n10993 & new_n11013;
  assign new_n11016 = ~new_n11014 & ~new_n11015;
  assign new_n11017 = n3006 & n5715;
  assign new_n11018 = ~n7061 & new_n11017;
  assign new_n11019 = n7061 & ~new_n11017;
  assign new_n11020 = ~new_n11018 & ~new_n11019;
  assign new_n11021 = ~new_n11016 & new_n11020;
  assign new_n11022 = new_n11016 & ~new_n11020;
  assign new_n11023 = ~new_n11021 & ~new_n11022;
  assign new_n11024 = ~new_n10622 & new_n10654;
  assign new_n11025 = ~new_n10620 & ~new_n11024;
  assign new_n11026 = ~new_n10803 & new_n10813;
  assign new_n11027 = ~new_n10802 & ~new_n11026;
  assign new_n11028 = new_n10787 & ~new_n10790;
  assign new_n11029 = ~new_n10791 & ~new_n11028;
  assign new_n11030_1 = new_n10805_1 & ~new_n10808;
  assign new_n11031 = ~new_n10809 & ~new_n11030_1;
  assign new_n11032 = ~new_n11029 & new_n11031;
  assign new_n11033 = new_n11029 & ~new_n11031;
  assign new_n11034 = ~new_n11032 & ~new_n11033;
  assign new_n11035 = new_n11027 & new_n11034;
  assign new_n11036 = ~new_n11027 & ~new_n11034;
  assign new_n11037 = ~new_n11035 & ~new_n11036;
  assign new_n11038 = n2057 & n11396;
  assign new_n11039 = n22 & n5586;
  assign new_n11040 = new_n11038 & ~new_n11039;
  assign new_n11041 = ~new_n11038 & new_n11039;
  assign new_n11042 = ~new_n11040 & ~new_n11041;
  assign new_n11043 = n1364 & n12263;
  assign new_n11044 = n353 & n4141;
  assign new_n11045 = ~new_n11043 & ~new_n11044;
  assign new_n11046 = new_n11043 & new_n11044;
  assign new_n11047 = ~new_n11045 & ~new_n11046;
  assign new_n11048 = n5167 & n8506;
  assign new_n11049 = n4122 & n5671;
  assign new_n11050 = new_n11048 & new_n11049;
  assign new_n11051 = ~new_n11048 & ~new_n11049;
  assign new_n11052 = ~new_n11050 & ~new_n11051;
  assign new_n11053 = new_n11047 & ~new_n11052;
  assign new_n11054 = ~new_n11047 & new_n11052;
  assign new_n11055 = ~new_n11053 & ~new_n11054;
  assign new_n11056 = ~new_n11042 & new_n11055;
  assign new_n11057_1 = new_n11042 & ~new_n11055;
  assign new_n11058_1 = ~new_n11056 & ~new_n11057_1;
  assign new_n11059 = new_n11037 & ~new_n11058_1;
  assign new_n11060 = ~new_n11037 & new_n11058_1;
  assign new_n11061_1 = ~new_n11059 & ~new_n11060;
  assign new_n11062 = new_n10898 & ~new_n10902;
  assign new_n11063 = ~new_n10900 & ~new_n11062;
  assign new_n11064 = new_n11061_1 & new_n11063;
  assign new_n11065 = ~new_n11061_1 & ~new_n11063;
  assign new_n11066 = ~new_n11064 & ~new_n11065;
  assign new_n11067 = new_n11025 & new_n11066;
  assign new_n11068 = ~new_n11025 & ~new_n11066;
  assign new_n11069 = ~new_n11067 & ~new_n11068;
  assign new_n11070 = new_n11023 & new_n11069;
  assign new_n11071 = ~new_n11023 & ~new_n11069;
  assign new_n11072 = ~new_n11070 & ~new_n11071;
  assign new_n11073 = ~new_n10977 & new_n11072;
  assign new_n11074 = new_n10977 & ~new_n11072;
  assign new_n11075 = ~new_n11073 & ~new_n11074;
  assign new_n11076 = ~new_n10976 & ~new_n11075;
  assign new_n11077_1 = new_n10976 & new_n11075;
  assign new_n11078 = ~new_n11076 & ~new_n11077_1;
  assign new_n11079 = ~new_n10937 & ~new_n10951;
  assign new_n11080 = ~new_n10938 & ~new_n11079;
  assign new_n11081 = ~new_n10828 & ~new_n10831;
  assign new_n11082 = n10908 & n11180;
  assign new_n11083 = new_n10707 & ~new_n10710;
  assign new_n11084 = ~new_n10711 & ~new_n11083;
  assign new_n11085 = ~new_n11082 & new_n11084;
  assign new_n11086 = new_n11082 & ~new_n11084;
  assign new_n11087 = ~new_n11085 & ~new_n11086;
  assign new_n11088 = ~new_n10715 & ~new_n10717;
  assign new_n11089 = ~new_n10718 & ~new_n11088;
  assign new_n11090 = new_n11087 & new_n11089;
  assign new_n11091 = ~new_n11087 & ~new_n11089;
  assign new_n11092 = ~new_n11090 & ~new_n11091;
  assign new_n11093 = n8139 & n12284;
  assign new_n11094 = n10560 & n12065;
  assign new_n11095 = new_n11093 & ~new_n11094;
  assign new_n11096 = ~new_n11093 & new_n11094;
  assign new_n11097 = ~new_n11095 & ~new_n11096;
  assign new_n11098 = n3311 & n6826;
  assign new_n11099 = n469 & n12003;
  assign new_n11100 = ~new_n11098 & ~new_n11099;
  assign new_n11101 = new_n11098 & new_n11099;
  assign new_n11102 = ~new_n11100 & ~new_n11101;
  assign new_n11103 = ~new_n11097 & new_n11102;
  assign new_n11104 = new_n11097 & ~new_n11102;
  assign new_n11105 = ~new_n11103 & ~new_n11104;
  assign new_n11106 = ~new_n11092 & new_n11105;
  assign new_n11107 = new_n11092 & ~new_n11105;
  assign new_n11108 = ~new_n11106 & ~new_n11107;
  assign new_n11109_1 = ~new_n10723 & ~new_n10727;
  assign new_n11110 = ~new_n10726 & ~new_n11109_1;
  assign new_n11111_1 = n3085 & n6409;
  assign new_n11112 = n12372 & n13201;
  assign new_n11113 = ~new_n11111_1 & ~new_n11112;
  assign new_n11114 = new_n11111_1 & new_n11112;
  assign new_n11115 = ~new_n11113 & ~new_n11114;
  assign new_n11116 = n3669 & n10805;
  assign new_n11117 = n124 & n5470;
  assign new_n11118 = new_n11116 & ~new_n11117;
  assign new_n11119 = ~new_n11116 & new_n11117;
  assign new_n11120 = ~new_n11118 & ~new_n11119;
  assign new_n11121 = ~new_n11115 & ~new_n11120;
  assign new_n11122 = new_n11115 & new_n11120;
  assign new_n11123 = ~new_n11121 & ~new_n11122;
  assign new_n11124 = ~new_n11110 & new_n11123;
  assign new_n11125 = new_n11110 & ~new_n11123;
  assign new_n11126 = ~new_n11124 & ~new_n11125;
  assign new_n11127 = ~new_n11108 & new_n11126;
  assign new_n11128 = new_n11108 & ~new_n11126;
  assign new_n11129 = ~new_n11127 & ~new_n11128;
  assign new_n11130 = new_n10819 & ~new_n10823;
  assign new_n11131 = ~new_n10821 & ~new_n11130;
  assign new_n11132 = new_n10722 & ~new_n10735;
  assign new_n11133 = ~new_n10734 & ~new_n11132;
  assign new_n11134 = new_n11131 & new_n11133;
  assign new_n11135 = ~new_n11131 & ~new_n11133;
  assign new_n11136 = ~new_n11134 & ~new_n11135;
  assign new_n11137 = new_n11129 & new_n11136;
  assign new_n11138 = ~new_n11129 & ~new_n11136;
  assign new_n11139 = ~new_n11137 & ~new_n11138;
  assign new_n11140_1 = new_n11081 & ~new_n11139;
  assign new_n11141 = ~new_n11081 & new_n11139;
  assign new_n11142 = ~new_n11140_1 & ~new_n11141;
  assign new_n11143 = new_n10626 & ~new_n10629;
  assign new_n11144 = ~new_n10630 & ~new_n11143;
  assign new_n11145 = ~new_n10636 & new_n10651;
  assign new_n11146 = ~new_n10635 & ~new_n11145;
  assign new_n11147_1 = ~new_n11144 & ~new_n11146;
  assign new_n11148 = new_n11144 & new_n11146;
  assign new_n11149 = ~new_n11147_1 & ~new_n11148;
  assign new_n11150 = n2771 & n12651;
  assign new_n11151 = ~n7161 & n8308;
  assign new_n11152 = n5214 & n7411;
  assign new_n11153 = new_n11151 & new_n11152;
  assign new_n11154 = ~new_n11151 & ~new_n11152;
  assign new_n11155 = ~new_n11153 & ~new_n11154;
  assign new_n11156 = new_n11150 & ~new_n11155;
  assign new_n11157 = ~new_n11150 & new_n11155;
  assign new_n11158 = ~new_n11156 & ~new_n11157;
  assign new_n11159 = n5568 & n6149;
  assign new_n11160 = n6168 & n11734;
  assign new_n11161 = ~n11411 & new_n11160;
  assign new_n11162 = n11411 & ~new_n11160;
  assign new_n11163 = ~new_n11161 & ~new_n11162;
  assign new_n11164 = ~new_n11159 & new_n11163;
  assign new_n11165 = new_n11159 & ~new_n11163;
  assign new_n11166 = ~new_n11164 & ~new_n11165;
  assign new_n11167 = ~new_n11158 & new_n11166;
  assign new_n11168 = new_n11158 & ~new_n11166;
  assign new_n11169 = ~new_n11167 & ~new_n11168;
  assign new_n11170 = ~new_n10640 & new_n10648;
  assign new_n11171 = ~new_n10639 & ~new_n11170;
  assign new_n11172 = n11411 & ~new_n10644;
  assign new_n11173 = ~new_n10643 & ~new_n11172;
  assign new_n11174 = new_n11171 & new_n11173;
  assign new_n11175 = ~new_n11171 & ~new_n11173;
  assign new_n11176 = ~new_n11174 & ~new_n11175;
  assign new_n11177 = ~new_n11169 & new_n11176;
  assign new_n11178 = new_n11169 & ~new_n11176;
  assign new_n11179 = ~new_n11177 & ~new_n11178;
  assign new_n11180_1 = new_n11149 & new_n11179;
  assign new_n11181 = ~new_n11149 & ~new_n11179;
  assign new_n11182 = ~new_n11180_1 & ~new_n11181;
  assign new_n11183 = ~new_n10705 & ~new_n10739;
  assign new_n11184 = ~new_n10703 & ~new_n11183;
  assign new_n11185 = n5801 & n12912;
  assign new_n11186 = n9475 & ~n10866;
  assign new_n11187 = n411 & n9041;
  assign new_n11188 = new_n11186 & ~new_n11187;
  assign new_n11189 = ~new_n11186 & new_n11187;
  assign new_n11190 = ~new_n11188 & ~new_n11189;
  assign new_n11191 = new_n11185 & ~new_n11190;
  assign new_n11192 = ~new_n11185 & new_n11190;
  assign new_n11193 = ~new_n11191 & ~new_n11192;
  assign new_n11194 = ~new_n11184 & new_n11193;
  assign new_n11195 = new_n11184 & ~new_n11193;
  assign new_n11196 = ~new_n11194 & ~new_n11195;
  assign new_n11197 = new_n11182 & new_n11196;
  assign new_n11198 = ~new_n11182 & ~new_n11196;
  assign new_n11199 = ~new_n11197 & ~new_n11198;
  assign new_n11200 = ~new_n11142 & new_n11199;
  assign new_n11201 = new_n11142 & ~new_n11199;
  assign new_n11202 = ~new_n11200 & ~new_n11201;
  assign new_n11203 = ~new_n10743 & ~new_n10746;
  assign new_n11204 = ~new_n10921 & ~new_n10933;
  assign new_n11205 = ~new_n10922 & ~new_n11204;
  assign new_n11206 = new_n11203 & new_n11205;
  assign new_n11207 = ~new_n11203 & ~new_n11205;
  assign new_n11208 = ~new_n11206 & ~new_n11207;
  assign new_n11209 = new_n11202 & ~new_n11208;
  assign new_n11210 = ~new_n11202 & new_n11208;
  assign new_n11211 = ~new_n11209 & ~new_n11210;
  assign new_n11212 = ~new_n11080 & new_n11211;
  assign new_n11213 = new_n11080 & ~new_n11211;
  assign new_n11214 = ~new_n11212 & ~new_n11213;
  assign new_n11215 = ~new_n11078 & new_n11214;
  assign new_n11216 = new_n11078 & ~new_n11214;
  assign new_n11217 = ~new_n11215 & ~new_n11216;
  assign new_n11218 = ~new_n10970 & ~new_n11217;
  assign new_n11219 = new_n10970 & new_n11217;
  assign n6683 = new_n11218 | new_n11219;
  assign new_n11221 = n7772 & n9528;
  assign new_n11222_1 = n7529 & n9669;
  assign new_n11223 = new_n10271 & ~new_n10274;
  assign new_n11224 = ~new_n10275 & ~new_n11223;
  assign new_n11225 = ~new_n11222_1 & new_n11224;
  assign new_n11226 = new_n11222_1 & ~new_n11224;
  assign new_n11227 = ~new_n11225 & ~new_n11226;
  assign new_n11228 = n8230 & n12853;
  assign new_n11229 = n7715 & n11891;
  assign new_n11230 = n2458 & n9531;
  assign new_n11231 = ~new_n11229 & ~new_n11230;
  assign new_n11232 = new_n11229 & new_n11230;
  assign new_n11233 = ~new_n11231 & ~new_n11232;
  assign new_n11234 = new_n11228 & ~new_n11233;
  assign new_n11235 = ~new_n11228 & new_n11233;
  assign new_n11236_1 = ~new_n11234 & ~new_n11235;
  assign new_n11237 = ~new_n11227 & new_n11236_1;
  assign new_n11238 = new_n11227 & ~new_n11236_1;
  assign new_n11239 = ~new_n11237 & ~new_n11238;
  assign new_n11240 = new_n11221 & new_n11239;
  assign new_n11241 = ~new_n11221 & ~new_n11239;
  assign new_n11242 = ~new_n10269 & new_n10279;
  assign new_n11243 = ~new_n10268 & ~new_n11242;
  assign new_n11244 = ~new_n11241 & new_n11243;
  assign new_n11245 = ~new_n11240 & ~new_n11244;
  assign new_n11246 = n7529 & n9528;
  assign new_n11247 = n7715 & n9669;
  assign new_n11248 = ~new_n11246 & ~new_n11247;
  assign new_n11249 = new_n11246 & new_n11247;
  assign new_n11250 = ~new_n11248 & ~new_n11249;
  assign new_n11251 = n2458 & n11891;
  assign new_n11252_1 = n8230 & n9531;
  assign new_n11253 = n6668 & n12853;
  assign new_n11254 = ~new_n11252_1 & ~new_n11253;
  assign new_n11255 = new_n11252_1 & new_n11253;
  assign new_n11256 = ~new_n11254 & ~new_n11255;
  assign new_n11257 = ~new_n11251 & ~new_n11256;
  assign new_n11258 = new_n11251 & new_n11256;
  assign new_n11259 = ~new_n11257 & ~new_n11258;
  assign new_n11260 = ~new_n11228 & ~new_n11232;
  assign new_n11261 = ~new_n11231 & ~new_n11260;
  assign new_n11262 = ~new_n11259 & ~new_n11261;
  assign new_n11263 = new_n11259 & new_n11261;
  assign new_n11264_1 = ~new_n11262 & ~new_n11263;
  assign new_n11265 = ~new_n11250 & ~new_n11264_1;
  assign new_n11266 = new_n11250 & new_n11264_1;
  assign new_n11267 = ~new_n11265 & ~new_n11266;
  assign new_n11268 = ~new_n11225 & ~new_n11236_1;
  assign new_n11269 = ~new_n11226 & ~new_n11268;
  assign new_n11270 = ~new_n11267 & ~new_n11269;
  assign new_n11271 = new_n11267 & new_n11269;
  assign new_n11272 = ~new_n11270 & ~new_n11271;
  assign new_n11273 = ~new_n11245 & ~new_n11272;
  assign new_n11274 = ~new_n11265 & ~new_n11269;
  assign new_n11275 = ~new_n11249 & ~new_n11274;
  assign new_n11276 = ~new_n11266 & new_n11275;
  assign new_n11277 = new_n11249 & new_n11274;
  assign new_n11278 = ~new_n11276 & ~new_n11277;
  assign new_n11279 = n7715 & n9528;
  assign new_n11280 = n7772 & n8522;
  assign new_n11281 = n6655 & n7529;
  assign new_n11282 = ~new_n11280 & ~new_n11281;
  assign new_n11283 = new_n11280 & new_n11281;
  assign new_n11284 = ~new_n11282 & ~new_n11283;
  assign new_n11285 = new_n11279 & ~new_n11284;
  assign new_n11286 = ~new_n11279 & new_n11284;
  assign new_n11287 = ~new_n11285 & ~new_n11286;
  assign new_n11288 = ~new_n11258 & ~new_n11261;
  assign new_n11289 = ~new_n11257 & ~new_n11288;
  assign new_n11290 = new_n11287 & ~new_n11289;
  assign new_n11291 = n2458 & n9669;
  assign new_n11292 = ~new_n11255 & ~new_n11291;
  assign new_n11293 = new_n11255 & new_n11291;
  assign new_n11294 = ~new_n11292 & ~new_n11293;
  assign new_n11295 = n7812 & n12853;
  assign new_n11296 = n6668 & n9531;
  assign new_n11297 = n8230 & n11891;
  assign new_n11298 = ~new_n11296 & ~new_n11297;
  assign new_n11299 = new_n11296 & new_n11297;
  assign new_n11300 = ~new_n11298 & ~new_n11299;
  assign new_n11301 = new_n11295 & ~new_n11300;
  assign new_n11302 = ~new_n11295 & new_n11300;
  assign new_n11303 = ~new_n11301 & ~new_n11302;
  assign new_n11304 = new_n11294 & new_n11303;
  assign new_n11305 = ~new_n11294 & ~new_n11303;
  assign new_n11306 = ~new_n11304 & ~new_n11305;
  assign new_n11307 = new_n11290 & new_n11306;
  assign new_n11308 = ~new_n11287 & new_n11289;
  assign new_n11309 = ~new_n11306 & new_n11308;
  assign new_n11310 = ~new_n11290 & ~new_n11306;
  assign new_n11311 = ~new_n11308 & ~new_n11310;
  assign new_n11312 = ~new_n11309 & ~new_n11311;
  assign new_n11313 = ~new_n11307 & ~new_n11312;
  assign new_n11314 = new_n11278 & ~new_n11313;
  assign new_n11315 = ~new_n11278 & new_n11313;
  assign new_n11316 = ~new_n11314 & ~new_n11315;
  assign new_n11317 = ~new_n11273 & new_n11316;
  assign new_n11318 = new_n11273 & ~new_n11316;
  assign new_n11319 = ~new_n11317 & ~new_n11318;
  assign new_n11320 = n6655 & n7772;
  assign new_n11321 = new_n11245 & new_n11272;
  assign new_n11322 = ~new_n11273 & ~new_n11321;
  assign new_n11323 = new_n11320 & new_n11322;
  assign new_n11324_1 = ~new_n11240 & ~new_n11241;
  assign new_n11325 = ~new_n11243 & ~new_n11324_1;
  assign new_n11326 = new_n11243 & new_n11324_1;
  assign new_n11327 = ~new_n11325 & ~new_n11326;
  assign new_n11328 = new_n10284 & new_n11327;
  assign new_n11329 = ~new_n11320 & ~new_n11322;
  assign new_n11330 = ~new_n11323 & ~new_n11329;
  assign new_n11331 = new_n11328 & new_n11330;
  assign new_n11332 = ~new_n11323 & ~new_n11331;
  assign new_n11333 = ~new_n11319 & new_n11332;
  assign new_n11334 = new_n11319 & ~new_n11332;
  assign new_n11335 = ~new_n11333 & ~new_n11334;
  assign new_n11336 = n11324 & new_n424;
  assign new_n11337 = n12348 & new_n11336;
  assign new_n11338 = ~n9216 & ~new_n11337;
  assign new_n11339 = ~new_n387 & new_n10333;
  assign new_n11340 = ~new_n11338 & ~new_n11339;
  assign new_n11341 = n854 & n8183;
  assign new_n11342 = ~new_n10333 & ~new_n11336;
  assign new_n11343 = ~n2068 & new_n387;
  assign new_n11344 = ~n12348 & new_n424;
  assign new_n11345 = ~new_n11343 & ~new_n11344;
  assign new_n11346 = ~new_n11342 & new_n11345;
  assign new_n11347 = ~new_n11341 & new_n11346;
  assign new_n11348 = new_n11341 & ~new_n11346;
  assign new_n11349 = ~new_n11347 & ~new_n11348;
  assign new_n11350_1 = new_n11340 & new_n11349;
  assign new_n11351 = n10142 & new_n11341;
  assign new_n11352 = ~n8183 & ~n10142;
  assign new_n11353 = n854 & ~new_n11352;
  assign new_n11354 = ~new_n11351 & new_n11353;
  assign new_n11355 = new_n10332 & new_n11354;
  assign new_n11356 = ~new_n10332 & ~new_n11354;
  assign new_n11357 = ~new_n11355 & ~new_n11356;
  assign new_n11358 = ~new_n11336 & ~new_n11341;
  assign new_n11359 = ~new_n10333 & ~new_n11358;
  assign new_n11360 = ~new_n11357 & new_n11359;
  assign new_n11361 = new_n11357 & ~new_n11359;
  assign new_n11362 = ~new_n11360 & ~new_n11361;
  assign new_n11363 = new_n424 & ~new_n11362;
  assign new_n11364 = ~new_n424 & new_n11362;
  assign new_n11365 = ~new_n11363 & ~new_n11364;
  assign new_n11366 = new_n10333 & ~new_n11341;
  assign new_n11367 = n12348 & ~new_n11366;
  assign new_n11368 = n8183 & new_n11336;
  assign new_n11369 = ~new_n11367 & ~new_n11368;
  assign new_n11370 = new_n11365 & new_n11369;
  assign new_n11371 = ~new_n11365 & ~new_n11369;
  assign new_n11372 = ~new_n11370 & ~new_n11371;
  assign new_n11373 = new_n11350_1 & ~new_n11372;
  assign new_n11374 = ~new_n11350_1 & new_n11372;
  assign new_n11375 = ~new_n11373 & ~new_n11374;
  assign new_n11376 = new_n384 & new_n11375;
  assign new_n11377 = ~new_n11340 & ~new_n11349;
  assign new_n11378 = ~new_n11350_1 & ~new_n11377;
  assign new_n11379 = new_n384 & new_n11337;
  assign new_n11380 = new_n11378 & new_n11379;
  assign new_n11381 = ~new_n11376 & ~new_n11380;
  assign new_n11382 = ~new_n11364 & ~new_n11369;
  assign new_n11383 = ~new_n11363 & ~new_n11382;
  assign new_n11384 = ~new_n10332 & ~new_n11351;
  assign new_n11385 = n11324 & new_n11351;
  assign new_n11386 = ~new_n11384 & ~new_n11385;
  assign new_n11387 = n854 & n10657;
  assign new_n11388 = ~new_n11354 & ~new_n11387;
  assign new_n11389 = new_n11354 & new_n11387;
  assign new_n11390 = ~new_n11388 & ~new_n11389;
  assign new_n11391 = ~new_n11386 & ~new_n11390;
  assign new_n11392 = new_n11386 & new_n11390;
  assign new_n11393 = ~new_n11391 & ~new_n11392;
  assign new_n11394 = new_n389_1 & new_n11393;
  assign new_n11395 = ~new_n389_1 & ~new_n11393;
  assign new_n11396_1 = ~new_n11394 & ~new_n11395;
  assign new_n11397 = ~new_n11355 & ~new_n11359;
  assign new_n11398 = ~new_n11356 & ~new_n11397;
  assign new_n11399 = new_n11396_1 & ~new_n11398;
  assign new_n11400 = ~new_n11396_1 & new_n11398;
  assign new_n11401 = ~new_n11399 & ~new_n11400;
  assign new_n11402 = ~new_n11383 & ~new_n11401;
  assign new_n11403 = new_n11383 & new_n11401;
  assign new_n11404 = ~new_n11402 & ~new_n11403;
  assign new_n11405 = new_n11373 & new_n11404;
  assign new_n11406 = ~new_n11373 & ~new_n11404;
  assign new_n11407 = ~new_n11405 & ~new_n11406;
  assign new_n11408 = ~new_n11381 & new_n11407;
  assign new_n11409 = new_n11381 & ~new_n11407;
  assign new_n11410 = ~new_n11408 & ~new_n11409;
  assign new_n11411_1 = n2295 & n12592;
  assign new_n11412 = n10168 & n13060;
  assign new_n11413 = ~new_n11411_1 & ~new_n11412;
  assign new_n11414 = new_n11411_1 & new_n11412;
  assign new_n11415 = ~new_n11413 & ~new_n11414;
  assign new_n11416 = n767 & n5189;
  assign new_n11417 = n8716 & n11537;
  assign new_n11418 = n834 & n951;
  assign new_n11419 = ~new_n11417 & ~new_n11418;
  assign new_n11420 = new_n11417 & new_n11418;
  assign new_n11421 = ~new_n11419 & ~new_n11420;
  assign new_n11422 = ~new_n11416 & ~new_n11421;
  assign new_n11423 = new_n11416 & new_n11421;
  assign new_n11424 = ~new_n11422 & ~new_n11423;
  assign new_n11425 = n5189 & n10168;
  assign new_n11426 = n767 & n8716;
  assign new_n11427 = new_n11425 & new_n11426;
  assign new_n11428 = n834 & n11537;
  assign new_n11429_1 = ~new_n11425 & ~new_n11426;
  assign new_n11430 = new_n11428 & ~new_n11429_1;
  assign new_n11431 = ~new_n11427 & ~new_n11430;
  assign new_n11432 = ~new_n11424 & new_n11431;
  assign new_n11433 = new_n11424 & ~new_n11431;
  assign new_n11434 = ~new_n11432 & ~new_n11433;
  assign new_n11435 = ~new_n11415 & ~new_n11434;
  assign new_n11436 = new_n11415 & new_n11434;
  assign new_n11437 = ~new_n11435 & ~new_n11436;
  assign new_n11438 = n12592 & n13060;
  assign new_n11439 = new_n10311 & ~new_n10314;
  assign new_n11440 = ~new_n10315 & ~new_n11439;
  assign new_n11441 = ~new_n11438 & new_n11440;
  assign new_n11442 = new_n11438 & ~new_n11440;
  assign new_n11443 = ~new_n11427 & ~new_n11429_1;
  assign new_n11444 = new_n11428 & ~new_n11443;
  assign new_n11445 = ~new_n11428 & new_n11443;
  assign new_n11446 = ~new_n11444 & ~new_n11445;
  assign new_n11447 = ~new_n11442 & new_n11446;
  assign new_n11448 = ~new_n11441 & ~new_n11447;
  assign new_n11449 = ~new_n11437 & ~new_n11448;
  assign new_n11450 = new_n11437 & new_n11448;
  assign new_n11451 = ~new_n11449 & ~new_n11450;
  assign new_n11452 = n2295 & n3178;
  assign new_n11453 = ~new_n11441 & ~new_n11442;
  assign new_n11454 = new_n11446 & ~new_n11453;
  assign new_n11455 = ~new_n11446 & new_n11453;
  assign new_n11456 = ~new_n11454 & ~new_n11455;
  assign new_n11457 = new_n11452 & new_n11456;
  assign new_n11458 = ~new_n11452 & ~new_n11456;
  assign new_n11459 = ~new_n10309 & new_n10319;
  assign new_n11460 = ~new_n10308 & ~new_n11459;
  assign new_n11461 = ~new_n11458 & new_n11460;
  assign new_n11462 = ~new_n11457 & ~new_n11461;
  assign new_n11463 = new_n11451 & ~new_n11462;
  assign new_n11464 = ~new_n11435 & new_n11448;
  assign new_n11465 = ~new_n11414 & ~new_n11464;
  assign new_n11466 = ~new_n11436 & new_n11465;
  assign new_n11467 = new_n11414 & new_n11464;
  assign new_n11468 = ~new_n11466 & ~new_n11467;
  assign new_n11469 = n2295 & n10168;
  assign new_n11470 = n2341 & n3178;
  assign new_n11471 = n1650 & n12592;
  assign new_n11472 = ~new_n11470 & ~new_n11471;
  assign new_n11473 = new_n11470 & new_n11471;
  assign new_n11474 = ~new_n11472 & ~new_n11473;
  assign new_n11475 = new_n11469 & ~new_n11474;
  assign new_n11476 = ~new_n11469 & new_n11474;
  assign new_n11477 = ~new_n11475 & ~new_n11476;
  assign new_n11478 = ~new_n11423 & new_n11431;
  assign new_n11479 = ~new_n11422 & ~new_n11478;
  assign new_n11480 = new_n11477 & ~new_n11479;
  assign new_n11481 = n767 & n13060;
  assign new_n11482 = new_n11420 & new_n11481;
  assign new_n11483 = ~new_n11420 & ~new_n11481;
  assign new_n11484_1 = ~new_n11482 & ~new_n11483;
  assign new_n11485 = n401 & n834;
  assign new_n11486 = n951 & n8716;
  assign new_n11487 = n5189 & n11537;
  assign new_n11488_1 = ~new_n11486 & ~new_n11487;
  assign new_n11489 = new_n11486 & new_n11487;
  assign new_n11490 = ~new_n11488_1 & ~new_n11489;
  assign new_n11491 = new_n11485 & ~new_n11490;
  assign new_n11492 = ~new_n11485 & new_n11490;
  assign new_n11493 = ~new_n11491 & ~new_n11492;
  assign new_n11494 = new_n11484_1 & new_n11493;
  assign new_n11495 = ~new_n11484_1 & ~new_n11493;
  assign new_n11496 = ~new_n11494 & ~new_n11495;
  assign new_n11497 = new_n11480 & new_n11496;
  assign new_n11498 = ~new_n11477 & new_n11479;
  assign new_n11499 = ~new_n11496 & new_n11498;
  assign new_n11500 = ~new_n11480 & ~new_n11496;
  assign new_n11501 = ~new_n11498 & ~new_n11500;
  assign new_n11502 = ~new_n11499 & ~new_n11501;
  assign new_n11503 = ~new_n11497 & ~new_n11502;
  assign new_n11504 = ~new_n11468 & ~new_n11503;
  assign new_n11505 = new_n11468 & new_n11503;
  assign new_n11506 = ~new_n11504 & ~new_n11505;
  assign new_n11507 = ~new_n11463 & ~new_n11506;
  assign new_n11508 = new_n11463 & new_n11506;
  assign new_n11509 = ~new_n11507 & ~new_n11508;
  assign new_n11510 = n1650 & n3178;
  assign new_n11511 = ~new_n11451 & new_n11462;
  assign new_n11512 = ~new_n11463 & ~new_n11511;
  assign new_n11513 = new_n11510 & new_n11512;
  assign new_n11514 = ~new_n11457 & ~new_n11458;
  assign new_n11515 = ~new_n11460 & ~new_n11514;
  assign new_n11516 = new_n11460 & new_n11514;
  assign new_n11517 = ~new_n11515 & ~new_n11516;
  assign new_n11518 = new_n10323 & new_n11517;
  assign new_n11519 = ~new_n11510 & ~new_n11512;
  assign new_n11520 = ~new_n11513 & ~new_n11519;
  assign new_n11521 = new_n11518 & new_n11520;
  assign new_n11522 = ~new_n11513 & ~new_n11521;
  assign new_n11523 = ~new_n11509 & new_n11522;
  assign new_n11524 = new_n11509 & ~new_n11522;
  assign new_n11525 = ~new_n11523 & ~new_n11524;
  assign new_n11526 = n8466 & n12579;
  assign new_n11527 = n8466 & n11222;
  assign new_n11528 = ~new_n10299 & ~new_n11527;
  assign new_n11529 = new_n10299 & new_n11527;
  assign new_n11530 = new_n10290 & ~new_n10293;
  assign new_n11531 = ~new_n10294 & ~new_n11530;
  assign new_n11532 = n510 & n2590;
  assign new_n11533 = n9 & n9591;
  assign new_n11534 = n2592 & n8290;
  assign new_n11535 = ~new_n11533 & ~new_n11534;
  assign new_n11536 = new_n11533 & new_n11534;
  assign new_n11537_1 = ~new_n11535 & ~new_n11536;
  assign new_n11538 = new_n11532 & ~new_n11537_1;
  assign new_n11539 = ~new_n11532 & new_n11537_1;
  assign new_n11540 = ~new_n11538 & ~new_n11539;
  assign new_n11541 = ~new_n11531 & ~new_n11540;
  assign new_n11542 = new_n11531 & new_n11540;
  assign new_n11543 = ~new_n11541 & ~new_n11542;
  assign new_n11544 = ~new_n11529 & ~new_n11543;
  assign new_n11545 = ~new_n11528 & ~new_n11544;
  assign new_n11546 = n5031 & n11222;
  assign new_n11547 = new_n11541 & new_n11546;
  assign new_n11548 = ~new_n11541 & ~new_n11546;
  assign new_n11549 = ~new_n11547 & ~new_n11548;
  assign new_n11550 = n2592 & n9591;
  assign new_n11551 = n510 & n11061;
  assign new_n11552 = n2590 & n8290;
  assign new_n11553 = ~new_n11551 & ~new_n11552;
  assign new_n11554 = new_n11551 & new_n11552;
  assign new_n11555 = ~new_n11553 & ~new_n11554;
  assign new_n11556 = new_n11550 & new_n11555;
  assign new_n11557 = ~new_n11550 & ~new_n11555;
  assign new_n11558 = ~new_n11556 & ~new_n11557;
  assign new_n11559 = new_n11532 & ~new_n11535;
  assign new_n11560 = ~new_n11536 & ~new_n11559;
  assign new_n11561 = ~new_n11558 & new_n11560;
  assign new_n11562 = new_n11558 & ~new_n11560;
  assign new_n11563 = ~new_n11561 & ~new_n11562;
  assign new_n11564 = ~new_n11549 & new_n11563;
  assign new_n11565 = new_n11549 & ~new_n11563;
  assign new_n11566 = ~new_n11564 & ~new_n11565;
  assign new_n11567 = ~new_n11545 & new_n11566;
  assign new_n11568 = new_n11545 & ~new_n11566;
  assign new_n11569 = ~new_n11567 & ~new_n11568;
  assign new_n11570 = new_n11526 & new_n11569;
  assign new_n11571 = ~new_n11528 & ~new_n11529;
  assign new_n11572 = new_n11543 & ~new_n11571;
  assign new_n11573 = ~new_n11543 & new_n11571;
  assign new_n11574_1 = ~new_n11572 & ~new_n11573;
  assign new_n11575 = new_n10303 & ~new_n11574_1;
  assign new_n11576 = ~new_n11526 & ~new_n11569;
  assign new_n11577 = ~new_n11570 & ~new_n11576;
  assign new_n11578 = new_n11575 & new_n11577;
  assign new_n11579 = ~new_n11570 & ~new_n11578;
  assign new_n11580 = n510 & n8768;
  assign new_n11581 = n8290 & n11061;
  assign new_n11582 = n2590 & n9591;
  assign new_n11583 = ~new_n11581 & ~new_n11582;
  assign new_n11584 = new_n11581 & new_n11582;
  assign new_n11585 = ~new_n11583 & ~new_n11584;
  assign new_n11586 = new_n11580 & ~new_n11585;
  assign new_n11587 = ~new_n11580 & new_n11585;
  assign new_n11588 = ~new_n11586 & ~new_n11587;
  assign new_n11589 = ~new_n11554 & new_n11588;
  assign new_n11590 = new_n11554 & ~new_n11588;
  assign new_n11591 = ~new_n11589 & ~new_n11590;
  assign new_n11592 = n9 & n11222;
  assign new_n11593 = n6023 & n8466;
  assign new_n11594 = n5031 & n12579;
  assign new_n11595 = ~new_n11593 & ~new_n11594;
  assign new_n11596 = new_n11593 & new_n11594;
  assign new_n11597 = ~new_n11595 & ~new_n11596;
  assign new_n11598 = new_n11592 & ~new_n11597;
  assign new_n11599 = ~new_n11592 & new_n11597;
  assign new_n11600 = ~new_n11598 & ~new_n11599;
  assign new_n11601 = ~new_n11556 & new_n11560;
  assign new_n11602 = ~new_n11557 & ~new_n11601;
  assign new_n11603 = ~new_n11600 & new_n11602;
  assign new_n11604 = new_n11600 & ~new_n11602;
  assign new_n11605 = ~new_n11603 & ~new_n11604;
  assign new_n11606 = new_n11591 & new_n11605;
  assign new_n11607 = ~new_n11591 & ~new_n11605;
  assign new_n11608 = ~new_n11606 & ~new_n11607;
  assign new_n11609 = ~new_n11547 & ~new_n11563;
  assign new_n11610 = ~new_n11548 & ~new_n11609;
  assign new_n11611 = ~new_n11608 & ~new_n11610;
  assign new_n11612 = new_n11608 & new_n11610;
  assign new_n11613 = ~new_n11611 & ~new_n11612;
  assign new_n11614 = new_n11568 & new_n11613;
  assign new_n11615 = ~new_n11568 & ~new_n11613;
  assign new_n11616 = ~new_n11614 & ~new_n11615;
  assign new_n11617 = ~new_n11579 & new_n11616;
  assign new_n11618 = new_n11579 & ~new_n11616;
  assign new_n11619 = ~new_n11617 & ~new_n11618;
  assign new_n11620 = ~new_n11525 & ~new_n11619;
  assign new_n11621 = new_n11525 & new_n11619;
  assign new_n11622 = ~new_n11620 & ~new_n11621;
  assign new_n11623 = ~new_n11575 & ~new_n11577;
  assign new_n11624 = ~new_n11578 & ~new_n11623;
  assign new_n11625 = ~new_n11518 & ~new_n11520;
  assign new_n11626 = ~new_n11521 & ~new_n11625;
  assign new_n11627 = ~new_n11624 & ~new_n11626;
  assign new_n11628 = new_n11624 & new_n11626;
  assign new_n11629 = ~new_n10323 & ~new_n11517;
  assign new_n11630 = ~new_n11518 & ~new_n11629;
  assign new_n11631 = ~new_n10303 & new_n11574_1;
  assign new_n11632 = ~new_n11575 & ~new_n11631;
  assign new_n11633 = ~new_n11630 & ~new_n11632;
  assign new_n11634_1 = new_n11630 & new_n11632;
  assign new_n11635 = ~new_n10287 & ~new_n10326;
  assign new_n11636 = ~new_n10327 & ~new_n11635;
  assign new_n11637 = ~new_n11634_1 & ~new_n11636;
  assign new_n11638 = ~new_n11633 & ~new_n11637;
  assign new_n11639 = ~new_n11628 & ~new_n11638;
  assign new_n11640 = ~new_n11627 & ~new_n11639;
  assign new_n11641 = ~new_n11622 & ~new_n11640;
  assign new_n11642 = new_n11622 & new_n11640;
  assign new_n11643 = ~new_n11641 & ~new_n11642;
  assign new_n11644 = new_n11410 & new_n11643;
  assign new_n11645 = ~new_n11410 & ~new_n11643;
  assign new_n11646 = ~new_n11644 & ~new_n11645;
  assign new_n11647 = new_n384 & ~new_n11380;
  assign new_n11648 = new_n11375 & ~new_n11647;
  assign new_n11649 = ~new_n11375 & new_n11647;
  assign new_n11650 = ~new_n11648 & ~new_n11649;
  assign new_n11651 = ~new_n11378 & ~new_n11379;
  assign new_n11652 = ~new_n11380 & ~new_n11651;
  assign new_n11653 = ~new_n11633 & ~new_n11634_1;
  assign new_n11654 = ~new_n11636 & ~new_n11653;
  assign new_n11655 = new_n11636 & new_n11653;
  assign new_n11656 = ~new_n11654 & ~new_n11655;
  assign new_n11657 = new_n11652 & new_n11656;
  assign new_n11658 = ~new_n11652 & ~new_n11656;
  assign new_n11659 = ~new_n10337 & ~new_n10341;
  assign new_n11660 = ~new_n10338 & ~new_n11659;
  assign new_n11661 = ~new_n11658 & ~new_n11660;
  assign new_n11662 = ~new_n11657 & ~new_n11661;
  assign new_n11663 = ~new_n11650 & ~new_n11662;
  assign new_n11664 = new_n11650 & new_n11662;
  assign new_n11665_1 = ~new_n11627 & ~new_n11628;
  assign new_n11666 = ~new_n11638 & new_n11665_1;
  assign new_n11667_1 = new_n11638 & ~new_n11665_1;
  assign new_n11668 = ~new_n11666 & ~new_n11667_1;
  assign new_n11669 = ~new_n11664 & ~new_n11668;
  assign new_n11670 = ~new_n11663 & ~new_n11669;
  assign new_n11671 = new_n11646 & new_n11670;
  assign new_n11672 = ~new_n11646 & ~new_n11670;
  assign new_n11673 = ~new_n11671 & ~new_n11672;
  assign new_n11674 = new_n11335 & ~new_n11673;
  assign new_n11675 = ~new_n11335 & new_n11673;
  assign new_n11676 = ~new_n11674 & ~new_n11675;
  assign new_n11677 = ~new_n11328 & ~new_n11330;
  assign new_n11678 = ~new_n11331 & ~new_n11677;
  assign new_n11679 = ~new_n11663 & ~new_n11664;
  assign new_n11680 = ~new_n11668 & new_n11679;
  assign new_n11681 = new_n11668 & ~new_n11679;
  assign new_n11682 = ~new_n11680 & ~new_n11681;
  assign new_n11683 = ~new_n11678 & ~new_n11682;
  assign new_n11684 = new_n11678 & new_n11682;
  assign new_n11685 = ~new_n10284 & ~new_n11327;
  assign new_n11686 = ~new_n11328 & ~new_n11685;
  assign new_n11687 = ~new_n11657 & ~new_n11658;
  assign new_n11688 = new_n11660 & ~new_n11687;
  assign new_n11689 = ~new_n11660 & new_n11687;
  assign new_n11690 = ~new_n11688 & ~new_n11689;
  assign new_n11691 = ~new_n11686 & ~new_n11690;
  assign new_n11692 = new_n11686 & new_n11690;
  assign new_n11693 = ~new_n10346 & ~new_n10349;
  assign new_n11694 = ~new_n10345 & ~new_n11693;
  assign new_n11695 = ~new_n11692 & new_n11694;
  assign new_n11696 = ~new_n11691 & ~new_n11695;
  assign new_n11697 = ~new_n11684 & ~new_n11696;
  assign new_n11698 = ~new_n11683 & ~new_n11697;
  assign new_n11699 = ~new_n11676 & new_n11698;
  assign new_n11700 = new_n11676 & ~new_n11698;
  assign n6862 = new_n11699 | new_n11700;
  assign new_n11702 = n8468 & n9216;
  assign new_n11703 = n11109 & n12348;
  assign new_n11704 = new_n10136 & ~new_n10139;
  assign new_n11705 = ~new_n10140 & ~new_n11704;
  assign new_n11706 = ~new_n11703 & new_n11705;
  assign new_n11707 = new_n11703 & ~new_n11705;
  assign new_n11708 = ~new_n11706 & ~new_n11707;
  assign new_n11709 = n2068 & n9906;
  assign new_n11710 = n6085 & n11324;
  assign new_n11711 = n5962 & n8183;
  assign new_n11712 = ~new_n11710 & ~new_n11711;
  assign new_n11713 = new_n11710 & new_n11711;
  assign new_n11714 = ~new_n11712 & ~new_n11713;
  assign new_n11715 = new_n11709 & ~new_n11714;
  assign new_n11716 = ~new_n11709 & new_n11714;
  assign new_n11717 = ~new_n11715 & ~new_n11716;
  assign new_n11718 = ~new_n11708 & new_n11717;
  assign new_n11719 = new_n11708 & ~new_n11717;
  assign new_n11720 = ~new_n11718 & ~new_n11719;
  assign new_n11721 = ~new_n11702 & ~new_n11720;
  assign new_n11722 = new_n11702 & new_n11720;
  assign new_n11723 = ~new_n10133 & ~new_n10144;
  assign new_n11724 = ~new_n10134 & ~new_n11723;
  assign new_n11725 = ~new_n11722 & new_n11724;
  assign new_n11726 = ~new_n11721 & ~new_n11725;
  assign new_n11727 = n2068 & n11109;
  assign new_n11728 = n8468 & n12348;
  assign new_n11729 = ~new_n11727 & ~new_n11728;
  assign new_n11730 = new_n11727 & new_n11728;
  assign new_n11731 = ~new_n11729 & ~new_n11730;
  assign new_n11732_1 = n9906 & n11324;
  assign new_n11733 = n6085 & n8183;
  assign new_n11734_1 = n5962 & n10142;
  assign new_n11735 = ~new_n11733 & ~new_n11734_1;
  assign new_n11736 = new_n11733 & new_n11734_1;
  assign new_n11737 = ~new_n11735 & ~new_n11736;
  assign new_n11738 = ~new_n11732_1 & ~new_n11737;
  assign new_n11739 = new_n11732_1 & new_n11737;
  assign new_n11740 = ~new_n11738 & ~new_n11739;
  assign new_n11741 = new_n11709 & ~new_n11712;
  assign new_n11742 = ~new_n11713 & ~new_n11741;
  assign new_n11743 = ~new_n11740 & ~new_n11742;
  assign new_n11744 = new_n11740 & new_n11742;
  assign new_n11745 = ~new_n11743 & ~new_n11744;
  assign new_n11746 = ~new_n11731 & new_n11745;
  assign new_n11747 = new_n11731 & ~new_n11745;
  assign new_n11748 = ~new_n11746 & ~new_n11747;
  assign new_n11749 = ~new_n11706 & ~new_n11717;
  assign new_n11750 = ~new_n11707 & ~new_n11749;
  assign new_n11751 = ~new_n11748 & new_n11750;
  assign new_n11752 = new_n11748 & ~new_n11750;
  assign new_n11753 = ~new_n11751 & ~new_n11752;
  assign new_n11754 = new_n11726 & new_n11753;
  assign new_n11755 = ~new_n11746 & ~new_n11750;
  assign new_n11756 = ~new_n11730 & ~new_n11755;
  assign new_n11757 = ~new_n11747 & new_n11756;
  assign new_n11758 = new_n11730 & new_n11755;
  assign new_n11759 = ~new_n11757 & ~new_n11758;
  assign new_n11760 = n1084 & n9216;
  assign new_n11761 = n2068 & n8468;
  assign new_n11762 = n6818 & n12348;
  assign new_n11763 = ~new_n11761 & ~new_n11762;
  assign new_n11764 = new_n11761 & new_n11762;
  assign new_n11765 = ~new_n11763 & ~new_n11764;
  assign new_n11766 = new_n11760 & ~new_n11765;
  assign new_n11767 = ~new_n11760 & new_n11765;
  assign new_n11768 = ~new_n11766 & ~new_n11767;
  assign new_n11769 = ~new_n11739 & new_n11742;
  assign new_n11770 = ~new_n11738 & ~new_n11769;
  assign new_n11771 = new_n11768 & ~new_n11770;
  assign new_n11772 = ~new_n11768 & new_n11770;
  assign new_n11773 = ~new_n11771 & ~new_n11772;
  assign new_n11774 = n11109 & n11324;
  assign new_n11775 = new_n11736 & new_n11774;
  assign new_n11776 = ~new_n11736 & ~new_n11774;
  assign new_n11777 = ~new_n11775 & ~new_n11776;
  assign new_n11778_1 = n8183 & n9906;
  assign new_n11779 = n6085 & n10142;
  assign new_n11780 = n5962 & n10657;
  assign new_n11781 = ~new_n11779 & ~new_n11780;
  assign new_n11782 = new_n11779 & new_n11780;
  assign new_n11783 = ~new_n11781 & ~new_n11782;
  assign new_n11784 = new_n11778_1 & ~new_n11783;
  assign new_n11785 = ~new_n11778_1 & new_n11783;
  assign new_n11786 = ~new_n11784 & ~new_n11785;
  assign new_n11787 = new_n11777 & new_n11786;
  assign new_n11788 = ~new_n11777 & ~new_n11786;
  assign new_n11789 = ~new_n11787 & ~new_n11788;
  assign new_n11790 = new_n11773 & new_n11789;
  assign new_n11791 = ~new_n11773 & ~new_n11789;
  assign new_n11792_1 = ~new_n11790 & ~new_n11791;
  assign new_n11793 = new_n11759 & new_n11792_1;
  assign new_n11794 = ~new_n11759 & ~new_n11792_1;
  assign new_n11795 = ~new_n11793 & ~new_n11794;
  assign new_n11796 = new_n11754 & ~new_n11795;
  assign new_n11797 = ~new_n11754 & new_n11795;
  assign new_n11798 = ~new_n11796 & ~new_n11797;
  assign new_n11799 = n6818 & n9216;
  assign new_n11800 = ~new_n11726 & ~new_n11753;
  assign new_n11801 = ~new_n11754 & ~new_n11800;
  assign new_n11802 = new_n11799 & new_n11801;
  assign new_n11803 = ~new_n11721 & ~new_n11722;
  assign new_n11804 = ~new_n11724 & ~new_n11803;
  assign new_n11805 = new_n11724 & new_n11803;
  assign new_n11806 = ~new_n11804 & ~new_n11805;
  assign new_n11807 = new_n10149 & ~new_n11806;
  assign new_n11808 = ~new_n11799 & ~new_n11801;
  assign new_n11809 = ~new_n11802 & ~new_n11808;
  assign new_n11810 = new_n11807 & new_n11809;
  assign new_n11811 = ~new_n11802 & ~new_n11810;
  assign new_n11812 = new_n11798 & ~new_n11811;
  assign new_n11813 = ~new_n11798 & new_n11811;
  assign new_n11814 = ~new_n11812 & ~new_n11813;
  assign new_n11815 = n3178 & n9300;
  assign new_n11816 = n1198 & n12592;
  assign new_n11817 = n2498 & n10168;
  assign new_n11818 = new_n11816 & new_n11817;
  assign new_n11819 = ~new_n11816 & ~new_n11817;
  assign new_n11820 = ~new_n11818 & ~new_n11819;
  assign new_n11821 = n767 & n5969;
  assign new_n11822 = n951 & n11058;
  assign new_n11823 = n1007 & n11537;
  assign new_n11824 = ~new_n11822 & ~new_n11823;
  assign new_n11825 = new_n11822 & new_n11823;
  assign new_n11826 = ~new_n11824 & ~new_n11825;
  assign new_n11827 = ~new_n11821 & ~new_n11826;
  assign new_n11828 = new_n11821 & new_n11826;
  assign new_n11829 = ~new_n11827 & ~new_n11828;
  assign new_n11830 = n5969 & n11537;
  assign new_n11831 = new_n10184 & new_n11830;
  assign new_n11832 = n767 & n1007;
  assign new_n11833 = n11058 & n11537;
  assign new_n11834 = n5969 & n10168;
  assign new_n11835_1 = ~new_n11833 & ~new_n11834;
  assign new_n11836 = new_n11832 & ~new_n11835_1;
  assign new_n11837 = ~new_n11831 & ~new_n11836;
  assign new_n11838 = ~new_n11829 & new_n11837;
  assign new_n11839 = new_n11829 & ~new_n11837;
  assign new_n11840 = ~new_n11838 & ~new_n11839;
  assign new_n11841 = ~new_n11820 & ~new_n11840;
  assign new_n11842 = new_n11820 & new_n11840;
  assign new_n11843 = ~new_n11841 & ~new_n11842;
  assign new_n11844 = n2498 & n12592;
  assign new_n11845 = new_n10198 & ~new_n10201;
  assign new_n11846 = ~new_n10202 & ~new_n11845;
  assign new_n11847 = ~new_n11844 & new_n11846;
  assign new_n11848 = new_n11844 & ~new_n11846;
  assign new_n11849 = ~new_n11831 & ~new_n11835_1;
  assign new_n11850 = ~new_n11832 & ~new_n11849;
  assign new_n11851 = new_n11832 & new_n11849;
  assign new_n11852 = ~new_n11850 & ~new_n11851;
  assign new_n11853 = ~new_n11848 & ~new_n11852;
  assign new_n11854 = ~new_n11847 & ~new_n11853;
  assign new_n11855 = ~new_n11843 & new_n11854;
  assign new_n11856 = new_n11843 & ~new_n11854;
  assign new_n11857 = ~new_n11855 & ~new_n11856;
  assign new_n11858 = n1198 & n3178;
  assign new_n11859 = ~new_n11847 & ~new_n11848;
  assign new_n11860 = ~new_n11852 & new_n11859;
  assign new_n11861 = new_n11852 & ~new_n11859;
  assign new_n11862 = ~new_n11860 & ~new_n11861;
  assign new_n11863 = new_n11858 & ~new_n11862;
  assign new_n11864 = ~new_n11858 & new_n11862;
  assign new_n11865 = ~new_n10195 & ~new_n10206;
  assign new_n11866 = ~new_n10196 & ~new_n11865;
  assign new_n11867 = ~new_n11864 & ~new_n11866;
  assign new_n11868 = ~new_n11863 & ~new_n11867;
  assign new_n11869 = ~new_n11857 & ~new_n11868;
  assign new_n11870 = new_n11857 & new_n11868;
  assign new_n11871 = ~new_n11869 & ~new_n11870;
  assign new_n11872 = new_n11815 & new_n11871;
  assign new_n11873 = ~new_n11863 & ~new_n11864;
  assign new_n11874 = ~new_n11866 & ~new_n11873;
  assign new_n11875 = new_n11866 & new_n11873;
  assign new_n11876 = ~new_n11874 & ~new_n11875;
  assign new_n11877 = new_n10210 & ~new_n11876;
  assign new_n11878 = ~new_n11815 & ~new_n11871;
  assign new_n11879_1 = ~new_n11872 & ~new_n11878;
  assign new_n11880 = new_n11877 & new_n11879_1;
  assign new_n11881 = ~new_n11872 & ~new_n11880;
  assign new_n11882_1 = n3178 & n11574;
  assign new_n11883 = n1198 & n10168;
  assign new_n11884 = n9300 & n12592;
  assign new_n11885 = ~new_n11883 & ~new_n11884;
  assign new_n11886 = n9300 & n10168;
  assign new_n11887 = new_n11816 & new_n11886;
  assign new_n11888 = ~new_n11885 & ~new_n11887;
  assign new_n11889 = ~new_n11882_1 & ~new_n11888;
  assign new_n11890 = new_n11882_1 & new_n11888;
  assign new_n11891_1 = ~new_n11889 & ~new_n11890;
  assign new_n11892 = ~new_n11828 & new_n11837;
  assign new_n11893 = ~new_n11827 & ~new_n11892;
  assign new_n11894 = ~new_n11891_1 & ~new_n11893;
  assign new_n11895_1 = new_n11891_1 & new_n11893;
  assign new_n11896 = ~new_n11894 & ~new_n11895_1;
  assign new_n11897 = n767 & n2498;
  assign new_n11898 = ~new_n11825 & ~new_n11897;
  assign new_n11899 = new_n11825 & new_n11897;
  assign new_n11900 = ~new_n11898 & ~new_n11899;
  assign new_n11901 = n951 & n1007;
  assign new_n11902 = n401 & n11058;
  assign new_n11903 = ~new_n11901 & ~new_n11902;
  assign new_n11904 = new_n11901 & new_n11902;
  assign new_n11905 = ~new_n11903 & ~new_n11904;
  assign new_n11906 = new_n11830 & ~new_n11905;
  assign new_n11907 = ~new_n11830 & new_n11905;
  assign new_n11908 = ~new_n11906 & ~new_n11907;
  assign new_n11909 = new_n11900 & new_n11908;
  assign new_n11910 = ~new_n11900 & ~new_n11908;
  assign new_n11911 = ~new_n11909 & ~new_n11910;
  assign new_n11912 = ~new_n11896 & new_n11911;
  assign new_n11913 = new_n11896 & ~new_n11911;
  assign new_n11914 = ~new_n11912 & ~new_n11913;
  assign new_n11915 = ~new_n11841 & new_n11854;
  assign new_n11916 = ~new_n11818 & ~new_n11915;
  assign new_n11917 = ~new_n11842 & new_n11916;
  assign new_n11918 = new_n11818 & new_n11915;
  assign new_n11919 = ~new_n11917 & ~new_n11918;
  assign new_n11920 = new_n11914 & new_n11919;
  assign new_n11921 = ~new_n11914 & ~new_n11919;
  assign new_n11922 = ~new_n11920 & ~new_n11921;
  assign new_n11923 = new_n11869 & new_n11922;
  assign new_n11924 = ~new_n11869 & ~new_n11922;
  assign new_n11925 = ~new_n11923 & ~new_n11924;
  assign new_n11926 = ~new_n11881 & new_n11925;
  assign new_n11927 = new_n11881 & ~new_n11925;
  assign new_n11928 = ~new_n11926 & ~new_n11927;
  assign new_n11929 = n2339 & n5031;
  assign new_n11930 = n9 & n9570;
  assign new_n11931 = ~new_n11929 & ~new_n11930;
  assign new_n11932 = new_n11929 & new_n11930;
  assign new_n11933 = ~new_n11931 & ~new_n11932;
  assign new_n11934 = n2592 & n12482;
  assign new_n11935 = n2590 & n7720;
  assign new_n11936 = n287 & n11061;
  assign new_n11937 = ~new_n11935 & ~new_n11936;
  assign new_n11938 = new_n11935 & new_n11936;
  assign new_n11939 = ~new_n11937 & ~new_n11938;
  assign new_n11940 = ~new_n11934 & ~new_n11939;
  assign new_n11941 = new_n11934 & new_n11939;
  assign new_n11942 = ~new_n11940 & ~new_n11941;
  assign new_n11943 = new_n10169 & new_n11935;
  assign new_n11944 = n9 & n12482;
  assign new_n11945 = n2592 & n7720;
  assign new_n11946 = n287 & n2590;
  assign new_n11947 = ~new_n11945 & ~new_n11946;
  assign new_n11948 = new_n11944 & ~new_n11947;
  assign new_n11949 = ~new_n11943 & ~new_n11948;
  assign new_n11950 = ~new_n11942 & new_n11949;
  assign new_n11951 = new_n11942 & ~new_n11949;
  assign new_n11952 = ~new_n11950 & ~new_n11951;
  assign new_n11953 = ~new_n11933 & ~new_n11952;
  assign new_n11954 = new_n11933 & new_n11952;
  assign new_n11955 = ~new_n11953 & ~new_n11954;
  assign new_n11956 = n5031 & n9570;
  assign new_n11957 = new_n10167 & ~new_n10170;
  assign new_n11958 = ~new_n10171 & ~new_n11957;
  assign new_n11959 = ~new_n11956 & new_n11958;
  assign new_n11960 = new_n11956 & ~new_n11958;
  assign new_n11961 = ~new_n11943 & ~new_n11947;
  assign new_n11962 = ~new_n11944 & ~new_n11961;
  assign new_n11963 = new_n11944 & new_n11961;
  assign new_n11964 = ~new_n11962 & ~new_n11963;
  assign new_n11965 = ~new_n11960 & ~new_n11964;
  assign new_n11966 = ~new_n11959 & ~new_n11965;
  assign new_n11967 = ~new_n11955 & ~new_n11966;
  assign new_n11968 = new_n11955 & new_n11966;
  assign new_n11969 = ~new_n11967 & ~new_n11968;
  assign new_n11970 = n2339 & n8466;
  assign new_n11971 = ~new_n11959 & new_n11965;
  assign new_n11972 = ~new_n11959 & ~new_n11960;
  assign new_n11973 = new_n11964 & ~new_n11972;
  assign new_n11974 = ~new_n11971 & ~new_n11973;
  assign new_n11975 = new_n11970 & ~new_n11974;
  assign new_n11976 = ~new_n11970 & new_n11974;
  assign new_n11977 = ~new_n10164 & ~new_n10175;
  assign new_n11978 = ~new_n10165 & ~new_n11977;
  assign new_n11979 = ~new_n11976 & ~new_n11978;
  assign new_n11980 = ~new_n11975 & ~new_n11979;
  assign new_n11981 = new_n11969 & ~new_n11980;
  assign new_n11982 = ~new_n11953 & new_n11966;
  assign new_n11983 = ~new_n11932 & ~new_n11982;
  assign new_n11984 = ~new_n11954 & new_n11983;
  assign new_n11985 = new_n11932 & new_n11982;
  assign new_n11986 = ~new_n11984 & ~new_n11985;
  assign new_n11987 = n9 & n2339;
  assign new_n11988 = n1307 & n5031;
  assign new_n11989 = ~new_n11987 & ~new_n11988;
  assign new_n11990 = new_n11987 & new_n11988;
  assign new_n11991 = ~new_n11989 & ~new_n11990;
  assign new_n11992 = ~new_n11941 & new_n11949;
  assign new_n11993 = ~new_n11940 & ~new_n11992;
  assign new_n11994 = new_n11991 & new_n11993;
  assign new_n11995 = ~new_n11991 & ~new_n11993;
  assign new_n11996 = ~new_n11994 & ~new_n11995;
  assign new_n11997 = n2590 & n12482;
  assign new_n11998 = n7720 & n11061;
  assign new_n11999 = n287 & n8768;
  assign new_n12000 = ~new_n11998 & ~new_n11999;
  assign new_n12001 = n7720 & n8768;
  assign new_n12002 = new_n11936 & new_n12001;
  assign new_n12003_1 = ~new_n12000 & ~new_n12002;
  assign new_n12004 = ~new_n11997 & ~new_n12003_1;
  assign new_n12005 = new_n11997 & new_n12003_1;
  assign new_n12006 = ~new_n12004 & ~new_n12005;
  assign new_n12007 = n2592 & n9570;
  assign new_n12008 = ~new_n11938 & ~new_n12007;
  assign new_n12009 = new_n11938 & new_n12007;
  assign new_n12010 = ~new_n12008 & ~new_n12009;
  assign new_n12011 = ~new_n12006 & new_n12010;
  assign new_n12012 = new_n12006 & ~new_n12010;
  assign new_n12013 = ~new_n12011 & ~new_n12012;
  assign new_n12014 = ~new_n11996 & ~new_n12013;
  assign new_n12015 = new_n11996 & new_n12013;
  assign new_n12016 = ~new_n12014 & ~new_n12015;
  assign new_n12017 = ~new_n11986 & new_n12016;
  assign new_n12018 = new_n11986 & ~new_n12016;
  assign new_n12019 = ~new_n12017 & ~new_n12018;
  assign new_n12020 = new_n11981 & new_n12019;
  assign new_n12021 = ~new_n11981 & ~new_n12019;
  assign new_n12022 = ~new_n12020 & ~new_n12021;
  assign new_n12023 = n1307 & n8466;
  assign new_n12024 = ~new_n11969 & new_n11980;
  assign new_n12025 = ~new_n11981 & ~new_n12024;
  assign new_n12026 = new_n12023 & new_n12025;
  assign new_n12027 = ~new_n11975 & ~new_n11976;
  assign new_n12028 = ~new_n11978 & ~new_n12027;
  assign new_n12029 = new_n11978 & new_n12027;
  assign new_n12030 = ~new_n12028 & ~new_n12029;
  assign new_n12031 = new_n10180 & ~new_n12030;
  assign new_n12032 = ~new_n12023 & ~new_n12025;
  assign new_n12033 = ~new_n12026 & ~new_n12032;
  assign new_n12034 = new_n12031 & new_n12033;
  assign new_n12035 = ~new_n12026 & ~new_n12034;
  assign new_n12036 = new_n12022 & ~new_n12035;
  assign new_n12037 = ~new_n12022 & new_n12035;
  assign new_n12038 = ~new_n12036 & ~new_n12037;
  assign new_n12039 = ~new_n11928 & ~new_n12038;
  assign new_n12040 = ~new_n12031 & ~new_n12033;
  assign new_n12041 = ~new_n12034 & ~new_n12040;
  assign new_n12042 = ~new_n11877 & ~new_n11879_1;
  assign new_n12043 = ~new_n11880 & ~new_n12042;
  assign new_n12044 = new_n12041 & new_n12043;
  assign new_n12045 = ~new_n12041 & ~new_n12043;
  assign new_n12046 = ~new_n10210 & new_n11876;
  assign new_n12047 = ~new_n11877 & ~new_n12046;
  assign new_n12048 = ~new_n10180 & new_n12030;
  assign new_n12049 = ~new_n12031 & ~new_n12048;
  assign new_n12050 = new_n12047 & new_n12049;
  assign new_n12051 = ~new_n12047 & ~new_n12049;
  assign new_n12052 = ~new_n10214 & ~new_n10225;
  assign new_n12053 = ~new_n10213 & ~new_n12052;
  assign new_n12054 = ~new_n12051 & ~new_n12053;
  assign new_n12055 = ~new_n12050 & ~new_n12054;
  assign new_n12056 = ~new_n12045 & ~new_n12055;
  assign new_n12057 = ~new_n12044 & ~new_n12056;
  assign new_n12058 = new_n12039 & new_n12057;
  assign new_n12059_1 = new_n11928 & new_n12038;
  assign new_n12060 = new_n12057 & ~new_n12059_1;
  assign new_n12061 = ~new_n12039 & ~new_n12060;
  assign new_n12062 = ~new_n12058 & ~new_n12061;
  assign new_n12063 = ~new_n12057 & new_n12059_1;
  assign new_n12064 = ~new_n12062 & ~new_n12063;
  assign new_n12065_1 = new_n11814 & ~new_n12064;
  assign new_n12066 = ~new_n11814 & new_n12064;
  assign new_n12067_1 = ~new_n11807 & ~new_n11809;
  assign new_n12068 = ~new_n11810 & ~new_n12067_1;
  assign new_n12069 = ~new_n12044 & ~new_n12045;
  assign new_n12070 = new_n12055 & ~new_n12069;
  assign new_n12071 = ~new_n12055 & new_n12069;
  assign new_n12072 = ~new_n12070 & ~new_n12071;
  assign new_n12073 = new_n12068 & new_n12072;
  assign new_n12074 = ~new_n12068 & ~new_n12072;
  assign new_n12075 = ~new_n10149 & new_n11806;
  assign new_n12076 = ~new_n11807 & ~new_n12075;
  assign new_n12077 = ~new_n12050 & ~new_n12051;
  assign new_n12078 = new_n12053 & ~new_n12077;
  assign new_n12079 = ~new_n12053 & new_n12077;
  assign new_n12080 = ~new_n12078 & ~new_n12079;
  assign new_n12081 = new_n12076 & new_n12080;
  assign new_n12082 = ~new_n12076 & ~new_n12080;
  assign new_n12083 = ~new_n10230 & ~new_n10243_1;
  assign new_n12084 = ~new_n10229 & ~new_n12083;
  assign new_n12085 = ~new_n12082 & ~new_n12084;
  assign new_n12086 = ~new_n12081 & ~new_n12085;
  assign new_n12087 = ~new_n12074 & ~new_n12086;
  assign new_n12088 = ~new_n12073 & ~new_n12087;
  assign new_n12089 = ~new_n12066 & ~new_n12088;
  assign new_n12090 = ~new_n12065_1 & ~new_n12089;
  assign new_n12091 = ~new_n11995 & ~new_n12013;
  assign new_n12092 = ~new_n11994 & ~new_n12091;
  assign new_n12093 = ~new_n11984 & ~new_n12016;
  assign new_n12094 = ~new_n11985 & ~new_n12093;
  assign new_n12095 = ~new_n11899 & new_n11908;
  assign new_n12096 = ~new_n11898 & ~new_n12095;
  assign new_n12097 = n287 & n4998;
  assign new_n12098 = n11574 & n12592;
  assign new_n12099 = new_n11882_1 & ~new_n11885;
  assign new_n12100 = ~new_n11887 & ~new_n12099;
  assign new_n12101 = ~new_n12098 & new_n12100;
  assign new_n12102 = new_n12098 & ~new_n12100;
  assign new_n12103 = ~new_n12101 & ~new_n12102;
  assign new_n12104 = ~new_n12097 & new_n12103;
  assign new_n12105 = new_n12097 & ~new_n12103;
  assign new_n12106 = ~new_n12104 & ~new_n12105;
  assign new_n12107 = new_n12096 & ~new_n12106;
  assign new_n12108 = ~new_n12096 & new_n12106;
  assign new_n12109 = ~new_n12107 & ~new_n12108;
  assign new_n12110 = new_n12094 & new_n12109;
  assign new_n12111 = ~new_n12094 & ~new_n12109;
  assign new_n12112 = ~new_n12110 & ~new_n12111;
  assign new_n12113 = ~new_n12092 & new_n12112;
  assign new_n12114 = new_n12092 & ~new_n12112;
  assign new_n12115 = ~new_n12113 & ~new_n12114;
  assign new_n12116 = n3409 & n7715;
  assign new_n12117 = n7113 & n7529;
  assign new_n12118 = new_n12116 & new_n12117;
  assign new_n12119 = ~new_n12116 & ~new_n12117;
  assign new_n12120 = ~new_n12118 & ~new_n12119;
  assign new_n12121 = n2458 & n10594;
  assign new_n12122 = n6668 & n10451;
  assign new_n12123 = n8230 & n9093;
  assign new_n12124 = ~new_n12122 & ~new_n12123;
  assign new_n12125 = new_n12122 & new_n12123;
  assign new_n12126 = ~new_n12124 & ~new_n12125;
  assign new_n12127 = n2458 & n9093;
  assign new_n12128 = n8230 & n10451;
  assign new_n12129 = new_n12127 & new_n12128;
  assign new_n12130 = ~new_n12127 & ~new_n12128;
  assign new_n12131 = n7715 & n10594;
  assign new_n12132 = ~new_n12130 & new_n12131;
  assign new_n12133 = ~new_n12129 & ~new_n12132;
  assign new_n12134 = ~new_n12126 & new_n12133;
  assign new_n12135 = new_n12126 & ~new_n12133;
  assign new_n12136 = ~new_n12134 & ~new_n12135;
  assign new_n12137 = ~new_n12121 & ~new_n12136;
  assign new_n12138 = new_n12121 & new_n12136;
  assign new_n12139 = ~new_n12137 & ~new_n12138;
  assign new_n12140 = ~new_n12120 & ~new_n12139;
  assign new_n12141 = n3409 & n7529;
  assign new_n12142 = new_n10105 & ~new_n10108;
  assign new_n12143 = ~new_n10109 & ~new_n12142;
  assign new_n12144 = ~new_n12141 & new_n12143;
  assign new_n12145 = new_n12141 & ~new_n12143;
  assign new_n12146 = ~new_n12129 & ~new_n12130;
  assign new_n12147 = ~new_n12131 & ~new_n12146;
  assign new_n12148 = new_n12131 & new_n12146;
  assign new_n12149 = ~new_n12147 & ~new_n12148;
  assign new_n12150 = ~new_n12145 & ~new_n12149;
  assign new_n12151 = ~new_n12144 & ~new_n12150;
  assign new_n12152 = ~new_n12140 & new_n12151;
  assign new_n12153 = new_n12118 & new_n12152;
  assign new_n12154 = new_n12120 & new_n12139;
  assign new_n12155 = ~new_n12118 & ~new_n12152;
  assign new_n12156 = ~new_n12154 & new_n12155;
  assign new_n12157 = n499 & n7772;
  assign new_n12158 = n7113 & n7715;
  assign new_n12159 = n1302 & n7529;
  assign new_n12160 = ~new_n12158 & ~new_n12159;
  assign new_n12161 = new_n12158 & new_n12159;
  assign new_n12162 = ~new_n12160 & ~new_n12161;
  assign new_n12163 = new_n12157 & ~new_n12162;
  assign new_n12164 = ~new_n12157 & new_n12162;
  assign new_n12165 = ~new_n12163 & ~new_n12164;
  assign new_n12166 = ~new_n12121 & ~new_n12135;
  assign new_n12167 = ~new_n12134 & ~new_n12166;
  assign new_n12168 = ~new_n12165 & new_n12167;
  assign new_n12169 = new_n12165 & ~new_n12167;
  assign new_n12170 = ~new_n12168 & ~new_n12169;
  assign new_n12171 = n2458 & n3409;
  assign new_n12172 = new_n12125 & new_n12171;
  assign new_n12173 = ~new_n12125 & ~new_n12171;
  assign new_n12174 = ~new_n12172 & ~new_n12173;
  assign new_n12175 = n8230 & n10594;
  assign new_n12176 = n6668 & n9093;
  assign new_n12177 = n7812 & n10451;
  assign new_n12178 = ~new_n12176 & ~new_n12177;
  assign new_n12179 = new_n12176 & new_n12177;
  assign new_n12180 = ~new_n12178 & ~new_n12179;
  assign new_n12181 = new_n12175 & ~new_n12180;
  assign new_n12182 = ~new_n12175 & new_n12180;
  assign new_n12183 = ~new_n12181 & ~new_n12182;
  assign new_n12184 = new_n12174 & new_n12183;
  assign new_n12185 = ~new_n12174 & ~new_n12183;
  assign new_n12186 = ~new_n12184 & ~new_n12185;
  assign new_n12187_1 = ~new_n12170 & ~new_n12186;
  assign new_n12188 = new_n12170 & new_n12186;
  assign new_n12189 = ~new_n12187_1 & ~new_n12188;
  assign new_n12190 = ~new_n12156 & ~new_n12189;
  assign new_n12191 = ~new_n12153 & ~new_n12190;
  assign new_n12192 = n11061 & n12482;
  assign new_n12193 = ~new_n12001 & ~new_n12192;
  assign new_n12194 = new_n12001 & new_n12192;
  assign new_n12195 = ~new_n12193 & ~new_n12194;
  assign new_n12196 = n9 & n1307;
  assign new_n12197 = n2339 & n2592;
  assign new_n12198 = ~new_n12196 & new_n12197;
  assign new_n12199 = new_n12196 & ~new_n12197;
  assign new_n12200 = ~new_n12198 & ~new_n12199;
  assign new_n12201 = ~new_n12195 & new_n12200;
  assign new_n12202 = new_n12195 & ~new_n12200;
  assign new_n12203 = ~new_n12201 & ~new_n12202;
  assign new_n12204 = new_n11997 & ~new_n12000;
  assign new_n12205 = ~new_n12002 & ~new_n12204;
  assign new_n12206 = n6843 & n8466;
  assign new_n12207 = n2590 & n9570;
  assign new_n12208 = ~new_n12206 & new_n12207;
  assign new_n12209 = new_n12206 & ~new_n12207;
  assign new_n12210 = ~new_n12208 & ~new_n12209;
  assign new_n12211 = new_n12205 & new_n12210;
  assign new_n12212 = ~new_n12205 & ~new_n12210;
  assign new_n12213 = ~new_n12211 & ~new_n12212;
  assign new_n12214 = new_n12203 & new_n12213;
  assign new_n12215 = ~new_n12203 & ~new_n12213;
  assign new_n12216 = ~new_n12214 & ~new_n12215;
  assign new_n12217 = new_n12006 & ~new_n12008;
  assign new_n12218 = ~new_n12009 & ~new_n12217;
  assign new_n12219 = new_n12216 & ~new_n12218;
  assign new_n12220 = ~new_n12216 & new_n12218;
  assign new_n12221 = ~new_n12219 & ~new_n12220;
  assign new_n12222 = ~new_n11895_1 & new_n11911;
  assign new_n12223 = ~new_n11894 & ~new_n12222;
  assign new_n12224 = new_n11830 & ~new_n11903;
  assign new_n12225 = ~new_n11904 & ~new_n12224;
  assign new_n12226 = ~new_n12223 & ~new_n12225;
  assign new_n12227 = new_n12223 & new_n12225;
  assign new_n12228 = ~new_n12226 & ~new_n12227;
  assign new_n12229 = ~new_n12221 & new_n12228;
  assign new_n12230 = new_n12221 & ~new_n12228;
  assign new_n12231 = ~new_n12229 & ~new_n12230;
  assign new_n12232 = new_n12191 & ~new_n12231;
  assign new_n12233 = ~new_n12191 & new_n12231;
  assign new_n12234 = ~new_n12232 & ~new_n12233;
  assign new_n12235 = n7772 & n11111;
  assign new_n12236 = n3409 & n8230;
  assign new_n12237 = new_n12235 & ~new_n12236;
  assign new_n12238 = ~new_n12235 & new_n12236;
  assign new_n12239 = ~new_n12237 & ~new_n12238;
  assign new_n12240 = n7812 & n9093;
  assign new_n12241 = n6668 & n10594;
  assign new_n12242 = ~new_n12240 & ~new_n12241;
  assign new_n12243 = new_n12240 & new_n12241;
  assign new_n12244 = ~new_n12242 & ~new_n12243;
  assign new_n12245 = ~new_n12239 & new_n12244;
  assign new_n12246 = new_n12239 & ~new_n12244;
  assign new_n12247 = ~new_n12245 & ~new_n12246;
  assign new_n12248 = ~new_n11990 & new_n12247;
  assign new_n12249 = new_n11990 & ~new_n12247;
  assign new_n12250 = ~new_n12248 & ~new_n12249;
  assign new_n12251 = ~new_n12234 & new_n12250;
  assign new_n12252 = new_n12234 & ~new_n12250;
  assign new_n12253 = ~new_n12251 & ~new_n12252;
  assign new_n12254 = new_n12115 & ~new_n12253;
  assign new_n12255 = ~new_n12115 & new_n12253;
  assign new_n12256 = ~new_n12254 & ~new_n12255;
  assign new_n12257 = ~new_n12020 & ~new_n12036;
  assign new_n12258 = ~new_n12140 & ~new_n12154;
  assign new_n12259 = ~new_n12151 & ~new_n12258;
  assign new_n12260 = new_n12151 & new_n12258;
  assign new_n12261 = ~new_n12259 & ~new_n12260;
  assign new_n12262 = n7113 & n7772;
  assign new_n12263_1 = ~new_n12144 & ~new_n12145;
  assign new_n12264 = ~new_n12149 & ~new_n12263_1;
  assign new_n12265 = new_n12149 & new_n12263_1;
  assign new_n12266 = ~new_n12264 & ~new_n12265;
  assign new_n12267 = new_n12262 & new_n12266;
  assign new_n12268 = ~new_n12262 & ~new_n12266;
  assign new_n12269 = ~new_n10102 & ~new_n10113_1;
  assign new_n12270 = ~new_n10103 & ~new_n12269;
  assign new_n12271 = ~new_n12268 & ~new_n12270;
  assign new_n12272 = ~new_n12267 & ~new_n12271;
  assign new_n12273 = new_n12261 & ~new_n12272;
  assign new_n12274 = ~new_n12153 & ~new_n12156;
  assign new_n12275 = new_n12189 & new_n12274;
  assign new_n12276 = ~new_n12189 & ~new_n12274;
  assign new_n12277 = ~new_n12275 & ~new_n12276;
  assign new_n12278 = new_n12273 & ~new_n12277;
  assign new_n12279 = n1302 & n7772;
  assign new_n12280 = ~new_n12261 & new_n12272;
  assign new_n12281 = ~new_n12273 & ~new_n12280;
  assign new_n12282 = new_n12279 & new_n12281;
  assign new_n12283 = new_n12267 & ~new_n12270;
  assign new_n12284_1 = new_n12268 & new_n12270;
  assign new_n12285 = new_n12272 & ~new_n12284_1;
  assign new_n12286 = ~new_n12283 & ~new_n12285;
  assign new_n12287 = new_n10118 & ~new_n12286;
  assign new_n12288 = ~new_n12279 & ~new_n12281;
  assign new_n12289_1 = ~new_n12282 & ~new_n12288;
  assign new_n12290 = new_n12287 & new_n12289_1;
  assign new_n12291 = ~new_n12282 & ~new_n12290;
  assign new_n12292 = ~new_n12273 & new_n12277;
  assign new_n12293 = ~new_n12278 & ~new_n12292;
  assign new_n12294 = ~new_n12291 & new_n12293;
  assign new_n12295 = ~new_n12278 & ~new_n12294;
  assign new_n12296 = new_n12257 & new_n12295;
  assign new_n12297 = ~new_n12257 & ~new_n12295;
  assign new_n12298 = ~new_n12296 & ~new_n12297;
  assign new_n12299 = new_n12256 & new_n12298;
  assign new_n12300 = ~new_n12256 & ~new_n12298;
  assign new_n12301 = ~new_n12299 & ~new_n12300;
  assign new_n12302 = ~new_n11923 & ~new_n11926;
  assign new_n12303 = new_n11760 & ~new_n11763;
  assign new_n12304 = ~new_n11764 & ~new_n12303;
  assign new_n12305 = new_n11914 & ~new_n11917;
  assign new_n12306_1 = ~new_n11918 & ~new_n12305;
  assign new_n12307 = ~new_n11772 & new_n11789;
  assign new_n12308 = ~new_n11771 & ~new_n12307;
  assign new_n12309 = n4419 & n11058;
  assign new_n12310 = n401 & n1007;
  assign new_n12311 = n3178 & n8859;
  assign new_n12312 = ~new_n12310 & new_n12311;
  assign new_n12313 = new_n12310 & ~new_n12311;
  assign new_n12314 = ~new_n12312 & ~new_n12313;
  assign new_n12315 = new_n12309 & new_n12314;
  assign new_n12316 = ~new_n12309 & ~new_n12314;
  assign new_n12317 = ~new_n12315 & ~new_n12316;
  assign new_n12318 = n951 & n5969;
  assign new_n12319 = n2498 & n11537;
  assign new_n12320 = ~new_n12318 & ~new_n12319;
  assign new_n12321 = new_n12318 & new_n12319;
  assign new_n12322 = ~new_n12320 & ~new_n12321;
  assign new_n12323 = n767 & n1198;
  assign new_n12324 = new_n11886 & ~new_n12323;
  assign new_n12325 = ~new_n11886 & new_n12323;
  assign new_n12326 = ~new_n12324 & ~new_n12325;
  assign new_n12327 = new_n12322 & new_n12326;
  assign new_n12328 = ~new_n12322 & ~new_n12326;
  assign new_n12329 = ~new_n12327 & ~new_n12328;
  assign new_n12330 = new_n12317 & ~new_n12329;
  assign new_n12331 = ~new_n12317 & new_n12329;
  assign new_n12332 = ~new_n12330 & ~new_n12331;
  assign new_n12333 = ~new_n12308 & ~new_n12332;
  assign new_n12334_1 = new_n12308 & new_n12332;
  assign new_n12335 = ~new_n12333 & ~new_n12334_1;
  assign new_n12336 = ~new_n11776 & ~new_n11786;
  assign new_n12337 = ~new_n11775 & ~new_n12336;
  assign new_n12338 = new_n11778_1 & ~new_n11781;
  assign new_n12339 = ~new_n11782 & ~new_n12338;
  assign new_n12340 = n2068 & n6818;
  assign new_n12341 = n1084 & n12348;
  assign new_n12342 = ~new_n12340 & new_n12341;
  assign new_n12343 = new_n12340 & ~new_n12341;
  assign new_n12344 = ~new_n12342 & ~new_n12343;
  assign new_n12345 = ~new_n12339 & ~new_n12344;
  assign new_n12346 = new_n12339 & new_n12344;
  assign new_n12347 = ~new_n12345 & ~new_n12346;
  assign new_n12348_1 = ~new_n12337 & ~new_n12347;
  assign new_n12349 = new_n12337 & new_n12347;
  assign new_n12350 = ~new_n12348_1 & ~new_n12349;
  assign new_n12351 = ~new_n12335 & new_n12350;
  assign new_n12352_1 = new_n12335 & ~new_n12350;
  assign new_n12353 = ~new_n12351 & ~new_n12352_1;
  assign new_n12354 = new_n12306_1 & new_n12353;
  assign new_n12355 = ~new_n12306_1 & ~new_n12353;
  assign new_n12356 = ~new_n12354 & ~new_n12355;
  assign new_n12357 = ~new_n12304 & new_n12356;
  assign new_n12358 = new_n12304 & ~new_n12356;
  assign new_n12359 = ~new_n12357 & ~new_n12358;
  assign new_n12360 = new_n12302 & new_n12359;
  assign new_n12361 = ~new_n12302 & ~new_n12359;
  assign new_n12362 = ~new_n12360 & ~new_n12361;
  assign new_n12363 = ~new_n11796 & ~new_n11812;
  assign new_n12364 = ~new_n11757 & ~new_n11792_1;
  assign new_n12365 = ~new_n11758 & ~new_n12364;
  assign new_n12366 = n4452 & n5962;
  assign new_n12367 = new_n12365 & new_n12366;
  assign new_n12368 = ~new_n12365 & ~new_n12366;
  assign new_n12369 = ~new_n12367 & ~new_n12368;
  assign new_n12370 = ~new_n12169 & ~new_n12186;
  assign new_n12371 = ~new_n12168 & ~new_n12370;
  assign new_n12372_1 = ~new_n12173 & ~new_n12183;
  assign new_n12373 = ~new_n12172 & ~new_n12372_1;
  assign new_n12374 = n1392 & n9216;
  assign new_n12375 = n6085 & n10657;
  assign new_n12376 = n9906 & n10142;
  assign new_n12377 = ~new_n12375 & ~new_n12376;
  assign new_n12378 = new_n12375 & new_n12376;
  assign new_n12379 = ~new_n12377 & ~new_n12378;
  assign new_n12380 = n8183 & n11109;
  assign new_n12381 = n8468 & n11324;
  assign new_n12382 = new_n12380 & ~new_n12381;
  assign new_n12383 = ~new_n12380 & new_n12381;
  assign new_n12384 = ~new_n12382 & ~new_n12383;
  assign new_n12385 = ~new_n12379 & ~new_n12384;
  assign new_n12386 = new_n12379 & new_n12384;
  assign new_n12387 = ~new_n12385 & ~new_n12386;
  assign new_n12388 = ~new_n12374 & new_n12387;
  assign new_n12389 = new_n12374 & ~new_n12387;
  assign new_n12390 = ~new_n12388 & ~new_n12389;
  assign new_n12391 = new_n12373 & new_n12390;
  assign new_n12392 = ~new_n12373 & ~new_n12390;
  assign new_n12393 = ~new_n12391 & ~new_n12392;
  assign new_n12394 = new_n12371 & ~new_n12393;
  assign new_n12395 = ~new_n12371 & new_n12393;
  assign new_n12396 = ~new_n12394 & ~new_n12395;
  assign new_n12397 = ~new_n12369 & ~new_n12396;
  assign new_n12398 = new_n12369 & new_n12396;
  assign new_n12399 = ~new_n12397 & ~new_n12398;
  assign new_n12400 = new_n12157 & ~new_n12160;
  assign new_n12401 = ~new_n12161 & ~new_n12400;
  assign new_n12402 = new_n12175 & ~new_n12178;
  assign new_n12403 = ~new_n12179 & ~new_n12402;
  assign new_n12404 = ~new_n12401 & new_n12403;
  assign new_n12405 = new_n12401 & ~new_n12403;
  assign new_n12406_1 = ~new_n12404 & ~new_n12405;
  assign new_n12407 = n1302 & n7715;
  assign new_n12408_1 = n499 & n7529;
  assign new_n12409 = n2458 & n7113;
  assign new_n12410 = new_n12408_1 & ~new_n12409;
  assign new_n12411 = ~new_n12408_1 & new_n12409;
  assign new_n12412 = ~new_n12410 & ~new_n12411;
  assign new_n12413 = new_n12407 & new_n12412;
  assign new_n12414 = ~new_n12407 & ~new_n12412;
  assign new_n12415 = ~new_n12413 & ~new_n12414;
  assign new_n12416 = new_n12406_1 & new_n12415;
  assign new_n12417 = ~new_n12406_1 & ~new_n12415;
  assign new_n12418 = ~new_n12416 & ~new_n12417;
  assign new_n12419 = ~new_n12399 & new_n12418;
  assign new_n12420 = new_n12399 & ~new_n12418;
  assign new_n12421 = ~new_n12419 & ~new_n12420;
  assign new_n12422 = new_n12363 & ~new_n12421;
  assign new_n12423 = ~new_n12363 & new_n12421;
  assign new_n12424 = ~new_n12422 & ~new_n12423;
  assign new_n12425 = ~new_n12362 & new_n12424;
  assign new_n12426 = new_n12362 & ~new_n12424;
  assign new_n12427 = ~new_n12425 & ~new_n12426;
  assign new_n12428 = ~new_n12061 & new_n12427;
  assign new_n12429 = new_n12061 & ~new_n12427;
  assign new_n12430 = ~new_n12428 & ~new_n12429;
  assign new_n12431 = ~new_n12301 & new_n12430;
  assign new_n12432 = new_n12301 & ~new_n12430;
  assign new_n12433 = ~new_n12431 & ~new_n12432;
  assign new_n12434 = new_n12090 & ~new_n12433;
  assign new_n12435 = ~new_n12090 & new_n12433;
  assign new_n12436 = ~new_n12434 & ~new_n12435;
  assign new_n12437 = new_n12291 & ~new_n12293;
  assign new_n12438 = ~new_n12294 & ~new_n12437;
  assign new_n12439 = new_n12066 & new_n12088;
  assign new_n12440 = new_n12065_1 & ~new_n12088;
  assign new_n12441 = ~new_n12090 & ~new_n12440;
  assign new_n12442 = ~new_n12439 & ~new_n12441;
  assign new_n12443 = ~new_n12438 & ~new_n12442;
  assign new_n12444 = new_n12438 & new_n12442;
  assign new_n12445 = ~new_n12287 & ~new_n12289_1;
  assign new_n12446 = ~new_n12290 & ~new_n12445;
  assign new_n12447 = ~new_n12073 & ~new_n12074;
  assign new_n12448 = new_n12086 & ~new_n12447;
  assign new_n12449 = ~new_n12086 & new_n12447;
  assign new_n12450 = ~new_n12448 & ~new_n12449;
  assign new_n12451 = ~new_n12446 & ~new_n12450;
  assign new_n12452 = new_n12446 & new_n12450;
  assign new_n12453 = ~new_n10118 & new_n12286;
  assign new_n12454 = ~new_n12287 & ~new_n12453;
  assign new_n12455 = ~new_n12081 & ~new_n12082;
  assign new_n12456 = new_n12084 & ~new_n12455;
  assign new_n12457 = ~new_n12084 & new_n12455;
  assign new_n12458 = ~new_n12456 & ~new_n12457;
  assign new_n12459 = ~new_n12454 & ~new_n12458;
  assign new_n12460 = new_n12454 & new_n12458;
  assign new_n12461 = ~new_n10248 & ~new_n10261;
  assign new_n12462 = ~new_n10247 & ~new_n12461;
  assign new_n12463_1 = ~new_n12460 & new_n12462;
  assign new_n12464 = ~new_n12459 & ~new_n12463_1;
  assign new_n12465 = ~new_n12452 & ~new_n12464;
  assign new_n12466 = ~new_n12451 & ~new_n12465;
  assign new_n12467 = ~new_n12444 & ~new_n12466;
  assign new_n12468 = ~new_n12443 & ~new_n12467;
  assign new_n12469 = new_n12436 & ~new_n12468;
  assign new_n12470 = ~new_n12436 & new_n12468;
  assign n7034 = ~new_n12469 & ~new_n12470;
  assign new_n12472 = ~new_n12459 & ~new_n12460;
  assign new_n12473 = new_n12462 & new_n12472;
  assign new_n12474 = ~new_n12462 & ~new_n12472;
  assign n7111 = new_n12473 | new_n12474;
  assign new_n12476 = n7529 & n7772;
  assign new_n12477 = n7772 & n11734;
  assign new_n12478 = ~n7529 & ~new_n12477;
  assign new_n12479 = ~n7715 & new_n12478;
  assign new_n12480 = n11734 & new_n12476;
  assign new_n12481 = ~n7715 & ~new_n12480;
  assign new_n12482_1 = ~new_n12478 & ~new_n12481;
  assign new_n12483 = n7715 & new_n12480;
  assign new_n12484 = new_n12482_1 & ~new_n12483;
  assign new_n12485 = ~new_n12479 & ~new_n12484;
  assign new_n12486 = new_n12476 & new_n12485;
  assign new_n12487 = n7529 & n11734;
  assign new_n12488 = n7715 & new_n12487;
  assign new_n12489 = ~n7715 & ~new_n12487;
  assign new_n12490 = n2458 & ~new_n12489;
  assign new_n12491 = ~new_n12488 & ~new_n12490;
  assign new_n12492 = ~n2458 & new_n12489;
  assign new_n12493 = new_n12491 & ~new_n12492;
  assign new_n12494 = n2458 & new_n12488;
  assign new_n12495 = ~new_n12493 & ~new_n12494;
  assign new_n12496 = n7772 & n12651;
  assign new_n12497 = ~new_n12482_1 & ~new_n12496;
  assign new_n12498 = new_n12482_1 & new_n12496;
  assign new_n12499 = ~new_n12497 & ~new_n12498;
  assign new_n12500 = new_n12495 & ~new_n12499;
  assign new_n12501 = ~new_n12495 & new_n12499;
  assign new_n12502 = ~new_n12500 & ~new_n12501;
  assign new_n12503_1 = new_n12486 & new_n12502;
  assign new_n12504 = n7411 & n7772;
  assign new_n12505 = n7715 & n11734;
  assign new_n12506 = n2458 & new_n12505;
  assign new_n12507 = ~n2458 & ~new_n12505;
  assign new_n12508 = n8230 & ~new_n12507;
  assign new_n12509 = ~new_n12506 & ~new_n12508;
  assign new_n12510 = ~n8230 & new_n12507;
  assign new_n12511 = new_n12509 & ~new_n12510;
  assign new_n12512 = n8230 & new_n12506;
  assign new_n12513 = ~new_n12511 & ~new_n12512;
  assign new_n12514 = n7529 & n12651;
  assign new_n12515_1 = new_n12491 & ~new_n12514;
  assign new_n12516 = ~new_n12491 & new_n12514;
  assign new_n12517 = ~new_n12515_1 & ~new_n12516;
  assign new_n12518 = new_n12513 & ~new_n12517;
  assign new_n12519 = ~new_n12513 & new_n12517;
  assign new_n12520 = ~new_n12518 & ~new_n12519;
  assign new_n12521 = ~new_n12504 & ~new_n12520;
  assign new_n12522 = new_n12504 & new_n12520;
  assign new_n12523 = ~new_n12521 & ~new_n12522;
  assign new_n12524 = ~new_n12495 & ~new_n12497;
  assign new_n12525 = ~new_n12498 & ~new_n12524;
  assign new_n12526 = ~new_n12523 & ~new_n12525;
  assign new_n12527 = new_n12523 & new_n12525;
  assign new_n12528 = ~new_n12526 & ~new_n12527;
  assign new_n12529 = new_n12503_1 & ~new_n12528;
  assign new_n12530 = ~new_n12503_1 & new_n12528;
  assign new_n12531 = ~new_n12529 & ~new_n12530;
  assign new_n12532 = ~new_n12486 & ~new_n12502;
  assign new_n12533 = ~new_n12503_1 & ~new_n12532;
  assign new_n12534 = n411 & n12348;
  assign new_n12535 = n9216 & n9475;
  assign new_n12536 = new_n12534 & new_n12535;
  assign new_n12537 = n6826 & n9216;
  assign new_n12538 = n9475 & n12348;
  assign new_n12539 = n411 & n2068;
  assign new_n12540 = ~new_n12538 & ~new_n12539;
  assign new_n12541 = new_n12538 & new_n12539;
  assign new_n12542 = ~new_n12540 & ~new_n12541;
  assign new_n12543 = new_n12537 & ~new_n12542;
  assign new_n12544 = ~new_n12537 & new_n12542;
  assign new_n12545 = ~new_n12543 & ~new_n12544;
  assign new_n12546 = new_n12536 & ~new_n12545;
  assign new_n12547 = ~new_n12536 & new_n12545;
  assign new_n12548 = ~new_n12546 & ~new_n12547;
  assign new_n12549 = n5031 & n8506;
  assign new_n12550 = n5536 & n8466;
  assign new_n12551 = new_n12549 & new_n12550;
  assign new_n12552 = n772 & n8466;
  assign new_n12553 = n5031 & n5536;
  assign new_n12554 = n9 & n8506;
  assign new_n12555 = ~new_n12553 & ~new_n12554;
  assign new_n12556 = new_n12553 & new_n12554;
  assign new_n12557 = ~new_n12555 & ~new_n12556;
  assign new_n12558 = new_n12552 & ~new_n12557;
  assign new_n12559 = ~new_n12552 & new_n12557;
  assign new_n12560 = ~new_n12558 & ~new_n12559;
  assign new_n12561 = new_n12551 & ~new_n12560;
  assign new_n12562 = ~new_n12551 & new_n12560;
  assign new_n12563 = ~new_n12561 & ~new_n12562;
  assign new_n12564 = n3085 & n12592;
  assign new_n12565 = n124 & n3178;
  assign new_n12566 = new_n12564 & new_n12565;
  assign new_n12567 = n3178 & n10805;
  assign new_n12568 = n124 & n12592;
  assign new_n12569 = n3085 & n10168;
  assign new_n12570 = ~new_n12568 & ~new_n12569;
  assign new_n12571 = new_n12568 & new_n12569;
  assign new_n12572 = ~new_n12570 & ~new_n12571;
  assign new_n12573 = new_n12567 & ~new_n12572;
  assign new_n12574 = ~new_n12567 & new_n12572;
  assign new_n12575 = ~new_n12573 & ~new_n12574;
  assign new_n12576 = new_n12566 & ~new_n12575;
  assign new_n12577 = ~new_n12566 & new_n12575;
  assign new_n12578 = ~new_n12576 & ~new_n12577;
  assign new_n12579_1 = ~new_n12563 & ~new_n12578;
  assign new_n12580 = new_n12563 & new_n12578;
  assign new_n12581 = ~new_n12579_1 & ~new_n12580;
  assign new_n12582 = ~new_n12549 & ~new_n12550;
  assign new_n12583 = ~new_n12551 & ~new_n12582;
  assign new_n12584 = new_n5652 & new_n12583;
  assign new_n12585 = ~new_n5652 & ~new_n12583;
  assign new_n12586 = ~new_n12564 & ~new_n12565;
  assign new_n12587 = ~new_n12566 & ~new_n12586;
  assign new_n12588 = ~new_n12585 & new_n12587;
  assign new_n12589 = ~new_n12584 & ~new_n12588;
  assign new_n12590 = ~new_n12581 & ~new_n12589;
  assign new_n12591 = new_n12581 & new_n12589;
  assign new_n12592_1 = ~new_n12590 & ~new_n12591;
  assign new_n12593 = ~new_n12548 & new_n12592_1;
  assign new_n12594 = new_n12548 & ~new_n12592_1;
  assign new_n12595 = ~new_n12534 & ~new_n12535;
  assign new_n12596 = ~new_n12536 & ~new_n12595;
  assign new_n12597 = ~new_n12584 & ~new_n12585;
  assign new_n12598 = new_n12587 & ~new_n12597;
  assign new_n12599 = ~new_n12587 & new_n12597;
  assign new_n12600 = ~new_n12598 & ~new_n12599;
  assign new_n12601 = ~new_n12596 & new_n12600;
  assign new_n12602 = new_n12596 & ~new_n12600;
  assign new_n12603 = ~new_n5656 & ~new_n12602;
  assign new_n12604 = ~new_n12601 & ~new_n12603;
  assign new_n12605_1 = ~new_n12594 & ~new_n12604;
  assign new_n12606 = ~new_n12593 & ~new_n12605_1;
  assign new_n12607 = n9216 & n12284;
  assign new_n12608 = new_n12537 & ~new_n12540;
  assign new_n12609 = ~new_n12541 & ~new_n12608;
  assign new_n12610 = ~new_n12607 & new_n12609;
  assign new_n12611 = new_n12607 & ~new_n12609;
  assign new_n12612 = ~new_n12610 & ~new_n12611;
  assign new_n12613 = n6826 & n12348;
  assign new_n12614 = n2068 & n9475;
  assign new_n12615 = n411 & n11324;
  assign new_n12616_1 = ~new_n12614 & ~new_n12615;
  assign new_n12617 = new_n12614 & new_n12615;
  assign new_n12618 = ~new_n12616_1 & ~new_n12617;
  assign new_n12619 = new_n12613 & ~new_n12618;
  assign new_n12620 = ~new_n12613 & new_n12618;
  assign new_n12621 = ~new_n12619 & ~new_n12620;
  assign new_n12622 = ~new_n12612 & new_n12621;
  assign new_n12623 = new_n12612 & ~new_n12621;
  assign new_n12624 = ~new_n12622 & ~new_n12623;
  assign new_n12625 = ~new_n12546 & ~new_n12624;
  assign new_n12626 = new_n12546 & new_n12624;
  assign new_n12627 = ~new_n12625 & ~new_n12626;
  assign new_n12628 = n2737 & n8466;
  assign new_n12629 = new_n12552 & ~new_n12555;
  assign new_n12630 = ~new_n12556 & ~new_n12629;
  assign new_n12631 = ~new_n12628 & new_n12630;
  assign new_n12632 = new_n12628 & ~new_n12630;
  assign new_n12633 = ~new_n12631 & ~new_n12632;
  assign new_n12634 = n772 & n5031;
  assign new_n12635 = n9 & n5536;
  assign new_n12636 = n2592 & n8506;
  assign new_n12637 = ~new_n12635 & ~new_n12636;
  assign new_n12638 = new_n12635 & new_n12636;
  assign new_n12639 = ~new_n12637 & ~new_n12638;
  assign new_n12640 = new_n12634 & ~new_n12639;
  assign new_n12641 = ~new_n12634 & new_n12639;
  assign new_n12642 = ~new_n12640 & ~new_n12641;
  assign new_n12643 = ~new_n12633 & new_n12642;
  assign new_n12644 = new_n12633 & ~new_n12642;
  assign new_n12645 = ~new_n12643 & ~new_n12644;
  assign new_n12646 = ~new_n12561 & ~new_n12645;
  assign new_n12647 = new_n12561 & new_n12645;
  assign new_n12648 = ~new_n12646 & ~new_n12647;
  assign new_n12649 = n3178 & n12263;
  assign new_n12650 = new_n12567 & ~new_n12570;
  assign new_n12651_1 = ~new_n12571 & ~new_n12650;
  assign new_n12652 = ~new_n12649 & new_n12651_1;
  assign new_n12653 = new_n12649 & ~new_n12651_1;
  assign new_n12654 = ~new_n12652 & ~new_n12653;
  assign new_n12655 = n10805 & n12592;
  assign new_n12656 = n124 & n10168;
  assign new_n12657 = n767 & n3085;
  assign new_n12658 = ~new_n12656 & ~new_n12657;
  assign new_n12659 = new_n12656 & new_n12657;
  assign new_n12660 = ~new_n12658 & ~new_n12659;
  assign new_n12661 = new_n12655 & ~new_n12660;
  assign new_n12662 = ~new_n12655 & new_n12660;
  assign new_n12663 = ~new_n12661 & ~new_n12662;
  assign new_n12664 = ~new_n12654 & new_n12663;
  assign new_n12665 = new_n12654 & ~new_n12663;
  assign new_n12666 = ~new_n12664 & ~new_n12665;
  assign new_n12667 = new_n12576 & new_n12666;
  assign new_n12668 = ~new_n12576 & ~new_n12666;
  assign new_n12669 = ~new_n12667 & ~new_n12668;
  assign new_n12670 = new_n12648 & new_n12669;
  assign new_n12671 = ~new_n12648 & ~new_n12669;
  assign new_n12672 = ~new_n12670 & ~new_n12671;
  assign new_n12673 = ~new_n12579_1 & ~new_n12589;
  assign new_n12674 = ~new_n12580 & ~new_n12673;
  assign new_n12675 = new_n12672 & new_n12674;
  assign new_n12676 = ~new_n12672 & ~new_n12674;
  assign new_n12677 = ~new_n12675 & ~new_n12676;
  assign new_n12678 = new_n12627 & ~new_n12677;
  assign new_n12679 = ~new_n12627 & new_n12677;
  assign new_n12680 = ~new_n12678 & ~new_n12679;
  assign new_n12681 = ~new_n12606 & ~new_n12680;
  assign new_n12682 = new_n12606 & new_n12680;
  assign new_n12683 = ~new_n12681 & ~new_n12682;
  assign new_n12684 = new_n12533 & new_n12683;
  assign new_n12685 = ~new_n12533 & ~new_n12683;
  assign new_n12686 = ~new_n12476 & ~new_n12485;
  assign new_n12687 = ~new_n12486 & ~new_n12686;
  assign new_n12688 = ~new_n12593 & ~new_n12594;
  assign new_n12689 = new_n12604 & ~new_n12688;
  assign new_n12690 = ~new_n12604 & new_n12688;
  assign new_n12691 = ~new_n12689 & ~new_n12690;
  assign new_n12692 = new_n12687 & ~new_n12691;
  assign new_n12693_1 = ~new_n12687 & new_n12691;
  assign new_n12694 = ~n7529 & new_n5659;
  assign new_n12695 = ~new_n12601 & ~new_n12602;
  assign new_n12696 = ~new_n5656 & new_n12695;
  assign new_n12697 = new_n5656 & ~new_n12695;
  assign new_n12698 = ~new_n12696 & ~new_n12697;
  assign new_n12699 = ~new_n12694 & new_n12698;
  assign new_n12700 = ~n7529 & ~n7772;
  assign new_n12701 = ~new_n5658 & new_n12476;
  assign new_n12702 = ~new_n12700 & ~new_n12701;
  assign new_n12703 = ~new_n12699 & new_n12702;
  assign new_n12704 = ~new_n12693_1 & new_n12703;
  assign new_n12705 = ~new_n12692 & ~new_n12704;
  assign new_n12706 = ~new_n12685 & ~new_n12705;
  assign new_n12707 = ~new_n12684 & ~new_n12706;
  assign new_n12708 = ~new_n12531 & new_n12707;
  assign new_n12709 = new_n12531 & ~new_n12707;
  assign new_n12710 = ~new_n12708 & ~new_n12709;
  assign new_n12711 = n469 & n9216;
  assign new_n12712 = n12284 & n12348;
  assign new_n12713 = new_n12613 & ~new_n12616_1;
  assign new_n12714 = ~new_n12617 & ~new_n12713;
  assign new_n12715 = ~new_n12712 & new_n12714;
  assign new_n12716 = new_n12712 & ~new_n12714;
  assign new_n12717 = ~new_n12715 & ~new_n12716;
  assign new_n12718 = n2068 & n6826;
  assign new_n12719 = n9475 & n11324;
  assign new_n12720 = n411 & n8183;
  assign new_n12721 = ~new_n12719 & ~new_n12720;
  assign new_n12722 = new_n12719 & new_n12720;
  assign new_n12723 = ~new_n12721 & ~new_n12722;
  assign new_n12724 = new_n12718 & ~new_n12723;
  assign new_n12725 = ~new_n12718 & new_n12723;
  assign new_n12726 = ~new_n12724 & ~new_n12725;
  assign new_n12727 = ~new_n12717 & new_n12726;
  assign new_n12728 = new_n12717 & ~new_n12726;
  assign new_n12729 = ~new_n12727 & ~new_n12728;
  assign new_n12730 = ~new_n12711 & ~new_n12729;
  assign new_n12731 = new_n12711 & new_n12729;
  assign new_n12732 = ~new_n12730 & ~new_n12731;
  assign new_n12733 = ~new_n12610 & ~new_n12621;
  assign new_n12734 = ~new_n12611 & ~new_n12733;
  assign new_n12735 = ~new_n12732 & new_n12734;
  assign new_n12736 = new_n12732 & ~new_n12734;
  assign new_n12737 = ~new_n12735 & ~new_n12736;
  assign new_n12738 = ~new_n12626 & ~new_n12737;
  assign new_n12739 = new_n12626 & new_n12737;
  assign new_n12740 = ~new_n12738 & ~new_n12739;
  assign new_n12741 = n8466 & n12408;
  assign new_n12742 = n2737 & n5031;
  assign new_n12743 = new_n12634 & ~new_n12637;
  assign new_n12744 = ~new_n12638 & ~new_n12743;
  assign new_n12745 = ~new_n12742 & new_n12744;
  assign new_n12746 = new_n12742 & ~new_n12744;
  assign new_n12747 = ~new_n12745 & ~new_n12746;
  assign new_n12748 = n9 & n772;
  assign new_n12749 = n2592 & n5536;
  assign new_n12750_1 = n2590 & n8506;
  assign new_n12751 = ~new_n12749 & ~new_n12750_1;
  assign new_n12752 = new_n12749 & new_n12750_1;
  assign new_n12753 = ~new_n12751 & ~new_n12752;
  assign new_n12754 = new_n12748 & ~new_n12753;
  assign new_n12755 = ~new_n12748 & new_n12753;
  assign new_n12756 = ~new_n12754 & ~new_n12755;
  assign new_n12757 = ~new_n12747 & new_n12756;
  assign new_n12758 = new_n12747 & ~new_n12756;
  assign new_n12759 = ~new_n12757 & ~new_n12758;
  assign new_n12760 = ~new_n12741 & ~new_n12759;
  assign new_n12761 = new_n12741 & new_n12759;
  assign new_n12762 = ~new_n12760 & ~new_n12761;
  assign new_n12763 = ~new_n12631 & ~new_n12642;
  assign new_n12764 = ~new_n12632 & ~new_n12763;
  assign new_n12765 = ~new_n12762 & new_n12764;
  assign new_n12766 = new_n12762 & ~new_n12764;
  assign new_n12767 = ~new_n12765 & ~new_n12766;
  assign new_n12768 = ~new_n12647 & ~new_n12767;
  assign new_n12769 = new_n12647 & new_n12767;
  assign new_n12770 = ~new_n12768 & ~new_n12769;
  assign new_n12771 = n353 & n3178;
  assign new_n12772 = n12263 & n12592;
  assign new_n12773 = new_n12655 & ~new_n12658;
  assign new_n12774 = ~new_n12659 & ~new_n12773;
  assign new_n12775 = ~new_n12772 & new_n12774;
  assign new_n12776 = new_n12772 & ~new_n12774;
  assign new_n12777 = ~new_n12775 & ~new_n12776;
  assign new_n12778 = n10168 & n10805;
  assign new_n12779 = n124 & n767;
  assign new_n12780 = n3085 & n11537;
  assign new_n12781 = ~new_n12779 & ~new_n12780;
  assign new_n12782 = new_n12779 & new_n12780;
  assign new_n12783 = ~new_n12781 & ~new_n12782;
  assign new_n12784 = new_n12778 & ~new_n12783;
  assign new_n12785 = ~new_n12778 & new_n12783;
  assign new_n12786 = ~new_n12784 & ~new_n12785;
  assign new_n12787 = ~new_n12777 & new_n12786;
  assign new_n12788 = new_n12777 & ~new_n12786;
  assign new_n12789 = ~new_n12787 & ~new_n12788;
  assign new_n12790 = ~new_n12771 & ~new_n12789;
  assign new_n12791 = new_n12771 & new_n12789;
  assign new_n12792 = ~new_n12790 & ~new_n12791;
  assign new_n12793 = ~new_n12652 & ~new_n12663;
  assign new_n12794 = ~new_n12653 & ~new_n12793;
  assign new_n12795 = ~new_n12792 & new_n12794;
  assign new_n12796 = new_n12792 & ~new_n12794;
  assign new_n12797 = ~new_n12795 & ~new_n12796;
  assign new_n12798 = ~new_n12667 & ~new_n12797;
  assign new_n12799 = new_n12667 & new_n12797;
  assign new_n12800 = ~new_n12798 & ~new_n12799;
  assign new_n12801 = new_n12770 & new_n12800;
  assign new_n12802 = ~new_n12770 & ~new_n12800;
  assign new_n12803 = ~new_n12801 & ~new_n12802;
  assign new_n12804 = ~new_n12671 & ~new_n12674;
  assign new_n12805 = ~new_n12670 & ~new_n12804;
  assign new_n12806 = new_n12803 & new_n12805;
  assign new_n12807 = ~new_n12803 & ~new_n12805;
  assign new_n12808 = ~new_n12806 & ~new_n12807;
  assign new_n12809 = ~new_n12740 & new_n12808;
  assign new_n12810 = new_n12740 & ~new_n12808;
  assign new_n12811 = ~new_n12809 & ~new_n12810;
  assign new_n12812 = ~new_n12606 & ~new_n12678;
  assign new_n12813 = ~new_n12679 & ~new_n12812;
  assign new_n12814 = new_n12811 & new_n12813;
  assign new_n12815 = ~new_n12811 & ~new_n12813;
  assign new_n12816 = ~new_n12814 & ~new_n12815;
  assign new_n12817 = ~new_n12710 & new_n12816;
  assign new_n12818 = ~new_n12709 & ~new_n12816;
  assign new_n12819 = ~new_n12708 & new_n12818;
  assign n7132 = new_n12817 | new_n12819;
  assign new_n12821 = ~new_n1350 & ~new_n1351;
  assign new_n12822 = new_n1395 & new_n12821;
  assign new_n12823 = ~new_n1395 & ~new_n12821;
  assign n7241 = ~new_n12822 & ~new_n12823;
  assign new_n12825 = ~new_n1382 & ~new_n1383;
  assign new_n12826 = ~new_n1387 & new_n12825;
  assign new_n12827 = new_n1387 & ~new_n12825;
  assign n7553 = new_n12826 | new_n12827;
  assign new_n12829 = ~new_n6040 & ~new_n6042;
  assign n7582 = new_n6043 | new_n12829;
  assign new_n12831 = ~new_n12684 & ~new_n12685;
  assign new_n12832 = new_n12705 & ~new_n12831;
  assign new_n12833 = ~new_n12705 & new_n12831;
  assign n7687 = ~new_n12832 & ~new_n12833;
  assign new_n12835 = ~new_n6030 & ~new_n6031;
  assign new_n12836 = new_n6055 & ~new_n12835;
  assign new_n12837 = ~new_n6055 & new_n12835;
  assign n7755 = new_n12836 | new_n12837;
  assign new_n12839_1 = ~new_n11691 & ~new_n11692;
  assign new_n12840 = new_n11694 & ~new_n12839_1;
  assign new_n12841 = ~new_n11694 & new_n12839_1;
  assign n7790 = ~new_n12840 & ~new_n12841;
  assign new_n12843 = ~new_n9323 & ~new_n9324;
  assign new_n12844 = new_n9347 & ~new_n12843;
  assign new_n12845 = ~new_n9347 & new_n12843;
  assign n7858 = ~new_n12844 & ~new_n12845;
  assign new_n12847 = ~new_n4861 & ~new_n4862_1;
  assign new_n12848 = new_n4916 & ~new_n12847;
  assign new_n12849 = ~new_n4916 & new_n12847;
  assign n7860 = ~new_n12848 & ~new_n12849;
  assign new_n12851 = ~new_n4011 & ~new_n4020;
  assign n7968 = ~new_n4021 & ~new_n12851;
  assign new_n12853_1 = ~new_n6022 & ~new_n6023_1;
  assign new_n12854 = new_n6057 & ~new_n12853_1;
  assign new_n12855 = ~new_n6057 & new_n12853_1;
  assign n8172 = new_n12854 | new_n12855;
  assign new_n12857 = ~new_n2609 & ~new_n2610;
  assign new_n12858 = new_n2654 & ~new_n12857;
  assign new_n12859 = ~new_n2654 & new_n12857;
  assign n8219 = new_n12858 | new_n12859;
  assign new_n12861 = ~new_n1981 & ~new_n1982_1;
  assign new_n12862 = new_n1996 & new_n12861;
  assign new_n12863 = ~new_n1996 & ~new_n12861;
  assign n8265 = ~new_n12862 & ~new_n12863;
  assign new_n12865 = ~new_n8663 & ~new_n8664;
  assign new_n12866 = new_n8666 & ~new_n12865;
  assign new_n12867 = ~new_n8666 & new_n12865;
  assign n8336 = ~new_n12866 & ~new_n12867;
  assign new_n12869 = ~new_n3505 & ~new_n3506;
  assign new_n12870 = ~new_n3516 & ~new_n12869;
  assign new_n12871 = new_n3516 & new_n12869;
  assign n8516 = ~new_n12870 & ~new_n12871;
  assign new_n12873 = ~new_n10961 & ~new_n10962;
  assign new_n12874 = ~new_n10966 & ~new_n12873;
  assign new_n12875 = new_n10966 & new_n12873;
  assign n8701 = ~new_n12874 & ~new_n12875;
  assign new_n12877 = ~n3006 & ~new_n9335;
  assign n9100 = ~new_n9343 & ~new_n12877;
  assign new_n12879 = ~new_n10955 & ~new_n10956;
  assign new_n12880 = ~new_n10968 & ~new_n12879;
  assign new_n12881 = new_n10968 & new_n12879;
  assign n9329 = new_n12880 | new_n12881;
  assign new_n12883 = ~new_n8635 & ~new_n8636;
  assign new_n12884 = ~new_n8680 & new_n12883;
  assign new_n12885 = new_n8680 & ~new_n12883;
  assign n9866 = new_n12884 | new_n12885;
  assign new_n12887 = n2252 & n10113;
  assign new_n12888 = n1757 & n4330;
  assign new_n12889 = ~new_n12887 & ~new_n12888;
  assign new_n12890 = new_n12887 & new_n12888;
  assign new_n12891 = ~new_n12889 & ~new_n12890;
  assign new_n12892 = ~new_n5429 & ~new_n5433;
  assign new_n12893 = ~new_n5432 & ~new_n12892;
  assign new_n12894 = n7659 & n10416;
  assign new_n12895 = n5729 & n11488;
  assign new_n12896 = n11030 & n12289;
  assign new_n12897 = ~new_n12895 & ~new_n12896;
  assign new_n12898 = new_n12895 & new_n12896;
  assign new_n12899 = ~new_n12897 & ~new_n12898;
  assign new_n12900 = new_n12894 & new_n12899;
  assign new_n12901 = ~new_n12894 & ~new_n12899;
  assign new_n12902 = ~new_n12900 & ~new_n12901;
  assign new_n12903 = ~new_n12893 & ~new_n12902;
  assign new_n12904 = new_n12893 & new_n12902;
  assign new_n12905 = ~new_n12903 & ~new_n12904;
  assign new_n12906 = ~new_n12891 & ~new_n12905;
  assign new_n12907 = new_n12891 & new_n12905;
  assign new_n12908 = ~new_n12906 & ~new_n12907;
  assign new_n12909 = ~new_n5427_1 & new_n5437;
  assign new_n12910 = ~new_n5426 & ~new_n12909;
  assign new_n12911 = new_n12908 & new_n12910;
  assign new_n12912_1 = ~new_n12908 & ~new_n12910;
  assign new_n12913 = ~new_n12911 & ~new_n12912_1;
  assign new_n12914 = ~new_n5441 & new_n5445;
  assign new_n12915 = ~new_n5442 & ~new_n12914;
  assign new_n12916 = new_n12913 & ~new_n12915;
  assign new_n12917 = ~new_n12906 & new_n12910;
  assign new_n12918 = ~new_n12890 & ~new_n12917;
  assign new_n12919 = ~new_n12907 & new_n12918;
  assign new_n12920 = new_n12890 & new_n12917;
  assign new_n12921 = ~new_n12919 & ~new_n12920;
  assign new_n12922 = n1757 & n2252;
  assign new_n12923 = n2482 & n5884;
  assign new_n12924 = n9747 & n10113;
  assign new_n12925 = ~new_n12923 & ~new_n12924;
  assign new_n12926 = new_n12923 & new_n12924;
  assign new_n12927 = ~new_n12925 & ~new_n12926;
  assign new_n12928 = new_n12922 & ~new_n12927;
  assign new_n12929 = ~new_n12922 & new_n12927;
  assign new_n12930 = ~new_n12928 & ~new_n12929;
  assign new_n12931 = ~new_n12893 & ~new_n12900;
  assign new_n12932 = ~new_n12901 & ~new_n12931;
  assign new_n12933 = new_n12930 & ~new_n12932;
  assign new_n12934 = n4330 & n10416;
  assign new_n12935 = new_n12898 & new_n12934;
  assign new_n12936 = ~new_n12898 & ~new_n12934;
  assign new_n12937 = ~new_n12935 & ~new_n12936;
  assign new_n12938 = n1982 & n5729;
  assign new_n12939 = n11488 & n12289;
  assign new_n12940 = n7659 & n11030;
  assign new_n12941 = ~new_n12939 & ~new_n12940;
  assign new_n12942 = new_n12939 & new_n12940;
  assign new_n12943 = ~new_n12941 & ~new_n12942;
  assign new_n12944 = new_n12938 & ~new_n12943;
  assign new_n12945 = ~new_n12938 & new_n12943;
  assign new_n12946 = ~new_n12944 & ~new_n12945;
  assign new_n12947 = new_n12937 & new_n12946;
  assign new_n12948 = ~new_n12937 & ~new_n12946;
  assign new_n12949 = ~new_n12947 & ~new_n12948;
  assign new_n12950 = new_n12933 & new_n12949;
  assign new_n12951 = ~new_n12930 & new_n12932;
  assign new_n12952 = ~new_n12949 & new_n12951;
  assign new_n12953 = ~new_n12933 & ~new_n12949;
  assign new_n12954 = ~new_n12951 & ~new_n12953;
  assign new_n12955 = ~new_n12952 & ~new_n12954;
  assign new_n12956 = ~new_n12950 & ~new_n12955;
  assign new_n12957 = new_n12921 & ~new_n12956;
  assign new_n12958 = ~new_n12921 & new_n12956;
  assign new_n12959 = ~new_n12957 & ~new_n12958;
  assign new_n12960 = ~new_n12916 & new_n12959;
  assign new_n12961 = new_n12916 & ~new_n12959;
  assign new_n12962 = ~new_n12960 & ~new_n12961;
  assign new_n12963 = n2482 & n9747;
  assign new_n12964 = ~new_n12913 & new_n12915;
  assign new_n12965_1 = ~new_n12916 & ~new_n12964;
  assign new_n12966 = new_n12963 & new_n12965_1;
  assign new_n12967 = ~new_n12963 & ~new_n12965_1;
  assign new_n12968_1 = ~new_n12966 & ~new_n12967;
  assign new_n12969 = new_n5450 & new_n12968_1;
  assign new_n12970 = ~new_n12966 & ~new_n12969;
  assign new_n12971 = ~new_n12962 & new_n12970;
  assign new_n12972 = new_n12962 & ~new_n12970;
  assign new_n12973 = ~new_n12971 & ~new_n12972;
  assign new_n12974 = ~new_n5560 & new_n5563;
  assign new_n12975 = ~new_n5559 & ~new_n12974;
  assign new_n12976 = n5065 & n11236;
  assign new_n12977 = n1636 & n4382;
  assign new_n12978 = ~new_n12976 & ~new_n12977;
  assign new_n12979 = new_n12976 & new_n12977;
  assign new_n12980 = ~new_n12978 & ~new_n12979;
  assign new_n12981 = n3130 & n4862;
  assign new_n12982 = n5920 & n9732;
  assign new_n12983 = n103 & n13058;
  assign new_n12984 = ~new_n12982 & ~new_n12983;
  assign new_n12985 = new_n12982 & new_n12983;
  assign new_n12986 = ~new_n12984 & ~new_n12985;
  assign new_n12987 = ~new_n12981 & ~new_n12986;
  assign new_n12988 = new_n12981 & new_n12986;
  assign new_n12989 = ~new_n12987 & ~new_n12988;
  assign new_n12990 = new_n5547 & ~new_n5550;
  assign new_n12991 = ~new_n5551 & ~new_n12990;
  assign new_n12992 = ~new_n12989 & new_n12991;
  assign new_n12993 = new_n12989 & ~new_n12991;
  assign new_n12994 = ~new_n12992 & ~new_n12993;
  assign new_n12995 = ~new_n12980 & ~new_n12994;
  assign new_n12996 = new_n12980 & new_n12994;
  assign new_n12997 = ~new_n12995 & ~new_n12996;
  assign new_n12998 = ~new_n5544 & ~new_n5555;
  assign new_n12999 = ~new_n5545 & ~new_n12998;
  assign new_n13000 = ~new_n12997 & ~new_n12999;
  assign new_n13001 = new_n12997 & new_n12999;
  assign new_n13002_1 = ~new_n13000 & ~new_n13001;
  assign new_n13003 = new_n12975 & ~new_n13002_1;
  assign new_n13004 = ~new_n12995 & ~new_n12999;
  assign new_n13005 = ~new_n12979 & ~new_n13004;
  assign new_n13006 = ~new_n12996 & new_n13005;
  assign new_n13007 = new_n12979 & new_n13004;
  assign new_n13008 = ~new_n13006 & ~new_n13007;
  assign new_n13009 = n4382 & n5065;
  assign new_n13010 = n8228 & n11835;
  assign new_n13011 = n443 & n11236;
  assign new_n13012 = ~new_n13010 & ~new_n13011;
  assign new_n13013 = new_n13010 & new_n13011;
  assign new_n13014 = ~new_n13012 & ~new_n13013;
  assign new_n13015 = new_n13009 & ~new_n13014;
  assign new_n13016 = ~new_n13009 & new_n13014;
  assign new_n13017 = ~new_n13015 & ~new_n13016;
  assign new_n13018 = ~new_n12988 & new_n12991;
  assign new_n13019 = ~new_n12987 & ~new_n13018;
  assign new_n13020 = new_n13017 & ~new_n13019;
  assign new_n13021 = n1636 & n3130;
  assign new_n13022 = new_n12985 & new_n13021;
  assign new_n13023 = ~new_n12985 & ~new_n13021;
  assign new_n13024 = ~new_n13022 & ~new_n13023;
  assign new_n13025 = n5320 & n13058;
  assign new_n13026 = n103 & n5920;
  assign new_n13027 = n4862 & n9732;
  assign new_n13028 = ~new_n13026 & ~new_n13027;
  assign new_n13029 = new_n13026 & new_n13027;
  assign new_n13030 = ~new_n13028 & ~new_n13029;
  assign new_n13031 = new_n13025 & ~new_n13030;
  assign new_n13032 = ~new_n13025 & new_n13030;
  assign new_n13033 = ~new_n13031 & ~new_n13032;
  assign new_n13034 = new_n13024 & new_n13033;
  assign new_n13035_1 = ~new_n13024 & ~new_n13033;
  assign new_n13036 = ~new_n13034 & ~new_n13035_1;
  assign new_n13037 = new_n13020 & new_n13036;
  assign new_n13038 = ~new_n13017 & new_n13019;
  assign new_n13039 = new_n13036 & ~new_n13038;
  assign new_n13040 = ~new_n13020 & ~new_n13039;
  assign new_n13041 = ~new_n13037 & ~new_n13040;
  assign new_n13042 = ~new_n13036 & new_n13038;
  assign new_n13043 = ~new_n13041 & ~new_n13042;
  assign new_n13044 = ~new_n13008 & new_n13043;
  assign new_n13045 = new_n13008 & ~new_n13043;
  assign new_n13046 = ~new_n13044 & ~new_n13045;
  assign new_n13047 = ~new_n13003 & ~new_n13046;
  assign new_n13048 = new_n13003 & new_n13046;
  assign new_n13049 = ~new_n13047 & ~new_n13048;
  assign new_n13050 = n443 & n8228;
  assign new_n13051 = ~new_n12975 & new_n13002_1;
  assign new_n13052 = ~new_n13003 & ~new_n13051;
  assign new_n13053 = new_n13050 & new_n13052;
  assign new_n13054 = ~new_n13050 & ~new_n13052;
  assign new_n13055 = ~new_n13053 & ~new_n13054;
  assign new_n13056 = new_n5568_1 & new_n13055;
  assign new_n13057 = ~new_n13053 & ~new_n13056;
  assign new_n13058_1 = ~new_n13049 & new_n13057;
  assign new_n13059 = new_n13049 & ~new_n13057;
  assign new_n13060_1 = ~new_n13058_1 & ~new_n13059;
  assign new_n13061 = ~new_n5589 & ~new_n5595;
  assign new_n13062 = n5684 & n8860;
  assign new_n13063 = n1916 & n4964;
  assign new_n13064 = ~new_n13062 & ~new_n13063;
  assign new_n13065 = new_n13062 & new_n13063;
  assign new_n13066 = ~new_n13064 & ~new_n13065;
  assign new_n13067 = n10162 & n10522;
  assign new_n13068 = n6392 & n10770;
  assign new_n13069 = n3769 & new_n13068;
  assign new_n13070 = ~new_n5577 & ~new_n13068;
  assign new_n13071 = ~new_n13069 & ~new_n13070;
  assign new_n13072 = ~new_n13067 & ~new_n13071;
  assign new_n13073 = new_n13067 & new_n13071;
  assign new_n13074 = ~new_n13072 & ~new_n13073;
  assign new_n13075 = new_n5577 & ~new_n5580;
  assign new_n13076 = ~new_n5581 & ~new_n13075;
  assign new_n13077 = ~new_n13074 & new_n13076;
  assign new_n13078 = new_n13074 & ~new_n13076;
  assign new_n13079 = ~new_n13077 & ~new_n13078;
  assign new_n13080 = ~new_n13066 & ~new_n13079;
  assign new_n13081 = new_n13066 & new_n13079;
  assign new_n13082 = ~new_n13080 & ~new_n13081;
  assign new_n13083 = ~new_n5575 & new_n5585;
  assign new_n13084 = ~new_n5574 & ~new_n13083;
  assign new_n13085 = ~new_n13082 & ~new_n13084;
  assign new_n13086 = new_n13082 & new_n13084;
  assign new_n13087 = ~new_n13085 & ~new_n13086;
  assign new_n13088 = new_n13061 & new_n13087;
  assign new_n13089 = ~new_n13080 & new_n13084;
  assign new_n13090 = ~new_n13065 & ~new_n13089;
  assign new_n13091 = ~new_n13081 & new_n13090;
  assign new_n13092 = new_n13065 & new_n13089;
  assign new_n13093 = ~new_n13091 & ~new_n13092;
  assign new_n13094 = n1916 & n5684;
  assign new_n13095 = n8940 & n11429;
  assign new_n13096 = n4964 & n7374;
  assign new_n13097 = ~new_n13095 & ~new_n13096;
  assign new_n13098 = new_n13095 & new_n13096;
  assign new_n13099 = ~new_n13097 & ~new_n13098;
  assign new_n13100 = new_n13094 & ~new_n13099;
  assign new_n13101 = ~new_n13094 & new_n13099;
  assign new_n13102 = ~new_n13100 & ~new_n13101;
  assign new_n13103 = ~new_n13073 & new_n13076;
  assign new_n13104 = ~new_n13072 & ~new_n13103;
  assign new_n13105 = ~new_n13102 & new_n13104;
  assign new_n13106 = new_n13102 & ~new_n13104;
  assign new_n13107 = ~new_n13105 & ~new_n13106;
  assign new_n13108 = ~n10162 & new_n13071;
  assign new_n13109 = n10162 & n10770;
  assign new_n13110 = ~new_n13071 & new_n13109;
  assign new_n13111 = ~new_n13108 & ~new_n13110;
  assign new_n13112 = n8860 & n10522;
  assign new_n13113 = new_n13069 & new_n13112;
  assign new_n13114 = ~new_n13069 & ~new_n13112;
  assign new_n13115 = ~new_n13113 & ~new_n13114;
  assign new_n13116 = new_n13111 & ~new_n13115;
  assign new_n13117 = ~new_n13111 & new_n13115;
  assign new_n13118 = ~new_n13116 & ~new_n13117;
  assign new_n13119 = new_n13107 & ~new_n13118;
  assign new_n13120 = ~new_n13107 & new_n13118;
  assign new_n13121 = ~new_n13119 & ~new_n13120;
  assign new_n13122 = ~new_n13093 & new_n13121;
  assign new_n13123 = new_n13093 & ~new_n13121;
  assign new_n13124 = ~new_n13122 & ~new_n13123;
  assign new_n13125 = ~new_n13088 & ~new_n13124;
  assign new_n13126 = new_n13088 & new_n13124;
  assign new_n13127 = ~new_n13125 & ~new_n13126;
  assign new_n13128 = n7374 & n8940;
  assign new_n13129 = ~new_n13061 & ~new_n13087;
  assign new_n13130 = ~new_n13088 & ~new_n13129;
  assign new_n13131 = new_n13128 & new_n13130;
  assign new_n13132 = ~new_n13128 & ~new_n13130;
  assign new_n13133 = ~new_n13131 & ~new_n13132;
  assign new_n13134 = new_n5599 & new_n13133;
  assign new_n13135 = ~new_n13131 & ~new_n13134;
  assign new_n13136 = ~new_n13127 & new_n13135;
  assign new_n13137 = new_n13127 & ~new_n13135;
  assign new_n13138 = ~new_n13136 & ~new_n13137;
  assign new_n13139 = ~new_n5620 & new_n5624;
  assign new_n13140 = ~new_n5621 & ~new_n13139;
  assign new_n13141 = n3076 & n6333;
  assign new_n13142 = n1912 & n11634;
  assign new_n13143 = ~new_n13141 & ~new_n13142;
  assign new_n13144 = new_n13141 & new_n13142;
  assign new_n13145 = ~new_n13143 & ~new_n13144;
  assign new_n13146 = n817 & n12750;
  assign new_n13147 = n3815 & n9620;
  assign new_n13148 = n761 & n5548;
  assign new_n13149 = ~new_n13147 & ~new_n13148;
  assign new_n13150 = new_n13147 & new_n13148;
  assign new_n13151 = ~new_n13149 & ~new_n13150;
  assign new_n13152 = ~new_n13146 & ~new_n13151;
  assign new_n13153 = new_n13146 & new_n13151;
  assign new_n13154 = ~new_n13152 & ~new_n13153;
  assign new_n13155 = ~new_n5608 & ~new_n5612;
  assign new_n13156 = ~new_n5611 & ~new_n13155;
  assign new_n13157 = ~new_n13154 & ~new_n13156;
  assign new_n13158 = new_n13154 & new_n13156;
  assign new_n13159 = ~new_n13157 & ~new_n13158;
  assign new_n13160 = ~new_n13145 & ~new_n13159;
  assign new_n13161 = new_n13145 & new_n13159;
  assign new_n13162 = ~new_n13160 & ~new_n13161;
  assign new_n13163 = ~new_n5605 & ~new_n5616;
  assign new_n13164 = ~new_n5606 & ~new_n13163;
  assign new_n13165 = ~new_n13162 & ~new_n13164;
  assign new_n13166 = new_n13162 & new_n13164;
  assign new_n13167 = ~new_n13165 & ~new_n13166;
  assign new_n13168 = ~new_n13140 & ~new_n13167;
  assign new_n13169 = ~new_n13160 & ~new_n13164;
  assign new_n13170 = ~new_n13144 & ~new_n13169;
  assign new_n13171 = ~new_n13161 & new_n13170;
  assign new_n13172 = new_n13144 & new_n13169;
  assign new_n13173 = ~new_n13171 & ~new_n13172;
  assign new_n13174 = n1912 & n3076;
  assign new_n13175 = n7974 & n9353;
  assign new_n13176 = n6333 & n8163;
  assign new_n13177 = ~new_n13175 & ~new_n13176;
  assign new_n13178 = new_n13175 & new_n13176;
  assign new_n13179 = ~new_n13177 & ~new_n13178;
  assign new_n13180 = new_n13174 & ~new_n13179;
  assign new_n13181 = ~new_n13174 & new_n13179;
  assign new_n13182 = ~new_n13180 & ~new_n13181;
  assign new_n13183 = ~new_n13153 & ~new_n13156;
  assign new_n13184 = ~new_n13152 & ~new_n13183;
  assign new_n13185 = new_n13182 & ~new_n13184;
  assign new_n13186 = n11634 & n12750;
  assign new_n13187 = new_n13150 & new_n13186;
  assign new_n13188 = ~new_n13150 & ~new_n13186;
  assign new_n13189 = ~new_n13187 & ~new_n13188;
  assign new_n13190 = n5548 & n5758;
  assign new_n13191 = n761 & n3815;
  assign new_n13192 = n817 & n9620;
  assign new_n13193 = ~new_n13191 & ~new_n13192;
  assign new_n13194 = new_n13191 & new_n13192;
  assign new_n13195 = ~new_n13193 & ~new_n13194;
  assign new_n13196 = new_n13190 & ~new_n13195;
  assign new_n13197 = ~new_n13190 & new_n13195;
  assign new_n13198 = ~new_n13196 & ~new_n13197;
  assign new_n13199 = new_n13189 & new_n13198;
  assign new_n13200 = ~new_n13189 & ~new_n13198;
  assign new_n13201_1 = ~new_n13199 & ~new_n13200;
  assign new_n13202 = new_n13185 & new_n13201_1;
  assign new_n13203 = ~new_n13182 & new_n13184;
  assign new_n13204 = ~new_n13201_1 & new_n13203;
  assign new_n13205 = ~new_n13185 & ~new_n13201_1;
  assign new_n13206 = ~new_n13203 & ~new_n13205;
  assign new_n13207 = ~new_n13204 & ~new_n13206;
  assign new_n13208 = ~new_n13202 & ~new_n13207;
  assign new_n13209 = new_n13173 & ~new_n13208;
  assign new_n13210 = ~new_n13173 & new_n13208;
  assign new_n13211 = ~new_n13209 & ~new_n13210;
  assign new_n13212 = ~new_n13168 & new_n13211;
  assign new_n13213 = new_n13168 & ~new_n13211;
  assign new_n13214 = ~new_n13212 & ~new_n13213;
  assign new_n13215 = n8163 & n9353;
  assign new_n13216 = new_n13140 & new_n13167;
  assign new_n13217 = ~new_n13168 & ~new_n13216;
  assign new_n13218 = new_n13215 & new_n13217;
  assign new_n13219 = ~new_n13215 & ~new_n13217;
  assign new_n13220 = ~new_n13218 & ~new_n13219;
  assign new_n13221 = new_n5629 & new_n13220;
  assign new_n13222 = ~new_n13218 & ~new_n13221;
  assign new_n13223 = ~new_n13214 & new_n13222;
  assign new_n13224 = new_n13214 & ~new_n13222;
  assign new_n13225 = ~new_n13223 & ~new_n13224;
  assign new_n13226 = ~new_n13138 & ~new_n13225;
  assign new_n13227 = ~new_n5599 & ~new_n13133;
  assign new_n13228 = ~new_n13134 & ~new_n13227;
  assign new_n13229 = ~new_n5629 & ~new_n13220;
  assign new_n13230 = ~new_n13221 & ~new_n13229;
  assign new_n13231 = new_n13228 & new_n13230;
  assign new_n13232 = ~new_n13228 & ~new_n13230;
  assign new_n13233 = ~new_n5631 & ~new_n5635;
  assign new_n13234 = ~new_n5632 & ~new_n13233;
  assign new_n13235 = ~new_n13232 & new_n13234;
  assign new_n13236 = ~new_n13231 & ~new_n13235;
  assign new_n13237 = new_n13226 & new_n13236;
  assign new_n13238 = new_n13138 & new_n13225;
  assign new_n13239 = new_n13236 & ~new_n13238;
  assign new_n13240 = ~new_n13226 & ~new_n13239;
  assign new_n13241 = ~new_n13237 & ~new_n13240;
  assign new_n13242 = ~new_n13236 & new_n13238;
  assign new_n13243 = ~new_n13241 & ~new_n13242;
  assign new_n13244 = new_n13060_1 & ~new_n13243;
  assign new_n13245 = ~new_n13060_1 & new_n13243;
  assign new_n13246 = ~new_n13244 & ~new_n13245;
  assign new_n13247 = ~new_n5568_1 & ~new_n13055;
  assign new_n13248 = ~new_n13056 & ~new_n13247;
  assign new_n13249 = ~new_n13231 & ~new_n13232;
  assign new_n13250 = ~new_n13234 & ~new_n13249;
  assign new_n13251 = ~new_n13231 & new_n13235;
  assign new_n13252 = ~new_n13250 & ~new_n13251;
  assign new_n13253 = new_n13248 & new_n13252;
  assign new_n13254 = ~new_n13248 & ~new_n13252;
  assign new_n13255 = ~new_n5639 & ~new_n5643;
  assign new_n13256 = ~new_n5640 & ~new_n13255;
  assign new_n13257 = ~new_n13254 & ~new_n13256;
  assign new_n13258 = ~new_n13253 & ~new_n13257;
  assign new_n13259 = new_n13246 & new_n13258;
  assign new_n13260 = ~new_n13246 & ~new_n13258;
  assign new_n13261 = ~new_n13259 & ~new_n13260;
  assign new_n13262 = new_n12973 & ~new_n13261;
  assign new_n13263 = ~new_n12973 & new_n13261;
  assign new_n13264 = ~new_n13262 & ~new_n13263;
  assign new_n13265 = ~new_n5450 & ~new_n12968_1;
  assign new_n13266 = ~new_n12969 & ~new_n13265;
  assign new_n13267 = ~new_n5538 & new_n5646;
  assign new_n13268 = ~new_n5537 & ~new_n13267;
  assign new_n13269 = new_n13266 & new_n13268;
  assign new_n13270 = ~new_n13266 & ~new_n13268;
  assign new_n13271 = ~new_n13253 & ~new_n13254;
  assign new_n13272 = new_n13256 & ~new_n13271;
  assign new_n13273 = ~new_n13256 & new_n13271;
  assign new_n13274 = ~new_n13272 & ~new_n13273;
  assign new_n13275 = ~new_n13270 & new_n13274;
  assign new_n13276 = ~new_n13269 & ~new_n13275;
  assign new_n13277 = new_n13264 & new_n13276;
  assign new_n13278 = ~new_n13264 & ~new_n13276;
  assign n9872 = new_n13277 | new_n13278;
  assign new_n13280 = ~new_n2637 & ~new_n2639;
  assign n10101 = ~new_n2640 & ~new_n13280;
  assign new_n13282 = ~new_n12443 & ~new_n12444;
  assign new_n13283 = ~new_n12466 & ~new_n13282;
  assign new_n13284 = new_n12466 & new_n13282;
  assign n10243 = ~new_n13283 & ~new_n13284;
  assign new_n13286 = ~new_n1989 & ~new_n1990;
  assign new_n13287 = ~new_n1994 & ~new_n13286;
  assign new_n13288 = new_n1994 & new_n13286;
  assign n10453 = new_n13287 | new_n13288;
  assign new_n13290 = new_n13111 & ~new_n13113;
  assign new_n13291 = ~new_n13114 & ~new_n13290;
  assign new_n13292 = ~new_n13244 & new_n13258;
  assign new_n13293 = ~new_n13245 & ~new_n13292;
  assign new_n13294 = new_n13291 & new_n13293;
  assign new_n13295 = ~new_n13291 & ~new_n13293;
  assign new_n13296 = ~new_n13294 & ~new_n13295;
  assign new_n13297 = ~new_n13006 & ~new_n13043;
  assign new_n13298 = ~new_n13007 & ~new_n13297;
  assign new_n13299 = n761 & n817;
  assign new_n13300 = n4075 & n8940;
  assign new_n13301 = ~new_n13299 & new_n13300;
  assign new_n13302 = new_n13299 & ~new_n13300;
  assign new_n13303 = ~new_n13301 & ~new_n13302;
  assign new_n13304 = new_n13298 & new_n13303;
  assign new_n13305 = ~new_n13298 & ~new_n13303;
  assign new_n13306 = ~new_n13304 & ~new_n13305;
  assign new_n13307 = n2482 & n10122;
  assign new_n13308 = new_n13025 & ~new_n13028;
  assign new_n13309 = ~new_n13029 & ~new_n13308;
  assign new_n13310 = ~new_n13307 & new_n13309;
  assign new_n13311 = new_n13307 & ~new_n13309;
  assign new_n13312 = ~new_n13310 & ~new_n13311;
  assign new_n13313 = n11236 & n11835;
  assign new_n13314 = n5729 & n8820;
  assign new_n13315 = new_n13313 & ~new_n13314;
  assign new_n13316 = ~new_n13313 & new_n13314;
  assign new_n13317 = ~new_n13315 & ~new_n13316;
  assign new_n13318 = n8860 & n10770;
  assign new_n13319 = n1916 & n10522;
  assign new_n13320 = ~new_n13318 & ~new_n13319;
  assign new_n13321 = new_n13318 & new_n13319;
  assign new_n13322 = ~new_n13320 & ~new_n13321;
  assign new_n13323 = ~new_n13317 & ~new_n13322;
  assign new_n13324 = new_n13317 & new_n13322;
  assign new_n13325 = ~new_n13323 & ~new_n13324;
  assign new_n13326 = n3130 & n5065;
  assign new_n13327 = n5548 & n12352;
  assign new_n13328 = ~new_n13326 & new_n13327;
  assign new_n13329 = new_n13326 & ~new_n13327;
  assign new_n13330 = ~new_n13328 & ~new_n13329;
  assign new_n13331 = n443 & n4382;
  assign new_n13332 = n3815 & n5758;
  assign new_n13333 = new_n13331 & ~new_n13332;
  assign new_n13334 = ~new_n13331 & new_n13332;
  assign new_n13335 = ~new_n13333 & ~new_n13334;
  assign new_n13336 = ~new_n13330 & new_n13335;
  assign new_n13337 = new_n13330 & ~new_n13335;
  assign new_n13338 = ~new_n13336 & ~new_n13337;
  assign new_n13339 = ~new_n13325 & new_n13338;
  assign new_n13340 = new_n13325 & ~new_n13338;
  assign new_n13341 = ~new_n13339 & ~new_n13340;
  assign new_n13342 = ~new_n13312 & new_n13341;
  assign new_n13343 = new_n13312 & ~new_n13341;
  assign new_n13344 = ~new_n13342 & ~new_n13343;
  assign new_n13345 = n4964 & n11429;
  assign new_n13346 = n5684 & n7374;
  assign new_n13347 = ~new_n13345 & new_n13346;
  assign new_n13348 = new_n13345 & ~new_n13346;
  assign new_n13349 = ~new_n13347 & ~new_n13348;
  assign new_n13350 = n1757 & n9747;
  assign new_n13351 = n5884 & n10113;
  assign new_n13352 = n1709 & n9353;
  assign new_n13353 = new_n13351 & new_n13352;
  assign new_n13354 = ~new_n13351 & ~new_n13352;
  assign new_n13355 = ~new_n13353 & ~new_n13354;
  assign new_n13356 = new_n13350 & ~new_n13355;
  assign new_n13357 = ~new_n13350 & new_n13355;
  assign new_n13358 = ~new_n13356 & ~new_n13357;
  assign new_n13359 = ~new_n13349 & ~new_n13358;
  assign new_n13360 = new_n13349 & new_n13358;
  assign new_n13361 = ~new_n13359 & ~new_n13360;
  assign new_n13362 = n7659 & n11488;
  assign new_n13363 = n1982 & n12289;
  assign new_n13364 = ~new_n13362 & ~new_n13363;
  assign new_n13365 = new_n13362 & new_n13363;
  assign new_n13366 = ~new_n13364 & ~new_n13365;
  assign new_n13367 = n4330 & n11030;
  assign new_n13368 = n2252 & n10416;
  assign new_n13369 = new_n13367 & ~new_n13368;
  assign new_n13370 = ~new_n13367 & new_n13368;
  assign new_n13371 = ~new_n13369 & ~new_n13370;
  assign new_n13372 = ~new_n13366 & ~new_n13371;
  assign new_n13373 = new_n13366 & new_n13371;
  assign new_n13374 = ~new_n13372 & ~new_n13373;
  assign new_n13375 = new_n13361 & new_n13374;
  assign new_n13376 = ~new_n13361 & ~new_n13374;
  assign new_n13377 = ~new_n13375 & ~new_n13376;
  assign new_n13378 = new_n13344 & new_n13377;
  assign new_n13379 = ~new_n13344 & ~new_n13377;
  assign new_n13380 = ~new_n13378 & ~new_n13379;
  assign new_n13381 = ~new_n12935 & new_n12946;
  assign new_n13382 = ~new_n12936 & ~new_n13381;
  assign new_n13383 = n9620 & n11634;
  assign new_n13384 = n3076 & n12750;
  assign new_n13385 = ~new_n13383 & ~new_n13384;
  assign new_n13386 = new_n13383 & new_n13384;
  assign new_n13387 = ~new_n13385 & ~new_n13386;
  assign new_n13388 = n6333 & n7974;
  assign new_n13389 = n1912 & n8163;
  assign new_n13390 = new_n13388 & ~new_n13389;
  assign new_n13391 = ~new_n13388 & new_n13389;
  assign new_n13392 = ~new_n13390 & ~new_n13391;
  assign new_n13393 = ~new_n13387 & new_n13392;
  assign new_n13394 = new_n13387 & ~new_n13392;
  assign new_n13395 = ~new_n13393 & ~new_n13394;
  assign new_n13396 = ~new_n13382 & new_n13395;
  assign new_n13397 = new_n13382 & ~new_n13395;
  assign new_n13398 = ~new_n13396 & ~new_n13397;
  assign new_n13399 = new_n13380 & new_n13398;
  assign new_n13400 = ~new_n13380 & ~new_n13398;
  assign new_n13401 = ~new_n13399 & ~new_n13400;
  assign new_n13402 = new_n13306 & ~new_n13401;
  assign new_n13403 = ~new_n13306 & new_n13401;
  assign new_n13404 = ~new_n13402 & ~new_n13403;
  assign new_n13405 = n5320 & n5920;
  assign new_n13406 = n5356 & n8228;
  assign new_n13407 = ~new_n13405 & new_n13406;
  assign new_n13408 = new_n13405 & ~new_n13406;
  assign new_n13409 = ~new_n13407 & ~new_n13408;
  assign new_n13410 = n103 & n4862;
  assign new_n13411 = n1636 & n9732;
  assign new_n13412 = ~new_n13410 & ~new_n13411;
  assign new_n13413 = new_n13410 & new_n13411;
  assign new_n13414 = ~new_n13412 & ~new_n13413;
  assign new_n13415 = ~new_n13409 & new_n13414;
  assign new_n13416 = new_n13409 & ~new_n13414;
  assign new_n13417 = ~new_n13415 & ~new_n13416;
  assign new_n13418 = n4743 & n13058;
  assign new_n13419 = new_n13111 & new_n13418;
  assign new_n13420 = ~new_n13111 & ~new_n13418;
  assign new_n13421 = ~new_n13419 & ~new_n13420;
  assign new_n13422 = ~new_n13187 & new_n13198;
  assign new_n13423 = ~new_n13188 & ~new_n13422;
  assign new_n13424 = ~new_n13421 & new_n13423;
  assign new_n13425 = new_n13421 & ~new_n13423;
  assign new_n13426 = ~new_n13424 & ~new_n13425;
  assign new_n13427 = new_n13417 & new_n13426;
  assign new_n13428 = ~new_n13417 & ~new_n13426;
  assign new_n13429 = ~new_n13427 & ~new_n13428;
  assign new_n13430 = new_n13404 & ~new_n13429;
  assign new_n13431 = ~new_n13404 & new_n13429;
  assign new_n13432 = ~new_n13430 & ~new_n13431;
  assign new_n13433 = ~new_n13240 & ~new_n13432;
  assign new_n13434 = new_n13240 & new_n13432;
  assign new_n13435 = ~new_n13433 & ~new_n13434;
  assign new_n13436 = new_n13206 & ~new_n13435;
  assign new_n13437 = ~new_n13206 & new_n13435;
  assign new_n13438 = ~new_n13436 & ~new_n13437;
  assign new_n13439 = new_n12922 & ~new_n12925;
  assign new_n13440 = ~new_n12926 & ~new_n13439;
  assign new_n13441 = ~new_n13438 & new_n13440;
  assign new_n13442 = new_n13438 & ~new_n13440;
  assign new_n13443 = ~new_n13441 & ~new_n13442;
  assign new_n13444 = ~new_n13126 & ~new_n13137;
  assign new_n13445 = ~new_n12919 & new_n12956;
  assign new_n13446 = ~new_n12920 & ~new_n13445;
  assign new_n13447 = n10162 & ~new_n13070;
  assign new_n13448 = ~new_n13069 & ~new_n13447;
  assign new_n13449 = new_n13190 & ~new_n13193;
  assign new_n13450 = ~new_n13194 & ~new_n13449;
  assign new_n13451 = ~new_n13448 & new_n13450;
  assign new_n13452 = new_n13448 & ~new_n13450;
  assign new_n13453 = ~new_n13451 & ~new_n13452;
  assign new_n13454 = ~new_n13040 & ~new_n13453;
  assign new_n13455 = new_n13040 & new_n13453;
  assign new_n13456 = ~new_n13454 & ~new_n13455;
  assign new_n13457 = new_n13446 & ~new_n13456;
  assign new_n13458 = ~new_n13446 & new_n13456;
  assign new_n13459 = ~new_n13457 & ~new_n13458;
  assign new_n13460 = new_n12954 & ~new_n13459;
  assign new_n13461 = ~new_n12954 & new_n13459;
  assign new_n13462 = ~new_n13460 & ~new_n13461;
  assign new_n13463 = new_n13444 & new_n13462;
  assign new_n13464 = ~new_n13444 & ~new_n13462;
  assign new_n13465 = ~new_n13463 & ~new_n13464;
  assign new_n13466 = ~new_n13443 & new_n13465;
  assign new_n13467 = new_n13443 & ~new_n13465;
  assign new_n13468 = ~new_n13466 & ~new_n13467;
  assign new_n13469 = ~new_n13296 & ~new_n13468;
  assign new_n13470 = new_n13296 & new_n13468;
  assign new_n13471 = ~new_n13469 & ~new_n13470;
  assign new_n13472 = ~new_n13262 & new_n13276;
  assign new_n13473 = ~new_n13263 & ~new_n13472;
  assign new_n13474 = ~new_n13048 & ~new_n13059;
  assign new_n13475 = ~new_n13091 & ~new_n13121;
  assign new_n13476 = ~new_n13092 & ~new_n13475;
  assign new_n13477 = new_n13094 & ~new_n13097;
  assign new_n13478 = ~new_n13098 & ~new_n13477;
  assign new_n13479 = ~new_n13106 & new_n13118;
  assign new_n13480 = ~new_n13105 & ~new_n13479;
  assign new_n13481 = new_n12938 & ~new_n12941;
  assign new_n13482 = ~new_n12942 & ~new_n13481;
  assign new_n13483 = new_n13009 & ~new_n13012;
  assign new_n13484 = ~new_n13013 & ~new_n13483;
  assign new_n13485 = ~new_n13482 & new_n13484;
  assign new_n13486 = new_n13482 & ~new_n13484;
  assign new_n13487 = ~new_n13485 & ~new_n13486;
  assign new_n13488 = new_n13480 & ~new_n13487;
  assign new_n13489 = ~new_n13480 & new_n13487;
  assign new_n13490 = ~new_n13488 & ~new_n13489;
  assign new_n13491 = ~new_n13478 & new_n13490;
  assign new_n13492 = new_n13478 & ~new_n13490;
  assign new_n13493 = ~new_n13491 & ~new_n13492;
  assign new_n13494 = new_n13476 & ~new_n13493;
  assign new_n13495 = ~new_n13476 & new_n13493;
  assign new_n13496 = ~new_n13494 & ~new_n13495;
  assign new_n13497 = ~new_n13474 & new_n13496;
  assign new_n13498 = new_n13474 & ~new_n13496;
  assign new_n13499 = ~new_n13497 & ~new_n13498;
  assign new_n13500 = ~new_n12961 & ~new_n12972;
  assign new_n13501 = ~new_n13023 & ~new_n13033;
  assign new_n13502 = ~new_n13022 & ~new_n13501;
  assign new_n13503 = ~new_n13500 & new_n13502;
  assign new_n13504 = new_n13500 & ~new_n13502;
  assign new_n13505 = ~new_n13503 & ~new_n13504;
  assign new_n13506 = ~new_n13213 & ~new_n13224;
  assign new_n13507 = ~new_n13171 & new_n13208;
  assign new_n13508 = ~new_n13172 & ~new_n13507;
  assign new_n13509 = new_n13174 & ~new_n13177;
  assign new_n13510 = ~new_n13178 & ~new_n13509;
  assign new_n13511 = ~new_n13508 & new_n13510;
  assign new_n13512 = new_n13508 & ~new_n13510;
  assign new_n13513 = ~new_n13511 & ~new_n13512;
  assign new_n13514 = new_n13506 & new_n13513;
  assign new_n13515 = ~new_n13506 & ~new_n13513;
  assign new_n13516 = ~new_n13514 & ~new_n13515;
  assign new_n13517 = new_n13505 & new_n13516;
  assign new_n13518 = ~new_n13505 & ~new_n13516;
  assign new_n13519 = ~new_n13517 & ~new_n13518;
  assign new_n13520 = new_n13499 & ~new_n13519;
  assign new_n13521 = ~new_n13499 & new_n13519;
  assign new_n13522 = ~new_n13520 & ~new_n13521;
  assign new_n13523 = ~new_n13473 & new_n13522;
  assign new_n13524 = new_n13473 & ~new_n13522;
  assign new_n13525 = ~new_n13523 & ~new_n13524;
  assign new_n13526 = new_n13471 & ~new_n13525;
  assign new_n13527 = ~new_n13471 & new_n13525;
  assign n10524 = ~new_n13526 & ~new_n13527;
  assign new_n13529 = new_n9337 & ~new_n9344;
  assign new_n13530 = ~new_n9341 & new_n13529;
  assign new_n13531 = new_n9341 & ~new_n13529;
  assign n10628 = new_n13530 | new_n13531;
  assign new_n13533 = n2482 & n7411;
  assign new_n13534 = n1757 & n11734;
  assign new_n13535 = n10416 & new_n13534;
  assign new_n13536 = ~n10416 & ~new_n13534;
  assign new_n13537 = ~new_n13535 & ~new_n13536;
  assign new_n13538 = n11030 & ~new_n13537;
  assign new_n13539 = ~n11030 & new_n13537;
  assign new_n13540 = ~new_n13538 & ~new_n13539;
  assign new_n13541 = n10113 & n12651;
  assign new_n13542 = n10416 & ~new_n10472;
  assign new_n13543 = ~new_n10471 & ~new_n13542;
  assign new_n13544 = ~new_n13541 & new_n13543;
  assign new_n13545 = new_n13541 & ~new_n13543;
  assign new_n13546 = ~new_n13544 & ~new_n13545;
  assign new_n13547 = ~new_n13540 & new_n13546;
  assign new_n13548 = new_n13540 & ~new_n13546;
  assign new_n13549 = ~new_n13547 & ~new_n13548;
  assign new_n13550 = ~new_n13533 & ~new_n13549;
  assign new_n13551 = new_n13533 & new_n13549;
  assign new_n13552 = ~new_n10476 & ~new_n10479;
  assign new_n13553 = ~new_n10480 & ~new_n13552;
  assign new_n13554 = ~new_n13551 & new_n13553;
  assign new_n13555 = ~new_n13550 & ~new_n13554;
  assign new_n13556 = n1757 & n12651;
  assign new_n13557 = n7411 & n10113;
  assign new_n13558 = ~new_n13556 & ~new_n13557;
  assign new_n13559 = new_n13556 & new_n13557;
  assign new_n13560 = ~new_n13558 & ~new_n13559;
  assign new_n13561 = n10416 & n11734;
  assign new_n13562 = n11030 & n11488;
  assign new_n13563 = ~n11030 & ~n11488;
  assign new_n13564 = ~new_n13562 & ~new_n13563;
  assign new_n13565 = new_n13561 & new_n13564;
  assign new_n13566 = ~new_n13561 & ~new_n13564;
  assign new_n13567 = n11030 & ~new_n13536;
  assign new_n13568 = ~new_n13535 & ~new_n13567;
  assign new_n13569 = ~new_n13566 & ~new_n13568;
  assign new_n13570 = ~new_n13565 & new_n13569;
  assign new_n13571 = ~new_n13565 & ~new_n13566;
  assign new_n13572 = new_n13568 & ~new_n13571;
  assign new_n13573 = ~new_n13570 & ~new_n13572;
  assign new_n13574 = ~new_n13560 & ~new_n13573;
  assign new_n13575 = new_n13560 & new_n13573;
  assign new_n13576 = ~new_n13574 & ~new_n13575;
  assign new_n13577 = ~new_n13540 & ~new_n13544;
  assign new_n13578 = ~new_n13545 & ~new_n13577;
  assign new_n13579 = ~new_n13576 & ~new_n13578;
  assign new_n13580 = new_n13576 & new_n13578;
  assign new_n13581 = ~new_n13579 & ~new_n13580;
  assign new_n13582 = new_n13555 & ~new_n13581;
  assign new_n13583 = ~new_n13565 & ~new_n13569;
  assign new_n13584 = n1757 & n7411;
  assign new_n13585 = ~n7161 & n10113;
  assign new_n13586 = n2482 & n6149;
  assign new_n13587 = ~new_n13585 & ~new_n13586;
  assign new_n13588 = new_n13585 & new_n13586;
  assign new_n13589 = ~new_n13587 & ~new_n13588;
  assign new_n13590 = new_n13584 & ~new_n13589;
  assign new_n13591 = ~new_n13584 & new_n13589;
  assign new_n13592 = ~new_n13590 & ~new_n13591;
  assign new_n13593 = ~new_n13583 & ~new_n13592;
  assign new_n13594 = new_n13583 & new_n13592;
  assign new_n13595 = ~new_n13593 & ~new_n13594;
  assign new_n13596 = n10416 & n12651;
  assign new_n13597 = new_n13562 & new_n13596;
  assign new_n13598 = ~new_n13562 & ~new_n13596;
  assign new_n13599 = ~new_n13597 & ~new_n13598;
  assign new_n13600 = n11030 & n11734;
  assign new_n13601 = n11488 & new_n13600;
  assign new_n13602 = ~n11488 & ~new_n13600;
  assign new_n13603 = ~new_n13601 & ~new_n13602;
  assign new_n13604 = ~n1982 & ~new_n13603;
  assign new_n13605 = n1982 & ~new_n13602;
  assign new_n13606 = ~new_n13601 & new_n13605;
  assign new_n13607 = ~new_n13604 & ~new_n13606;
  assign new_n13608 = ~new_n13599 & ~new_n13607;
  assign new_n13609 = ~new_n13598 & new_n13607;
  assign new_n13610 = ~new_n13597 & new_n13609;
  assign new_n13611 = ~new_n13608 & ~new_n13610;
  assign new_n13612 = ~new_n13595 & new_n13611;
  assign new_n13613 = new_n13595 & ~new_n13611;
  assign new_n13614 = ~new_n13612 & ~new_n13613;
  assign new_n13615 = new_n13559 & ~new_n13614;
  assign new_n13616 = ~new_n13559 & new_n13614;
  assign new_n13617 = ~new_n13615 & ~new_n13616;
  assign new_n13618 = ~new_n13574 & ~new_n13578;
  assign new_n13619 = ~new_n13575 & ~new_n13618;
  assign new_n13620 = ~new_n13617 & new_n13619;
  assign new_n13621 = new_n13617 & ~new_n13619;
  assign new_n13622 = ~new_n13620 & ~new_n13621;
  assign new_n13623 = ~new_n13582 & ~new_n13622;
  assign new_n13624 = new_n13582 & new_n13622;
  assign new_n13625 = ~new_n13623 & ~new_n13624;
  assign new_n13626 = n2482 & ~n7161;
  assign new_n13627 = ~new_n13555 & new_n13581;
  assign new_n13628 = ~new_n13582 & ~new_n13627;
  assign new_n13629 = new_n13626 & new_n13628;
  assign new_n13630 = ~new_n13550 & ~new_n13551;
  assign new_n13631 = ~new_n13553 & ~new_n13630;
  assign new_n13632 = new_n13553 & new_n13630;
  assign new_n13633 = ~new_n13631 & ~new_n13632;
  assign new_n13634 = new_n10486 & ~new_n13633;
  assign new_n13635 = ~new_n13626 & ~new_n13628;
  assign new_n13636 = ~new_n13629 & ~new_n13635;
  assign new_n13637 = new_n13634 & new_n13636;
  assign new_n13638 = ~new_n13629 & ~new_n13637;
  assign new_n13639 = new_n13625 & ~new_n13638;
  assign new_n13640 = ~new_n13625 & new_n13638;
  assign new_n13641 = ~new_n13639 & ~new_n13640;
  assign new_n13642 = n469 & n11236;
  assign new_n13643 = n4382 & n12284;
  assign new_n13644 = ~new_n13642 & ~new_n13643;
  assign new_n13645 = new_n13642 & new_n13643;
  assign new_n13646 = ~new_n13644 & ~new_n13645;
  assign new_n13647 = n3130 & n6826;
  assign new_n13648 = n9475 & n9732;
  assign new_n13649 = n103 & n411;
  assign new_n13650 = ~new_n13648 & ~new_n13649;
  assign new_n13651 = new_n13648 & new_n13649;
  assign new_n13652 = ~new_n13650 & ~new_n13651;
  assign new_n13653 = ~new_n13647 & ~new_n13652;
  assign new_n13654 = new_n13647 & new_n13652;
  assign new_n13655 = ~new_n13653 & ~new_n13654;
  assign new_n13656 = n4382 & n6826;
  assign new_n13657 = n3130 & n9475;
  assign new_n13658 = new_n13656 & new_n13657;
  assign new_n13659 = n411 & n9732;
  assign new_n13660 = ~new_n13656 & ~new_n13657;
  assign new_n13661 = new_n13659 & ~new_n13660;
  assign new_n13662 = ~new_n13658 & ~new_n13661;
  assign new_n13663 = ~new_n13655 & new_n13662;
  assign new_n13664 = new_n13655 & ~new_n13662;
  assign new_n13665 = ~new_n13663 & ~new_n13664;
  assign new_n13666 = ~new_n13646 & ~new_n13665;
  assign new_n13667 = new_n13646 & new_n13665;
  assign new_n13668 = ~new_n13666 & ~new_n13667;
  assign new_n13669 = n11236 & n12284;
  assign new_n13670 = new_n10494 & ~new_n10497;
  assign new_n13671 = ~new_n10498 & ~new_n13670;
  assign new_n13672 = ~new_n13669 & new_n13671;
  assign new_n13673 = new_n13669 & ~new_n13671;
  assign new_n13674 = ~new_n13658 & ~new_n13660;
  assign new_n13675 = new_n13659 & ~new_n13674;
  assign new_n13676 = ~new_n13659 & new_n13674;
  assign new_n13677 = ~new_n13675 & ~new_n13676;
  assign new_n13678 = ~new_n13673 & new_n13677;
  assign new_n13679 = ~new_n13672 & ~new_n13678;
  assign new_n13680 = ~new_n13668 & ~new_n13679;
  assign new_n13681 = new_n13668 & new_n13679;
  assign new_n13682 = ~new_n13680 & ~new_n13681;
  assign new_n13683 = n469 & n8228;
  assign new_n13684 = ~new_n13672 & ~new_n13673;
  assign new_n13685 = new_n13677 & ~new_n13684;
  assign new_n13686 = ~new_n13677 & new_n13684;
  assign new_n13687 = ~new_n13685 & ~new_n13686;
  assign new_n13688 = new_n13683 & new_n13687;
  assign new_n13689 = ~new_n13683 & ~new_n13687;
  assign new_n13690 = ~new_n10492 & new_n10502;
  assign new_n13691 = ~new_n10491 & ~new_n13690;
  assign new_n13692 = ~new_n13689 & new_n13691;
  assign new_n13693 = ~new_n13688 & ~new_n13692;
  assign new_n13694 = new_n13682 & ~new_n13693;
  assign new_n13695 = ~new_n13666 & new_n13679;
  assign new_n13696 = ~new_n13645 & ~new_n13695;
  assign new_n13697 = ~new_n13667 & new_n13696;
  assign new_n13698 = new_n13645 & new_n13695;
  assign new_n13699 = ~new_n13697 & ~new_n13698;
  assign new_n13700 = n469 & n4382;
  assign new_n13701 = n8228 & n11180;
  assign new_n13702 = n11236 & n12065;
  assign new_n13703 = ~new_n13701 & ~new_n13702;
  assign new_n13704 = new_n13701 & new_n13702;
  assign new_n13705 = ~new_n13703 & ~new_n13704;
  assign new_n13706 = new_n13700 & ~new_n13705;
  assign new_n13707 = ~new_n13700 & new_n13705;
  assign new_n13708 = ~new_n13706 & ~new_n13707;
  assign new_n13709 = ~new_n13654 & new_n13662;
  assign new_n13710 = ~new_n13653 & ~new_n13709;
  assign new_n13711 = new_n13708 & ~new_n13710;
  assign new_n13712 = n3130 & n12284;
  assign new_n13713 = ~new_n13651 & ~new_n13712;
  assign new_n13714 = new_n13651 & new_n13712;
  assign new_n13715 = ~new_n13713 & ~new_n13714;
  assign new_n13716 = n411 & n5320;
  assign new_n13717 = n103 & n9475;
  assign new_n13718 = n6826 & n9732;
  assign new_n13719 = ~new_n13717 & ~new_n13718;
  assign new_n13720 = new_n13717 & new_n13718;
  assign new_n13721 = ~new_n13719 & ~new_n13720;
  assign new_n13722 = new_n13716 & ~new_n13721;
  assign new_n13723 = ~new_n13716 & new_n13721;
  assign new_n13724 = ~new_n13722 & ~new_n13723;
  assign new_n13725 = new_n13715 & new_n13724;
  assign new_n13726 = ~new_n13715 & ~new_n13724;
  assign new_n13727 = ~new_n13725 & ~new_n13726;
  assign new_n13728 = new_n13711 & new_n13727;
  assign new_n13729 = ~new_n13708 & new_n13710;
  assign new_n13730 = ~new_n13727 & new_n13729;
  assign new_n13731 = ~new_n13711 & ~new_n13727;
  assign new_n13732 = ~new_n13729 & ~new_n13731;
  assign new_n13733 = ~new_n13730 & ~new_n13732;
  assign new_n13734 = ~new_n13728 & ~new_n13733;
  assign new_n13735 = new_n13699 & ~new_n13734;
  assign new_n13736 = ~new_n13699 & new_n13734;
  assign new_n13737 = ~new_n13735 & ~new_n13736;
  assign new_n13738 = ~new_n13694 & new_n13737;
  assign new_n13739 = new_n13694 & ~new_n13737;
  assign new_n13740 = ~new_n13738 & ~new_n13739;
  assign new_n13741 = n8228 & n12065;
  assign new_n13742 = ~new_n13682 & new_n13693;
  assign new_n13743 = ~new_n13694 & ~new_n13742;
  assign new_n13744 = new_n13741 & new_n13743;
  assign new_n13745 = ~new_n13688 & ~new_n13689;
  assign new_n13746 = ~new_n13691 & ~new_n13745;
  assign new_n13747 = new_n13691 & new_n13745;
  assign new_n13748 = ~new_n13746 & ~new_n13747;
  assign new_n13749 = new_n10507 & new_n13748;
  assign new_n13750 = ~new_n13741 & ~new_n13743;
  assign new_n13751 = ~new_n13744 & ~new_n13750;
  assign new_n13752 = new_n13749 & new_n13751;
  assign new_n13753 = ~new_n13744 & ~new_n13752;
  assign new_n13754 = ~new_n13740 & new_n13753;
  assign new_n13755 = new_n13740 & ~new_n13753;
  assign new_n13756 = ~new_n13754 & ~new_n13755;
  assign new_n13757 = n4964 & n12408;
  assign new_n13758 = n2737 & n5684;
  assign new_n13759 = ~new_n13757 & ~new_n13758;
  assign new_n13760 = new_n13757 & new_n13758;
  assign new_n13761 = ~new_n13759 & ~new_n13760;
  assign new_n13762 = n772 & n10522;
  assign new_n13763 = n5536 & n10770;
  assign new_n13764 = n8506 & new_n13763;
  assign new_n13765 = n8506 & n10770;
  assign new_n13766 = ~new_n13763 & ~new_n13765;
  assign new_n13767 = ~new_n13764 & ~new_n13766;
  assign new_n13768 = ~new_n13762 & ~new_n13767;
  assign new_n13769 = new_n13762 & new_n13767;
  assign new_n13770 = ~new_n13768 & ~new_n13769;
  assign new_n13771 = n772 & n5684;
  assign new_n13772 = n5536 & n10522;
  assign new_n13773 = new_n13771 & new_n13772;
  assign new_n13774 = ~new_n13771 & ~new_n13772;
  assign new_n13775 = new_n13765 & ~new_n13774;
  assign new_n13776 = ~new_n13773 & ~new_n13775;
  assign new_n13777 = ~new_n13770 & new_n13776;
  assign new_n13778 = new_n13770 & ~new_n13776;
  assign new_n13779 = ~new_n13777 & ~new_n13778;
  assign new_n13780 = ~new_n13761 & ~new_n13779;
  assign new_n13781 = new_n13761 & new_n13779;
  assign new_n13782 = ~new_n13780 & ~new_n13781;
  assign new_n13783 = n2737 & n4964;
  assign new_n13784 = new_n10515 & ~new_n10518;
  assign new_n13785 = ~new_n10519 & ~new_n13784;
  assign new_n13786 = ~new_n13783 & new_n13785;
  assign new_n13787 = new_n13783 & ~new_n13785;
  assign new_n13788 = ~new_n13773 & ~new_n13774;
  assign new_n13789 = new_n13765 & ~new_n13788;
  assign new_n13790 = ~new_n13765 & new_n13788;
  assign new_n13791 = ~new_n13789 & ~new_n13790;
  assign new_n13792 = ~new_n13787 & new_n13791;
  assign new_n13793 = ~new_n13786 & ~new_n13792;
  assign new_n13794 = ~new_n13782 & ~new_n13793;
  assign new_n13795 = new_n13782 & new_n13793;
  assign new_n13796 = ~new_n13794 & ~new_n13795;
  assign new_n13797 = n8940 & n12408;
  assign new_n13798 = ~new_n13786 & ~new_n13787;
  assign new_n13799 = new_n13791 & ~new_n13798;
  assign new_n13800 = ~new_n13791 & new_n13798;
  assign new_n13801 = ~new_n13799 & ~new_n13800;
  assign new_n13802 = new_n13797 & new_n13801;
  assign new_n13803 = ~new_n13797 & ~new_n13801;
  assign new_n13804 = ~new_n10513 & new_n10523;
  assign new_n13805 = ~new_n10512 & ~new_n13804;
  assign new_n13806 = ~new_n13803 & new_n13805;
  assign new_n13807 = ~new_n13802 & ~new_n13806;
  assign new_n13808 = new_n13796 & ~new_n13807;
  assign new_n13809 = ~new_n13780 & new_n13793;
  assign new_n13810 = ~new_n13760 & ~new_n13809;
  assign new_n13811 = ~new_n13781 & new_n13810;
  assign new_n13812 = new_n13760 & new_n13809;
  assign new_n13813 = ~new_n13811 & ~new_n13812;
  assign new_n13814 = n5684 & n12408;
  assign new_n13815 = n8940 & n11350;
  assign new_n13816 = n4964 & n9846;
  assign new_n13817 = ~new_n13815 & ~new_n13816;
  assign new_n13818 = new_n13815 & new_n13816;
  assign new_n13819 = ~new_n13817 & ~new_n13818;
  assign new_n13820 = new_n13814 & ~new_n13819;
  assign new_n13821 = ~new_n13814 & new_n13819;
  assign new_n13822 = ~new_n13820 & ~new_n13821;
  assign new_n13823 = ~new_n13769 & new_n13776;
  assign new_n13824 = ~new_n13768 & ~new_n13823;
  assign new_n13825 = ~new_n13822 & new_n13824;
  assign new_n13826 = new_n13822 & ~new_n13824;
  assign new_n13827 = ~new_n13825 & ~new_n13826;
  assign new_n13828 = ~n772 & new_n13767;
  assign new_n13829 = n772 & n10770;
  assign new_n13830 = ~new_n13767 & new_n13829;
  assign new_n13831 = ~new_n13828 & ~new_n13830;
  assign new_n13832 = n2737 & n10522;
  assign new_n13833 = new_n13764 & new_n13832;
  assign new_n13834 = ~new_n13764 & ~new_n13832;
  assign new_n13835 = ~new_n13833 & ~new_n13834;
  assign new_n13836 = new_n13831 & ~new_n13835;
  assign new_n13837 = ~new_n13831 & new_n13835;
  assign new_n13838 = ~new_n13836 & ~new_n13837;
  assign new_n13839 = new_n13827 & ~new_n13838;
  assign new_n13840 = ~new_n13827 & new_n13838;
  assign new_n13841 = ~new_n13839 & ~new_n13840;
  assign new_n13842 = ~new_n13813 & new_n13841;
  assign new_n13843 = new_n13813 & ~new_n13841;
  assign new_n13844 = ~new_n13842 & ~new_n13843;
  assign new_n13845 = ~new_n13808 & ~new_n13844;
  assign new_n13846 = new_n13808 & new_n13844;
  assign new_n13847 = ~new_n13845 & ~new_n13846;
  assign new_n13848 = n8940 & n9846;
  assign new_n13849 = ~new_n13796 & new_n13807;
  assign new_n13850 = ~new_n13808 & ~new_n13849;
  assign new_n13851 = new_n13848 & new_n13850;
  assign new_n13852 = ~new_n13802 & ~new_n13803;
  assign new_n13853 = new_n13805 & new_n13852;
  assign new_n13854 = ~new_n13805 & ~new_n13852;
  assign new_n13855 = ~new_n13853 & ~new_n13854;
  assign new_n13856 = new_n10528 & new_n13855;
  assign new_n13857 = ~new_n13848 & ~new_n13850;
  assign new_n13858 = ~new_n13851 & ~new_n13857;
  assign new_n13859 = new_n13856 & new_n13858;
  assign new_n13860 = ~new_n13851 & ~new_n13859;
  assign new_n13861 = ~new_n13847 & new_n13860;
  assign new_n13862 = new_n13847 & ~new_n13860;
  assign new_n13863 = ~new_n13861 & ~new_n13862;
  assign new_n13864 = n353 & n6333;
  assign new_n13865 = n1912 & n12263;
  assign new_n13866 = ~new_n13864 & ~new_n13865;
  assign new_n13867 = new_n13864 & new_n13865;
  assign new_n13868 = ~new_n13866 & ~new_n13867;
  assign new_n13869 = n10805 & n12750;
  assign new_n13870 = n124 & n9620;
  assign new_n13871 = n761 & n3085;
  assign new_n13872 = ~new_n13870 & ~new_n13871;
  assign new_n13873 = new_n13870 & new_n13871;
  assign new_n13874 = ~new_n13872 & ~new_n13873;
  assign new_n13875 = new_n13869 & new_n13874;
  assign new_n13876 = ~new_n13869 & ~new_n13874;
  assign new_n13877 = ~new_n13875 & ~new_n13876;
  assign new_n13878 = n1912 & n10805;
  assign new_n13879 = n124 & n12750;
  assign new_n13880 = new_n13878 & new_n13879;
  assign new_n13881 = ~new_n13878 & ~new_n13879;
  assign new_n13882 = n3085 & n9620;
  assign new_n13883 = ~new_n13881 & new_n13882;
  assign new_n13884 = ~new_n13880 & ~new_n13883;
  assign new_n13885 = ~new_n13877 & new_n13884;
  assign new_n13886 = new_n13877 & ~new_n13884;
  assign new_n13887 = ~new_n13885 & ~new_n13886;
  assign new_n13888 = ~new_n13868 & ~new_n13887;
  assign new_n13889 = new_n13868 & new_n13887;
  assign new_n13890 = ~new_n13888 & ~new_n13889;
  assign new_n13891 = n6333 & n12263;
  assign new_n13892 = new_n10536 & ~new_n10539;
  assign new_n13893 = ~new_n10540 & ~new_n13892;
  assign new_n13894 = ~new_n13891 & new_n13893;
  assign new_n13895 = new_n13891 & ~new_n13893;
  assign new_n13896 = ~new_n13880 & ~new_n13881;
  assign new_n13897 = ~new_n13882 & ~new_n13896;
  assign new_n13898 = new_n13882 & new_n13896;
  assign new_n13899 = ~new_n13897 & ~new_n13898;
  assign new_n13900 = ~new_n13895 & ~new_n13899;
  assign new_n13901 = ~new_n13894 & ~new_n13900;
  assign new_n13902 = ~new_n13890 & new_n13901;
  assign new_n13903 = new_n13890 & ~new_n13901;
  assign new_n13904 = ~new_n13902 & ~new_n13903;
  assign new_n13905 = n353 & n9353;
  assign new_n13906 = ~new_n13894 & ~new_n13895;
  assign new_n13907 = ~new_n13899 & new_n13906;
  assign new_n13908 = new_n13899 & ~new_n13906;
  assign new_n13909 = ~new_n13907 & ~new_n13908;
  assign new_n13910 = new_n13905 & ~new_n13909;
  assign new_n13911 = ~new_n13905 & new_n13909;
  assign new_n13912 = ~new_n10534 & new_n10544;
  assign new_n13913 = ~new_n10533 & ~new_n13912;
  assign new_n13914 = ~new_n13911 & new_n13913;
  assign new_n13915 = ~new_n13910 & ~new_n13914;
  assign new_n13916 = ~new_n13904 & ~new_n13915;
  assign new_n13917 = ~new_n13888 & new_n13901;
  assign new_n13918 = ~new_n13867 & ~new_n13917;
  assign new_n13919 = ~new_n13889 & new_n13918;
  assign new_n13920 = new_n13867 & new_n13917;
  assign new_n13921 = ~new_n13919 & ~new_n13920;
  assign new_n13922 = n353 & n1912;
  assign new_n13923 = n9353 & n11396;
  assign new_n13924 = n22 & n6333;
  assign new_n13925 = ~new_n13923 & ~new_n13924;
  assign new_n13926 = new_n13923 & new_n13924;
  assign new_n13927 = ~new_n13925 & ~new_n13926;
  assign new_n13928 = new_n13922 & ~new_n13927;
  assign new_n13929 = ~new_n13922 & new_n13927;
  assign new_n13930 = ~new_n13928 & ~new_n13929;
  assign new_n13931 = ~new_n13875 & new_n13884;
  assign new_n13932 = ~new_n13876 & ~new_n13931;
  assign new_n13933 = new_n13930 & ~new_n13932;
  assign new_n13934 = n12263 & n12750;
  assign new_n13935 = new_n13873 & new_n13934;
  assign new_n13936 = ~new_n13873 & ~new_n13934;
  assign new_n13937 = ~new_n13935 & ~new_n13936;
  assign new_n13938 = n3085 & n5758;
  assign new_n13939 = n124 & n761;
  assign new_n13940 = n9620 & n10805;
  assign new_n13941 = ~new_n13939 & ~new_n13940;
  assign new_n13942 = new_n13939 & new_n13940;
  assign new_n13943 = ~new_n13941 & ~new_n13942;
  assign new_n13944 = new_n13938 & ~new_n13943;
  assign new_n13945 = ~new_n13938 & new_n13943;
  assign new_n13946 = ~new_n13944 & ~new_n13945;
  assign new_n13947 = new_n13937 & new_n13946;
  assign new_n13948 = ~new_n13937 & ~new_n13946;
  assign new_n13949 = ~new_n13947 & ~new_n13948;
  assign new_n13950 = new_n13933 & new_n13949;
  assign new_n13951 = ~new_n13930 & new_n13932;
  assign new_n13952 = ~new_n13949 & new_n13951;
  assign new_n13953 = ~new_n13933 & ~new_n13949;
  assign new_n13954 = ~new_n13951 & ~new_n13953;
  assign new_n13955 = ~new_n13952 & ~new_n13954;
  assign new_n13956 = ~new_n13950 & ~new_n13955;
  assign new_n13957 = ~new_n13921 & ~new_n13956;
  assign new_n13958 = new_n13921 & new_n13956;
  assign new_n13959 = ~new_n13957 & ~new_n13958;
  assign new_n13960 = ~new_n13916 & ~new_n13959;
  assign new_n13961 = new_n13916 & new_n13959;
  assign new_n13962 = ~new_n13960 & ~new_n13961;
  assign new_n13963 = n22 & n9353;
  assign new_n13964 = new_n13904 & new_n13915;
  assign new_n13965 = ~new_n13916 & ~new_n13964;
  assign new_n13966 = new_n13963 & new_n13965;
  assign new_n13967 = ~new_n13910 & ~new_n13911;
  assign new_n13968 = new_n13913 & new_n13967;
  assign new_n13969 = ~new_n13913 & ~new_n13967;
  assign new_n13970 = ~new_n13968 & ~new_n13969;
  assign new_n13971 = new_n10548 & new_n13970;
  assign new_n13972 = ~new_n13963 & ~new_n13965;
  assign new_n13973 = ~new_n13966 & ~new_n13972;
  assign new_n13974 = new_n13971 & new_n13973;
  assign new_n13975 = ~new_n13966 & ~new_n13974;
  assign new_n13976 = ~new_n13962 & new_n13975;
  assign new_n13977 = new_n13962 & ~new_n13975;
  assign new_n13978 = ~new_n13976 & ~new_n13977;
  assign new_n13979 = ~new_n13863 & ~new_n13978;
  assign new_n13980 = ~new_n13971 & ~new_n13973;
  assign new_n13981 = ~new_n13974 & ~new_n13980;
  assign new_n13982 = ~new_n13856 & ~new_n13858;
  assign new_n13983 = ~new_n13859 & ~new_n13982;
  assign new_n13984 = new_n13981 & new_n13983;
  assign new_n13985 = ~new_n13981 & ~new_n13983;
  assign new_n13986 = ~new_n10528 & ~new_n13855;
  assign new_n13987 = ~new_n13856 & ~new_n13986;
  assign new_n13988 = ~new_n10548 & ~new_n13970;
  assign new_n13989 = ~new_n13971 & ~new_n13988;
  assign new_n13990 = new_n13987 & new_n13989;
  assign new_n13991 = ~new_n13987 & ~new_n13989;
  assign new_n13992 = ~new_n10552 & ~new_n10555;
  assign new_n13993 = ~new_n10551 & ~new_n13992;
  assign new_n13994 = ~new_n13991 & ~new_n13993;
  assign new_n13995 = ~new_n13990 & ~new_n13994;
  assign new_n13996 = ~new_n13985 & ~new_n13995;
  assign new_n13997 = ~new_n13984 & ~new_n13996;
  assign new_n13998 = new_n13979 & new_n13997;
  assign new_n13999 = new_n13863 & new_n13978;
  assign new_n14000 = ~new_n13997 & new_n13999;
  assign new_n14001 = ~new_n13979 & ~new_n13997;
  assign new_n14002 = ~new_n13999 & ~new_n14001;
  assign new_n14003 = ~new_n14000 & ~new_n14002;
  assign new_n14004 = ~new_n13998 & ~new_n14003;
  assign new_n14005 = new_n13756 & new_n14004;
  assign new_n14006 = ~new_n13756 & ~new_n14004;
  assign new_n14007 = ~new_n14005 & ~new_n14006;
  assign new_n14008 = ~new_n13749 & ~new_n13751;
  assign new_n14009 = ~new_n13752 & ~new_n14008;
  assign new_n14010 = ~new_n10507 & ~new_n13748;
  assign new_n14011 = ~new_n13749 & ~new_n14010;
  assign new_n14012 = ~new_n13990 & ~new_n13991;
  assign new_n14013 = new_n13993 & ~new_n14012;
  assign new_n14014 = ~new_n13993 & new_n14012;
  assign new_n14015 = ~new_n14013 & ~new_n14014;
  assign new_n14016 = ~new_n14011 & ~new_n14015;
  assign new_n14017 = new_n14011 & new_n14015;
  assign new_n14018 = ~new_n10559 & ~new_n10563;
  assign new_n14019 = ~new_n10560_1 & ~new_n14018;
  assign new_n14020 = ~new_n14017 & ~new_n14019;
  assign new_n14021 = ~new_n14016 & ~new_n14020;
  assign new_n14022 = new_n14009 & new_n14021;
  assign new_n14023 = ~new_n14009 & ~new_n14021;
  assign new_n14024 = ~new_n13984 & ~new_n13985;
  assign new_n14025 = new_n13995 & ~new_n14024;
  assign new_n14026 = ~new_n13995 & new_n14024;
  assign new_n14027 = ~new_n14025 & ~new_n14026;
  assign new_n14028 = ~new_n14023 & new_n14027;
  assign new_n14029 = ~new_n14022 & ~new_n14028;
  assign new_n14030 = ~new_n14007 & new_n14029;
  assign new_n14031 = new_n14007 & ~new_n14029;
  assign new_n14032 = ~new_n14030 & ~new_n14031;
  assign new_n14033 = ~new_n13641 & ~new_n14032;
  assign new_n14034 = ~new_n13634 & ~new_n13636;
  assign new_n14035 = ~new_n13637 & ~new_n14034;
  assign new_n14036 = ~new_n10486 & new_n13633;
  assign new_n14037 = ~new_n13634 & ~new_n14036;
  assign new_n14038 = ~new_n14016 & ~new_n14017;
  assign new_n14039 = new_n14019 & ~new_n14038;
  assign new_n14040 = ~new_n14019 & new_n14038;
  assign new_n14041 = ~new_n14039 & ~new_n14040;
  assign new_n14042 = ~new_n14037 & new_n14041;
  assign new_n14043 = new_n14037 & ~new_n14041;
  assign new_n14044 = ~new_n10469 & ~new_n10567;
  assign new_n14045 = ~new_n10568 & ~new_n14044;
  assign new_n14046 = ~new_n14043 & new_n14045;
  assign new_n14047 = ~new_n14042 & ~new_n14046;
  assign new_n14048 = new_n14035 & new_n14047;
  assign new_n14049 = ~new_n14035 & ~new_n14047;
  assign new_n14050 = ~new_n14022 & ~new_n14023;
  assign new_n14051 = new_n14027 & new_n14050;
  assign new_n14052 = ~new_n14027 & ~new_n14050;
  assign new_n14053 = ~new_n14051 & ~new_n14052;
  assign new_n14054 = ~new_n14049 & new_n14053;
  assign new_n14055 = ~new_n14048 & ~new_n14054;
  assign new_n14056 = new_n14033 & new_n14055;
  assign new_n14057 = new_n13641 & new_n14032;
  assign new_n14058 = ~new_n14055 & new_n14057;
  assign new_n14059 = ~new_n14033 & ~new_n14055;
  assign new_n14060 = ~new_n14057 & ~new_n14059;
  assign new_n14061 = ~new_n14058 & ~new_n14060;
  assign n10736 = ~new_n14056 & ~new_n14061;
  assign new_n14063 = ~new_n1378 & ~new_n1380;
  assign n10797 = ~new_n1381 & ~new_n14063;
  assign new_n14065 = ~new_n8653 & ~new_n8654;
  assign new_n14066 = new_n8668 & ~new_n14065;
  assign new_n14067 = ~new_n8668 & new_n14065;
  assign n11057 = ~new_n14066 & ~new_n14067;
  assign new_n14069 = ~new_n12692 & ~new_n12693_1;
  assign new_n14070 = ~new_n12703 & ~new_n14069;
  assign new_n14071 = new_n12703 & new_n14069;
  assign n11077 = ~new_n14070 & ~new_n14071;
  assign new_n14073 = ~new_n6038 & ~new_n6039;
  assign new_n14074 = new_n6053 & ~new_n14073;
  assign new_n14075 = ~new_n6053 & new_n14073;
  assign n11140 = new_n14074 | new_n14075;
  assign new_n14077 = ~new_n8645 & ~new_n8646;
  assign new_n14078 = new_n8670 & ~new_n14077;
  assign new_n14079 = ~new_n8670 & new_n14077;
  assign n11147 = ~new_n14078 & ~new_n14079;
  assign new_n14081 = ~new_n14006 & ~new_n14029;
  assign new_n14082 = ~new_n14005 & ~new_n14081;
  assign new_n14083 = ~new_n13697 & new_n13734;
  assign new_n14084 = ~new_n13698 & ~new_n14083;
  assign new_n14085 = ~new_n13597 & ~new_n13609;
  assign new_n14086 = ~new_n13954 & ~new_n14085;
  assign new_n14087 = new_n13954 & new_n14085;
  assign new_n14088 = ~new_n14086 & ~new_n14087;
  assign new_n14089 = ~new_n13732 & new_n14088;
  assign new_n14090 = new_n13732 & ~new_n14088;
  assign new_n14091 = ~new_n14089 & ~new_n14090;
  assign new_n14092 = new_n14084 & ~new_n14091;
  assign new_n14093 = ~new_n14084 & new_n14091;
  assign new_n14094 = ~new_n14092 & ~new_n14093;
  assign new_n14095 = ~new_n13739 & ~new_n13755;
  assign new_n14096 = ~new_n13846 & ~new_n13862;
  assign new_n14097 = ~new_n14095 & new_n14096;
  assign new_n14098 = new_n14095 & ~new_n14096;
  assign new_n14099 = ~new_n14097 & ~new_n14098;
  assign new_n14100 = ~new_n13919 & new_n13956;
  assign new_n14101 = ~new_n13920 & ~new_n14100;
  assign new_n14102 = ~new_n13961 & ~new_n13977;
  assign new_n14103 = new_n14101 & new_n14102;
  assign new_n14104 = ~new_n14101 & ~new_n14102;
  assign new_n14105 = ~new_n14103 & ~new_n14104;
  assign new_n14106 = new_n14099 & ~new_n14105;
  assign new_n14107 = ~new_n14099 & new_n14105;
  assign new_n14108 = ~new_n14106 & ~new_n14107;
  assign new_n14109 = ~new_n14094 & new_n14108;
  assign new_n14110 = new_n14094 & ~new_n14108;
  assign new_n14111 = ~new_n14109 & ~new_n14110;
  assign new_n14112 = new_n14082 & new_n14111;
  assign new_n14113 = ~new_n14082 & ~new_n14111;
  assign new_n14114 = ~new_n14112 & ~new_n14113;
  assign new_n14115 = n772 & ~new_n13766;
  assign new_n14116 = ~new_n13764 & ~new_n14115;
  assign new_n14117 = ~new_n13935 & new_n13946;
  assign new_n14118 = ~new_n13936 & ~new_n14117;
  assign new_n14119 = ~new_n13714 & new_n13724;
  assign new_n14120 = ~new_n13713 & ~new_n14119;
  assign new_n14121 = n4964 & n11350;
  assign new_n14122 = n5684 & n9846;
  assign new_n14123 = ~new_n14121 & ~new_n14122;
  assign new_n14124 = new_n14121 & new_n14122;
  assign new_n14125 = ~new_n14123 & ~new_n14124;
  assign new_n14126 = n4122 & n8940;
  assign new_n14127 = n469 & n3130;
  assign new_n14128 = n4382 & n12065;
  assign new_n14129 = ~new_n14127 & new_n14128;
  assign new_n14130 = new_n14127 & ~new_n14128;
  assign new_n14131 = ~new_n14129 & ~new_n14130;
  assign new_n14132 = ~new_n14126 & new_n14131;
  assign new_n14133 = new_n14126 & ~new_n14131;
  assign new_n14134 = ~new_n14132 & ~new_n14133;
  assign new_n14135 = ~new_n14125 & new_n14134;
  assign new_n14136 = new_n14125 & ~new_n14134;
  assign new_n14137 = ~new_n14135 & ~new_n14136;
  assign new_n14138 = new_n13814 & ~new_n13817;
  assign new_n14139 = ~new_n13818 & ~new_n14138;
  assign new_n14140 = n6333 & n11396;
  assign new_n14141 = n22 & n1912;
  assign new_n14142 = new_n14140 & ~new_n14141;
  assign new_n14143 = ~new_n14140 & new_n14141;
  assign new_n14144 = ~new_n14142 & ~new_n14143;
  assign new_n14145 = new_n14139 & new_n14144;
  assign new_n14146 = ~new_n14139 & ~new_n14144;
  assign new_n14147 = ~new_n14145 & ~new_n14146;
  assign new_n14148 = ~new_n14137 & new_n14147;
  assign new_n14149 = new_n14137 & ~new_n14147;
  assign new_n14150 = ~new_n14148 & ~new_n14149;
  assign new_n14151 = n411 & n4743;
  assign new_n14152 = n11488 & n11734;
  assign new_n14153 = ~n1982 & new_n14152;
  assign new_n14154 = n1982 & ~new_n14152;
  assign new_n14155 = ~new_n14153 & ~new_n14154;
  assign new_n14156 = new_n14151 & new_n14155;
  assign new_n14157 = ~new_n14151 & ~new_n14155;
  assign new_n14158 = ~new_n14156 & ~new_n14157;
  assign new_n14159 = n3085 & n12352;
  assign new_n14160 = n9353 & n12372;
  assign new_n14161 = ~new_n14159 & new_n14160;
  assign new_n14162 = new_n14159 & ~new_n14160;
  assign new_n14163 = ~new_n14161 & ~new_n14162;
  assign new_n14164 = n7411 & n10416;
  assign new_n14165 = n11030 & n12651;
  assign new_n14166 = ~new_n14164 & new_n14165;
  assign new_n14167 = new_n14164 & ~new_n14165;
  assign new_n14168 = ~new_n14166 & ~new_n14167;
  assign new_n14169 = ~new_n14163 & new_n14168;
  assign new_n14170 = new_n14163 & ~new_n14168;
  assign new_n14171 = ~new_n14169 & ~new_n14170;
  assign new_n14172 = new_n14158 & new_n14171;
  assign new_n14173 = ~new_n14158 & ~new_n14171;
  assign new_n14174 = ~new_n14172 & ~new_n14173;
  assign new_n14175 = new_n13700 & ~new_n13703;
  assign new_n14176 = ~new_n13704 & ~new_n14175;
  assign new_n14177 = new_n14174 & new_n14176;
  assign new_n14178 = ~new_n14174 & ~new_n14176;
  assign new_n14179 = ~new_n14177 & ~new_n14178;
  assign new_n14180 = ~new_n14150 & new_n14179;
  assign new_n14181 = new_n14150 & ~new_n14179;
  assign new_n14182 = ~new_n14180 & ~new_n14181;
  assign new_n14183 = new_n14120 & ~new_n14182;
  assign new_n14184 = ~new_n14120 & new_n14182;
  assign new_n14185 = ~new_n14183 & ~new_n14184;
  assign new_n14186 = ~new_n13616 & ~new_n13619;
  assign new_n14187 = ~new_n13615 & ~new_n14186;
  assign new_n14188 = ~new_n14185 & new_n14187;
  assign new_n14189 = new_n14185 & ~new_n14187;
  assign new_n14190 = ~new_n14188 & ~new_n14189;
  assign new_n14191 = ~new_n14118 & ~new_n14190;
  assign new_n14192 = new_n14118 & new_n14190;
  assign new_n14193 = ~new_n14191 & ~new_n14192;
  assign new_n14194 = ~new_n13594 & new_n13611;
  assign new_n14195 = ~new_n13593 & ~new_n14194;
  assign new_n14196 = ~new_n13826 & new_n13838;
  assign new_n14197 = ~new_n13825 & ~new_n14196;
  assign new_n14198 = n11180 & n11236;
  assign new_n14199 = n103 & n6826;
  assign new_n14200 = n9732 & n12284;
  assign new_n14201 = ~new_n14199 & new_n14200;
  assign new_n14202 = new_n14199 & ~new_n14200;
  assign new_n14203 = ~new_n14201 & ~new_n14202;
  assign new_n14204 = n761 & n10805;
  assign new_n14205 = n124 & n5758;
  assign new_n14206 = ~new_n14204 & ~new_n14205;
  assign new_n14207 = new_n14204 & new_n14205;
  assign new_n14208 = ~new_n14206 & ~new_n14207;
  assign new_n14209 = ~new_n14203 & new_n14208;
  assign new_n14210 = new_n14203 & ~new_n14208;
  assign new_n14211 = ~new_n14209 & ~new_n14210;
  assign new_n14212 = ~new_n14198 & new_n14211;
  assign new_n14213 = new_n14198 & ~new_n14211;
  assign new_n14214 = ~new_n14212 & ~new_n14213;
  assign new_n14215 = ~new_n14197 & new_n14214;
  assign new_n14216 = new_n14197 & ~new_n14214;
  assign new_n14217 = ~new_n14215 & ~new_n14216;
  assign new_n14218 = new_n14195 & new_n14217;
  assign new_n14219 = ~new_n14195 & ~new_n14217;
  assign new_n14220 = ~new_n14218 & ~new_n14219;
  assign new_n14221 = ~new_n13922 & ~new_n13926;
  assign new_n14222 = ~new_n13925 & ~new_n14221;
  assign new_n14223 = ~new_n13601 & ~new_n13605;
  assign new_n14224 = new_n14222 & new_n14223;
  assign new_n14225 = ~new_n14222 & ~new_n14223;
  assign new_n14226 = ~new_n14224 & ~new_n14225;
  assign new_n14227 = new_n13716 & ~new_n13719;
  assign new_n14228 = ~new_n13720 & ~new_n14227;
  assign new_n14229 = n9620 & n12263;
  assign new_n14230 = n353 & n12750;
  assign new_n14231 = ~new_n14229 & ~new_n14230;
  assign new_n14232 = new_n14229 & new_n14230;
  assign new_n14233 = ~new_n14231 & ~new_n14232;
  assign new_n14234 = n2737 & n10770;
  assign new_n14235 = n10522 & n12408;
  assign new_n14236 = new_n14234 & ~new_n14235;
  assign new_n14237 = ~new_n14234 & new_n14235;
  assign new_n14238 = ~new_n14236 & ~new_n14237;
  assign new_n14239 = ~new_n14233 & new_n14238;
  assign new_n14240 = new_n14233 & ~new_n14238;
  assign new_n14241 = ~new_n14239 & ~new_n14240;
  assign new_n14242 = ~new_n13831 & new_n14241;
  assign new_n14243 = new_n13831 & ~new_n14241;
  assign new_n14244 = ~new_n14242 & ~new_n14243;
  assign new_n14245 = new_n14228 & ~new_n14244;
  assign new_n14246 = ~new_n14228 & new_n14244;
  assign new_n14247 = ~new_n14245 & ~new_n14246;
  assign new_n14248 = new_n13938 & ~new_n13941;
  assign new_n14249 = ~new_n13942 & ~new_n14248;
  assign new_n14250 = new_n13584 & ~new_n13587;
  assign new_n14251 = ~new_n13588 & ~new_n14250;
  assign new_n14252 = n5320 & n9475;
  assign new_n14253 = n8228 & n12912;
  assign new_n14254 = ~new_n14252 & new_n14253;
  assign new_n14255 = new_n14252 & ~new_n14253;
  assign new_n14256 = ~new_n14254 & ~new_n14255;
  assign new_n14257 = new_n14251 & ~new_n14256;
  assign new_n14258 = ~new_n14251 & new_n14256;
  assign new_n14259 = ~new_n14257 & ~new_n14258;
  assign new_n14260 = n6149 & n10113;
  assign new_n14261 = n8820 & ~new_n14260;
  assign new_n14262 = ~n8820 & new_n14260;
  assign new_n14263 = ~new_n14261 & ~new_n14262;
  assign new_n14264 = n2482 & n5715;
  assign new_n14265 = n1757 & ~n7161;
  assign new_n14266 = ~new_n14264 & new_n14265;
  assign new_n14267 = new_n14264 & ~new_n14265;
  assign new_n14268 = ~new_n14266 & ~new_n14267;
  assign new_n14269 = ~new_n14263 & ~new_n14268;
  assign new_n14270 = new_n14263 & new_n14268;
  assign new_n14271 = ~new_n14269 & ~new_n14270;
  assign new_n14272 = new_n14259 & ~new_n14271;
  assign new_n14273 = ~new_n14259 & new_n14271;
  assign new_n14274 = ~new_n14272 & ~new_n14273;
  assign new_n14275 = ~new_n14249 & new_n14274;
  assign new_n14276 = new_n14249 & ~new_n14274;
  assign new_n14277 = ~new_n14275 & ~new_n14276;
  assign new_n14278 = new_n14247 & new_n14277;
  assign new_n14279 = ~new_n14247 & ~new_n14277;
  assign new_n14280 = ~new_n14278 & ~new_n14279;
  assign new_n14281 = new_n14226 & ~new_n14280;
  assign new_n14282 = ~new_n14226 & new_n14280;
  assign new_n14283 = ~new_n14281 & ~new_n14282;
  assign new_n14284 = ~new_n14220 & ~new_n14283;
  assign new_n14285 = new_n14220 & new_n14283;
  assign new_n14286 = ~new_n14284 & ~new_n14285;
  assign new_n14287 = ~new_n14193 & new_n14286;
  assign new_n14288 = new_n14193 & ~new_n14286;
  assign new_n14289 = ~new_n14287 & ~new_n14288;
  assign new_n14290 = ~new_n13811 & ~new_n13841;
  assign new_n14291 = ~new_n13812 & ~new_n14290;
  assign new_n14292 = new_n13831 & ~new_n13833;
  assign new_n14293 = ~new_n13834 & ~new_n14292;
  assign new_n14294 = ~new_n14291 & ~new_n14293;
  assign new_n14295 = new_n14291 & new_n14293;
  assign new_n14296 = ~new_n14294 & ~new_n14295;
  assign new_n14297 = new_n14289 & ~new_n14296;
  assign new_n14298 = ~new_n14289 & new_n14296;
  assign new_n14299 = ~new_n14297 & ~new_n14298;
  assign new_n14300 = ~new_n14116 & new_n14299;
  assign new_n14301 = new_n14116 & ~new_n14299;
  assign new_n14302 = ~new_n14300 & ~new_n14301;
  assign new_n14303 = new_n14002 & ~new_n14302;
  assign new_n14304 = ~new_n14002 & new_n14302;
  assign new_n14305 = ~new_n14303 & ~new_n14304;
  assign new_n14306 = ~new_n13624 & ~new_n13639;
  assign new_n14307 = new_n14305 & new_n14306;
  assign new_n14308 = ~new_n14305 & ~new_n14306;
  assign new_n14309 = ~new_n14307 & ~new_n14308;
  assign new_n14310 = new_n14114 & ~new_n14309;
  assign new_n14311 = ~new_n14114 & new_n14309;
  assign new_n14312 = ~new_n14310 & ~new_n14311;
  assign new_n14313 = ~new_n14060 & ~new_n14312;
  assign new_n14314 = new_n14060 & new_n14312;
  assign n11252 = new_n14313 | new_n14314;
  assign new_n14316 = ~new_n1965 & ~new_n1966;
  assign new_n14317 = new_n2000 & ~new_n14316;
  assign new_n14318 = ~new_n2000 & new_n14316;
  assign n11264 = ~new_n14317 & ~new_n14318;
  assign new_n14320 = ~new_n5533 & ~new_n5534;
  assign new_n14321 = new_n4109 & ~new_n14320;
  assign new_n14322 = ~new_n4109 & new_n14320;
  assign n11484 = ~new_n14321 & ~new_n14322;
  assign new_n14324 = ~new_n11508 & ~new_n11524;
  assign new_n14325 = ~new_n11293 & new_n11303;
  assign new_n14326 = ~new_n11292 & ~new_n14325;
  assign new_n14327 = ~new_n11311 & new_n14326;
  assign new_n14328 = new_n11311 & ~new_n14326;
  assign new_n14329 = ~new_n14327 & ~new_n14328;
  assign new_n14330 = ~new_n11395 & new_n11398;
  assign new_n14331 = ~new_n11394 & ~new_n14330;
  assign new_n14332 = ~n10657 & ~new_n11351;
  assign new_n14333 = new_n11353 & ~new_n14332;
  assign new_n14334 = ~new_n11345 & new_n11384;
  assign new_n14335 = new_n11345 & ~new_n11384;
  assign new_n14336 = ~new_n14334 & ~new_n14335;
  assign new_n14337 = new_n14333 & new_n14336;
  assign new_n14338 = ~new_n14333 & ~new_n14336;
  assign new_n14339 = ~new_n14337 & ~new_n14338;
  assign new_n14340 = new_n11391 & new_n14339;
  assign new_n14341 = ~new_n11391 & ~new_n14339;
  assign new_n14342 = ~new_n14340 & ~new_n14341;
  assign new_n14343 = new_n14331 & ~new_n14342;
  assign new_n14344 = ~new_n14331 & new_n14342;
  assign new_n14345 = ~new_n14343 & ~new_n14344;
  assign new_n14346 = ~new_n14329 & ~new_n14345;
  assign new_n14347 = new_n14329 & new_n14345;
  assign new_n14348 = ~new_n14346 & ~new_n14347;
  assign new_n14349 = ~new_n386 & new_n14348;
  assign new_n14350 = new_n386 & ~new_n14348;
  assign new_n14351 = ~new_n14349 & ~new_n14350;
  assign new_n14352 = new_n14324 & ~new_n14351;
  assign new_n14353 = ~new_n14324 & new_n14351;
  assign new_n14354 = ~new_n14352 & ~new_n14353;
  assign new_n14355 = new_n11279 & ~new_n11282;
  assign new_n14356 = ~new_n11283 & ~new_n14355;
  assign new_n14357 = ~new_n14354 & new_n14356;
  assign new_n14358 = new_n14354 & ~new_n14356;
  assign new_n14359 = ~new_n14357 & ~new_n14358;
  assign new_n14360 = ~new_n11621 & ~new_n11640;
  assign new_n14361 = ~new_n11620 & ~new_n14360;
  assign new_n14362 = n5031 & n6023;
  assign new_n14363 = n9 & n12579;
  assign new_n14364 = n2666 & n8466;
  assign new_n14365 = new_n14363 & ~new_n14364;
  assign new_n14366 = ~new_n14363 & new_n14364;
  assign new_n14367 = ~new_n14365 & ~new_n14366;
  assign new_n14368 = n9591 & n11061;
  assign new_n14369 = n2592 & n11222;
  assign new_n14370 = new_n14368 & ~new_n14369;
  assign new_n14371 = ~new_n14368 & new_n14369;
  assign new_n14372 = ~new_n14370 & ~new_n14371;
  assign new_n14373 = ~new_n14367 & ~new_n14372;
  assign new_n14374 = new_n14367 & new_n14372;
  assign new_n14375 = ~new_n14373 & ~new_n14374;
  assign new_n14376 = ~new_n14362 & new_n14375;
  assign new_n14377 = new_n14362 & ~new_n14375;
  assign new_n14378 = ~new_n14376 & ~new_n14377;
  assign new_n14379 = new_n11590 & ~new_n14378;
  assign new_n14380 = ~new_n11590 & new_n14378;
  assign new_n14381 = ~new_n14379 & ~new_n14380;
  assign new_n14382 = ~new_n14361 & new_n14381;
  assign new_n14383 = new_n14361 & ~new_n14381;
  assign new_n14384 = ~new_n14382 & ~new_n14383;
  assign new_n14385 = new_n14359 & ~new_n14384;
  assign new_n14386 = ~new_n14359 & new_n14384;
  assign new_n14387 = ~new_n14385 & ~new_n14386;
  assign new_n14388 = ~new_n11614 & ~new_n11617;
  assign new_n14389 = ~new_n11402 & ~new_n11408;
  assign new_n14390 = ~new_n11405 & new_n14389;
  assign new_n14391 = new_n14388 & ~new_n14390;
  assign new_n14392 = ~new_n14388 & new_n14390;
  assign new_n14393 = ~new_n14391 & ~new_n14392;
  assign new_n14394 = new_n11469 & ~new_n11472;
  assign new_n14395 = ~new_n11473 & ~new_n14394;
  assign new_n14396 = new_n11485 & ~new_n11488_1;
  assign new_n14397 = ~new_n11489 & ~new_n14396;
  assign new_n14398 = ~new_n14395 & new_n14397;
  assign new_n14399 = new_n14395 & ~new_n14397;
  assign new_n14400 = ~new_n14398 & ~new_n14399;
  assign new_n14401 = n510 & n4998;
  assign new_n14402 = ~new_n11482 & new_n11493;
  assign new_n14403 = ~new_n11483 & ~new_n14402;
  assign new_n14404 = n2341 & n12592;
  assign new_n14405 = new_n11501 & new_n14404;
  assign new_n14406 = ~new_n11501 & ~new_n14404;
  assign new_n14407 = ~new_n14405 & ~new_n14406;
  assign new_n14408 = new_n14403 & ~new_n14407;
  assign new_n14409 = ~new_n14403 & new_n14407;
  assign new_n14410 = ~new_n14408 & ~new_n14409;
  assign new_n14411 = new_n14401 & new_n14410;
  assign new_n14412 = ~new_n14401 & ~new_n14410;
  assign new_n14413 = ~new_n14411 & ~new_n14412;
  assign new_n14414 = new_n14400 & ~new_n14413;
  assign new_n14415 = ~new_n14400 & new_n14413;
  assign new_n14416 = ~new_n14414 & ~new_n14415;
  assign new_n14417 = ~new_n11466 & new_n11503;
  assign new_n14418 = ~new_n11467 & ~new_n14417;
  assign new_n14419 = n951 & n5189;
  assign new_n14420 = n767 & n2295;
  assign new_n14421 = ~new_n14419 & ~new_n14420;
  assign new_n14422 = new_n14419 & new_n14420;
  assign new_n14423 = ~new_n14421 & ~new_n14422;
  assign new_n14424 = n401 & n8716;
  assign new_n14425 = n3178 & n12693;
  assign new_n14426 = ~new_n14424 & new_n14425;
  assign new_n14427 = new_n14424 & ~new_n14425;
  assign new_n14428 = ~new_n14426 & ~new_n14427;
  assign new_n14429 = ~new_n14423 & new_n14428;
  assign new_n14430 = new_n14423 & ~new_n14428;
  assign new_n14431 = ~new_n14429 & ~new_n14430;
  assign new_n14432 = n834 & n4419;
  assign new_n14433 = n11537 & n13060;
  assign new_n14434 = n1650 & n10168;
  assign new_n14435 = new_n14433 & ~new_n14434;
  assign new_n14436 = ~new_n14433 & new_n14434;
  assign new_n14437 = ~new_n14435 & ~new_n14436;
  assign new_n14438 = new_n14432 & new_n14437;
  assign new_n14439 = ~new_n14432 & ~new_n14437;
  assign new_n14440 = ~new_n14438 & ~new_n14439;
  assign new_n14441 = new_n14431 & new_n14440;
  assign new_n14442 = ~new_n14431 & ~new_n14440;
  assign new_n14443 = ~new_n14441 & ~new_n14442;
  assign new_n14444 = new_n11612 & ~new_n14443;
  assign new_n14445 = ~new_n11612 & new_n14443;
  assign new_n14446 = ~new_n14444 & ~new_n14445;
  assign new_n14447 = new_n14418 & new_n14446;
  assign new_n14448 = ~new_n14418 & ~new_n14446;
  assign new_n14449 = ~new_n14447 & ~new_n14448;
  assign new_n14450 = n389 & n9216;
  assign new_n14451 = n854 & n4452;
  assign new_n14452 = ~new_n14450 & ~new_n14451;
  assign new_n14453 = new_n14450 & new_n14451;
  assign new_n14454 = ~new_n14452 & ~new_n14453;
  assign new_n14455 = new_n14449 & ~new_n14454;
  assign new_n14456 = ~new_n14449 & new_n14454;
  assign new_n14457 = ~new_n14455 & ~new_n14456;
  assign new_n14458 = ~new_n14416 & new_n14457;
  assign new_n14459 = new_n14416 & ~new_n14457;
  assign new_n14460 = ~new_n14458 & ~new_n14459;
  assign new_n14461 = new_n14393 & ~new_n14460;
  assign new_n14462 = ~new_n14393 & new_n14460;
  assign new_n14463 = ~new_n14461 & ~new_n14462;
  assign new_n14464 = ~new_n11645 & ~new_n11670;
  assign new_n14465 = ~new_n11644 & ~new_n14464;
  assign new_n14466 = new_n14463 & new_n14465;
  assign new_n14467 = ~new_n14463 & ~new_n14465;
  assign new_n14468 = ~new_n14466 & ~new_n14467;
  assign new_n14469 = new_n14387 & new_n14468;
  assign new_n14470 = ~new_n14387 & ~new_n14468;
  assign new_n14471 = ~new_n14469 & ~new_n14470;
  assign new_n14472 = ~new_n11318 & ~new_n11334;
  assign new_n14473 = ~new_n11276 & new_n11313;
  assign new_n14474 = ~new_n11277 & ~new_n14473;
  assign new_n14475 = new_n11592 & ~new_n11595;
  assign new_n14476 = ~new_n11596 & ~new_n14475;
  assign new_n14477 = ~new_n11591 & ~new_n11603;
  assign new_n14478 = ~new_n11604 & ~new_n14477;
  assign new_n14479 = ~new_n14476 & ~new_n14478;
  assign new_n14480 = new_n14476 & new_n14478;
  assign new_n14481 = ~new_n14479 & ~new_n14480;
  assign new_n14482 = n6655 & n7715;
  assign new_n14483 = n2458 & n9528;
  assign new_n14484 = new_n14482 & ~new_n14483;
  assign new_n14485 = ~new_n14482 & new_n14483;
  assign new_n14486 = ~new_n14484 & ~new_n14485;
  assign new_n14487 = n6668 & n11891;
  assign new_n14488 = n8230 & n9669;
  assign new_n14489 = ~new_n14487 & ~new_n14488;
  assign new_n14490 = new_n14487 & new_n14488;
  assign new_n14491 = ~new_n14489 & ~new_n14490;
  assign new_n14492 = n7529 & n8522;
  assign new_n14493 = n7812 & n9531;
  assign new_n14494 = new_n14492 & new_n14493;
  assign new_n14495 = ~new_n14492 & ~new_n14493;
  assign new_n14496 = ~new_n14494 & ~new_n14495;
  assign new_n14497 = new_n14491 & ~new_n14496;
  assign new_n14498 = ~new_n14491 & new_n14496;
  assign new_n14499 = ~new_n14497 & ~new_n14498;
  assign new_n14500 = ~new_n14486 & new_n14499;
  assign new_n14501 = new_n14486 & ~new_n14499;
  assign new_n14502 = ~new_n14500 & ~new_n14501;
  assign new_n14503 = ~new_n11295 & ~new_n11299;
  assign new_n14504 = ~new_n11298 & ~new_n14503;
  assign new_n14505 = n5427 & n7772;
  assign new_n14506 = new_n14504 & new_n14505;
  assign new_n14507 = ~new_n14504 & ~new_n14505;
  assign new_n14508 = ~new_n14506 & ~new_n14507;
  assign new_n14509 = new_n14502 & new_n14508;
  assign new_n14510 = ~new_n14502 & ~new_n14508;
  assign new_n14511 = ~new_n14509 & ~new_n14510;
  assign new_n14512 = ~new_n14481 & new_n14511;
  assign new_n14513 = new_n14481 & ~new_n14511;
  assign new_n14514 = ~new_n14512 & ~new_n14513;
  assign new_n14515 = new_n14474 & new_n14514;
  assign new_n14516 = ~new_n14474 & ~new_n14514;
  assign new_n14517 = ~new_n14515 & ~new_n14516;
  assign new_n14518 = n8290 & n8768;
  assign new_n14519 = new_n11580 & ~new_n11583;
  assign new_n14520 = ~new_n11584 & ~new_n14519;
  assign new_n14521 = ~new_n14518 & ~new_n14520;
  assign new_n14522 = new_n14518 & new_n14520;
  assign new_n14523 = ~new_n14521 & ~new_n14522;
  assign new_n14524 = ~new_n14517 & new_n14523;
  assign new_n14525 = new_n14517 & ~new_n14523;
  assign new_n14526 = ~new_n14524 & ~new_n14525;
  assign new_n14527 = new_n14472 & new_n14526;
  assign new_n14528 = ~new_n14472 & ~new_n14526;
  assign new_n14529 = ~new_n14527 & ~new_n14528;
  assign new_n14530 = ~new_n11674 & ~new_n11698;
  assign new_n14531 = ~new_n11675 & ~new_n14530;
  assign new_n14532 = ~new_n14529 & new_n14531;
  assign new_n14533 = new_n14529 & ~new_n14531;
  assign new_n14534 = ~new_n14532 & ~new_n14533;
  assign new_n14535 = ~new_n14471 & ~new_n14534;
  assign new_n14536 = new_n14471 & new_n14534;
  assign n11667 = new_n14535 | new_n14536;
  assign new_n14538 = ~new_n4895 & ~new_n4896;
  assign new_n14539 = ~new_n4900 & new_n14538;
  assign new_n14540 = new_n4900 & ~new_n14538;
  assign n11732 = ~new_n14539 & ~new_n14540;
  assign new_n14542 = ~new_n13269 & ~new_n13270;
  assign new_n14543 = new_n13274 & new_n14542;
  assign new_n14544 = ~new_n13274 & ~new_n14542;
  assign n11778 = ~new_n14543 & ~new_n14544;
  assign new_n14546 = ~new_n1985 & ~new_n1987;
  assign n11792 = ~new_n1988 & ~new_n14546;
  assign new_n14548 = ~new_n14048 & ~new_n14049;
  assign new_n14549 = new_n14053 & ~new_n14548;
  assign new_n14550 = ~new_n14053 & new_n14548;
  assign n11879 = new_n14549 | new_n14550;
  assign new_n14552 = ~new_n2617 & ~new_n2618;
  assign new_n14553 = ~new_n2652 & ~new_n14552;
  assign new_n14554 = new_n2652 & new_n14552;
  assign n11882 = new_n14553 | new_n14554;
  assign new_n14556 = new_n10458 & ~new_n10462;
  assign new_n14557 = new_n10467 & ~new_n14556;
  assign new_n14558 = new_n10462 & ~new_n10466;
  assign n11895 = ~new_n14557 & ~new_n14558;
  assign new_n14560 = ~new_n12451 & ~new_n12452;
  assign new_n14561 = new_n12464 & ~new_n14560;
  assign new_n14562 = ~new_n12451 & new_n12465;
  assign n12059 = new_n14561 | new_n14562;
  assign new_n14564 = ~new_n14042 & ~new_n14043;
  assign new_n14565 = new_n14045 & new_n14564;
  assign new_n14566 = ~new_n14045 & ~new_n14564;
  assign n12067 = new_n14565 | new_n14566;
  assign new_n14568 = ~new_n5287 & ~new_n5288;
  assign new_n14569 = ~new_n5292 & new_n14568;
  assign new_n14570 = new_n5292 & ~new_n14568;
  assign n12187 = new_n14569 | new_n14570;
  assign new_n14572 = ~new_n9582 & ~new_n9583;
  assign new_n14573 = ~new_n9584 & ~new_n14572;
  assign new_n14574 = new_n9584 & new_n14572;
  assign n12334 = new_n14573 | new_n14574;
  assign new_n14576 = ~n7161 & n7772;
  assign new_n14577 = ~new_n12521 & ~new_n12525;
  assign new_n14578 = ~new_n12522 & ~new_n14577;
  assign new_n14579 = n7411 & n7529;
  assign new_n14580 = n7715 & n12651;
  assign new_n14581 = ~new_n14579 & ~new_n14580;
  assign new_n14582 = new_n14579 & new_n14580;
  assign new_n14583 = ~new_n14581 & ~new_n14582;
  assign new_n14584 = n2458 & n11734;
  assign new_n14585 = n6668 & n8230;
  assign new_n14586 = ~n6668 & ~n8230;
  assign new_n14587 = ~new_n14585 & ~new_n14586;
  assign new_n14588 = new_n14584 & new_n14587;
  assign new_n14589 = ~new_n14584 & ~new_n14587;
  assign new_n14590 = ~new_n12509 & ~new_n14589;
  assign new_n14591 = ~new_n14588 & new_n14590;
  assign new_n14592 = ~new_n14588 & ~new_n14589;
  assign new_n14593 = new_n12509 & ~new_n14592;
  assign new_n14594 = ~new_n14591 & ~new_n14593;
  assign new_n14595 = ~new_n14583 & ~new_n14594;
  assign new_n14596 = new_n14583 & new_n14594;
  assign new_n14597 = ~new_n14595 & ~new_n14596;
  assign new_n14598 = ~new_n12513 & ~new_n12515_1;
  assign new_n14599 = ~new_n12516 & ~new_n14598;
  assign new_n14600 = ~new_n14597 & new_n14599;
  assign new_n14601 = new_n14597 & ~new_n14599;
  assign new_n14602 = ~new_n14600 & ~new_n14601;
  assign new_n14603 = ~new_n14578 & new_n14602;
  assign new_n14604 = new_n14578 & ~new_n14602;
  assign new_n14605 = ~new_n14603 & ~new_n14604;
  assign new_n14606 = new_n14576 & new_n14605;
  assign new_n14607 = ~new_n14576 & ~new_n14605;
  assign new_n14608 = ~new_n14606 & ~new_n14607;
  assign new_n14609 = new_n12529 & new_n14608;
  assign new_n14610 = ~new_n14606 & ~new_n14609;
  assign new_n14611 = ~new_n14588 & ~new_n14590;
  assign new_n14612 = n7411 & n7715;
  assign new_n14613 = ~n7161 & n7529;
  assign new_n14614 = n6149 & n7772;
  assign new_n14615 = ~new_n14613 & ~new_n14614;
  assign new_n14616 = new_n14613 & new_n14614;
  assign new_n14617 = ~new_n14615 & ~new_n14616;
  assign new_n14618 = new_n14612 & ~new_n14617;
  assign new_n14619 = ~new_n14612 & new_n14617;
  assign new_n14620 = ~new_n14618 & ~new_n14619;
  assign new_n14621 = ~new_n14611 & ~new_n14620;
  assign new_n14622 = new_n14611 & new_n14620;
  assign new_n14623 = ~new_n14621 & ~new_n14622;
  assign new_n14624 = n2458 & n12651;
  assign new_n14625 = new_n14585 & new_n14624;
  assign new_n14626 = ~new_n14585 & ~new_n14624;
  assign new_n14627 = ~new_n14625 & ~new_n14626;
  assign new_n14628 = n8230 & n11734;
  assign new_n14629 = ~n6668 & ~new_n14628;
  assign new_n14630 = ~n7812 & new_n14629;
  assign new_n14631 = n11734 & new_n14585;
  assign new_n14632 = ~n7812 & ~new_n14631;
  assign new_n14633 = ~new_n14629 & ~new_n14632;
  assign new_n14634 = n7812 & new_n14631;
  assign new_n14635 = new_n14633 & ~new_n14634;
  assign new_n14636 = ~new_n14630 & ~new_n14635;
  assign new_n14637 = ~new_n14627 & ~new_n14636;
  assign new_n14638 = new_n14627 & new_n14636;
  assign new_n14639 = ~new_n14637 & ~new_n14638;
  assign new_n14640 = new_n14623 & ~new_n14639;
  assign new_n14641 = ~new_n14623 & new_n14639;
  assign new_n14642 = ~new_n14640 & ~new_n14641;
  assign new_n14643 = new_n14582 & ~new_n14642;
  assign new_n14644 = ~new_n14582 & new_n14642;
  assign new_n14645 = ~new_n14643 & ~new_n14644;
  assign new_n14646 = ~new_n14595 & ~new_n14599;
  assign new_n14647 = ~new_n14596 & ~new_n14646;
  assign new_n14648 = ~new_n14645 & ~new_n14647;
  assign new_n14649 = new_n14645 & new_n14647;
  assign new_n14650 = ~new_n14648 & ~new_n14649;
  assign new_n14651 = new_n14603 & ~new_n14650;
  assign new_n14652 = ~new_n14603 & new_n14650;
  assign new_n14653 = ~new_n14651 & ~new_n14652;
  assign new_n14654 = ~new_n14610 & new_n14653;
  assign new_n14655 = new_n14610 & ~new_n14653;
  assign new_n14656 = ~new_n14654 & ~new_n14655;
  assign new_n14657 = ~new_n12731 & new_n12734;
  assign new_n14658 = ~new_n12730 & ~new_n14657;
  assign new_n14659 = n469 & n12348;
  assign new_n14660 = n2068 & n12284;
  assign new_n14661 = ~new_n14659 & ~new_n14660;
  assign new_n14662 = new_n14659 & new_n14660;
  assign new_n14663 = ~new_n14661 & ~new_n14662;
  assign new_n14664 = n6826 & n11324;
  assign new_n14665 = n8183 & n9475;
  assign new_n14666 = n411 & n10142;
  assign new_n14667 = ~new_n14665 & ~new_n14666;
  assign new_n14668 = new_n14665 & new_n14666;
  assign new_n14669 = ~new_n14667 & ~new_n14668;
  assign new_n14670 = new_n14664 & new_n14669;
  assign new_n14671 = ~new_n14664 & ~new_n14669;
  assign new_n14672 = ~new_n14670 & ~new_n14671;
  assign new_n14673 = new_n12718 & ~new_n12721;
  assign new_n14674 = ~new_n12722 & ~new_n14673;
  assign new_n14675 = ~new_n14672 & new_n14674;
  assign new_n14676 = new_n14672 & ~new_n14674;
  assign new_n14677 = ~new_n14675 & ~new_n14676;
  assign new_n14678 = ~new_n14663 & ~new_n14677;
  assign new_n14679 = new_n14663 & new_n14677;
  assign new_n14680 = ~new_n14678 & ~new_n14679;
  assign new_n14681 = ~new_n12715 & ~new_n12726;
  assign new_n14682 = ~new_n12716 & ~new_n14681;
  assign new_n14683 = ~new_n14680 & ~new_n14682;
  assign new_n14684 = new_n14680 & new_n14682;
  assign new_n14685 = ~new_n14683 & ~new_n14684;
  assign new_n14686 = new_n14658 & ~new_n14685;
  assign new_n14687 = ~new_n14678 & ~new_n14682;
  assign new_n14688 = ~new_n14662 & ~new_n14687;
  assign new_n14689 = ~new_n14679 & new_n14688;
  assign new_n14690 = new_n14662 & new_n14687;
  assign new_n14691 = ~new_n14689 & ~new_n14690;
  assign new_n14692 = n9216 & n11180;
  assign new_n14693 = n469 & n2068;
  assign new_n14694 = n12065 & n12348;
  assign new_n14695 = ~new_n14693 & ~new_n14694;
  assign new_n14696 = new_n14693 & new_n14694;
  assign new_n14697 = ~new_n14695 & ~new_n14696;
  assign new_n14698 = new_n14692 & ~new_n14697;
  assign new_n14699 = ~new_n14692 & new_n14697;
  assign new_n14700 = ~new_n14698 & ~new_n14699;
  assign new_n14701 = ~new_n14670 & new_n14674;
  assign new_n14702 = ~new_n14671 & ~new_n14701;
  assign new_n14703 = new_n14700 & ~new_n14702;
  assign new_n14704 = n11324 & n12284;
  assign new_n14705 = ~new_n14668 & ~new_n14704;
  assign new_n14706 = new_n14668 & new_n14704;
  assign new_n14707 = ~new_n14705 & ~new_n14706;
  assign new_n14708 = n6826 & n8183;
  assign new_n14709 = n9475 & n10142;
  assign new_n14710 = n411 & n10657;
  assign new_n14711 = ~new_n14709 & ~new_n14710;
  assign new_n14712 = new_n14709 & new_n14710;
  assign new_n14713 = ~new_n14711 & ~new_n14712;
  assign new_n14714 = new_n14708 & ~new_n14713;
  assign new_n14715 = ~new_n14708 & new_n14713;
  assign new_n14716 = ~new_n14714 & ~new_n14715;
  assign new_n14717 = new_n14707 & new_n14716;
  assign new_n14718 = ~new_n14707 & ~new_n14716;
  assign new_n14719 = ~new_n14717 & ~new_n14718;
  assign new_n14720 = new_n14703 & new_n14719;
  assign new_n14721 = ~new_n14700 & new_n14702;
  assign new_n14722 = new_n14719 & ~new_n14721;
  assign new_n14723 = ~new_n14703 & ~new_n14722;
  assign new_n14724 = ~new_n14720 & ~new_n14723;
  assign new_n14725 = ~new_n14719 & new_n14721;
  assign new_n14726 = ~new_n14724 & ~new_n14725;
  assign new_n14727 = ~new_n14691 & ~new_n14726;
  assign new_n14728 = new_n14691 & new_n14726;
  assign new_n14729 = ~new_n14727 & ~new_n14728;
  assign new_n14730 = ~new_n14686 & new_n14729;
  assign new_n14731 = new_n14686 & ~new_n14729;
  assign new_n14732 = ~new_n14730 & ~new_n14731;
  assign new_n14733 = n9216 & n12065;
  assign new_n14734 = ~new_n14658 & new_n14685;
  assign new_n14735 = ~new_n14686 & ~new_n14734;
  assign new_n14736 = new_n14733 & new_n14735;
  assign new_n14737 = ~new_n14733 & ~new_n14735;
  assign new_n14738 = ~new_n14736 & ~new_n14737;
  assign new_n14739 = new_n12739 & new_n14738;
  assign new_n14740 = ~new_n14736 & ~new_n14739;
  assign new_n14741 = ~new_n14732 & new_n14740;
  assign new_n14742 = new_n14732 & ~new_n14740;
  assign new_n14743 = ~new_n14741 & ~new_n14742;
  assign new_n14744 = ~new_n12761 & new_n12764;
  assign new_n14745 = ~new_n12760 & ~new_n14744;
  assign new_n14746 = n5031 & n12408;
  assign new_n14747 = n9 & n2737;
  assign new_n14748 = ~new_n14746 & ~new_n14747;
  assign new_n14749 = new_n14746 & new_n14747;
  assign new_n14750 = ~new_n14748 & ~new_n14749;
  assign new_n14751 = n772 & n2592;
  assign new_n14752 = n2590 & n5536;
  assign new_n14753 = n8506 & n11061;
  assign new_n14754 = ~new_n14752 & ~new_n14753;
  assign new_n14755 = new_n14752 & new_n14753;
  assign new_n14756 = ~new_n14754 & ~new_n14755;
  assign new_n14757 = new_n14751 & new_n14756;
  assign new_n14758 = ~new_n14751 & ~new_n14756;
  assign new_n14759 = ~new_n14757 & ~new_n14758;
  assign new_n14760 = new_n12748 & ~new_n12751;
  assign new_n14761 = ~new_n12752 & ~new_n14760;
  assign new_n14762 = ~new_n14759 & new_n14761;
  assign new_n14763 = new_n14759 & ~new_n14761;
  assign new_n14764 = ~new_n14762 & ~new_n14763;
  assign new_n14765 = ~new_n14750 & ~new_n14764;
  assign new_n14766 = new_n14750 & new_n14764;
  assign new_n14767 = ~new_n14765 & ~new_n14766;
  assign new_n14768 = ~new_n12745 & ~new_n12756;
  assign new_n14769 = ~new_n12746 & ~new_n14768;
  assign new_n14770 = ~new_n14767 & ~new_n14769;
  assign new_n14771 = new_n14767 & new_n14769;
  assign new_n14772 = ~new_n14770 & ~new_n14771;
  assign new_n14773 = new_n14745 & ~new_n14772;
  assign new_n14774 = ~new_n14765 & ~new_n14769;
  assign new_n14775 = ~new_n14749 & ~new_n14774;
  assign new_n14776 = ~new_n14766 & new_n14775;
  assign new_n14777 = new_n14749 & new_n14774;
  assign new_n14778 = ~new_n14776 & ~new_n14777;
  assign new_n14779 = n8466 & n11350;
  assign new_n14780 = n9 & n12408;
  assign new_n14781 = n5031 & n9846;
  assign new_n14782 = ~new_n14780 & ~new_n14781;
  assign new_n14783 = new_n14780 & new_n14781;
  assign new_n14784 = ~new_n14782 & ~new_n14783;
  assign new_n14785 = new_n14779 & ~new_n14784;
  assign new_n14786 = ~new_n14779 & new_n14784;
  assign new_n14787 = ~new_n14785 & ~new_n14786;
  assign new_n14788 = ~new_n14757 & new_n14761;
  assign new_n14789 = ~new_n14758 & ~new_n14788;
  assign new_n14790 = new_n14787 & ~new_n14789;
  assign new_n14791 = n2592 & n2737;
  assign new_n14792 = new_n14755 & new_n14791;
  assign new_n14793 = ~new_n14755 & ~new_n14791;
  assign new_n14794 = ~new_n14792 & ~new_n14793;
  assign new_n14795 = n772 & n2590;
  assign new_n14796 = n5536 & n11061;
  assign new_n14797 = n8506 & n8768;
  assign new_n14798 = ~new_n14796 & ~new_n14797;
  assign new_n14799 = new_n14796 & new_n14797;
  assign new_n14800 = ~new_n14798 & ~new_n14799;
  assign new_n14801 = new_n14795 & ~new_n14800;
  assign new_n14802 = ~new_n14795 & new_n14800;
  assign new_n14803 = ~new_n14801 & ~new_n14802;
  assign new_n14804 = new_n14794 & new_n14803;
  assign new_n14805 = ~new_n14794 & ~new_n14803;
  assign new_n14806 = ~new_n14804 & ~new_n14805;
  assign new_n14807 = new_n14790 & new_n14806;
  assign new_n14808 = ~new_n14787 & new_n14789;
  assign new_n14809 = new_n14806 & ~new_n14808;
  assign new_n14810 = ~new_n14790 & ~new_n14809;
  assign new_n14811 = ~new_n14807 & ~new_n14810;
  assign new_n14812 = ~new_n14806 & new_n14808;
  assign new_n14813 = ~new_n14811 & ~new_n14812;
  assign new_n14814 = ~new_n14778 & new_n14813;
  assign new_n14815 = new_n14778 & ~new_n14813;
  assign new_n14816 = ~new_n14814 & ~new_n14815;
  assign new_n14817 = ~new_n14773 & ~new_n14816;
  assign new_n14818 = new_n14773 & new_n14816;
  assign new_n14819 = ~new_n14817 & ~new_n14818;
  assign new_n14820 = n8466 & n9846;
  assign new_n14821 = ~new_n14745 & new_n14772;
  assign new_n14822 = ~new_n14773 & ~new_n14821;
  assign new_n14823 = new_n14820 & new_n14822;
  assign new_n14824 = ~new_n14820 & ~new_n14822;
  assign new_n14825 = ~new_n14823 & ~new_n14824;
  assign new_n14826 = new_n12769 & new_n14825;
  assign new_n14827 = ~new_n14823 & ~new_n14826;
  assign new_n14828 = ~new_n14819 & new_n14827;
  assign new_n14829 = new_n14819 & ~new_n14827;
  assign new_n14830 = ~new_n14828 & ~new_n14829;
  assign new_n14831 = ~new_n12791 & new_n12794;
  assign new_n14832 = ~new_n12790 & ~new_n14831;
  assign new_n14833 = n353 & n12592;
  assign new_n14834 = n10168 & n12263;
  assign new_n14835 = ~new_n14833 & ~new_n14834;
  assign new_n14836 = new_n14833 & new_n14834;
  assign new_n14837 = ~new_n14835 & ~new_n14836;
  assign new_n14838 = n767 & n10805;
  assign new_n14839 = n124 & n11537;
  assign new_n14840 = n951 & n3085;
  assign new_n14841 = ~new_n14839 & ~new_n14840;
  assign new_n14842 = new_n14839 & new_n14840;
  assign new_n14843 = ~new_n14841 & ~new_n14842;
  assign new_n14844 = new_n14838 & new_n14843;
  assign new_n14845 = ~new_n14838 & ~new_n14843;
  assign new_n14846 = ~new_n14844 & ~new_n14845;
  assign new_n14847 = new_n12778 & ~new_n12781;
  assign new_n14848 = ~new_n12782 & ~new_n14847;
  assign new_n14849 = ~new_n14846 & new_n14848;
  assign new_n14850 = new_n14846 & ~new_n14848;
  assign new_n14851 = ~new_n14849 & ~new_n14850;
  assign new_n14852 = ~new_n14837 & ~new_n14851;
  assign new_n14853 = new_n14837 & new_n14851;
  assign new_n14854 = ~new_n14852 & ~new_n14853;
  assign new_n14855 = ~new_n12775 & ~new_n12786;
  assign new_n14856 = ~new_n12776 & ~new_n14855;
  assign new_n14857 = ~new_n14854 & ~new_n14856;
  assign new_n14858 = new_n14854 & new_n14856;
  assign new_n14859 = ~new_n14857 & ~new_n14858;
  assign new_n14860 = new_n14832 & ~new_n14859;
  assign new_n14861 = ~new_n14852 & ~new_n14856;
  assign new_n14862 = ~new_n14836 & ~new_n14861;
  assign new_n14863 = ~new_n14853 & new_n14862;
  assign new_n14864 = new_n14836 & new_n14861;
  assign new_n14865 = ~new_n14863 & ~new_n14864;
  assign new_n14866 = n3178 & n11396;
  assign new_n14867 = n353 & n10168;
  assign new_n14868 = n22 & n12592;
  assign new_n14869 = ~new_n14867 & ~new_n14868;
  assign new_n14870 = new_n14867 & new_n14868;
  assign new_n14871 = ~new_n14869 & ~new_n14870;
  assign new_n14872 = new_n14866 & ~new_n14871;
  assign new_n14873 = ~new_n14866 & new_n14871;
  assign new_n14874 = ~new_n14872 & ~new_n14873;
  assign new_n14875 = ~new_n14844 & new_n14848;
  assign new_n14876 = ~new_n14845 & ~new_n14875;
  assign new_n14877 = new_n14874 & ~new_n14876;
  assign new_n14878 = n767 & n12263;
  assign new_n14879 = new_n14842 & new_n14878;
  assign new_n14880 = ~new_n14842 & ~new_n14878;
  assign new_n14881 = ~new_n14879 & ~new_n14880;
  assign new_n14882 = n10805 & n11537;
  assign new_n14883 = n124 & n951;
  assign new_n14884 = n401 & n3085;
  assign new_n14885 = ~new_n14883 & ~new_n14884;
  assign new_n14886 = new_n14883 & new_n14884;
  assign new_n14887 = ~new_n14885 & ~new_n14886;
  assign new_n14888 = new_n14882 & ~new_n14887;
  assign new_n14889 = ~new_n14882 & new_n14887;
  assign new_n14890 = ~new_n14888 & ~new_n14889;
  assign new_n14891 = new_n14881 & new_n14890;
  assign new_n14892 = ~new_n14881 & ~new_n14890;
  assign new_n14893 = ~new_n14891 & ~new_n14892;
  assign new_n14894 = new_n14877 & new_n14893;
  assign new_n14895 = ~new_n14874 & new_n14876;
  assign new_n14896 = new_n14893 & ~new_n14895;
  assign new_n14897 = ~new_n14877 & ~new_n14896;
  assign new_n14898 = ~new_n14894 & ~new_n14897;
  assign new_n14899 = ~new_n14893 & new_n14895;
  assign new_n14900 = ~new_n14898 & ~new_n14899;
  assign new_n14901 = ~new_n14865 & new_n14900;
  assign new_n14902 = new_n14865 & ~new_n14900;
  assign new_n14903 = ~new_n14901 & ~new_n14902;
  assign new_n14904 = ~new_n14860 & ~new_n14903;
  assign new_n14905 = new_n14860 & new_n14903;
  assign new_n14906 = ~new_n14904 & ~new_n14905;
  assign new_n14907 = n22 & n3178;
  assign new_n14908 = ~new_n14832 & new_n14859;
  assign new_n14909 = ~new_n14860 & ~new_n14908;
  assign new_n14910 = new_n14907 & new_n14909;
  assign new_n14911 = ~new_n14907 & ~new_n14909;
  assign new_n14912 = ~new_n14910 & ~new_n14911;
  assign new_n14913 = new_n12799 & new_n14912;
  assign new_n14914 = ~new_n14910 & ~new_n14913;
  assign new_n14915 = ~new_n14906 & new_n14914;
  assign new_n14916 = new_n14906 & ~new_n14914;
  assign new_n14917 = ~new_n14915 & ~new_n14916;
  assign new_n14918 = new_n14830 & new_n14917;
  assign new_n14919 = ~new_n14830 & ~new_n14917;
  assign new_n14920 = ~new_n14918 & ~new_n14919;
  assign new_n14921 = ~new_n12799 & ~new_n14912;
  assign new_n14922 = ~new_n14913 & ~new_n14921;
  assign new_n14923 = ~new_n12802 & ~new_n12805;
  assign new_n14924 = ~new_n12801 & ~new_n14923;
  assign new_n14925 = ~new_n14922 & new_n14924;
  assign new_n14926 = new_n14922 & ~new_n14924;
  assign new_n14927 = ~new_n12769 & ~new_n14825;
  assign new_n14928 = ~new_n14826 & ~new_n14927;
  assign new_n14929 = ~new_n14926 & ~new_n14928;
  assign new_n14930 = ~new_n14925 & ~new_n14929;
  assign new_n14931 = new_n14920 & ~new_n14930;
  assign new_n14932 = ~new_n14920 & new_n14930;
  assign new_n14933 = ~new_n14931 & ~new_n14932;
  assign new_n14934 = new_n14743 & ~new_n14933;
  assign new_n14935 = ~new_n14743 & new_n14933;
  assign new_n14936 = ~new_n14934 & ~new_n14935;
  assign new_n14937 = ~new_n12739 & ~new_n14738;
  assign new_n14938 = ~new_n14739 & ~new_n14937;
  assign new_n14939 = ~new_n14925 & ~new_n14926;
  assign new_n14940 = ~new_n14928 & ~new_n14939;
  assign new_n14941 = new_n14928 & new_n14939;
  assign new_n14942 = ~new_n14940 & ~new_n14941;
  assign new_n14943 = new_n14938 & new_n14942;
  assign new_n14944 = ~new_n14938 & ~new_n14942;
  assign new_n14945 = ~new_n12810 & ~new_n12813;
  assign new_n14946 = ~new_n12809 & ~new_n14945;
  assign new_n14947 = ~new_n14944 & new_n14946;
  assign new_n14948 = ~new_n14943 & ~new_n14947;
  assign new_n14949 = new_n14936 & new_n14948;
  assign new_n14950 = ~new_n14936 & ~new_n14948;
  assign new_n14951 = ~new_n14949 & ~new_n14950;
  assign new_n14952 = new_n14656 & ~new_n14951;
  assign new_n14953 = ~new_n14656 & new_n14951;
  assign new_n14954 = ~new_n14952 & ~new_n14953;
  assign new_n14955 = ~new_n12529 & ~new_n14608;
  assign new_n14956 = ~new_n14609 & ~new_n14955;
  assign new_n14957 = ~new_n12708 & ~new_n12818;
  assign new_n14958 = new_n14956 & new_n14957;
  assign new_n14959 = ~new_n14956 & ~new_n14957;
  assign new_n14960 = new_n14943 & new_n14946;
  assign new_n14961 = new_n14944 & ~new_n14946;
  assign new_n14962 = new_n14948 & ~new_n14961;
  assign new_n14963 = ~new_n14960 & ~new_n14962;
  assign new_n14964 = ~new_n14959 & ~new_n14963;
  assign new_n14965 = ~new_n14958 & ~new_n14964;
  assign new_n14966 = ~new_n14954 & ~new_n14965;
  assign new_n14967 = new_n14954 & new_n14965;
  assign n12406 = new_n14966 | new_n14967;
  assign new_n14969 = ~new_n7794 & ~new_n7795;
  assign new_n14970 = new_n7825 & new_n14969;
  assign new_n14971 = ~new_n7825 & ~new_n14969;
  assign n12463 = new_n14970 | new_n14971;
  assign new_n14973 = ~new_n12694 & new_n12702;
  assign new_n14974 = ~new_n12698 & new_n14973;
  assign new_n14975 = new_n12698 & ~new_n14973;
  assign n12503 = ~new_n14974 & ~new_n14975;
  assign new_n14977 = ~new_n7336 & ~new_n7337;
  assign new_n14978 = new_n7359 & ~new_n14977;
  assign new_n14979 = ~new_n7359 & new_n14977;
  assign n12515 = ~new_n14978 & ~new_n14979;
  assign new_n14981 = ~new_n14958 & ~new_n14959;
  assign new_n14982 = new_n14963 & ~new_n14981;
  assign new_n14983 = ~new_n14963 & new_n14981;
  assign n12616 = ~new_n14982 & ~new_n14983;
  assign new_n14985 = ~new_n11683 & ~new_n11684;
  assign new_n14986 = new_n11696 & ~new_n14985;
  assign new_n14987 = ~new_n11696 & new_n14985;
  assign n12839 = new_n14986 | new_n14987;
  assign new_n14989 = ~new_n4909 & ~new_n4910;
  assign new_n14990 = new_n4914 & ~new_n14989;
  assign new_n14991 = ~new_n4914 & new_n14989;
  assign n12968 = ~new_n14990 & ~new_n14991;
  assign new_n14993 = ~new_n5283 & ~new_n5285;
  assign n13002 = ~new_n5286 & ~new_n14993;
  assign new_n14995 = ~new_n14953 & ~new_n14965;
  assign new_n14996 = ~new_n14952 & ~new_n14995;
  assign new_n14997 = ~new_n14731 & ~new_n14742;
  assign new_n14998 = ~new_n14689 & ~new_n14726;
  assign new_n14999 = ~new_n14690 & ~new_n14998;
  assign new_n15000 = n411 & n4452;
  assign new_n15001 = n8230 & n12651;
  assign new_n15002 = n2458 & n7411;
  assign new_n15003 = new_n15001 & ~new_n15002;
  assign new_n15004 = ~new_n15001 & new_n15002;
  assign new_n15005 = ~new_n15003 & ~new_n15004;
  assign new_n15006 = new_n14612 & ~new_n14615;
  assign new_n15007 = ~new_n14616 & ~new_n15006;
  assign new_n15008 = ~new_n15005 & new_n15007;
  assign new_n15009 = new_n15005 & ~new_n15007;
  assign new_n15010 = ~new_n15008 & ~new_n15009;
  assign new_n15011 = n6149 & n7529;
  assign new_n15012 = ~n7161 & n7715;
  assign new_n15013 = ~new_n15011 & ~new_n15012;
  assign new_n15014 = new_n15011 & new_n15012;
  assign new_n15015 = ~new_n15013 & ~new_n15014;
  assign new_n15016 = new_n14633 & new_n15015;
  assign new_n15017 = ~new_n14633 & ~new_n15015;
  assign new_n15018 = ~new_n15016 & ~new_n15017;
  assign new_n15019 = new_n15010 & new_n15018;
  assign new_n15020 = ~new_n15010 & ~new_n15018;
  assign new_n15021 = ~new_n15019 & ~new_n15020;
  assign new_n15022 = ~new_n14626 & new_n14636;
  assign new_n15023 = ~new_n14625 & ~new_n15022;
  assign new_n15024 = ~new_n15021 & ~new_n15023;
  assign new_n15025 = new_n15021 & new_n15023;
  assign new_n15026 = ~new_n15024 & ~new_n15025;
  assign new_n15027 = ~new_n14622 & new_n14639;
  assign new_n15028 = ~new_n14621 & ~new_n15027;
  assign new_n15029 = new_n15026 & ~new_n15028;
  assign new_n15030 = ~new_n15026 & new_n15028;
  assign new_n15031 = ~new_n15029 & ~new_n15030;
  assign new_n15032 = ~new_n15000 & new_n15031;
  assign new_n15033 = new_n15000 & ~new_n15031;
  assign new_n15034 = ~new_n15032 & ~new_n15033;
  assign new_n15035 = new_n14999 & ~new_n15034;
  assign new_n15036 = ~new_n14999 & new_n15034;
  assign new_n15037 = ~new_n15035 & ~new_n15036;
  assign new_n15038 = n9475 & n10657;
  assign new_n15039 = n6826 & n10142;
  assign new_n15040 = ~new_n15038 & ~new_n15039;
  assign new_n15041 = new_n15038 & new_n15039;
  assign new_n15042 = ~new_n15040 & ~new_n15041;
  assign new_n15043 = ~new_n15037 & new_n15042;
  assign new_n15044 = new_n15037 & ~new_n15042;
  assign new_n15045 = ~new_n15043 & ~new_n15044;
  assign new_n15046 = new_n14795 & ~new_n14798;
  assign new_n15047 = ~new_n14799 & ~new_n15046;
  assign new_n15048 = new_n14779 & ~new_n14782;
  assign new_n15049 = ~new_n14783 & ~new_n15048;
  assign new_n15050 = ~new_n15047 & new_n15049;
  assign new_n15051 = new_n15047 & ~new_n15049;
  assign new_n15052 = ~new_n15050 & ~new_n15051;
  assign new_n15053 = ~new_n15045 & new_n15052;
  assign new_n15054 = new_n15045 & ~new_n15052;
  assign new_n15055 = ~new_n15053 & ~new_n15054;
  assign new_n15056 = new_n14997 & new_n15055;
  assign new_n15057 = ~new_n14997 & ~new_n15055;
  assign new_n15058 = ~new_n15056 & ~new_n15057;
  assign new_n15059 = ~new_n14919 & new_n14930;
  assign new_n15060 = ~new_n14918 & ~new_n15059;
  assign new_n15061 = ~new_n14905 & ~new_n14916;
  assign new_n15062 = ~new_n14863 & ~new_n14900;
  assign new_n15063 = ~new_n14864 & ~new_n15062;
  assign new_n15064 = n951 & n10805;
  assign new_n15065 = n353 & n767;
  assign new_n15066 = new_n15064 & ~new_n15065;
  assign new_n15067 = ~new_n15064 & new_n15065;
  assign new_n15068 = ~new_n15066 & ~new_n15067;
  assign new_n15069 = n124 & n401;
  assign new_n15070 = n11537 & n12263;
  assign new_n15071 = ~new_n15069 & ~new_n15070;
  assign new_n15072 = new_n15069 & new_n15070;
  assign new_n15073 = ~new_n15071 & ~new_n15072;
  assign new_n15074 = ~new_n15068 & new_n15073;
  assign new_n15075 = new_n15068 & ~new_n15073;
  assign new_n15076 = ~new_n15074 & ~new_n15075;
  assign new_n15077 = n3085 & n4419;
  assign new_n15078 = n3178 & n12372;
  assign new_n15079 = ~new_n15077 & new_n15078;
  assign new_n15080 = new_n15077 & ~new_n15078;
  assign new_n15081 = ~new_n15079 & ~new_n15080;
  assign new_n15082 = ~new_n15076 & new_n15081;
  assign new_n15083 = new_n15076 & ~new_n15081;
  assign new_n15084 = ~new_n15082 & ~new_n15083;
  assign new_n15085 = new_n15063 & ~new_n15084;
  assign new_n15086 = ~new_n15063 & new_n15084;
  assign new_n15087 = ~new_n15085 & ~new_n15086;
  assign new_n15088 = new_n15061 & ~new_n15087;
  assign new_n15089 = ~new_n15061 & new_n15087;
  assign new_n15090 = ~new_n15088 & ~new_n15089;
  assign new_n15091 = new_n14692 & ~new_n14695;
  assign new_n15092 = ~new_n14696 & ~new_n15091;
  assign new_n15093 = new_n14723 & new_n15092;
  assign new_n15094 = ~new_n14723 & ~new_n15092;
  assign new_n15095 = ~new_n15093 & ~new_n15094;
  assign new_n15096 = ~new_n14706 & new_n14716;
  assign new_n15097 = ~new_n14705 & ~new_n15096;
  assign new_n15098 = n469 & n11324;
  assign new_n15099 = new_n14708 & ~new_n14711;
  assign new_n15100 = ~new_n14712 & ~new_n15099;
  assign new_n15101 = n2068 & n12065;
  assign new_n15102 = n11180 & n12348;
  assign new_n15103 = ~new_n15101 & new_n15102;
  assign new_n15104 = new_n15101 & ~new_n15102;
  assign new_n15105 = ~new_n15103 & ~new_n15104;
  assign new_n15106 = ~new_n15100 & ~new_n15105;
  assign new_n15107 = new_n15100 & new_n15105;
  assign new_n15108 = ~new_n15106 & ~new_n15107;
  assign new_n15109 = ~new_n15098 & new_n15108;
  assign new_n15110 = new_n15098 & ~new_n15108;
  assign new_n15111 = ~new_n15109 & ~new_n15110;
  assign new_n15112 = ~new_n15097 & new_n15111;
  assign new_n15113 = new_n15097 & ~new_n15111;
  assign new_n15114 = ~new_n15112 & ~new_n15113;
  assign new_n15115 = n9216 & n12912;
  assign new_n15116 = n8183 & n12284;
  assign new_n15117 = new_n15115 & new_n15116;
  assign new_n15118 = ~new_n15115 & ~new_n15116;
  assign new_n15119 = ~new_n15117 & ~new_n15118;
  assign new_n15120 = new_n15114 & ~new_n15119;
  assign new_n15121 = ~new_n15114 & new_n15119;
  assign new_n15122 = ~new_n15120 & ~new_n15121;
  assign new_n15123 = ~new_n15095 & ~new_n15122;
  assign new_n15124 = new_n15095 & new_n15122;
  assign new_n15125 = ~new_n15123 & ~new_n15124;
  assign new_n15126 = ~new_n15090 & new_n15125;
  assign new_n15127 = new_n15090 & ~new_n15125;
  assign new_n15128 = ~new_n15126 & ~new_n15127;
  assign new_n15129 = new_n15060 & new_n15128;
  assign new_n15130 = ~new_n15060 & ~new_n15128;
  assign new_n15131 = ~new_n15129 & ~new_n15130;
  assign new_n15132 = new_n15058 & ~new_n15131;
  assign new_n15133 = ~new_n15058 & new_n15131;
  assign new_n15134 = ~new_n15132 & ~new_n15133;
  assign new_n15135 = ~new_n14818 & ~new_n14829;
  assign new_n15136 = ~new_n14651 & ~new_n14654;
  assign new_n15137 = new_n15135 & new_n15136;
  assign new_n15138 = ~new_n15135 & ~new_n15136;
  assign new_n15139 = ~new_n15137 & ~new_n15138;
  assign new_n15140 = n4122 & n8466;
  assign new_n15141 = n2590 & n2737;
  assign new_n15142 = new_n15140 & ~new_n15141;
  assign new_n15143 = ~new_n15140 & new_n15141;
  assign new_n15144 = ~new_n15142 & ~new_n15143;
  assign new_n15145 = n9 & n9846;
  assign new_n15146 = n5031 & n11350;
  assign new_n15147 = ~new_n15145 & ~new_n15146;
  assign new_n15148 = new_n15145 & new_n15146;
  assign new_n15149 = ~new_n15147 & ~new_n15148;
  assign new_n15150 = ~new_n15144 & new_n15149;
  assign new_n15151 = new_n15144 & ~new_n15149;
  assign new_n15152 = ~new_n15150 & ~new_n15151;
  assign new_n15153 = n4998 & n8506;
  assign new_n15154 = n2592 & n12408;
  assign new_n15155 = ~new_n15153 & new_n15154;
  assign new_n15156 = new_n15153 & ~new_n15154;
  assign new_n15157 = ~new_n15155 & ~new_n15156;
  assign new_n15158 = n5536 & n8768;
  assign new_n15159 = n772 & n11061;
  assign new_n15160 = new_n15158 & ~new_n15159;
  assign new_n15161 = ~new_n15158 & new_n15159;
  assign new_n15162 = ~new_n15160 & ~new_n15161;
  assign new_n15163 = ~new_n15157 & ~new_n15162;
  assign new_n15164 = new_n15157 & new_n15162;
  assign new_n15165 = ~new_n15163 & ~new_n15164;
  assign new_n15166 = new_n14866 & ~new_n14869;
  assign new_n15167 = ~new_n14870 & ~new_n15166;
  assign new_n15168 = new_n15165 & new_n15167;
  assign new_n15169 = ~new_n15165 & ~new_n15167;
  assign new_n15170 = ~new_n15168 & ~new_n15169;
  assign new_n15171 = ~new_n15152 & new_n15170;
  assign new_n15172 = new_n15152 & ~new_n15170;
  assign new_n15173 = ~new_n15171 & ~new_n15172;
  assign new_n15174 = new_n14882 & ~new_n14885;
  assign new_n15175 = ~new_n14886 & ~new_n15174;
  assign new_n15176 = n22 & n10168;
  assign new_n15177 = n11396 & n12592;
  assign new_n15178 = ~new_n15176 & new_n15177;
  assign new_n15179 = new_n15176 & ~new_n15177;
  assign new_n15180 = ~new_n15178 & ~new_n15179;
  assign new_n15181 = new_n15175 & ~new_n15180;
  assign new_n15182 = ~new_n15175 & new_n15180;
  assign new_n15183 = ~new_n15181 & ~new_n15182;
  assign new_n15184 = ~new_n14879 & new_n14890;
  assign new_n15185 = ~new_n14880 & ~new_n15184;
  assign new_n15186 = ~new_n15183 & ~new_n15185;
  assign new_n15187 = new_n15183 & new_n15185;
  assign new_n15188 = ~new_n15186 & ~new_n15187;
  assign new_n15189 = ~new_n15173 & new_n15188;
  assign new_n15190 = new_n15173 & ~new_n15188;
  assign new_n15191 = ~new_n15189 & ~new_n15190;
  assign new_n15192 = ~new_n14776 & ~new_n14813;
  assign new_n15193 = ~new_n14777 & ~new_n15192;
  assign new_n15194 = new_n14897 & new_n15193;
  assign new_n15195 = ~new_n14897 & ~new_n15193;
  assign new_n15196 = ~new_n15194 & ~new_n15195;
  assign new_n15197 = new_n15191 & new_n15196;
  assign new_n15198 = ~new_n15191 & ~new_n15196;
  assign new_n15199 = ~new_n15197 & ~new_n15198;
  assign new_n15200 = new_n14810 & ~new_n15199;
  assign new_n15201 = ~new_n14810 & new_n15199;
  assign new_n15202 = ~new_n15200 & ~new_n15201;
  assign new_n15203 = ~new_n14643 & new_n14647;
  assign new_n15204 = ~new_n14644 & ~new_n15203;
  assign new_n15205 = ~new_n14792 & new_n14803;
  assign new_n15206 = ~new_n14793 & ~new_n15205;
  assign new_n15207 = n6668 & n11734;
  assign new_n15208 = n5715 & n7772;
  assign new_n15209 = ~n7812 & new_n15208;
  assign new_n15210 = n7812 & ~new_n15208;
  assign new_n15211 = ~new_n15209 & ~new_n15210;
  assign new_n15212 = ~new_n15207 & new_n15211;
  assign new_n15213 = new_n15207 & ~new_n15211;
  assign new_n15214 = ~new_n15212 & ~new_n15213;
  assign new_n15215 = new_n15206 & new_n15214;
  assign new_n15216 = ~new_n15206 & ~new_n15214;
  assign new_n15217 = ~new_n15215 & ~new_n15216;
  assign new_n15218 = ~new_n15204 & ~new_n15217;
  assign new_n15219 = new_n15204 & new_n15217;
  assign new_n15220 = ~new_n15218 & ~new_n15219;
  assign new_n15221 = ~new_n15202 & new_n15220;
  assign new_n15222 = new_n15202 & ~new_n15220;
  assign new_n15223 = ~new_n15221 & ~new_n15222;
  assign new_n15224 = ~new_n15139 & ~new_n15223;
  assign new_n15225 = new_n15139 & new_n15223;
  assign new_n15226 = ~new_n15224 & ~new_n15225;
  assign new_n15227 = ~new_n14934 & new_n14948;
  assign new_n15228 = ~new_n14935 & ~new_n15227;
  assign new_n15229 = new_n15226 & new_n15228;
  assign new_n15230 = ~new_n15226 & ~new_n15228;
  assign new_n15231 = ~new_n15229 & ~new_n15230;
  assign new_n15232 = new_n15134 & ~new_n15231;
  assign new_n15233 = ~new_n15134 & new_n15231;
  assign new_n15234 = ~new_n15232 & ~new_n15233;
  assign new_n15235 = ~new_n14996 & ~new_n15234;
  assign new_n15236 = new_n14996 & new_n15234;
  assign n13035 = new_n15235 | new_n15236;
endmodule


