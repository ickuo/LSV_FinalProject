// Benchmark "top" written by ABC on Sun Dec 21 18:12:47 2025

module top ( 
    n11, n21, n29, n40, n45, n50, n52, n54, n56, n58, n71, n77, n82, n86,
    n87, n94, n107, n117, n138, n143, n153, n155, n156, n159, n200, n219,
    n220, n222, n223, n243, n244, n246, n251, n254, n262, n268, n273, n284,
    n288, n293, n299, n300, n307, n310, n312, n314, n315, n318, n341, n344,
    n346, n374, n376, n380, n391, n392, n399, n408, n409, n416, n420, n430,
    n477, n478, n487, n489, n502, n506, n507, n510, n545, n559, n560, n561,
    n567, n574, n581, n582, n589, n593, n598, n600, n607, n608, n609, n626,
    n641, n645, n663, n671, n676, n690, n695, n701, n710, n727, n729, n734,
    n742, n743, n755, n769, n775, n778, n779, n787, n790, n823, n831, n832,
    n839, n849, n879, n882, n885, n905, n920, n936, n947, n953, n961, n969,
    n980, n984, n986, n992, n997, n1023, n1040, n1044, n1054, n1061, n1071,
    n1095, n1103, n1114, n1121, n1138, n1152, n1154, n1156, n1164, n1172,
    n1175, n1187, n1191, n1193, n1205, n1225, n1227, n1239, n1246, n1250,
    n1263, n1278, n1281, n1283, n1286, n1289, n1299, n1301, n1305, n1345,
    n1346, n1350, n1361, n1386, n1387, n1389, n1393, n1401, n1411, n1415,
    n1418, n1428, n1435, n1438, n1443, n1446, n1448, n1463, n1470, n1474,
    n1476, n1500, n1502, n1506, n1516, n1520, n1521, n1523, n1536, n1566,
    n1569, n1576, n1586, n1592, n1609, n1613, n1616, n1626, n1627, n1644,
    n1647, n1656, n1750, n1753,
    n22, n23, n27, n30, n85, n112, n126, n130, n161, n164, n173, n181,
    n184, n216, n230, n233, n247, n275, n292, n301, n304, n337, n352, n362,
    n364, n370, n378, n396, n417, n428, n453, n457, n460, n497, n498, n501,
    n509, n516, n517, n534, n553, n585, n595, n597, n625, n638, n640, n669,
    n693, n714, n719, n726, n773, n782, n794, n821, n842, n894, n916, n918,
    n952, n990, n1006, n1017, n1042, n1050, n1051, n1058, n1060, n1063,
    n1065, n1177, n1186, n1195, n1209, n1211, n1231, n1234, n1253, n1285,
    n1288, n1292, n1296, n1302, n1306, n1320, n1322, n1337, n1359, n1368,
    n1375, n1391, n1420, n1421, n1427, n1527, n1534, n1547, n1548, n1588,
    n1594, n1632, n1639, n1645, n1687, n1729, n1738, n1752  );
  input  n11, n21, n29, n40, n45, n50, n52, n54, n56, n58, n71, n77, n82,
    n86, n87, n94, n107, n117, n138, n143, n153, n155, n156, n159, n200,
    n219, n220, n222, n223, n243, n244, n246, n251, n254, n262, n268, n273,
    n284, n288, n293, n299, n300, n307, n310, n312, n314, n315, n318, n341,
    n344, n346, n374, n376, n380, n391, n392, n399, n408, n409, n416, n420,
    n430, n477, n478, n487, n489, n502, n506, n507, n510, n545, n559, n560,
    n561, n567, n574, n581, n582, n589, n593, n598, n600, n607, n608, n609,
    n626, n641, n645, n663, n671, n676, n690, n695, n701, n710, n727, n729,
    n734, n742, n743, n755, n769, n775, n778, n779, n787, n790, n823, n831,
    n832, n839, n849, n879, n882, n885, n905, n920, n936, n947, n953, n961,
    n969, n980, n984, n986, n992, n997, n1023, n1040, n1044, n1054, n1061,
    n1071, n1095, n1103, n1114, n1121, n1138, n1152, n1154, n1156, n1164,
    n1172, n1175, n1187, n1191, n1193, n1205, n1225, n1227, n1239, n1246,
    n1250, n1263, n1278, n1281, n1283, n1286, n1289, n1299, n1301, n1305,
    n1345, n1346, n1350, n1361, n1386, n1387, n1389, n1393, n1401, n1411,
    n1415, n1418, n1428, n1435, n1438, n1443, n1446, n1448, n1463, n1470,
    n1474, n1476, n1500, n1502, n1506, n1516, n1520, n1521, n1523, n1536,
    n1566, n1569, n1576, n1586, n1592, n1609, n1613, n1616, n1626, n1627,
    n1644, n1647, n1656, n1750, n1753;
  output n22, n23, n27, n30, n85, n112, n126, n130, n161, n164, n173, n181,
    n184, n216, n230, n233, n247, n275, n292, n301, n304, n337, n352, n362,
    n364, n370, n378, n396, n417, n428, n453, n457, n460, n497, n498, n501,
    n509, n516, n517, n534, n553, n585, n595, n597, n625, n638, n640, n669,
    n693, n714, n719, n726, n773, n782, n794, n821, n842, n894, n916, n918,
    n952, n990, n1006, n1017, n1042, n1050, n1051, n1058, n1060, n1063,
    n1065, n1177, n1186, n1195, n1209, n1211, n1231, n1234, n1253, n1285,
    n1288, n1292, n1296, n1302, n1306, n1320, n1322, n1337, n1359, n1368,
    n1375, n1391, n1420, n1421, n1427, n1527, n1534, n1547, n1548, n1588,
    n1594, n1632, n1639, n1645, n1687, n1729, n1738, n1752;
  wire new_n316, new_n317, new_n318_1, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337_1, new_n338, new_n339, new_n340, new_n341_1,
    new_n342, new_n343, new_n344_1, new_n345, new_n346_1, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352_1, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362_1, new_n363, new_n364_1, new_n365, new_n366, new_n367,
    new_n368, new_n369, new_n370_1, new_n371, new_n372, new_n373,
    new_n374_1, new_n375, new_n376_1, new_n377, new_n378_1, new_n379,
    new_n380_1, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391_1, new_n392_1,
    new_n393, new_n394, new_n395, new_n396_1, new_n397, new_n398,
    new_n399_1, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408_1, new_n409_1, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416_1, new_n417_1,
    new_n418, new_n419, new_n420_1, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428_1, new_n429, new_n430_1,
    new_n431, new_n432, new_n433, new_n434, new_n435, new_n436, new_n437,
    new_n438, new_n439, new_n440, new_n441, new_n442, new_n443, new_n444,
    new_n445, new_n446, new_n447, new_n448, new_n449, new_n450, new_n451,
    new_n452, new_n453_1, new_n454, new_n455, new_n456, new_n457_1,
    new_n458, new_n459, new_n460_1, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477_1,
    new_n478_1, new_n479, new_n480, new_n481, new_n482, new_n483, new_n484,
    new_n485, new_n486, new_n487_1, new_n488, new_n489_1, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497_1,
    new_n498_1, new_n499, new_n500, new_n501_1, new_n502_1, new_n503,
    new_n504, new_n505, new_n506_1, new_n507_1, new_n508, new_n509_1,
    new_n510_1, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516_1, new_n517_1, new_n518, new_n519, new_n520, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534_1, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545_1, new_n546, new_n547, new_n548, new_n551,
    new_n553_1, new_n554, new_n556, new_n557, new_n558, new_n559_1,
    new_n560_1, new_n561_1, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567_1, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574_1, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581_1, new_n582_1, new_n583, new_n584, new_n585_1,
    new_n586, new_n587, new_n588, new_n589_1, new_n590, new_n591, new_n592,
    new_n593_1, new_n594, new_n595_1, new_n596, new_n597_1, new_n598_1,
    new_n599, new_n600_1, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607_1, new_n608_1, new_n609_1, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625_1,
    new_n626_1, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638_1, new_n639,
    new_n640_1, new_n641_1, new_n642, new_n643, new_n644, new_n645_1,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663_1, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669_1, new_n670, new_n671_1, new_n672,
    new_n673, new_n674, new_n675, new_n676_1, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690_1, new_n691, new_n692,
    new_n693_1, new_n694, new_n695_1, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701_1, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710_1, new_n711, new_n712,
    new_n713, new_n714_1, new_n715, new_n716, new_n717, new_n718,
    new_n719_1, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726_1, new_n727_1, new_n728, new_n729_1, new_n730, new_n731,
    new_n732, new_n733, new_n734_1, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742_1, new_n743_1, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755_1, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769_1, new_n770, new_n771, new_n772,
    new_n773_1, new_n774, new_n775_1, new_n776, new_n777, new_n778_1,
    new_n779_1, new_n780, new_n781, new_n782_1, new_n783, new_n784,
    new_n785, new_n786, new_n787_1, new_n788, new_n789, new_n790_1,
    new_n791, new_n792, new_n793, new_n794_1, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821_1, new_n822, new_n823_1, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831_1,
    new_n832_1, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839_1, new_n840, new_n841, new_n842_1, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849_1, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879_1,
    new_n880, new_n881, new_n882_1, new_n883, new_n885_1, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894_1,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905_1, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916_1,
    new_n917, new_n918_1, new_n919, new_n920_1, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936_1, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947_1, new_n948, new_n949, new_n950, new_n951,
    new_n952_1, new_n953_1, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961_1, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969_1, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980_1, new_n981, new_n982, new_n983, new_n984_1,
    new_n985, new_n986_1, new_n987, new_n988, new_n989, new_n990_1,
    new_n991, new_n992_1, new_n993, new_n994, new_n995, new_n996,
    new_n997_1, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006_1, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017_1, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1025, new_n1026, new_n1027, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040_1, new_n1041, new_n1042_1, new_n1043,
    new_n1044_1, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050_1, new_n1051_1, new_n1052, new_n1053, new_n1054_1, new_n1055,
    new_n1056, new_n1057, new_n1058_1, new_n1059, new_n1060_1, new_n1061_1,
    new_n1062, new_n1063_1, new_n1064, new_n1065_1, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071_1, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095_1, new_n1096, new_n1097,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103_1,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114_1, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1127, new_n1128, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138_1, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1149, new_n1150, new_n1151,
    new_n1152_1, new_n1153, new_n1155, new_n1156_1, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164_1, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172_1, new_n1173, new_n1174, new_n1175_1, new_n1176, new_n1177_1,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186_1, new_n1187_1, new_n1188, new_n1189,
    new_n1190, new_n1191_1, new_n1192, new_n1193_1, new_n1194, new_n1195_1,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205_1, new_n1206, new_n1207,
    new_n1208, new_n1209_1, new_n1210, new_n1211_1, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225_1,
    new_n1226, new_n1227_1, new_n1228, new_n1229, new_n1230, new_n1231_1,
    new_n1233, new_n1234_1, new_n1236, new_n1238, new_n1239_1, new_n1240,
    new_n1241, new_n1244, new_n1245, new_n1246_1, new_n1247, new_n1248,
    new_n1250_1, new_n1251, new_n1252, new_n1254, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263_1,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278_1, new_n1279, new_n1280, new_n1281_1,
    new_n1282, new_n1283_1, new_n1284, new_n1285_1, new_n1286_1, new_n1287,
    new_n1288_1, new_n1289_1, new_n1290, new_n1291, new_n1292_1, new_n1293,
    new_n1294, new_n1295, new_n1296_1, new_n1297, new_n1298, new_n1299_1,
    new_n1300, new_n1301_1, new_n1302_1, new_n1303, new_n1304, new_n1305_1,
    new_n1306_1, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320_1, new_n1321, new_n1322_1, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337_1, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345_1, new_n1346_1, new_n1347,
    new_n1348, new_n1349, new_n1350_1, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359_1,
    new_n1360, new_n1361_1, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368_1, new_n1369, new_n1371, new_n1372,
    new_n1374, new_n1375_1, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386_1,
    new_n1387_1, new_n1388, new_n1389_1, new_n1390, new_n1391_1, new_n1392,
    new_n1393_1, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401_1, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411_1, new_n1412, new_n1413, new_n1414, new_n1415_1, new_n1416,
    new_n1417, new_n1418_1, new_n1419, new_n1420_1, new_n1421_1, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427_1, new_n1428_1,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435_1, new_n1436, new_n1437, new_n1438_1, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443_1, new_n1444, new_n1445, new_n1446_1,
    new_n1447, new_n1448_1, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463_1, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470_1,
    new_n1471, new_n1472, new_n1473, new_n1474_1, new_n1475, new_n1476_1,
    new_n1477, new_n1478, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500_1,
    new_n1501, new_n1502_1, new_n1503, new_n1504, new_n1505, new_n1507,
    new_n1508, new_n1509, new_n1510, new_n1511, new_n1512, new_n1513,
    new_n1514, new_n1515, new_n1516_1, new_n1517, new_n1518, new_n1519,
    new_n1520_1, new_n1521_1, new_n1522, new_n1523_1, new_n1524, new_n1525,
    new_n1526, new_n1527_1, new_n1528, new_n1529, new_n1530, new_n1531,
    new_n1532, new_n1533, new_n1534_1, new_n1535, new_n1536_1, new_n1537,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545, new_n1546, new_n1547_1, new_n1548_1, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1558, new_n1559, new_n1560, new_n1561,
    new_n1562, new_n1563, new_n1564, new_n1565, new_n1566_1, new_n1567,
    new_n1568, new_n1569_1, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576_1, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586_1, new_n1587, new_n1588_1, new_n1589, new_n1590, new_n1591,
    new_n1592_1, new_n1593, new_n1594_1, new_n1595, new_n1596, new_n1597,
    new_n1598, new_n1599, new_n1600, new_n1601, new_n1602, new_n1603,
    new_n1604, new_n1605, new_n1606, new_n1607, new_n1608, new_n1609_1,
    new_n1610, new_n1611, new_n1612, new_n1613_1, new_n1614, new_n1615,
    new_n1616_1, new_n1618, new_n1620, new_n1622, new_n1623, new_n1624,
    new_n1625, new_n1627_1, new_n1629, new_n1631, new_n1633, new_n1634,
    new_n1635, new_n1637, new_n1639_1, new_n1641, new_n1642, new_n1643,
    new_n1644_1, new_n1645_1, new_n1646, new_n1647_1, new_n1648, new_n1649,
    new_n1650, new_n1651, new_n1652, new_n1653, new_n1654, new_n1655,
    new_n1656_1, new_n1657, new_n1658, new_n1659, new_n1660, new_n1661,
    new_n1662, new_n1663, new_n1664, new_n1665, new_n1666, new_n1667,
    new_n1668, new_n1669, new_n1670, new_n1671, new_n1672, new_n1673,
    new_n1674, new_n1675, new_n1676, new_n1677, new_n1678, new_n1679,
    new_n1680, new_n1681, new_n1682, new_n1683, new_n1684, new_n1685,
    new_n1686, new_n1687_1, new_n1688, new_n1689, new_n1690, new_n1691,
    new_n1692, new_n1693, new_n1694, new_n1695, new_n1696, new_n1697,
    new_n1698, new_n1699, new_n1700, new_n1701, new_n1702, new_n1703,
    new_n1704, new_n1705, new_n1706, new_n1707, new_n1708, new_n1709,
    new_n1710, new_n1711, new_n1712, new_n1713, new_n1714, new_n1715,
    new_n1716, new_n1717, new_n1718, new_n1719, new_n1720, new_n1722,
    new_n1723, new_n1724, new_n1726, new_n1728, new_n1730, new_n1732,
    new_n1733, new_n1734, new_n1735, new_n1737, new_n1739, new_n1740,
    new_n1741, new_n1742, new_n1744, new_n1745, new_n1746;
  assign new_n316 = n11 & n984;
  assign new_n317 = ~n220 & n1239;
  assign new_n318_1 = ~new_n316 & ~new_n317;
  assign new_n319 = ~n1263 & new_n318_1;
  assign new_n320 = n1263 & ~new_n318_1;
  assign new_n321 = ~new_n319 & ~new_n320;
  assign new_n322 = ~n391 & n1239;
  assign new_n323 = ~new_n316 & ~new_n322;
  assign new_n324 = ~n346 & new_n323;
  assign new_n325 = n346 & ~new_n323;
  assign new_n326 = ~n905 & n1239;
  assign new_n327 = ~new_n316 & ~new_n326;
  assign new_n328 = ~n399 & new_n327;
  assign new_n329 = n399 & ~new_n327;
  assign new_n330 = ~new_n328 & ~new_n329;
  assign new_n331 = n1239 & ~n1278;
  assign new_n332 = ~new_n316 & ~new_n331;
  assign new_n333 = ~n980 & new_n332;
  assign new_n334 = new_n330 & new_n333;
  assign new_n335 = ~new_n328 & ~new_n334;
  assign new_n336 = ~new_n325 & ~new_n335;
  assign new_n337_1 = ~new_n324 & ~new_n336;
  assign new_n338 = n980 & ~new_n332;
  assign new_n339 = new_n330 & ~new_n338;
  assign new_n340 = ~new_n333 & new_n339;
  assign new_n341_1 = ~new_n324 & ~new_n325;
  assign new_n342 = new_n340 & new_n341_1;
  assign new_n343 = n1239 & ~n1435;
  assign new_n344_1 = ~new_n316 & ~new_n343;
  assign new_n345 = ~n318 & new_n344_1;
  assign new_n346_1 = n318 & ~new_n344_1;
  assign new_n347 = n1239 & n1474;
  assign new_n348 = ~n1239 & n1506;
  assign new_n349 = ~new_n347 & ~new_n348;
  assign new_n350 = n1592 & new_n349;
  assign new_n351 = ~n1592 & ~new_n349;
  assign new_n352_1 = n58 & n1239;
  assign new_n353 = ~n1239 & n1443;
  assign new_n354 = ~new_n352_1 & ~new_n353;
  assign new_n355 = ~n1616 & ~new_n354;
  assign new_n356 = n1616 & new_n354;
  assign new_n357 = n598 & n1239;
  assign new_n358 = ~n1239 & n1647;
  assign new_n359 = ~new_n357 & ~new_n358;
  assign new_n360 = ~n1446 & ~new_n359;
  assign new_n361 = n1239 & n1415;
  assign new_n362_1 = ~n1239 & n1246;
  assign new_n363 = ~new_n361 & ~new_n362_1;
  assign new_n364_1 = ~n1345 & ~new_n363;
  assign new_n365 = n1446 & new_n359;
  assign new_n366 = new_n364_1 & ~new_n365;
  assign new_n367 = ~new_n360 & ~new_n366;
  assign new_n368 = ~new_n356 & ~new_n367;
  assign new_n369 = ~new_n355 & ~new_n368;
  assign new_n370_1 = ~new_n351 & new_n369;
  assign new_n371 = ~new_n350 & ~new_n370_1;
  assign new_n372 = ~new_n346_1 & new_n371;
  assign new_n373 = ~new_n345 & ~new_n372;
  assign new_n374_1 = n1345 & new_n363;
  assign new_n375 = ~new_n364_1 & ~new_n374_1;
  assign new_n376_1 = ~new_n355 & ~new_n356;
  assign new_n377 = ~new_n360 & ~new_n365;
  assign new_n378_1 = new_n376_1 & new_n377;
  assign new_n379 = new_n375 & new_n378_1;
  assign new_n380_1 = ~new_n345 & ~new_n346_1;
  assign new_n381 = ~new_n350 & ~new_n351;
  assign new_n382 = new_n380_1 & new_n381;
  assign new_n383 = new_n379 & new_n382;
  assign new_n384 = n1239 & n1350;
  assign new_n385 = n262 & ~n1239;
  assign new_n386 = ~new_n384 & ~new_n385;
  assign new_n387 = ~n1301 & ~new_n386;
  assign new_n388 = n1301 & new_n386;
  assign new_n389 = ~new_n387 & ~new_n388;
  assign new_n390 = n676 & n1239;
  assign new_n391_1 = n1154 & ~n1239;
  assign new_n392_1 = ~new_n390 & ~new_n391_1;
  assign new_n393 = n1566 & new_n392_1;
  assign new_n394 = ~n1566 & ~new_n392_1;
  assign new_n395 = ~new_n393 & ~new_n394;
  assign new_n396_1 = new_n389 & new_n395;
  assign new_n397 = n251 & n1239;
  assign new_n398 = n1172 & ~n1239;
  assign new_n399_1 = ~new_n397 & ~new_n398;
  assign new_n400 = ~n408 & ~new_n399_1;
  assign new_n401 = n408 & new_n399_1;
  assign new_n402 = n1239 & n1516;
  assign new_n403 = n710 & ~n1239;
  assign new_n404 = ~new_n402 & ~new_n403;
  assign new_n405 = n1476 & new_n404;
  assign new_n406 = ~n1476 & ~new_n404;
  assign new_n407 = n790 & n1239;
  assign new_n408_1 = ~n1239 & n1521;
  assign new_n409_1 = ~new_n407 & ~new_n408_1;
  assign new_n410 = ~n823 & ~new_n409_1;
  assign new_n411 = n823 & new_n409_1;
  assign new_n412 = n1239 & n1576;
  assign new_n413 = ~n1239 & n1283;
  assign new_n414 = ~new_n412 & ~new_n413;
  assign new_n415 = ~n153 & ~new_n414;
  assign new_n416_1 = n153 & new_n414;
  assign new_n417_1 = n82 & n1239;
  assign new_n418 = n1061 & ~n1239;
  assign new_n419 = ~new_n417_1 & ~new_n418;
  assign new_n420_1 = ~n1401 & ~new_n419;
  assign new_n421 = ~new_n416_1 & new_n420_1;
  assign new_n422 = ~new_n415 & ~new_n421;
  assign new_n423 = ~new_n411 & ~new_n422;
  assign new_n424 = ~new_n410 & ~new_n423;
  assign new_n425 = ~new_n406 & new_n424;
  assign new_n426 = ~new_n405 & ~new_n425;
  assign new_n427 = ~new_n401 & new_n426;
  assign new_n428_1 = ~new_n400 & ~new_n427;
  assign new_n429 = n645 & n1239;
  assign new_n430_1 = n87 & ~n1239;
  assign new_n431 = ~new_n429 & ~new_n430_1;
  assign new_n432 = ~n374 & ~new_n431;
  assign new_n433 = n374 & new_n431;
  assign new_n434 = ~new_n432 & ~new_n433;
  assign new_n435 = n268 & n1239;
  assign new_n436 = n600 & ~n1239;
  assign new_n437 = ~new_n435 & ~new_n436;
  assign new_n438 = ~n567 & ~new_n437;
  assign new_n439 = n567 & new_n437;
  assign new_n440 = ~new_n438 & ~new_n439;
  assign new_n441 = new_n434 & new_n440;
  assign new_n442 = n1239 & n1393;
  assign new_n443 = n254 & ~n1239;
  assign new_n444 = ~new_n442 & ~new_n443;
  assign new_n445 = n1463 & new_n444;
  assign new_n446 = ~n1463 & ~new_n444;
  assign new_n447 = ~new_n445 & ~new_n446;
  assign new_n448 = n312 & n1239;
  assign new_n449 = n307 & ~n1239;
  assign new_n450 = ~new_n448 & ~new_n449;
  assign new_n451 = ~n222 & ~new_n450;
  assign new_n452 = n222 & new_n450;
  assign new_n453_1 = ~new_n451 & ~new_n452;
  assign new_n454 = n1239 & n1609;
  assign new_n455 = n54 & ~n1239;
  assign new_n456 = ~new_n454 & ~new_n455;
  assign new_n457_1 = n608 & new_n456;
  assign new_n458 = ~n608 & ~new_n456;
  assign new_n459 = ~new_n457_1 & ~new_n458;
  assign new_n460_1 = n310 & n1239;
  assign new_n461 = n1175 & ~n1239;
  assign new_n462 = ~new_n460_1 & ~new_n461;
  assign new_n463 = n1071 & new_n462;
  assign new_n464 = ~n1071 & ~new_n462;
  assign new_n465 = ~new_n463 & ~new_n464;
  assign new_n466 = new_n459 & new_n465;
  assign new_n467 = n219 & n1239;
  assign new_n468 = n409 & ~n1239;
  assign new_n469 = ~new_n467 & ~new_n468;
  assign new_n470 = n45 & new_n469;
  assign new_n471 = ~n45 & ~new_n469;
  assign new_n472 = ~new_n470 & ~new_n471;
  assign new_n473 = n1239 & n1569;
  assign new_n474 = ~n1239 & n1250;
  assign new_n475 = ~new_n473 & ~new_n474;
  assign new_n476 = ~n695 & ~new_n475;
  assign new_n477_1 = n510 & ~n1239;
  assign new_n478_1 = ~n1205 & new_n477_1;
  assign new_n479 = n695 & new_n475;
  assign new_n480 = new_n478_1 & ~new_n479;
  assign new_n481 = ~new_n476 & ~new_n480;
  assign new_n482 = new_n472 & ~new_n481;
  assign new_n483 = new_n466 & new_n482;
  assign new_n484 = ~new_n464 & ~new_n471;
  assign new_n485 = ~new_n463 & ~new_n484;
  assign new_n486 = ~new_n457_1 & new_n485;
  assign new_n487_1 = ~new_n458 & ~new_n486;
  assign new_n488 = ~new_n483 & new_n487_1;
  assign new_n489_1 = ~n510 & ~n1239;
  assign new_n490 = n1205 & new_n489_1;
  assign new_n491 = ~new_n478_1 & ~new_n490;
  assign new_n492 = ~new_n476 & ~new_n479;
  assign new_n493 = new_n472 & new_n492;
  assign new_n494 = new_n491 & new_n493;
  assign new_n495 = new_n465 & new_n494;
  assign new_n496 = new_n459 & new_n495;
  assign new_n497_1 = n545 & new_n496;
  assign new_n498_1 = new_n488 & ~new_n497_1;
  assign new_n499 = new_n453_1 & ~new_n498_1;
  assign new_n500 = new_n447 & new_n499;
  assign new_n501_1 = new_n441 & new_n500;
  assign new_n502_1 = ~new_n445 & new_n451;
  assign new_n503 = ~new_n446 & ~new_n502_1;
  assign new_n504 = ~new_n439 & ~new_n503;
  assign new_n505 = ~new_n438 & ~new_n504;
  assign new_n506_1 = ~new_n433 & ~new_n505;
  assign new_n507_1 = ~new_n432 & ~new_n506_1;
  assign new_n508 = ~new_n501_1 & new_n507_1;
  assign new_n509_1 = n1401 & new_n419;
  assign new_n510_1 = ~new_n420_1 & ~new_n509_1;
  assign new_n511 = ~new_n410 & ~new_n411;
  assign new_n512 = ~new_n415 & ~new_n416_1;
  assign new_n513 = new_n511 & new_n512;
  assign new_n514 = new_n510_1 & new_n513;
  assign new_n515 = ~new_n400 & ~new_n401;
  assign new_n516_1 = ~new_n405 & ~new_n406;
  assign new_n517_1 = new_n515 & new_n516_1;
  assign new_n518 = new_n514 & new_n517_1;
  assign new_n519 = ~new_n508 & new_n518;
  assign new_n520 = new_n428_1 & ~new_n519;
  assign new_n521 = n244 & n1239;
  assign new_n522 = n641 & ~n1239;
  assign new_n523 = ~new_n521 & ~new_n522;
  assign new_n524 = ~n293 & ~new_n523;
  assign new_n525 = n293 & new_n523;
  assign new_n526 = ~new_n524 & ~new_n525;
  assign new_n527 = ~new_n520 & new_n526;
  assign new_n528 = n1239 & n1289;
  assign new_n529 = n1193 & ~n1239;
  assign new_n530 = ~new_n528 & ~new_n529;
  assign new_n531 = n920 & new_n530;
  assign new_n532 = ~n920 & ~new_n530;
  assign new_n533 = ~new_n531 & ~new_n532;
  assign new_n534_1 = new_n527 & new_n533;
  assign new_n535 = new_n396_1 & new_n534_1;
  assign new_n536 = ~new_n524 & ~new_n532;
  assign new_n537 = ~new_n531 & ~new_n536;
  assign new_n538 = ~new_n394 & ~new_n537;
  assign new_n539 = ~new_n393 & ~new_n538;
  assign new_n540 = ~new_n388 & new_n539;
  assign new_n541 = ~new_n387 & ~new_n540;
  assign new_n542 = ~new_n535 & new_n541;
  assign new_n543 = new_n383 & ~new_n542;
  assign new_n544 = new_n373 & ~new_n543;
  assign new_n545_1 = new_n342 & ~new_n544;
  assign new_n546 = new_n337_1 & ~new_n545_1;
  assign new_n547 = new_n321 & new_n546;
  assign new_n548 = ~new_n321 & ~new_n546;
  assign n22 = new_n547 | new_n548;
  assign n30 = n1361 | ~n1387;
  assign new_n551 = new_n520 & ~new_n526;
  assign n112 = ~new_n527 & ~new_n551;
  assign new_n553_1 = n1520 & n1613;
  assign new_n554 = n284 & n574;
  assign n126 = ~new_n553_1 | ~new_n554;
  assign new_n556 = n156 & ~n559;
  assign new_n557 = n986 & ~new_n556;
  assign new_n558 = n559 & n589;
  assign new_n559_1 = n156 & ~n986;
  assign new_n560_1 = ~new_n558 & new_n559_1;
  assign new_n561_1 = ~new_n557 & ~new_n560_1;
  assign new_n562 = ~n727 & n1239;
  assign new_n563 = ~new_n316 & ~new_n562;
  assign new_n564 = n40 & ~n1239;
  assign new_n565 = n1239 & ~n1263;
  assign new_n566 = ~new_n564 & ~new_n565;
  assign new_n567_1 = new_n563 & ~new_n566;
  assign new_n568 = ~n94 & n1239;
  assign new_n569 = ~new_n316 & ~new_n568;
  assign new_n570 = n489 & ~n1239;
  assign new_n571 = ~n346 & n1239;
  assign new_n572 = ~new_n570 & ~new_n571;
  assign new_n573 = new_n569 & ~new_n572;
  assign new_n574_1 = ~new_n567_1 & ~new_n573;
  assign new_n575 = ~new_n563 & new_n566;
  assign new_n576 = ~new_n574_1 & ~new_n575;
  assign new_n577 = ~new_n569 & new_n572;
  assign new_n578 = new_n574_1 & ~new_n575;
  assign new_n579 = ~new_n577 & new_n578;
  assign new_n580 = ~n787 & n1239;
  assign new_n581_1 = ~new_n316 & ~new_n580;
  assign new_n582_1 = n1164 & ~n1239;
  assign new_n583 = ~n399 & n1239;
  assign new_n584 = ~new_n582_1 & ~new_n583;
  assign new_n585_1 = new_n581_1 & ~new_n584;
  assign new_n586 = ~n609 & n1239;
  assign new_n587 = ~new_n316 & ~new_n586;
  assign new_n588 = n71 & ~n1239;
  assign new_n589_1 = ~n980 & n1239;
  assign new_n590 = ~new_n588 & ~new_n589_1;
  assign new_n591 = new_n587 & ~new_n590;
  assign new_n592 = ~new_n585_1 & ~new_n591;
  assign new_n593_1 = ~new_n581_1 & new_n584;
  assign new_n594 = ~new_n592 & ~new_n593_1;
  assign new_n595_1 = ~n839 & n1239;
  assign new_n596 = ~new_n316 & ~new_n595_1;
  assign new_n597_1 = ~n1239 & n1523;
  assign new_n598_1 = ~n318 & n1239;
  assign new_n599 = ~new_n597_1 & ~new_n598_1;
  assign new_n600_1 = ~new_n596 & new_n599;
  assign new_n601 = ~new_n587 & new_n590;
  assign new_n602 = new_n592 & ~new_n593_1;
  assign new_n603 = ~new_n601 & new_n602;
  assign new_n604 = n953 & n1239;
  assign new_n605 = ~new_n348 & ~new_n604;
  assign new_n606 = ~n1239 & n1305;
  assign new_n607_1 = n1239 & ~n1592;
  assign new_n608_1 = ~new_n606 & ~new_n607_1;
  assign new_n609_1 = ~new_n605 & ~new_n608_1;
  assign new_n610 = new_n596 & ~new_n599;
  assign new_n611 = ~new_n609_1 & ~new_n610;
  assign new_n612 = n52 & n1239;
  assign new_n613 = ~new_n353 & ~new_n612;
  assign new_n614 = ~n1239 & n1418;
  assign new_n615 = n1239 & ~n1616;
  assign new_n616 = ~new_n614 & ~new_n615;
  assign new_n617 = new_n613 & new_n616;
  assign new_n618 = new_n605 & new_n608_1;
  assign new_n619 = ~new_n617 & ~new_n618;
  assign new_n620 = ~new_n613 & ~new_n616;
  assign new_n621 = n1239 & n1428;
  assign new_n622 = ~new_n358 & ~new_n621;
  assign new_n623 = n1156 & ~n1239;
  assign new_n624 = n1239 & ~n1446;
  assign new_n625_1 = ~new_n623 & ~new_n624;
  assign new_n626_1 = ~new_n622 & ~new_n625_1;
  assign new_n627 = n607 & n1239;
  assign new_n628 = ~new_n362_1 & ~new_n627;
  assign new_n629 = n969 & ~n1239;
  assign new_n630 = n1239 & ~n1345;
  assign new_n631 = ~new_n629 & ~new_n630;
  assign new_n632 = ~new_n628 & ~new_n631;
  assign new_n633 = ~new_n626_1 & ~new_n632;
  assign new_n634 = new_n622 & new_n625_1;
  assign new_n635 = ~new_n633 & ~new_n634;
  assign new_n636 = ~new_n620 & ~new_n635;
  assign new_n637 = new_n619 & ~new_n636;
  assign new_n638_1 = new_n611 & ~new_n637;
  assign new_n639 = new_n603 & ~new_n638_1;
  assign new_n640_1 = ~new_n600_1 & new_n639;
  assign new_n641_1 = ~new_n594 & ~new_n640_1;
  assign new_n642 = new_n579 & ~new_n641_1;
  assign new_n643 = ~new_n576 & ~new_n642;
  assign new_n644 = new_n611 & ~new_n620;
  assign new_n645_1 = ~new_n634 & new_n644;
  assign new_n646 = new_n579 & new_n603;
  assign new_n647 = new_n645_1 & new_n646;
  assign new_n648 = new_n628 & new_n631;
  assign new_n649 = ~new_n600_1 & ~new_n648;
  assign new_n650 = new_n619 & new_n649;
  assign new_n651 = new_n633 & new_n650;
  assign new_n652 = n734 & n1239;
  assign new_n653 = ~new_n398 & ~new_n652;
  assign new_n654 = n1152 & ~n1239;
  assign new_n655 = ~n408 & n1239;
  assign new_n656 = ~new_n654 & ~new_n655;
  assign new_n657 = ~new_n653 & ~new_n656;
  assign new_n658 = new_n653 & new_n656;
  assign new_n659 = ~new_n657 & ~new_n658;
  assign new_n660 = n1239 & n1586;
  assign new_n661 = ~new_n403 & ~new_n660;
  assign new_n662 = ~n1239 & n1386;
  assign new_n663_1 = n1239 & ~n1476;
  assign new_n664 = ~new_n662 & ~new_n663_1;
  assign new_n665 = ~new_n661 & ~new_n664;
  assign new_n666 = n77 & n1239;
  assign new_n667 = ~new_n408_1 & ~new_n666;
  assign new_n668 = n882 & ~n1239;
  assign new_n669_1 = ~n823 & n1239;
  assign new_n670 = ~new_n668 & ~new_n669_1;
  assign new_n671_1 = ~new_n667 & ~new_n670;
  assign new_n672 = n344 & n1239;
  assign new_n673 = ~new_n418 & ~new_n672;
  assign new_n674 = n1227 & ~n1239;
  assign new_n675 = n1239 & ~n1401;
  assign new_n676_1 = ~new_n674 & ~new_n675;
  assign new_n677 = new_n673 & new_n676_1;
  assign new_n678 = ~new_n671_1 & ~new_n677;
  assign new_n679 = ~new_n665 & new_n678;
  assign new_n680 = new_n659 & new_n679;
  assign new_n681 = n273 & n1239;
  assign new_n682 = ~new_n391_1 & ~new_n681;
  assign new_n683 = n507 & ~n1239;
  assign new_n684 = n1239 & ~n1566;
  assign new_n685 = ~new_n683 & ~new_n684;
  assign new_n686 = new_n682 & new_n685;
  assign new_n687 = n376 & n1239;
  assign new_n688 = ~new_n385 & ~new_n687;
  assign new_n689 = n779 & ~n1239;
  assign new_n690_1 = n1239 & ~n1301;
  assign new_n691 = ~new_n689 & ~new_n690_1;
  assign new_n692 = ~new_n688 & ~new_n691;
  assign new_n693_1 = ~new_n682 & ~new_n685;
  assign new_n694 = ~new_n692 & ~new_n693_1;
  assign new_n695_1 = new_n688 & new_n691;
  assign new_n696 = new_n694 & ~new_n695_1;
  assign new_n697 = ~new_n686 & new_n696;
  assign new_n698 = n1114 & n1239;
  assign new_n699 = ~new_n413 & ~new_n698;
  assign new_n700 = ~n1239 & n1627;
  assign new_n701_1 = ~n153 & n1239;
  assign new_n702 = ~new_n700 & ~new_n701_1;
  assign new_n703 = new_n699 & new_n702;
  assign new_n704 = n288 & n1239;
  assign new_n705 = ~new_n436 & ~new_n704;
  assign new_n706 = n936 & ~n1239;
  assign new_n707 = ~n567 & n1239;
  assign new_n708 = ~new_n706 & ~new_n707;
  assign new_n709 = ~new_n705 & ~new_n708;
  assign new_n710_1 = n1239 & n1753;
  assign new_n711 = ~new_n430_1 & ~new_n710_1;
  assign new_n712 = n755 & ~n1239;
  assign new_n713 = ~n374 & n1239;
  assign new_n714_1 = ~new_n712 & ~new_n713;
  assign new_n715 = new_n711 & new_n714_1;
  assign new_n716 = new_n709 & new_n715;
  assign new_n717 = ~new_n703 & ~new_n716;
  assign new_n718 = new_n697 & new_n717;
  assign new_n719_1 = n50 & n1239;
  assign new_n720 = ~new_n522 & ~new_n719_1;
  assign new_n721 = ~n1239 & n1448;
  assign new_n722 = ~n293 & n1239;
  assign new_n723 = ~new_n721 & ~new_n722;
  assign new_n724 = new_n720 & new_n723;
  assign new_n725 = n885 & n1239;
  assign new_n726_1 = ~new_n529 & ~new_n725;
  assign new_n727_1 = n107 & ~n1239;
  assign new_n728 = ~n920 & n1239;
  assign new_n729_1 = ~new_n727_1 & ~new_n728;
  assign new_n730 = ~new_n726_1 & ~new_n729_1;
  assign new_n731 = ~new_n720 & ~new_n723;
  assign new_n732 = ~new_n730 & ~new_n731;
  assign new_n733 = new_n726_1 & new_n729_1;
  assign new_n734_1 = new_n732 & ~new_n733;
  assign new_n735 = ~new_n724 & new_n734_1;
  assign new_n736 = new_n667 & new_n670;
  assign new_n737 = ~new_n699 & ~new_n702;
  assign new_n738 = ~new_n673 & ~new_n676_1;
  assign new_n739 = ~new_n737 & ~new_n738;
  assign new_n740 = new_n661 & new_n664;
  assign new_n741 = new_n739 & ~new_n740;
  assign new_n742_1 = ~new_n736 & new_n741;
  assign new_n743_1 = new_n735 & new_n742_1;
  assign new_n744 = new_n718 & new_n743_1;
  assign new_n745 = new_n705 & new_n708;
  assign new_n746 = n416 & n1239;
  assign new_n747 = ~new_n443 & ~new_n746;
  assign new_n748 = n159 & ~n1239;
  assign new_n749 = n1239 & ~n1463;
  assign new_n750 = ~new_n748 & ~new_n749;
  assign new_n751 = new_n747 & new_n750;
  assign new_n752 = ~new_n715 & ~new_n751;
  assign new_n753 = ~new_n745 & new_n752;
  assign new_n754 = n506 & n1239;
  assign new_n755_1 = ~new_n449 & ~new_n754;
  assign new_n756 = n243 & ~n1239;
  assign new_n757 = ~n222 & n1239;
  assign new_n758 = ~new_n756 & ~new_n757;
  assign new_n759 = new_n755_1 & new_n758;
  assign new_n760 = n392 & n1239;
  assign new_n761 = ~new_n455 & ~new_n760;
  assign new_n762 = n742 & ~n1239;
  assign new_n763 = ~n608 & n1239;
  assign new_n764 = ~new_n762 & ~new_n763;
  assign new_n765 = ~new_n761 & ~new_n764;
  assign new_n766 = n671 & n1239;
  assign new_n767 = ~new_n461 & ~new_n766;
  assign new_n768 = n341 & ~n1239;
  assign new_n769_1 = ~n1071 & n1239;
  assign new_n770 = ~new_n768 & ~new_n769_1;
  assign new_n771 = new_n767 & new_n770;
  assign new_n772 = n778 & n1239;
  assign new_n773_1 = ~new_n474 & ~new_n772;
  assign new_n774 = n502 & ~n1239;
  assign new_n775_1 = ~n695 & n1239;
  assign new_n776 = ~new_n774 & ~new_n775_1;
  assign new_n777 = ~new_n773_1 & ~new_n776;
  assign new_n778_1 = ~n729 & new_n489_1;
  assign new_n779_1 = n690 & ~new_n778_1;
  assign new_n780 = n729 & new_n477_1;
  assign new_n781 = ~new_n779_1 & ~new_n780;
  assign new_n782_1 = ~new_n777 & new_n781;
  assign new_n783 = n29 & n1239;
  assign new_n784 = ~new_n468 & ~new_n783;
  assign new_n785 = n849 & ~n1239;
  assign new_n786 = ~n45 & n1239;
  assign new_n787_1 = ~new_n785 & ~new_n786;
  assign new_n788 = new_n784 & new_n787_1;
  assign new_n789 = new_n773_1 & new_n776;
  assign new_n790_1 = ~new_n788 & ~new_n789;
  assign new_n791 = ~new_n782_1 & new_n790_1;
  assign new_n792 = ~new_n767 & ~new_n770;
  assign new_n793 = ~new_n784 & ~new_n787_1;
  assign new_n794_1 = ~new_n792 & ~new_n793;
  assign new_n795 = ~new_n791 & new_n794_1;
  assign new_n796 = ~new_n771 & ~new_n795;
  assign new_n797 = ~new_n765 & ~new_n796;
  assign new_n798 = new_n761 & new_n764;
  assign new_n799 = ~new_n797 & ~new_n798;
  assign new_n800 = ~new_n759 & new_n799;
  assign new_n801 = ~new_n755_1 & ~new_n758;
  assign new_n802 = ~new_n747 & ~new_n750;
  assign new_n803 = ~new_n801 & ~new_n802;
  assign new_n804 = ~new_n800 & new_n803;
  assign new_n805 = new_n753 & ~new_n804;
  assign new_n806 = ~new_n711 & ~new_n714_1;
  assign new_n807 = ~new_n709 & ~new_n806;
  assign new_n808 = ~new_n805 & new_n807;
  assign new_n809 = new_n744 & ~new_n808;
  assign new_n810 = new_n680 & new_n809;
  assign new_n811 = ~new_n694 & ~new_n695_1;
  assign new_n812 = ~new_n732 & ~new_n733;
  assign new_n813 = ~new_n703 & ~new_n739;
  assign new_n814 = ~new_n671_1 & ~new_n813;
  assign new_n815 = ~new_n736 & ~new_n814;
  assign new_n816 = ~new_n740 & new_n815;
  assign new_n817 = ~new_n657 & ~new_n665;
  assign new_n818 = ~new_n816 & new_n817;
  assign new_n819 = ~new_n658 & new_n735;
  assign new_n820 = ~new_n818 & new_n819;
  assign new_n821_1 = ~new_n812 & ~new_n820;
  assign new_n822 = new_n697 & ~new_n821_1;
  assign new_n823_1 = ~new_n811 & ~new_n822;
  assign n1306 = new_n810 | ~new_n823_1;
  assign new_n825 = new_n651 & n1306;
  assign new_n826 = new_n647 & new_n825;
  assign new_n827 = new_n643 & ~new_n826;
  assign new_n828 = n1239 & ~n1299;
  assign new_n829 = ~new_n316 & ~new_n828;
  assign new_n830 = n879 & ~n1239;
  assign new_n831_1 = ~n769 & n1239;
  assign new_n832_1 = ~new_n830 & ~new_n831_1;
  assign new_n833 = new_n829 & ~new_n832_1;
  assign new_n834 = ~n86 & n1239;
  assign new_n835 = ~new_n316 & ~new_n834;
  assign new_n836 = n561 & ~n1239;
  assign new_n837 = ~n138 & n1239;
  assign new_n838 = ~new_n836 & ~new_n837;
  assign new_n839_1 = new_n835 & ~new_n838;
  assign new_n840 = ~new_n833 & ~new_n839_1;
  assign new_n841 = n1239 & ~n1502;
  assign new_n842_1 = ~new_n316 & ~new_n841;
  assign new_n843 = n143 & ~n1239;
  assign new_n844 = ~n626 & n1239;
  assign new_n845 = ~new_n843 & ~new_n844;
  assign new_n846 = new_n842_1 & new_n845;
  assign new_n847 = ~new_n842_1 & ~new_n845;
  assign new_n848 = ~new_n846 & ~new_n847;
  assign new_n849_1 = new_n840 & ~new_n848;
  assign new_n850 = ~new_n829 & new_n832_1;
  assign new_n851 = ~n223 & n1239;
  assign new_n852 = ~new_n316 & ~new_n851;
  assign new_n853 = n300 & ~n1239;
  assign new_n854 = n1239 & ~n1470;
  assign new_n855 = ~new_n853 & ~new_n854;
  assign new_n856 = ~new_n852 & new_n855;
  assign new_n857 = ~new_n835 & new_n838;
  assign new_n858 = ~new_n856 & ~new_n857;
  assign new_n859 = new_n852 & ~new_n855;
  assign new_n860 = n663 & ~n1239;
  assign new_n861 = n1239 & ~n1656;
  assign new_n862 = ~new_n860 & ~new_n861;
  assign new_n863 = new_n316 & new_n862;
  assign new_n864 = ~new_n859 & ~new_n863;
  assign new_n865 = ~new_n316 & ~new_n862;
  assign new_n866 = new_n864 & ~new_n865;
  assign new_n867 = new_n858 & new_n866;
  assign new_n868 = ~new_n850 & new_n867;
  assign new_n869 = new_n849_1 & new_n868;
  assign new_n870 = ~new_n827 & new_n869;
  assign new_n871 = ~n1656 & ~new_n845;
  assign new_n872 = new_n841 & ~new_n871;
  assign new_n873 = new_n845 & new_n862;
  assign new_n874 = ~new_n850 & ~new_n873;
  assign new_n875 = ~new_n316 & new_n874;
  assign new_n876 = ~new_n872 & new_n875;
  assign new_n877 = new_n840 & ~new_n876;
  assign new_n878 = new_n858 & ~new_n877;
  assign new_n879_1 = ~new_n859 & ~new_n878;
  assign new_n880 = ~new_n870 & new_n879_1;
  assign new_n881 = new_n561_1 & ~new_n880;
  assign new_n882_1 = n589 & n986;
  assign new_n883 = ~new_n557 & ~new_n882_1;
  assign n161 = new_n881 | ~new_n883;
  assign new_n885_1 = new_n370_1 & ~new_n379;
  assign new_n886 = ~new_n350 & ~new_n885_1;
  assign new_n887 = new_n370_1 & new_n542;
  assign new_n888 = new_n886 & ~new_n887;
  assign new_n889 = ~new_n380_1 & new_n888;
  assign new_n890 = new_n380_1 & ~new_n888;
  assign n164 = new_n889 | new_n890;
  assign new_n892 = ~new_n333 & ~new_n338;
  assign new_n893 = ~new_n544 & ~new_n892;
  assign new_n894_1 = new_n544 & new_n892;
  assign n181 = new_n893 | new_n894_1;
  assign new_n896 = ~n477 & n1239;
  assign new_n897 = ~new_n316 & ~new_n896;
  assign new_n898 = n769 & ~new_n897;
  assign new_n899 = ~n769 & new_n897;
  assign new_n900 = ~new_n898 & ~new_n899;
  assign new_n901 = ~n1191 & n1239;
  assign new_n902 = ~new_n316 & ~new_n901;
  assign new_n903 = ~n626 & new_n902;
  assign new_n904 = n626 & ~new_n902;
  assign new_n905_1 = ~new_n903 & ~new_n904;
  assign new_n906 = ~n430 & n1239;
  assign new_n907 = ~new_n316 & ~new_n906;
  assign new_n908 = ~n1656 & new_n907;
  assign new_n909 = n1656 & ~new_n907;
  assign new_n910 = ~new_n908 & ~new_n909;
  assign new_n911 = ~new_n324 & ~new_n328;
  assign new_n912 = new_n321 & ~new_n325;
  assign new_n913 = ~new_n911 & new_n912;
  assign new_n914 = ~new_n324 & new_n912;
  assign new_n915 = new_n340 & ~new_n544;
  assign new_n916_1 = ~new_n334 & ~new_n915;
  assign new_n917 = new_n914 & ~new_n916_1;
  assign new_n918_1 = ~new_n913 & ~new_n917;
  assign new_n919 = ~new_n319 & new_n918_1;
  assign new_n920_1 = new_n910 & ~new_n919;
  assign new_n921 = ~new_n908 & ~new_n920_1;
  assign new_n922 = new_n905_1 & ~new_n921;
  assign new_n923 = ~new_n903 & ~new_n922;
  assign new_n924 = new_n900 & new_n923;
  assign new_n925 = ~new_n900 & ~new_n923;
  assign n216 = new_n924 | new_n925;
  assign new_n927 = new_n447 & ~new_n452;
  assign new_n928 = new_n440 & ~new_n451;
  assign new_n929 = new_n927 & new_n928;
  assign new_n930 = new_n505 & ~new_n929;
  assign new_n931 = ~new_n447 & ~new_n451;
  assign new_n932 = ~new_n927 & ~new_n931;
  assign new_n933 = ~new_n434 & ~new_n440;
  assign new_n934 = ~new_n441 & ~new_n933;
  assign new_n935 = new_n503 & ~new_n934;
  assign new_n936_1 = ~new_n503 & new_n934;
  assign new_n937 = ~new_n935 & ~new_n936_1;
  assign new_n938 = ~new_n932 & new_n937;
  assign new_n939 = new_n932 & ~new_n937;
  assign new_n940 = ~new_n938 & ~new_n939;
  assign new_n941 = new_n930 & new_n940;
  assign new_n942 = ~new_n930 & ~new_n940;
  assign new_n943 = ~new_n941 & ~new_n942;
  assign new_n944 = ~new_n488 & new_n943;
  assign new_n945 = ~new_n447 & new_n452;
  assign new_n946 = ~new_n927 & ~new_n945;
  assign new_n947_1 = new_n505 & ~new_n946;
  assign new_n948 = ~new_n505 & new_n946;
  assign new_n949 = ~new_n947_1 & ~new_n948;
  assign new_n950 = ~new_n937 & new_n949;
  assign new_n951 = new_n937 & ~new_n949;
  assign new_n952_1 = new_n488 & ~new_n951;
  assign new_n953_1 = ~new_n950 & new_n952_1;
  assign new_n954 = ~n545 & ~new_n953_1;
  assign new_n955 = ~new_n944 & new_n954;
  assign new_n956 = new_n488 & ~new_n496;
  assign new_n957 = new_n943 & ~new_n956;
  assign new_n958 = ~new_n496 & new_n953_1;
  assign new_n959 = n545 & ~new_n958;
  assign new_n960 = ~new_n957 & new_n959;
  assign new_n961_1 = ~new_n955 & ~new_n960;
  assign new_n962 = ~new_n459 & ~new_n465;
  assign new_n963 = ~new_n466 & ~new_n962;
  assign new_n964 = ~new_n476 & new_n490;
  assign new_n965 = ~new_n479 & ~new_n964;
  assign new_n966 = ~new_n491 & new_n965;
  assign new_n967 = new_n491 & ~new_n965;
  assign new_n968 = ~new_n966 & ~new_n967;
  assign new_n969_1 = ~new_n963 & ~new_n968;
  assign new_n970 = new_n963 & new_n968;
  assign new_n971 = ~new_n969_1 & ~new_n970;
  assign new_n972 = ~new_n471 & ~new_n482;
  assign new_n973 = new_n490 & ~new_n972;
  assign new_n974 = ~new_n490 & ~new_n494;
  assign new_n975 = new_n972 & new_n974;
  assign new_n976 = ~new_n973 & ~new_n975;
  assign new_n977 = ~new_n971 & new_n976;
  assign new_n978 = new_n971 & ~new_n976;
  assign new_n979 = ~new_n977 & ~new_n978;
  assign new_n980_1 = ~new_n472 & ~new_n492;
  assign new_n981 = ~new_n493 & ~new_n980_1;
  assign new_n982 = ~new_n482 & new_n484;
  assign new_n983 = ~new_n463 & ~new_n982;
  assign new_n984_1 = ~new_n495 & ~new_n983;
  assign new_n985 = new_n981 & new_n984_1;
  assign new_n986_1 = ~new_n981 & ~new_n984_1;
  assign new_n987 = ~new_n985 & ~new_n986_1;
  assign new_n988 = ~new_n979 & new_n987;
  assign new_n989 = new_n979 & ~new_n987;
  assign new_n990_1 = ~new_n988 & ~new_n989;
  assign new_n991 = n545 & new_n990_1;
  assign new_n992_1 = new_n478_1 & ~new_n963;
  assign new_n993 = ~new_n478_1 & new_n963;
  assign new_n994 = ~new_n992_1 & ~new_n993;
  assign new_n995 = new_n470 & ~new_n481;
  assign new_n996 = new_n471 & new_n481;
  assign new_n997_1 = ~new_n995 & ~new_n996;
  assign new_n998 = new_n994 & new_n997_1;
  assign new_n999 = ~new_n994 & ~new_n997_1;
  assign new_n1000 = ~new_n998 & ~new_n999;
  assign new_n1001 = new_n491 & new_n981;
  assign new_n1002 = ~new_n491 & ~new_n981;
  assign new_n1003 = ~new_n1001 & ~new_n1002;
  assign new_n1004 = new_n983 & new_n1003;
  assign new_n1005 = ~new_n983 & ~new_n1003;
  assign new_n1006_1 = ~new_n1004 & ~new_n1005;
  assign new_n1007 = new_n1000 & new_n1006_1;
  assign new_n1008 = ~new_n1000 & ~new_n1006_1;
  assign new_n1009 = ~new_n1007 & ~new_n1008;
  assign new_n1010 = ~n545 & new_n1009;
  assign new_n1011 = ~new_n991 & ~new_n1010;
  assign new_n1012 = ~new_n961_1 & new_n1011;
  assign new_n1013 = new_n961_1 & ~new_n1011;
  assign n233 = ~new_n1012 & ~new_n1013;
  assign new_n1015 = ~new_n508 & new_n510_1;
  assign new_n1016 = ~new_n420_1 & ~new_n1015;
  assign new_n1017_1 = new_n512 & ~new_n1016;
  assign new_n1018 = ~new_n415 & ~new_n1017_1;
  assign new_n1019 = new_n511 & ~new_n1018;
  assign new_n1020 = ~new_n410 & ~new_n1019;
  assign new_n1021 = ~new_n516_1 & new_n1020;
  assign new_n1022 = new_n516_1 & ~new_n1020;
  assign n247 = ~new_n1021 & ~new_n1022;
  assign n304 = n420 & n832;
  assign new_n1025 = new_n335 & ~new_n915;
  assign new_n1026 = new_n341_1 & ~new_n1025;
  assign new_n1027 = ~new_n341_1 & new_n1025;
  assign n364 = ~new_n1026 & ~new_n1027;
  assign new_n1029 = new_n425 & new_n508;
  assign new_n1030 = ~new_n405 & new_n514;
  assign new_n1031 = ~new_n426 & ~new_n1030;
  assign new_n1032 = ~new_n1029 & ~new_n1031;
  assign new_n1033 = ~new_n515 & new_n1032;
  assign new_n1034 = new_n515 & ~new_n1032;
  assign n370 = new_n1033 | new_n1034;
  assign new_n1036 = n1239 & ~n1500;
  assign new_n1037 = ~new_n316 & ~new_n1036;
  assign new_n1038 = n138 & ~new_n1037;
  assign new_n1039 = new_n900 & new_n905_1;
  assign new_n1040_1 = ~new_n899 & ~new_n903;
  assign new_n1041 = ~new_n898 & ~new_n1040_1;
  assign new_n1042_1 = ~new_n1039 & ~new_n1041;
  assign new_n1043 = new_n910 & ~new_n1042_1;
  assign new_n1044_1 = ~n138 & new_n1037;
  assign new_n1045 = ~new_n908 & ~new_n1041;
  assign new_n1046 = ~new_n1042_1 & ~new_n1045;
  assign new_n1047 = ~new_n1044_1 & ~new_n1046;
  assign new_n1048 = ~new_n1043 & new_n1047;
  assign new_n1049 = ~new_n1038 & ~new_n1048;
  assign new_n1050_1 = ~new_n900 & ~new_n905_1;
  assign new_n1051_1 = ~new_n1039 & ~new_n1050_1;
  assign new_n1052 = ~new_n905_1 & new_n910;
  assign new_n1053 = new_n905_1 & new_n908;
  assign new_n1054_1 = ~new_n903 & ~new_n1053;
  assign new_n1055 = ~n582 & n1239;
  assign new_n1056 = ~new_n316 & ~new_n1055;
  assign new_n1057 = ~n1470 & new_n1056;
  assign new_n1058_1 = n1470 & ~new_n1056;
  assign new_n1059 = ~new_n1057 & ~new_n1058_1;
  assign new_n1060_1 = ~new_n1038 & ~new_n1044_1;
  assign new_n1061_1 = new_n1059 & new_n1060_1;
  assign new_n1062 = ~new_n1059 & ~new_n1060_1;
  assign new_n1063_1 = ~new_n1061_1 & ~new_n1062;
  assign new_n1064 = ~new_n1054_1 & new_n1063_1;
  assign new_n1065_1 = new_n1054_1 & ~new_n1063_1;
  assign new_n1066 = ~new_n1064 & ~new_n1065_1;
  assign new_n1067 = new_n909 & ~new_n1041;
  assign new_n1068 = ~new_n909 & ~new_n1042_1;
  assign new_n1069 = ~new_n1067 & ~new_n1068;
  assign new_n1070 = ~new_n1066 & new_n1069;
  assign new_n1071_1 = new_n1066 & ~new_n1069;
  assign new_n1072 = ~new_n1070 & ~new_n1071_1;
  assign new_n1073 = new_n1052 & new_n1072;
  assign new_n1074 = ~new_n1052 & ~new_n1072;
  assign new_n1075 = ~new_n1073 & ~new_n1074;
  assign new_n1076 = new_n1051_1 & new_n1075;
  assign new_n1077 = ~new_n1051_1 & ~new_n1075;
  assign new_n1078 = ~new_n1076 & ~new_n1077;
  assign new_n1079 = new_n1049 & ~new_n1078;
  assign new_n1080 = ~new_n1049 & new_n1078;
  assign new_n1081 = ~new_n1079 & ~new_n1080;
  assign new_n1082 = ~new_n919 & new_n1081;
  assign new_n1083 = ~new_n910 & ~new_n1051_1;
  assign new_n1084 = new_n910 & new_n1051_1;
  assign new_n1085 = ~new_n1083 & ~new_n1084;
  assign new_n1086 = new_n908 & ~new_n1042_1;
  assign new_n1087 = ~new_n1045 & ~new_n1086;
  assign new_n1088 = ~new_n1038 & ~new_n1047;
  assign new_n1089 = new_n1087 & new_n1088;
  assign new_n1090 = ~new_n1087 & ~new_n1088;
  assign new_n1091 = ~new_n1089 & ~new_n1090;
  assign new_n1092 = new_n1066 & new_n1091;
  assign new_n1093 = ~new_n1066 & ~new_n1091;
  assign new_n1094 = ~new_n1092 & ~new_n1093;
  assign new_n1095_1 = new_n1085 & ~new_n1094;
  assign new_n1096 = ~new_n1085 & new_n1094;
  assign new_n1097 = ~new_n1095_1 & ~new_n1096;
  assign new_n1098 = new_n919 & new_n1097;
  assign new_n1099 = ~new_n1082 & ~new_n1098;
  assign new_n1100 = ~new_n920_1 & new_n1045;
  assign new_n1101 = ~new_n1042_1 & ~new_n1100;
  assign new_n1102 = new_n1060_1 & new_n1101;
  assign new_n1103_1 = ~new_n1044_1 & ~new_n1057;
  assign new_n1104 = ~new_n1102 & new_n1103_1;
  assign new_n1105 = ~new_n1058_1 & ~new_n1104;
  assign new_n1106 = n156 & n200;
  assign new_n1107 = n986 & new_n1106;
  assign new_n1108 = ~n487 & new_n1107;
  assign new_n1109 = n156 & n487;
  assign new_n1110 = ~new_n1107 & new_n1109;
  assign new_n1111 = ~new_n1108 & ~new_n1110;
  assign new_n1112 = new_n1105 & ~new_n1111;
  assign new_n1113 = ~n986 & ~new_n1106;
  assign new_n1114_1 = new_n1109 & new_n1113;
  assign new_n1115 = ~new_n1109 & ~new_n1113;
  assign new_n1116 = ~new_n1114_1 & ~new_n1115;
  assign new_n1117 = ~new_n1105 & ~new_n1116;
  assign new_n1118 = ~new_n1112 & ~new_n1117;
  assign new_n1119 = ~new_n1099 & new_n1118;
  assign new_n1120 = new_n1099 & ~new_n1118;
  assign n378 = new_n1119 | new_n1120;
  assign new_n1122 = ~new_n338 & ~new_n544;
  assign new_n1123 = ~new_n333 & ~new_n1122;
  assign new_n1124 = ~new_n330 & new_n1123;
  assign new_n1125 = new_n330 & ~new_n1123;
  assign n396 = ~new_n1124 & ~new_n1125;
  assign new_n1127 = ~new_n1105 & ~new_n1111;
  assign new_n1128 = new_n1105 & new_n1116;
  assign n428 = ~new_n1127 & ~new_n1128;
  assign new_n1130 = ~new_n1107 & ~new_n1113;
  assign new_n1131 = new_n1105 & ~new_n1130;
  assign new_n1132 = ~new_n1105 & new_n1130;
  assign n453 = ~new_n1131 & ~new_n1132;
  assign new_n1134 = new_n526 & new_n533;
  assign new_n1135 = new_n538 & ~new_n1134;
  assign new_n1136 = ~new_n393 & ~new_n1135;
  assign new_n1137 = new_n520 & new_n538;
  assign new_n1138_1 = new_n1136 & ~new_n1137;
  assign new_n1139 = ~new_n389 & new_n1138_1;
  assign new_n1140 = new_n389 & ~new_n1138_1;
  assign n517 = new_n1139 | new_n1140;
  assign new_n1142 = new_n375 & ~new_n542;
  assign new_n1143 = ~new_n364_1 & ~new_n1142;
  assign new_n1144 = new_n377 & ~new_n1143;
  assign new_n1145 = ~new_n360 & ~new_n1144;
  assign new_n1146 = ~new_n376_1 & new_n1145;
  assign new_n1147 = new_n376_1 & ~new_n1145;
  assign n534 = ~new_n1146 & ~new_n1147;
  assign new_n1149 = n487 & new_n1106;
  assign new_n1150 = n986 & ~new_n1149;
  assign new_n1151 = ~n200 & ~n487;
  assign new_n1152_1 = new_n559_1 & ~new_n1151;
  assign new_n1153 = new_n1105 & ~new_n1152_1;
  assign n553 = new_n1150 | new_n1153;
  assign new_n1155 = n545 & new_n491;
  assign new_n1156_1 = ~n545 & ~new_n491;
  assign n597 = ~new_n1155 & ~new_n1156_1;
  assign new_n1158 = ~new_n537 & ~new_n1134;
  assign new_n1159 = ~new_n389 & ~new_n395;
  assign new_n1160 = ~new_n396_1 & ~new_n1159;
  assign new_n1161 = ~new_n524 & ~new_n533;
  assign new_n1162 = new_n524 & new_n533;
  assign new_n1163 = ~new_n1161 & ~new_n1162;
  assign new_n1164_1 = new_n1160 & new_n1163;
  assign new_n1165 = ~new_n1160 & ~new_n1163;
  assign new_n1166 = ~new_n1164_1 & ~new_n1165;
  assign new_n1167 = new_n1136 & new_n1166;
  assign new_n1168 = ~new_n1136 & ~new_n1166;
  assign new_n1169 = ~new_n1167 & ~new_n1168;
  assign new_n1170 = new_n1158 & ~new_n1169;
  assign new_n1171 = ~new_n1158 & new_n1169;
  assign new_n1172_1 = ~new_n1170 & ~new_n1171;
  assign new_n1173 = ~new_n520 & ~new_n1172_1;
  assign new_n1174 = new_n524 & ~new_n532;
  assign new_n1175_1 = ~new_n525 & new_n531;
  assign new_n1176 = new_n525 & ~new_n531;
  assign new_n1177_1 = ~new_n1175_1 & ~new_n1176;
  assign new_n1178 = ~new_n1174 & new_n1177_1;
  assign new_n1179 = ~new_n1160 & new_n1178;
  assign new_n1180 = new_n1160 & ~new_n1178;
  assign new_n1181 = ~new_n1179 & ~new_n1180;
  assign new_n1182 = ~new_n539 & new_n1181;
  assign new_n1183 = new_n539 & ~new_n1181;
  assign new_n1184 = ~new_n1182 & ~new_n1183;
  assign new_n1185 = new_n520 & ~new_n1184;
  assign new_n1186_1 = ~new_n1173 & ~new_n1185;
  assign new_n1187_1 = new_n426 & new_n510_1;
  assign new_n1188 = ~new_n426 & ~new_n510_1;
  assign new_n1189 = ~new_n1187_1 & ~new_n1188;
  assign new_n1190 = ~new_n511 & ~new_n512;
  assign new_n1191_1 = ~new_n513 & ~new_n1190;
  assign new_n1192 = ~new_n415 & ~new_n420_1;
  assign new_n1193_1 = ~new_n421 & ~new_n1192;
  assign new_n1194 = ~new_n1191_1 & new_n1193_1;
  assign new_n1195_1 = new_n1191_1 & ~new_n1193_1;
  assign new_n1196 = ~new_n1194 & ~new_n1195_1;
  assign new_n1197 = ~new_n515 & ~new_n516_1;
  assign new_n1198 = ~new_n517_1 & ~new_n1197;
  assign new_n1199 = new_n424 & new_n1198;
  assign new_n1200 = ~new_n424 & ~new_n1198;
  assign new_n1201 = ~new_n1199 & ~new_n1200;
  assign new_n1202 = ~new_n1196 & new_n1201;
  assign new_n1203 = new_n1196 & ~new_n1201;
  assign new_n1204 = ~new_n1202 & ~new_n1203;
  assign new_n1205_1 = ~new_n1189 & new_n1204;
  assign new_n1206 = new_n1189 & ~new_n1204;
  assign new_n1207 = ~new_n1205_1 & ~new_n1206;
  assign new_n1208 = new_n508 & ~new_n1207;
  assign new_n1209_1 = ~new_n1030 & new_n1189;
  assign new_n1210 = ~new_n509_1 & ~new_n514;
  assign new_n1211_1 = new_n424 & new_n1210;
  assign new_n1212 = ~new_n424 & new_n509_1;
  assign new_n1213 = ~new_n1211_1 & ~new_n1212;
  assign new_n1214 = ~new_n1191_1 & ~new_n1198;
  assign new_n1215 = new_n1191_1 & new_n1198;
  assign new_n1216 = ~new_n1214 & ~new_n1215;
  assign new_n1217 = ~new_n415 & new_n509_1;
  assign new_n1218 = ~new_n416_1 & ~new_n1217;
  assign new_n1219 = ~new_n1216 & new_n1218;
  assign new_n1220 = new_n1216 & ~new_n1218;
  assign new_n1221 = ~new_n1219 & ~new_n1220;
  assign new_n1222 = ~new_n1213 & new_n1221;
  assign new_n1223 = new_n1213 & ~new_n1221;
  assign new_n1224 = ~new_n1222 & ~new_n1223;
  assign new_n1225_1 = new_n1209_1 & new_n1224;
  assign new_n1226 = ~new_n1209_1 & ~new_n1224;
  assign new_n1227_1 = ~new_n1225_1 & ~new_n1226;
  assign new_n1228 = ~new_n508 & ~new_n1227_1;
  assign new_n1229 = ~new_n1208 & ~new_n1228;
  assign new_n1230 = new_n1186_1 & ~new_n1229;
  assign new_n1231_1 = ~new_n1186_1 & new_n1229;
  assign n625 = new_n1230 | new_n1231_1;
  assign new_n1233 = n1438 & n1536;
  assign new_n1234_1 = n315 & n997;
  assign n669 = ~new_n1233 | ~new_n1234_1;
  assign new_n1236 = ~new_n512 & new_n1016;
  assign n693 = ~new_n1017_1 & ~new_n1236;
  assign new_n1238 = new_n498_1 & new_n505;
  assign new_n1239_1 = ~new_n930 & ~new_n1238;
  assign new_n1240 = ~new_n434 & new_n1239_1;
  assign new_n1241 = new_n434 & ~new_n1239_1;
  assign n714 = new_n1240 | new_n1241;
  assign n719 = n1225 | n1361;
  assign new_n1244 = ~new_n478_1 & ~new_n1155;
  assign new_n1245 = new_n492 & ~new_n1244;
  assign new_n1246_1 = ~new_n476 & ~new_n1245;
  assign new_n1247 = ~new_n472 & new_n1246_1;
  assign new_n1248 = new_n472 & ~new_n1246_1;
  assign n794 = ~new_n1247 & ~new_n1248;
  assign new_n1250_1 = ~new_n355 & ~new_n1147;
  assign new_n1251 = ~new_n381 & new_n1250_1;
  assign new_n1252 = new_n381 & ~new_n1250_1;
  assign n894 = ~new_n1251 & ~new_n1252;
  assign new_n1254 = ~new_n910 & new_n919;
  assign n916 = ~new_n920_1 & ~new_n1254;
  assign new_n1256 = n1239 & ~new_n316;
  assign new_n1257 = n246 & ~n1389;
  assign new_n1258 = ~n246 & n1389;
  assign new_n1259 = ~new_n1257 & ~new_n1258;
  assign new_n1260 = n56 & new_n1259;
  assign new_n1261 = ~n56 & ~new_n1259;
  assign new_n1262 = ~new_n1260 & ~new_n1261;
  assign new_n1263_1 = new_n1256 & new_n1262;
  assign new_n1264 = new_n828 & new_n842_1;
  assign new_n1265 = new_n829 & new_n841;
  assign new_n1266 = ~new_n1264 & ~new_n1265;
  assign new_n1267 = ~new_n835 & new_n852;
  assign new_n1268 = new_n835 & new_n851;
  assign new_n1269 = ~new_n1267 & ~new_n1268;
  assign new_n1270 = ~new_n1266 & new_n1269;
  assign new_n1271 = new_n1266 & ~new_n1269;
  assign new_n1272 = ~new_n1270 & ~new_n1271;
  assign new_n1273 = ~new_n1263_1 & new_n1272;
  assign new_n1274 = new_n1263_1 & ~new_n1272;
  assign new_n1275 = ~new_n1273 & ~new_n1274;
  assign new_n1276 = new_n673 & ~new_n699;
  assign new_n1277 = ~new_n673 & new_n699;
  assign new_n1278_1 = ~new_n1276 & ~new_n1277;
  assign new_n1279 = new_n661 & new_n1278_1;
  assign new_n1280 = ~new_n661 & ~new_n1278_1;
  assign new_n1281_1 = ~new_n1279 & ~new_n1280;
  assign new_n1282 = new_n653 & new_n682;
  assign new_n1283_1 = ~new_n653 & ~new_n682;
  assign new_n1284 = ~new_n1282 & ~new_n1283_1;
  assign new_n1285_1 = n1121 & ~n1239;
  assign new_n1286_1 = n560 & n1239;
  assign new_n1287 = ~new_n1285_1 & ~new_n1286_1;
  assign new_n1288_1 = ~new_n667 & new_n1287;
  assign new_n1289_1 = new_n667 & ~new_n1287;
  assign new_n1290 = ~new_n1288_1 & ~new_n1289_1;
  assign new_n1291 = ~new_n1284 & new_n1290;
  assign new_n1292_1 = new_n1284 & ~new_n1290;
  assign new_n1293 = ~new_n1291 & ~new_n1292_1;
  assign new_n1294 = new_n688 & new_n726_1;
  assign new_n1295 = ~new_n688 & ~new_n726_1;
  assign new_n1296_1 = ~new_n1294 & ~new_n1295;
  assign new_n1297 = new_n720 & new_n1296_1;
  assign new_n1298 = ~new_n720 & ~new_n1296_1;
  assign new_n1299_1 = ~new_n1297 & ~new_n1298;
  assign new_n1300 = new_n1293 & ~new_n1299_1;
  assign new_n1301_1 = ~new_n1293 & new_n1299_1;
  assign new_n1302_1 = ~new_n1300 & ~new_n1301_1;
  assign new_n1303 = ~new_n1281_1 & new_n1302_1;
  assign new_n1304 = new_n1281_1 & ~new_n1302_1;
  assign new_n1305_1 = ~new_n1303 & ~new_n1304;
  assign new_n1306_1 = ~new_n1275 & ~new_n1305_1;
  assign new_n1307 = n299 & ~n1239;
  assign new_n1308 = n1044 & n1239;
  assign new_n1309 = ~new_n1307 & ~new_n1308;
  assign new_n1310 = new_n784 & ~new_n1309;
  assign new_n1311 = ~new_n784 & new_n1309;
  assign new_n1312 = ~new_n1310 & ~new_n1311;
  assign new_n1313 = new_n711 & new_n755_1;
  assign new_n1314 = ~new_n711 & ~new_n755_1;
  assign new_n1315 = ~new_n1313 & ~new_n1314;
  assign new_n1316 = new_n1312 & ~new_n1315;
  assign new_n1317 = ~new_n1312 & new_n1315;
  assign new_n1318 = ~new_n1316 & ~new_n1317;
  assign new_n1319 = n1239 & ~n1411;
  assign new_n1320_1 = ~new_n489_1 & ~new_n1319;
  assign new_n1321 = ~new_n773_1 & new_n1320_1;
  assign new_n1322_1 = new_n773_1 & ~new_n1320_1;
  assign new_n1323 = ~new_n1321 & ~new_n1322_1;
  assign new_n1324 = new_n705 & new_n747;
  assign new_n1325 = ~new_n705 & ~new_n747;
  assign new_n1326 = ~new_n1324 & ~new_n1325;
  assign new_n1327 = new_n1323 & ~new_n1326;
  assign new_n1328 = ~new_n1323 & new_n1326;
  assign new_n1329 = ~new_n1327 & ~new_n1328;
  assign new_n1330 = new_n761 & new_n767;
  assign new_n1331 = ~new_n761 & ~new_n767;
  assign new_n1332 = ~new_n1330 & ~new_n1331;
  assign new_n1333 = new_n1329 & ~new_n1332;
  assign new_n1334 = ~new_n1329 & new_n1332;
  assign new_n1335 = ~new_n1333 & ~new_n1334;
  assign new_n1336 = ~new_n1318 & ~new_n1335;
  assign new_n1337_1 = new_n1318 & new_n1335;
  assign new_n1338 = ~new_n1336 & ~new_n1337_1;
  assign new_n1339 = new_n581_1 & new_n586;
  assign new_n1340 = new_n580 & new_n587;
  assign new_n1341 = ~new_n1339 & ~new_n1340;
  assign new_n1342 = new_n596 & new_n1341;
  assign new_n1343 = ~new_n596 & ~new_n1341;
  assign new_n1344 = ~new_n1342 & ~new_n1343;
  assign new_n1345_1 = new_n562 & new_n569;
  assign new_n1346_1 = new_n563 & new_n568;
  assign new_n1347 = ~new_n1345_1 & ~new_n1346_1;
  assign new_n1348 = new_n622 & new_n628;
  assign new_n1349 = ~new_n622 & ~new_n628;
  assign new_n1350_1 = ~new_n1348 & ~new_n1349;
  assign new_n1351 = ~new_n1347 & new_n1350_1;
  assign new_n1352 = new_n1347 & ~new_n1350_1;
  assign new_n1353 = ~new_n1351 & ~new_n1352;
  assign new_n1354 = n1103 & ~n1239;
  assign new_n1355 = n1023 & n1239;
  assign new_n1356 = ~new_n1354 & ~new_n1355;
  assign new_n1357 = ~new_n613 & new_n1356;
  assign new_n1358 = new_n613 & ~new_n1356;
  assign new_n1359_1 = ~new_n1357 & ~new_n1358;
  assign new_n1360 = new_n605 & new_n1359_1;
  assign new_n1361_1 = ~new_n605 & ~new_n1359_1;
  assign new_n1362 = ~new_n1360 & ~new_n1361_1;
  assign new_n1363 = new_n1353 & ~new_n1362;
  assign new_n1364 = ~new_n1353 & new_n1362;
  assign new_n1365 = ~new_n1363 & ~new_n1364;
  assign new_n1366 = ~new_n1344 & ~new_n1365;
  assign new_n1367 = new_n1344 & new_n1365;
  assign new_n1368_1 = ~new_n1366 & ~new_n1367;
  assign new_n1369 = new_n1338 & new_n1368_1;
  assign n1375 = ~new_n1306_1 | ~new_n1369;
  assign new_n1371 = n743 & n1095;
  assign new_n1372 = n478 & n581;
  assign n1752 = ~new_n1371 | ~new_n1372;
  assign new_n1374 = n1054 & n1286;
  assign new_n1375_1 = n593 & n1040;
  assign n1594 = ~new_n1374 | ~new_n1375_1;
  assign new_n1377 = ~n1752 & ~n1594;
  assign new_n1378 = ~n126 & new_n1377;
  assign new_n1379 = ~n669 & new_n1378;
  assign new_n1380 = ~n1375 & new_n1379;
  assign new_n1381 = n559 & ~n1239;
  assign new_n1382 = ~n487 & n1239;
  assign new_n1383 = ~new_n1381 & ~new_n1382;
  assign new_n1384 = new_n862 & ~new_n1383;
  assign new_n1385 = ~new_n862 & new_n1383;
  assign new_n1386_1 = ~new_n1384 & ~new_n1385;
  assign new_n1387_1 = ~n1239 & n1346;
  assign new_n1388 = ~n831 & n1239;
  assign new_n1389_1 = ~new_n1387_1 & ~new_n1388;
  assign new_n1390 = new_n838 & new_n845;
  assign new_n1391_1 = ~new_n838 & ~new_n845;
  assign new_n1392 = ~new_n1390 & ~new_n1391_1;
  assign new_n1393_1 = ~new_n1389_1 & new_n1392;
  assign new_n1394 = new_n1389_1 & ~new_n1392;
  assign new_n1395 = ~new_n1393_1 & ~new_n1394;
  assign new_n1396 = new_n1386_1 & new_n1395;
  assign new_n1397 = ~new_n1386_1 & ~new_n1395;
  assign new_n1398 = ~new_n1396 & ~new_n1397;
  assign new_n1399 = n589 & ~n1239;
  assign new_n1400 = ~n200 & n1239;
  assign new_n1401_1 = ~new_n1399 & ~new_n1400;
  assign new_n1402 = new_n832_1 & new_n855;
  assign new_n1403 = ~new_n832_1 & ~new_n855;
  assign new_n1404 = ~new_n1402 & ~new_n1403;
  assign new_n1405 = ~new_n1401_1 & new_n1404;
  assign new_n1406 = new_n1401_1 & ~new_n1404;
  assign new_n1407 = ~new_n1405 & ~new_n1406;
  assign new_n1408 = new_n1398 & new_n1407;
  assign new_n1409 = ~new_n1398 & ~new_n1407;
  assign new_n1410 = ~new_n1408 & ~new_n1409;
  assign new_n1411_1 = new_n685 & new_n691;
  assign new_n1412 = ~new_n685 & ~new_n691;
  assign new_n1413 = ~new_n1411_1 & ~new_n1412;
  assign new_n1414 = new_n664 & new_n670;
  assign new_n1415_1 = ~new_n664 & ~new_n670;
  assign new_n1416 = ~new_n1414 & ~new_n1415_1;
  assign new_n1417 = ~new_n1413 & new_n1416;
  assign new_n1418_1 = new_n1413 & ~new_n1416;
  assign new_n1419 = ~new_n1417 & ~new_n1418_1;
  assign new_n1420_1 = n947 & n1239;
  assign new_n1421_1 = ~n1239 & ~n1750;
  assign new_n1422 = ~new_n1420_1 & ~new_n1421_1;
  assign new_n1423 = ~new_n676_1 & new_n1422;
  assign new_n1424 = new_n676_1 & ~new_n1422;
  assign new_n1425 = ~new_n1423 & ~new_n1424;
  assign new_n1426 = new_n656 & new_n702;
  assign new_n1427_1 = ~new_n656 & ~new_n702;
  assign new_n1428_1 = ~new_n1426 & ~new_n1427_1;
  assign new_n1429 = new_n1425 & new_n1428_1;
  assign new_n1430 = ~new_n1425 & ~new_n1428_1;
  assign new_n1431 = ~new_n1429 & ~new_n1430;
  assign new_n1432 = ~new_n723 & new_n729_1;
  assign new_n1433 = new_n723 & ~new_n729_1;
  assign new_n1434 = ~new_n1432 & ~new_n1433;
  assign new_n1435_1 = ~new_n1431 & new_n1434;
  assign new_n1436 = new_n1431 & ~new_n1434;
  assign new_n1437 = ~new_n1435_1 & ~new_n1436;
  assign new_n1438_1 = ~new_n1419 & new_n1437;
  assign new_n1439 = new_n1419 & ~new_n1437;
  assign new_n1440 = ~new_n1438_1 & ~new_n1439;
  assign new_n1441 = ~new_n1410 & new_n1440;
  assign new_n1442 = new_n566 & new_n572;
  assign new_n1443_1 = ~new_n566 & ~new_n572;
  assign new_n1444 = ~new_n1442 & ~new_n1443_1;
  assign new_n1445 = new_n599 & ~new_n608_1;
  assign new_n1446_1 = ~new_n599 & new_n608_1;
  assign new_n1447 = ~new_n1445 & ~new_n1446_1;
  assign new_n1448_1 = new_n584 & new_n590;
  assign new_n1449 = ~new_n584 & ~new_n590;
  assign new_n1450 = ~new_n1448_1 & ~new_n1449;
  assign new_n1451 = new_n1447 & ~new_n1450;
  assign new_n1452 = ~new_n1447 & new_n1450;
  assign new_n1453 = ~new_n1451 & ~new_n1452;
  assign new_n1454 = ~new_n1444 & ~new_n1453;
  assign new_n1455 = new_n1444 & new_n1453;
  assign new_n1456 = ~new_n1454 & ~new_n1455;
  assign new_n1457 = new_n616 & new_n631;
  assign new_n1458 = ~new_n616 & ~new_n631;
  assign new_n1459 = ~new_n1457 & ~new_n1458;
  assign new_n1460 = n21 & n1239;
  assign new_n1461 = ~n1239 & ~n1644;
  assign new_n1462 = ~new_n1460 & ~new_n1461;
  assign new_n1463_1 = ~new_n625_1 & new_n1462;
  assign new_n1464 = new_n625_1 & ~new_n1462;
  assign new_n1465 = ~new_n1463_1 & ~new_n1464;
  assign new_n1466 = ~new_n1459 & new_n1465;
  assign new_n1467 = new_n1459 & ~new_n1465;
  assign new_n1468 = ~new_n1466 & ~new_n1467;
  assign new_n1469 = new_n1456 & new_n1468;
  assign new_n1470_1 = ~new_n1456 & ~new_n1468;
  assign new_n1471 = ~new_n1469 & ~new_n1470_1;
  assign new_n1472 = new_n764 & ~new_n770;
  assign new_n1473 = ~new_n764 & new_n770;
  assign new_n1474_1 = ~new_n1472 & ~new_n1473;
  assign new_n1475 = new_n750 & new_n758;
  assign new_n1476_1 = ~new_n750 & ~new_n758;
  assign new_n1477 = ~new_n1475 & ~new_n1476_1;
  assign new_n1478 = new_n1474_1 & new_n1477;
  assign new_n1479 = ~new_n1474_1 & ~new_n1477;
  assign new_n1480 = ~new_n1478 & ~new_n1479;
  assign new_n1481 = n1138 & n1239;
  assign new_n1482 = ~n155 & ~n1239;
  assign new_n1483 = ~new_n1481 & ~new_n1482;
  assign new_n1484 = ~new_n1480 & new_n1483;
  assign new_n1485 = new_n1480 & ~new_n1483;
  assign new_n1486 = ~new_n1484 & ~new_n1485;
  assign new_n1487 = n1205 & n1239;
  assign new_n1488 = ~n729 & ~n1239;
  assign new_n1489 = ~new_n1487 & ~new_n1488;
  assign new_n1490 = new_n787_1 & ~new_n1489;
  assign new_n1491 = ~new_n787_1 & new_n1489;
  assign new_n1492 = ~new_n1490 & ~new_n1491;
  assign new_n1493 = new_n708 & new_n714_1;
  assign new_n1494 = ~new_n708 & ~new_n714_1;
  assign new_n1495 = ~new_n1493 & ~new_n1494;
  assign new_n1496 = ~new_n1492 & new_n1495;
  assign new_n1497 = new_n1492 & ~new_n1495;
  assign new_n1498 = ~new_n1496 & ~new_n1497;
  assign new_n1499 = new_n776 & new_n1498;
  assign new_n1500_1 = ~new_n776 & ~new_n1498;
  assign new_n1501 = ~new_n1499 & ~new_n1500_1;
  assign new_n1502_1 = ~new_n1486 & new_n1501;
  assign new_n1503 = new_n1486 & ~new_n1501;
  assign new_n1504 = ~new_n1502_1 & ~new_n1503;
  assign new_n1505 = ~new_n1471 & ~new_n1504;
  assign n1322 = ~new_n1441 | ~new_n1505;
  assign new_n1507 = ~n775 & n1626;
  assign new_n1508 = n775 & ~n1626;
  assign new_n1509 = ~new_n1507 & ~new_n1508;
  assign new_n1510 = n430 & new_n1509;
  assign new_n1511 = ~n430 & ~new_n1509;
  assign new_n1512 = ~new_n1510 & ~new_n1511;
  assign new_n1513 = new_n1256 & new_n1512;
  assign new_n1514 = new_n897 & new_n901;
  assign new_n1515 = new_n896 & new_n902;
  assign new_n1516_1 = ~new_n1514 & ~new_n1515;
  assign new_n1517 = new_n1036 & new_n1056;
  assign new_n1518 = new_n1037 & new_n1055;
  assign new_n1519 = ~new_n1517 & ~new_n1518;
  assign new_n1520_1 = ~new_n1516_1 & new_n1519;
  assign new_n1521_1 = new_n1516_1 & ~new_n1519;
  assign new_n1522 = ~new_n1520_1 & ~new_n1521_1;
  assign new_n1523_1 = ~new_n1513 & new_n1522;
  assign new_n1524 = new_n1513 & ~new_n1522;
  assign new_n1525 = ~new_n1523_1 & ~new_n1524;
  assign new_n1526 = new_n469 & new_n475;
  assign new_n1527_1 = ~new_n469 & ~new_n475;
  assign new_n1528 = ~new_n1526 & ~new_n1527_1;
  assign new_n1529 = new_n437 & new_n450;
  assign new_n1530 = ~new_n437 & ~new_n450;
  assign new_n1531 = ~new_n1529 & ~new_n1530;
  assign new_n1532 = ~new_n1528 & new_n1531;
  assign new_n1533 = new_n1528 & ~new_n1531;
  assign new_n1534_1 = ~new_n1532 & ~new_n1533;
  assign new_n1535 = ~new_n456 & new_n462;
  assign new_n1536_1 = new_n456 & ~new_n462;
  assign new_n1537 = ~new_n1535 & ~new_n1536_1;
  assign new_n1538 = n1239 & n1281;
  assign new_n1539 = ~new_n1307 & ~new_n1538;
  assign new_n1540 = ~n961 & n1239;
  assign new_n1541 = ~new_n489_1 & ~new_n1540;
  assign new_n1542 = ~new_n1539 & new_n1541;
  assign new_n1543 = new_n1539 & ~new_n1541;
  assign new_n1544 = ~new_n1542 & ~new_n1543;
  assign new_n1545 = new_n431 & new_n444;
  assign new_n1546 = ~new_n431 & ~new_n444;
  assign new_n1547_1 = ~new_n1545 & ~new_n1546;
  assign new_n1548_1 = new_n1544 & new_n1547_1;
  assign new_n1549 = ~new_n1544 & ~new_n1547_1;
  assign new_n1550 = ~new_n1548_1 & ~new_n1549;
  assign new_n1551 = new_n1537 & ~new_n1550;
  assign new_n1552 = ~new_n1537 & new_n1550;
  assign new_n1553 = ~new_n1551 & ~new_n1552;
  assign new_n1554 = ~new_n1534_1 & ~new_n1553;
  assign new_n1555 = new_n1534_1 & new_n1553;
  assign new_n1556 = ~new_n1554 & ~new_n1555;
  assign new_n1557 = ~new_n1525 & ~new_n1556;
  assign new_n1558 = n117 & n1239;
  assign new_n1559 = ~new_n1354 & ~new_n1558;
  assign new_n1560 = new_n359 & ~new_n1559;
  assign new_n1561 = ~new_n359 & new_n1559;
  assign new_n1562 = ~new_n1560 & ~new_n1561;
  assign new_n1563 = new_n344_1 & new_n349;
  assign new_n1564 = ~new_n344_1 & ~new_n349;
  assign new_n1565 = ~new_n1563 & ~new_n1564;
  assign new_n1566_1 = new_n1562 & ~new_n1565;
  assign new_n1567 = ~new_n1562 & new_n1565;
  assign new_n1568 = ~new_n1566_1 & ~new_n1567;
  assign new_n1569_1 = new_n354 & new_n363;
  assign new_n1570 = ~new_n354 & ~new_n363;
  assign new_n1571 = ~new_n1569_1 & ~new_n1570;
  assign new_n1572 = new_n327 & new_n331;
  assign new_n1573 = new_n326 & new_n332;
  assign new_n1574 = ~new_n1572 & ~new_n1573;
  assign new_n1575 = new_n318_1 & new_n322;
  assign new_n1576_1 = new_n317 & new_n323;
  assign new_n1577 = ~new_n1575 & ~new_n1576_1;
  assign new_n1578 = new_n1574 & new_n1577;
  assign new_n1579 = ~new_n1574 & ~new_n1577;
  assign new_n1580 = ~new_n1578 & ~new_n1579;
  assign new_n1581 = new_n1571 & ~new_n1580;
  assign new_n1582 = ~new_n1571 & new_n1580;
  assign new_n1583 = ~new_n1581 & ~new_n1582;
  assign new_n1584 = ~new_n1568 & ~new_n1583;
  assign new_n1585 = new_n1568 & new_n1583;
  assign new_n1586_1 = ~new_n1584 & ~new_n1585;
  assign new_n1587 = new_n404 & new_n409_1;
  assign new_n1588_1 = ~new_n404 & ~new_n409_1;
  assign new_n1589 = ~new_n1587 & ~new_n1588_1;
  assign new_n1590 = n314 & n1239;
  assign new_n1591 = ~new_n1285_1 & ~new_n1590;
  assign new_n1592_1 = ~new_n419 & new_n1591;
  assign new_n1593 = new_n419 & ~new_n1591;
  assign new_n1594_1 = ~new_n1592_1 & ~new_n1593;
  assign new_n1595 = ~new_n1589 & new_n1594_1;
  assign new_n1596 = new_n1589 & ~new_n1594_1;
  assign new_n1597 = ~new_n1595 & ~new_n1596;
  assign new_n1598 = new_n399_1 & new_n414;
  assign new_n1599 = ~new_n399_1 & ~new_n414;
  assign new_n1600 = ~new_n1598 & ~new_n1599;
  assign new_n1601 = ~new_n1597 & new_n1600;
  assign new_n1602 = new_n1597 & ~new_n1600;
  assign new_n1603 = ~new_n1601 & ~new_n1602;
  assign new_n1604 = new_n386 & new_n530;
  assign new_n1605 = ~new_n386 & ~new_n530;
  assign new_n1606 = ~new_n1604 & ~new_n1605;
  assign new_n1607 = new_n523 & new_n1606;
  assign new_n1608 = ~new_n523 & ~new_n1606;
  assign new_n1609_1 = ~new_n1607 & ~new_n1608;
  assign new_n1610 = new_n392_1 & new_n1609_1;
  assign new_n1611 = ~new_n392_1 & ~new_n1609_1;
  assign new_n1612 = ~new_n1610 & ~new_n1611;
  assign new_n1613_1 = ~new_n1603 & new_n1612;
  assign new_n1614 = new_n1603 & ~new_n1612;
  assign new_n1615 = ~new_n1613_1 & ~new_n1614;
  assign new_n1616_1 = new_n1586_1 & new_n1615;
  assign n1288 = ~new_n1557 | ~new_n1616_1;
  assign new_n1618 = ~n1322 & ~n1288;
  assign n918 = ~new_n1380 | ~new_n1618;
  assign new_n1620 = ~new_n511 & new_n1018;
  assign n952 = ~new_n1019 & ~new_n1620;
  assign new_n1622 = ~new_n1044_1 & ~new_n1101;
  assign new_n1623 = ~new_n1038 & ~new_n1622;
  assign new_n1624 = ~new_n1059 & ~new_n1623;
  assign new_n1625 = new_n1059 & new_n1623;
  assign n990 = ~new_n1624 & ~new_n1625;
  assign new_n1627_1 = ~new_n453_1 & new_n498_1;
  assign n1006 = ~new_n499 & ~new_n1627_1;
  assign new_n1629 = n380 & ~n1361;
  assign n1050 = ~n701 | ~new_n1629;
  assign new_n1631 = ~new_n377 & new_n1143;
  assign n1051 = ~new_n1144 & ~new_n1631;
  assign new_n1633 = ~new_n471 & ~new_n1248;
  assign new_n1634 = ~new_n465 & new_n1633;
  assign new_n1635 = new_n465 & ~new_n1633;
  assign n1058 = ~new_n1634 & ~new_n1635;
  assign new_n1637 = ~new_n527 & ~new_n1163;
  assign n1060 = ~new_n534_1 & ~new_n1637;
  assign new_n1639_1 = new_n508 & ~new_n510_1;
  assign n1063 = ~new_n1015 & ~new_n1639_1;
  assign new_n1641 = new_n373 & ~new_n383;
  assign new_n1642 = new_n335 & ~new_n340;
  assign new_n1643 = new_n325 & ~new_n1642;
  assign new_n1644_1 = new_n324 & new_n1642;
  assign new_n1645_1 = ~new_n1643 & ~new_n1644_1;
  assign new_n1646 = ~new_n321 & ~new_n341_1;
  assign new_n1647_1 = ~new_n914 & ~new_n1646;
  assign new_n1648 = ~new_n330 & ~new_n333;
  assign new_n1649 = ~new_n334 & ~new_n1648;
  assign new_n1650 = ~new_n1647_1 & new_n1649;
  assign new_n1651 = new_n1647_1 & ~new_n1649;
  assign new_n1652 = ~new_n1650 & ~new_n1651;
  assign new_n1653 = new_n1645_1 & new_n1652;
  assign new_n1654 = ~new_n1645_1 & ~new_n1652;
  assign new_n1655 = ~new_n1653 & ~new_n1654;
  assign new_n1656_1 = ~new_n1641 & new_n1655;
  assign new_n1657 = ~new_n542 & new_n1656_1;
  assign new_n1658 = ~new_n334 & new_n911;
  assign new_n1659 = ~new_n336 & ~new_n1658;
  assign new_n1660 = ~new_n330 & new_n338;
  assign new_n1661 = ~new_n339 & ~new_n1660;
  assign new_n1662 = new_n1647_1 & ~new_n1661;
  assign new_n1663 = ~new_n1647_1 & new_n1661;
  assign new_n1664 = ~new_n1662 & ~new_n1663;
  assign new_n1665 = ~new_n1659 & new_n1664;
  assign new_n1666 = new_n1659 & ~new_n1664;
  assign new_n1667 = ~new_n1665 & ~new_n1666;
  assign new_n1668 = new_n373 & ~new_n1667;
  assign new_n1669 = ~new_n373 & new_n1655;
  assign new_n1670 = ~new_n1668 & ~new_n1669;
  assign new_n1671 = new_n542 & ~new_n1670;
  assign new_n1672 = new_n1641 & ~new_n1667;
  assign new_n1673 = ~new_n1671 & ~new_n1672;
  assign new_n1674 = ~new_n1657 & new_n1673;
  assign new_n1675 = new_n371 & new_n375;
  assign new_n1676 = ~new_n371 & ~new_n375;
  assign new_n1677 = ~new_n1675 & ~new_n1676;
  assign new_n1678 = ~new_n360 & ~new_n364_1;
  assign new_n1679 = ~new_n366 & ~new_n1678;
  assign new_n1680 = ~new_n380_1 & ~new_n381;
  assign new_n1681 = ~new_n382 & ~new_n1680;
  assign new_n1682 = new_n1679 & ~new_n1681;
  assign new_n1683 = ~new_n1679 & new_n1681;
  assign new_n1684 = ~new_n1682 & ~new_n1683;
  assign new_n1685 = ~new_n376_1 & ~new_n377;
  assign new_n1686 = ~new_n378_1 & ~new_n1685;
  assign new_n1687_1 = new_n369 & ~new_n1686;
  assign new_n1688 = ~new_n369 & new_n1686;
  assign new_n1689 = ~new_n1687_1 & ~new_n1688;
  assign new_n1690 = ~new_n1684 & new_n1689;
  assign new_n1691 = new_n1684 & ~new_n1689;
  assign new_n1692 = ~new_n1690 & ~new_n1691;
  assign new_n1693 = ~new_n1677 & new_n1692;
  assign new_n1694 = new_n1677 & ~new_n1692;
  assign new_n1695 = ~new_n1693 & ~new_n1694;
  assign new_n1696 = new_n542 & ~new_n1695;
  assign new_n1697 = new_n375 & new_n886;
  assign new_n1698 = ~new_n1676 & ~new_n1697;
  assign new_n1699 = new_n369 & new_n374_1;
  assign new_n1700 = ~new_n369 & ~new_n374_1;
  assign new_n1701 = ~new_n1699 & ~new_n1700;
  assign new_n1702 = ~new_n379 & new_n1701;
  assign new_n1703 = ~new_n360 & new_n374_1;
  assign new_n1704 = ~new_n365 & ~new_n1703;
  assign new_n1705 = new_n1681 & new_n1704;
  assign new_n1706 = ~new_n1681 & ~new_n1704;
  assign new_n1707 = ~new_n1705 & ~new_n1706;
  assign new_n1708 = ~new_n1686 & new_n1707;
  assign new_n1709 = new_n1686 & ~new_n1707;
  assign new_n1710 = ~new_n1708 & ~new_n1709;
  assign new_n1711 = ~new_n1702 & new_n1710;
  assign new_n1712 = new_n1702 & ~new_n1710;
  assign new_n1713 = ~new_n1711 & ~new_n1712;
  assign new_n1714 = new_n1698 & new_n1713;
  assign new_n1715 = ~new_n1698 & ~new_n1713;
  assign new_n1716 = ~new_n1714 & ~new_n1715;
  assign new_n1717 = ~new_n542 & ~new_n1716;
  assign new_n1718 = ~new_n1696 & ~new_n1717;
  assign new_n1719 = new_n1674 & ~new_n1718;
  assign new_n1720 = ~new_n1674 & new_n1718;
  assign n1065 = new_n1719 | new_n1720;
  assign new_n1722 = ~new_n500 & new_n503;
  assign new_n1723 = ~new_n440 & new_n1722;
  assign new_n1724 = new_n440 & ~new_n1722;
  assign n1195 = ~new_n1723 & ~new_n1724;
  assign new_n1726 = ~new_n905_1 & new_n921;
  assign n1302 = ~new_n922 & ~new_n1726;
  assign new_n1728 = ~new_n1060_1 & ~new_n1101;
  assign n1391 = ~new_n1102 & ~new_n1728;
  assign new_n1730 = ~new_n492 & new_n1244;
  assign n1420 = ~new_n1245 & ~new_n1730;
  assign new_n1732 = ~new_n451 & new_n498_1;
  assign new_n1733 = ~new_n452 & ~new_n1732;
  assign new_n1734 = new_n447 & new_n1733;
  assign new_n1735 = ~new_n447 & ~new_n1733;
  assign n1427 = ~new_n1734 & ~new_n1735;
  assign new_n1737 = ~new_n375 & new_n542;
  assign n1527 = ~new_n1142 & ~new_n1737;
  assign new_n1739 = n545 & new_n495;
  assign new_n1740 = ~new_n983 & ~new_n1739;
  assign new_n1741 = new_n459 & new_n1740;
  assign new_n1742 = ~new_n459 & ~new_n1740;
  assign n1639 = new_n1741 | new_n1742;
  assign new_n1744 = ~new_n534_1 & ~new_n537;
  assign new_n1745 = ~new_n395 & ~new_n1744;
  assign new_n1746 = new_n395 & new_n1744;
  assign n1687 = new_n1745 | new_n1746;
  assign n275 = ~n992;
  assign n23 = n346;
  assign n27 = n947;
  assign n85 = n153;
  assign n130 = n1592;
  assign n173 = n823;
  assign n184 = n420;
  assign n230 = n831;
  assign n292 = n408;
  assign n301 = n318;
  assign n337 = n626;
  assign n352 = n1463;
  assign n362 = n30;
  assign n417 = n399;
  assign n457 = n161;
  assign n460 = n21;
  assign n497 = n1656;
  assign n498 = n293;
  assign n501 = n200;
  assign n509 = n769;
  assign n516 = n1187;
  assign n585 = n553;
  assign n595 = n1301;
  assign n638 = n420;
  assign n640 = n1345;
  assign n726 = n275;
  assign n773 = n980;
  assign n782 = n222;
  assign n821 = n374;
  assign n842 = n1205;
  assign n1017 = n1476;
  assign n1042 = n1566;
  assign n1177 = n487;
  assign n1186 = n553;
  assign n1209 = n1071;
  assign n1211 = n161;
  assign n1231 = n1470;
  assign n1234 = n608;
  assign n1253 = n1050;
  assign n1285 = n1401;
  assign n1292 = n1616;
  assign n1296 = n275;
  assign n1320 = n1263;
  assign n1337 = n1138;
  assign n1359 = n453;
  assign n1368 = n420;
  assign n1421 = n695;
  assign n1534 = n920;
  assign n1547 = n420;
  assign n1548 = n567;
  assign n1588 = n428;
  assign n1632 = n553;
  assign n1645 = n1446;
  assign n1729 = n138;
  assign n1738 = n45;
endmodule


