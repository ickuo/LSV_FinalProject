// Benchmark "top" written by ABC on Sun Dec 21 18:06:36 2025

module top ( 
    n0, n2, n17, n18, n23, n27, n29, n37, n43, n58, n59, n70, n75, n84,
    n90, n91, n107, n130, n133, n137, n169, n174, n179, n187, n194, n196,
    n210, n211, n214, n226, n234, n237, n238, n249, n256, n260, n272, n278,
    n281, n289, n292,
    n24, n26, n61, n66, n73, n80, n81, n86, n88, n89, n94, n98, n104, n123,
    n129, n145, n151, n160, n164, n168, n199, n212, n213, n217, n221, n246,
    n253, n261, n265, n286, n304, n310  );
  input  n0, n2, n17, n18, n23, n27, n29, n37, n43, n58, n59, n70, n75,
    n84, n90, n91, n107, n130, n133, n137, n169, n174, n179, n187, n194,
    n196, n210, n211, n214, n226, n234, n237, n238, n249, n256, n260, n272,
    n278, n281, n289, n292;
  output n24, n26, n61, n66, n73, n80, n81, n86, n88, n89, n94, n98, n104,
    n123, n129, n145, n151, n160, n164, n168, n199, n212, n213, n217, n221,
    n246, n253, n261, n265, n286, n304, n310;
  wire new_n74, new_n75_1, new_n76, new_n77, new_n78, new_n79, new_n80_1,
    new_n81_1, new_n82, new_n83, new_n84_1, new_n85, new_n86_1, new_n87,
    new_n88_1, new_n89_1, new_n90_1, new_n91_1, new_n92, new_n93,
    new_n94_1, new_n95, new_n96, new_n97, new_n98_1, new_n99, new_n100,
    new_n101, new_n102, new_n103, new_n104_1, new_n105, new_n106,
    new_n107_1, new_n108, new_n109, new_n110, new_n111, new_n112, new_n113,
    new_n114, new_n115, new_n116, new_n117, new_n118, new_n119, new_n120,
    new_n121, new_n122, new_n123_1, new_n124, new_n125, new_n126, new_n127,
    new_n128, new_n129_1, new_n130_1, new_n131, new_n132, new_n133_1,
    new_n134, new_n135, new_n136, new_n137_1, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145_1, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151_1, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n158, new_n159, new_n160_1, new_n161,
    new_n162, new_n163, new_n164_1, new_n165, new_n166, new_n167,
    new_n168_1, new_n169_1, new_n170, new_n171, new_n172, new_n173,
    new_n174_1, new_n175, new_n176, new_n177, new_n178, new_n179_1,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187_1, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194_1, new_n195, new_n196_1, new_n197, new_n198, new_n199_1,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210_1, new_n211_1, new_n212_1,
    new_n213_1, new_n214_1, new_n215, new_n216, new_n217_1, new_n218,
    new_n219, new_n220, new_n221_1, new_n222, new_n223, new_n224, new_n225,
    new_n226_1, new_n227, new_n228, new_n229, new_n230, new_n231, new_n232,
    new_n233, new_n234_1, new_n235, new_n236, new_n237_1, new_n238_1,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246_1, new_n247, new_n248, new_n249_1, new_n250, new_n251,
    new_n252, new_n253_1, new_n254, new_n255, new_n256_1, new_n257,
    new_n258, new_n259, new_n260_1, new_n261_1, new_n262, new_n263,
    new_n264, new_n265_1, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272_1, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278_1, new_n279, new_n280, new_n281_1, new_n282, new_n283,
    new_n284, new_n285, new_n286_1, new_n287, new_n288, new_n289_1,
    new_n290, new_n291, new_n292_1, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304_1, new_n305, new_n306, new_n308, new_n309, new_n310_1,
    new_n311, new_n312, new_n313, new_n314, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n346, new_n347, new_n348, new_n350, new_n351,
    new_n352, new_n353, new_n355, new_n356, new_n357, new_n358, new_n360,
    new_n361, new_n362, new_n363, new_n365, new_n366, new_n367, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n375, new_n376, new_n377,
    new_n378, new_n380, new_n381, new_n382, new_n383, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n391, new_n392, new_n393, new_n394,
    new_n396, new_n397, new_n398, new_n400, new_n401, new_n402, new_n404,
    new_n405, new_n406, new_n408, new_n409, new_n410, new_n412, new_n413,
    new_n414, new_n416, new_n417, new_n418, new_n419, new_n421, new_n422,
    new_n423, new_n425, new_n426, new_n427, new_n429, new_n430, new_n431,
    new_n432, new_n434, new_n435, new_n436, new_n438, new_n439, new_n440,
    new_n442, new_n443, new_n444, new_n446, new_n447, new_n448, new_n450,
    new_n451, new_n452, new_n454, new_n455, new_n456, new_n458, new_n459,
    new_n460;
  assign new_n74 = n133 & n281;
  assign new_n75_1 = ~n27 & ~n194;
  assign new_n76 = n27 & n194;
  assign new_n77 = ~new_n75_1 & ~new_n76;
  assign new_n78 = ~new_n74 & ~new_n77;
  assign new_n79 = new_n74 & new_n77;
  assign new_n80_1 = ~new_n78 & ~new_n79;
  assign new_n81_1 = ~n187 & n211;
  assign new_n82 = n187 & ~n211;
  assign new_n83 = ~new_n81_1 & ~new_n82;
  assign new_n84_1 = new_n80_1 & ~new_n83;
  assign new_n85 = ~new_n80_1 & new_n83;
  assign new_n86_1 = ~new_n84_1 & ~new_n85;
  assign new_n87 = ~n249 & n289;
  assign new_n88_1 = n249 & ~n289;
  assign new_n89_1 = ~new_n87 & ~new_n88_1;
  assign new_n90_1 = n107 & n214;
  assign new_n91_1 = ~n107 & ~n214;
  assign new_n92 = ~new_n90_1 & ~new_n91_1;
  assign new_n93 = new_n89_1 & new_n92;
  assign new_n94_1 = ~new_n89_1 & ~new_n92;
  assign new_n95 = ~new_n93 & ~new_n94_1;
  assign new_n96 = ~n174 & n210;
  assign new_n97 = n174 & ~n210;
  assign new_n98_1 = ~new_n96 & ~new_n97;
  assign new_n99 = n59 & n169;
  assign new_n100 = ~n59 & ~n169;
  assign new_n101 = ~new_n99 & ~new_n100;
  assign new_n102 = new_n98_1 & new_n101;
  assign new_n103 = ~new_n98_1 & ~new_n101;
  assign new_n104_1 = ~new_n102 & ~new_n103;
  assign new_n105 = new_n95 & new_n104_1;
  assign new_n106 = ~new_n95 & ~new_n104_1;
  assign new_n107_1 = ~new_n105 & ~new_n106;
  assign new_n108 = new_n86_1 & new_n107_1;
  assign new_n109 = ~new_n86_1 & ~new_n107_1;
  assign new_n110 = ~new_n108 & ~new_n109;
  assign new_n111 = ~n130 & n256;
  assign new_n112 = n130 & ~n256;
  assign new_n113 = ~new_n111 & ~new_n112;
  assign new_n114 = n23 & n43;
  assign new_n115 = ~n23 & ~n43;
  assign new_n116 = ~new_n114 & ~new_n115;
  assign new_n117 = new_n113 & new_n116;
  assign new_n118 = ~new_n113 & ~new_n116;
  assign new_n119 = ~new_n117 & ~new_n118;
  assign new_n120 = n226 & n281;
  assign new_n121 = ~n137 & ~n260;
  assign new_n122 = n137 & n260;
  assign new_n123_1 = ~new_n121 & ~new_n122;
  assign new_n124 = ~new_n120 & new_n123_1;
  assign new_n125 = new_n120 & ~new_n123_1;
  assign new_n126 = ~new_n124 & ~new_n125;
  assign new_n127 = new_n119 & ~new_n126;
  assign new_n128 = ~new_n119 & new_n126;
  assign new_n129_1 = ~new_n127 & ~new_n128;
  assign new_n130_1 = ~n90 & n237;
  assign new_n131 = n90 & ~n237;
  assign new_n132 = ~new_n130_1 & ~new_n131;
  assign new_n133_1 = n2 & n70;
  assign new_n134 = ~n2 & ~n70;
  assign new_n135 = ~new_n133_1 & ~new_n134;
  assign new_n136 = new_n132 & new_n135;
  assign new_n137_1 = ~new_n132 & ~new_n135;
  assign new_n138 = ~new_n136 & ~new_n137_1;
  assign new_n139 = ~n0 & n179;
  assign new_n140 = n0 & ~n179;
  assign new_n141 = ~new_n139 & ~new_n140;
  assign new_n142 = new_n138 & ~new_n141;
  assign new_n143 = ~new_n138 & new_n141;
  assign new_n144 = ~new_n142 & ~new_n143;
  assign new_n145_1 = ~new_n129_1 & new_n144;
  assign new_n146 = new_n129_1 & ~new_n144;
  assign new_n147 = ~new_n145_1 & ~new_n146;
  assign new_n148 = new_n110 & new_n147;
  assign new_n149 = n84 & n281;
  assign new_n150 = ~n196 & ~n272;
  assign new_n151_1 = n196 & n272;
  assign new_n152 = ~new_n150 & ~new_n151_1;
  assign new_n153 = ~new_n149 & ~new_n152;
  assign new_n154 = new_n149 & new_n152;
  assign new_n155 = ~new_n153 & ~new_n154;
  assign new_n156 = ~n29 & n75;
  assign new_n157 = n29 & ~n75;
  assign new_n158 = ~new_n156 & ~new_n157;
  assign new_n159 = new_n155 & ~new_n158;
  assign new_n160_1 = ~new_n155 & new_n158;
  assign new_n161 = ~new_n159 & ~new_n160_1;
  assign new_n162 = new_n95 & new_n119;
  assign new_n163 = ~new_n95 & ~new_n119;
  assign new_n164_1 = ~new_n162 & ~new_n163;
  assign new_n165 = new_n161 & new_n164_1;
  assign new_n166 = ~new_n161 & ~new_n164_1;
  assign new_n167 = ~new_n165 & ~new_n166;
  assign new_n168_1 = n58 & n281;
  assign new_n169_1 = ~n234 & ~n278;
  assign new_n170 = n234 & n278;
  assign new_n171 = ~new_n169_1 & ~new_n170;
  assign new_n172 = ~new_n168_1 & new_n171;
  assign new_n173 = new_n168_1 & ~new_n171;
  assign new_n174_1 = ~new_n172 & ~new_n173;
  assign new_n175 = new_n104_1 & ~new_n174_1;
  assign new_n176 = ~new_n104_1 & new_n174_1;
  assign new_n177 = ~new_n175 & ~new_n176;
  assign new_n178 = ~n17 & n238;
  assign new_n179_1 = n17 & ~n238;
  assign new_n180 = ~new_n178 & ~new_n179_1;
  assign new_n181 = new_n138 & ~new_n180;
  assign new_n182 = ~new_n138 & new_n180;
  assign new_n183 = ~new_n181 & ~new_n182;
  assign new_n184 = ~new_n177 & new_n183;
  assign new_n185 = new_n177 & ~new_n183;
  assign new_n186 = ~new_n184 & ~new_n185;
  assign new_n187_1 = ~new_n167 & ~new_n186;
  assign new_n188 = ~n23 & n249;
  assign new_n189 = n23 & ~n249;
  assign new_n190 = ~new_n188 & ~new_n189;
  assign new_n191 = ~n272 & n278;
  assign new_n192 = n272 & ~n278;
  assign new_n193 = ~new_n191 & ~new_n192;
  assign new_n194_1 = n137 & n194;
  assign new_n195 = ~n137 & ~n194;
  assign new_n196_1 = ~new_n194_1 & ~new_n195;
  assign new_n197 = new_n193 & new_n196_1;
  assign new_n198 = ~new_n193 & ~new_n196_1;
  assign new_n199_1 = ~new_n197 & ~new_n198;
  assign new_n200 = ~new_n190 & new_n199_1;
  assign new_n201 = new_n190 & ~new_n199_1;
  assign new_n202 = ~new_n200 & ~new_n201;
  assign new_n203 = ~n234 & n260;
  assign new_n204 = n234 & ~n260;
  assign new_n205 = ~new_n203 & ~new_n204;
  assign new_n206 = n27 & n196;
  assign new_n207 = ~n27 & ~n196;
  assign new_n208 = ~new_n206 & ~new_n207;
  assign new_n209 = new_n205 & new_n208;
  assign new_n210_1 = ~new_n205 & ~new_n208;
  assign new_n211_1 = ~new_n209 & ~new_n210_1;
  assign new_n212_1 = n91 & n281;
  assign new_n213_1 = ~n210 & ~n237;
  assign new_n214_1 = n210 & n237;
  assign new_n215 = ~new_n213_1 & ~new_n214_1;
  assign new_n216 = ~new_n212_1 & ~new_n215;
  assign new_n217_1 = new_n212_1 & new_n215;
  assign new_n218 = ~new_n216 & ~new_n217_1;
  assign new_n219 = new_n211_1 & new_n218;
  assign new_n220 = ~new_n211_1 & ~new_n218;
  assign new_n221_1 = ~new_n219 & ~new_n220;
  assign new_n222 = new_n202 & new_n221_1;
  assign new_n223 = ~new_n202 & ~new_n221_1;
  assign new_n224 = ~new_n222 & ~new_n223;
  assign new_n225 = n281 & n292;
  assign new_n226_1 = ~n59 & ~n90;
  assign new_n227 = n59 & n90;
  assign new_n228 = ~new_n226_1 & ~new_n227;
  assign new_n229 = ~new_n225 & ~new_n228;
  assign new_n230 = new_n225 & new_n228;
  assign new_n231 = ~new_n229 & ~new_n230;
  assign new_n232 = ~n43 & n214;
  assign new_n233 = n43 & ~n214;
  assign new_n234_1 = ~new_n232 & ~new_n233;
  assign new_n235 = new_n231 & ~new_n234_1;
  assign new_n236 = ~new_n231 & new_n234_1;
  assign new_n237_1 = ~new_n235 & ~new_n236;
  assign new_n238_1 = ~n75 & n211;
  assign new_n239 = n75 & ~n211;
  assign new_n240 = ~new_n238_1 & ~new_n239;
  assign new_n241 = n0 & n17;
  assign new_n242 = ~n0 & ~n17;
  assign new_n243 = ~new_n241 & ~new_n242;
  assign new_n244 = new_n240 & new_n243;
  assign new_n245 = ~new_n240 & ~new_n243;
  assign new_n246_1 = ~new_n244 & ~new_n245;
  assign new_n247 = ~n187 & n238;
  assign new_n248 = n187 & ~n238;
  assign new_n249_1 = ~new_n247 & ~new_n248;
  assign new_n250 = n29 & n179;
  assign new_n251 = ~n29 & ~n179;
  assign new_n252 = ~new_n250 & ~new_n251;
  assign new_n253_1 = new_n249_1 & new_n252;
  assign new_n254 = ~new_n249_1 & ~new_n252;
  assign new_n255 = ~new_n253_1 & ~new_n254;
  assign new_n256_1 = new_n246_1 & new_n255;
  assign new_n257 = ~new_n246_1 & ~new_n255;
  assign new_n258 = ~new_n256_1 & ~new_n257;
  assign new_n259 = new_n237_1 & new_n258;
  assign new_n260_1 = ~new_n237_1 & ~new_n258;
  assign new_n261_1 = ~new_n259 & ~new_n260_1;
  assign new_n262 = ~new_n224 & new_n261_1;
  assign new_n263 = n18 & n281;
  assign new_n264 = ~n2 & ~n169;
  assign new_n265_1 = n2 & n169;
  assign new_n266 = ~new_n264 & ~new_n265_1;
  assign new_n267 = ~new_n263 & ~new_n266;
  assign new_n268 = new_n263 & new_n266;
  assign new_n269 = ~new_n267 & ~new_n268;
  assign new_n270 = ~n256 & n289;
  assign new_n271 = n256 & ~n289;
  assign new_n272_1 = ~new_n270 & ~new_n271;
  assign new_n273 = new_n269 & ~new_n272_1;
  assign new_n274 = ~new_n269 & new_n272_1;
  assign new_n275 = ~new_n273 & ~new_n274;
  assign new_n276 = new_n211_1 & new_n246_1;
  assign new_n277 = ~new_n211_1 & ~new_n246_1;
  assign new_n278_1 = ~new_n276 & ~new_n277;
  assign new_n279 = new_n275 & new_n278_1;
  assign new_n280 = ~new_n275 & ~new_n278_1;
  assign new_n281_1 = ~new_n279 & ~new_n280;
  assign new_n282 = n37 & n281;
  assign new_n283 = ~n70 & ~n174;
  assign new_n284 = n70 & n174;
  assign new_n285 = ~new_n283 & ~new_n284;
  assign new_n286_1 = ~new_n282 & ~new_n285;
  assign new_n287 = new_n282 & new_n285;
  assign new_n288 = ~new_n286_1 & ~new_n287;
  assign new_n289_1 = ~n107 & n130;
  assign new_n290 = n107 & ~n130;
  assign new_n291 = ~new_n289_1 & ~new_n290;
  assign new_n292_1 = new_n288 & ~new_n291;
  assign new_n293 = ~new_n288 & new_n291;
  assign new_n294 = ~new_n292_1 & ~new_n293;
  assign new_n295 = new_n199_1 & new_n255;
  assign new_n296 = ~new_n199_1 & ~new_n255;
  assign new_n297 = ~new_n295 & ~new_n296;
  assign new_n298 = new_n294 & new_n297;
  assign new_n299 = ~new_n294 & ~new_n297;
  assign new_n300 = ~new_n298 & ~new_n299;
  assign new_n301 = ~new_n281_1 & ~new_n300;
  assign new_n302 = new_n262 & new_n301;
  assign new_n303 = new_n187_1 & new_n302;
  assign new_n304_1 = new_n148 & new_n303;
  assign new_n305 = n59 & ~new_n304_1;
  assign new_n306 = ~n59 & new_n304_1;
  assign n24 = new_n305 | new_n306;
  assign new_n308 = ~new_n224 & ~new_n261_1;
  assign new_n309 = new_n281_1 & ~new_n300;
  assign new_n310_1 = new_n308 & new_n309;
  assign new_n311 = new_n187_1 & new_n310_1;
  assign new_n312 = new_n148 & new_n311;
  assign new_n313 = n169 & ~new_n312;
  assign new_n314 = ~n169 & new_n312;
  assign n26 = new_n313 | new_n314;
  assign new_n316 = ~new_n110 & new_n147;
  assign new_n317 = new_n187_1 & new_n316;
  assign new_n318 = new_n262 & new_n317;
  assign new_n319 = new_n309 & new_n318;
  assign new_n320 = ~n17 & ~new_n319;
  assign new_n321 = n17 & new_n319;
  assign n61 = ~new_n320 & ~new_n321;
  assign new_n323 = ~new_n281_1 & new_n300;
  assign new_n324 = new_n167 & new_n186;
  assign new_n325 = new_n316 & new_n324;
  assign new_n326 = new_n262 & new_n325;
  assign new_n327 = new_n323 & new_n326;
  assign new_n328 = ~n29 & ~new_n327;
  assign new_n329 = n29 & new_n327;
  assign n66 = ~new_n328 & ~new_n329;
  assign new_n331 = new_n224 & ~new_n261_1;
  assign new_n332 = ~new_n167 & new_n186;
  assign new_n333 = ~new_n110 & ~new_n147;
  assign new_n334 = new_n332 & new_n333;
  assign new_n335 = new_n331 & new_n334;
  assign new_n336 = new_n309 & new_n335;
  assign new_n337 = n260 & ~new_n336;
  assign new_n338 = ~n260 & new_n336;
  assign n73 = new_n337 | new_n338;
  assign new_n340 = new_n308 & new_n323;
  assign new_n341 = new_n187_1 & new_n340;
  assign new_n342 = new_n148 & new_n341;
  assign new_n343 = n174 & ~new_n342;
  assign new_n344 = ~n174 & new_n342;
  assign n80 = new_n343 | new_n344;
  assign new_n346 = new_n303 & new_n333;
  assign new_n347 = n90 & new_n346;
  assign new_n348 = ~n90 & ~new_n346;
  assign n81 = ~new_n347 & ~new_n348;
  assign new_n350 = new_n325 & new_n331;
  assign new_n351 = new_n309 & new_n350;
  assign new_n352 = n196 & ~new_n351;
  assign new_n353 = ~n196 & new_n351;
  assign n86 = new_n352 | new_n353;
  assign new_n355 = new_n324 & new_n340;
  assign new_n356 = new_n148 & new_n355;
  assign new_n357 = n107 & ~new_n356;
  assign new_n358 = ~n107 & new_n356;
  assign n88 = new_n357 | new_n358;
  assign new_n360 = new_n302 & new_n324;
  assign new_n361 = new_n333 & new_n360;
  assign new_n362 = n43 & ~new_n361;
  assign new_n363 = ~n43 & new_n361;
  assign n89 = new_n362 | new_n363;
  assign new_n365 = new_n323 & new_n335;
  assign new_n366 = n137 & ~new_n365;
  assign new_n367 = ~n137 & new_n365;
  assign n94 = new_n366 | new_n367;
  assign new_n369 = new_n148 & new_n332;
  assign new_n370 = new_n331 & new_n369;
  assign new_n371 = new_n309 & new_n370;
  assign new_n372 = n27 & ~new_n371;
  assign new_n373 = ~n27 & new_n371;
  assign n98 = new_n372 | new_n373;
  assign new_n375 = new_n310_1 & new_n324;
  assign new_n376 = new_n148 & new_n375;
  assign new_n377 = n289 & ~new_n376;
  assign new_n378 = ~n289 & new_n376;
  assign n104 = new_n377 | new_n378;
  assign new_n380 = new_n262 & new_n369;
  assign new_n381 = new_n309 & new_n380;
  assign new_n382 = ~n211 & ~new_n381;
  assign new_n383 = n211 & new_n381;
  assign n123 = ~new_n382 & ~new_n383;
  assign new_n385 = new_n301 & new_n331;
  assign new_n386 = new_n187_1 & new_n385;
  assign new_n387 = new_n148 & new_n386;
  assign new_n388 = n210 & ~new_n387;
  assign new_n389 = ~n210 & new_n387;
  assign n129 = new_n388 | new_n389;
  assign new_n391 = new_n317 & new_n331;
  assign new_n392 = new_n323 & new_n391;
  assign new_n393 = ~n278 & ~new_n392;
  assign new_n394 = n278 & new_n392;
  assign n145 = ~new_n393 & ~new_n394;
  assign new_n396 = new_n309 & new_n391;
  assign new_n397 = n234 & ~new_n396;
  assign new_n398 = ~n234 & new_n396;
  assign n151 = new_n397 | new_n398;
  assign new_n400 = new_n333 & new_n341;
  assign new_n401 = ~n70 & ~new_n400;
  assign new_n402 = n70 & new_n400;
  assign n160 = ~new_n401 & ~new_n402;
  assign new_n404 = new_n311 & new_n333;
  assign new_n405 = n2 & new_n404;
  assign new_n406 = ~n2 & ~new_n404;
  assign n164 = ~new_n405 & ~new_n406;
  assign new_n408 = new_n333 & new_n355;
  assign new_n409 = ~n130 & ~new_n408;
  assign new_n410 = n130 & new_n408;
  assign n168 = ~new_n409 & ~new_n410;
  assign new_n412 = new_n323 & new_n380;
  assign new_n413 = ~n187 & ~new_n412;
  assign new_n414 = n187 & new_n412;
  assign n199 = ~new_n413 & ~new_n414;
  assign new_n416 = new_n324 & new_n385;
  assign new_n417 = new_n333 & new_n416;
  assign new_n418 = ~n23 & ~new_n417;
  assign new_n419 = n23 & new_n417;
  assign n212 = ~new_n418 & ~new_n419;
  assign new_n421 = new_n309 & new_n326;
  assign new_n422 = ~n75 & ~new_n421;
  assign new_n423 = n75 & new_n421;
  assign n213 = ~new_n422 & ~new_n423;
  assign new_n425 = new_n333 & new_n375;
  assign new_n426 = n256 & new_n425;
  assign new_n427 = ~n256 & ~new_n425;
  assign n217 = ~new_n426 & ~new_n427;
  assign new_n429 = new_n262 & new_n334;
  assign new_n430 = new_n323 & new_n429;
  assign new_n431 = ~n179 & ~new_n430;
  assign new_n432 = n179 & new_n430;
  assign n221 = ~new_n431 & ~new_n432;
  assign new_n434 = new_n148 & new_n416;
  assign new_n435 = n249 & ~new_n434;
  assign new_n436 = ~n249 & new_n434;
  assign n246 = new_n435 | new_n436;
  assign new_n438 = new_n323 & new_n350;
  assign new_n439 = n272 & ~new_n438;
  assign new_n440 = ~n272 & new_n438;
  assign n253 = new_n439 | new_n440;
  assign new_n442 = new_n309 & new_n429;
  assign new_n443 = ~n0 & ~new_n442;
  assign new_n444 = n0 & new_n442;
  assign n261 = ~new_n443 & ~new_n444;
  assign new_n446 = new_n323 & new_n370;
  assign new_n447 = n194 & ~new_n446;
  assign new_n448 = ~n194 & new_n446;
  assign n265 = new_n447 | new_n448;
  assign new_n450 = new_n318 & new_n323;
  assign new_n451 = n238 & new_n450;
  assign new_n452 = ~n238 & ~new_n450;
  assign n286 = ~new_n451 & ~new_n452;
  assign new_n454 = new_n148 & new_n360;
  assign new_n455 = n214 & ~new_n454;
  assign new_n456 = ~n214 & new_n454;
  assign n304 = new_n455 | new_n456;
  assign new_n458 = new_n333 & new_n386;
  assign new_n459 = ~n237 & ~new_n458;
  assign new_n460 = n237 & new_n458;
  assign n310 = ~new_n459 & ~new_n460;
endmodule


