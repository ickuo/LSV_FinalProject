// Benchmark "top" written by ABC on Sun Dec 21 18:06:00 2025

module top ( 
    n1, n4, n15, n21, n23, n28, n37, n38, n45, n52, n53, n60, n75, n79,
    n83, n87, n95, n105, n114, n117, n122, n152, n155, n160, n162, n168,
    n183, n187, n194, n198, n206, n215, n218, n227, n228, n231, n242, n269,
    n276, n278, n280,
    n3, n32, n40, n47, n50, n54, n72, n81, n86, n91, n97, n99, n111, n139,
    n154, n176, n185, n191, n197, n200, n205, n208, n211, n214, n220, n243,
    n248, n254, n262, n265, n273, n283  );
  input  n1, n4, n15, n21, n23, n28, n37, n38, n45, n52, n53, n60, n75,
    n79, n83, n87, n95, n105, n114, n117, n122, n152, n155, n160, n162,
    n168, n183, n187, n194, n198, n206, n215, n218, n227, n228, n231, n242,
    n269, n276, n278, n280;
  output n3, n32, n40, n47, n50, n54, n72, n81, n86, n91, n97, n99, n111,
    n139, n154, n176, n185, n191, n197, n200, n205, n208, n211, n214, n220,
    n243, n248, n254, n262, n265, n273, n283;
  wire new_n74, new_n75_1, new_n76, new_n77, new_n78, new_n79_1, new_n80,
    new_n81_1, new_n82, new_n83_1, new_n84, new_n85, new_n86_1, new_n87_1,
    new_n88, new_n89, new_n90, new_n91_1, new_n92, new_n93, new_n94,
    new_n95_1, new_n96, new_n97_1, new_n98, new_n99_1, new_n100, new_n101,
    new_n102, new_n103, new_n104, new_n105_1, new_n106, new_n107, new_n108,
    new_n109, new_n110, new_n111_1, new_n112, new_n113, new_n114_1,
    new_n115, new_n116, new_n117_1, new_n118, new_n119, new_n120, new_n121,
    new_n122_1, new_n123, new_n124, new_n125, new_n126, new_n127, new_n128,
    new_n129, new_n130, new_n131, new_n132, new_n133, new_n134, new_n135,
    new_n136, new_n137, new_n138, new_n139_1, new_n140, new_n141, new_n142,
    new_n143, new_n144, new_n145, new_n146, new_n147, new_n148, new_n149,
    new_n150, new_n151, new_n152_1, new_n153, new_n154_1, new_n155_1,
    new_n156, new_n157, new_n158, new_n159, new_n160_1, new_n161,
    new_n162_1, new_n163, new_n164, new_n165, new_n166, new_n167,
    new_n168_1, new_n169, new_n170, new_n171, new_n172, new_n173, new_n174,
    new_n175, new_n176_1, new_n177, new_n178, new_n179, new_n180, new_n181,
    new_n182, new_n183_1, new_n184, new_n185_1, new_n186, new_n187_1,
    new_n188, new_n189, new_n190, new_n191_1, new_n192, new_n193,
    new_n194_1, new_n195, new_n196, new_n197_1, new_n198_1, new_n199,
    new_n200_1, new_n201, new_n202, new_n203, new_n204, new_n205_1,
    new_n206_1, new_n207, new_n208_1, new_n209, new_n210, new_n211_1,
    new_n212, new_n213, new_n214_1, new_n215_1, new_n216, new_n217,
    new_n218_1, new_n219, new_n220_1, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227_1, new_n228_1, new_n229,
    new_n230, new_n231_1, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242_1,
    new_n243_1, new_n244, new_n245, new_n246, new_n247, new_n248_1,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254_1, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262_1,
    new_n263, new_n264, new_n265_1, new_n266, new_n267, new_n268,
    new_n269_1, new_n270, new_n271, new_n272, new_n273_1, new_n274,
    new_n275, new_n276_1, new_n277, new_n278_1, new_n279, new_n280_1,
    new_n281, new_n282, new_n283_1, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n308, new_n309,
    new_n310, new_n311, new_n312, new_n313, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n324, new_n325,
    new_n326, new_n327, new_n328, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n343, new_n344, new_n345, new_n346, new_n347, new_n348, new_n349,
    new_n351, new_n352, new_n353, new_n354, new_n355, new_n357, new_n358,
    new_n359, new_n361, new_n362, new_n363, new_n364, new_n366, new_n367,
    new_n368, new_n369, new_n370, new_n372, new_n373, new_n374, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n382, new_n383, new_n384,
    new_n386, new_n387, new_n388, new_n390, new_n391, new_n392, new_n393,
    new_n395, new_n396, new_n397, new_n399, new_n400, new_n401, new_n402,
    new_n404, new_n405, new_n406, new_n408, new_n409, new_n410, new_n412,
    new_n413, new_n414, new_n415, new_n417, new_n418, new_n419, new_n421,
    new_n422, new_n423, new_n425, new_n426, new_n427, new_n429, new_n430,
    new_n431, new_n433, new_n434, new_n435, new_n437, new_n438, new_n439,
    new_n441, new_n442, new_n443, new_n445, new_n446, new_n447, new_n449,
    new_n450, new_n451, new_n453, new_n454, new_n455, new_n457, new_n458,
    new_n459;
  assign new_n74 = ~n194 & n280;
  assign new_n75_1 = n194 & ~n280;
  assign new_n76 = ~new_n74 & ~new_n75_1;
  assign new_n77 = n21 & n37;
  assign new_n78 = ~n21 & ~n37;
  assign new_n79_1 = ~new_n77 & ~new_n78;
  assign new_n80 = new_n76 & new_n79_1;
  assign new_n81_1 = ~new_n76 & ~new_n79_1;
  assign new_n82 = ~new_n80 & ~new_n81_1;
  assign new_n83_1 = ~n122 & n276;
  assign new_n84 = n122 & ~n276;
  assign new_n85 = ~new_n83_1 & ~new_n84;
  assign new_n86_1 = n75 & n79;
  assign new_n87_1 = ~n75 & ~n79;
  assign new_n88 = ~new_n86_1 & ~new_n87_1;
  assign new_n89 = ~new_n85 & new_n88;
  assign new_n90 = new_n85 & ~new_n88;
  assign new_n91_1 = ~new_n89 & ~new_n90;
  assign new_n92 = ~new_n82 & new_n91_1;
  assign new_n93 = new_n82 & ~new_n91_1;
  assign new_n94 = ~new_n92 & ~new_n93;
  assign new_n95_1 = n4 & n60;
  assign new_n96 = ~n160 & n227;
  assign new_n97_1 = n160 & ~n227;
  assign new_n98 = ~new_n96 & ~new_n97_1;
  assign new_n99_1 = n105 & n152;
  assign new_n100 = ~n105 & ~n152;
  assign new_n101 = ~new_n99_1 & ~new_n100;
  assign new_n102 = new_n98 & new_n101;
  assign new_n103 = ~new_n98 & ~new_n101;
  assign new_n104 = ~new_n102 & ~new_n103;
  assign new_n105_1 = new_n95_1 & new_n104;
  assign new_n106 = ~new_n95_1 & ~new_n104;
  assign new_n107 = ~new_n105_1 & ~new_n106;
  assign new_n108 = new_n94 & new_n107;
  assign new_n109 = ~new_n94 & ~new_n107;
  assign new_n110 = ~new_n108 & ~new_n109;
  assign new_n111_1 = n4 & n198;
  assign new_n112 = ~new_n104 & ~new_n111_1;
  assign new_n113 = new_n104 & new_n111_1;
  assign new_n114_1 = ~new_n112 & ~new_n113;
  assign new_n115 = ~n83 & n155;
  assign new_n116 = n83 & ~n155;
  assign new_n117_1 = ~new_n115 & ~new_n116;
  assign new_n118 = n23 & n53;
  assign new_n119 = ~n23 & ~n53;
  assign new_n120 = ~new_n118 & ~new_n119;
  assign new_n121 = new_n117_1 & new_n120;
  assign new_n122_1 = ~new_n117_1 & ~new_n120;
  assign new_n123 = ~new_n121 & ~new_n122_1;
  assign new_n124 = ~n162 & n215;
  assign new_n125 = n162 & ~n215;
  assign new_n126 = ~new_n124 & ~new_n125;
  assign new_n127 = n15 & n28;
  assign new_n128 = ~n15 & ~n28;
  assign new_n129 = ~new_n127 & ~new_n128;
  assign new_n130 = ~new_n126 & new_n129;
  assign new_n131 = new_n126 & ~new_n129;
  assign new_n132 = ~new_n130 & ~new_n131;
  assign new_n133 = ~new_n123 & new_n132;
  assign new_n134 = new_n123 & ~new_n132;
  assign new_n135 = ~new_n133 & ~new_n134;
  assign new_n136 = new_n114_1 & ~new_n135;
  assign new_n137 = ~new_n114_1 & new_n135;
  assign new_n138 = ~new_n136 & ~new_n137;
  assign new_n139_1 = new_n110 & ~new_n138;
  assign new_n140 = n4 & n114;
  assign new_n141 = ~new_n123 & ~new_n140;
  assign new_n142 = new_n123 & new_n140;
  assign new_n143 = ~new_n141 & ~new_n142;
  assign new_n144 = ~n242 & n278;
  assign new_n145 = n242 & ~n278;
  assign new_n146 = ~new_n144 & ~new_n145;
  assign new_n147 = n52 & n87;
  assign new_n148 = ~n52 & ~n87;
  assign new_n149 = ~new_n147 & ~new_n148;
  assign new_n150 = new_n146 & new_n149;
  assign new_n151 = ~new_n146 & ~new_n149;
  assign new_n152_1 = ~new_n150 & ~new_n151;
  assign new_n153 = ~n187 & n228;
  assign new_n154_1 = n187 & ~n228;
  assign new_n155_1 = ~new_n153 & ~new_n154_1;
  assign new_n156 = n45 & n95;
  assign new_n157 = ~n45 & ~n95;
  assign new_n158 = ~new_n156 & ~new_n157;
  assign new_n159 = ~new_n155_1 & new_n158;
  assign new_n160_1 = new_n155_1 & ~new_n158;
  assign new_n161 = ~new_n159 & ~new_n160_1;
  assign new_n162_1 = ~new_n152_1 & new_n161;
  assign new_n163 = new_n152_1 & ~new_n161;
  assign new_n164 = ~new_n162_1 & ~new_n163;
  assign new_n165 = new_n143 & ~new_n164;
  assign new_n166 = ~new_n143 & new_n164;
  assign new_n167 = ~new_n165 & ~new_n166;
  assign new_n168_1 = new_n139_1 & new_n167;
  assign new_n169 = n4 & n117;
  assign new_n170 = ~n162 & n183;
  assign new_n171 = n162 & ~n183;
  assign new_n172 = ~new_n170 & ~new_n171;
  assign new_n173 = n45 & n75;
  assign new_n174 = ~n45 & ~n75;
  assign new_n175 = ~new_n173 & ~new_n174;
  assign new_n176_1 = new_n172 & new_n175;
  assign new_n177 = ~new_n172 & ~new_n175;
  assign new_n178 = ~new_n176_1 & ~new_n177;
  assign new_n179 = ~new_n169 & ~new_n178;
  assign new_n180 = new_n169 & new_n178;
  assign new_n181 = ~new_n179 & ~new_n180;
  assign new_n182 = ~n206 & n215;
  assign new_n183_1 = n206 & ~n215;
  assign new_n184 = ~new_n182 & ~new_n183_1;
  assign new_n185_1 = n122 & n187;
  assign new_n186 = ~n122 & ~n187;
  assign new_n187_1 = ~new_n185_1 & ~new_n186;
  assign new_n188 = new_n184 & new_n187_1;
  assign new_n189 = ~new_n184 & ~new_n187_1;
  assign new_n190 = ~new_n188 & ~new_n189;
  assign new_n191_1 = ~n194 & n242;
  assign new_n192 = n194 & ~n242;
  assign new_n193 = ~new_n191_1 & ~new_n192;
  assign new_n194_1 = n53 & n105;
  assign new_n195 = ~n53 & ~n105;
  assign new_n196 = ~new_n194_1 & ~new_n195;
  assign new_n197_1 = ~new_n193 & new_n196;
  assign new_n198_1 = new_n193 & ~new_n196;
  assign new_n199 = ~new_n197_1 & ~new_n198_1;
  assign new_n200_1 = ~new_n190 & new_n199;
  assign new_n201 = new_n190 & ~new_n199;
  assign new_n202 = ~new_n200_1 & ~new_n201;
  assign new_n203 = new_n181 & ~new_n202;
  assign new_n204 = ~new_n181 & new_n202;
  assign new_n205_1 = ~new_n203 & ~new_n204;
  assign new_n206_1 = n4 & n269;
  assign new_n207 = ~new_n82 & ~new_n206_1;
  assign new_n208_1 = new_n82 & new_n206_1;
  assign new_n209 = ~new_n207 & ~new_n208_1;
  assign new_n210 = ~n183 & n206;
  assign new_n211_1 = n183 & ~n206;
  assign new_n212 = ~new_n210 & ~new_n211_1;
  assign new_n213 = n1 & n38;
  assign new_n214_1 = ~n1 & ~n38;
  assign new_n215_1 = ~new_n213 & ~new_n214_1;
  assign new_n216 = ~new_n212 & new_n215_1;
  assign new_n217 = new_n212 & ~new_n215_1;
  assign new_n218_1 = ~new_n216 & ~new_n217;
  assign new_n219 = ~new_n152_1 & new_n218_1;
  assign new_n220_1 = new_n152_1 & ~new_n218_1;
  assign new_n221 = ~new_n219 & ~new_n220_1;
  assign new_n222 = new_n209 & ~new_n221;
  assign new_n223 = ~new_n209 & new_n221;
  assign new_n224 = ~new_n222 & ~new_n223;
  assign new_n225 = ~new_n205_1 & new_n224;
  assign new_n226 = ~n83 & n227;
  assign new_n227_1 = n83 & ~n227;
  assign new_n228_1 = ~new_n226 & ~new_n227_1;
  assign new_n229 = n21 & n52;
  assign new_n230 = ~n21 & ~n52;
  assign new_n231_1 = ~new_n229 & ~new_n230;
  assign new_n232 = ~new_n228_1 & new_n231_1;
  assign new_n233 = new_n228_1 & ~new_n231_1;
  assign new_n234 = ~new_n232 & ~new_n233;
  assign new_n235 = ~new_n178 & new_n234;
  assign new_n236 = new_n178 & ~new_n234;
  assign new_n237 = ~new_n235 & ~new_n236;
  assign new_n238 = n4 & n231;
  assign new_n239 = ~n95 & n276;
  assign new_n240 = n95 & ~n276;
  assign new_n241 = ~new_n239 & ~new_n240;
  assign new_n242_1 = n15 & n38;
  assign new_n243_1 = ~n15 & ~n38;
  assign new_n244 = ~new_n242_1 & ~new_n243_1;
  assign new_n245 = new_n241 & new_n244;
  assign new_n246 = ~new_n241 & ~new_n244;
  assign new_n247 = ~new_n245 & ~new_n246;
  assign new_n248_1 = new_n238 & new_n247;
  assign new_n249 = ~new_n238 & ~new_n247;
  assign new_n250 = ~new_n248_1 & ~new_n249;
  assign new_n251 = new_n237 & new_n250;
  assign new_n252 = ~new_n237 & ~new_n250;
  assign new_n253 = ~new_n251 & ~new_n252;
  assign new_n254_1 = n4 & n218;
  assign new_n255 = ~n79 & n228;
  assign new_n256 = n79 & ~n228;
  assign new_n257 = ~new_n255 & ~new_n256;
  assign new_n258 = n1 & n28;
  assign new_n259 = ~n1 & ~n28;
  assign new_n260 = ~new_n258 & ~new_n259;
  assign new_n261 = new_n257 & new_n260;
  assign new_n262_1 = ~new_n257 & ~new_n260;
  assign new_n263 = ~new_n261 & ~new_n262_1;
  assign new_n264 = ~new_n254_1 & new_n263;
  assign new_n265_1 = new_n254_1 & ~new_n263;
  assign new_n266 = ~new_n264 & ~new_n265_1;
  assign new_n267 = ~n278 & n280;
  assign new_n268 = n278 & ~n280;
  assign new_n269_1 = ~new_n267 & ~new_n268;
  assign new_n270 = n23 & n152;
  assign new_n271 = ~n23 & ~n152;
  assign new_n272 = ~new_n270 & ~new_n271;
  assign new_n273_1 = ~new_n269_1 & new_n272;
  assign new_n274 = new_n269_1 & ~new_n272;
  assign new_n275 = ~new_n273_1 & ~new_n274;
  assign new_n276_1 = ~new_n190 & new_n275;
  assign new_n277 = new_n190 & ~new_n275;
  assign new_n278_1 = ~new_n276_1 & ~new_n277;
  assign new_n279 = new_n266 & ~new_n278_1;
  assign new_n280_1 = ~new_n266 & new_n278_1;
  assign new_n281 = ~new_n279 & ~new_n280_1;
  assign new_n282 = new_n253 & ~new_n281;
  assign new_n283_1 = n4 & n168;
  assign new_n284 = ~new_n247 & ~new_n283_1;
  assign new_n285 = new_n247 & new_n283_1;
  assign new_n286 = ~new_n284 & ~new_n285;
  assign new_n287 = ~n155 & n160;
  assign new_n288 = n155 & ~n160;
  assign new_n289 = ~new_n287 & ~new_n288;
  assign new_n290 = n37 & n87;
  assign new_n291 = ~n37 & ~n87;
  assign new_n292 = ~new_n290 & ~new_n291;
  assign new_n293 = ~new_n289 & new_n292;
  assign new_n294 = new_n289 & ~new_n292;
  assign new_n295 = ~new_n293 & ~new_n294;
  assign new_n296 = ~new_n263 & new_n295;
  assign new_n297 = new_n263 & ~new_n295;
  assign new_n298 = ~new_n296 & ~new_n297;
  assign new_n299 = new_n286 & ~new_n298;
  assign new_n300 = ~new_n286 & new_n298;
  assign new_n301 = ~new_n299 & ~new_n300;
  assign new_n302 = new_n282 & ~new_n301;
  assign new_n303 = new_n225 & new_n302;
  assign new_n304 = new_n168_1 & new_n303;
  assign new_n305 = ~n278 & ~new_n304;
  assign new_n306 = n278 & new_n304;
  assign n3 = ~new_n305 & ~new_n306;
  assign new_n308 = ~new_n205_1 & ~new_n224;
  assign new_n309 = new_n301 & new_n308;
  assign new_n310 = new_n282 & new_n309;
  assign new_n311 = new_n168_1 & new_n310;
  assign new_n312 = ~n228 & ~new_n311;
  assign new_n313 = n228 & new_n311;
  assign n32 = ~new_n312 & ~new_n313;
  assign new_n315 = ~new_n253 & new_n281;
  assign new_n316 = new_n139_1 & ~new_n167;
  assign new_n317 = new_n205_1 & ~new_n301;
  assign new_n318 = new_n224 & new_n317;
  assign new_n319 = new_n316 & new_n318;
  assign new_n320 = new_n315 & new_n319;
  assign new_n321 = n183 & ~new_n320;
  assign new_n322 = ~n183 & new_n320;
  assign n40 = new_n321 | new_n322;
  assign new_n324 = new_n225 & new_n301;
  assign new_n325 = new_n316 & new_n324;
  assign new_n326 = new_n315 & new_n325;
  assign new_n327 = n38 & ~new_n326;
  assign new_n328 = ~n38 & new_n326;
  assign n47 = new_n327 | new_n328;
  assign new_n330 = new_n253 & new_n281;
  assign new_n331 = new_n324 & new_n330;
  assign new_n332 = new_n168_1 & new_n331;
  assign new_n333 = ~n87 & ~new_n332;
  assign new_n334 = n87 & new_n332;
  assign n50 = ~new_n333 & ~new_n334;
  assign new_n336 = ~new_n110 & ~new_n167;
  assign new_n337 = new_n138 & new_n336;
  assign new_n338 = new_n309 & new_n330;
  assign new_n339 = new_n337 & new_n338;
  assign new_n340 = n160 & ~new_n339;
  assign new_n341 = ~n160 & new_n339;
  assign n54 = new_n340 | new_n341;
  assign new_n343 = new_n110 & new_n138;
  assign new_n344 = ~new_n167 & new_n343;
  assign new_n345 = ~new_n224 & new_n317;
  assign new_n346 = new_n315 & new_n345;
  assign new_n347 = new_n344 & new_n346;
  assign new_n348 = ~n162 & ~new_n347;
  assign new_n349 = n162 & new_n347;
  assign n72 = ~new_n348 & ~new_n349;
  assign new_n351 = ~new_n138 & new_n336;
  assign new_n352 = new_n318 & new_n330;
  assign new_n353 = new_n351 & new_n352;
  assign new_n354 = n194 & ~new_n353;
  assign new_n355 = ~n194 & new_n353;
  assign n81 = new_n354 | new_n355;
  assign new_n357 = new_n331 & new_n351;
  assign new_n358 = n37 & ~new_n357;
  assign new_n359 = ~n37 & new_n357;
  assign n86 = new_n358 | new_n359;
  assign new_n361 = new_n302 & new_n308;
  assign new_n362 = new_n337 & new_n361;
  assign new_n363 = n152 & ~new_n362;
  assign new_n364 = ~n152 & new_n362;
  assign n91 = new_n363 | new_n364;
  assign new_n366 = new_n167 & new_n343;
  assign new_n367 = new_n330 & new_n345;
  assign new_n368 = new_n366 & new_n367;
  assign new_n369 = n53 & new_n368;
  assign new_n370 = ~n53 & ~new_n368;
  assign n97 = ~new_n369 & ~new_n370;
  assign new_n372 = new_n303 & new_n351;
  assign new_n373 = n280 & ~new_n372;
  assign new_n374 = ~n280 & new_n372;
  assign n99 = new_n373 | new_n374;
  assign new_n376 = ~new_n301 & new_n315;
  assign new_n377 = new_n308 & new_n376;
  assign new_n378 = new_n366 & new_n377;
  assign new_n379 = n83 & ~new_n378;
  assign new_n380 = ~n83 & new_n378;
  assign n111 = new_n379 | new_n380;
  assign new_n382 = new_n338 & new_n366;
  assign new_n383 = n155 & ~new_n382;
  assign new_n384 = ~n155 & new_n382;
  assign n139 = new_n383 | new_n384;
  assign new_n386 = new_n282 & new_n319;
  assign new_n387 = n206 & ~new_n386;
  assign new_n388 = ~n206 & new_n386;
  assign n154 = new_n387 | new_n388;
  assign new_n390 = new_n309 & new_n315;
  assign new_n391 = new_n168_1 & new_n390;
  assign new_n392 = ~n95 & ~new_n391;
  assign new_n393 = n95 & new_n391;
  assign n176 = ~new_n392 & ~new_n393;
  assign new_n395 = new_n351 & new_n390;
  assign new_n396 = n276 & ~new_n395;
  assign new_n397 = ~n276 & new_n395;
  assign n185 = new_n396 | new_n397;
  assign new_n399 = new_n282 & new_n345;
  assign new_n400 = new_n344 & new_n399;
  assign new_n401 = ~n215 & ~new_n400;
  assign new_n402 = n215 & new_n400;
  assign n191 = ~new_n401 & ~new_n402;
  assign new_n404 = new_n168_1 & new_n352;
  assign new_n405 = ~n242 & ~new_n404;
  assign new_n406 = n242 & new_n404;
  assign n197 = ~new_n405 & ~new_n406;
  assign new_n408 = new_n361 & new_n366;
  assign new_n409 = n23 & ~new_n408;
  assign new_n410 = ~n23 & new_n408;
  assign n200 = new_n409 | new_n410;
  assign new_n412 = new_n225 & new_n376;
  assign new_n413 = new_n351 & new_n412;
  assign new_n414 = ~n21 & ~new_n413;
  assign new_n415 = n21 & new_n413;
  assign n205 = ~new_n414 & ~new_n415;
  assign new_n417 = new_n168_1 & new_n412;
  assign new_n418 = ~n52 & ~new_n417;
  assign new_n419 = n52 & new_n417;
  assign n208 = ~new_n418 & ~new_n419;
  assign new_n421 = new_n351 & new_n399;
  assign new_n422 = n122 & ~new_n421;
  assign new_n423 = ~n122 & new_n421;
  assign n211 = new_n422 | new_n423;
  assign new_n425 = new_n168_1 & new_n399;
  assign new_n426 = ~n187 & ~new_n425;
  assign new_n427 = n187 & new_n425;
  assign n214 = ~new_n426 & ~new_n427;
  assign new_n429 = new_n337 & new_n377;
  assign new_n430 = ~n227 & ~new_n429;
  assign new_n431 = n227 & new_n429;
  assign n220 = ~new_n430 & ~new_n431;
  assign new_n433 = new_n168_1 & new_n346;
  assign new_n434 = ~n45 & ~new_n433;
  assign new_n435 = n45 & new_n433;
  assign n243 = ~new_n434 & ~new_n435;
  assign new_n437 = new_n344 & new_n390;
  assign new_n438 = n15 & ~new_n437;
  assign new_n439 = ~n15 & new_n437;
  assign n248 = new_n438 | new_n439;
  assign new_n441 = new_n310 & new_n344;
  assign new_n442 = n28 & ~new_n441;
  assign new_n443 = ~n28 & new_n441;
  assign n254 = new_n442 | new_n443;
  assign new_n445 = new_n282 & new_n325;
  assign new_n446 = n1 & ~new_n445;
  assign new_n447 = ~n1 & new_n445;
  assign n262 = new_n446 | new_n447;
  assign new_n449 = new_n310 & new_n351;
  assign new_n450 = n79 & ~new_n449;
  assign new_n451 = ~n79 & new_n449;
  assign n265 = new_n450 | new_n451;
  assign new_n453 = new_n346 & new_n351;
  assign new_n454 = n75 & ~new_n453;
  assign new_n455 = ~n75 & new_n453;
  assign n273 = new_n454 | new_n455;
  assign new_n457 = new_n337 & new_n367;
  assign new_n458 = ~n105 & ~new_n457;
  assign new_n459 = n105 & new_n457;
  assign n283 = ~new_n458 & ~new_n459;
endmodule


