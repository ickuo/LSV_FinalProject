module top( n59 , n74 , n85 , n145 , n161 , n228 , n232 , n272 , n330 , 
n388 , n400 , n402 , n407 , n434 , n435 , n476 , n520 , n579 , n582 , 
n599 , n648 , n653 , n660 , n674 , n676 , n728 , n730 , n757 , n794 , 
n819 , n844 , n881 , n964 , n997 , n1007 , n1055 , n1067 , n1087 , n1117 , 
n1119 , n1123 , n1125 , n1134 , n1183 , n1187 , n1244 , n1271 , n1275 , n1282 , 
n1298 , n1308 , n1367 , n1382 , n1411 , n1428 , n1512 , n1543 , n1588 , n1613 , 
n1660 , n1676 , n1679 , n1692 , n1778 , n1779 , n1806 , n1833 , n1858 , n1900 , 
n1901 , n1904 , n1905 , n1924 , n1948 , n1956 , n1960 , n1970 , n1987 , n2004 , 
n2029 , n2073 , n2157 , n2163 , n2188 , n2192 , n2220 , n2232 , n2301 , n2303 , 
n2310 , n2311 , n2387 , n2408 , n2450 , n2516 , n2521 , n2536 , n2551 , n2567 , 
n2582 , n2586 , n2628 , n2666 , n2673 , n2747 , n2753 , n2801 , n2853 , n2886 , 
n2903 , n2906 , n3034 , n3055 , n3073 , n3105 , n3112 , n3121 , n3141 , n3156 , 
n3238 , n3241 , n3302 , n3329 , n3333 , n3366 , n3413 , n3414 , n3430 , n3439 , 
n3498 , n3529 , n3542 , n3546 , n3566 , n3584 , n3652 , n3659 , n3662 );
    input n59 , n74 , n145 , n161 , n228 , n272 , n330 , n388 , n400 , 
n402 , n407 , n434 , n435 , n476 , n520 , n579 , n582 , n648 , n653 , 
n660 , n674 , n728 , n730 , n757 , n794 , n819 , n844 , n881 , n997 , 
n1055 , n1067 , n1087 , n1117 , n1119 , n1123 , n1125 , n1134 , n1183 , n1187 , 
n1244 , n1271 , n1275 , n1282 , n1298 , n1308 , n1367 , n1382 , n1411 , n1428 , 
n1512 , n1543 , n1588 , n1613 , n1660 , n1676 , n1679 , n1692 , n1778 , n1779 , 
n1806 , n1833 , n1858 , n1900 , n1901 , n1904 , n1905 , n1924 , n1948 , n1956 , 
n1960 , n1970 , n1987 , n2004 , n2029 , n2073 , n2157 , n2163 , n2188 , n2220 , 
n2232 , n2301 , n2303 , n2310 , n2311 , n2387 , n2408 , n2450 , n2516 , n2521 , 
n2536 , n2551 , n2567 , n2582 , n2628 , n2666 , n2753 , n2801 , n2853 , n2906 , 
n3034 , n3073 , n3105 , n3141 , n3156 , n3238 , n3302 , n3329 , n3333 , n3366 , 
n3413 , n3414 , n3430 , n3439 , n3498 , n3529 , n3542 , n3546 , n3566 , n3652 , 
n3659 , n3662 ;
    output n85 , n232 , n599 , n676 , n964 , n1007 , n2192 , n2586 , n2673 , 
n2747 , n2886 , n2903 , n3055 , n3112 , n3121 , n3241 , n3584 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , 
n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , 
n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , 
n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , 
n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , 
n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , 
n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
n70 , n71 , n72 , n73 , n75 , n76 , n77 , n78 , n79 , n80 , 
n81 , n82 , n83 , n84 , n86 , n87 , n88 , n89 , n90 , n91 , 
n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , 
n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , 
n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , 
n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , 
n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , 
n142 , n143 , n144 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , 
n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n162 , n163 , 
n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , 
n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , 
n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , 
n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , 
n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , 
n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , 
n224 , n225 , n226 , n227 , n229 , n230 , n231 , n233 , n234 , n235 , 
n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , 
n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , 
n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , 
n266 , n267 , n268 , n269 , n270 , n271 , n273 , n274 , n275 , n276 , 
n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , 
n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , 
n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
n327 , n328 , n329 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , 
n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , 
n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , 
n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , 
n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , 
n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , 
n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , 
n399 , n401 , n403 , n404 , n405 , n406 , n408 , n409 , n410 , n411 , 
n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , 
n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , 
n432 , n433 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , 
n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , 
n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , 
n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , 
n474 , n475 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , 
n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , 
n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , 
n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , 
n515 , n516 , n517 , n518 , n519 , n521 , n522 , n523 , n524 , n525 , 
n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , 
n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , 
n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , 
n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , 
n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , 
n576 , n577 , n578 , n580 , n581 , n583 , n584 , n585 , n586 , n587 , 
n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , 
n598 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , 
n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , 
n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , 
n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , 
n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n649 , 
n650 , n651 , n652 , n654 , n655 , n656 , n657 , n658 , n659 , n661 , 
n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , 
n672 , n673 , n675 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , 
n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , 
n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , 
n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , 
n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , 
n724 , n725 , n726 , n727 , n729 , n731 , n732 , n733 , n734 , n735 , 
n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , 
n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , 
n756 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , 
n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , 
n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , 
n787 , n788 , n789 , n790 , n791 , n792 , n793 , n795 , n796 , n797 , 
n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , 
n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , 
n818 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , 
n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , 
n839 , n840 , n841 , n842 , n843 , n845 , n846 , n847 , n848 , n849 , 
n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
n880 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , 
n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , 
n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , 
n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , 
n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , 
n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , 
n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , 
n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , 
n961 , n962 , n963 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , 
n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , 
n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , 
n992 , n993 , n994 , n995 , n996 , n998 , n999 , n1000 , n1001 , n1002 , 
n1003 , n1004 , n1005 , n1006 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , 
n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , 
n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , 
n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , 
n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , 
n1054 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , 
n1065 , n1066 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , 
n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , 
n1086 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , 
n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , 
n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , 
n1118 , n1120 , n1121 , n1122 , n1124 , n1126 , n1127 , n1128 , n1129 , n1130 , 
n1131 , n1132 , n1133 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , 
n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , 
n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , 
n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , 
n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , 
n1182 , n1184 , n1185 , n1186 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , 
n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , 
n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , 
n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , 
n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , 
n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , 
n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , 
n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , 
n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1272 , n1273 , n1274 , n1276 , 
n1277 , n1278 , n1279 , n1280 , n1281 , n1283 , n1284 , n1285 , n1286 , n1287 , 
n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , 
n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1309 , 
n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1368 , n1369 , n1370 , 
n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , 
n1381 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , 
n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , 
n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1412 , 
n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , 
n1423 , n1424 , n1425 , n1426 , n1427 , n1429 , n1430 , n1431 , n1432 , n1433 , 
n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , 
n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , 
n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , 
n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , 
n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , 
n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , 
n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , 
n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1513 , n1514 , 
n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , 
n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , 
n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1544 , n1545 , 
n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , 
n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , 
n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , 
n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , 
n1586 , n1587 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , 
n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , 
n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1614 , n1615 , n1616 , n1617 , 
n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , 
n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , 
n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , 
n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , 
n1658 , n1659 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , 
n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1677 , n1678 , n1680 , 
n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , 
n1691 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , 
n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , 
n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , 
n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , 
n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , 
n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , 
n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , 
n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , 
n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1780 , n1781 , n1782 , n1783 , 
n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , 
n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , 
n1804 , n1805 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , 
n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , 
n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1834 , n1835 , 
n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , 
n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , 
n1856 , n1857 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , 
n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , 
n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , 
n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , 
n1897 , n1898 , n1899 , n1902 , n1903 , n1906 , n1907 , n1908 , n1909 , n1910 , 
n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , 
n1921 , n1922 , n1923 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , 
n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , 
n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1949 , n1950 , n1951 , n1952 , 
n1953 , n1954 , n1955 , n1957 , n1958 , n1959 , n1961 , n1962 , n1963 , n1964 , 
n1965 , n1966 , n1967 , n1968 , n1969 , n1971 , n1972 , n1973 , n1974 , n1975 , 
n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , 
n1986 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , 
n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2005 , n2006 , n2007 , 
n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , 
n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , 
n2028 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , 
n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , 
n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , 
n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , 
n2069 , n2070 , n2071 , n2072 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2158 , n2159 , n2160 , 
n2161 , n2162 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , 
n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , 
n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2189 , n2190 , n2191 , n2193 , 
n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , 
n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , 
n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2221 , n2222 , n2223 , n2224 , 
n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2233 , n2234 , n2235 , 
n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , 
n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , 
n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , 
n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , 
n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , 
n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , 
n2296 , n2297 , n2298 , n2299 , n2300 , n2302 , n2304 , n2305 , n2306 , n2307 , 
n2308 , n2309 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2388 , n2389 , n2390 , 
n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2409 , n2410 , n2411 , 
n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , 
n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , 
n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , 
n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2451 , n2452 , 
n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , 
n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , 
n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , 
n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , 
n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , 
n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , 
n2513 , n2514 , n2515 , n2517 , n2518 , n2519 , n2520 , n2522 , n2523 , n2524 , 
n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , 
n2535 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , 
n2546 , n2547 , n2548 , n2549 , n2550 , n2552 , n2553 , n2554 , n2555 , n2556 , 
n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , 
n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , 
n2578 , n2579 , n2580 , n2581 , n2583 , n2584 , n2585 , n2587 , n2588 , n2589 , 
n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2629 , n2630 , 
n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , 
n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , 
n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
n2661 , n2662 , n2663 , n2664 , n2665 , n2667 , n2668 , n2669 , n2670 , n2671 , 
n2672 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , 
n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , 
n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , 
n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , 
n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , 
n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , 
n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , 
n2743 , n2744 , n2745 , n2746 , n2748 , n2749 , n2750 , n2751 , n2752 , n2754 , 
n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , 
n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , 
n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , 
n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , 
n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2802 , n2803 , n2804 , n2805 , 
n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , 
n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , 
n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , 
n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , 
n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2854 , n2855 , n2856 , 
n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , 
n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , 
n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2887 , 
n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , 
n2898 , n2899 , n2900 , n2901 , n2902 , n2904 , n2905 , n2907 , n2908 , n2909 , 
n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
n3030 , n3031 , n3032 , n3033 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , 
n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , 
n3051 , n3052 , n3053 , n3054 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , 
n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , 
n3072 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , 
n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , 
n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , 
n3103 , n3104 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3113 , n3114 , 
n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3122 , n3123 , n3124 , n3125 , 
n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , 
n3136 , n3137 , n3138 , n3139 , n3140 , n3142 , n3143 , n3144 , n3145 , n3146 , 
n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3157 , 
n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , 
n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , 
n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , 
n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , 
n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , 
n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , 
n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , 
n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , 
n3239 , n3240 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
n3300 , n3301 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , 
n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , 
n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3330 , n3331 , 
n3332 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , 
n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , 
n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , 
n3363 , n3364 , n3365 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , 
n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , 
n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , 
n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , 
n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3415 , 
n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , 
n3426 , n3427 , n3428 , n3429 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , 
n3437 , n3438 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , 
n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , 
n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , 
n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , 
n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , 
n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , 
n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , 
n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , 
n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , 
n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
n3540 , n3541 , n3543 , n3544 , n3545 , n3547 , n3548 , n3549 , n3550 , n3551 , 
n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , 
n3562 , n3563 , n3564 , n3565 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , 
n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , 
n3583 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , 
n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , 
n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , 
n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , 
n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , 
n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , 
n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3653 , n3654 , 
n3655 , n3656 , n3657 , n3658 , n3660 , n3661 , n3663 , n3664 , n3665 , n3666 , 
n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , 
n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 ;
    xnor g0 ( n1263 , n465 , n2462 );
    and g1 ( n1723 , n131 , n2185 );
    and g2 ( n1267 , n2204 , n1937 );
    xnor g3 ( n2164 , n2619 , n831 );
    not g4 ( n3417 , n2157 );
    not g5 ( n1716 , n2481 );
    or g6 ( n3544 , n2429 , n840 );
    and g7 ( n1699 , n614 , n622 );
    xor g8 ( n1133 , n2773 , n301 );
    or g9 ( n355 , n2062 , n1396 );
    xnor g10 ( n42 , n661 , n1376 );
    or g11 ( n1409 , n3446 , n2963 );
    xnor g12 ( n1196 , n2947 , n3462 );
    or g13 ( n1105 , n1499 , n1587 );
    or g14 ( n3245 , n726 , n2329 );
    xnor g15 ( n3650 , n824 , n99 );
    xnor g16 ( n3459 , n1978 , n1106 );
    or g17 ( n1830 , n487 , n554 );
    not g18 ( n1509 , n2516 );
    or g19 ( n1867 , n3093 , n2102 );
    nor g20 ( n1018 , n1070 , n2344 );
    not g21 ( n441 , n1858 );
    xnor g22 ( n1483 , n3174 , n3609 );
    and g23 ( n1001 , n1755 , n1472 );
    not g24 ( n1746 , n3225 );
    and g25 ( n1727 , n246 , n3435 );
    and g26 ( n262 , n2267 , n1830 );
    and g27 ( n966 , n1702 , n2087 );
    and g28 ( n336 , n1375 , n1894 );
    and g29 ( n886 , n6 , n2068 );
    or g30 ( n195 , n1887 , n220 );
    or g31 ( n2391 , n2449 , n3450 );
    or g32 ( n1374 , n3332 , n387 );
    xnor g33 ( n2786 , n543 , n377 );
    xnor g34 ( n2464 , n464 , n2885 );
    nor g35 ( n2402 , n2410 , n3442 );
    not g36 ( n2968 , n3414 );
    or g37 ( n2706 , n1052 , n521 );
    xnor g38 ( n1090 , n1366 , n2354 );
    xnor g39 ( n3154 , n2723 , n2752 );
    or g40 ( n2815 , n1987 , n2701 );
    and g41 ( n1591 , n1500 , n346 );
    or g42 ( n2692 , n2535 , n1413 );
    or g43 ( n2456 , n1115 , n2481 );
    xnor g44 ( n1293 , n3144 , n787 );
    or g45 ( n775 , n3028 , n3217 );
    or g46 ( n3438 , n487 , n329 );
    and g47 ( n2361 , n1591 , n247 );
    and g48 ( n2951 , n2301 , n330 );
    or g49 ( n1455 , n2573 , n1861 );
    and g50 ( n2070 , n3223 , n2740 );
    xnor g51 ( n1827 , n3628 , n1893 );
    or g52 ( n2806 , n925 , n453 );
    xnor g53 ( n2970 , n1609 , n1263 );
    xnor g54 ( n2807 , n874 , n3295 );
    and g55 ( n2864 , n2319 , n2167 );
    not g56 ( n3221 , n2042 );
    xnor g57 ( n981 , n1069 , n185 );
    or g58 ( n1057 , n1428 , n1476 );
    xnor g59 ( n2348 , n2800 , n3117 );
    not g60 ( n189 , n435 );
    xor g61 ( n2609 , n314 , n538 );
    or g62 ( n3385 , n957 , n1314 );
    xnor g63 ( n3378 , n148 , n1694 );
    or g64 ( n2530 , n1851 , n2074 );
    xnor g65 ( n3545 , n2297 , n748 );
    and g66 ( n1043 , n3310 , n1242 );
    xnor g67 ( n1675 , n2617 , n2312 );
    xnor g68 ( n3274 , n2829 , n2676 );
    and g69 ( n2638 , n1883 , n1392 );
    or g70 ( n2026 , n23 , n1907 );
    not g71 ( n1144 , n1121 );
    xnor g72 ( n244 , n2263 , n1269 );
    or g73 ( n106 , n1256 , n1515 );
    and g74 ( n3 , n2105 , n80 );
    or g75 ( n733 , n2615 , n1802 );
    and g76 ( n2789 , n1660 , n1055 );
    xnor g77 ( n1605 , n2064 , n30 );
    xnor g78 ( n736 , n2650 , n16 );
    and g79 ( n2007 , n2452 , n2929 );
    nor g80 ( n1268 , n1431 , n3007 );
    and g81 ( n902 , n3666 , n380 );
    or g82 ( n1750 , n1428 , n2153 );
    or g83 ( n2427 , n2617 , n2312 );
    xnor g84 ( n1668 , n1010 , n101 );
    or g85 ( n1886 , n2535 , n2233 );
    and g86 ( n2984 , n817 , n2277 );
    and g87 ( n3167 , n1646 , n2373 );
    and g88 ( n1249 , n1429 , n113 );
    and g89 ( n3503 , n806 , n1370 );
    or g90 ( n3619 , n1405 , n2397 );
    or g91 ( n1480 , n362 , n513 );
    or g92 ( n2566 , n412 , n3682 );
    and g93 ( n792 , n1913 , n711 );
    not g94 ( n2589 , n2823 );
    xnor g95 ( n2193 , n600 , n1014 );
    nor g96 ( n1358 , n3247 , n2095 );
    or g97 ( n2708 , n615 , n146 );
    or g98 ( n888 , n1361 , n331 );
    xnor g99 ( n3109 , n2041 , n1749 );
    or g100 ( n2927 , n2753 , n2225 );
    xnor g101 ( n412 , n3099 , n3076 );
    or g102 ( n3296 , n3550 , n955 );
    or g103 ( n2629 , n3268 , n1228 );
    or g104 ( n1417 , n2569 , n220 );
    or g105 ( n2895 , n1596 , n18 );
    xnor g106 ( n1027 , n3178 , n3383 );
    xnor g107 ( n1478 , n2009 , n2122 );
    xnor g108 ( n1861 , n2062 , n1383 );
    or g109 ( n3435 , n1774 , n89 );
    xnor g110 ( n3206 , n2979 , n1715 );
    or g111 ( n1704 , n3415 , n431 );
    xnor g112 ( n245 , n3032 , n1953 );
    xnor g113 ( n2538 , n1856 , n2782 );
    and g114 ( n341 , n3222 , n721 );
    xnor g115 ( n1651 , n3002 , n1818 );
    or g116 ( n2255 , n1871 , n1413 );
    or g117 ( n1434 , n3441 , n1687 );
    or g118 ( n2269 , n1388 , n3626 );
    not g119 ( n3326 , n1244 );
    and g120 ( n3672 , n486 , n2135 );
    and g121 ( n1468 , n646 , n1850 );
    or g122 ( n3374 , n2956 , n41 );
    or g123 ( n3364 , n2362 , n3275 );
    or g124 ( n1094 , n2236 , n970 );
    or g125 ( n3015 , n1073 , n2294 );
    or g126 ( n3533 , n1144 , n3589 );
    not g127 ( n3335 , n559 );
    and g128 ( n271 , n1639 , n625 );
    or g129 ( n3018 , n561 , n1421 );
    or g130 ( n2312 , n1596 , n1235 );
    not g131 ( n3229 , n1439 );
    xnor g132 ( n2639 , n1336 , n2978 );
    nor g133 ( n2834 , n198 , n765 );
    xnor g134 ( n3151 , n2089 , n167 );
    or g135 ( n369 , n2753 , n254 );
    or g136 ( n421 , n633 , n1961 );
    xnor g137 ( n2561 , n1547 , n1486 );
    xnor g138 ( n2552 , n3619 , n780 );
    not g139 ( n498 , n2287 );
    or g140 ( n1525 , n2569 , n2010 );
    not g141 ( n1129 , n3219 );
    or g142 ( n105 , n2267 , n1830 );
    xnor g143 ( n2747 , n2657 , n672 );
    not g144 ( n2571 , n2273 );
    or g145 ( n1086 , n2616 , n1300 );
    and g146 ( n3279 , n1299 , n52 );
    not g147 ( n3293 , n434 );
    and g148 ( n780 , n2368 , n3512 );
    or g149 ( n3211 , n1744 , n1669 );
    not g150 ( n3009 , n736 );
    or g151 ( n3523 , n925 , n3267 );
    and g152 ( n1228 , n1081 , n2065 );
    or g153 ( n1394 , n2457 , n1555 );
    or g154 ( n1114 , n1586 , n2701 );
    xnor g155 ( n431 , n2966 , n159 );
    or g156 ( n903 , n2112 , n315 );
    or g157 ( n2746 , n3621 , n1427 );
    nor g158 ( n2040 , n1954 , n2857 );
    or g159 ( n474 , n1135 , n1822 );
    and g160 ( n1583 , n1798 , n3132 );
    or g161 ( n2703 , n588 , n2822 );
    or g162 ( n1163 , n3417 , n1707 );
    not g163 ( n372 , n1994 );
    and g164 ( n116 , n1670 , n2887 );
    and g165 ( n782 , n1882 , n809 );
    or g166 ( n3656 , n1785 , n2543 );
    and g167 ( n923 , n12 , n194 );
    xnor g168 ( n1671 , n2769 , n217 );
    and g169 ( n2583 , n3506 , n795 );
    xnor g170 ( n169 , n2371 , n1690 );
    or g171 ( n112 , n3646 , n282 );
    not g172 ( n2108 , n526 );
    xnor g173 ( n3487 , n1489 , n3483 );
    not g174 ( n787 , n297 );
    not g175 ( n1992 , n2188 );
    or g176 ( n3369 , n2697 , n1381 );
    xnor g177 ( n1489 , n2813 , n384 );
    or g178 ( n1287 , n1520 , n1377 );
    or g179 ( n191 , n1552 , n453 );
    or g180 ( n3400 , n3581 , n2537 );
    xnor g181 ( n1974 , n251 , n2472 );
    and g182 ( n2687 , n208 , n1156 );
    and g183 ( n403 , n1187 , n407 );
    or g184 ( n1909 , n2163 , n2870 );
    or g185 ( n868 , n1170 , n445 );
    and g186 ( n2208 , n1858 , n730 );
    xnor g187 ( n2503 , n901 , n1567 );
    not g188 ( n3633 , n3146 );
    and g189 ( n3224 , n2098 , n1597 );
    xnor g190 ( n3127 , n2084 , n357 );
    or g191 ( n102 , n2509 , n1019 );
    and g192 ( n383 , n2950 , n1329 );
    or g193 ( n385 , n2163 , n2162 );
    not g194 ( n3428 , n2370 );
    not g195 ( n2517 , n1298 );
    or g196 ( n909 , n3460 , n2077 );
    nor g197 ( n2884 , n467 , n2394 );
    xnor g198 ( n455 , n1387 , n3209 );
    or g199 ( n1081 , n1216 , n149 );
    or g200 ( n449 , n1632 , n1619 );
    or g201 ( n291 , n700 , n1437 );
    or g202 ( n321 , n751 , n195 );
    not g203 ( n2707 , n807 );
    or g204 ( n908 , n942 , n690 );
    or g205 ( n1364 , n1170 , n649 );
    and g206 ( n2636 , n753 , n2476 );
    nor g207 ( n3370 , n2257 , n158 );
    and g208 ( n1028 , n3629 , n3097 );
    nor g209 ( n1229 , n1111 , n3377 );
    and g210 ( n632 , n2286 , n25 );
    not g211 ( n2768 , n912 );
    and g212 ( n6 , n3325 , n1703 );
    and g213 ( n3660 , n1884 , n1823 );
    xnor g214 ( n3112 , n1881 , n754 );
    nor g215 ( n3437 , n544 , n3346 );
    or g216 ( n684 , n2389 , n2076 );
    and g217 ( n3045 , n318 , n2890 );
    and g218 ( n2610 , n2388 , n171 );
    or g219 ( n772 , n791 , n71 );
    or g220 ( n975 , n1987 , n1950 );
    or g221 ( n2240 , n1887 , n645 );
    and g222 ( n3303 , n1448 , n3635 );
    xor g223 ( n921 , n587 , n3291 );
    xnor g224 ( n3527 , n1300 , n2616 );
    and g225 ( n1349 , n2249 , n804 );
    or g226 ( n3622 , n3370 , n3276 );
    or g227 ( n2098 , n1211 , n2015 );
    and g228 ( n3587 , n908 , n2336 );
    or g229 ( n751 , n1054 , n3318 );
    or g230 ( n1595 , n204 , n1658 );
    not g231 ( n2399 , n1078 );
    or g232 ( n1702 , n3248 , n1243 );
    or g233 ( n694 , n1953 , n2731 );
    xnor g234 ( n2159 , n2331 , n827 );
    or g235 ( n1639 , n3096 , n955 );
    xnor g236 ( n1432 , n2525 , n1725 );
    and g237 ( n280 , n480 , n1816 );
    and g238 ( n1811 , n2609 , n3284 );
    or g239 ( n3421 , n173 , n1235 );
    nor g240 ( n3092 , n3395 , n2104 );
    or g241 ( n1281 , n2081 , n1468 );
    xnor g242 ( n2277 , n3339 , n508 );
    xnor g243 ( n2847 , n2721 , n650 );
    xnor g244 ( n2132 , n3488 , n127 );
    and g245 ( n3040 , n133 , n2761 );
    and g246 ( n1621 , n942 , n690 );
    or g247 ( n1717 , n2553 , n2968 );
    nor g248 ( n3654 , n2321 , n2049 );
    xnor g249 ( n516 , n2702 , n3457 );
    xnor g250 ( n1686 , n1267 , n2155 );
    and g251 ( n3564 , n3479 , n2308 );
    not g252 ( n363 , n672 );
    and g253 ( n1376 , n1401 , n3317 );
    xnor g254 ( n1451 , n1710 , n2799 );
    nor g255 ( n1115 , n2908 , n2415 );
    xnor g256 ( n3356 , n621 , n3052 );
    and g257 ( n1377 , n2966 , n1807 );
    nor g258 ( n2083 , n202 , n2055 );
    or g259 ( n1101 , n2753 , n1145 );
    or g260 ( n1020 , n636 , n1876 );
    or g261 ( n2560 , n555 , n1461 );
    or g262 ( n1714 , n2819 , n2010 );
    or g263 ( n61 , n3468 , n2006 );
    xnor g264 ( n1748 , n1885 , n3610 );
    xnor g265 ( n159 , n1807 , n1520 );
    or g266 ( n1039 , n1428 , n3560 );
    or g267 ( n3005 , n1248 , n306 );
    or g268 ( n2907 , n988 , n2431 );
    and g269 ( n638 , n736 , n2370 );
    xnor g270 ( n3628 , n752 , n319 );
    xor g271 ( n3636 , n2729 , n1539 );
    and g272 ( n3257 , n373 , n951 );
    or g273 ( n3605 , n2096 , n3267 );
    xnor g274 ( n265 , n3494 , n1082 );
    or g275 ( n3122 , n3096 , n34 );
    or g276 ( n3218 , n778 , n3482 );
    and g277 ( n2496 , n1756 , n47 );
    not g278 ( n1795 , n569 );
    or g279 ( n2207 , n1222 , n2137 );
    or g280 ( n2379 , n2220 , n2912 );
    not g281 ( n1413 , n1956 );
    xnor g282 ( n30 , n2600 , n522 );
    or g283 ( n2675 , n2290 , n1986 );
    or g284 ( n1594 , n3271 , n1891 );
    xnor g285 ( n2216 , n94 , n3445 );
    not g286 ( n1205 , n1906 );
    or g287 ( n2376 , n128 , n2186 );
    and g288 ( n829 , n1213 , n909 );
    not g289 ( n2459 , n1765 );
    not g290 ( n3520 , n3383 );
    or g291 ( n2299 , n2465 , n2244 );
    xnor g292 ( n2455 , n54 , n1808 );
    or g293 ( n480 , n3334 , n3368 );
    or g294 ( n1674 , n173 , n1921 );
    or g295 ( n1885 , n1540 , n3152 );
    and g296 ( n591 , n3441 , n1687 );
    or g297 ( n269 , n540 , n1489 );
    xnor g298 ( n2351 , n1566 , n1148 );
    not g299 ( n2705 , n1670 );
    or g300 ( n2961 , n2059 , n347 );
    xnor g301 ( n276 , n3298 , n102 );
    or g302 ( n615 , n2648 , n1015 );
    and g303 ( n1541 , n398 , n2460 );
    or g304 ( n1657 , n251 , n2720 );
    xnor g305 ( n706 , n3492 , n2755 );
    and g306 ( n1070 , n223 , n2997 );
    or g307 ( n3286 , n173 , n189 );
    or g308 ( n2172 , n1784 , n79 );
    nor g309 ( n2620 , n1611 , n1583 );
    xnor g310 ( n307 , n2518 , n1036 );
    or g311 ( n738 , n1926 , n1110 );
    not g312 ( n46 , n3351 );
    or g313 ( n132 , n2291 , n1334 );
    and g314 ( n2949 , n779 , n1022 );
    and g315 ( n1504 , n1604 , n1826 );
    or g316 ( n354 , n2163 , n3480 );
    not g317 ( n2201 , n820 );
    and g318 ( n2426 , n1843 , n2094 );
    xnor g319 ( n3042 , n2532 , n399 );
    xnor g320 ( n326 , n3129 , n3172 );
    xnor g321 ( n3277 , n1316 , n598 );
    or g322 ( n689 , n3243 , n780 );
    and g323 ( n313 , n1928 , n26 );
    xnor g324 ( n232 , n2907 , n1839 );
    and g325 ( n1953 , n1208 , n57 );
    and g326 ( n436 , n1301 , n1630 );
    or g327 ( n3418 , n3202 , n18 );
    and g328 ( n1023 , n969 , n542 );
    or g329 ( n1157 , n1946 , n1149 );
    and g330 ( n1642 , n1435 , n1610 );
    xnor g331 ( n472 , n356 , n833 );
    not g332 ( n173 , n2801 );
    xnor g333 ( n2087 , n2252 , n84 );
    and g334 ( n2161 , n1202 , n3308 );
    or g335 ( n166 , n735 , n32 );
    xnor g336 ( n207 , n2835 , n2719 );
    and g337 ( n1063 , n2611 , n2252 );
    or g338 ( n3027 , n1513 , n1137 );
    and g339 ( n2384 , n1309 , n624 );
    xnor g340 ( n69 , n531 , n3004 );
    or g341 ( n2997 , n196 , n3165 );
    or g342 ( n3317 , n2782 , n67 );
    xnor g343 ( n574 , n440 , n1895 );
    not g344 ( n1898 , n2567 );
    not g345 ( n577 , n274 );
    and g346 ( n837 , n579 , n2906 );
    not g347 ( n3318 , n1779 );
    or g348 ( n887 , n2686 , n3130 );
    xnor g349 ( n662 , n1591 , n756 );
    and g350 ( n2162 , n2305 , n13 );
    or g351 ( n325 , n1084 , n2550 );
    and g352 ( n651 , n924 , n3299 );
    and g353 ( n3131 , n1700 , n2606 );
    or g354 ( n3629 , n2480 , n3496 );
    or g355 ( n3124 , n2213 , n524 );
    not g356 ( n1237 , n2636 );
    and g357 ( n762 , n1284 , n325 );
    or g358 ( n2534 , n1251 , n789 );
    or g359 ( n2191 , n1952 , n2278 );
    not g360 ( n2131 , n1755 );
    and g361 ( n704 , n1172 , n3470 );
    or g362 ( n915 , n3202 , n34 );
    xnor g363 ( n501 , n2958 , n259 );
    xnor g364 ( n1753 , n2365 , n1752 );
    and g365 ( n375 , n3472 , n1936 );
    and g366 ( n1759 , n751 , n195 );
    not g367 ( n1720 , n954 );
    and g368 ( n1210 , n3242 , n3136 );
    or g369 ( n1098 , n3343 , n2848 );
    or g370 ( n3616 , n1792 , n3664 );
    and g371 ( n1989 , n3074 , n693 );
    not g372 ( n1209 , n3145 );
    not g373 ( n2492 , n56 );
    or g374 ( n1464 , n2780 , n420 );
    or g375 ( n3623 , n631 , n163 );
    or g376 ( n1294 , n3094 , n2041 );
    or g377 ( n2957 , n398 , n2460 );
    and g378 ( n505 , n2973 , n2816 );
    or g379 ( n1226 , n1631 , n3267 );
    xnor g380 ( n1712 , n154 , n455 );
    or g381 ( n3501 , n712 , n2251 );
    xnor g382 ( n37 , n3567 , n1976 );
    or g383 ( n2554 , n2163 , n1922 );
    nor g384 ( n9 , n2753 , n2620 );
    or g385 ( n317 , n377 , n2812 );
    or g386 ( n2093 , n154 , n1677 );
    and g387 ( n2591 , n1542 , n630 );
    or g388 ( n2901 , n1405 , n1801 );
    or g389 ( n2067 , n3248 , n1648 );
    and g390 ( n2134 , n394 , n929 );
    and g391 ( n2034 , n1901 , n1117 );
    xnor g392 ( n2229 , n2053 , n1357 );
    or g393 ( n473 , n2772 , n2824 );
    not g394 ( n1805 , n2426 );
    or g395 ( n1392 , n441 , n1648 );
    or g396 ( n3436 , n3645 , n1728 );
    and g397 ( n927 , n2772 , n2824 );
    or g398 ( n3137 , n2895 , n1854 );
    not g399 ( n760 , n2566 );
    or g400 ( n1824 , n38 , n1235 );
    or g401 ( n1188 , n2463 , n3234 );
    xnor g402 ( n3143 , n1435 , n3282 );
    not g403 ( n1707 , n3498 );
    not g404 ( n1617 , n2845 );
    not g405 ( n1015 , n476 );
    xnor g406 ( n3576 , n732 , n2036 );
    or g407 ( n237 , n1569 , n1246 );
    or g408 ( n14 , n2002 , n1398 );
    or g409 ( n188 , n3272 , n1334 );
    or g410 ( n3664 , n1987 , n3500 );
    and g411 ( n764 , n1313 , n1350 );
    and g412 ( n1312 , n1104 , n3393 );
    xnor g413 ( n99 , n182 , n23 );
    or g414 ( n1771 , n2109 , n1714 );
    xnor g415 ( n2885 , n3588 , n3153 );
    or g416 ( n2604 , n1987 , n3644 );
    xnor g417 ( n109 , n2075 , n209 );
    xnor g418 ( n2020 , n2348 , n2470 );
    or g419 ( n2771 , n1166 , n249 );
    not g420 ( n3316 , n238 );
    xnor g421 ( n3170 , n839 , n1437 );
    or g422 ( n631 , n2696 , n955 );
    or g423 ( n3539 , n925 , n1658 );
    and g424 ( n2963 , n2288 , n237 );
    xnor g425 ( n3163 , n589 , n2416 );
    and g426 ( n3062 , n1287 , n1356 );
    or g427 ( n2109 , n457 , n645 );
    and g428 ( n2943 , n1133 , n174 );
    and g429 ( n3562 , n2245 , n2961 );
    xnor g430 ( n1049 , n2015 , n1261 );
    or g431 ( n1633 , n1884 , n1823 );
    or g432 ( n1600 , n2790 , n2846 );
    and g433 ( n1127 , n939 , n3164 );
    or g434 ( n192 , n3455 , n1605 );
    not g435 ( n2236 , n2259 );
    or g436 ( n3115 , n937 , n3641 );
    or g437 ( n290 , n451 , n1060 );
    not g438 ( n3083 , n1335 );
    or g439 ( n3006 , n3398 , n3660 );
    not g440 ( n53 , n1134 );
    xnor g441 ( n3462 , n1231 , n3015 );
    or g442 ( n2637 , n2079 , n2825 );
    and g443 ( n3208 , n2564 , n1237 );
    not g444 ( n2664 , n1117 );
    and g445 ( n553 , n1349 , n2482 );
    not g446 ( n718 , n810 );
    xnor g447 ( n2261 , n2496 , n390 );
    or g448 ( n219 , n457 , n3318 );
    or g449 ( n425 , n1683 , n1171 );
    xnor g450 ( n1612 , n1883 , n1392 );
    or g451 ( n1503 , n2030 , n1138 );
    or g452 ( n3102 , n1372 , n2712 );
    and g453 ( n977 , n1958 , n515 );
    xnor g454 ( n941 , n3562 , n656 );
    or g455 ( n45 , n2946 , n1334 );
    or g456 ( n1000 , n3248 , n1868 );
    and g457 ( n3671 , n2513 , n2708 );
    or g458 ( n1636 , n530 , n1759 );
    and g459 ( n777 , n2544 , n3001 );
    or g460 ( n73 , n82 , n1355 );
    not g461 ( n2186 , n757 );
    xnor g462 ( n1385 , n1395 , n472 );
    or g463 ( n2377 , n910 , n2684 );
    or g464 ( n2656 , n806 , n1370 );
    or g465 ( n1076 , n185 , n1056 );
    nor g466 ( n3410 , n1105 , n3547 );
    nor g467 ( n266 , n1814 , n1015 );
    not g468 ( n1006 , n3576 );
    and g469 ( n2278 , n3600 , n3627 );
    and g470 ( n1207 , n1927 , n1726 );
    or g471 ( n1516 , n1310 , n329 );
    and g472 ( n1785 , n1825 , n1266 );
    or g473 ( n160 , n1307 , n24 );
    xnor g474 ( n122 , n1504 , n2282 );
    xnor g475 ( n3281 , n2284 , n926 );
    or g476 ( n1135 , n3631 , n257 );
    or g477 ( n2227 , n2634 , n3071 );
    not g478 ( n2595 , n1925 );
    xor g479 ( n3106 , n1064 , n181 );
    nor g480 ( n3521 , n1650 , n3424 );
    and g481 ( n255 , n186 , n175 );
    xnor g482 ( n1178 , n2315 , n176 );
    or g483 ( n80 , n1195 , n3103 );
    or g484 ( n1781 , n3394 , n3452 );
    and g485 ( n2966 , n1221 , n180 );
    or g486 ( n769 , n1236 , n2153 );
    not g487 ( n2819 , n1806 );
    or g488 ( n2052 , n3040 , n553 );
    not g489 ( n2971 , n3677 );
    and g490 ( n3358 , n2920 , n2645 );
    or g491 ( n2204 , n3516 , n222 );
    and g492 ( n2322 , n3583 , n1008 );
    or g493 ( n2063 , n3255 , n1334 );
    or g494 ( n617 , n2231 , n2524 );
    or g495 ( n124 , n856 , n1545 );
    xnor g496 ( n1203 , n323 , n1142 );
    and g497 ( n8 , n295 , n1959 );
    or g498 ( n2891 , n2984 , n2488 );
    nor g499 ( n1946 , n1002 , n2424 );
    and g500 ( n1608 , n2419 , n3168 );
    or g501 ( n2723 , n2517 , n3290 );
    not g502 ( n1146 , n147 );
    and g503 ( n767 , n675 , n1188 );
    and g504 ( n3070 , n2944 , n1896 );
    and g505 ( n3392 , n848 , n2771 );
    and g506 ( n2659 , n2662 , n2531 );
    or g507 ( n985 , n2648 , n649 );
    and g508 ( n1403 , n2084 , n357 );
    or g509 ( n1104 , n1165 , n1805 );
    xnor g510 ( n618 , n3205 , n2754 );
    not g511 ( n3228 , n168 );
    xnor g512 ( n251 , n3357 , n1775 );
    and g513 ( n2175 , n2422 , n334 );
    or g514 ( n2782 , n466 , n2397 );
    or g515 ( n558 , n1596 , n955 );
    or g516 ( n497 , n1112 , n111 );
    and g517 ( n1562 , n1711 , n1763 );
    or g518 ( n2421 , n6 , n2068 );
    xnor g519 ( n20 , n3404 , n1820 );
    xnor g520 ( n2041 , n1545 , n3530 );
    xnor g521 ( n3280 , n459 , n863 );
    or g522 ( n2218 , n2833 , n3289 );
    or g523 ( n1131 , n1011 , n1233 );
    or g524 ( n2002 , n3326 , n24 );
    xnor g525 ( n2945 , n2181 , n3487 );
    nor g526 ( n1514 , n1748 , n1892 );
    or g527 ( n3220 , n3255 , n2074 );
    or g528 ( n3639 , n3503 , n3513 );
    and g529 ( n874 , n3077 , n2165 );
    or g530 ( n522 , n2535 , n554 );
    and g531 ( n2420 , n3565 , n302 );
    not g532 ( n3669 , n2724 );
    and g533 ( n3185 , n1773 , n2737 );
    and g534 ( n2870 , n1105 , n3547 );
    not g535 ( n211 , n2226 );
    and g536 ( n755 , n888 , n1418 );
    or g537 ( n41 , n1987 , n2475 );
    not g538 ( n456 , n336 );
    nor g539 ( n815 , n1436 , n3008 );
    or g540 ( n1343 , n1646 , n2373 );
    or g541 ( n2230 , n487 , n2186 );
    and g542 ( n1089 , n2121 , n1739 );
    or g543 ( n3192 , n441 , n1243 );
    or g544 ( n860 , n828 , n2530 );
    or g545 ( n3097 , n865 , n1085 );
    xnor g546 ( n150 , n1941 , n1050 );
    or g547 ( n1825 , n51 , n3361 );
    or g548 ( n66 , n1971 , n3461 );
    or g549 ( n151 , n1533 , n1452 );
    or g550 ( n974 , n716 , n2807 );
    xnor g551 ( n2417 , n1002 , n3100 );
    or g552 ( n1866 , n2993 , n1624 );
    or g553 ( n3216 , n2036 , n732 );
    or g554 ( n3271 , n128 , n554 );
    xnor g555 ( n744 , n1823 , n3088 );
    xnor g556 ( n3033 , n3396 , n811 );
    xnor g557 ( n1366 , n3470 , n2964 );
    and g558 ( n3254 , n502 , n2053 );
    or g559 ( n3451 , n499 , n1454 );
    xnor g560 ( n964 , n3607 , n3042 );
    and g561 ( n1010 , n1563 , n488 );
    and g562 ( n3548 , n698 , n2132 );
    or g563 ( n1415 , n897 , n1707 );
    or g564 ( n108 , n3211 , n3131 );
    or g565 ( n1582 , n1631 , n2968 );
    or g566 ( n439 , n2443 , n2644 );
    or g567 ( n938 , n1435 , n1610 );
    or g568 ( n2173 , n2648 , n2830 );
    or g569 ( n1844 , n1865 , n1930 );
    or g570 ( n3382 , n2850 , n3239 );
    xnor g571 ( n250 , n1727 , n2726 );
    not g572 ( n2413 , n2559 );
    not g573 ( n925 , n1679 );
    or g574 ( n2442 , n1073 , n802 );
    and g575 ( n961 , n1288 , n428 );
    or g576 ( n174 , n1514 , n3478 );
    and g577 ( n2178 , n46 , n2571 );
    or g578 ( n833 , n3615 , n3275 );
    not g579 ( n1524 , n1154 );
    not g580 ( n426 , n285 );
    and g581 ( n2918 , n1547 , n241 );
    or g582 ( n1286 , n487 , n1413 );
    or g583 ( n1471 , n1547 , n241 );
    and g584 ( n1466 , n1985 , n3400 );
    and g585 ( n2665 , n2527 , n2969 );
    and g586 ( n2527 , n3376 , n717 );
    nor g587 ( n2934 , n2691 , n1968 );
    and g588 ( n2225 , n1794 , n3113 );
    or g589 ( n2316 , n1788 , n1754 );
    or g590 ( n3491 , n3272 , n3275 );
    and g591 ( n2526 , n1764 , n135 );
    and g592 ( n3443 , n1869 , n498 );
    not g593 ( n2894 , n3536 );
    and g594 ( n1003 , n1767 , n2333 );
    xnor g595 ( n371 , n3223 , n2992 );
    xnor g596 ( n2892 , n1579 , n603 );
    or g597 ( n898 , n2615 , n2233 );
    or g598 ( n1985 , n2044 , n119 );
    xnor g599 ( n2481 , n1529 , n2976 );
    or g600 ( n123 , n629 , n2765 );
    and g601 ( n2614 , n2284 , n1061 );
    or g602 ( n1345 , n737 , n1627 );
    xnor g603 ( n3390 , n3444 , n1279 );
    or g604 ( n171 , n1725 , n2330 );
    or g605 ( n1777 , n3098 , n396 );
    or g606 ( n2981 , n419 , n2834 );
    or g607 ( n3327 , n945 , n3672 );
    or g608 ( n1773 , n2230 , n11 );
    xnor g609 ( n3003 , n2748 , n1929 );
    or g610 ( n2146 , n2596 , n767 );
    nor g611 ( n252 , n3644 , n1402 );
    or g612 ( n2588 , n1964 , n2381 );
    or g613 ( n2335 , n2445 , n3003 );
    xnor g614 ( n1775 , n3418 , n1554 );
    or g615 ( n1988 , n2096 , n2968 );
    and g616 ( n3557 , n3617 , n382 );
    nor g617 ( n552 , n3291 , n587 );
    and g618 ( n2829 , n1365 , n1704 );
    and g619 ( n2724 , n3009 , n3428 );
    or g620 ( n175 , n1295 , n1168 );
    or g621 ( n573 , n3202 , n189 );
    xnor g622 ( n3482 , n499 , n2174 );
    and g623 ( n485 , n1145 , n849 );
    not g624 ( n931 , n3171 );
    or g625 ( n1966 , n3404 , n138 );
    or g626 ( n2539 , n1803 , n3061 );
    not g627 ( n2024 , n1733 );
    and g628 ( n589 , n3667 , n2661 );
    or g629 ( n2694 , n3078 , n3443 );
    not g630 ( n2340 , n3018 );
    or g631 ( n1250 , n2163 , n702 );
    or g632 ( n1052 , n1307 , n2750 );
    and g633 ( n1110 , n1364 , n1191 );
    or g634 ( n2653 , n531 , n3678 );
    not g635 ( n2080 , n929 );
    xnor g636 ( n2495 , n2710 , n3508 );
    not g637 ( n13 , n1562 );
    or g638 ( n3647 , n2797 , n775 );
    or g639 ( n1876 , n1428 , n2289 );
    and g640 ( n1167 , n2568 , n944 );
    or g641 ( n2206 , n2271 , n2866 );
    or g642 ( n2286 , n188 , n1709 );
    xnor g643 ( n1261 , n1211 , n1466 );
    or g644 ( n616 , n2100 , n3374 );
    or g645 ( n853 , n352 , n800 );
    xnor g646 ( n894 , n2132 , n698 );
    or g647 ( n564 , n534 , n2032 );
    nor g648 ( n1107 , n3182 , n2478 );
    not g649 ( n1995 , n1799 );
    or g650 ( n322 , n915 , n3421 );
    xor g651 ( n3252 , n2271 , n1304 );
    not g652 ( n3345 , n941 );
    xnor g653 ( n1817 , n1687 , n507 );
    or g654 ( n1175 , n2220 , n2603 );
    and g655 ( n2444 , n677 , n2938 );
    xnor g656 ( n3367 , n3211 , n396 );
    or g657 ( n2598 , n466 , n3318 );
    xnor g658 ( n2404 , n2002 , n2110 );
    and g659 ( n2181 , n1862 , n3525 );
    or g660 ( n1739 , n2829 , n1600 );
    or g661 ( n1910 , n2819 , n3634 );
    not g662 ( n3272 , n3439 );
    or g663 ( n951 , n626 , n3228 );
    and g664 ( n3581 , n2044 , n119 );
    nor g665 ( n607 , n77 , n491 );
    nor g666 ( n2871 , n3106 , n2832 );
    or g667 ( n928 , n3546 , n3130 );
    or g668 ( n1899 , n952 , n928 );
    not g669 ( n1361 , n1120 );
    not g670 ( n2940 , n417 );
    xnor g671 ( n2199 , n1533 , n2168 );
    xnor g672 ( n1687 , n2824 , n2412 );
    nor g673 ( n2506 , n1428 , n2406 );
    and g674 ( n3273 , n627 , n403 );
    or g675 ( n3618 , n3257 , n936 );
    or g676 ( n2843 , n3053 , n270 );
    and g677 ( n297 , n3156 , n1948 );
    not g678 ( n2104 , n1949 );
    not g679 ( n3331 , n1428 );
    or g680 ( n481 , n2569 , n3634 );
    or g681 ( n2114 , n533 , n3597 );
    or g682 ( n3031 , n1690 , n1957 );
    or g683 ( n2403 , n2544 , n3001 );
    and g684 ( n2038 , n1340 , n2003 );
    and g685 ( n1476 , n770 , n3266 );
    xnor g686 ( n1185 , n1473 , n3372 );
    or g687 ( n1643 , n413 , n3190 );
    or g688 ( n2925 , n2994 , n1811 );
    and g689 ( n1215 , n555 , n1461 );
    xnor g690 ( n1618 , n3301 , n274 );
    nor g691 ( n3191 , n2178 , n3555 );
    and g692 ( n800 , n1793 , n3115 );
    xnor g693 ( n1044 , n1150 , n3135 );
    not g694 ( n137 , n337 );
    and g695 ( n2461 , n1456 , n3474 );
    not g696 ( n1407 , n2861 );
    xnor g697 ( n3338 , n3259 , n1557 );
    not g698 ( n2013 , n685 );
    or g699 ( n3425 , n3587 , n2455 );
    and g700 ( n201 , n356 , n833 );
    xnor g701 ( n1936 , n1854 , n3535 );
    xnor g702 ( n1069 , n2451 , n1478 );
    or g703 ( n870 , n1596 , n2712 );
    and g704 ( n1977 , n344 , n1177 );
    not g705 ( n318 , n2365 );
    nor g706 ( n1695 , n1743 , n1289 );
    xnor g707 ( n1940 , n1309 , n624 );
    or g708 ( n2494 , n410 , n620 );
    xnor g709 ( n2751 , n983 , n3591 );
    xnor g710 ( n2991 , n1265 , n1911 );
    xnor g711 ( n2863 , n168 , n3337 );
    or g712 ( n2584 , n359 , n2054 );
    and g713 ( n1487 , n879 , n1292 );
    or g714 ( n2219 , n3202 , n955 );
    xnor g715 ( n3559 , n2612 , n2883 );
    or g716 ( n1630 , n2515 , n3166 );
    and g717 ( n2937 , n1834 , n3350 );
    and g718 ( n1788 , n2597 , n1296 );
    xnor g719 ( n2669 , n557 , n2563 );
    or g720 ( n1944 , n128 , n1138 );
    and g721 ( n3020 , n2195 , n187 );
    or g722 ( n1079 , n2163 , n1663 );
    xnor g723 ( n361 , n1994 , n76 );
    or g724 ( n3492 , n2844 , n880 );
    and g725 ( n3626 , n2958 , n259 );
    or g726 ( n1530 , n1399 , n1277 );
    not g727 ( n3634 , n3329 );
    xnor g728 ( n1304 , n1052 , n521 );
    and g729 ( n1870 , n45 , n2315 );
    not g730 ( n2648 , n1271 );
    and g731 ( n1820 , n3380 , n689 );
    or g732 ( n1430 , n2946 , n1509 );
    nor g733 ( n940 , n1252 , n3026 );
    xnor g734 ( n158 , n2171 , n3464 );
    or g735 ( n1965 , n2220 , n3443 );
    and g736 ( n3347 , n862 , n317 );
    xnor g737 ( n491 , n1162 , n1655 );
    or g738 ( n2896 , n1391 , n2622 );
    not g739 ( n2362 , n1901 );
    or g740 ( n3354 , n1073 , n3267 );
    or g741 ( n234 , n851 , n2186 );
    xnor g742 ( n1559 , n1121 , n1632 );
    xnor g743 ( n1068 , n534 , n665 );
    nor g744 ( n2005 , n1925 , n1339 );
    or g745 ( n1080 , n1014 , n600 );
    or g746 ( n1816 , n1508 , n215 );
    xnor g747 ( n834 , n2414 , n2787 );
    or g748 ( n2356 , n2422 , n334 );
    or g749 ( n2061 , n128 , n329 );
    xnor g750 ( n1412 , n3306 , n2962 );
    or g751 ( n1810 , n3279 , n3236 );
    nor g752 ( n2367 , n3537 , n2694 );
    or g753 ( n2079 , n27 , n3290 );
    and g754 ( n3149 , n342 , n699 );
    or g755 ( n11 , n851 , n2489 );
    or g756 ( n2288 , n2187 , n2352 );
    or g757 ( n1980 , n204 , n24 );
    xnor g758 ( n673 , n2087 , n3561 );
    not g759 ( n2349 , n1375 );
    or g760 ( n2454 , n2674 , n2361 );
    or g761 ( n2721 , n2134 , n3285 );
    or g762 ( n1832 , n656 , n3562 );
    not g763 ( n2908 , n3616 );
    and g764 ( n2585 , n151 , n884 );
    xnor g765 ( n2412 , n2772 , n2060 );
    and g766 ( n2926 , n778 , n3482 );
    xnor g767 ( n3269 , n79 , n1784 );
    or g768 ( n1846 , n1568 , n229 );
    and g769 ( n789 , n1141 , n2909 );
    or g770 ( n56 , n918 , n1049 );
    or g771 ( n3330 , n3293 , n2233 );
    and g772 ( n1637 , n523 , n2316 );
    or g773 ( n754 , n2589 , n92 );
    not g774 ( n1558 , n2195 );
    or g775 ( n2704 , n701 , n1482 );
    or g776 ( n890 , n1886 , n225 );
    xnor g777 ( n1051 , n2969 , n3084 );
    nor g778 ( n3165 , n2468 , n460 );
    not g779 ( n2750 , n1613 );
    xnor g780 ( n65 , n565 , n3307 );
    xnor g781 ( n2411 , n3394 , n3452 );
    and g782 ( n919 , n166 , n1571 );
    or g783 ( n2787 , n27 , n1992 );
    not g784 ( n360 , n829 );
    xnor g785 ( n3361 , n1959 , n1072 );
    not g786 ( n1887 , n1308 );
    or g787 ( n3011 , n2818 , n3111 );
    not g788 ( n2177 , n3354 );
    xnor g789 ( n1317 , n1371 , n3 );
    or g790 ( n683 , n2535 , n1138 );
    xnor g791 ( n2865 , n1786 , n3170 );
    and g792 ( n511 , n1864 , n2618 );
    xnor g793 ( n2824 , n663 , n3527 );
    or g794 ( n2423 , n1944 , n103 );
    or g795 ( n2550 , n1428 , n2607 );
    or g796 ( n2121 , n58 , n3264 );
    xnor g797 ( n756 , n247 , n2674 );
    and g798 ( n1120 , n1382 , n435 );
    or g799 ( n3432 , n128 , n3546 );
    xnor g800 ( n3055 , n1223 , n2628 );
    or g801 ( n1703 , n129 , n2794 );
    and g802 ( n3225 , n2262 , n1776 );
    or g803 ( n2353 , n1941 , n2229 );
    and g804 ( n1892 , n462 , n21 );
    or g805 ( n433 , n2175 , n2685 );
    xnor g806 ( n1393 , n1270 , n800 );
    or g807 ( n605 , n758 , n1438 );
    or g808 ( n1305 , n1425 , n2028 );
    not g809 ( n1059 , n2738 );
    or g810 ( n2 , n2598 , n1501 );
    xnor g811 ( n420 , n144 , n42 );
    or g812 ( n1577 , n2163 , n2278 );
    and g813 ( n2468 , n417 , n136 );
    and g814 ( n2929 , n474 , n320 );
    and g815 ( n2619 , n2377 , n1080 );
    and g816 ( n3409 , n2306 , n210 );
    xnor g817 ( n532 , n3350 , n2169 );
    or g818 ( n1071 , n3671 , n1653 );
    and g819 ( n3572 , n2109 , n1714 );
    or g820 ( n381 , n1428 , n829 );
    and g821 ( n3461 , n726 , n2329 );
    nor g822 ( n1580 , n116 , n3628 );
    and g823 ( n3509 , n1462 , n2176 );
    or g824 ( n930 , n10 , n1116 );
    xnor g825 ( n2741 , n1561 , n2940 );
    nor g826 ( n416 , n651 , n2248 );
    or g827 ( n1849 , n2014 , n705 );
    and g828 ( n2036 , n1434 , n1672 );
    and g829 ( n3234 , n2914 , n821 );
    and g830 ( n404 , n439 , n287 );
    xnor g831 ( n176 , n45 , n632 );
    or g832 ( n3077 , n1764 , n135 );
    or g833 ( n2700 , n2612 , n2067 );
    or g834 ( n356 , n2291 , n2074 );
    and g835 ( n2511 , n3353 , n1745 );
    and g836 ( n1978 , n2215 , n2988 );
    xnor g837 ( n818 , n2308 , n2982 );
    or g838 ( n2133 , n31 , n299 );
    xnor g839 ( n1881 , n1650 , n706 );
    xnor g840 ( n3445 , n744 , n1737 );
    or g841 ( n2710 , n1814 , n3152 );
    and g842 ( n956 , n1214 , n2287 );
    nor g843 ( n2254 , n1200 , n168 );
    nor g844 ( n2339 , n2973 , n2816 );
    and g845 ( n2211 , n1345 , n3213 );
    or g846 ( n2480 , n2553 , n2750 );
    nor g847 ( n2967 , n1962 , n2779 );
    or g848 ( n1024 , n659 , n2127 );
    and g849 ( n3188 , n2091 , n529 );
    or g850 ( n1927 , n517 , n1330 );
    or g851 ( n3393 , n2150 , n634 );
    and g852 ( n922 , n3091 , n687 );
    or g853 ( n3250 , n1320 , n1994 );
    and g854 ( n571 , n3394 , n3452 );
    or g855 ( n2877 , n3259 , n2000 );
    or g856 ( n2797 , n2631 , n2398 );
    not g857 ( n793 , n3273 );
    not g858 ( n2632 , n1989 );
    xnor g859 ( n49 , n3320 , n1981 );
    or g860 ( n3014 , n1363 , n2528 );
    xnor g861 ( n2900 , n868 , n604 );
    and g862 ( n3215 , n2266 , n619 );
    xnor g863 ( n869 , n2730 , n2158 );
    xnor g864 ( n2006 , n1501 , n741 );
    or g865 ( n442 , n173 , n2671 );
    or g866 ( n3301 , n1509 , n1446 );
    xnor g867 ( n364 , n3506 , n2295 );
    xnor g868 ( n3307 , n1550 , n1615 );
    xnor g869 ( n1968 , n460 , n1318 );
    or g870 ( n1649 , n1661 , n2010 );
    or g871 ( n1700 , n3303 , n3545 );
    or g872 ( n156 , n1999 , n155 );
    or g873 ( n3600 , n1695 , n495 );
    or g874 ( n398 , n53 , n3318 );
    or g875 ( n1399 , n38 , n955 );
    or g876 ( n2396 , n2535 , n329 );
    and g877 ( n2798 , n1824 , n2037 );
    or g878 ( n3463 , n3048 , n893 );
    or g879 ( n3474 , n1077 , n1487 );
    and g880 ( n2930 , n3257 , n936 );
    and g881 ( n119 , n2838 , n747 );
    or g882 ( n2992 , n1319 , n2197 );
    and g883 ( n3449 , n1096 , n1550 );
    or g884 ( n604 , n2517 , n1992 );
    or g885 ( n3638 , n3326 , n802 );
    not g886 ( n3538 , n2709 );
    and g887 ( n2158 , n1914 , n948 );
    and g888 ( n2439 , n1633 , n3006 );
    or g889 ( n3108 , n60 , n2614 );
    and g890 ( n157 , n1211 , n2015 );
    xnor g891 ( n1303 , n2350 , n2743 );
    and g892 ( n976 , n2353 , n996 );
    xnor g893 ( n1848 , n3185 , n3392 );
    or g894 ( n295 , n2291 , n1243 );
    or g895 ( n761 , n1249 , n2899 );
    or g896 ( n1614 , n2163 , n2400 );
    nor g897 ( n235 , n3063 , n3128 );
    or g898 ( n850 , n1902 , n1475 );
    or g899 ( n15 , n654 , n2461 );
    not g900 ( n382 , n2651 );
    nor g901 ( n2033 , n2944 , n1896 );
    or g902 ( n33 , n1719 , n1017 );
    xnor g903 ( n2726 , n1161 , n893 );
    xnor g904 ( n3035 , n2324 , n1934 );
    xnor g905 ( n2599 , n82 , n834 );
    not g906 ( n200 , n1602 );
    and g907 ( n3455 , n3288 , n1831 );
    not g908 ( n783 , n1241 );
    or g909 ( n1565 , n1622 , n1521 );
    or g910 ( n2809 , n3248 , n3275 );
    and g911 ( n3173 , n3185 , n43 );
    or g912 ( n1831 , n1787 , n3082 );
    not g913 ( n603 , n403 );
    and g914 ( n2059 , n2107 , n2991 );
    not g915 ( n3555 , n932 );
    xnor g916 ( n1934 , n3011 , n857 );
    or g917 ( n2576 , n1883 , n1392 );
    or g918 ( n1786 , n3550 , n34 );
    xnor g919 ( n1745 , n3442 , n2410 );
    or g920 ( n726 , n1073 , n453 );
    not g921 ( n1868 , n145 );
    nor g922 ( n905 , n132 , n2428 );
    and g923 ( n3673 , n1376 , n661 );
    or g924 ( n572 , n3282 , n1642 );
    and g925 ( n1348 , n3075 , n3364 );
    not g926 ( n1354 , n702 );
    not g927 ( n2712 , n997 );
    and g928 ( n3064 , n1302 , n1458 );
    xnor g929 ( n2382 , n1944 , n2255 );
    not g930 ( n802 , n1282 );
    and g931 ( n2081 , n1549 , n1341 );
    or g932 ( n1173 , n722 , n1608 );
    xnor g933 ( n1615 , n1096 , n1804 );
    and g934 ( n3404 , n2320 , n2860 );
    or g935 ( n3024 , n2990 , n2599 );
    not g936 ( n288 , n3565 );
    xnor g937 ( n2904 , n2072 , n249 );
    or g938 ( n3288 , n3438 , n3330 );
    and g939 ( n39 , n1803 , n3061 );
    and g940 ( n2502 , n3271 , n1891 );
    xnor g941 ( n912 , n3283 , n987 );
    or g942 ( n3198 , n1591 , n247 );
    not g943 ( n1511 , n2240 );
    not g944 ( n1164 , n361 );
    and g945 ( n139 , n2895 , n1854 );
    xnor g946 ( n1532 , n2493 , n1423 );
    or g947 ( n3116 , n2517 , n1015 );
    or g948 ( n2513 , n1440 , n2425 );
    or g949 ( n1177 , n2527 , n2969 );
    or g950 ( n1919 , n646 , n1850 );
    or g951 ( n93 , n2660 , n1712 );
    and g952 ( n1906 , n1173 , n1325 );
    and g953 ( n620 , n2239 , n93 );
    or g954 ( n735 , n3615 , n1868 );
    xnor g955 ( n2275 , n898 , n1328 );
    not g956 ( n487 , n1960 );
    nor g957 ( n549 , n785 , n3515 );
    xnor g958 ( n1491 , n1582 , n982 );
    xnor g959 ( n2563 , n1899 , n617 );
    or g960 ( n1896 , n338 , n3447 );
    not g961 ( n1534 , n3065 );
    or g962 ( n2451 , n2569 , n645 );
    xnor g963 ( n691 , n870 , n1482 );
    or g964 ( n864 , n1584 , n608 );
    or g965 ( n2082 , n2409 , n2406 );
    xnor g966 ( n1942 , n3412 , n2954 );
    xnor g967 ( n2212 , n695 , n244 );
    xnor g968 ( n85 , n340 , n2854 );
    and g969 ( n1518 , n1771 , n2774 );
    not g970 ( n2074 , n272 );
    xnor g971 ( n1346 , n1850 , n2842 );
    and g972 ( n3065 , n2016 , n1982 );
    or g973 ( n1517 , n173 , n34 );
    or g974 ( n1549 , n835 , n3251 );
    not g975 ( n3649 , n1339 );
    or g976 ( n1579 , n2291 , n1868 );
    and g977 ( n2469 , n983 , n986 );
    and g978 ( n1269 , n1480 , n425 );
    or g979 ( n1191 , n2517 , n445 );
    xnor g980 ( n1747 , n2796 , n3620 );
    nor g981 ( n3204 , n2399 , n3196 );
    xnor g982 ( n2273 , n2006 , n2633 );
    xnor g983 ( n838 , n2280 , n378 );
    xnor g984 ( n2246 , n1830 , n509 );
    or g985 ( n696 , n466 , n1801 );
    or g986 ( n3630 , n2331 , n2749 );
    not g987 ( n331 , n1790 );
    and g988 ( n2153 , n2811 , n3636 );
    not g989 ( n1603 , n1167 );
    or g990 ( n675 , n2901 , n1265 );
    xnor g991 ( n3592 , n647 , n3431 );
    or g992 ( n3558 , n3598 , n1182 );
    and g993 ( n545 , n3177 , n256 );
    and g994 ( n231 , n2656 , n3639 );
    or g995 ( n867 , n1987 , n2651 );
    and g996 ( n1136 , n206 , n2471 );
    and g997 ( n2051 , n2321 , n2049 );
    and g998 ( n2197 , n2133 , n752 );
    and g999 ( n1834 , n1065 , n447 );
    and g1000 ( n3663 , n148 , n1694 );
    not g1001 ( n2294 , n161 );
    xnor g1002 ( n2091 , n11 , n2540 );
    and g1003 ( n2762 , n2889 , n858 );
    or g1004 ( n1193 , n2741 , n567 );
    or g1005 ( n1311 , n2084 , n357 );
    xnor g1006 ( n2681 , n1440 , n2425 );
    or g1007 ( n3357 , n173 , n2712 );
    not g1008 ( n3349 , n2034 );
    nor g1009 ( n233 , n3459 , n2566 );
    or g1010 ( n2846 , n2753 , n2039 );
    xnor g1011 ( n1999 , n913 , n1477 );
    xnor g1012 ( n2673 , n2618 , n1331 );
    xnor g1013 ( n1884 , n503 , n3675 );
    not g1014 ( n3352 , n2136 );
    or g1015 ( n2383 , n2233 , n3432 );
    and g1016 ( n1972 , n3430 , n648 );
    not g1017 ( n2415 , n1732 );
    or g1018 ( n484 , n836 , n2608 );
    xnor g1019 ( n1232 , n451 , n75 );
    and g1020 ( n2042 , n579 , n59 );
    xnor g1021 ( n3570 , n1518 , n1323 );
    or g1022 ( n370 , n2220 , n2709 );
    xnor g1023 ( n2470 , n9 , n2323 );
    xnor g1024 ( n598 , n2221 , n713 );
    and g1025 ( n2883 , n281 , n1034 );
    not g1026 ( n466 , n579 );
    or g1027 ( n1606 , n663 , n3199 );
    and g1028 ( n669 , n1512 , n730 );
    or g1029 ( n286 , n1018 , n3315 );
    xnor g1030 ( n1912 , n1525 , n3225 );
    xnor g1031 ( n611 , n670 , n3319 );
    or g1032 ( n1181 , n209 , n607 );
    xnor g1033 ( n127 , n1135 , n1822 );
    or g1034 ( n1141 , n3091 , n687 );
    or g1035 ( n236 , n16 , n2650 );
    or g1036 ( n797 , n1641 , n340 );
    xnor g1037 ( n1172 , n690 , n667 );
    not g1038 ( n978 , n734 );
    and g1039 ( n2463 , n2901 , n1265 );
    or g1040 ( n2422 , n3615 , n2664 );
    xnor g1041 ( n1799 , n567 , n125 );
    or g1042 ( n2791 , n204 , n2968 );
    xnor g1043 ( n79 , n3321 , n3434 );
    or g1044 ( n3452 , n2946 , n1648 );
    or g1045 ( n3323 , n3153 , n2022 );
    or g1046 ( n3059 , n1518 , n818 );
    xor g1047 ( n1301 , n943 , n935 );
    and g1048 ( n3270 , n3319 , n670 );
    not g1049 ( n866 , n2178 );
    xnor g1050 ( n633 , n1194 , n2131 );
    or g1051 ( n593 , n639 , n525 );
    and g1052 ( n1447 , n465 , n2462 );
    or g1053 ( n2491 , n905 , n3469 );
    xnor g1054 ( n831 , n1290 , n3656 );
    or g1055 ( n3164 , n351 , n1278 );
    or g1056 ( n367 , n1451 , n1681 );
    or g1057 ( n1882 , n1054 , n3634 );
    xnor g1058 ( n2015 , n215 , n1272 );
    nor g1059 ( n2333 , n3546 , n422 );
    or g1060 ( n2737 , n1503 , n2756 );
    nor g1061 ( n2631 , n1091 , n837 );
    nor g1062 ( n1611 , n2017 , n3577 );
    or g1063 ( n2559 , n1552 , n802 );
    xnor g1064 ( n1318 , n2468 , n196 );
    or g1065 ( n2910 , n2298 , n2659 );
    nor g1066 ( n550 , n643 , n2978 );
    not g1067 ( n1857 , n2039 );
    and g1068 ( n3048 , n1161 , n1727 );
    or g1069 ( n865 , n204 , n2294 );
    xnor g1070 ( n2948 , n2580 , n468 );
    and g1071 ( n3123 , n3101 , n3327 );
    and g1072 ( n2447 , n1134 , n74 );
    or g1073 ( n2773 , n1540 , n3290 );
    xnor g1074 ( n1673 , n765 , n2035 );
    xor g1075 ( n507 , n3441 , n1043 );
    or g1076 ( n1095 , n2710 , n3508 );
    or g1077 ( n2627 , n3546 , n1724 );
    and g1078 ( n212 , n517 , n1330 );
    or g1079 ( n2346 , n851 , n329 );
    or g1080 ( n1065 , n2626 , n1517 );
    or g1081 ( n3200 , n940 , n784 );
    not g1082 ( n2200 , n2372 );
    and g1083 ( n2370 , n2391 , n1354 );
    or g1084 ( n1264 , n2696 , n1235 );
    and g1085 ( n471 , n3486 , n973 );
    and g1086 ( n924 , n1543 , n2450 );
    xnor g1087 ( n1545 , n442 , n1678 );
    and g1088 ( n3321 , n2179 , n3066 );
    and g1089 ( n2763 , n56 , n574 );
    or g1090 ( n25 , n3375 , n2141 );
    xnor g1091 ( n3535 , n2895 , n1592 );
    and g1092 ( n1918 , n3543 , n3205 );
    and g1093 ( n1964 , n2874 , n2434 );
    or g1094 ( n2008 , n956 , n1965 );
    or g1095 ( n2327 , n680 , n3254 );
    nor g1096 ( n2542 , n1027 , n3622 );
    xnor g1097 ( n2338 , n1977 , n1903 );
    or g1098 ( n1420 , n91 , n3149 );
    or g1099 ( n3394 , n3272 , n1868 );
    nor g1100 ( n3159 , n3045 , n411 );
    and g1101 ( n2471 , n963 , n825 );
    or g1102 ( n12 , n2030 , n2489 );
    or g1103 ( n1404 , n1428 , n1879 );
    or g1104 ( n2524 , n1428 , n3478 );
    or g1105 ( n2092 , n441 , n2074 );
    xnor g1106 ( n319 , n3416 , n3147 );
    not g1107 ( n953 , n48 );
    or g1108 ( n3552 , n3550 , n1921 );
    xnor g1109 ( n1251 , n2795 , n920 );
    xnor g1110 ( n340 , n2973 , n2972 );
    and g1111 ( n2888 , n3237 , n54 );
    xnor g1112 ( n3580 , n2520 , n307 );
    or g1113 ( n1242 , n1688 , n2212 );
    and g1114 ( n1880 , n1380 , n3099 );
    not g1115 ( n2990 , n2607 );
    and g1116 ( n3528 , n1643 , n761 );
    or g1117 ( n1797 , n827 , n328 );
    or g1118 ( n3574 , n3202 , n1235 );
    or g1119 ( n1113 , n3550 , n18 );
    or g1120 ( n1776 , n541 , n479 );
    and g1121 ( n2257 , n1274 , n1457 );
    and g1122 ( n1557 , n3613 , n3118 );
    or g1123 ( n2838 , n1639 , n625 );
    xor g1124 ( n3074 , n2461 , n654 );
    xnor g1125 ( n83 , n1683 , n316 );
    and g1126 ( n2727 , n696 , n1979 );
    or g1127 ( n1369 , n2220 , n1558 );
    xnor g1128 ( n1915 , n858 , n3659 );
    or g1129 ( n1074 , n3138 , n2063 );
    and g1130 ( n1220 , n3298 , n102 );
    not g1131 ( n1689 , n3151 );
    not g1132 ( n3396 , n1627 );
    and g1133 ( n1555 , n1150 , n3135 );
    not g1134 ( n220 , n2906 );
    and g1135 ( n2879 , n540 , n1489 );
    xor g1136 ( n1213 , n789 , n1251 );
    and g1137 ( n3239 , n3277 , n576 );
    or g1138 ( n2690 , n1609 , n1447 );
    or g1139 ( n2936 , n855 , n1885 );
    or g1140 ( n3489 , n2070 , n2932 );
    or g1141 ( n1925 , n764 , n878 );
    xnor g1142 ( n144 , n722 , n2097 );
    not g1143 ( n581 , n1900 );
    nor g1144 ( n3460 , n896 , n178 );
    or g1145 ( n2196 , n2060 , n927 );
    and g1146 ( n260 , n1210 , n3200 );
    or g1147 ( n3567 , n2615 , n2186 );
    xnor g1148 ( n3383 , n2135 , n3085 );
    or g1149 ( n2779 , n2090 , n339 );
    or g1150 ( n3068 , n3248 , n2664 );
    or g1151 ( n292 , n684 , n762 );
    or g1152 ( n483 , n1069 , n2279 );
    not g1153 ( n944 , n1476 );
    not g1154 ( n77 , n2075 );
    xnor g1155 ( n2621 , n3200 , n265 );
    xnor g1156 ( n743 , n2136 , n3355 );
    xnor g1157 ( n1330 , n3030 , n368 );
    or g1158 ( n2965 , n107 , n2557 );
    or g1159 ( n469 , n184 , n2164 );
    and g1160 ( n1744 , n3576 , n1335 );
    or g1161 ( n3194 , n280 , n2209 );
    or g1162 ( n3606 , n182 , n824 );
    or g1163 ( n1623 , n1702 , n2087 );
    and g1164 ( n2295 , n1657 , n2588 );
    xnor g1165 ( n3107 , n2219 , n2634 );
    and g1166 ( n2498 , n2560 , n405 );
    or g1167 ( n3266 , n19 , n1879 );
    or g1168 ( n855 , n897 , n3290 );
    and g1169 ( n1441 , n1451 , n1681 );
    and g1170 ( n2573 , n1513 , n1137 );
    and g1171 ( n2821 , n1720 , n2658 );
    not g1172 ( n2691 , n1548 );
    and g1173 ( n1889 , n566 , n430 );
    xor g1174 ( n1718 , n2537 , n596 );
    xnor g1175 ( n306 , n2970 , n852 );
    or g1176 ( n1277 , n581 , n1921 );
    or g1177 ( n3308 , n895 , n3092 );
    or g1178 ( n3320 , n1307 , n3267 );
    and g1179 ( n1922 , n658 , n2810 );
    or g1180 ( n2018 , n1026 , n2155 );
    not g1181 ( n3485 , n1843 );
    xnor g1182 ( n16 , n1936 , n1465 );
    and g1183 ( n2790 , n941 , n810 );
    or g1184 ( n828 , n3272 , n1243 );
    xnor g1185 ( n2972 , n2816 , n662 );
    and g1186 ( n1544 , n1941 , n2229 );
    not g1187 ( n1230 , n2759 );
    xnor g1188 ( n1762 , n3336 , n65 );
    xnor g1189 ( n3291 , n2274 , n1450 );
    or g1190 ( n1442 , n3546 , n3166 );
    xnor g1191 ( n943 , n3676 , n2318 );
    and g1192 ( n1533 , n2957 , n2862 );
    or g1193 ( n227 , n1631 , n24 );
    xnor g1194 ( n2430 , n1277 , n2915 );
    or g1195 ( n3640 , n1912 , n459 );
    xnor g1196 ( n1398 , n2718 , n3278 );
    nor g1197 ( n134 , n505 , n662 );
    xnor g1198 ( n1875 , n1410 , n2487 );
    or g1199 ( n2167 , n2995 , n1066 );
    nor g1200 ( n1419 , n97 , n1529 );
    or g1201 ( n3284 , n3549 , n422 );
    or g1202 ( n619 , n224 , n3159 );
    xnor g1203 ( n2640 , n1637 , n2783 );
    or g1204 ( n1025 , n179 , n214 );
    xnor g1205 ( n2586 , n147 , n397 );
    or g1206 ( n3019 , n3212 , n2203 );
    or g1207 ( n142 , n3473 , n3363 );
    xor g1208 ( n2235 , n1791 , n2386 );
    or g1209 ( n2336 , n3086 , n1621 );
    xnor g1210 ( n2828 , n3661 , n2574 );
    xnor g1211 ( n3182 , n1743 , n3608 );
    or g1212 ( n3171 , n1307 , n453 );
    and g1213 ( n3406 , n2477 , n2442 );
    not g1214 ( n3355 , n2208 );
    and g1215 ( n1902 , n1180 , n3359 );
    xor g1216 ( n1359 , n202 , n3390 );
    xnor g1217 ( n586 , n2213 , n1685 );
    or g1218 ( n1951 , n1923 , n546 );
    or g1219 ( n1208 , n1649 , n2817 );
    or g1220 ( n3093 , n2946 , n2664 );
    or g1221 ( n242 , n2804 , n2766 );
    xnor g1222 ( n2066 , n1624 , n3150 );
    xnor g1223 ( n1539 , n1346 , n1207 );
    xnor g1224 ( n0 , n71 , n1068 );
    xnor g1225 ( n1072 , n295 , n861 );
    and g1226 ( n1130 , n1271 , n2188 );
    or g1227 ( n406 , n3062 , n2520 );
    xnor g1228 ( n2252 , n3397 , n2411 );
    or g1229 ( n2868 , n3185 , n43 );
    or g1230 ( n3052 , n1405 , n3634 );
    and g1231 ( n1194 , n105 , n990 );
    and g1232 ( n901 , n1654 , n2194 );
    not g1233 ( n208 , n3224 );
    or g1234 ( n389 , n2350 , n719 );
    xnor g1235 ( n1452 , n2880 , n2902 );
    or g1236 ( n1982 , n1379 , n782 );
    and g1237 ( n2078 , n3279 , n3236 );
    xnor g1238 ( n3233 , n2749 , n2159 );
    xnor g1239 ( n2485 , n1388 , n501 );
    or g1240 ( n996 , n1050 , n1544 );
    or g1241 ( n2597 , n3326 , n2968 );
    xnor g1242 ( n2274 , n43 , n1848 );
    or g1243 ( n40 , n1887 , n3318 );
    xnor g1244 ( n100 , n1349 , n3040 );
    and g1245 ( n2668 , n856 , n1545 );
    or g1246 ( n2822 , n3615 , n1334 );
    or g1247 ( n2392 , n683 , n2490 );
    xnor g1248 ( n3362 , n1958 , n575 );
    not g1249 ( n1156 , n3109 );
    or g1250 ( n2364 , n2946 , n1868 );
    nor g1251 ( n1701 , n2882 , n2734 );
    and g1252 ( n2369 , n2759 , n2115 );
    and g1253 ( n2276 , n514 , n308 );
    and g1254 ( n1550 , n3647 , n2960 );
    or g1255 ( n3433 , n897 , n1015 );
    or g1256 ( n1426 , n3417 , n649 );
    xnor g1257 ( n3219 , n526 , n2383 );
    not g1258 ( n1372 , n1382 );
    and g1259 ( n3511 , n2328 , n1005 );
    and g1260 ( n639 , n1344 , n2974 );
    nor g1261 ( n294 , n438 , n518 );
    xnor g1262 ( n2859 , n1622 , n1902 );
    not g1263 ( n2247 , n3514 );
    or g1264 ( n3419 , n1349 , n2482 );
    nor g1265 ( n1102 , n1860 , n2436 );
    xnor g1266 ( n1352 , n795 , n364 );
    or g1267 ( n916 , n759 , n1877 );
    xnor g1268 ( n1938 , n135 , n1668 );
    xnor g1269 ( n3292 , n206 , n2471 );
    and g1270 ( n2625 , n2061 , n1045 );
    or g1271 ( n1218 , n94 , n2519 );
    xnor g1272 ( n1323 , n1337 , n2507 );
    or g1273 ( n3138 , n2362 , n1648 );
    xnor g1274 ( n1655 , n1790 , n1361 );
    and g1275 ( n827 , n578 , n2120 );
    xnor g1276 ( n2735 , n160 , n1699 );
    or g1277 ( n2649 , n2517 , n2830 );
    and g1278 ( n2448 , n846 , n2602 );
    or g1279 ( n2878 , n1958 , n515 );
    or g1280 ( n1709 , n2946 , n1243 );
    and g1281 ( n75 , n3262 , n1099 );
    and g1282 ( n3309 , n1821 , n816 );
    and g1283 ( n1548 , n200 , n1995 );
    and g1284 ( n2214 , n1832 , n1857 );
    not g1285 ( n222 , n3161 );
    xnor g1286 ( n1749 , n3094 , n280 );
    or g1287 ( n117 , n575 , n977 );
    or g1288 ( n1 , n1887 , n3634 );
    or g1289 ( n1265 , n2819 , n1573 );
    or g1290 ( n3665 , n457 , n1801 );
    xnor g1291 ( n986 , n3433 , n2900 );
    and g1292 ( n1515 , n2598 , n1501 );
    and g1293 ( n1182 , n2079 , n2825 );
    not g1294 ( n3583 , n1313 );
    and g1295 ( n2616 , n3680 , n366 );
    or g1296 ( n3512 , n3052 , n1040 );
    or g1297 ( n1856 , n1054 , n1573 );
    and g1298 ( n2603 , n2216 , n165 );
    and g1299 ( n2043 , n1753 , n1974 );
    and g1300 ( n3258 , n1620 , n261 );
    or g1301 ( n2332 , n1631 , n2294 );
    and g1302 ( n859 , n2700 , n1498 );
    or g1303 ( n463 , n1473 , n2346 );
    or g1304 ( n1916 , n713 , n560 );
    or g1305 ( n3551 , n2595 , n3649 );
    and g1306 ( n1482 , n2427 , n548 );
    and g1307 ( n583 , n950 , n2207 );
    and g1308 ( n968 , n2855 , n28 );
    xnor g1309 ( n742 , n3138 , n2063 );
    not g1310 ( n1921 , n1055 );
    xnor g1311 ( n2672 , n3177 , n3528 );
    and g1312 ( n2596 , n2378 , n2688 );
    or g1313 ( n2260 , n868 , n604 );
    or g1314 ( n2380 , n1307 , n2294 );
    or g1315 ( n1758 , n139 , n1592 );
    and g1316 ( n3586 , n350 , n2302 );
    or g1317 ( n180 , n3039 , n650 );
    nor g1318 ( n3549 , n2181 , n3139 );
    and g1319 ( n2475 , n953 , n2201 );
    and g1320 ( n184 , n3621 , n1427 );
    not g1321 ( n27 , n1411 );
    or g1322 ( n1467 , n3230 , n3409 );
    xnor g1323 ( n199 , n2477 , n3240 );
    or g1324 ( n3285 , n2220 , n3440 );
    and g1325 ( n2473 , n3630 , n1797 );
    not g1326 ( n3290 , n1692 );
    or g1327 ( n1510 , n2545 , n609 );
    xnor g1328 ( n2964 , n1172 , n489 );
    or g1329 ( n816 , n3673 , n144 );
    or g1330 ( n1782 , n3638 , n1028 );
    not g1331 ( n329 , n674 );
    xnor g1332 ( n2772 , n3193 , n1612 );
    and g1333 ( n3223 , n1095 , n1075 );
    xnor g1334 ( n273 , n994 , n1575 );
    and g1335 ( n2418 , n2617 , n2312 );
    nor g1336 ( n1578 , n569 , n685 );
    or g1337 ( n2646 , n160 , n2160 );
    or g1338 ( n1945 , n1575 , n470 );
    not g1339 ( n2696 , n3662 );
    or g1340 ( n3658 , n1572 , n1174 );
    and g1341 ( n2352 , n386 , n283 );
    or g1342 ( n2243 , n1661 , n1573 );
    nor g1343 ( n544 , n2281 , n264 );
    xnor g1344 ( n1329 , n2465 , n1227 );
    xnor g1345 ( n667 , n942 , n3086 );
    not g1346 ( n851 , n1119 );
    xnor g1347 ( n2861 , n178 , n896 );
    or g1348 ( n284 , n3 , n1371 );
    or g1349 ( n3125 , n401 , n3297 );
    and g1350 ( n3471 , n1576 , n1975 );
    nor g1351 ( n2323 , n1987 , n3249 );
    or g1352 ( n35 , n1552 , n3267 );
    or g1353 ( n26 , n2619 , n1863 );
    xnor g1354 ( n335 , n2329 , n2942 );
    xnor g1355 ( n1421 , n2160 , n2735 );
    and g1356 ( n3251 , n1305 , n3014 );
    and g1357 ( n1154 , n3537 , n2694 );
    and g1358 ( n240 , n275 , n142 );
    or g1359 ( n68 , n1987 , n1705 );
    or g1360 ( n913 , n3326 , n3267 );
    and g1361 ( n3360 , n2518 , n3541 );
    or g1362 ( n1370 , n876 , n1175 );
    or g1363 ( n541 , n53 , n3634 );
    and g1364 ( n2039 , n3345 , n718 );
    xnor g1365 ( n2954 , n1691 , n2066 );
    not g1366 ( n2671 , n2450 );
    or g1367 ( n3515 , n2928 , n1705 );
    xnor g1368 ( n183 , n3514 , n807 );
    not g1369 ( n3448 , n2851 );
    and g1370 ( n1592 , n3658 , n2299 );
    and g1371 ( n652 , n1784 , n79 );
    xnor g1372 ( n2978 , n1673 , n3402 );
    xnor g1373 ( n125 , n2741 , n823 );
    or g1374 ( n3025 , n581 , n189 );
    or g1375 ( n1061 , n641 , n2627 );
    or g1376 ( n1672 , n1043 , n591 );
    xnor g1377 ( n656 , n2688 , n2654 );
    or g1378 ( n2452 , n294 , n570 );
    or g1379 ( n1855 , n1870 , n632 );
    or g1380 ( n880 , n1987 , n2444 );
    not g1381 ( n1259 , n2145 );
    or g1382 ( n3479 , n1887 , n1801 );
    xnor g1383 ( n1179 , n3122 , n1195 );
    not g1384 ( n3196 , n803 );
    not g1385 ( n1667 , n902 );
    not g1386 ( n655 , n2769 );
    or g1387 ( n1458 , n2325 , n1580 );
    or g1388 ( n630 , n53 , n645 );
    or g1389 ( n578 , n335 , n3206 );
    nor g1390 ( n418 , n2493 , n3157 );
    or g1391 ( n2601 , n1741 , n2130 );
    xnor g1392 ( n2031 , n541 , n768 );
    or g1393 ( n2933 , n2163 , n2724 );
    or g1394 ( n2341 , n2317 , n3663 );
    xnor g1395 ( n3588 , n3638 , n3235 );
    or g1396 ( n243 , n1871 , n1138 );
    and g1397 ( n1765 , n1972 , n2042 );
    and g1398 ( n496 , n289 , n2601 );
    or g1399 ( n450 , n814 , n3067 );
    xnor g1400 ( n748 , n2792 , n69 );
    and g1401 ( n1433 , n3018 , n2845 );
    and g1402 ( n1877 , n3606 , n2026 );
    and g1403 ( n2102 , n828 , n2530 );
    xnor g1404 ( n3232 , n1344 , n3322 );
    xnor g1405 ( n628 , n428 , n1288 );
    or g1406 ( n2378 , n2819 , n1801 );
    not g1407 ( n3017 , n394 );
    or g1408 ( n1034 , n2578 , n602 );
    or g1409 ( n2358 , n3181 , n2182 );
    xnor g1410 ( n3236 , n2317 , n3378 );
    xnor g1411 ( n3470 , n3650 , n2503 );
    and g1412 ( n1640 , n3138 , n2063 );
    xnor g1413 ( n384 , n1607 , n3046 );
    xnor g1414 ( n2783 , n2602 , n512 );
    and g1415 ( n2565 , n1666 , n248 );
    xnor g1416 ( n2886 , n2814 , n3044 );
    or g1417 ( n2363 , n729 , n2689 );
    and g1418 ( n89 , n3467 , n3218 );
    and g1419 ( n3534 , n1616 , n277 );
    xnor g1420 ( n1143 , n1548 , n1968 );
    and g1421 ( n863 , n2390 , n3176 );
    or g1422 ( n3531 , n227 , n1991 );
    not g1423 ( n204 , n2303 );
    and g1424 ( n347 , n1966 , n2071 );
    or g1425 ( n23 , n2517 , n1707 );
    nor g1426 ( n1984 , n181 , n1064 );
    xnor g1427 ( n567 , n2758 , n1031 );
    and g1428 ( n2435 , n1231 , n3015 );
    or g1429 ( n3372 , n487 , n1138 );
    or g1430 ( n1933 , n2533 , n2625 );
    and g1431 ( n3553 , n1285 , n2154 );
    and g1432 ( n3012 , n1152 , n2704 );
    or g1433 ( n1563 , n766 , n1220 );
    or g1434 ( n3222 , n2432 , n2927 );
    or g1435 ( n2529 , n35 , n1196 );
    and g1436 ( n3577 , n1042 , n2146 );
    or g1437 ( n708 , n2806 , n1582 );
    xnor g1438 ( n1290 , n404 , n1721 );
    or g1439 ( n1142 , n2553 , n2294 );
    or g1440 ( n3091 , n1540 , n1707 );
    xnor g1441 ( n2641 , n3401 , n729 );
    or g1442 ( n2923 , n2295 , n2583 );
    xnor g1443 ( n3030 , n615 , n2681 );
    nor g1444 ( n3458 , n658 , n2810 );
    and g1445 ( n3189 , n3110 , n3304 );
    or g1446 ( n2044 , n3096 , n189 );
    or g1447 ( n2099 , n3192 , n1640 );
    and g1448 ( n190 , n2555 , n1337 );
    and g1449 ( n67 , n1856 , n1 );
    nor g1450 ( n478 , n3457 , n312 );
    or g1451 ( n1103 , n2371 , n3604 );
    and g1452 ( n3683 , n2151 , n426 );
    or g1453 ( n2958 , n773 , n216 );
    not g1454 ( n1073 , n2408 );
    or g1455 ( n113 , n3357 , n55 );
    xnor g1456 ( n229 , n2226 , n2198 );
    xnor g1457 ( n2532 , n3674 , n3493 );
    and g1458 ( n2259 , n123 , n2506 );
    or g1459 ( n2810 , n235 , n2870 );
    and g1460 ( n2270 , n452 , n2730 );
    not g1461 ( n3510 , n2675 );
    xnor g1462 ( n3608 , n1352 , n2217 );
    or g1463 ( n281 , n2364 , n3339 );
    or g1464 ( n796 , n1226 , n2048 );
    nor g1465 ( n714 , n3163 , n657 );
    xnor g1466 ( n2171 , n1451 , n2483 );
    and g1467 ( n2678 , n3567 , n2784 );
    and g1468 ( n357 , n2123 , n73 );
    or g1469 ( n3175 , n1899 , n557 );
    and g1470 ( n1139 , n427 , n2341 );
    and g1471 ( n2145 , n2247 , n2707 );
    or g1472 ( n2587 , n1284 , n325 );
    and g1473 ( n3646 , n2549 , n1147 );
    and g1474 ( n524 , n2663 , n1206 );
    or g1475 ( n804 , n2282 , n805 );
    or g1476 ( n1150 , n2030 , n554 );
    xnor g1477 ( n3169 , n3395 , n895 );
    and g1478 ( n1601 , n2804 , n2766 );
    and g1479 ( n750 , n1584 , n608 );
    nor g1480 ( n2290 , n565 , n3336 );
    and g1481 ( n3079 , n915 , n3421 );
    xnor g1482 ( n3536 , n2840 , n2760 );
    xnor g1483 ( n920 , n2558 , n976 );
    and g1484 ( n3023 , n651 , n2248 );
    not g1485 ( n2556 , n3628 );
    or g1486 ( n309 , n2477 , n2442 );
    or g1487 ( n2140 , n2952 , n3100 );
    and g1488 ( n178 , n3425 , n50 );
    and g1489 ( n1733 , n1471 , n2238 );
    not g1490 ( n2946 , n3073 );
    xnor g1491 ( n1328 , n1616 , n277 );
    or g1492 ( n2068 , n2359 , n1644 );
    xnor g1493 ( n3128 , n2974 , n3232 );
    not g1494 ( n2830 , n1183 );
    xnor g1495 ( n1913 , n1761 , n3021 );
    xnor g1496 ( n270 , n2430 , n628 );
    or g1497 ( n3505 , n2744 , n635 );
    and g1498 ( n1222 , n2529 , n120 );
    or g1499 ( n1554 , n1372 , n34 );
    and g1500 ( n813 , n2166 , n3162 );
    xnor g1501 ( n3114 , n2499 , n3184 );
    or g1502 ( n304 , n2719 , n2572 );
    and g1503 ( n2578 , n2364 , n3339 );
    or g1504 ( n3351 , n1479 , n2512 );
    or g1505 ( n965 , n3661 , n2574 );
    and g1506 ( n891 , n669 , n2827 );
    not g1507 ( n677 , n3684 );
    or g1508 ( n1766 , n471 , n900 );
    or g1509 ( n1853 , n3220 , n743 );
    nor g1510 ( n1665 , n3172 , n3129 );
    and g1511 ( n3056 , n2646 , n3571 );
    and g1512 ( n2973 , n1189 , n1025 );
    xnor g1513 ( n3094 , n1264 , n573 );
    xnor g1514 ( n3044 , n527 , n3333 );
    or g1515 ( n2267 , n1310 , n1138 );
    or g1516 ( n2156 , n502 , n2053 );
    not g1517 ( n1798 , n358 );
    and g1518 ( n701 , n870 , n1198 );
    or g1519 ( n415 , n2553 , n453 );
    and g1520 ( n2899 , n413 , n3190 );
    and g1521 ( n1602 , n1594 , n1153 );
    xnor g1522 ( n2825 , n1384 , n98 );
    xnor g1523 ( n58 , n3062 , n3580 );
    not g1524 ( n970 , n1003 );
    and g1525 ( n2592 , n1878 , n647 );
    nor g1526 ( n2893 , n1118 , n2486 );
    and g1527 ( n692 , n874 , n3429 );
    xnor g1528 ( n2386 , n2527 , n1051 );
    and g1529 ( n3363 , n1659 , n1444 );
    xnor g1530 ( n1729 , n2565 , n3646 );
    xnor g1531 ( n3160 , n1593 , n3602 );
    not g1532 ( n2952 , n1002 );
    and g1533 ( n3440 , n3017 , n2080 );
    xnor g1534 ( n3184 , n1137 , n1535 );
    or g1535 ( n278 , n2437 , n3408 );
    xnor g1536 ( n3597 , n786 , n2786 );
    and g1537 ( n2622 , n2437 , n3408 );
    and g1538 ( n2314 , n1533 , n1452 );
    xnor g1539 ( n1698 , n3230 , n1897 );
    or g1540 ( n2983 , n3032 , n1671 );
    not g1541 ( n2875 , n1346 );
    and g1542 ( n2840 , n2732 , n2891 );
    and g1543 ( n1845 , n1518 , n818 );
    xnor g1544 ( n3625 , n546 , n2069 );
    or g1545 ( n2466 , n183 , n1410 );
    and g1546 ( n1587 , n2492 , n1038 );
    or g1547 ( n680 , n2517 , n3152 );
    xnor g1548 ( n1796 , n2613 , n1222 );
    xnor g1549 ( n1961 , n1391 , n1560 );
    xor g1550 ( n3133 , n2394 , n467 );
    or g1551 ( n1198 , n581 , n1235 );
    or g1552 ( n3069 , n3392 , n3173 );
    and g1553 ( n1459 , n1269 , n2263 );
    and g1554 ( n1171 , n362 , n513 );
    or g1555 ( n3585 , n2275 , n3518 );
    or g1556 ( n624 , n3255 , n3275 );
    or g1557 ( n502 , n1170 , n3290 );
    and g1558 ( n2577 , n2585 , n2917 );
    not g1559 ( n3132 , n2214 );
    or g1560 ( n2897 , n897 , n3152 );
    not g1561 ( n554 , n3105 );
    xnor g1562 ( n3486 , n2675 , n3269 );
    or g1563 ( n3002 , n3255 , n1509 );
    and g1564 ( n3144 , n2447 , n655 );
    or g1565 ( n3420 , n2161 , n1412 );
    or g1566 ( n729 , n2030 , n1413 );
    or g1567 ( n1967 , n3550 , n1235 );
    xnor g1568 ( n2902 , n219 , n2118 );
    or g1569 ( n1152 , n870 , n1198 );
    or g1570 ( n2306 , n2297 , n2792 );
    and g1571 ( n3591 , n1574 , n88 );
    and g1572 ( n2374 , n2297 , n2792 );
    or g1573 ( n3183 , n252 , n2655 );
    or g1574 ( n131 , n2855 , n28 );
    and g1575 ( n1017 , n191 , n1109 );
    nor g1576 ( n2409 , n3517 , n2265 );
    and g1577 ( n1879 , n2056 , n2808 );
    and g1578 ( n2284 , n1768 , n2523 );
    or g1579 ( n1221 , n2721 , n2047 );
    not g1580 ( n1368 , n1207 );
    or g1581 ( n3054 , n3616 , n1732 );
    or g1582 ( n2623 , n2220 , n891 );
    or g1583 ( n575 , n38 , n2671 );
    xnor g1584 ( n2749 , n155 , n1519 );
    or g1585 ( n973 , n844 , n2264 );
    not g1586 ( n2344 , n3160 );
    not g1587 ( n3666 , n1124 );
    or g1588 ( n1693 , n1270 , n3399 );
    xnor g1589 ( n2223 , n335 , n1537 );
    xnor g1590 ( n1012 , n6 , n1062 );
    and g1591 ( n393 , n2356 , n433 );
    or g1592 ( n2477 , n1552 , n2750 );
    not g1593 ( n845 , n3563 );
    or g1594 ( n3028 , n220 , n2484 );
    or g1595 ( n551 , n1878 , n647 );
    xnor g1596 ( n2155 , n3236 , n2635 );
    xnor g1597 ( n1808 , n3237 , n1023 );
    or g1598 ( n140 , n2158 , n2270 );
    or g1599 ( n989 , n2163 , n2492 );
    and g1600 ( n1462 , n708 , n2358 );
    xnor g1601 ( n1291 , n1835 , n273 );
    and g1602 ( n63 , n1485 , n3175 );
    or g1603 ( n2836 , n1231 , n3015 );
    xnor g1604 ( n2760 , n2067 , n3559 );
    or g1605 ( n2757 , n441 , n1334 );
    xnor g1606 ( n634 , n3330 , n1760 );
    or g1607 ( n3172 , n3326 , n453 );
    not g1608 ( n3371 , n2629 );
    and g1609 ( n2054 , n556 , n3382 );
    and g1610 ( n332 , n1097 , n279 );
    or g1611 ( n1564 , n1428 , n2077 );
    nor g1612 ( n177 , n78 , n1338 );
    or g1613 ( n2179 , n1096 , n1550 );
    xnor g1614 ( n1223 , n238 , n1209 );
    xnor g1615 ( n699 , n2173 , n2351 );
    or g1616 ( n1914 , n2600 , n522 );
    or g1617 ( n3497 , n2025 , n777 );
    nor g1618 ( n2027 , n2056 , n2808 );
    xnor g1619 ( n774 , n2109 , n1874 );
    or g1620 ( n1446 , n2291 , n2220 );
    not g1621 ( n1865 , n565 );
    or g1622 ( n3341 , n1769 , n2069 );
    xor g1623 ( n2405 , n936 , n1012 );
    xnor g1624 ( n1314 , n743 , n2106 );
    and g1625 ( n3199 , n2616 , n1300 );
    xnor g1626 ( n2986 , n828 , n3093 );
    nor g1627 ( n2431 , n511 , n3000 );
    or g1628 ( n10 , n2504 , n381 );
    or g1629 ( n82 , n3417 , n1015 );
    and g1630 ( n2611 , n242 , n3041 );
    xnor g1631 ( n2285 , n2544 , n2025 );
    or g1632 ( n2165 , n2526 , n1668 );
    xnor g1633 ( n2160 , n1196 , n454 );
    xnor g1634 ( n399 , n3437 , n233 );
    xnor g1635 ( n2876 , n533 , n3212 );
    xnor g1636 ( n256 , n1198 , n691 );
    or g1637 ( n3086 , n2648 , n3152 );
    and g1638 ( n2345 , n481 , n1696 );
    xnor g1639 ( n1031 , n2396 , n1127 );
    or g1640 ( n1937 , n1736 , n3668 );
    or g1641 ( n2419 , n787 , n213 );
    and g1642 ( n479 , n3197 , n642 );
    xnor g1643 ( n896 , n687 , n376 );
    and g1644 ( n2287 , n1218 , n2124 );
    or g1645 ( n1337 , n2819 , n3318 );
    and g1646 ( n2110 , n156 , n162 );
    and g1647 ( n2012 , n3062 , n2520 );
    xnor g1648 ( n809 , n1381 , n606 );
    and g1649 ( n2182 , n2806 , n1582 );
    xnor g1650 ( n22 , n1398 , n2404 );
    or g1651 ( n906 , n1310 , n2186 );
    xnor g1652 ( n2788 , n2019 , n1559 );
    xnor g1653 ( n768 , n3197 , n642 );
    or g1654 ( n621 , n457 , n2397 );
    not g1655 ( n31 , n3147 );
    xnor g1656 ( n3177 , n401 , n2828 );
    and g1657 ( n3243 , n3619 , n1910 );
    and g1658 ( n1843 , n1960 , n653 );
    or g1659 ( n2238 , n1486 , n2918 );
    and g1660 ( n3276 , n962 , n1114 );
    or g1661 ( n2375 , n323 , n2210 );
    and g1662 ( n1815 , n1722 , n2234 );
    and g1663 ( n3322 , n1294 , n3194 );
    xnor g1664 ( n2544 , n2240 , n2872 );
    not g1665 ( n3207 , n2680 );
    xnor g1666 ( n654 , n840 , n1378 );
    or g1667 ( n592 , n1871 , n329 );
    xnor g1668 ( n1585 , n1882 , n1379 );
    or g1669 ( n3481 , n3524 , n857 );
    or g1670 ( n540 , n2376 , n243 );
    not g1671 ( n64 , n924 );
    nor g1672 ( n1460 , n1113 , n2021 );
    nor g1673 ( n3493 , n3465 , n2005 );
    xnor g1674 ( n785 , n2500 , n3563 );
    xnor g1675 ( n907 , n1314 , n2101 );
    xor g1676 ( n3627 , n532 , n3215 );
    or g1677 ( n835 , n27 , n649 );
    nor g1678 ( n2505 , n379 , n3411 );
    not g1679 ( n1479 , n1860 );
    and g1680 ( n239 , n1124 , n610 );
    or g1681 ( n71 , n638 , n2933 );
    or g1682 ( n3635 , n2367 , n1283 );
    not g1683 ( n1864 , n881 );
    xnor g1684 ( n1997 , n2460 , n854 );
    xnor g1685 ( n3431 , n1878 , n1020 );
    xnor g1686 ( n1004 , n566 , n430 );
    xnor g1687 ( n678 , n2211 , n3114 );
    and g1688 ( n1445 , n2350 , n719 );
    not g1689 ( n1678 , n2789 );
    or g1690 ( n2549 , n219 , n2880 );
    xnor g1691 ( n91 , n1728 , n613 );
    or g1692 ( n2839 , n75 , n1262 );
    or g1693 ( n2793 , n1269 , n2263 );
    or g1694 ( n1732 , n3145 , n3316 );
    xnor g1695 ( n3179 , n2963 , n3446 );
    and g1696 ( n374 , n3412 , n1691 );
    nor g1697 ( n2184 , n3273 , n1108 );
    or g1698 ( n462 , n2558 , n2795 );
    or g1699 ( n1556 , n2881 , n2541 );
    not g1700 ( n1200 , n626 );
    and g1701 ( n1118 , n284 , n2335 );
    xnor g1702 ( n3453 , n3183 , n1888 );
    xnor g1703 ( n529 , n3072 , n2904 );
    or g1704 ( n1756 , n2396 , n2758 );
    or g1705 ( n1019 , n3546 , n3315 );
    or g1706 ( n3375 , n1851 , n2664 );
    or g1707 ( n3145 , n802 , n2508 );
    xnor g1708 ( n226 , n2455 , n2113 );
    and g1709 ( n2289 , n3133 , n2082 );
    and g1710 ( n2141 , n188 , n1709 );
    and g1711 ( n3494 , n3648 , n2593 );
    nor g1712 ( n528 , n167 , n2089 );
    not g1713 ( n740 , n1389 );
    xnor g1714 ( n98 , n1584 , n608 );
    and g1715 ( n1688 , n104 , n919 );
    or g1716 ( n3174 , n2030 , n2186 );
    nor g1717 ( n429 , n3081 , n2925 );
    or g1718 ( n601 , n38 , n189 );
    xnor g1719 ( n1626 , n3277 , n2850 );
    and g1720 ( n875 , n3320 , n2856 );
    and g1721 ( n635 , n631 , n163 );
    or g1722 ( n103 , n1310 , n554 );
    xnor g1723 ( n3464 , n3162 , n2166 );
    not g1724 ( n1100 , n737 );
    xnor g1725 ( n2174 , n707 , n450 );
    and g1726 ( n531 , n551 , n3294 );
    and g1727 ( n1653 , n1568 , n229 );
    or g1728 ( n2319 , n493 , n913 );
    or g1729 ( n2579 , n2163 , n1587 );
    and g1730 ( n359 , n1494 , n1916 );
    or g1731 ( n2118 , n1405 , n2010 );
    and g1732 ( n185 , n1565 , n850 );
    not g1733 ( n1527 , n390 );
    or g1734 ( n2606 , n1448 , n3635 );
    or g1735 ( n410 , n3191 , n1101 );
    xnor g1736 ( n1629 , n1168 , n2739 );
    xnor g1737 ( n54 , n1415 , n1538 );
    and g1738 ( n90 , n2539 , n36 );
    and g1739 ( n1677 , n3209 , n1387 );
    nor g1740 ( n4 , n998 , n1406 );
    or g1741 ( n1486 , n1552 , n2968 );
    or g1742 ( n182 , n1170 , n2830 );
    xnor g1743 ( n3598 , n1926 , n2728 );
    and g1744 ( n911 , n2357 , n1279 );
    not g1745 ( n217 , n2447 );
    or g1746 ( n2647 , n1204 , n3314 );
    xnor g1747 ( n2674 , n806 , n2764 );
    or g1748 ( n2266 , n2849 , n1352 );
    not g1749 ( n801 , n2476 );
    xor g1750 ( n3483 , n540 , n3037 );
    xnor g1751 ( n1387 , n1151 , n894 );
    or g1752 ( n3186 , n966 , n2610 );
    or g1753 ( n570 , n1428 , n2811 );
    or g1754 ( n1126 , n2163 , n495 );
    and g1755 ( n2939 , n1912 , n459 );
    xnor g1756 ( n1522 , n1363 , n2334 );
    xnor g1757 ( n892 , n519 , n62 );
    and g1758 ( n458 , n798 , n304 );
    or g1759 ( n2602 , n3326 , n1658 );
    nor g1760 ( n2985 , n1460 , n2162 );
    not g1761 ( n3391 , n2779 );
    xnor g1762 ( n1357 , n502 , n680 );
    and g1763 ( n1088 , n2864 , n2718 );
    xor g1764 ( n1279 , n63 , n3338 );
    or g1765 ( n2523 , n468 , n1963 );
    xnor g1766 ( n2263 , n2530 , n2986 );
    xnor g1767 ( n459 , n818 , n3570 );
    xnor g1768 ( n840 , n3399 , n1393 );
    xnor g1769 ( n1682 , n1891 , n2826 );
    and g1770 ( n2487 , n2637 , n3558 );
    xnor g1771 ( n527 , n524 , n586 );
    nor g1772 ( n1973 , n1505 , n2103 );
    or g1773 ( n1270 , n3293 , n2186 );
    not g1774 ( n3590 , n3682 );
    xnor g1775 ( n3090 , n3343 , n2848 );
    or g1776 ( n2028 , n3417 , n1992 );
    or g1777 ( n2032 , n1859 , n2977 );
    or g1778 ( n1159 , n1078 , n803 );
    xnor g1779 ( n2755 , n1581 , n2125 );
    or g1780 ( n2210 , n204 , n802 );
    and g1781 ( n1469 , n359 , n2054 );
    and g1782 ( n1091 , n3430 , n74 );
    or g1783 ( n1943 , n592 , n3405 );
    or g1784 ( n2916 , n2027 , n1404 );
    or g1785 ( n258 , n2163 , n2882 );
    or g1786 ( n427 , n148 , n1694 );
    or g1787 ( n3095 , n342 , n699 );
    not g1788 ( n1289 , n3608 );
    not g1789 ( n3667 , n3056 );
    or g1790 ( n530 , n466 , n2010 );
    xnor g1791 ( n3677 , n1997 , n1293 );
    and g1792 ( n94 , n3253 , n841 );
    xnor g1793 ( n3611 , n3539 , n2250 );
    xnor g1794 ( n3532 , n3653 , n724 );
    or g1795 ( n2835 , n2553 , n3267 );
    not g1796 ( n1763 , n2400 );
    xnor g1797 ( n2976 , n2797 , n995 );
    nor g1798 ( n3674 , n1852 , n478 );
    xnor g1799 ( n732 , n3604 , n169 );
    nor g1800 ( n2683 , n1301 , n1630 );
    and g1801 ( n1947 , n3351 , n2273 );
    or g1802 ( n1784 , n1842 , n2604 );
    and g1803 ( n2111 , n2213 , n524 );
    xnor g1804 ( n1383 , n1396 , n664 );
    and g1805 ( n822 , n14 , n3407 );
    and g1806 ( n1991 , n3539 , n2250 );
    xnor g1807 ( n1760 , n3438 , n1787 );
    or g1808 ( n3472 , n3550 , n2712 );
    xnor g1809 ( n2168 , n630 , n535 );
    or g1810 ( n1731 , n1364 , n1191 );
    or g1811 ( n2969 , n792 , n3214 );
    or g1812 ( n3397 , n1851 , n1334 );
    or g1813 ( n3324 , n1753 , n1974 );
    and g1814 ( n3046 , n192 , n3585 );
    or g1815 ( n3670 , n3096 , n18 );
    and g1816 ( n3212 , n278 , n2896 );
    xnor g1817 ( n2302 , n2332 , n1241 );
    or g1818 ( n2458 , n1987 , n3276 );
    or g1819 ( n2317 , n1851 , n1509 );
    or g1820 ( n848 , n2072 , n3072 );
    or g1821 ( n2660 , n1947 , n2785 );
    or g1822 ( n47 , n1127 , n1829 );
    xor g1823 ( n3554 , n3450 , n2449 );
    xnor g1824 ( n138 , n1224 , n3087 );
    or g1825 ( n990 , n2692 , n262 );
    and g1826 ( n3415 , n2570 , n1977 );
    nor g1827 ( n1436 , n234 , n432 );
    xnor g1828 ( n253 , n2091 , n3347 );
    nor g1829 ( n1499 , n1895 , n440 );
    xnor g1830 ( n1276 , n2241 , n179 );
    and g1831 ( n2528 , n1425 , n2028 );
    or g1832 ( n3104 , n959 , n190 );
    or g1833 ( n2796 , n2362 , n1868 );
    and g1834 ( n3201 , n2781 , n140 );
    nor g1835 ( n3556 , n3283 , n1253 );
    and g1836 ( n569 , n2567 , n520 );
    and g1837 ( n2166 , n1782 , n605 );
    not g1838 ( n1658 , n330 );
    xnor g1839 ( n1812 , n2892 , n1686 );
    and g1840 ( n2203 , n533 , n3597 );
    or g1841 ( n3340 , n45 , n2315 );
    xnor g1842 ( n1046 , n2917 , n2585 );
    and g1843 ( n739 , n160 , n2160 );
    or g1844 ( n1751 , n1309 , n624 );
    and g1845 ( n3038 , n3029 , n3676 );
    xnor g1846 ( n599 , n2049 , n2581 );
    not g1847 ( n2776 , n2444 );
    and g1848 ( n1570 , n2443 , n2644 );
    xnor g1849 ( n606 , n1481 , n2716 );
    xnor g1850 ( n1439 , n1949 , n3169 );
    not g1851 ( n1408 , n1264 );
    or g1852 ( n126 , n581 , n2671 );
    nor g1853 ( n1952 , n3215 , n532 );
    or g1854 ( n1890 , n1540 , n649 );
    or g1855 ( n2292 , n874 , n3429 );
    or g1856 ( n1184 , n3528 , n545 );
    nor g1857 ( n2050 , n770 , n3266 );
    xnor g1858 ( n2758 , n2253 , n3485 );
    and g1859 ( n1350 , n1920 , n3379 );
    or g1860 ( n717 , n1556 , n1581 );
    or g1861 ( n3213 , n1589 , n3035 );
    or g1862 ( n2308 , n53 , n2397 );
    not g1863 ( n1422 , n3557 );
    not g1864 ( n2291 , n1512 );
    xnor g1865 ( n2695 , n2107 , n347 );
    or g1866 ( n2366 , n1417 , n2565 );
    xnor g1867 ( n854 , n398 , n3490 );
    or g1868 ( n2226 , n1170 , n1015 );
    or g1869 ( n3111 , n2163 , n651 );
    not g1870 ( n1138 , n3413 );
    or g1871 ( n1211 , n3096 , n1235 );
    or g1872 ( n1189 , n1342 , n2241 );
    not g1873 ( n1801 , n648 );
    xnor g1874 ( n1219 , n89 , n2898 );
    or g1875 ( n626 , n1546 , n2458 );
    or g1876 ( n1498 , n2474 , n2883 );
    not g1877 ( n2938 , n3683 );
    or g1878 ( n753 , n1326 , n3229 );
    or g1879 ( n747 , n310 , n271 );
    and g1880 ( n790 , n2791 , n409 );
    and g1881 ( n3162 , n2959 , n3323 );
    xnor g1882 ( n679 , n2061 , n1045 );
    and g1883 ( n1050 , n3057 , n916 );
    or g1884 ( n3454 , n1405 , n1573 );
    xnor g1885 ( n1506 , n2510 , n2014 );
    xnor g1886 ( n2748 , n3670 , n2941 );
    xnor g1887 ( n378 , n588 , n2822 );
    or g1888 ( n1212 , n3506 , n795 );
    or g1889 ( n1822 , n2505 , n1502 );
    or g1890 ( n1285 , n698 , n2132 );
    and g1891 ( n2446 , n3340 , n1855 );
    and g1892 ( n803 , n2148 , n333 );
    or g1893 ( n1231 , n925 , n2750 );
    not g1894 ( n3377 , n1682 );
    and g1895 ( n311 , n2796 , n3620 );
    xnor g1896 ( n1662 , n1659 , n1444 );
    or g1897 ( n2365 , n3550 , n2671 );
    and g1898 ( n3297 , n3661 , n2574 );
    or g1899 ( n1501 , n1661 , n220 );
    or g1900 ( n959 , n1405 , n645 );
    xnor g1901 ( n500 , n1553 , n3532 );
    and g1902 ( n1873 , n3568 , n1562 );
    and g1903 ( n3158 , n2699 , n2227 );
    and g1904 ( n3047 , n960 , n3538 );
    xnor g1905 ( n2989 , n1717 , n1980 );
    xnor g1906 ( n2011 , n1291 , n458 );
    and g1907 ( n1375 , n2301 , n2666 );
    xnor g1908 ( n2932 , n1923 , n3625 );
    or g1909 ( n1161 , n3458 , n2554 );
    xnor g1910 ( n2300 , n1412 , n2161 );
    or g1911 ( n2239 , n3321 , n3120 );
    or g1912 ( n210 , n2374 , n69 );
    xnor g1913 ( n2837 , n3116 , n1004 );
    xnor g1914 ( n2728 , n1364 , n1191 );
    or g1915 ( n640 , n1680 , n2384 );
    not g1916 ( n3379 , n2745 );
    xnor g1917 ( n3561 , n1702 , n2610 );
    and g1918 ( n55 , n3418 , n1554 );
    xnor g1919 ( n1465 , n3472 , n1186 );
    or g1920 ( n2568 , n2522 , n226 );
    and g1921 ( n3386 , n3343 , n2848 );
    or g1922 ( n3310 , n104 , n919 );
    xnor g1923 ( n2613 , n3523 , n2349 );
    or g1924 ( n825 , n1395 , n201 );
    and g1925 ( n1508 , n3334 , n3368 );
    or g1926 ( n1757 , n1481 , n2716 );
    or g1927 ( n2520 , n3142 , n623 );
    or g1928 ( n88 , n3116 , n1889 );
    and g1929 ( n2244 , n1572 , n1174 );
    or g1930 ( n3016 , n307 , n2012 );
    xnor g1931 ( n1715 , n2176 , n1462 );
    xnor g1932 ( n3241 , n912 , n1449 );
    xnor g1933 ( n3675 , n1139 , n240 );
    nor g1934 ( n2994 , n538 , n314 );
    xnor g1935 ( n3147 , n1163 , n2495 );
    not g1936 ( n1307 , n2582 );
    xnor g1937 ( n1609 , n3421 , n2919 );
    xnor g1938 ( n3643 , n555 , n3187 );
    or g1939 ( n296 , n583 , n595 );
    or g1940 ( n3637 , n2725 , n2752 );
    or g1941 ( n2941 , n2696 , n34 );
    or g1942 ( n1568 , n1898 , n445 );
    or g1943 ( n1224 , n2819 , n2397 );
    or g1944 ( n3226 , n2220 , n78 );
    or g1945 ( n95 , n3209 , n1387 );
    or g1946 ( n2574 , n38 , n34 );
    not g1947 ( n3157 , n1423 );
    or g1948 ( n386 , n983 , n986 );
    nor g1949 ( n395 , n3064 , n490 );
    and g1950 ( n1037 , n3404 , n138 );
    xnor g1951 ( n2318 , n3029 , n437 );
    or g1952 ( n585 , n3123 , n3233 );
    and g1953 ( n1026 , n2892 , n1267 );
    xnor g1954 ( n3342 , n1605 , n3455 );
    and g1955 ( n2371 , n2576 , n843 );
    or g1956 ( n2543 , n2220 , n3469 );
    not g1957 ( n2124 , n2603 );
    xnor g1958 ( n2919 , n915 , n3102 );
    not g1959 ( n3096 , n1543 );
    or g1960 ( n1794 , n2402 , n485 );
    or g1961 ( n2570 , n2775 , n799 );
    and g1962 ( n871 , n2710 , n3508 );
    and g1963 ( n328 , n2331 , n2749 );
    and g1964 ( n342 , n1731 , n738 );
    xnor g1965 ( n1935 , n2480 , n865 );
    xnor g1966 ( n3684 , n3233 , n3123 );
    not g1967 ( n1772 , n2863 );
    and g1968 ( n3518 , n3455 , n1605 );
    xnor g1969 ( n2069 , n986 , n2751 );
    or g1970 ( n1284 , n2108 , n2383 );
    or g1971 ( n1014 , n177 , n547 );
    and g1972 ( n716 , n231 , n2008 );
    not g1973 ( n3246 , n597 );
    or g1974 ( n1153 , n563 , n2502 );
    xnor g1975 ( n629 , n3517 , n3381 );
    or g1976 ( n1273 , n2743 , n1445 );
    and g1977 ( n935 , n3250 , n2119 );
    nor g1978 ( n2928 , n519 , n392 );
    not g1979 ( n3063 , n2687 );
    xnor g1980 ( n2106 , n3220 , n712 );
    or g1981 ( n2617 , n38 , n2712 );
    xnor g1982 ( n2546 , n751 , n530 );
    not g1983 ( n3499 , n302 );
    xnor g1984 ( n971 , n1296 , n1939 );
    or g1985 ( n784 , n2753 , n2372 );
    or g1986 ( n2064 , n487 , n2489 );
    xnor g1987 ( n2739 , n1765 , n1906 );
    xnor g1988 ( n3584 , n2823 , n92 );
    or g1989 ( n344 , n2665 , n3084 );
    not g1990 ( n2234 , n3358 );
    and g1991 ( n1423 , n1470 , n1360 );
    xnor g1992 ( n3568 , n2021 , n1113 );
    nor g1993 ( n1319 , n3147 , n3416 );
    not g1994 ( n1851 , n728 );
    or g1995 ( n1572 , n38 , n18 );
    nor g1996 ( n2501 , n3546 , n3008 );
    or g1997 ( n2017 , n2569 , n1801 );
    or g1998 ( n2221 , n1661 , n1801 );
    or g1999 ( n2120 , n1537 , n808 );
    and g2000 ( n2987 , n3258 , n1791 );
    and g2001 ( n2445 , n3 , n1371 );
    or g2002 ( n623 , n2220 , n2745 );
    or g2003 ( n642 , n1661 , n2397 );
    xnor g2004 ( n3513 , n1764 , n1938 );
    and g2005 ( n2715 , n1556 , n1581 );
    and g2006 ( n181 , n3005 , n484 );
    or g2007 ( n3376 , n3426 , n2715 );
    or g2008 ( n1097 , n3237 , n54 );
    xnor g2009 ( n984 , n2717 , n1827 );
    not g2010 ( n18 , n1067 );
    and g2011 ( n3478 , n3207 , n2296 );
    not g2012 ( n2535 , n2232 );
    xnor g2013 ( n2130 , n633 , n2667 );
    or g2014 ( n92 , n797 , n2863 );
    and g2015 ( n2268 , n3587 , n2455 );
    xnor g2016 ( n2483 , n1681 , n1158 );
    or g2017 ( n366 , n2757 , n311 );
    and g2018 ( n495 , n3182 , n2478 );
    and g2019 ( n2467 , n2491 , n2639 );
    xnor g2020 ( n2996 , n306 , n1030 );
    not g2021 ( n561 , n3644 );
    or g2022 ( n3244 , n1661 , n3634 );
    and g2023 ( n791 , n1343 , n979 );
    xnor g2024 ( n3081 , n496 , n361 );
    and g2025 ( n1166 , n2072 , n3072 );
    xnor g2026 ( n3610 , n855 , n315 );
    or g2027 ( n310 , n2696 , n2671 );
    or g2028 ( n3148 , n3595 , n436 );
    or g2029 ( n3339 , n1851 , n1648 );
    or g2030 ( n3651 , n2284 , n1061 );
    or g2031 ( n2869 , n581 , n955 );
    or g2032 ( n1813 , n3002 , n1348 );
    or g2033 ( n246 , n2142 , n2485 );
    xnor g2034 ( n2354 , n2145 , n1204 );
    or g2035 ( n2742 , n12 , n194 );
    xnor g2036 ( n2903 , n1766 , n1915 );
    or g2037 ( n697 , n2652 , n3184 );
    or g2038 ( n1280 , n1595 , n2514 );
    or g2039 ( n2453 , n695 , n1459 );
    nor g2040 ( n1362 , n2023 , n2322 );
    or g2041 ( n486 , n1710 , n2799 );
    nor g2042 ( n636 , n3133 , n2082 );
    or g2043 ( n283 , n3591 , n2469 );
    xnor g2044 ( n1477 , n493 , n2995 );
    xnor g2045 ( n982 , n2806 , n3181 );
    and g2046 ( n3037 , n3657 , n115 );
    or g2047 ( n2410 , n1054 , n2397 );
    or g2048 ( n3101 , n486 , n2135 );
    and g2049 ( n2202 , n3163 , n657 );
    xnor g2050 ( n2823 , n3257 , n2405 );
    or g2051 ( n1165 , n2535 , n2489 );
    or g2052 ( n2373 , n2237 , n1250 );
    or g2053 ( n465 , n2696 , n18 );
    or g2054 ( n2761 , n2970 , n141 );
    or g2055 ( n1507 , n193 , n887 );
    or g2056 ( n2443 , n1701 , n989 );
    and g2057 ( n1941 , n365 , n1849 );
    or g2058 ( n622 , n1981 , n875 );
    nor g2059 ( n2150 , n2309 , n2426 );
    or g2060 ( n3328 , n715 , n3586 );
    or g2061 ( n17 , n2220 , n2467 );
    xnor g2062 ( n2307 , n3161 , n3516 );
    or g2063 ( n430 , n1170 , n1992 );
    or g2064 ( n3504 , n1987 , n1983 );
    or g2065 ( n969 , n901 , n3650 );
    or g2066 ( n2688 , n2569 , n1573 );
    or g2067 ( n2014 , n1170 , n3152 );
    xnor g2068 ( n1897 , n1238 , n2948 );
    or g2069 ( n2457 , n2615 , n329 );
    xnor g2070 ( n72 , n3616 , n1716 );
    and g2071 ( n721 , n469 , n2746 );
    and g2072 ( n1713 , n3385 , n3477 );
    not g2073 ( n1472 , n1194 );
    xnor g2074 ( n3530 , n856 , n3158 );
    or g2075 ( n991 , n231 , n2008 );
    and g2076 ( n2514 , n415 , n1988 );
    and g2077 ( n3029 , n463 , n2624 );
    xnor g2078 ( n3681 , n1803 , n3061 );
    or g2079 ( n707 , n671 , n1750 );
    not g2080 ( n1802 , n653 );
    and g2081 ( n705 , n2510 , n1890 );
    and g2082 ( n1950 , n2340 , n1617 );
    and g2083 ( n2956 , n48 , n820 );
    or g2084 ( n2820 , n2748 , n755 );
    or g2085 ( n884 , n2168 , n2314 );
    and g2086 ( n3282 , n3231 , n1933 );
    nor g2087 ( n1742 , n3422 , n1673 );
    and g2088 ( n312 , n1089 , n2702 );
    or g2089 ( n2055 , n1873 , n385 );
    and g2090 ( n3259 , n1507 , n2501 );
    or g2091 ( n1711 , n2865 , n2038 );
    or g2092 ( n1494 , n2221 , n1316 );
    not g2093 ( n1315 , n765 );
    xnor g2094 ( n899 , n1522 , n3127 );
    not g2095 ( n2955 , n3582 );
    or g2096 ( n2136 , n3272 , n1509 );
    or g2097 ( n514 , n793 , n2433 );
    or g2098 ( n2393 , n350 , n2302 );
    and g2099 ( n933 , n1649 , n2817 );
    or g2100 ( n2909 , n922 , n332 );
    xnor g2101 ( n811 , n737 , n1443 );
    or g2102 ( n798 , n2835 , n2326 );
    or g2103 ( n980 , n1897 , n1128 );
    xnor g2104 ( n2842 , n646 , n2081 );
    xnor g2105 ( n1911 , n2901 , n3234 );
    not g2106 ( n2920 , n1913 );
    and g2107 ( n3153 , n1866 , n1374 );
    nor g2108 ( n724 , n1428 , n2438 );
    and g2109 ( n2780 , n3533 , n449 );
    xnor g2110 ( n512 , n846 , n2498 );
    xnor g2111 ( n1839 , n1762 , n2551 );
    and g2112 ( n437 , n2114 , n3019 );
    or g2113 ( n2105 , n3122 , n3574 );
    xnor g2114 ( n1058 , n313 , n947 );
    or g2115 ( n2250 , n1073 , n2968 );
    and g2116 ( n3180 , n1103 , n3031 );
    and g2117 ( n534 , n3108 , n3651 );
    xnor g2118 ( n1955 , n336 , n583 );
    not g2119 ( n490 , n1306 );
    xnor g2120 ( n1607 , n452 , n869 );
    or g2121 ( n2960 , n1419 , n3033 );
    or g2122 ( n373 , n2254 , n1453 );
    or g2123 ( n2076 , n3546 , n2369 );
    xnor g2124 ( n1931 , n28 , n3344 );
    or g2125 ( n2541 , n2753 , n3208 );
    and g2126 ( n538 , n269 , n873 );
    or g2127 ( n1683 , n1851 , n3275 );
    xor g2128 ( n518 , n1330 , n2343 );
    xnor g2129 ( n2343 , n517 , n2831 );
    and g2130 ( n230 , n130 , n1159 );
    or g2131 ( n2441 , n1987 , n285 );
    and g2132 ( n563 , n938 , n572 );
    or g2133 ( n163 , n1372 , n1921 );
    or g2134 ( n846 , n2096 , n453 );
    or g2135 ( n1461 , n2096 , n1658 );
    xnor g2136 ( n1893 , n116 , n2325 );
    and g2137 ( n2522 , n1414 , n2647 );
    or g2138 ( n1292 , n3347 , n3188 );
    or g2139 ( n877 , n3354 , n2955 );
    xnor g2140 ( n3021 , n1696 , n1155 );
    xnor g2141 ( n2942 , n726 , n1971 );
    or g2142 ( n2241 , n2088 , n68 );
    xnor g2143 ( n48 , n822 , n971 );
    nor g2144 ( n1842 , n1983 , n1201 );
    and g2145 ( n546 , n1647 , n2337 );
    xnor g2146 ( n719 , n3456 , n1730 );
    nor g2147 ( n1738 , n2609 , n3284 );
    and g2148 ( n2881 , n2300 , n2636 );
    and g2149 ( n2112 , n855 , n1885 );
    or g2150 ( n391 , n3601 , n2916 );
    or g2151 ( n1669 , n2220 , n1327 );
    and g2152 ( n700 , n839 , n1786 );
    xnor g2153 ( n954 , n2659 , n2298 );
    nor g2154 ( n2999 , n3023 , n1718 );
    and g2155 ( n2882 , n3023 , n1718 );
    or g2156 ( n588 , n2291 , n1648 );
    xnor g2157 ( n3563 , n2464 , n1532 );
    not g2158 ( n2734 , n1049 );
    or g2159 ( n3679 , n1441 , n1158 );
    xor g2160 ( n962 , n158 , n2257 );
    and g2161 ( n826 , n137 , n1689 );
    or g2162 ( n2802 , n1635 , n2043 );
    or g2163 ( n979 , n3167 , n3281 );
    or g2164 ( n2249 , n3552 , n1504 );
    or g2165 ( n475 , n2452 , n2929 );
    not g2166 ( n3134 , n326 );
    and g2167 ( n3447 , n769 , n984 );
    xnor g2168 ( n686 , n191 , n1109 );
    not g2169 ( n2293 , n420 );
    and g2170 ( n1344 , n1408 , n763 );
    or g2171 ( n129 , n3204 , n1497 );
    and g2172 ( n2745 , n2894 , n1488 );
    or g2173 ( n1195 , n2696 , n2712 );
    and g2174 ( n3187 , n2479 , n1280 );
    or g2175 ( n2785 , n2753 , n2178 );
    and g2176 ( n2077 , n1407 , n1603 );
    not g2177 ( n645 , n1948 );
    and g2178 ( n2912 , n1431 , n3007 );
    and g2179 ( n264 , n1978 , n1024 );
    and g2180 ( n1454 , n707 , n450 );
    or g2181 ( n488 , n3298 , n102 );
    xnor g2182 ( n2056 , n7 , n1090 );
    or g2183 ( n2618 , n3403 , n1223 );
    or g2184 ( n2245 , n2107 , n2991 );
    xnor g2185 ( n2979 , n3605 , n2989 );
    not g2186 ( n213 , n3144 );
    xnor g2187 ( n1959 , n2685 , n2803 );
    or g2188 ( n320 , n3488 , n904 );
    not g2189 ( n38 , n1660 );
    xnor g2190 ( n1331 , n3000 , n881 );
    or g2191 ( n1774 , n3410 , n1909 );
    or g2192 ( n2832 , n2893 , n1663 );
    or g2193 ( n950 , n2613 , n1837 );
    and g2194 ( n1863 , n3656 , n1290 );
    and g2195 ( n610 , n585 , n2776 );
    or g2196 ( n1975 , n2979 , n3509 );
    or g2197 ( n3661 , n173 , n18 );
    and g2198 ( n1336 , n3246 , n2777 );
    xnor g2199 ( n1979 , n1714 , n774 );
    and g2200 ( n3129 , n1628 , n1225 );
    xnor g2201 ( n3190 , n3025 , n1675 );
    xnor g2202 ( n2217 , n3045 , n224 );
    or g2203 ( n287 , n3553 , n1570 );
    and g2204 ( n1840 , n1074 , n2099 );
    and g2205 ( n197 , n358 , n2214 );
    xnor g2206 ( n1272 , n3334 , n3368 );
    not g2207 ( n443 , n3208 );
    xnor g2208 ( n600 , n3553 , n3624 );
    or g2209 ( n994 , n2553 , n24 );
    or g2210 ( n133 , n3511 , n3227 );
    not g2211 ( n1488 , n3047 );
    or g2212 ( n3080 , n733 , n923 );
    or g2213 ( n1414 , n1259 , n1366 );
    and g2214 ( n2493 , n931 , n2951 );
    or g2215 ( n1628 , n846 , n2602 );
    and g2216 ( n499 , n475 , n1836 );
    and g2217 ( n343 , n35 , n1196 );
    or g2218 ( n414 , n3287 , n527 );
    xnor g2219 ( n1296 , n1461 , n3643 );
    or g2220 ( n1694 , n2946 , n3275 );
    or g2221 ( n1029 , n2819 , n645 );
    or g2222 ( n666 , n2892 , n1267 );
    nor g2223 ( n1619 , n1121 , n2019 );
    and g2224 ( n1238 , n391 , n2653 );
    or g2225 ( n1926 , n897 , n1992 );
    or g2226 ( n1258 , n2669 , n3360 );
    xnor g2227 ( n2654 , n2378 , n767 );
    not g2228 ( n2486 , n2996 );
    not g2229 ( n1770 , n2599 );
    xnor g2230 ( n2279 , n1910 , n2552 );
    not g2231 ( n198 , n838 );
    or g2232 ( n1493 , n1527 , n1783 );
    or g2233 ( n664 , n1495 , n1039 );
    nor g2234 ( n338 , n327 , n1827 );
    or g2235 ( n3599 , n2615 , n2489 );
    or g2236 ( n2744 , n3202 , n2671 );
    and g2237 ( n2651 , n568 , n740 );
    or g2238 ( n843 , n3193 , n2638 );
    or g2239 ( n3473 , n441 , n2664 );
    xnor g2240 ( n1721 , n3482 , n778 );
    xnor g2241 ( n2472 , n2720 , n1964 );
    xnor g2242 ( n2845 , n1406 , n998 );
    and g2243 ( n2605 , n1999 , n155 );
    or g2244 ( n2719 , n204 , n2750 );
    xnor g2245 ( n1998 , n2950 , n3012 );
    xnor g2246 ( n368 , n835 , n3251 );
    and g2247 ( n904 , n1135 , n1822 );
    xnor g2248 ( n1313 , n859 , n1000 );
    or g2249 ( n1147 , n2118 , n2935 );
    xnor g2250 ( n2764 , n1370 , n3513 );
    or g2251 ( n799 , n2753 , n2821 );
    and g2252 ( n1761 , n2584 , n1254 );
    xnor g2253 ( n3295 , n3429 , n3592 );
    or g2254 ( n1225 , n2448 , n2498 );
    xnor g2255 ( n1321 , n1812 , n324 );
    xnor g2256 ( n2547 , n2784 , n37 );
    or g2257 ( n1634 , n456 , n946 );
    and g2258 ( n3039 , n2721 , n2047 );
    or g2259 ( n548 , n3025 , n2418 );
    and g2260 ( n1957 , n2371 , n3604 );
    or g2261 ( n713 , n53 , n1573 );
    xnor g2262 ( n2826 , n3271 , n563 );
    not g2263 ( n345 , n1111 );
    xnor g2264 ( n2917 , n1417 , n1729 );
    or g2265 ( n248 , n3244 , n2591 );
    or g2266 ( n3596 , n2934 , n1993 );
    not g2267 ( n1338 , n3361 );
    xnor g2268 ( n2169 , n1834 , n3265 );
    or g2269 ( n452 , n851 , n2233 );
    nor g2270 ( n1295 , n1765 , n1205 );
    or g2271 ( n3050 , n1824 , n2037 );
    xor g2272 ( n193 , n234 , n432 );
    or g2273 ( n2580 , n2683 , n594 );
    not g2274 ( n1235 , n2029 );
    and g2275 ( n519 , n1634 , n296 );
    xnor g2276 ( n2633 , n3468 , n2347 );
    and g2277 ( n1217 , n1033 , n1184 );
    xnor g2278 ( n3668 , n1430 , n1990 );
    or g2279 ( n1363 , n1898 , n1015 );
    xnor g2280 ( n107 , n721 , n2643 );
    or g2281 ( n1969 , n2166 , n3162 );
    or g2282 ( n1836 , n3655 , n2007 );
    or g2283 ( n3135 , n3293 , n2489 );
    or g2284 ( n521 , n1552 , n2294 );
    and g2285 ( n1342 , n3010 , n2965 );
    and g2286 ( n2684 , n1014 , n600 );
    and g2287 ( n823 , n389 , n1273 );
    not g2288 ( n327 , n2717 );
    not g2289 ( n1243 , n2073 );
    or g2290 ( n2624 , n3372 , n143 );
    and g2291 ( n1474 , n2429 , n840 );
    nor g2292 ( n876 , n2216 , n165 );
    or g2293 ( n1247 , n1491 , n203 );
    or g2294 ( n1473 , n2535 , n2186 );
    and g2295 ( n1379 , n61 , n423 );
    or g2296 ( n3467 , n404 , n2926 );
    and g2297 ( n3312 , n2558 , n2795 );
    and g2298 ( n1335 , n681 , n1524 );
    or g2299 ( n2852 , n838 , n1315 );
    or g2300 ( n223 , n972 , n1324 );
    or g2301 ( n2357 , n1347 , n3444 );
    or g2302 ( n1854 , n581 , n34 );
    xnor g2303 ( n2075 , n3574 , n1179 );
    or g2304 ( n2931 , n191 , n1109 );
    and g2305 ( n1389 , n749 , n205 );
    xnor g2306 ( n3278 , n2864 , n2949 );
    or g2307 ( n1641 , n2657 , n363 );
    or g2308 ( n672 , n1526 , n3654 );
    or g2309 ( n3657 , n444 , n1312 );
    xnor g2310 ( n2676 , n1600 , n58 );
    not g2311 ( n445 , n660 );
    or g2312 ( n1033 , n3177 , n256 );
    or g2313 ( n1917 , n1967 , n1048 );
    or g2314 ( n2119 , n745 , n170 );
    and g2315 ( n3446 , n3126 , n1390 );
    and g2316 ( n3161 , n2208 , n3352 );
    or g2317 ( n3242 , n3222 , n721 );
    and g2318 ( n3082 , n3438 , n3330 );
    or g2319 ( n889 , n3265 , n2937 );
    or g2320 ( n1351 , n3012 , n383 );
    nor g2321 ( n3466 , n1120 , n1790 );
    or g2322 ( n1202 , n2313 , n1949 );
    or g2323 ( n3181 , n1073 , n1658 );
    nor g2324 ( n2088 , n892 , n1047 );
    or g2325 ( n3026 , n424 , n2225 );
    xnor g2326 ( n533 , n2346 , n1185 );
    xnor g2327 ( n3506 , n3296 , n121 );
    xnor g2328 ( n2462 , n126 , n3526 );
    and g2329 ( n3119 , n2861 , n1167 );
    not g2330 ( n1008 , n1350 );
    or g2331 ( n1042 , n2378 , n2688 );
    and g2332 ( n814 , n337 , n3151 );
    xnor g2333 ( n3084 , n2047 , n2847 );
    or g2334 ( n503 , n3248 , n1509 );
    or g2335 ( n2600 , n1310 , n1413 );
    xnor g2336 ( n3624 , n2644 , n2443 );
    xnor g2337 ( n1266 , n2428 , n132 );
    not g2338 ( n2548 , n2951 );
    xnor g2339 ( n2512 , n195 , n2546 );
    or g2340 ( n1457 , n418 , n2464 );
    not g2341 ( n2321 , n1588 );
    not g2342 ( n3304 , n3440 );
    or g2343 ( n1099 , n999 , n2577 );
    or g2344 ( n3613 , n1133 , n174 );
    or g2345 ( n2264 , n1819 , n1260 );
    and g2346 ( n1755 , n1119 , n653 );
    xnor g2347 ( n1664 , n2804 , n2766 );
    xnor g2348 ( n781 , n2079 , n3598 );
    or g2349 ( n1234 , n465 , n2462 );
    and g2350 ( n559 , n1534 , n3579 );
    xnor g2351 ( n3319 , n1 , n2538 );
    or g2352 ( n3682 , n2768 , n1449 );
    and g2353 ( n2142 , n1774 , n89 );
    or g2354 ( n3645 , n1170 , n1707 );
    or g2355 ( n3468 , n1054 , n645 );
    or g2356 ( n2398 , n2753 , n1860 );
    and g2357 ( n3265 , n1212 , n2923 );
    and g2358 ( n659 , n326 , n3557 );
    not g2359 ( n1529 , n775 );
    or g2360 ( n153 , n3615 , n1243 );
    not g2361 ( n349 , n1090 );
    and g2362 ( n2025 , n1757 , n3369 );
    and g2363 ( n776 , n1899 , n557 );
    and g2364 ( n3008 , n193 , n887 );
    or g2365 ( n883 , n714 , n3384 );
    or g2366 ( n2071 , n1820 , n1037 );
    xnor g2367 ( n3060 , n1452 , n2199 );
    or g2368 ( n1456 , n1240 , n2274 );
    or g2369 ( n1740 , n3270 , n2971 );
    and g2370 ( n432 , n727 , n2116 );
    not g2371 ( n1054 , n3430 );
    or g2372 ( n2194 , n2173 , n3140 );
    or g2373 ( n362 , n3272 , n2664 );
    not g2374 ( n348 , n1366 );
    not g2375 ( n3540 , n153 );
    and g2376 ( n3043 , n3238 , n2188 );
    or g2377 ( n2889 , n3659 , n1766 );
    and g2378 ( n504 , n3422 , n1673 );
    xor g2379 ( n3085 , n486 , n945 );
    or g2380 ( n2766 , n3272 , n1648 );
    and g2381 ( n1288 , n2878 , n117 );
    xnor g2382 ( n1610 , n1886 , n2562 );
    and g2383 ( n1192 , n2640 , n1389 );
    and g2384 ( n305 , n3311 , n3124 );
    or g2385 ( n3256 , n2555 , n1337 );
    or g2386 ( n734 , n27 , n3152 );
    xnor g2387 ( n926 , n1061 , n60 );
    xnor g2388 ( n1685 , n3621 , n2913 );
    xnor g2389 ( n121 , n2626 , n1517 );
    or g2390 ( n681 , n1723 , n3051 );
    not g2391 ( n830 , n899 );
    xnor g2392 ( n537 , n1568 , n3671 );
    or g2393 ( n2107 , n2569 , n2397 );
    or g2394 ( n2147 , n489 , n704 );
    xnor g2395 ( n1828 , n634 , n1789 );
    not g2396 ( n1648 , n407 );
    or g2397 ( n114 , n1142 , n1996 );
    and g2398 ( n298 , n503 , n1139 );
    or g2399 ( n2009 , n53 , n1801 );
    and g2400 ( n644 , n3544 , n510 );
    xnor g2401 ( n2187 , n3543 , n618 );
    or g2402 ( n2679 , n580 , n3495 );
    and g2403 ( n1581 , n3373 , n2421 );
    and g2404 ( n352 , n1270 , n3399 );
    xnor g2405 ( n316 , n362 , n513 );
    xnor g2406 ( n2540 , n2230 , n1503 );
    xnor g2407 ( n993 , n1312 , n1416 );
    or g2408 ( n873 , n3037 , n2879 );
    and g2409 ( n301 , n2936 , n903 );
    and g2410 ( n2689 , n3401 , n3599 );
    or g2411 ( n824 , n897 , n649 );
    and g2412 ( n2730 , n1656 , n2924 );
    or g2413 ( n1523 , n3096 , n2163 );
    or g2414 ( n821 , n3454 , n3475 );
    xnor g2415 ( n2643 , n3222 , n1058 );
    xnor g2416 ( n999 , n2031 , n3614 );
    or g2417 ( n3525 , n2967 , n1593 );
    xnor g2418 ( n2851 , n1326 , n1439 );
    or g2419 ( n1928 , n3656 , n1290 );
    or g2420 ( n2626 , n1372 , n18 );
    xnor g2421 ( n3607 , n2020 , n500 );
    and g2422 ( n1598 , n1623 , n3186 );
    nor g2423 ( n1546 , n962 , n1114 );
    and g2424 ( n2725 , n2723 , n2897 );
    xnor g2425 ( n2224 , n620 , n3036 );
    xnor g2426 ( n1553 , n1706 , n3013 );
    xnor g2427 ( n358 , n3577 , n2017 );
    or g2428 ( n779 , n2791 , n409 );
    or g2429 ( n1604 , n3263 , n3286 );
    and g2430 ( n1093 , n835 , n3251 );
    nor g2431 ( n3078 , n2276 , n1931 );
    xnor g2432 ( n3237 , n1890 , n1506 );
    and g2433 ( n1128 , n3230 , n3409 );
    nor g2434 ( n2023 , n1000 , n859 );
    or g2435 ( n3384 , n1987 , n2202 );
    or g2436 ( n52 , n1430 , n96 );
    and g2437 ( n3264 , n2829 , n1600 );
    xnor g2438 ( n444 , n2376 , n243 );
    and g2439 ( n3098 , n3211 , n3131 );
    not g2440 ( n457 , n3141 );
    not g2441 ( n3051 , n1817 );
    not g2442 ( n293 , n2332 );
    or g2443 ( n1625 , n2518 , n3541 );
    xnor g2444 ( n893 , n766 , n276 );
    xnor g2445 ( n1850 , n229 , n537 );
    and g2446 ( n2047 , n1777 , n108 );
    xnor g2447 ( n3076 , n1380 , n3274 );
    and g2448 ( n992 , n3263 , n3286 );
    or g2449 ( n2497 , n1908 , n1217 );
    and g2450 ( n2716 , n2 , n106 );
    and g2451 ( n587 , n2841 , n2407 );
    xnor g2452 ( n32 , n3192 , n742 );
    and g2453 ( n3336 , n3054 , n2456 );
    or g2454 ( n737 , n2045 , n2623 );
    not g2455 ( n3255 , n1676 );
    or g2456 ( n447 , n3296 , n2980 );
    not g2457 ( n1780 , n2115 );
    or g2458 ( n1841 , n1428 , n3070 );
    nor g2459 ( n19 , n7 , n349 );
    or g2460 ( n3298 , n2033 , n1841 );
    and g2461 ( n1622 , n3256 , n3104 );
    and g2462 ( n914 , n2741 , n567 );
    not g2463 ( n2096 , n3302 );
    and g2464 ( n1819 , n2551 , n2907 );
    or g2465 ( n1620 , n3521 , n2755 );
    not g2466 ( n2309 , n1165 );
    and g2467 ( n2754 , n2260 , n1016 );
    and g2468 ( n3205 , n1098 , n720 );
    and g2469 ( n3053 , n2748 , n755 );
    not g2470 ( n972 , n2468 );
    xnor g2471 ( n857 , n1284 , n2722 );
    xnor g2472 ( n1252 , n2780 , n2293 );
    or g2473 ( n958 , n2958 , n259 );
    and g2474 ( n929 , n3216 , n2304 );
    or g2475 ( n1551 , n2272 , n1068 );
    and g2476 ( n1186 , n2733 , n1351 );
    nor g2477 ( n525 , n3322 , n2360 );
    and g2478 ( n670 , n2983 , n694 );
    and g2479 ( n2993 , n2375 , n114 );
    not g2480 ( n1783 , n2496 );
    nor g2481 ( n641 , n921 , n3148 );
    or g2482 ( n1920 , n2760 , n2840 );
    or g2483 ( n1502 , n3546 , n1111 );
    xnor g2484 ( n2525 , n3068 , n1664 );
    not g2485 ( n2849 , n3045 );
    and g2486 ( n2775 , n954 , n1815 );
    xnor g2487 ( n3434 , n1712 , n2660 );
    or g2488 ( n2733 , n2950 , n1329 );
    or g2489 ( n1425 , n27 , n445 );
    not g2490 ( n2857 , n461 );
    or g2491 ( n2816 , n549 , n2815 );
    not g2492 ( n3423 , n1385 );
    or g2493 ( n323 , n1631 , n2750 );
    xnor g2494 ( n725 , n2373 , n3281 );
    or g2495 ( n1041 , n482 , n2078 );
    or g2496 ( n3648 , n812 , n1219 );
    and g2497 ( n2385 , n588 , n2822 );
    and g2498 ( n1246 , n2187 , n2352 );
    xnor g2499 ( n676 , n797 , n1772 );
    and g2500 ( n214 , n1342 , n2241 );
    and g2501 ( n820 , n2953 , n1667 );
    or g2502 ( n723 , n3223 , n2740 );
    and g2503 ( n1262 , n451 , n1060 );
    or g2504 ( n1075 , n1163 , n871 );
    xnor g2505 ( n1092 , n12 , n194 );
    xnor g2506 ( n1397 , n2277 , n1199 );
    not g2507 ( n2814 , n3578 );
    or g2508 ( n241 , n925 , n24 );
    or g2509 ( n3195 , n1834 , n3350 );
    and g2510 ( n602 , n1781 , n3575 );
    not g2511 ( n506 , n442 );
    xnor g2512 ( n2113 , n3587 , n87 );
    or g2513 ( n2117 , n863 , n2939 );
    or g2514 ( n3359 , n2243 , n3564 );
    and g2515 ( n1255 , n3618 , n2256 );
    or g2516 ( n1332 , n2499 , n2211 );
    or g2517 ( n1435 , n128 , n2489 );
    or g2518 ( n247 , n2040 , n369 );
    xnor g2519 ( n1496 , n1070 , n3160 );
    not g2520 ( n1650 , n1255 );
    or g2521 ( n3066 , n3449 , n678 );
    or g2522 ( n2533 , n1310 , n2233 );
    or g2523 ( n3609 , n3293 , n1138 );
    or g2524 ( n1005 , n2430 , n961 );
    and g2525 ( n1116 , n534 , n2032 );
    xnor g2526 ( n1923 , n1169 , n734 );
    and g2527 ( n861 , n917 , n81 );
    not g2528 ( n3579 , n1708 );
    xnor g2529 ( n314 , n2130 , n1122 );
    and g2530 ( n2129 , n2534 , n360 );
    nor g2531 ( n988 , n1864 , n2618 );
    not g2532 ( n205 , n2475 );
    not g2533 ( n2890 , n1752 );
    xnor g2534 ( n3381 , n1149 , n2417 );
    or g2535 ( n1390 , n2754 , n1918 );
    or g2536 ( n1047 , n29 , n2202 );
    not g2537 ( n299 , n3416 );
    or g2538 ( n2947 , n1631 , n802 );
    and g2539 ( n745 , n421 , n1872 );
    nor g2540 ( n1236 , n2729 , n1539 );
    or g2541 ( n2342 , n2869 , n2798 );
    xor g2542 ( n3411 , n1610 , n3143 );
    and g2543 ( n7 , n1409 , n2086 );
    and g2544 ( n1438 , n3638 , n1028 );
    xnor g2545 ( n2097 , n1608 , n3060 );
    not g2546 ( n1804 , n678 );
    or g2547 ( n493 , n1631 , n453 );
    and g2548 ( n2844 , n3684 , n3683 );
    or g2549 ( n1169 , n1814 , n3290 );
    and g2550 ( n302 , n236 , n3669 );
    not g2551 ( n949 , n230 );
    or g2552 ( n2072 , n3293 , n1413 );
    xnor g2553 ( n722 , n3203 , n3221 );
    or g2554 ( n2634 , n1372 , n2671 );
    or g2555 ( n1575 , n204 , n3267 );
    or g2556 ( n709 , n1403 , n1522 );
    xnor g2557 ( n847 , n685 , n1795 );
    not g2558 ( n1038 , n574 );
    nor g2559 ( n3117 , n2149 , n1160 );
    and g2560 ( n1976 , n1693 , n853 );
    xnor g2561 ( n324 , n562 , n1424 );
    and g2562 ( n1790 , n506 , n2789 );
    or g2563 ( n3041 , n3068 , n1601 );
    and g2564 ( n685 , n1130 , n211 );
    and g2565 ( n1681 , n2931 , n33 );
    and g2566 ( n3398 , n1810 , n1041 );
    xnor g2567 ( n3004 , n3678 , n2916 );
    or g2568 ( n1241 , n2553 , n802 );
    or g2569 ( n1470 , n3412 , n1691 );
    or g2570 ( n1666 , n1542 , n630 );
    not g2571 ( n3217 , n1618 );
    or g2572 ( n580 , n2517 , n649 );
    or g2573 ( n1597 , n1466 , n157 );
    and g2574 ( n2297 , n1257 , n2292 );
    or g2575 ( n1325 , n832 , n3060 );
    not g2576 ( n2590 , n491 );
    not g2577 ( n849 , n1745 );
    and g2578 ( n339 , n1493 , n1828 );
    xnor g2579 ( n2898 , n1774 , n2485 );
    and g2580 ( n2818 , n64 , n3022 );
    or g2581 ( n963 , n356 , n833 );
    and g2582 ( n3071 , n2219 , n1674 );
    xnor g2583 ( n155 , n409 , n172 );
    xnor g2584 ( n1730 , n1516 , n351 );
    or g2585 ( n2476 , n3448 , n230 );
    or g2586 ( n727 , n3567 , n2784 );
    or g2587 ( n1574 , n566 , n430 );
    xnor g2588 ( n2736 , n2065 , n3388 );
    or g2589 ( n2414 , n1814 , n445 );
    xnor g2590 ( n947 , n688 , n1219 );
    xnor g2591 ( n2507 , n2555 , n959 );
    or g2592 ( n2127 , n1987 , n2873 );
    and g2593 ( n3395 , n2126 , n1746 );
    not g2594 ( n51 , n78 );
    xnor g2595 ( n576 , n1521 , n2859 );
    and g2596 ( n3099 , n3210 , n616 );
    and g2597 ( n3140 , n1566 , n1148 );
    or g2598 ( n1427 , n2511 , n86 );
    xnor g2599 ( n2974 , n491 , n109 );
    and g2600 ( n2143 , n735 , n32 );
    not g2601 ( n3424 , n3492 );
    xnor g2602 ( n2281 , n1089 , n516 );
    nor g2603 ( n671 , n2811 , n3636 );
    xnor g2604 ( n390 , n103 , n2382 );
    or g2605 ( n2148 , n3309 , n44 );
    nor g2606 ( n1852 , n1089 , n2702 );
    or g2607 ( n1481 , n466 , n645 );
    not g2608 ( n1140 , n3333 );
    or g2609 ( n3262 , n2585 , n2917 );
    and g2610 ( n812 , n688 , n313 );
    nor g2611 ( n2359 , n2851 , n949 );
    or g2612 ( n2988 , n1880 , n3274 );
    or g2613 ( n1365 , n2570 , n1977 );
    and g2614 ( n2756 , n2230 , n11 );
    nor g2615 ( n408 , n2773 , n301 );
    xnor g2616 ( n786 , n3599 , n2641 );
    or g2617 ( n3519 , n1733 , n3371 );
    not g2618 ( n3248 , n2536 );
    not g2619 ( n3560 , n3024 );
    or g2620 ( n2368 , n621 , n1029 );
    xnor g2621 ( n932 , n809 , n1585 );
    or g2622 ( n2508 , n1307 , n1987 );
    nor g2623 ( n3118 , n1428 , n2943 );
    nor g2624 ( n3314 , n2145 , n348 );
    or g2625 ( n303 , n2864 , n2718 );
    and g2626 ( n2743 , n1943 , n890 );
    nor g2627 ( n1736 , n885 , n3161 );
    xnor g2628 ( n1062 , n2068 , n539 );
    and g2629 ( n2183 , n483 , n1076 );
    or g2630 ( n3168 , n1697 , n1997 );
    nor g2631 ( n3268 , n1484 , n448 );
    xnor g2632 ( n1569 , n2825 , n781 );
    and g2633 ( n2500 , n3519 , n1176 );
    or g2634 ( n1045 , n1871 , n1802 );
    and g2635 ( n647 , n746 , n1094 );
    or g2636 ( n3429 , n2871 , n354 );
    or g2637 ( n566 , n2648 , n445 );
    and g2638 ( n2488 , n1531 , n2205 );
    and g2639 ( n1475 , n1622 , n1521 );
    or g2640 ( n3197 , n1887 , n1573 );
    or g2641 ( n872 , n1140 , n2814 );
    or g2642 ( n746 , n1010 , n477 );
    or g2643 ( n409 , n2096 , n24 );
    and g2644 ( n1907 , n182 , n824 );
    nor g2645 ( n446 , n2491 , n2639 );
    and g2646 ( n806 , n2575 , n221 );
    xnor g2647 ( n1431 , n3146 , n1321 );
    and g2648 ( n1705 , n892 , n1047 );
    or g2649 ( n135 , n1973 , n1079 );
    xnor g2650 ( n1333 , n183 , n1875 );
    and g2651 ( n154 , n1332 , n697 );
    xnor g2652 ( n3350 , n256 , n2672 );
    not g2653 ( n568 , n2640 );
    and g2654 ( n2867 , n3261 , n3313 );
    or g2655 ( n3508 , n27 , n2830 );
    nor g2656 ( n1386 , n3600 , n3627 );
    nor g2657 ( n595 , n336 , n2736 );
    and g2658 ( n2850 , n3059 , n1492 );
    xnor g2659 ( n3061 , n733 , n1092 );
    and g2660 ( n3120 , n2660 , n1712 );
    and g2661 ( n945 , n367 , n3679 );
    or g2662 ( n2320 , n2009 , n2451 );
    and g2663 ( n1388 , n2682 , n3451 );
    and g2664 ( n3524 , n3011 , n2324 );
    not g2665 ( n3089 , n187 );
    not g2666 ( n2094 , n2253 );
    or g2667 ( n3655 , n1229 , n2228 );
    not g2668 ( n34 , n2853 );
    or g2669 ( n118 , n3546 , n379 );
    or g2670 ( n1656 , n1616 , n277 );
    or g2671 ( n1384 , n2648 , n1707 );
    and g2672 ( n1670 , n1411 , n3498 );
    not g2673 ( n3444 , n2055 );
    and g2674 ( n3422 , n3540 , n2034 );
    xnor g2675 ( n460 , n1828 , n2261 );
    nor g2676 ( n492 , n3633 , n1321 );
    or g2677 ( n164 , n2723 , n2897 );
    and g2678 ( n2189 , n3468 , n2006 );
    or g2679 ( n547 , n2220 , n3612 );
    xnor g2680 ( n596 , n2044 , n119 );
    and g2681 ( n203 , n458 , n1291 );
    or g2682 ( n3575 , n3397 , n571 );
    or g2683 ( n2478 , n1984 , n3480 );
    or g2684 ( n1395 , n2362 , n1509 );
    nor g2685 ( n477 , n2259 , n1003 );
    or g2686 ( n36 , n2246 , n39 );
    or g2687 ( n216 , n1428 , n3447 );
    or g2688 ( n2215 , n1380 , n3099 );
    and g2689 ( n934 , n1717 , n3605 );
    xnor g2690 ( n1737 , n3273 , n2433 );
    or g2691 ( n1206 , n3183 , n668 );
    xnor g2692 ( n3537 , n1723 , n1817 );
    and g2693 ( n1160 , n3259 , n2000 );
    or g2694 ( n1132 , n1987 , n902 );
    and g2695 ( n470 , n994 , n1835 );
    or g2696 ( n3680 , n2796 , n3620 );
    nor g2697 ( n2686 , n2547 , n644 );
    not g2698 ( n2313 , n3395 );
    xnor g2699 ( n2594 , n906 , n683 );
    and g2700 ( n2381 , n251 , n2720 );
    and g2701 ( n2855 , n2139 , n1013 );
    not g2702 ( n1809 , n1881 );
    xnor g2703 ( n172 , n2791 , n2867 );
    or g2704 ( n2575 , n5 , n250 );
    or g2705 ( n2555 , n457 , n3634 );
    xnor g2706 ( n2537 , n163 , n3573 );
    xnor g2707 ( n765 , n3668 , n2307 );
    or g2708 ( n1449 , n1146 , n397 );
    not g2709 ( n2126 , n1525 );
    and g2710 ( n96 , n2092 , n3491 );
    xnor g2711 ( n1064 , n2482 , n100 );
    not g2712 ( n3603 , n1159 );
    xnor g2713 ( n3457 , n1339 , n1322 );
    or g2714 ( n1032 , n652 , n3510 );
    xnor g2715 ( n396 , n3409 , n1698 );
    xnor g2716 ( n858 , n668 , n3453 );
    xnor g2717 ( n1837 , n2302 , n2401 );
    or g2718 ( n515 , n1596 , n1921 );
    and g2719 ( n1355 , n2414 , n2787 );
    xnor g2720 ( n1168 , n999 , n1046 );
    xnor g2721 ( n1391 , n1286 , n2594 );
    nor g2722 ( n637 , n891 , n3423 );
    and g2723 ( n2222 , n1411 , n476 );
    not g2724 ( n3049 , n891 );
    or g2725 ( n1401 , n1856 , n1 );
    or g2726 ( n3405 , n1310 , n1802 );
    or g2727 ( n3441 , n2809 , n1840 );
    and g2728 ( n2437 , n2742 , n3080 );
    not g2729 ( n1145 , n3353 );
    or g2730 ( n942 , n1898 , n3290 );
    and g2731 ( n590 , n601 , n558 );
    xnor g2732 ( n3412 , n3171 , n2548 );
    nor g2733 ( n2360 , n1344 , n2974 );
    xnor g2734 ( n1521 , n1029 , n3356 );
    and g2735 ( n1860 , n1091 , n837 );
    or g2736 ( n862 , n543 , n786 );
    not g2737 ( n2030 , n582 );
    and g2738 ( n2717 , n1368 , n2875 );
    or g2739 ( n1793 , n3174 , n3609 );
    or g2740 ( n3305 , n1161 , n1727 );
    and g2741 ( n612 , n1424 , n562 );
    xnor g2742 ( n2101 , n957 , n393 );
    or g2743 ( n2848 , n1898 , n1707 );
    not g2744 ( n3203 , n1972 );
    or g2745 ( n1248 , n3670 , n2941 );
    xnor g2746 ( n3402 , n3422 , n1713 );
    or g2747 ( n2808 , n2884 , n2289 );
    or g2748 ( n2781 , n452 , n2730 );
    or g2749 ( n3514 , n1540 , n1992 );
    and g2750 ( n5 , n3494 , n2058 );
    xnor g2751 ( n2416 , n2736 , n1955 );
    and g2752 ( n1339 , n406 , n3016 );
    xnor g2753 ( n2065 , n3289 , n1932 );
    and g2754 ( n2209 , n3094 , n2041 );
    xnor g2755 ( n2738 , n644 , n2547 );
    or g2756 ( n1302 , n2057 , n2556 );
    or g2757 ( n3334 , n2696 , n189 );
    and g2758 ( n2048 , n1011 , n1233 );
    nor g2759 ( n3249 , n1665 , n2873 );
    not g2760 ( n1324 , n460 );
    xnor g2761 ( n1007 , n2264 , n2170 );
    and g2762 ( n2474 , n2612 , n2067 );
    xnor g2763 ( n3344 , n2855 , n2439 );
    and g2764 ( n1066 , n493 , n913 );
    xnor g2765 ( n2998 , n1639 , n310 );
    or g2766 ( n337 , n345 , n1682 );
    xnor g2767 ( n101 , n1003 , n2259 );
    xnor g2768 ( n2428 , n907 , n597 );
    not g2769 ( n1353 , n589 );
    or g2770 ( n2804 , n441 , n1868 );
    xnor g2771 ( n3150 , n2993 , n3332 );
    xnor g2772 ( n1124 , n2473 , n22 );
    or g2773 ( n168 , n134 , n2339 );
    or g2774 ( n625 , n3202 , n1921 );
    and g2775 ( n805 , n3552 , n1504 );
    or g2776 ( n1872 , n90 , n3569 );
    xnor g2777 ( n2089 , n1799 , n1602 );
    xnor g2778 ( n3573 , n631 , n2744 );
    not g2779 ( n2661 , n1735 );
    xnor g2780 ( n76 , n1001 , n745 );
    or g2781 ( n2350 , n1871 , n2489 );
    or g2782 ( n2765 , n395 , n3070 );
    and g2783 ( n3315 , n1496 , n3596 );
    and g2784 ( n143 , n1473 , n2346 );
    xnor g2785 ( n147 , n3258 , n2235 );
    or g2786 ( n1971 , n1631 , n1658 );
    and g2787 ( n712 , n1751 , n640 );
    or g2788 ( n1826 , n2693 , n992 );
    xnor g2789 ( n2713 , n305 , n2778 );
    xnor g2790 ( n1410 , n699 , n2767 );
    or g2791 ( n2242 , n906 , n1286 );
    nor g2792 ( n2090 , n390 , n2496 );
    not g2793 ( n1573 , n59 );
    or g2794 ( n3253 , n1424 , n562 );
    xnor g2795 ( n957 , n153 , n3349 );
    or g2796 ( n423 , n2347 , n2189 );
    and g2797 ( n2701 , n785 , n3515 );
    xnor g2798 ( n1903 , n2570 , n431 );
    or g2799 ( n542 , n1567 , n2975 );
    or g2800 ( n1616 , n2030 , n329 );
    and g2801 ( n2866 , n1052 , n521 );
    and g2802 ( n832 , n722 , n1608 );
    and g2803 ( n379 , n2369 , n353 );
    xnor g2804 ( n2562 , n592 , n3405 );
    not g2805 ( n3516 , n885 );
    or g2806 ( n771 , n3011 , n2324 );
    or g2807 ( n698 , n2999 , n258 );
    and g2808 ( n711 , n3420 , n443 );
    or g2809 ( n614 , n3320 , n2856 );
    or g2810 ( n2390 , n696 , n1979 );
    xnor g2811 ( n3526 , n601 , n558 );
    and g2812 ( n1002 , n1463 , n978 );
    not g2813 ( n1310 , n400 );
    and g2814 ( n1437 , n3137 , n1758 );
    xnor g2815 ( n1036 , n3541 , n2669 );
    or g2816 ( n2484 , n1054 , n2753 );
    and g2817 ( n2001 , n2423 , n1645 );
    and g2818 ( n1327 , n1006 , n3083 );
    or g2819 ( n1011 , n925 , n2968 );
    or g2820 ( n2434 , n126 , n590 );
    xnor g2821 ( n2944 , n3064 , n1306 );
    xnor g2822 ( n687 , n2229 , n150 );
    xnor g2823 ( n440 , n3109 , n3224 );
    nor g2824 ( n2515 , n496 , n1164 );
    or g2825 ( n279 , n1023 , n2888 );
    and g2826 ( n2670 , n1944 , n103 );
    and g2827 ( n597 , n70 , n731 );
    xnor g2828 ( n1939 , n2597 , n1754 );
    not g2829 ( n2569 , n1970 );
    or g2830 ( n2395 , n3102 , n3079 );
    xnor g2831 ( n1593 , n444 , n993 );
    xor g2832 ( n1201 , n2856 , n49 );
    or g2833 ( n277 , n3293 , n1802 );
    xnor g2834 ( n2449 , n1048 , n300 );
    not g2835 ( n2397 , n1904 );
    not g2836 ( n995 , n3033 );
    or g2837 ( n856 , n1372 , n955 );
    or g2838 ( n1316 , n2569 , n3318 );
    or g2839 ( n1490 , n528 , n826 );
    or g2840 ( n2995 , n2553 , n1658 );
    or g2841 ( n1180 , n3479 , n2308 );
    not g2842 ( n2304 , n1327 );
    or g2843 ( n817 , n3248 , n1334 );
    and g2844 ( n2811 , n438 , n518 );
    and g2845 ( n1204 , n2466 , n1239 );
    and g2846 ( n387 , n2993 , n1624 );
    or g2847 ( n1874 , n1405 , n3318 );
    xnor g2848 ( n2722 , n325 , n684 );
    and g2849 ( n2950 , n965 , n3125 );
    or g2850 ( n1022 , n790 , n2867 );
    or g2851 ( n70 , n295 , n1959 );
    or g2852 ( n2053 , n897 , n2830 );
    or g2853 ( n1485 , n776 , n617 );
    or g2854 ( n2702 , n197 , n1847 );
    not g2855 ( n1540 , n794 );
    or g2856 ( n2195 , n3049 , n1385 );
    or g2857 ( n2699 , n2219 , n1674 );
    or g2858 ( n3300 , n2947 , n2435 );
    or g2859 ( n3126 , n3543 , n3205 );
    not g2860 ( n136 , n1561 );
    and g2861 ( n1260 , n1762 , n2085 );
    or g2862 ( n1396 , n788 , n118 );
    xnor g2863 ( n3427 , n2352 , n2187 );
    and g2864 ( n3469 , n3612 , n842 );
    or g2865 ( n2429 , n851 , n1413 );
    and g2866 ( n224 , n3324 , n2802 );
    xnor g2867 ( n2644 , n2929 , n2355 );
    not g2868 ( n1443 , n3035 );
    nor g2869 ( n1084 , n3043 , n2222 );
    xnor g2870 ( n3337 , n1200 , n1453 );
    xnor g2871 ( n646 , n1426 , n2705 );
    or g2872 ( n1652 , n813 , n2171 );
    xnor g2873 ( n2915 , n1399 , n2545 );
    and g2874 ( n2794 , n3198 , n2454 );
    or g2875 ( n2058 , n1268 , n2379 );
    not g2876 ( n3260 , n1954 );
    or g2877 ( n517 , n1814 , n1707 );
    and g2878 ( n196 , n1193 , n2905 );
    or g2879 ( n1807 , n2642 , n370 );
    and g2880 ( n1908 , n1967 , n1048 );
    and g2881 ( n3142 , n3536 , n3047 );
    and g2882 ( n2697 , n1481 , n2716 );
    or g2883 ( n2324 , n2921 , n1129 );
    not g2884 ( n2887 , n1426 );
    xnor g2885 ( n2170 , n3486 , n844 );
    and g2886 ( n2022 , n3588 , n464 );
    and g2887 ( n2406 , n629 , n2765 );
    xnor g2888 ( n1158 , n1491 , n2011 );
    xor g2889 ( n2248 , n625 , n2998 );
    not g2890 ( n3589 , n2019 );
    nor g2891 ( n2677 , n1713 , n1742 );
    and g2892 ( n836 , n2820 , n2843 );
    and g2893 ( n3631 , n3024 , n899 );
    and g2894 ( n2642 , n1638 , n3189 );
    or g2895 ( n167 , n128 , n1413 );
    and g2896 ( n377 , n2242 , n2392 );
    xnor g2897 ( n1789 , n1165 , n2426 );
    xnor g2898 ( n1214 , n1931 , n2276 );
    nor g2899 ( n1706 , n2163 , n2985 );
    or g2900 ( n1013 , n240 , n298 );
    xnor g2901 ( n535 , n1542 , n3244 );
    xnor g2902 ( n2813 , n2246 , n3681 );
    xnor g2903 ( n3547 , n2687 , n3128 );
    xnor g2904 ( n1416 , n2275 , n3342 );
    or g2905 ( n3399 , n2615 , n1138 );
    and g2906 ( n3500 , n1599 , n2413 );
    not g2907 ( n2190 , n2821 );
    or g2908 ( n2103 , n1358 , n1922 );
    xnor g2909 ( n2355 , n2452 , n3655 );
    or g2910 ( n3325 , n3594 , n2858 );
    or g2911 ( n1440 , n3417 , n445 );
    and g2912 ( n2650 , n1917 , n2497 );
    or g2913 ( n1240 , n851 , n554 );
    nor g2914 ( n3013 , n2220 , n1362 );
    or g2915 ( n939 , n1516 , n3456 );
    xnor g2916 ( n482 , n3473 , n1662 );
    not g2917 ( n842 , n1266 );
    or g2918 ( n3353 , n866 , n932 );
    and g2919 ( n1663 , n1505 , n2103 );
    or g2920 ( n2921 , n1921 , n1523 );
    or g2921 ( n1016 , n3433 , n152 );
    and g2922 ( n3387 , n579 , n3329 );
    or g2923 ( n1645 , n2255 , n2670 );
    or g2924 ( n351 , n2535 , n1802 );
    xnor g2925 ( n1450 , n1240 , n1487 );
    or g2926 ( n3380 , n3619 , n1910 );
    or g2927 ( n333 , n3260 , n461 );
    or g2928 ( n657 , n4 , n1950 );
    xnor g2929 ( n2581 , n2713 , n1588 );
    and g2930 ( n526 , n3331 , n266 );
    and g2931 ( n1986 , n1844 , n3307 );
    not g2932 ( n882 , n584 );
    and g2933 ( n448 , n2393 , n3328 );
    or g2934 ( n257 , n1428 , n438 );
    xnor g2935 ( n215 , n1674 , n3107 );
    and g2936 ( n1151 , n3027 , n1455 );
    or g2937 ( n2016 , n1882 , n809 );
    not g2938 ( n411 , n1352 );
    xnor g2939 ( n2334 , n1425 , n2028 );
    not g2940 ( n649 , n520 );
    not g2941 ( n946 , n2736 );
    and g2942 ( n2630 , n2002 , n1398 );
    and g2943 ( n3621 , n497 , n2494 );
    and g2944 ( n2752 , n2156 , n2327 );
    and g2945 ( n2980 , n2626 , n1517 );
    xnor g2946 ( n1162 , n515 , n3362 );
    or g2947 ( n2328 , n1288 , n428 );
    or g2948 ( n3209 , n3020 , n3226 );
    xnor g2949 ( n539 , n1448 , n2152 );
    xnor g2950 ( n464 , n1719 , n686 );
    xnor g2951 ( n3388 , n448 , n1484 );
    xnor g2952 ( n1453 , n2794 , n3484 );
    or g2953 ( n720 , n985 , n3386 );
    not g2954 ( n3275 , n730 );
    xnor g2955 ( n2667 , n1961 , n90 );
    or g2956 ( n206 , n2291 , n2664 );
    or g2957 ( n2862 , n3490 , n1541 );
    or g2958 ( n2388 , n2525 , n1178 );
    or g2959 ( n3067 , n3546 , n826 );
    and g2960 ( n766 , n958 , n2269 );
    or g2961 ( n2612 , n1851 , n1868 );
    xnor g2962 ( n1949 , n576 , n1626 );
    not g2963 ( n1962 , n2001 );
    not g2964 ( n2854 , n1641 );
    nor g2965 ( n2237 , n3554 , n2191 );
    xnor g2966 ( n650 , n1646 , n725 );
    xnor g2967 ( n983 , n985 , n3090 );
    or g2968 ( n3543 , n1540 , n1015 );
    or g2969 ( n2128 , n1150 , n3135 );
    xnor g2970 ( n1818 , n3075 , n3364 );
    and g2971 ( n1371 , n703 , n1181 );
    xnor g2972 ( n3442 , n1708 , n3065 );
    and g2973 ( n1077 , n1240 , n2274 );
    xnor g2974 ( n3036 , n410 , n1112 );
    not g2975 ( n643 , n1336 );
    not g2976 ( n2777 , n907 );
    or g2977 ( n2531 , n2345 , n2183 );
    or g2978 ( n2271 , n925 , n802 );
    and g2979 ( n2347 , n321 , n1636 );
    and g2980 ( n146 , n1440 , n2425 );
    or g2981 ( n2769 , n457 , n220 );
    or g2982 ( n2407 , n437 , n3038 );
    and g2983 ( n2975 , n901 , n3650 );
    xnor g2984 ( n1053 , n1011 , n1233 );
    or g2985 ( n693 , n552 , n1724 );
    or g2986 ( n3477 , n393 , n1528 );
    and g2987 ( n263 , n3183 , n668 );
    and g2988 ( n1400 , n2062 , n1396 );
    or g2989 ( n1547 , n1307 , n1658 );
    or g2990 ( n148 , n3272 , n2074 );
    not g2991 ( n1373 , n3189 );
    and g2992 ( n461 , n1464 , n2200 );
    or g2993 ( n703 , n2075 , n2590 );
    xnor g2994 ( n2135 , n3206 , n2223 );
    xnor g2995 ( n2911 , n1733 , n2629 );
    or g2996 ( n308 , n2184 , n744 );
    not g2997 ( n128 , n402 );
    or g2998 ( n3313 , n1980 , n934 );
    xnor g2999 ( n1060 , n1912 , n3280 );
    and g3000 ( n2021 , n3476 , n291 );
    or g3001 ( n937 , n2615 , n1413 );
    and g3002 ( n3155 , n444 , n1312 );
    or g3003 ( n1576 , n1462 , n2176 );
    or g3004 ( n2682 , n707 , n450 );
    not g3005 ( n3615 , n1187 );
    xnor g3006 ( n1381 , n2817 , n2283 );
    xnor g3007 ( n2805 , n188 , n1709 );
    nor g3008 ( n3346 , n1978 , n1024 );
    not g3009 ( n3283 , n2100 );
    xnor g3010 ( n1994 , n3597 , n2876 );
    or g3011 ( n350 , n1073 , n2750 );
    xnor g3012 ( n238 , n3028 , n1618 );
    xnor g3013 ( n1929 , n755 , n270 );
    or g3014 ( n682 , n3401 , n3599 );
    or g3015 ( n1883 , n3255 , n1868 );
    or g3016 ( n917 , n206 , n2471 );
    or g3017 ( n1257 , n692 , n3592 );
    not g3018 ( n763 , n573 );
    or g3019 ( n275 , n1659 , n1444 );
    and g3020 ( n2557 , n305 , n883 );
    not g3021 ( n1930 , n3336 );
    not g3022 ( n3022 , n3299 );
    xnor g3023 ( n218 , n3263 , n2693 );
    not g3024 ( n2740 , n2992 );
    or g3025 ( n2213 , n1433 , n975 );
    and g3026 ( n536 , n309 , n3593 );
    and g3027 ( n2330 , n2525 , n1178 );
    xnor g3028 ( n2913 , n1427 , n2164 );
    xnor g3029 ( n1838 , n413 , n1249 );
    not g3030 ( n2553 , n1125 );
    or g3031 ( n1584 , n3417 , n3152 );
    xor g3032 ( n1030 , n1248 , n836 );
    xnor g3033 ( n1696 , n138 , n20 );
    or g3034 ( n2792 , n1107 , n1126 );
    and g3035 ( n3601 , n531 , n3678 );
    xnor g3036 ( n454 , n35 , n536 );
    or g3037 ( n3032 , n1661 , n3318 );
    or g3038 ( n3571 , n1699 , n739 );
    and g3039 ( n2251 , n3220 , n743 );
    or g3040 ( n2693 , n1372 , n1235 );
    and g3041 ( n3100 , n1951 , n3341 );
    or g3042 ( n86 , n2753 , n485 );
    or g3043 ( n3496 , n2096 , n802 );
    or g3044 ( n878 , n2220 , n2322 );
    or g3045 ( n2139 , n503 , n1139 );
    and g3046 ( n758 , n1131 , n796 );
    and g3047 ( n3348 , n3659 , n1766 );
    xnor g3048 ( n2125 , n1556 , n3426 );
    or g3049 ( n1821 , n1376 , n661 );
    and g3050 ( n1040 , n621 , n1029 );
    not g3051 ( n2436 , n2512 );
    and g3052 ( n2400 , n288 , n3499 );
    xnor g3053 ( n1520 , n791 , n0 );
    or g3054 ( n2545 , n1596 , n2671 );
    nor g3055 ( n1495 , n2607 , n1770 );
    or g3056 ( n3210 , n2338 , n3556 );
    or g3057 ( n3146 , n504 , n2677 );
    xnor g3058 ( n752 , n2837 , n847 );
    or g3059 ( n2326 , n2096 , n2294 );
    not g3060 ( n2296 , n2129 );
    and g3061 ( n810 , n2910 , n2190 );
    and g3062 ( n2282 , n1530 , n1510 );
    and g3063 ( n3365 , n2600 , n522 );
    or g3064 ( n1791 , n239 , n1132 );
    xnor g3065 ( n1932 , n3354 , n3582 );
    xnor g3066 ( n2680 , n1892 , n1748 );
    or g3067 ( n2977 , n3546 , n1989 );
    or g3068 ( n1895 , n3096 , n2712 );
    and g3069 ( n141 , n3511 , n3227 );
    or g3070 ( n21 , n3312 , n976 );
    or g3071 ( n3311 , n1685 , n2111 );
    or g3072 ( n2655 , n1987 , n2340 );
    xnor g3073 ( n2482 , n1753 , n1800 );
    not g3074 ( n3612 , n1825 );
    or g3075 ( n3632 , n3319 , n670 );
    xnor g3076 ( n967 , n415 , n1595 );
    xnor g3077 ( n665 , n2032 , n10 );
    or g3078 ( n2440 , n3046 , n1197 );
    nor g3079 ( n2045 , n669 , n2827 );
    and g3080 ( n1963 , n2580 , n1238 );
    xnor g3081 ( n3306 , n2279 , n981 );
    nor g3082 ( n3287 , n3333 , n3578 );
    or g3083 ( n2924 , n898 , n3534 );
    not g3084 ( n2564 , n2300 );
    and g3085 ( n900 , n844 , n2264 );
    or g3086 ( n2154 , n1151 , n3548 );
    xnor g3087 ( n2720 , n2869 , n2258 );
    and g3088 ( n2812 , n543 , n786 );
    or g3089 ( n513 , n2946 , n2074 );
    xnor g3090 ( n1954 , n3309 , n1629 );
    not g3091 ( n1402 , n1421 );
    and g3092 ( n715 , n2836 , n3300 );
    xnor g3093 ( n1082 , n2058 , n250 );
    or g3094 ( n3593 , n3240 , n3406 );
    xnor g3095 ( n2152 , n3635 , n3545 );
    or g3096 ( n1958 , n173 , n955 );
    and g3097 ( n584 , n15 , n2632 );
    not g3098 ( n3152 , n2311 );
    or g3099 ( n2510 , n2648 , n3290 );
    xnor g3100 ( n3408 , n2457 , n1044 );
    or g3101 ( n3230 , n1386 , n1577 );
    or g3102 ( n998 , n1307 , n2968 );
    or g3103 ( n50 , n87 , n2268 );
    nor g3104 ( n773 , n769 , n984 );
    or g3105 ( n2774 , n1874 , n3572 );
    not g3106 ( n24 , n2666 );
    and g3107 ( n2652 , n2499 , n2211 );
    or g3108 ( n1492 , n1323 , n1845 );
    or g3109 ( n1444 , n3255 , n1243 );
    and g3110 ( n807 , n864 , n2138 );
    and g3111 ( n2873 , n3134 , n1422 );
    xnor g3112 ( n1823 , n32 , n1021 );
    or g3113 ( n1174 , n1596 , n34 );
    or g3114 ( n688 , n446 , n17 );
    or g3115 ( n1380 , n1192 , n867 );
    or g3116 ( n608 , n1898 , n2830 );
    and g3117 ( n3582 , n293 , n783 );
    and g3118 ( n1993 , n1143 , n1490 );
    or g3119 ( n267 , n1172 , n3470 );
    and g3120 ( n2518 , n772 , n1551 );
    xnor g3121 ( n84 , n2611 , n2446 );
    and g3122 ( n2049 , n872 , n414 );
    or g3123 ( n3263 , n3202 , n2712 );
    xnor g3124 ( n2685 , n1680 , n1940 );
    and g3125 ( n910 , n95 , n2093 );
    and g3126 ( n2331 , n3245 , n66 );
    not g3127 ( n1552 , n2301 );
    and g3128 ( n417 , n1833 , n3105 );
    nor g3129 ( n3653 , n3546 , n815 );
    or g3130 ( n1513 , n416 , n1009 );
    and g3131 ( n3480 , n3106 , n2832 );
    and g3132 ( n562 , n2852 , n2981 );
    xnor g3133 ( n2714 , n1060 , n1232 );
    or g3134 ( n3678 , n429 , n1442 );
    not g3135 ( n2519 , n3445 );
    and g3136 ( n1056 , n1069 , n2279 );
    not g3137 ( n1869 , n1214 );
    and g3138 ( n1567 , n3436 , n2679 );
    and g3139 ( n1690 , n473 , n2196 );
    and g3140 ( n2490 , n906 , n1286 );
    not g3141 ( n1347 , n202 );
    xnor g3142 ( n663 , n3375 , n2805 );
    and g3143 ( n209 , n124 , n1536 );
    not g3144 ( n2265 , n3381 );
    and g3145 ( n2770 , n2009 , n2451 );
    or g3146 ( n2874 , n601 , n558 );
    or g3147 ( n1429 , n3418 , n1554 );
    or g3148 ( n1561 , n1310 , n2489 );
    and g3149 ( n2935 , n219 , n2880 );
    and g3150 ( n1983 , n3500 , n3252 );
    or g3151 ( n1239 , n2487 , n3058 );
    xnor g3152 ( n187 , n1651 , n3292 );
    and g3153 ( n1632 , n2403 , n3497 );
    or g3154 ( n2959 , n3588 , n464 );
    or g3155 ( n2663 , n263 , n2224 );
    and g3156 ( n557 , n930 , n564 );
    not g3157 ( n2198 , n1130 );
    xnor g3158 ( n1112 , n910 , n2193 );
    and g3159 ( n1743 , n3419 , n2052 );
    or g3160 ( n3010 , n305 , n883 );
    and g3161 ( n3495 , n3645 , n1728 );
    and g3162 ( n1792 , n2380 , n2559 );
    and g3163 ( n282 , n1417 , n2565 );
    and g3164 ( n3507 , n1190 , n2440 );
    or g3165 ( n365 , n2510 , n1890 );
    or g3166 ( n1659 , n2362 , n1334 );
    or g3167 ( n839 , n581 , n18 );
    or g3168 ( n3110 , n673 , n3180 );
    or g3169 ( n1728 , n897 , n445 );
    and g3170 ( n2060 , n2793 , n2453 );
    or g3171 ( n960 , n1397 , n1598 );
    and g3172 ( n1278 , n1516 , n3456 );
    or g3173 ( n1035 , n2280 , n2385 );
    or g3174 ( n3176 , n2031 , n2727 );
    not g3175 ( n1814 , n3238 );
    or g3176 ( n2460 , n1405 , n220 );
    xnor g3177 ( n2401 , n350 , n715 );
    or g3178 ( n1283 , n2220 , n1154 );
    nor g3179 ( n1697 , n297 , n3144 );
    or g3180 ( n3072 , n2615 , n554 );
    xnor g3181 ( n508 , n2364 , n602 );
    and g3182 ( n2858 , n129 , n2794 );
    xnor g3183 ( n3001 , n1671 , n245 );
    and g3184 ( n467 , n2140 , n1157 );
    or g3185 ( n3476 , n839 , n1786 );
    xnor g3186 ( n3121 , n412 , n3590 );
    and g3187 ( n3488 , n355 , n1734 );
    and g3188 ( n1137 , n771 , n3481 );
    or g3189 ( n3578 , n2762 , n3348 );
    or g3190 ( n1710 , n3326 , n2294 );
    not g3191 ( n2305 , n3568 );
    and g3192 ( n1769 , n1923 , n546 );
    not g3193 ( n380 , n610 );
    xnor g3194 ( n2778 , n883 , n107 );
    or g3195 ( n1722 , n3021 , n1761 );
    or g3196 ( n690 , n1540 , n445 );
    not g3197 ( n1463 , n1169 );
    or g3198 ( n948 , n2064 , n3365 );
    or g3199 ( n3057 , n2649 , n1415 );
    or g3200 ( n936 , n2542 , n2441 );
    and g3201 ( n111 , n410 , n620 );
    or g3202 ( n2205 , n2446 , n1063 );
    xor g3203 ( n353 , n2533 , n679 );
    xnor g3204 ( n695 , n2757 , n1747 );
    xnor g3205 ( n1990 , n2092 , n3491 );
    and g3206 ( n2149 , n2877 , n1557 );
    xnor g3207 ( n2711 , n919 , n2212 );
    xnor g3208 ( n1484 , n241 , n2561 );
    and g3209 ( n1752 , n322 , n2395 );
    xnor g3210 ( n3113 , n559 , n2788 );
    xnor g3211 ( n62 , n1942 , n2911 );
    or g3212 ( n710 , n2949 , n1088 );
    not g3213 ( n1631 , n2310 );
    not g3214 ( n1334 , n388 );
    or g3215 ( n1009 , n2163 , n3023 );
    or g3216 ( n1096 , n1102 , n1083 );
    xnor g3217 ( n1306 , n2932 , n371 );
    or g3218 ( n1340 , n3472 , n1936 );
    or g3219 ( n3193 , n3248 , n2074 );
    not g3220 ( n97 , n2797 );
    not g3221 ( n453 , n1087 );
    nor g3222 ( n2509 , n1496 , n3596 );
    xnor g3223 ( n1021 , n735 , n83 );
    xnor g3224 ( n3332 , n1226 , n1053 );
    or g3225 ( n221 , n3494 , n2058 );
    or g3226 ( n3407 , n2630 , n2110 );
    not g3227 ( n2645 , n711 );
    xnor g3228 ( n795 , n3190 , n1838 );
    not g3229 ( n44 , n1629 );
    and g3230 ( n3103 , n3122 , n3574 );
    and g3231 ( n543 , n2128 , n1394 );
    xnor g3232 ( n1122 , n3507 , n3201 );
    or g3233 ( n556 , n3277 , n576 );
    or g3234 ( n2084 , n1814 , n649 );
    xnor g3235 ( n394 , n3180 , n673 );
    or g3236 ( n1256 , n1887 , n2010 );
    and g3237 ( n2176 , n494 , n1945 );
    xnor g3238 ( n1109 , n2326 , n207 );
    not g3239 ( n2000 , n63 );
    or g3240 ( n1083 , n2753 , n46 );
    and g3241 ( n1326 , n290 , n2839 );
    xnor g3242 ( n1199 , n817 , n2488 );
    or g3243 ( n401 , n3550 , n189 );
    and g3244 ( n2231 , n2680 , n2129 );
    xnor g3245 ( n376 , n3091 , n332 );
    nor g3246 ( n1526 , n2713 , n2051 );
    or g3247 ( n2280 , n2362 , n1243 );
    xnor g3248 ( n741 , n2598 , n1256 );
    xnor g3249 ( n3604 , n1178 , n1432 );
    or g3250 ( n2905 , n823 , n914 );
    xor g3251 ( n987 , n1253 , n2338 );
    or g3252 ( n3642 , n3546 , n1993 );
    or g3253 ( n3075 , n3615 , n2074 );
    xnor g3254 ( n43 , n937 , n1483 );
    or g3255 ( n1627 , n3301 , n577 );
    or g3256 ( n2228 , n3546 , n137 );
    or g3257 ( n2729 , n1814 , n2830 );
    xnor g3258 ( n1505 , n1118 , n2996 );
    and g3259 ( n1297 , n3446 , n2963 );
    or g3260 ( n1341 , n1093 , n3030 );
    xnor g3261 ( n2394 , n1333 , n3179 );
    or g3262 ( n1734 , n664 , n1400 );
    xnor g3263 ( n852 , n3227 , n3511 );
    or g3264 ( n2784 , n851 , n1138 );
    not g3265 ( n2233 , n3366 );
    and g3266 ( n1764 , n3463 , n3305 );
    and g3267 ( n560 , n2221 , n1316 );
    or g3268 ( n2262 , n3197 , n642 );
    or g3269 ( n165 , n492 , n2912 );
    xnor g3270 ( n3087 , n3665 , n3454 );
    or g3271 ( n2256 , n2930 , n1012 );
    not g3272 ( n2489 , n3566 );
    and g3273 ( n87 , n267 , n2147 );
    not g3274 ( n3403 , n2628 );
    or g3275 ( n749 , n971 , n822 );
    and g3276 ( n1691 , n877 , n2218 );
    not g3277 ( n627 , n1579 );
    or g3278 ( n2086 , n1297 , n1333 );
    and g3279 ( n2372 , n1252 , n3026 );
    not g3280 ( n1320 , n1001 );
    xnor g3281 ( n509 , n2267 , n2692 );
    or g3282 ( n1309 , n2362 , n2074 );
    nor g3283 ( n1859 , n3074 , n693 );
    and g3284 ( n759 , n2649 , n1415 );
    or g3285 ( n1654 , n1566 , n1148 );
    and g3286 ( n438 , n3560 , n830 );
    not g3287 ( n1684 , n2493 );
    and g3288 ( n3641 , n3174 , n3609 );
    or g3289 ( n405 , n1215 , n3187 );
    and g3290 ( n1829 , n2396 , n2758 );
    or g3291 ( n594 , n3546 , n436 );
    xnor g3292 ( n2019 , n3677 , n611 );
    or g3293 ( n2732 , n817 , n2277 );
    or g3294 ( n2037 , n1596 , n189 );
    or g3295 ( n2337 , n1578 , n2837 );
    and g3296 ( n702 , n3554 , n2191 );
    or g3297 ( n2558 , n1540 , n2830 );
    and g3298 ( n334 , n2144 , n1813 );
    xnor g3299 ( n3565 , n2038 , n2865 );
    or g3300 ( n3401 , n3293 , n554 );
    and g3301 ( n1111 , n379 , n3411 );
    and g3302 ( n2731 , n3032 , n1671 );
    and g3303 ( n2137 , n2613 , n1837 );
    xnor g3304 ( n2095 , n3003 , n1317 );
    or g3305 ( n2698 , n458 , n1291 );
    xor g3306 ( n770 , n226 , n2522 );
    or g3307 ( n3007 , n550 , n2467 );
    or g3308 ( n468 , n2050 , n1057 );
    and g3309 ( n952 , n2738 , n584 );
    xnor g3310 ( n179 , n1210 , n2621 );
    not g3311 ( n268 , n1638 );
    or g3312 ( n2185 , n2439 , n968 );
    or g3313 ( n2914 , n3665 , n1224 );
    not g3314 ( n2615 , n228 );
    and g3315 ( n2922 , n2868 , n3069 );
    xnor g3316 ( n2635 , n3279 , n482 );
    and g3317 ( n2062 , n2587 , n292 );
    or g3318 ( n1536 , n3158 , n2668 );
    or g3319 ( n1542 , n1887 , n2397 );
    and g3320 ( n1996 , n323 , n2210 );
    or g3321 ( n289 , n3201 , n3507 );
    not g3322 ( n3267 , n2387 );
    nor g3323 ( n788 , n2369 , n353 );
    xnor g3324 ( n3000 , n2415 , n72 );
    or g3325 ( n2860 , n2122 , n2770 );
    or g3326 ( n60 , n3119 , n1564 );
    or g3327 ( n2465 , n581 , n2712 );
    xnor g3328 ( n1735 , n1837 , n1796 );
    or g3329 ( n1148 , n1898 , n3152 );
    or g3330 ( n841 , n612 , n1812 );
    or g3331 ( n1299 , n2092 , n3491 );
    or g3332 ( n1245 , n3546 , n1811 );
    or g3333 ( n2315 , n1851 , n1243 );
    or g3334 ( n81 , n1136 , n1651 );
    or g3335 ( n2003 , n375 , n1186 );
    or g3336 ( n565 , n3389 , n3504 );
    xnor g3337 ( n3594 , n231 , n3502 );
    nor g3338 ( n29 , n1353 , n2416 );
    not g3339 ( n3550 , n3542 );
    or g3340 ( n1647 , n1795 , n2013 );
    and g3341 ( n1537 , n2698 , n1247 );
    not g3342 ( n1253 , n3374 );
    and g3343 ( n3416 , n1846 , n1071 );
    xnor g3344 ( n1560 , n3408 , n2437 );
    and g3345 ( n3644 , n1983 , n1201 );
    xnor g3346 ( n3602 , n2001 , n2779 );
    or g3347 ( n2046 , n3539 , n2250 );
    not g3348 ( n3247 , n593 );
    and g3349 ( n1085 , n2480 , n3496 );
    xnor g3350 ( n274 , n2921 , n3219 );
    or g3351 ( n731 , n861 , n8 );
    or g3352 ( n2253 , n2030 , n2233 );
    nor g3353 ( n2432 , n1794 , n3113 );
    xnor g3354 ( n1149 , n1569 , n3427 );
    and g3355 ( n3178 , n1969 , n1652 );
    xnor g3356 ( n2795 , n2897 , n3154 );
    or g3357 ( n1768 , n2580 , n1238 );
    or g3358 ( n115 , n3155 , n1416 );
    or g3359 ( n1274 , n1684 , n1423 );
    not g3360 ( n3139 , n3487 );
    not g3361 ( n2424 , n3100 );
    or g3362 ( n1566 , n3417 , n3290 );
    xnor g3363 ( n1624 , n3496 , n1935 );
    or g3364 ( n57 , n40 , n933 );
    or g3365 ( n130 , n255 , n2714 );
    and g3366 ( n2325 , n1919 , n1281 );
    nor g3367 ( n424 , n3335 , n2788 );
    or g3368 ( n2151 , n3178 , n3520 );
    or g3369 ( n2880 , n2819 , n220 );
    and g3370 ( n1300 , n860 , n1867 );
    and g3371 ( n2709 , n268 , n1373 );
    and g3372 ( n419 , n1853 , n3501 );
    xnor g3373 ( n1322 , n2595 , n1359 );
    xnor g3374 ( n2718 , n1988 , n967 );
    xnor g3375 ( n2856 , n2442 , n199 );
    and g3376 ( n2799 , n2046 , n3531 );
    and g3377 ( n668 , n1032 , n2172 );
    and g3378 ( n3517 , n723 , n3489 );
    or g3379 ( n1680 , n441 , n1509 );
    xnor g3380 ( n1519 , n1999 , n3471 );
    and g3381 ( n3130 , n1059 , n882 );
    or g3382 ( n1254 , n1469 , n3306 );
    and g3383 ( n315 , n164 , n3637 );
    not g3384 ( n918 , n2882 );
    not g3385 ( n2658 , n1815 );
    xnor g3386 ( n1538 , n2649 , n1877 );
    or g3387 ( n1360 , n374 , n2066 );
    or g3388 ( n2479 , n415 , n1988 );
    not g3389 ( n1661 , n3156 );
    or g3390 ( n2144 , n3075 , n3364 );
    xnor g3391 ( n658 , n593 , n2095 );
    not g3392 ( n392 , n62 );
    and g3393 ( n895 , n3640 , n2117 );
    and g3394 ( n2272 , n791 , n71 );
    xnor g3395 ( n1708 , n3001 , n2285 );
    and g3396 ( n202 , n1625 , n1258 );
    or g3397 ( n523 , n2597 , n1296 );
    xnor g3398 ( n2283 , n1649 , n40 );
    or g3399 ( n2329 , n3326 , n2750 );
    xnor g3400 ( n1155 , n481 , n2183 );
    or g3401 ( n3617 , n2783 , n1637 );
    and g3402 ( n1448 , n974 , n991 );
    or g3403 ( n2817 , n53 , n220 );
    xnor g3404 ( n3426 , n3131 , n3367 );
    or g3405 ( n3456 , n487 , n2233 );
    nor g3406 ( n3595 , n935 , n943 );
    or g3407 ( n3490 , n457 , n2010 );
    or g3408 ( n510 , n1474 , n2922 );
    or g3409 ( n3231 , n2061 , n1045 );
    xnor g3410 ( n1800 , n1974 , n1635 );
    not g3411 ( n1599 , n2380 );
    xnor g3412 ( n613 , n3645 , n580 );
    xnor g3413 ( n2192 , n3459 , n760 );
    and g3414 ( n2433 , n666 , n2018 );
    xnor g3415 ( n1719 , n227 , n3611 );
    xnor g3416 ( n3088 , n1884 , n3398 );
    not g3417 ( n1405 , n3529 );
    xnor g3418 ( n104 , n2809 , n1840 );
    not g3419 ( n1170 , n2521 );
    and g3420 ( n413 , n3050 , n2342 );
    and g3421 ( n285 , n1027 , n3622 );
    or g3422 ( n162 , n3471 , n2605 );
    and g3423 ( n1197 , n1607 , n2813 );
    and g3424 ( n249 , n682 , n2363 );
    xnor g3425 ( n2258 , n1824 , n2037 );
    xnor g3426 ( n2767 , n342 , n91 );
    and g3427 ( n489 , n3095 , n1420 );
    or g3428 ( n2499 , n637 , n1369 );
    not g3429 ( n897 , n1367 );
    or g3430 ( n2138 , n1384 , n750 );
    or g3431 ( n1590 , n2386 , n2987 );
    not g3432 ( n1108 , n2433 );
    and g3433 ( n1724 , n921 , n3148 );
    or g3434 ( n1356 , n2966 , n1807 );
    or g3435 ( n3343 , n3417 , n2830 );
    or g3436 ( n1767 , n2945 , n286 );
    xnor g3437 ( n3227 , n3552 , n122 );
    and g3438 ( n3465 , n3551 , n1359 );
    xnor g3439 ( n1638 , n1598 , n1397 );
    nor g3440 ( n3522 , n1143 , n1490 );
    xnor g3441 ( n1227 , n1572 , n1174 );
    or g3442 ( n259 , n3522 , n3642 );
    not g3443 ( n254 , n333 );
    and g3444 ( n661 , n3632 , n1740 );
    or g3445 ( n3261 , n1717 , n3605 );
    not g3446 ( n1894 , n3523 );
    or g3447 ( n2662 , n481 , n1696 );
    or g3448 ( n1418 , n3466 , n1162 );
    or g3449 ( n778 , n2763 , n2579 );
    and g3450 ( n3475 , n3665 , n1224 );
    xnor g3451 ( n1106 , n1024 , n2281 );
    xnor g3452 ( n2035 , n838 , n419 );
    and g3453 ( n1528 , n957 , n1314 );
    xnor g3454 ( n28 , n104 , n2711 );
    nor g3455 ( n2504 , n1213 , n909 );
    or g3456 ( n1787 , n2030 , n1802 );
    and g3457 ( n3368 , n3623 , n3505 );
    and g3458 ( n2572 , n2835 , n2326 );
    and g3459 ( n2827 , n1187 , n2516 );
    and g3460 ( n885 , n1676 , n1117 );
    or g3461 ( n3136 , n1058 , n341 );
    xnor g3462 ( n2657 , n1342 , n1276 );
    or g3463 ( n3541 , n2420 , n1614 );
    or g3464 ( n2180 , n3258 , n1791 );
    and g3465 ( n808 , n335 , n3206 );
    xnor g3466 ( n2298 , n2991 , n2695 );
    xnor g3467 ( n3235 , n1028 , n758 );
    and g3468 ( n3569 , n633 , n1961 );
    or g3469 ( n1500 , n265 , n260 );
    and g3470 ( n2100 , n1590 , n2180 );
    nor g3471 ( n1589 , n1100 , n3396 );
    and g3472 ( n225 , n592 , n3405 );
    not g3473 ( n1888 , n2224 );
    not g3474 ( n1596 , n3034 );
    xnor g3475 ( n3676 , n529 , n253 );
    not g3476 ( n2010 , n74 );
    xnor g3477 ( n2803 , n2422 , n334 );
    or g3478 ( n2425 , n1898 , n1992 );
    not g3479 ( n2872 , n3387 );
    and g3480 ( n1121 , n3387 , n1511 );
    or g3481 ( n879 , n2091 , n529 );
    or g3482 ( n3620 , n3255 , n1648 );
    or g3483 ( n3373 , n539 , n886 );
    and g3484 ( n1635 , n1234 , n2690 );
    xnor g3485 ( n3484 , n129 , n3594 );
    and g3486 ( n451 , n2366 , n112 );
    xnor g3487 ( n1048 , n1329 , n1998 );
    or g3488 ( n1233 , n1073 , n24 );
    and g3489 ( n2389 , n1230 , n1780 );
    and g3490 ( n2115 , n1833 , n3366 );
    and g3491 ( n2607 , n3043 , n2222 );
    nor g3492 ( n2833 , n2177 , n3582 );
    xnor g3493 ( n300 , n1967 , n1217 );
    not g3494 ( n1216 , n1484 );
    and g3495 ( n78 , n1558 , n3089 );
    xnor g3496 ( n1891 , n719 , n1303 );
    not g3497 ( n2057 , n116 );
    xnor g3498 ( n3614 , n696 , n1979 );
    and g3499 ( n3166 , n3081 , n2925 );
    xnor g3500 ( n428 , n3286 , n218 );
    xnor g3501 ( n1378 , n2429 , n2922 );
    or g3502 ( n1862 , n2001 , n3391 );
    or g3503 ( n346 , n1210 , n3200 );
    xnor g3504 ( n2962 , n2054 , n359 );
    xnor g3505 ( n1535 , n1513 , n1861 );
    not g3506 ( n955 , n1905 );
    or g3507 ( n1190 , n1607 , n2813 );
    xnor g3508 ( n2982 , n3479 , n2243 );
    or g3509 ( n1176 , n110 , n1942 );
    and g3510 ( n1741 , n3201 , n3507 );
    and g3511 ( n1981 , n2706 , n2206 );
    not g3512 ( n149 , n448 );
    nor g3513 ( n2800 , n911 , n2083 );
    or g3514 ( n2841 , n3029 , n3676 );
    and g3515 ( n3058 , n183 , n1410 );
    nor g3516 ( n1586 , n2500 , n845 );
    and g3517 ( n2608 , n1248 , n306 );
    and g3518 ( n2831 , n1311 , n709 );
    or g3519 ( n120 , n536 , n343 );
    or g3520 ( n3240 , n925 , n2294 );
    xnor g3521 ( n1078 , n2714 , n255 );
    nor g3522 ( n3389 , n3500 , n3252 );
    and g3523 ( n2759 , n402 , n653 );
    and g3524 ( n1646 , n1467 , n980 );
    and g3525 ( n1725 , n1086 , n1606 );
    xnor g3526 ( n1406 , n1735 , n3056 );
    or g3527 ( n1726 , n2831 , n212 );
    or g3528 ( n1847 , n2753 , n1583 );
    nor g3529 ( n2438 , n408 , n2943 );
    or g3530 ( n194 , n3293 , n329 );
    or g3531 ( n2116 , n2678 , n1976 );
    or g3532 ( n2953 , n22 , n2473 );
    or g3533 ( n3294 , n2592 , n1020 );
    or g3534 ( n261 , n1255 , n3492 );
    and g3535 ( n1424 , n2703 , n1035 );
    or g3536 ( n555 , n204 , n453 );
    and g3537 ( n3450 , n3195 , n889 );
    or g3538 ( n1803 , n1871 , n2186 );
    or g3539 ( n494 , n994 , n1835 );
    or g3540 ( n1644 , n2753 , n801 );
    not g3541 ( n1871 , n1833 );
    or g3542 ( n2085 , n2551 , n2907 );
    and g3543 ( n609 , n1399 , n1277 );
    or g3544 ( n2123 , n2414 , n2787 );
    or g3545 ( n2593 , n688 , n313 );
    or g3546 ( n1878 , n1738 , n1245 );
    or g3547 ( n1571 , n83 , n2143 );
    or g3548 ( n1497 , n2753 , n3603 );
    or g3549 ( n1531 , n2611 , n2252 );
    or g3550 ( n1835 , n2096 , n2750 );
    nor g3551 ( n170 , n1001 , n372 );
    or g3552 ( n3214 , n2753 , n3358 );
    xnor g3553 ( n3502 , n2008 , n2807 );
    xnor g3554 ( n3289 , n2210 , n1203 );
    and g3555 ( n1754 , n303 , n710 );
    and g3556 ( n3299 , n3662 , n1055 );
    or g3557 ( n2122 , n457 , n1573 );
    nor g3558 ( n110 , n2024 , n2629 );
    or g3559 ( n397 , n1809 , n754 );
    not g3560 ( n3202 , n1123 );
    or g3561 ( n186 , n2459 , n1906 );
    and g3562 ( n152 , n868 , n604 );
    and g3563 ( n422 , n2945 , n286 );
endmodule
