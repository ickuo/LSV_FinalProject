module top( n1 , n3 , n10 , n15 , n18 , n20 , n29 , n31 , n33 , 
n42 , n43 , n49 , n52 , n69 , n71 , n73 , n75 , n76 , n91 , 
n96 , n101 , n103 , n107 , n112 , n114 , n116 , n117 , n133 , n135 , 
n139 , n149 , n152 , n164 , n165 , n180 , n197 , n200 , n219 , n226 , 
n227 , n228 , n233 , n235 , n256 , n257 , n263 , n282 , n284 , n285 , 
n292 , n293 , n297 , n303 , n313 , n321 , n325 , n326 , n330 , n334 , 
n336 , n337 , n351 , n359 , n373 , n379 , n398 , n399 , n409 , n413 , 
n422 , n434 , n438 , n446 , n459 , n462 , n463 , n473 , n477 , n484 , 
n492 , n498 , n503 , n507 , n516 , n519 , n524 , n526 , n531 , n555 , 
n559 , n575 , n580 , n582 , n587 , n601 , n604 , n617 , n636 , n644 , 
n647 , n652 , n675 , n676 , n680 , n687 , n691 , n703 , n705 , n709 , 
n710 , n712 , n718 , n720 , n749 , n751 , n754 , n757 , n762 , n770 , 
n774 , n775 , n784 , n785 , n789 , n796 , n803 , n805 , n810 , n812 , 
n818 , n834 , n838 , n842 , n854 , n858 , n863 , n873 , n877 , n886 , 
n889 , n895 , n897 , n912 , n915 , n924 , n926 , n928 , n932 , n941 , 
n945 , n949 , n953 , n954 , n958 , n960 , n963 , n966 , n971 , n974 , 
n983 , n984 , n986 , n991 , n1013 , n1015 , n1027 , n1049 , n1051 , n1061 , 
n1062 , n1063 , n1084 , n1086 , n1094 , n1105 , n1113 , n1114 , n1116 , n1122 , 
n1130 , n1136 , n1143 , n1144 , n1145 , n1150 , n1151 , n1161 , n1163 , n1178 , 
n1179 , n1201 , n1204 , n1216 , n1219 , n1229 , n1233 , n1235 , n1238 , n1241 , 
n1253 , n1260 , n1266 , n1268 , n1274 , n1276 , n1277 , n1287 , n1297 , n1301 , 
n1305 , n1309 , n1314 , n1328 , n1332 , n1338 , n1347 , n1352 , n1360 , n1366 , 
n1372 , n1392 , n1393 , n1395 , n1403 , n1405 , n1418 , n1428 , n1434 , n1458 , 
n1461 , n1470 , n1481 , n1491 , n1499 , n1503 , n1504 , n1506 , n1514 , n1533 , 
n1544 , n1548 , n1549 , n1558 , n1559 , n1576 , n1583 , n1585 , n1615 , n1616 , 
n1625 , n1629 , n1631 , n1632 , n1648 , n1660 , n1661 , n1662 , n1666 , n1679 , 
n1682 , n1688 , n1696 , n1703 , n1719 , n1728 , n1731 , n1735 , n1736 , n1741 , 
n1743 , n1757 , n1758 , n1765 , n1766 , n1771 , n1774 , n1778 , n1779 , n1794 , 
n1805 , n1807 , n1809 , n1814 , n1821 , n1827 , n1829 , n1831 , n1838 , n1841 , 
n1852 , n1855 , n1861 , n1862 , n1869 , n1873 , n1879 , n1880 , n1886 , n1889 , 
n1892 , n1896 , n1897 , n1906 , n1912 , n1924 , n1925 , n1926 , n1932 , n1933 , 
n1936 , n1938 , n1940 , n1944 , n1947 , n1952 , n1953 , n1954 , n1958 , n1966 , 
n1991 , n2015 , n2025 , n2026 , n2029 , n2037 , n2043 , n2049 , n2051 , n2052 , 
n2061 , n2066 , n2093 , n2094 , n2102 , n2106 , n2116 , n2119 , n2121 , n2133 , 
n2144 , n2149 , n2157 , n2159 , n2170 , n2185 , n2189 , n2194 , n2195 , n2196 , 
n2210 , n2211 , n2212 , n2213 , n2222 , n2233 , n2236 , n2243 , n2257 , n2266 , 
n2281 , n2289 , n2304 , n2311 , n2315 , n2322 , n2352 , n2353 , n2358 , n2379 , 
n2414 , n2424 , n2430 , n2431 , n2436 , n2437 , n2443 , n2445 , n2446 , n2448 , 
n2449 , n2457 , n2459 , n2463 , n2467 , n2469 , n2470 , n2473 , n2477 , n2479 , 
n2482 , n2487 , n2491 , n2498 , n2516 , n2527 , n2529 , n2532 , n2533 , n2550 , 
n2561 , n2563 , n2564 , n2569 , n2584 , n2587 , n2589 , n2590 , n2592 , n2606 , 
n2613 , n2615 , n2616 , n2622 , n2628 , n2638 , n2644 , n2648 , n2650 , n2658 , 
n2685 , n2699 , n2703 , n2705 , n2706 , n2722 , n2731 , n2738 , n2768 , n2775 , 
n2780 , n2784 , n2788 , n2801 , n2803 , n2813 , n2820 , n2833 , n2839 , n2840 , 
n2848 , n2856 , n2865 , n2870 , n2872 , n2873 , n2888 , n2893 , n2896 , n2910 , 
n2918 , n2919 , n2925 , n2933 , n2938 , n2945 , n2954 , n2955 , n2967 , n2968 , 
n2975 , n2979 , n2984 , n2985 , n2986 , n2991 , n2995 , n3000 , n3002 , n3014 , 
n3016 , n3020 , n3027 , n3030 , n3031 , n3034 , n3048 , n3051 , n3060 , n3063 , 
n3087 , n3097 , n3101 , n3107 , n3115 , n3119 , n3124 , n3131 , n3137 , n3152 , 
n3155 , n3157 , n3171 , n3173 , n3189 , n3203 , n3208 , n3213 , n3215 , n3217 , 
n3220 , n3221 , n3224 , n3225 , n3227 , n3233 , n3236 , n3255 , n3258 , n3261 , 
n3268 , n3272 , n3279 , n3296 , n3303 , n3308 , n3310 , n3323 , n3336 , n3339 , 
n3355 , n3370 , n3373 , n3382 , n3390 , n3393 , n3399 , n3402 , n3416 , n3422 , 
n3423 , n3426 , n3427 , n3430 , n3434 , n3439 , n3441 , n3460 , n3471 , n3474 , 
n3477 , n3481 , n3484 , n3511 , n3512 , n3519 , n3528 , n3530 , n3547 , n3548 , 
n3551 , n3553 , n3563 , n3571 , n3574 , n3580 , n3581 , n3584 , n3598 , n3600 , 
n3603 , n3606 , n3608 , n3614 , n3621 , n3624 , n3629 , n3631 , n3633 , n3634 , 
n3643 , n3646 , n3648 , n3658 , n3663 , n3686 , n3691 , n3693 , n3696 , n3708 , 
n3711 , n3712 , n3713 , n3718 , n3726 , n3731 , n3739 , n3747 , n3749 , n3752 , 
n3754 , n3772 , n3782 , n3787 , n3808 , n3809 , n3810 , n3815 , n3819 , n3825 , 
n3836 , n3852 , n3856 , n3860 , n3867 , n3871 , n3873 , n3885 , n3897 , n3905 , 
n3914 );
    input n3 , n10 , n15 , n18 , n29 , n31 , n33 , n42 , n43 , 
n71 , n73 , n75 , n76 , n91 , n96 , n101 , n103 , n112 , n116 , 
n117 , n133 , n139 , n149 , n152 , n164 , n165 , n180 , n197 , n219 , 
n226 , n227 , n228 , n233 , n256 , n257 , n263 , n282 , n284 , n285 , 
n293 , n303 , n321 , n325 , n337 , n351 , n359 , n373 , n379 , n398 , 
n409 , n413 , n422 , n434 , n438 , n446 , n459 , n462 , n473 , n477 , 
n492 , n498 , n503 , n507 , n516 , n519 , n526 , n555 , n580 , n582 , 
n601 , n604 , n617 , n644 , n652 , n675 , n676 , n680 , n687 , n691 , 
n703 , n705 , n709 , n710 , n712 , n718 , n720 , n754 , n757 , n762 , 
n770 , n774 , n775 , n789 , n796 , n803 , n805 , n810 , n818 , n838 , 
n842 , n854 , n858 , n863 , n877 , n886 , n889 , n895 , n912 , n915 , 
n924 , n926 , n928 , n941 , n945 , n949 , n953 , n954 , n960 , n966 , 
n971 , n974 , n984 , n986 , n991 , n1013 , n1015 , n1027 , n1049 , n1051 , 
n1061 , n1062 , n1063 , n1086 , n1113 , n1114 , n1116 , n1130 , n1136 , n1144 , 
n1145 , n1150 , n1151 , n1163 , n1178 , n1179 , n1201 , n1216 , n1219 , n1229 , 
n1233 , n1253 , n1274 , n1276 , n1287 , n1305 , n1309 , n1314 , n1328 , n1332 , 
n1338 , n1347 , n1352 , n1360 , n1366 , n1372 , n1392 , n1393 , n1395 , n1403 , 
n1418 , n1428 , n1434 , n1470 , n1481 , n1491 , n1499 , n1506 , n1514 , n1533 , 
n1544 , n1548 , n1549 , n1559 , n1576 , n1583 , n1585 , n1615 , n1629 , n1631 , 
n1648 , n1661 , n1662 , n1666 , n1679 , n1688 , n1703 , n1719 , n1728 , n1731 , 
n1736 , n1743 , n1757 , n1758 , n1765 , n1766 , n1774 , n1778 , n1779 , n1794 , 
n1805 , n1807 , n1809 , n1814 , n1821 , n1827 , n1829 , n1831 , n1838 , n1841 , 
n1852 , n1861 , n1862 , n1873 , n1879 , n1880 , n1886 , n1892 , n1897 , n1906 , 
n1924 , n1925 , n1926 , n1932 , n1933 , n1938 , n1940 , n1944 , n1947 , n1954 , 
n1958 , n1966 , n1991 , n2026 , n2037 , n2043 , n2049 , n2051 , n2052 , n2061 , 
n2066 , n2102 , n2116 , n2119 , n2121 , n2133 , n2144 , n2149 , n2157 , n2170 , 
n2189 , n2194 , n2195 , n2196 , n2210 , n2211 , n2213 , n2222 , n2236 , n2243 , 
n2257 , n2266 , n2281 , n2289 , n2311 , n2322 , n2353 , n2358 , n2414 , n2424 , 
n2430 , n2431 , n2436 , n2437 , n2443 , n2445 , n2446 , n2448 , n2449 , n2457 , 
n2459 , n2463 , n2467 , n2469 , n2470 , n2473 , n2477 , n2479 , n2482 , n2487 , 
n2491 , n2498 , n2516 , n2527 , n2529 , n2533 , n2563 , n2564 , n2569 , n2587 , 
n2589 , n2590 , n2606 , n2613 , n2615 , n2616 , n2622 , n2628 , n2638 , n2644 , 
n2648 , n2658 , n2685 , n2699 , n2703 , n2705 , n2706 , n2722 , n2731 , n2738 , 
n2768 , n2775 , n2780 , n2784 , n2788 , n2813 , n2820 , n2848 , n2856 , n2865 , 
n2872 , n2893 , n2896 , n2910 , n2918 , n2919 , n2925 , n2933 , n2938 , n2945 , 
n2954 , n2955 , n2967 , n2968 , n2979 , n2984 , n2985 , n2986 , n2991 , n2995 , 
n3002 , n3016 , n3020 , n3027 , n3030 , n3034 , n3048 , n3051 , n3060 , n3063 , 
n3097 , n3101 , n3107 , n3119 , n3124 , n3137 , n3152 , n3155 , n3171 , n3189 , 
n3203 , n3208 , n3213 , n3215 , n3217 , n3220 , n3221 , n3224 , n3227 , n3233 , 
n3236 , n3255 , n3258 , n3261 , n3268 , n3272 , n3279 , n3296 , n3303 , n3308 , 
n3310 , n3323 , n3370 , n3373 , n3382 , n3390 , n3393 , n3399 , n3402 , n3416 , 
n3422 , n3423 , n3426 , n3427 , n3430 , n3434 , n3439 , n3441 , n3460 , n3471 , 
n3474 , n3477 , n3481 , n3484 , n3511 , n3512 , n3519 , n3528 , n3530 , n3547 , 
n3553 , n3571 , n3574 , n3581 , n3598 , n3600 , n3606 , n3608 , n3614 , n3621 , 
n3624 , n3629 , n3631 , n3633 , n3634 , n3643 , n3648 , n3658 , n3686 , n3693 , 
n3708 , n3711 , n3712 , n3713 , n3718 , n3726 , n3731 , n3739 , n3747 , n3749 , 
n3752 , n3754 , n3772 , n3787 , n3808 , n3809 , n3810 , n3815 , n3819 , n3825 , 
n3836 , n3852 , n3856 , n3860 , n3867 , n3871 , n3873 , n3885 , n3897 , n3905 , 
n3914 ;
    output n1 , n20 , n49 , n52 , n69 , n107 , n114 , n135 , n200 , 
n235 , n292 , n297 , n313 , n326 , n330 , n334 , n336 , n399 , n463 , 
n484 , n524 , n531 , n559 , n575 , n587 , n636 , n647 , n749 , n751 , 
n784 , n785 , n812 , n834 , n873 , n897 , n932 , n958 , n963 , n983 , 
n1084 , n1094 , n1105 , n1122 , n1143 , n1161 , n1204 , n1235 , n1238 , n1241 , 
n1260 , n1266 , n1268 , n1277 , n1297 , n1301 , n1405 , n1458 , n1461 , n1503 , 
n1504 , n1558 , n1616 , n1625 , n1632 , n1660 , n1682 , n1696 , n1735 , n1741 , 
n1771 , n1855 , n1869 , n1889 , n1896 , n1912 , n1936 , n1952 , n1953 , n2015 , 
n2025 , n2029 , n2093 , n2094 , n2106 , n2159 , n2185 , n2212 , n2233 , n2304 , 
n2315 , n2352 , n2379 , n2532 , n2550 , n2561 , n2584 , n2592 , n2650 , n2801 , 
n2803 , n2833 , n2839 , n2840 , n2870 , n2873 , n2888 , n2975 , n3000 , n3014 , 
n3031 , n3087 , n3115 , n3131 , n3157 , n3173 , n3225 , n3336 , n3339 , n3355 , 
n3548 , n3551 , n3563 , n3580 , n3584 , n3603 , n3646 , n3663 , n3691 , n3696 , 
n3782 ;
    wire n0 , n2 , n4 , n5 , n6 , n7 , n8 , n9 , n11 , 
n12 , n13 , n14 , n16 , n17 , n19 , n21 , n22 , n23 , n24 , 
n25 , n26 , n27 , n28 , n30 , n32 , n34 , n35 , n36 , n37 , 
n38 , n39 , n40 , n41 , n44 , n45 , n46 , n47 , n48 , n50 , 
n51 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , 
n62 , n63 , n64 , n65 , n66 , n67 , n68 , n70 , n72 , n74 , 
n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , 
n87 , n88 , n89 , n90 , n92 , n93 , n94 , n95 , n97 , n98 , 
n99 , n100 , n102 , n104 , n105 , n106 , n108 , n109 , n110 , n111 , 
n113 , n115 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , 
n126 , n127 , n128 , n129 , n130 , n131 , n132 , n134 , n136 , n137 , 
n138 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , 
n150 , n151 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
n161 , n162 , n163 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , 
n173 , n174 , n175 , n176 , n177 , n178 , n179 , n181 , n182 , n183 , 
n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , 
n194 , n195 , n196 , n198 , n199 , n201 , n202 , n203 , n204 , n205 , 
n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , 
n216 , n217 , n218 , n220 , n221 , n222 , n223 , n224 , n225 , n229 , 
n230 , n231 , n232 , n234 , n236 , n237 , n238 , n239 , n240 , n241 , 
n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , 
n252 , n253 , n254 , n255 , n258 , n259 , n260 , n261 , n262 , n264 , 
n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , 
n275 , n276 , n277 , n278 , n279 , n280 , n281 , n283 , n286 , n287 , 
n288 , n289 , n290 , n291 , n294 , n295 , n296 , n298 , n299 , n300 , 
n301 , n302 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , 
n312 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n322 , n323 , 
n324 , n327 , n328 , n329 , n331 , n332 , n333 , n335 , n338 , n339 , 
n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
n350 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n360 , n361 , 
n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , 
n372 , n374 , n375 , n376 , n377 , n378 , n380 , n381 , n382 , n383 , 
n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , 
n394 , n395 , n396 , n397 , n400 , n401 , n402 , n403 , n404 , n405 , 
n406 , n407 , n408 , n410 , n411 , n412 , n414 , n415 , n416 , n417 , 
n418 , n419 , n420 , n421 , n423 , n424 , n425 , n426 , n427 , n428 , 
n429 , n430 , n431 , n432 , n433 , n435 , n436 , n437 , n439 , n440 , 
n441 , n442 , n443 , n444 , n445 , n447 , n448 , n449 , n450 , n451 , 
n452 , n453 , n454 , n455 , n456 , n457 , n458 , n460 , n461 , n464 , 
n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n474 , n475 , 
n476 , n478 , n479 , n480 , n481 , n482 , n483 , n485 , n486 , n487 , 
n488 , n489 , n490 , n491 , n493 , n494 , n495 , n496 , n497 , n499 , 
n500 , n501 , n502 , n504 , n505 , n506 , n508 , n509 , n510 , n511 , 
n512 , n513 , n514 , n515 , n517 , n518 , n520 , n521 , n522 , n523 , 
n525 , n527 , n528 , n529 , n530 , n532 , n533 , n534 , n535 , n536 , 
n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , 
n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n556 , n557 , 
n558 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , 
n569 , n570 , n571 , n572 , n573 , n574 , n576 , n577 , n578 , n579 , 
n581 , n583 , n584 , n585 , n586 , n588 , n589 , n590 , n591 , n592 , 
n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n602 , n603 , 
n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
n615 , n616 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , 
n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , 
n637 , n638 , n639 , n640 , n641 , n642 , n643 , n645 , n646 , n648 , 
n649 , n650 , n651 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
n670 , n671 , n672 , n673 , n674 , n677 , n678 , n679 , n681 , n682 , 
n683 , n684 , n685 , n686 , n688 , n689 , n690 , n692 , n693 , n694 , 
n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n704 , n706 , 
n707 , n708 , n711 , n713 , n714 , n715 , n716 , n717 , n719 , n721 , 
n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , 
n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , 
n742 , n743 , n744 , n745 , n746 , n747 , n748 , n750 , n752 , n753 , 
n755 , n756 , n758 , n759 , n760 , n761 , n763 , n764 , n765 , n766 , 
n767 , n768 , n769 , n771 , n772 , n773 , n776 , n777 , n778 , n779 , 
n780 , n781 , n782 , n783 , n786 , n787 , n788 , n790 , n791 , n792 , 
n793 , n794 , n795 , n797 , n798 , n799 , n800 , n801 , n802 , n804 , 
n806 , n807 , n808 , n809 , n811 , n813 , n814 , n815 , n816 , n817 , 
n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , 
n829 , n830 , n831 , n832 , n833 , n835 , n836 , n837 , n839 , n840 , 
n841 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , 
n852 , n853 , n855 , n856 , n857 , n859 , n860 , n861 , n862 , n864 , 
n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n874 , n875 , 
n876 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n887 , 
n888 , n890 , n891 , n892 , n893 , n894 , n896 , n898 , n899 , n900 , 
n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , 
n911 , n913 , n914 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , 
n923 , n925 , n927 , n929 , n930 , n931 , n933 , n934 , n935 , n936 , 
n937 , n938 , n939 , n940 , n942 , n943 , n944 , n946 , n947 , n948 , 
n950 , n951 , n952 , n955 , n956 , n957 , n959 , n961 , n962 , n964 , 
n965 , n967 , n968 , n969 , n970 , n972 , n973 , n975 , n976 , n977 , 
n978 , n979 , n980 , n981 , n982 , n985 , n987 , n988 , n989 , n990 , 
n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , 
n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , 
n1012 , n1014 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , 
n1024 , n1025 , n1026 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , 
n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , 
n1045 , n1046 , n1047 , n1048 , n1050 , n1052 , n1053 , n1054 , n1055 , n1056 , 
n1057 , n1058 , n1059 , n1060 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
n1080 , n1081 , n1082 , n1083 , n1085 , n1087 , n1088 , n1089 , n1090 , n1091 , 
n1092 , n1093 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , 
n1103 , n1104 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1115 , 
n1117 , n1118 , n1119 , n1120 , n1121 , n1123 , n1124 , n1125 , n1126 , n1127 , 
n1128 , n1129 , n1131 , n1132 , n1133 , n1134 , n1135 , n1137 , n1138 , n1139 , 
n1140 , n1141 , n1142 , n1146 , n1147 , n1148 , n1149 , n1152 , n1153 , n1154 , 
n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1162 , n1164 , n1165 , n1166 , 
n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , 
n1177 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , 
n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , 
n1199 , n1200 , n1202 , n1203 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , 
n1211 , n1212 , n1213 , n1214 , n1215 , n1217 , n1218 , n1220 , n1221 , n1222 , 
n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1230 , n1231 , n1232 , n1234 , 
n1236 , n1237 , n1239 , n1240 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , 
n1248 , n1249 , n1250 , n1251 , n1252 , n1254 , n1255 , n1256 , n1257 , n1258 , 
n1259 , n1261 , n1262 , n1263 , n1264 , n1265 , n1267 , n1269 , n1270 , n1271 , 
n1272 , n1273 , n1275 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , 
n1285 , n1286 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , 
n1296 , n1298 , n1299 , n1300 , n1302 , n1303 , n1304 , n1306 , n1307 , n1308 , 
n1310 , n1311 , n1312 , n1313 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , 
n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1329 , n1330 , n1331 , 
n1333 , n1334 , n1335 , n1336 , n1337 , n1339 , n1340 , n1341 , n1342 , n1343 , 
n1344 , n1345 , n1346 , n1348 , n1349 , n1350 , n1351 , n1353 , n1354 , n1355 , 
n1356 , n1357 , n1358 , n1359 , n1361 , n1362 , n1363 , n1364 , n1365 , n1367 , 
n1368 , n1369 , n1370 , n1371 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , 
n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , 
n1389 , n1390 , n1391 , n1394 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , 
n1402 , n1404 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , 
n1414 , n1415 , n1416 , n1417 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , 
n1425 , n1426 , n1427 , n1429 , n1430 , n1431 , n1432 , n1433 , n1435 , n1436 , 
n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , 
n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , 
n1457 , n1459 , n1460 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , 
n1469 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
n1480 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , 
n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1500 , n1501 , n1502 , 
n1505 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1515 , n1516 , 
n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , 
n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1534 , n1535 , n1536 , n1537 , 
n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1545 , n1546 , n1547 , n1550 , 
n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1560 , n1561 , n1562 , 
n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , 
n1573 , n1574 , n1575 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1584 , 
n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , 
n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , 
n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1617 , 
n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1626 , n1627 , n1628 , 
n1630 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , 
n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1649 , n1650 , n1651 , n1652 , 
n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1663 , n1664 , n1665 , 
n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , 
n1677 , n1678 , n1680 , n1681 , n1683 , n1684 , n1685 , n1686 , n1687 , n1689 , 
n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1697 , n1698 , n1699 , n1700 , 
n1701 , n1702 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , 
n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1720 , n1721 , n1722 , 
n1723 , n1724 , n1725 , n1726 , n1727 , n1729 , n1730 , n1732 , n1733 , n1734 , 
n1737 , n1738 , n1739 , n1740 , n1742 , n1744 , n1745 , n1746 , n1747 , n1748 , 
n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1759 , n1760 , 
n1761 , n1762 , n1763 , n1764 , n1767 , n1768 , n1769 , n1770 , n1772 , n1773 , 
n1775 , n1776 , n1777 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , 
n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1795 , n1796 , n1797 , 
n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1806 , n1808 , n1810 , 
n1811 , n1812 , n1813 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1822 , 
n1823 , n1824 , n1825 , n1826 , n1828 , n1830 , n1832 , n1833 , n1834 , n1835 , 
n1836 , n1837 , n1839 , n1840 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , 
n1848 , n1849 , n1850 , n1851 , n1853 , n1854 , n1856 , n1857 , n1858 , n1859 , 
n1860 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1870 , n1871 , n1872 , 
n1874 , n1875 , n1876 , n1877 , n1878 , n1881 , n1882 , n1883 , n1884 , n1885 , 
n1887 , n1888 , n1890 , n1891 , n1893 , n1894 , n1895 , n1898 , n1899 , n1900 , 
n1901 , n1902 , n1903 , n1904 , n1905 , n1907 , n1908 , n1909 , n1910 , n1911 , 
n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , 
n1923 , n1927 , n1928 , n1929 , n1930 , n1931 , n1934 , n1935 , n1937 , n1939 , 
n1941 , n1942 , n1943 , n1945 , n1946 , n1948 , n1949 , n1950 , n1951 , n1955 , 
n1956 , n1957 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1967 , 
n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , 
n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , 
n1988 , n1989 , n1990 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , 
n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , 
n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2016 , n2017 , n2018 , n2019 , 
n2020 , n2021 , n2022 , n2023 , n2024 , n2027 , n2028 , n2030 , n2031 , n2032 , 
n2033 , n2034 , n2035 , n2036 , n2038 , n2039 , n2040 , n2041 , n2042 , n2044 , 
n2045 , n2046 , n2047 , n2048 , n2050 , n2053 , n2054 , n2055 , n2056 , n2057 , 
n2058 , n2059 , n2060 , n2062 , n2063 , n2064 , n2065 , n2067 , n2068 , n2069 , 
n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
n2090 , n2091 , n2092 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , 
n2103 , n2104 , n2105 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , 
n2114 , n2115 , n2117 , n2118 , n2120 , n2122 , n2123 , n2124 , n2125 , n2126 , 
n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2134 , n2135 , n2136 , n2137 , 
n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2145 , n2146 , n2147 , n2148 , 
n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2158 , n2160 , n2161 , 
n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2171 , n2172 , 
n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , 
n2183 , n2184 , n2186 , n2187 , n2188 , n2190 , n2191 , n2192 , n2193 , n2197 , 
n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , 
n2208 , n2209 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , 
n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , 
n2234 , n2235 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2244 , n2245 , 
n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , 
n2256 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2267 , 
n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , 
n2278 , n2279 , n2280 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , 
n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
n2300 , n2301 , n2302 , n2303 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , 
n2312 , n2313 , n2314 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2323 , 
n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , 
n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , 
n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2354 , n2355 , 
n2356 , n2357 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , 
n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , 
n2377 , n2378 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , 
n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , 
n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , 
n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2415 , n2416 , n2417 , n2418 , 
n2419 , n2420 , n2421 , n2422 , n2423 , n2425 , n2426 , n2427 , n2428 , n2429 , 
n2432 , n2433 , n2434 , n2435 , n2438 , n2439 , n2440 , n2441 , n2442 , n2444 , 
n2447 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2458 , n2460 , 
n2461 , n2462 , n2464 , n2465 , n2466 , n2468 , n2471 , n2472 , n2474 , n2475 , 
n2476 , n2478 , n2480 , n2481 , n2483 , n2484 , n2485 , n2486 , n2488 , n2489 , 
n2490 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2499 , n2500 , n2501 , 
n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , 
n2512 , n2513 , n2514 , n2515 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , 
n2523 , n2524 , n2525 , n2526 , n2528 , n2530 , n2531 , n2534 , n2535 , n2536 , 
n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , 
n2547 , n2548 , n2549 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , 
n2558 , n2559 , n2560 , n2562 , n2565 , n2566 , n2567 , n2568 , n2570 , n2571 , 
n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , 
n2582 , n2583 , n2585 , n2586 , n2588 , n2591 , n2593 , n2594 , n2595 , n2596 , 
n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2607 , 
n2608 , n2609 , n2610 , n2611 , n2612 , n2614 , n2617 , n2618 , n2619 , n2620 , 
n2621 , n2623 , n2624 , n2625 , n2626 , n2627 , n2629 , n2630 , n2631 , n2632 , 
n2633 , n2634 , n2635 , n2636 , n2637 , n2639 , n2640 , n2641 , n2642 , n2643 , 
n2645 , n2646 , n2647 , n2649 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , 
n2657 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , 
n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , 
n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2686 , n2687 , n2688 , 
n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , 
n2700 , n2701 , n2702 , n2704 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , 
n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2723 , 
n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2732 , n2733 , n2734 , 
n2735 , n2736 , n2737 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , 
n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , 
n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , 
n2766 , n2767 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2776 , n2777 , 
n2778 , n2779 , n2781 , n2782 , n2783 , n2785 , n2786 , n2787 , n2789 , n2790 , 
n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , 
n2802 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , 
n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2821 , n2822 , n2823 , n2824 , 
n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2834 , n2835 , 
n2836 , n2837 , n2838 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , 
n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2857 , n2858 , n2859 , 
n2860 , n2861 , n2862 , n2863 , n2864 , n2866 , n2867 , n2868 , n2869 , n2871 , 
n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , 
n2884 , n2885 , n2886 , n2887 , n2889 , n2890 , n2891 , n2892 , n2894 , n2895 , 
n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , 
n2907 , n2908 , n2909 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , 
n2920 , n2921 , n2922 , n2923 , n2924 , n2926 , n2927 , n2928 , n2929 , n2930 , 
n2931 , n2932 , n2934 , n2935 , n2936 , n2937 , n2939 , n2940 , n2941 , n2942 , 
n2943 , n2944 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , 
n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , 
n2966 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2976 , n2977 , n2978 , 
n2980 , n2981 , n2982 , n2983 , n2987 , n2988 , n2989 , n2990 , n2992 , n2993 , 
n2994 , n2996 , n2997 , n2998 , n2999 , n3001 , n3003 , n3004 , n3005 , n3006 , 
n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3015 , n3017 , n3018 , 
n3019 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3028 , n3029 , n3032 , 
n3033 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , 
n3044 , n3045 , n3046 , n3047 , n3049 , n3050 , n3052 , n3053 , n3054 , n3055 , 
n3056 , n3057 , n3058 , n3059 , n3061 , n3062 , n3064 , n3065 , n3066 , n3067 , 
n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , 
n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3088 , 
n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3098 , n3099 , 
n3100 , n3102 , n3103 , n3104 , n3105 , n3106 , n3108 , n3109 , n3110 , n3111 , 
n3112 , n3113 , n3114 , n3116 , n3117 , n3118 , n3120 , n3121 , n3122 , n3123 , 
n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3132 , n3133 , n3134 , n3135 , 
n3136 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , 
n3147 , n3148 , n3149 , n3150 , n3151 , n3153 , n3154 , n3156 , n3158 , n3159 , 
n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
n3170 , n3172 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , 
n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3190 , n3191 , n3192 , 
n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , 
n3204 , n3205 , n3206 , n3207 , n3209 , n3210 , n3211 , n3212 , n3214 , n3216 , 
n3218 , n3219 , n3222 , n3223 , n3226 , n3228 , n3229 , n3230 , n3231 , n3232 , 
n3234 , n3235 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , 
n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , 
n3256 , n3257 , n3259 , n3260 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , 
n3269 , n3270 , n3271 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3280 , 
n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , 
n3291 , n3292 , n3293 , n3294 , n3295 , n3297 , n3298 , n3299 , n3300 , n3301 , 
n3302 , n3304 , n3305 , n3306 , n3307 , n3309 , n3311 , n3312 , n3313 , n3314 , 
n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3324 , n3325 , 
n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , 
n3337 , n3338 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , 
n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3356 , n3357 , n3358 , 
n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , 
n3369 , n3371 , n3372 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , 
n3381 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3391 , n3392 , 
n3394 , n3395 , n3396 , n3397 , n3398 , n3400 , n3401 , n3403 , n3404 , n3405 , 
n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , 
n3417 , n3418 , n3419 , n3420 , n3421 , n3424 , n3425 , n3428 , n3429 , n3431 , 
n3432 , n3433 , n3435 , n3436 , n3437 , n3438 , n3440 , n3442 , n3443 , n3444 , 
n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , 
n3455 , n3456 , n3457 , n3458 , n3459 , n3461 , n3462 , n3463 , n3464 , n3465 , 
n3466 , n3467 , n3468 , n3469 , n3470 , n3472 , n3473 , n3475 , n3476 , n3478 , 
n3479 , n3480 , n3482 , n3483 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , 
n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3520 , n3521 , n3522 , n3523 , 
n3524 , n3525 , n3526 , n3527 , n3529 , n3531 , n3532 , n3533 , n3534 , n3535 , 
n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , 
n3546 , n3549 , n3550 , n3552 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
n3560 , n3561 , n3562 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , 
n3572 , n3573 , n3575 , n3576 , n3577 , n3578 , n3579 , n3582 , n3583 , n3585 , 
n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , 
n3596 , n3597 , n3599 , n3601 , n3602 , n3604 , n3605 , n3607 , n3609 , n3610 , 
n3611 , n3612 , n3613 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3622 , 
n3623 , n3625 , n3626 , n3627 , n3628 , n3630 , n3632 , n3635 , n3636 , n3637 , 
n3638 , n3639 , n3640 , n3641 , n3642 , n3644 , n3645 , n3647 , n3649 , n3650 , 
n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3659 , n3660 , n3661 , 
n3662 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , 
n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , 
n3683 , n3684 , n3685 , n3687 , n3688 , n3689 , n3690 , n3692 , n3694 , n3695 , 
n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , 
n3707 , n3709 , n3710 , n3714 , n3715 , n3716 , n3717 , n3719 , n3720 , n3721 , 
n3722 , n3723 , n3724 , n3725 , n3727 , n3728 , n3729 , n3730 , n3732 , n3733 , 
n3734 , n3735 , n3736 , n3737 , n3738 , n3740 , n3741 , n3742 , n3743 , n3744 , 
n3745 , n3746 , n3748 , n3750 , n3751 , n3753 , n3755 , n3756 , n3757 , n3758 , 
n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , 
n3769 , n3770 , n3771 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
n3780 , n3781 , n3783 , n3784 , n3785 , n3786 , n3788 , n3789 , n3790 , n3791 , 
n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , 
n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3811 , n3812 , n3813 , n3814 , 
n3816 , n3817 , n3818 , n3820 , n3821 , n3822 , n3823 , n3824 , n3826 , n3827 , 
n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3837 , n3838 , 
n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , 
n3849 , n3850 , n3851 , n3853 , n3854 , n3855 , n3857 , n3858 , n3859 , n3861 , 
n3862 , n3863 , n3864 , n3865 , n3866 , n3868 , n3869 , n3870 , n3872 , n3874 , 
n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , 
n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , 
n3896 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3906 , n3907 , 
n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3915 , n3916 , n3917 , n3918 , 
n3919 ;
    and g0 ( n2113 , n1673 , n680 );
    or g1 ( n3601 , n470 , n474 );
    not g2 ( n913 , n3097 );
    nor g3 ( n2042 , n2348 , n3844 );
    not g4 ( n2073 , n3027 );
    nor g5 ( n3165 , n842 , n404 );
    not g6 ( n2319 , n285 );
    or g7 ( n647 , n1946 , n1345 );
    and g8 ( n2932 , n1188 , n877 );
    and g9 ( n2410 , n693 , n2683 );
    and g10 ( n3671 , n1864 , n228 );
    nor g11 ( n1056 , n3323 , n2374 );
    nor g12 ( n2057 , n874 , n3659 );
    or g13 ( n2039 , n3460 , n3449 );
    and g14 ( n891 , n1692 , n2196 );
    or g15 ( n2829 , n516 , n1101 );
    not g16 ( n921 , n3856 );
    and g17 ( n2252 , n2708 , n1921 );
    or g18 ( n657 , n889 , n2929 );
    not g19 ( n2695 , n2457 );
    and g20 ( n1568 , n643 , n2437 );
    nor g21 ( n2660 , n821 , n2339 );
    and g22 ( n1039 , n763 , n3901 );
    not g23 ( n181 , n3527 );
    nor g24 ( n1680 , n3534 , n3496 );
    or g25 ( n260 , n2311 , n1898 );
    buf g26 ( n1207 , n3900 );
    not g27 ( n1252 , n1794 );
    not g28 ( n747 , n3379 );
    nor g29 ( n1485 , n379 , n1574 );
    and g30 ( n756 , n3615 , n3094 );
    not g31 ( n2777 , n3427 );
    and g32 ( n1607 , n3196 , n2729 );
    or g33 ( n1379 , n1481 , n1101 );
    or g34 ( n1337 , n3327 , n1460 );
    or g35 ( n1896 , n1383 , n3702 );
    nor g36 ( n956 , n2613 , n3202 );
    or g37 ( n1106 , n2569 , n3169 );
    nor g38 ( n499 , n2995 , n3733 );
    nor g39 ( n781 , n2979 , n3707 );
    or g40 ( n2973 , n3711 , n3707 );
    and g41 ( n3757 , n396 , n1170 );
    and g42 ( n1536 , n608 , n459 );
    not g43 ( n3372 , n838 );
    not g44 ( n3480 , n1627 );
    or g45 ( n3607 , n1464 , n2916 );
    or g46 ( n1810 , n2588 , n3701 );
    nor g47 ( n1222 , n3891 , n1540 );
    or g48 ( n63 , n757 , n1131 );
    or g49 ( n2095 , n926 , n2607 );
    nor g50 ( n1763 , n2820 , n115 );
    or g51 ( n2877 , n2527 , n2996 );
    and g52 ( n979 , n279 , n1136 );
    or g53 ( n3408 , n1852 , n3903 );
    not g54 ( n3733 , n76 );
    not g55 ( n669 , n1403 );
    or g56 ( n521 , n2823 , n2598 );
    nor g57 ( n309 , n2761 , n217 );
    nor g58 ( n3915 , n351 , n380 );
    and g59 ( n3207 , n1647 , n1648 );
    or g60 ( n1155 , n2857 , n1459 );
    and g61 ( n2165 , n1489 , n666 );
    nor g62 ( n3637 , n2189 , n1124 );
    and g63 ( n2709 , n2331 , n1666 );
    and g64 ( n2696 , n679 , n2139 );
    or g65 ( n3542 , n3193 , n3649 );
    not g66 ( n2798 , n3308 );
    and g67 ( n2920 , n2713 , n3477 );
    and g68 ( n1509 , n655 , n1839 );
    nor g69 ( n885 , n3784 , n3661 );
    not g70 ( n1505 , n2332 );
    not g71 ( n2834 , n3528 );
    nor g72 ( n3147 , n1313 , n802 );
    not g73 ( n3893 , n1666 );
    or g74 ( n439 , n1868 , n3083 );
    and g75 ( n386 , n483 , n2942 );
    and g76 ( n2174 , n3659 , n3443 );
    or g77 ( n1488 , n366 , n2930 );
    or g78 ( n1118 , n2515 , n3573 );
    nor g79 ( n2948 , n1437 , n3452 );
    and g80 ( n1980 , n1893 , n1066 );
    not g81 ( n2759 , n3633 );
    or g82 ( n3720 , n1631 , n2996 );
    and g83 ( n1273 , n2456 , n2449 );
    or g84 ( n301 , n133 , n908 );
    and g85 ( n1983 , n1613 , n327 );
    or g86 ( n3248 , n2232 , n2135 );
    and g87 ( n1280 , n1096 , n38 );
    or g88 ( n1937 , n257 , n295 );
    and g89 ( n216 , n3902 , n709 );
    or g90 ( n911 , n710 , n1898 );
    nor g91 ( n1317 , n1808 , n1139 );
    nor g92 ( n3453 , n2165 , n342 );
    not g93 ( n2147 , n2671 );
    or g94 ( n423 , n2442 , n2117 );
    not g95 ( n2393 , n3506 );
    and g96 ( n3098 , n1895 , n3358 );
    and g97 ( n1290 , n3672 , n2006 );
    nor g98 ( n319 , n3372 , n38 );
    and g99 ( n99 , n1635 , n316 );
    or g100 ( n1630 , n753 , n2456 );
    and g101 ( n1212 , n684 , n7 );
    not g102 ( n401 , n2859 );
    and g103 ( n1005 , n1388 , n666 );
    nor g104 ( n2369 , n2494 , n287 );
    nor g105 ( n3229 , n3434 , n1922 );
    and g106 ( n839 , n597 , n2969 );
    and g107 ( n1848 , n142 , n2633 );
    nor g108 ( n3831 , n2516 , n2607 );
    and g109 ( n1663 , n2392 , n1371 );
    and g110 ( n2623 , n1598 , n2700 );
    or g111 ( n1942 , n1040 , n14 );
    not g112 ( n338 , n3385 );
    nor g113 ( n1571 , n2116 , n3622 );
    or g114 ( n472 , n966 , n3692 );
    and g115 ( n1976 , n3167 , n94 );
    and g116 ( n1882 , n1370 , n3309 );
    not g117 ( n24 , n1675 );
    not g118 ( n892 , n924 );
    or g119 ( n2106 , n1793 , n2244 );
    or g120 ( n3577 , n2590 , n2810 );
    not g121 ( n3597 , n3101 );
    nor g122 ( n2626 , n2133 , n1554 );
    not g123 ( n2756 , n818 );
    nor g124 ( n3820 , n3609 , n1356 );
    not g125 ( n3883 , n1524 );
    and g126 ( n3175 , n2455 , n2979 );
    not g127 ( n1011 , n2408 );
    and g128 ( n1721 , n476 , n1439 );
    not g129 ( n2032 , n3379 );
    not g130 ( n478 , n1779 );
    or g131 ( n3774 , n2915 , n1525 );
    not g132 ( n1490 , n2257 );
    and g133 ( n90 , n1125 , n1306 );
    and g134 ( n2802 , n1016 , n2202 );
    and g135 ( n1507 , n3078 , n2822 );
    not g136 ( n475 , n3203 );
    and g137 ( n3527 , n3607 , n1185 );
    and g138 ( n1919 , n1031 , n3845 );
    and g139 ( n3751 , n2860 , n3217 );
    nor g140 ( n1335 , n1916 , n1974 );
    and g141 ( n239 , n1384 , n1430 );
    and g142 ( n2328 , n2757 , n3574 );
    not g143 ( n3500 , n3439 );
    not g144 ( n2494 , n259 );
    or g145 ( n3888 , n1782 , n682 );
    and g146 ( n160 , n3210 , n3526 );
    and g147 ( n539 , n696 , n3068 );
    not g148 ( n1257 , n1544 );
    nor g149 ( n1464 , n3642 , n1528 );
    nor g150 ( n3084 , n225 , n3596 );
    or g151 ( n489 , n1134 , n1212 );
    or g152 ( n2239 , n2196 , n509 );
    buf g153 ( n3379 , n3666 );
    or g154 ( n1804 , n705 , n2032 );
    not g155 ( n1823 , n2991 );
    and g156 ( n349 , n2951 , n1627 );
    nor g157 ( n2503 , n2431 , n1993 );
    and g158 ( n639 , n1582 , n1467 );
    nor g159 ( n952 , n2533 , n2607 );
    or g160 ( n3322 , n3189 , n1165 );
    nor g161 ( n840 , n3625 , n429 );
    nor g162 ( n1959 , n3279 , n792 );
    or g163 ( n702 , n1328 , n3449 );
    or g164 ( n2779 , n3905 , n1207 );
    nor g165 ( n642 , n3063 , n3486 );
    or g166 ( n2143 , n2470 , n3910 );
    not g167 ( n1249 , n1761 );
    nor g168 ( n3145 , n3382 , n3184 );
    and g169 ( n2458 , n2153 , n1080 );
    not g170 ( n1692 , n149 );
    not g171 ( n3514 , n229 );
    not g172 ( n2280 , n434 );
    not g173 ( n3909 , n2868 );
    and g174 ( n2885 , n2769 , n3504 );
    or g175 ( n1369 , n1276 , n3505 );
    not g176 ( n1715 , n75 );
    nor g177 ( n573 , n3848 , n2665 );
    and g178 ( n2455 , n2921 , n3143 );
    or g179 ( n2240 , n3165 , n2076 );
    nor g180 ( n2117 , n1559 , n722 );
    nor g181 ( n3454 , n2435 , n3223 );
    or g182 ( n2594 , n2775 , n1207 );
    nor g183 ( n3623 , n1809 , n1554 );
    nor g184 ( n3118 , n31 , n3153 );
    or g185 ( n1741 , n2340 , n1399 );
    and g186 ( n903 , n1984 , n3577 );
    not g187 ( n1193 , n1305 );
    and g188 ( n1068 , n3284 , n3393 );
    or g189 ( n2212 , n309 , n875 );
    not g190 ( n914 , n3710 );
    not g191 ( n501 , n2589 );
    nor g192 ( n3562 , n1940 , n2607 );
    nor g193 ( n1822 , n3523 , n585 );
    not g194 ( n2761 , n1883 );
    nor g195 ( n1964 , n346 , n3139 );
    and g196 ( n611 , n262 , n2666 );
    or g197 ( n286 , n1513 , n864 );
    or g198 ( n3156 , n1114 , n1188 );
    or g199 ( n2734 , n3089 , n3201 );
    or g200 ( n1467 , n1794 , n150 );
    and g201 ( n2520 , n546 , n3677 );
    not g202 ( n1796 , n895 );
    nor g203 ( n3420 , n3756 , n78 );
    not g204 ( n772 , n1027 );
    or g205 ( n3641 , n245 , n3469 );
    not g206 ( n888 , n1428 );
    and g207 ( n2282 , n2629 , n3718 );
    and g208 ( n2580 , n2980 , n832 );
    not g209 ( n3133 , n91 );
    not g210 ( n3575 , n877 );
    or g211 ( n2476 , n2141 , n2493 );
    and g212 ( n170 , n1373 , n3392 );
    or g213 ( n833 , n668 , n2339 );
    or g214 ( n3425 , n3740 , n3673 );
    nor g215 ( n3110 , n3790 , n2486 );
    nor g216 ( n1157 , n51 , n2870 );
    not g217 ( n2701 , n1631 );
    and g218 ( n1420 , n1860 , n3026 );
    and g219 ( n1498 , n1462 , n1680 );
    or g220 ( n444 , n2759 , n513 );
    and g221 ( n2010 , n3483 , n525 );
    or g222 ( n857 , n2563 , n3742 );
    and g223 ( n451 , n3114 , n475 );
    or g224 ( n343 , n2812 , n2394 );
    not g225 ( n1601 , n2974 );
    and g226 ( n244 , n509 , n718 );
    not g227 ( n2295 , n2170 );
    and g228 ( n225 , n3256 , n1505 );
    or g229 ( n1256 , n1107 , n3846 );
    not g230 ( n105 , n1279 );
    or g231 ( n275 , n3699 , n1487 );
    not g232 ( n1510 , n303 );
    not g233 ( n3865 , n706 );
    or g234 ( n1124 , n532 , n2363 );
    and g235 ( n566 , n2494 , n1839 );
    or g236 ( n2277 , n1703 , n3466 );
    nor g237 ( n1609 , n3504 , n1640 );
    and g238 ( n1356 , n2761 , n3618 );
    or g239 ( n759 , n863 , n3449 );
    and g240 ( n3565 , n3475 , n2450 );
    or g241 ( n1411 , n659 , n223 );
    and g242 ( n1557 , n2167 , n2459 );
    or g243 ( n2976 , n3860 , n2607 );
    and g244 ( n261 , n1893 , n1423 );
    nor g245 ( n1180 , n1906 , n2234 );
    or g246 ( n2679 , n1886 , n1916 );
    not g247 ( n468 , n3002 );
    buf g248 ( n1898 , n1694 );
    not g249 ( n1537 , n3581 );
    nor g250 ( n746 , n3433 , n3417 );
    and g251 ( n2545 , n2256 , n2954 );
    not g252 ( n178 , n2625 );
    or g253 ( n1468 , n2119 , n1916 );
    nor g254 ( n1240 , n1347 , n1028 );
    and g255 ( n2495 , n340 , n1343 );
    and g256 ( n2292 , n3169 , n519 );
    or g257 ( n1082 , n1325 , n824 );
    not g258 ( n2652 , n2946 );
    or g259 ( n2983 , n3512 , n3169 );
    not g260 ( n177 , n498 );
    or g261 ( n155 , n3107 , n1916 );
    not g262 ( n1702 , n2479 );
    or g263 ( n738 , n3815 , n2929 );
    and g264 ( n2712 , n1033 , n1879 );
    or g265 ( n844 , n2270 , n343 );
    or g266 ( n2218 , n3749 , n3015 );
    not g267 ( n602 , n3468 );
    or g268 ( n631 , n652 , n2629 );
    and g269 ( n3191 , n929 , n362 );
    and g270 ( n2826 , n685 , n1872 );
    or g271 ( n3529 , n3020 , n3262 );
    nor g272 ( n2286 , n3136 , n3721 );
    and g273 ( n3833 , n3228 , n89 );
    or g274 ( n3343 , n2210 , n1620 );
    not g275 ( n1859 , n1043 );
    not g276 ( n2632 , n635 );
    nor g277 ( n977 , n1480 , n3136 );
    nor g278 ( n2943 , n790 , n2764 );
    nor g279 ( n1330 , n1774 , n1554 );
    not g280 ( n2345 , n2651 );
    not g281 ( n3421 , n2780 );
    nor g282 ( n851 , n3547 , n1943 );
    or g283 ( n3285 , n103 , n3887 );
    and g284 ( n2389 , n3522 , n120 );
    not g285 ( n627 , n666 );
    and g286 ( n3117 , n1404 , n3796 );
    nor g287 ( n3388 , n3600 , n2152 );
    not g288 ( n1768 , n2281 );
    or g289 ( n2771 , n3168 , n1658 );
    and g290 ( n1874 , n2599 , n3757 );
    and g291 ( n579 , n902 , n1036 );
    nor g292 ( n1282 , n98 , n370 );
    nor g293 ( n970 , n2457 , n831 );
    or g294 ( n878 , n1924 , n3604 );
    and g295 ( n1184 , n3086 , n523 );
    or g296 ( n1139 , n1377 , n1529 );
    or g297 ( n834 , n1905 , n2676 );
    nor g298 ( n3401 , n2236 , n491 );
    not g299 ( n1010 , n832 );
    not g300 ( n982 , n3460 );
    not g301 ( n893 , n2651 );
    or g302 ( n1461 , n1157 , n1876 );
    or g303 ( n511 , n1994 , n181 );
    and g304 ( n2475 , n2074 , n788 );
    or g305 ( n3582 , n1111 , n2314 );
    not g306 ( n2524 , n3918 );
    nor g307 ( n194 , n3847 , n494 );
    or g308 ( n1264 , n3380 , n816 );
    or g309 ( n3187 , n1728 , n3910 );
    not g310 ( n1597 , n3344 );
    and g311 ( n3864 , n2631 , n469 );
    nor g312 ( n1076 , n2437 , n643 );
    not g313 ( n3539 , n3220 );
    not g314 ( n3684 , n2875 );
    or g315 ( n1016 , n1488 , n2522 );
    and g316 ( n3361 , n1441 , n1430 );
    and g317 ( n2354 , n1750 , n1963 );
    or g318 ( n697 , n149 , n3903 );
    or g319 ( n529 , n1229 , n3491 );
    and g320 ( n2380 , n2280 , n3571 );
    or g321 ( n1262 , n2712 , n3482 );
    and g322 ( n2300 , n3653 , n3735 );
    or g323 ( n3086 , n409 , n249 );
    not g324 ( n3803 , n2448 );
    and g325 ( n1586 , n3010 , n2828 );
    nor g326 ( n766 , n1250 , n3389 );
    or g327 ( n3259 , n617 , n3742 );
    and g328 ( n1599 , n3800 , n2067 );
    not g329 ( n3400 , n3181 );
    or g330 ( n3656 , n398 , n32 );
    and g331 ( n981 , n145 , n1683 );
    not g332 ( n909 , n1686 );
    nor g333 ( n3837 , n473 , n281 );
    or g334 ( n313 , n900 , n549 );
    not g335 ( n1775 , n2705 );
    and g336 ( n2711 , n2384 , n2547 );
    or g337 ( n56 , n555 , n2800 );
    not g338 ( n1265 , n178 );
    and g339 ( n2333 , n3498 , n310 );
    and g340 ( n2710 , n1030 , n248 );
    or g341 ( n1696 , n2369 , n1509 );
    and g342 ( n542 , n238 , n1873 );
    and g343 ( n1915 , n650 , n1211 );
    and g344 ( n3105 , n3483 , n848 );
    and g345 ( n3061 , n1851 , n1402 );
    and g346 ( n2279 , n510 , n3051 );
    and g347 ( n2676 , n3316 , n3462 );
    or g348 ( n2347 , n1102 , n3103 );
    and g349 ( n2858 , n3125 , n1634 );
    or g350 ( n972 , n1668 , n3795 );
    and g351 ( n1645 , n2423 , n3106 );
    and g352 ( n2741 , n482 , n976 );
    nor g353 ( n3620 , n339 , n3306 );
    and g354 ( n577 , n1996 , n2128 );
    not g355 ( n2713 , n351 );
    not g356 ( n2485 , n2946 );
    and g357 ( n339 , n363 , n1412 );
    nor g358 ( n1633 , n1280 , n1588 );
    or g359 ( n1522 , n1352 , n237 );
    or g360 ( n1973 , n1901 , n2082 );
    not g361 ( n3142 , n2616 );
    and g362 ( n2670 , n3510 , n3329 );
    nor g363 ( n2355 , n395 , n2158 );
    nor g364 ( n3412 , n645 , n600 );
    and g365 ( n707 , n2285 , n415 );
    or g366 ( n1613 , n3739 , n312 );
    nor g367 ( n1099 , n16 , n130 );
    nor g368 ( n794 , n2380 , n190 );
    and g369 ( n3462 , n2277 , n771 );
    or g370 ( n682 , n520 , n795 );
    or g371 ( n1732 , n2954 , n2256 );
    and g372 ( n2821 , n1465 , n1672 );
    or g373 ( n3349 , n572 , n244 );
    buf g374 ( n831 , n2607 );
    and g375 ( n3302 , n620 , n2083 );
    and g376 ( n3918 , n1476 , n3337 );
    or g377 ( n2861 , n1662 , n138 );
    and g378 ( n930 , n1702 , n1688 );
    nor g379 ( n1077 , n3367 , n1359 );
    or g380 ( n958 , n158 , n3695 );
    or g381 ( n3313 , n2644 , n908 );
    nor g382 ( n2842 , n497 , n246 );
    or g383 ( n1632 , n2562 , n1120 );
    not g384 ( n2903 , n3836 );
    or g385 ( n3763 , n241 , n1678 );
    nor g386 ( n371 , n2102 , n2607 );
    not g387 ( n2836 , n1390 );
    or g388 ( n3074 , n2445 , n3692 );
    nor g389 ( n1453 , n2044 , n2754 );
    or g390 ( n734 , n2729 , n2818 );
    not g391 ( n2502 , n712 );
    or g392 ( n3174 , n1704 , n2198 );
    nor g393 ( n3771 , n2780 , n867 );
    and g394 ( n1032 , n2441 , n1940 );
    nor g395 ( n2489 , n2142 , n1117 );
    not g396 ( n3853 , n3379 );
    or g397 ( n3289 , n3229 , n209 );
    and g398 ( n1364 , n1824 , n3617 );
    and g399 ( n1612 , n2008 , n625 );
    and g400 ( n662 , n3417 , n3376 );
    not g401 ( n3374 , n1341 );
    and g402 ( n3661 , n2398 , n1339 );
    or g403 ( n565 , n1366 , n2712 );
    nor g404 ( n2804 , n3651 , n2555 );
    and g405 ( n435 , n2288 , n3519 );
    nor g406 ( n1564 , n3393 , n3683 );
    or g407 ( n1034 , n3137 , n2027 );
    nor g408 ( n1900 , n101 , n868 );
    not g409 ( n3760 , n597 );
    nor g410 ( n2373 , n3035 , n2179 );
    not g411 ( n356 , n1708 );
    and g412 ( n1390 , n1025 , n3177 );
    nor g413 ( n514 , n1274 , n1828 );
    nor g414 ( n1132 , n3768 , n187 );
    nor g415 ( n1671 , n1813 , n111 );
    and g416 ( n1397 , n1556 , n2510 );
    or g417 ( n1238 , n1776 , n2837 );
    or g418 ( n3797 , n2773 , n291 );
    or g419 ( n2620 , n3679 , n874 );
    or g420 ( n246 , n2681 , n3661 );
    and g421 ( n1656 , n2178 , n1724 );
    or g422 ( n1866 , n789 , n1101 );
    and g423 ( n2115 , n1245 , n1085 );
    nor g424 ( n1221 , n73 , n1197 );
    or g425 ( n640 , n3 , n761 );
    and g426 ( n3346 , n901 , n1110 );
    or g427 ( n2693 , n1501 , n2265 );
    and g428 ( n3889 , n2127 , n3752 );
    not g429 ( n238 , n3236 );
    or g430 ( n326 , n1160 , n1448 );
    or g431 ( n1628 , n1436 , n3302 );
    not g432 ( n2493 , n1387 );
    not g433 ( n3179 , n1341 );
    and g434 ( n661 , n3662 , n3067 );
    nor g435 ( n2667 , n593 , n506 );
    not g436 ( n2548 , n1314 );
    nor g437 ( n1911 , n3606 , n2317 );
    nor g438 ( n2474 , n2191 , n480 );
    and g439 ( n3326 , n518 , n1428 );
    or g440 ( n3901 , n970 , n1564 );
    and g441 ( n1318 , n3833 , n1734 );
    or g442 ( n1634 , n1309 , n3692 );
    not g443 ( n596 , n1287 );
    or g444 ( n2339 , n243 , n3275 );
    or g445 ( n2023 , n3401 , n231 );
    or g446 ( n1378 , n966 , n715 );
    or g447 ( n391 , n2467 , n1898 );
    and g448 ( n3817 , n787 , n104 );
    not g449 ( n144 , n695 );
    and g450 ( n1739 , n2028 , n247 );
    not g451 ( n3158 , n676 );
    or g452 ( n2231 , n3373 , n1916 );
    not g453 ( n2217 , n264 );
    nor g454 ( n980 , n2107 , n904 );
    or g455 ( n383 , n3117 , n384 );
    nor g456 ( n3451 , n1408 , n2948 );
    nor g457 ( n93 , n3504 , n2551 );
    or g458 ( n1621 , n3307 , n1857 );
    or g459 ( n951 , n1219 , n1382 );
    or g460 ( n534 , n3063 , n827 );
    nor g461 ( n2131 , n948 , n3546 );
    not g462 ( n2970 , n923 );
    and g463 ( n22 , n2406 , n567 );
    not g464 ( n1640 , n1729 );
    nor g465 ( n2642 , n2985 , n596 );
    or g466 ( n2894 , n2662 , n1447 );
    and g467 ( n3854 , n2988 , n2973 );
    and g468 ( n1432 , n2324 , n3295 );
    not g469 ( n3698 , n497 );
    or g470 ( n3341 , n2150 , n5 );
    or g471 ( n2942 , n117 , n893 );
    nor g472 ( n3389 , n257 , n3879 );
    not g473 ( n594 , n984 );
    nor g474 ( n2399 , n2023 , n1142 );
    or g475 ( n35 , n2660 , n2733 );
    not g476 ( n2600 , n2995 );
    and g477 ( n3524 , n1923 , n1407 );
    nor g478 ( n1239 , n3480 , n3319 );
    not g479 ( n2177 , n3744 );
    or g480 ( n2392 , n2051 , n3449 );
    not g481 ( n836 , n1983 );
    and g482 ( n2076 , n3636 , n2037 );
    not g483 ( n2337 , n2371 );
    and g484 ( n1686 , n3386 , n332 );
    nor g485 ( n2972 , n680 , n205 );
    not g486 ( n2956 , n3379 );
    or g487 ( n2274 , n1061 , n1188 );
    and g488 ( n776 , n933 , n804 );
    not g489 ( n2951 , n1341 );
    nor g490 ( n1887 , n578 , n1109 );
    and g491 ( n2602 , n1893 , n1125 );
    and g492 ( n1357 , n835 , n830 );
    not g493 ( n3479 , n3512 );
    and g494 ( n3561 , n448 , n2816 );
    and g495 ( n3081 , n65 , n1008 );
    and g496 ( n452 , n3483 , n2332 );
    not g497 ( n3092 , n3387 );
    and g498 ( n1228 , n186 , n1611 );
    and g499 ( n3023 , n1684 , n1271 );
    or g500 ( n668 , n2699 , n1930 );
    or g501 ( n910 , n810 , n1188 );
    or g502 ( n3688 , n709 , n2996 );
    or g503 ( n2822 , n1794 , n3903 );
    or g504 ( n506 , n1234 , n700 );
    not g505 ( n1433 , n2482 );
    and g506 ( n3767 , n2625 , n1707 );
    or g507 ( n504 , n2287 , n2989 );
    not g508 ( n3288 , n2946 );
    or g509 ( n3572 , n1186 , n826 );
    not g510 ( n3352 , n2984 );
    nor g511 ( n1141 , n274 , n1726 );
    and g512 ( n1354 , n3451 , n2751 );
    or g513 ( n2905 , n2760 , n1283 );
    or g514 ( n2755 , n1836 , n914 );
    nor g515 ( n3916 , n1202 , n3445 );
    or g516 ( n3723 , n2848 , n509 );
    and g517 ( n2164 , n454 , n1285 );
    nor g518 ( n2757 , n1641 , n1728 );
    or g519 ( n2214 , n507 , n908 );
    or g520 ( n704 , n1049 , n3232 );
    nor g521 ( n1469 , n1236 , n166 );
    and g522 ( n2142 , n2330 , n3869 );
    or g523 ( n3635 , n403 , n3573 );
    not g524 ( n850 , n2788 );
    nor g525 ( n1111 , n810 , n2891 );
    nor g526 ( n2501 , n1531 , n919 );
    or g527 ( n1511 , n1938 , n3449 );
    and g528 ( n564 , n3816 , n1369 );
    or g529 ( n2383 , n1798 , n1097 );
    and g530 ( n3304 , n74 , n1872 );
    or g531 ( n2160 , n608 , n1473 );
    not g532 ( n62 , n3379 );
    and g533 ( n3586 , n2769 , n1364 );
    and g534 ( n1154 , n2544 , n470 );
    not g535 ( n3298 , n3469 );
    not g536 ( n3079 , n133 );
    or g537 ( n3342 , n2691 , n2855 );
    and g538 ( n425 , n2879 , n2519 );
    not g539 ( n2565 , n1360 );
    and g540 ( n3790 , n1041 , n3644 );
    nor g541 ( n1429 , n438 , n3133 );
    nor g542 ( n1856 , n3675 , n993 );
    and g543 ( n1190 , n937 , n3088 );
    nor g544 ( n2866 , n670 , n2258 );
    nor g545 ( n2045 , n3004 , n203 );
    nor g546 ( n442 , n3151 , n2572 );
    or g547 ( n901 , n2254 , n3257 );
    or g548 ( n3347 , n3608 , n2939 );
    or g549 ( n2083 , n2443 , n3142 );
    or g550 ( n1237 , n2149 , n3887 );
    not g551 ( n2556 , n691 );
    nor g552 ( n862 , n3398 , n2399 );
    and g553 ( n2253 , n2846 , n1522 );
    or g554 ( n3824 , n2685 , n571 );
    nor g555 ( n2808 , n1098 , n959 );
    or g556 ( n540 , n1757 , n3903 );
    and g557 ( n2960 , n3114 , n789 );
    and g558 ( n1681 , n3851 , n3774 );
    and g559 ( n864 , n1763 , n2519 );
    not g560 ( n882 , n1332 );
    or g561 ( n2453 , n3220 , n3887 );
    nor g562 ( n1126 , n3631 , n2084 );
    and g563 ( n779 , n2625 , n1517 );
    not g564 ( n3231 , n580 );
    or g565 ( n388 , n2616 , n3692 );
    and g566 ( n3324 , n2268 , n669 );
    nor g567 ( n544 , n2467 , n819 );
    not g568 ( n3536 , n2195 );
    nor g569 ( n461 , n2333 , n3298 );
    nor g570 ( n2535 , n2289 , n439 );
    not g571 ( n1647 , n1958 );
    nor g572 ( n1890 , n1592 , n3425 );
    or g573 ( n822 , n1890 , n2943 );
    or g574 ( n3077 , n1808 , n992 );
    or g575 ( n1244 , n3787 , n1101 );
    not g576 ( n1128 , n2031 );
    and g577 ( n1801 , n1074 , n3441 );
    and g578 ( n3832 , n312 , n3739 );
    or g579 ( n874 , n2626 , n2807 );
    not g580 ( n430 , n2946 );
    and g581 ( n493 , n562 , n629 );
    not g582 ( n2481 , n2639 );
    not g583 ( n2022 , n139 );
    or g584 ( n154 , n3227 , n908 );
    and g585 ( n1123 , n3758 , n1128 );
    or g586 ( n1215 , n971 , n3262 );
    nor g587 ( n1918 , n1765 , n2397 );
    or g588 ( n751 , n1689 , n306 );
    and g589 ( n3610 , n2109 , n1150 );
    nor g590 ( n2088 , n3643 , n1324 );
    and g591 ( n3319 , n1468 , n2829 );
    or g592 ( n1996 , n3160 , n1832 );
    not g593 ( n3773 , n2919 );
    nor g594 ( n1484 , n622 , n1667 );
    and g595 ( n3330 , n1796 , n1831 );
    and g596 ( n2107 , n3075 , n1569 );
    and g597 ( n1373 , n3801 , n734 );
    and g598 ( n623 , n733 , n1960 );
    and g599 ( n2114 , n989 , n71 );
    nor g600 ( n1950 , n2196 , n3503 );
    not g601 ( n3777 , n705 );
    nor g602 ( n3537 , n1441 , n1384 );
    not g603 ( n2331 , n2463 );
    and g604 ( n3630 , n2625 , n2723 );
    and g605 ( n591 , n3687 , n2722 );
    nor g606 ( n2278 , n1038 , n2539 );
    not g607 ( n867 , n637 );
    or g608 ( n1035 , n2545 , n591 );
    or g609 ( n814 , n576 , n1187 );
    and g610 ( n1627 , n1001 , n3824 );
    and g611 ( n3895 , n2779 , n540 );
    not g612 ( n1816 , n2946 );
    not g613 ( n3099 , n2336 );
    not g614 ( n3785 , n2933 );
    nor g615 ( n393 , n28 , n1072 );
    nor g616 ( n3241 , n2925 , n2607 );
    and g617 ( n800 , n1962 , n473 );
    nor g618 ( n3784 , n3312 , n860 );
    and g619 ( n1930 , n2793 , n3852 );
    or g620 ( n2811 , n615 , n3324 );
    and g621 ( n1319 , n9 , n2356 );
    nor g622 ( n2044 , n3681 , n1939 );
    not g623 ( n1849 , n2520 );
    not g624 ( n2665 , n2946 );
    and g625 ( n916 , n3774 , n1611 );
    and g626 ( n1858 , n961 , n364 );
    nor g627 ( n1465 , n2308 , n393 );
    nor g628 ( n3049 , n774 , n849 );
    not g629 ( n3083 , n1754 );
    nor g630 ( n2690 , n3028 , n3470 );
    nor g631 ( n659 , n3856 , n610 );
    and g632 ( n1160 , n437 , n707 );
    not g633 ( n2596 , n1966 );
    or g634 ( n484 , n1152 , n2164 );
    and g635 ( n1387 , n2776 , n2557 );
    and g636 ( n355 , n3091 , n2537 );
    and g637 ( n3640 , n1983 , n2861 );
    nor g638 ( n700 , n872 , n3172 );
    and g639 ( n2408 , n3375 , n383 );
    or g640 ( n817 , n774 , n1898 );
    or g641 ( n1936 , n26 , n3513 );
    not g642 ( n2806 , n1892 );
    and g643 ( n1368 , n2608 , n1585 );
    nor g644 ( n2242 , n117 , n1566 );
    and g645 ( n3585 , n3156 , n3343 );
    not g646 ( n491 , n3897 );
    or g647 ( n2404 , n1144 , n893 );
    or g648 ( n1271 , n2459 , n3692 );
    nor g649 ( n2068 , n2734 , n558 );
    and g650 ( n2797 , n259 , n1090 );
    not g651 ( n1037 , n3426 );
    nor g652 ( n2655 , n1091 , n2306 );
    nor g653 ( n3595 , n1774 , n2944 );
    nor g654 ( n1218 , n3360 , n2769 );
    nor g655 ( n230 , n1530 , n2474 );
    not g656 ( n3033 , n3624 );
    not g657 ( n792 , n945 );
    nor g658 ( n1785 , n1971 , n808 );
    not g659 ( n1574 , n718 );
    and g660 ( n1071 , n3515 , n315 );
    nor g661 ( n2471 , n1900 , n3465 );
    nor g662 ( n767 , n1411 , n3244 );
    nor g663 ( n1065 , n85 , n2485 );
    and g664 ( n3724 , n545 , n1897 );
    and g665 ( n1623 , n251 , n1886 );
    and g666 ( n1676 , n1993 , n2431 );
    and g667 ( n61 , n1729 , n525 );
    or g668 ( n350 , n1491 , n3466 );
    or g669 ( n3496 , n1135 , n981 );
    not g670 ( n496 , n2946 );
    or g671 ( n3805 , n233 , n222 );
    and g672 ( n2666 , n2976 , n63 );
    and g673 ( n830 , n2635 , n744 );
    nor g674 ( n2438 , n1579 , n3612 );
    and g675 ( n1008 , n350 , n1519 );
    nor g676 ( n942 , n3790 , n1348 );
    nor g677 ( n2158 , n2646 , n1950 );
    or g678 ( n3031 , n658 , n2904 );
    not g679 ( n2898 , n3379 );
    or g680 ( n2205 , n1199 , n876 );
    and g681 ( n1899 , n122 , n3722 );
    or g682 ( n1787 , n3509 , n1141 );
    buf g683 ( n908 , n3887 );
    or g684 ( n3526 , n2243 , n2701 );
    and g685 ( n3041 , n3250 , n3914 );
    or g686 ( n2324 , n2933 , n1916 );
    or g687 ( n2517 , n3528 , n1188 );
    nor g688 ( n1956 , n2063 , n862 );
    or g689 ( n28 , n1420 , n3363 );
    or g690 ( n741 , n3614 , n2996 );
    and g691 ( n1497 , n973 , n2762 );
    and g692 ( n3294 , n3520 , n3905 );
    or g693 ( n742 , n2431 , n3742 );
    and g694 ( n1279 , n1949 , n2038 );
    or g695 ( n2462 , n1997 , n2497 );
    not g696 ( n1296 , n1593 );
    not g697 ( n1331 , n3349 );
    and g698 ( n826 , n275 , n2068 );
    and g699 ( n3573 , n814 , n1064 );
    and g700 ( n46 , n2720 , n832 );
    nor g701 ( n768 , n3468 , n944 );
    not g702 ( n3328 , n2658 );
    not g703 ( n2653 , n2648 );
    not g704 ( n3403 , n2910 );
    not g705 ( n3900 , n3887 );
    nor g706 ( n1482 , n3177 , n1025 );
    and g707 ( n2619 , n1860 , n455 );
    and g708 ( n998 , n759 , n2694 );
    or g709 ( n610 , n1069 , n3760 );
    nor g710 ( n2209 , n216 , n2641 );
    or g711 ( n1587 , n242 , n85 );
    or g712 ( n2040 , n1548 , n509 );
    nor g713 ( n685 , n1151 , n2747 );
    and g714 ( n220 , n3694 , n329 );
    nor g715 ( n3167 , n2669 , n382 );
    or g716 ( n2464 , n3159 , n632 );
    and g717 ( n1109 , n3133 , n438 );
    or g718 ( n3228 , n1287 , n1916 );
    or g719 ( n1080 , n2960 , n451 );
    not g720 ( n1843 , n1612 );
    or g721 ( n3038 , n1482 , n714 );
    or g722 ( n2724 , n858 , n295 );
    nor g723 ( n2505 , n401 , n3045 );
    nor g724 ( n3876 , n569 , n2181 );
    and g725 ( n3847 , n1574 , n379 );
    and g726 ( n3494 , n2625 , n264 );
    not g727 ( n3404 , n467 );
    not g728 ( n1808 , n2968 );
    and g729 ( n3843 , n278 , n738 );
    or g730 ( n1791 , n1915 , n341 );
    and g731 ( n3197 , n2980 , n2656 );
    or g732 ( n2304 , n898 , n2434 );
    or g733 ( n2742 , n282 , n761 );
    or g734 ( n283 , n1690 , n3746 );
    and g735 ( n1362 , n3357 , n3808 );
    not g736 ( n3689 , n1100 );
    not g737 ( n3566 , n2439 );
    or g738 ( n1869 , n3676 , n1005 );
    nor g739 ( n3702 , n2111 , n467 );
    not g740 ( n1734 , n2111 );
    nor g741 ( n2599 , n2617 , n3407 );
    or g742 ( n1302 , n957 , n642 );
    not g743 ( n2860 , n3887 );
    or g744 ( n1565 , n2211 , n3692 );
    nor g745 ( n59 , n3282 , n3418 );
    or g746 ( n1923 , n3190 , n2182 );
    and g747 ( n2412 , n437 , n3095 );
    or g748 ( n3076 , n226 , n1207 );
    or g749 ( n1534 , n3441 , n3887 );
    nor g750 ( n2914 , n1837 , n3535 );
    or g751 ( n1967 , n321 , n761 );
    or g752 ( n1541 , n2991 , n1188 );
    nor g753 ( n1383 , n3833 , n1716 );
    or g754 ( n3078 , n842 , n2996 );
    or g755 ( n1987 , n1392 , n1456 );
    and g756 ( n3518 , n234 , n1205 );
    and g757 ( n1582 , n3526 , n2259 );
    and g758 ( n2456 , n1910 , n2130 );
    or g759 ( n625 , n1533 , n2162 );
    or g760 ( n2890 , n1395 , n3015 );
    nor g761 ( n1017 , n2384 , n3046 );
    and g762 ( n693 , n910 , n939 );
    and g763 ( n3504 , n2814 , n2069 );
    nor g764 ( n3904 , n1368 , n1918 );
    or g765 ( n1205 , n2463 , n761 );
    not g766 ( n3721 , n1341 );
    not g767 ( n3186 , n2166 );
    not g768 ( n2864 , n1013 );
    or g769 ( n2796 , n3427 , n2607 );
    or g770 ( n3210 , n3411 , n1362 );
    and g771 ( n3839 , n2247 , n3728 );
    or g772 ( n3765 , n3881 , n2410 );
    or g773 ( n815 , n371 , n956 );
    and g774 ( n3862 , n3076 , n2047 );
    and g775 ( n2987 , n1572 , n2862 );
    and g776 ( n2499 , n346 , n2079 );
    and g777 ( n1194 , n1089 , n2460 );
    nor g778 ( n426 , n2529 , n2765 );
    nor g779 ( n381 , n144 , n254 );
    and g780 ( n3616 , n36 , n2762 );
    and g781 ( n2055 , n1987 , n3270 );
    not g782 ( n2360 , n1341 );
    and g783 ( n615 , n2268 , n1338 );
    nor g784 ( n2175 , n3912 , n3765 );
    not g785 ( n3178 , n3063 );
    not g786 ( n1960 , n3476 );
    not g787 ( n44 , n2774 );
    nor g788 ( n3300 , n3710 , n1164 );
    or g789 ( n1710 , n2425 , n1455 );
    nor g790 ( n1206 , n1061 , n2806 );
    or g791 ( n2226 , n1130 , n2607 );
    and g792 ( n424 , n1893 , n2853 );
    or g793 ( n1990 , n407 , n3667 );
    not g794 ( n433 , n1661 );
    or g795 ( n3502 , n1544 , n2607 );
    or g796 ( n3182 , n3390 , n3910 );
    and g797 ( n269 , n2625 , n1618 );
    or g798 ( n114 , n2570 , n2541 );
    and g799 ( n1754 , n1323 , n677 );
    and g800 ( n3168 , n433 , n2955 );
    or g801 ( n849 , n1753 , n3732 );
    or g802 ( n1486 , n1778 , n1898 );
    nor g803 ( n111 , n42 , n146 );
    or g804 ( n52 , n3211 , n1333 );
    and g805 ( n1867 , n3021 , n1304 );
    or g806 ( n1110 , n2738 , n11 );
    and g807 ( n3919 , n1711 , n1780 );
    and g808 ( n922 , n1035 , n1732 );
    and g809 ( n169 , n177 , n2049 );
    or g810 ( n1301 , n255 , n1042 );
    or g811 ( n3431 , n2335 , n2411 );
    and g812 ( n211 , n3266 , n3476 );
    nor g813 ( n204 , n1779 , n3161 );
    not g814 ( n3318 , n3593 );
    or g815 ( n2272 , n152 , n1445 );
    or g816 ( n2478 , n3034 , n1929 );
    and g817 ( n1606 , n639 , n2037 );
    nor g818 ( n267 , n2300 , n2735 );
    and g819 ( n1416 , n719 , n964 );
    nor g820 ( n2168 , n1182 , n3725 );
    and g821 ( n3008 , n3483 , n1773 );
    and g822 ( n1832 , n1628 , n3347 );
    not g823 ( n1730 , n2946 );
    and g824 ( n2183 , n1759 , n1506 );
    not g825 ( n3516 , n3817 );
    and g826 ( n215 , n3483 , n1167 );
    not g827 ( n403 , n233 );
    and g828 ( n648 , n903 , n1849 );
    not g829 ( n545 , n519 );
    not g830 ( n1670 , n2498 );
    nor g831 ( n1018 , n2998 , n3482 );
    or g832 ( n2433 , n462 , n1101 );
    nor g833 ( n19 , n3856 , n831 );
    or g834 ( n1103 , n2655 , n3558 );
    or g835 ( n3714 , n2242 , n1020 );
    nor g836 ( n129 , n2052 , n1878 );
    nor g837 ( n2847 , n1083 , n2192 );
    or g838 ( n2005 , n2266 , n761 );
    nor g839 ( n1406 , n3571 , n831 );
    not g840 ( n3455 , n2469 );
    not g841 ( n600 , n2946 );
    or g842 ( n281 , n1962 , n2579 );
    not g843 ( n277 , n3 );
    and g844 ( n729 , n2990 , n472 );
    nor g845 ( n2125 , n1942 , n1337 );
    or g846 ( n3017 , n986 , n3853 );
    not g847 ( n2542 , n2439 );
    and g848 ( n2669 , n2944 , n1774 );
    nor g849 ( n2085 , n2552 , n1440 );
    or g850 ( n1504 , n2310 , n1594 );
    or g851 ( n1096 , n3372 , n80 );
    or g852 ( n2028 , n426 , n2746 );
    or g853 ( n3691 , n1755 , n894 );
    or g854 ( n1291 , n1999 , n1322 );
    nor g855 ( n1455 , n459 , n2160 );
    and g856 ( n1738 , n2769 , n2306 );
    and g857 ( n2434 , n2665 , n1255 );
    nor g858 ( n3866 , n3814 , n1512 );
    and g859 ( n218 , n1828 , n1274 );
    and g860 ( n3405 , n2625 , n2461 );
    or g861 ( n557 , n3809 , n3650 );
    not g862 ( n3506 , n2364 );
    not g863 ( n1761 , n2103 );
    nor g864 ( n3467 , n1721 , n551 );
    or g865 ( n2163 , n2498 , n3887 );
    or g866 ( n2621 , n3885 , n908 );
    not g867 ( n3546 , n568 );
    not g868 ( n2793 , n912 );
    not g869 ( n3345 , n3379 );
    not g870 ( n1197 , n2731 );
    or g871 ( n3532 , n526 , n3053 );
    not g872 ( n311 , n3107 );
    and g873 ( n1707 , n3044 , n2404 );
    and g874 ( n1914 , n188 , n3859 );
    not g875 ( n2152 , n1051 );
    nor g876 ( n1234 , n3273 , n3714 );
    not g877 ( n3043 , n3380 );
    nor g878 ( n3730 , n462 , n2827 );
    or g879 ( n2007 , n3248 , n1740 );
    or g880 ( n3602 , n1429 , n3864 );
    and g881 ( n2736 , n3841 , n1004 );
    not g882 ( n827 , n3658 );
    or g883 ( n3151 , n2175 , n1217 );
    and g884 ( n134 , n430 , n1789 );
    or g885 ( n976 , n3747 , n3202 );
    or g886 ( n474 , n3830 , n2484 );
    nor g887 ( n3559 , n588 , n129 );
    buf g888 ( n1277 , n1143 );
    and g889 ( n119 , n39 , n3643 );
    and g890 ( n1917 , n792 , n3279 );
    or g891 ( n936 , n3390 , n2017 );
    and g892 ( n2691 , n1373 , n732 );
    and g893 ( n572 , n761 , n379 );
    or g894 ( n358 , n949 , n3015 );
    or g895 ( n1343 , n164 , n1073 );
    or g896 ( n1292 , n2512 , n859 );
    nor g897 ( n3368 , n1104 , n2568 );
    nor g898 ( n1002 , n398 , n1257 );
    and g899 ( n143 , n3765 , n537 );
    or g900 ( n2678 , n1880 , n2996 );
    nor g901 ( n3740 , n227 , n3597 );
    buf g902 ( n1893 , n2769 );
    not g903 ( n3612 , n2946 );
    not g904 ( n612 , n3137 );
    or g905 ( n1500 , n1418 , n2716 );
    not g906 ( n1143 , n1701 );
    or g907 ( n3680 , n1629 , n3692 );
    or g908 ( n1324 , n39 , n3275 );
    and g909 ( n2386 , n3483 , n1686 );
    not g910 ( n279 , n3310 );
    or g911 ( n2966 , n2477 , n571 );
    or g912 ( n677 , n3430 , n3047 );
    not g913 ( n1045 , n2215 );
    or g914 ( n193 , n2183 , n2640 );
    and g915 ( n1793 , n437 , n1435 );
    and g916 ( n1603 , n2162 , n1533 );
    not g917 ( n777 , n3296 );
    or g918 ( n399 , n2412 , n3913 );
    not g919 ( n1489 , n1397 );
    not g920 ( n2351 , n2266 );
    or g921 ( n537 , n3912 , n2410 );
    and g922 ( n1965 , n2586 , n2381 );
    nor g923 ( n1764 , n3207 , n1003 );
    and g924 ( n1350 , n1074 , n2073 );
    or g925 ( n2427 , n3621 , n369 );
    and g926 ( n2538 , n1304 , n2248 );
    not g927 ( n2000 , n17 );
    not g928 ( n276 , n1431 );
    or g929 ( n3589 , n492 , n1898 );
    or g930 ( n330 , n3704 , n3105 );
    and g931 ( n1480 , n2624 , n711 );
    nor g932 ( n1543 , n1585 , n2810 );
    and g933 ( n2762 , n554 , n1516 );
    and g934 ( n679 , n3639 , n3601 );
    and g935 ( n2791 , n437 , n527 );
    or g936 ( n3823 , n1662 , n761 );
    or g937 ( n3663 , n1819 , n68 );
    or g938 ( n298 , n3831 , n3655 );
    and g939 ( n2978 , n2464 , n3086 );
    nor g940 ( n1040 , n284 , n563 );
    and g941 ( n1075 , n481 , n2013 );
    and g942 ( n208 , n955 , n3705 );
    or g943 ( n82 , n1398 , n344 );
    or g944 ( n1588 , n2097 , n577 );
    and g945 ( n1263 , n3879 , n257 );
    and g946 ( n2275 , n3660 , n1991 );
    and g947 ( n341 , n1043 , n2312 );
    buf g948 ( n3548 , n1701 );
    or g949 ( n3472 , n1944 , n3015 );
    not g950 ( n2141 , n3061 );
    and g951 ( n3185 , n2391 , n999 );
    nor g952 ( n1093 , n1743 , n406 );
    and g953 ( n717 , n3209 , n2326 );
    or g954 ( n1740 , n3564 , n2882 );
    nor g955 ( n2585 , n218 , n3821 );
    or g956 ( n1299 , n2443 , n3466 );
    not g957 ( n32 , n2906 );
    or g958 ( n1138 , n675 , n1207 );
    or g959 ( n2260 , n46 , n1645 );
    not g960 ( n1868 , n152 );
    and g961 ( n2748 , n1546 , n2656 );
    nor g962 ( n1326 , n2491 , n3703 );
    or g963 ( n89 , n2985 , n302 );
    not g964 ( n2136 , n2176 );
    and g965 ( n16 , n55 , n127 );
    or g966 ( n2884 , n1998 , n1623 );
    or g967 ( n2766 , n3085 , n1749 );
    nor g968 ( n3377 , n829 , n40 );
    or g969 ( n198 , n2853 , n90 );
    not g970 ( n2293 , n1418 );
    and g971 ( n3333 , n1596 , n2483 );
    not g972 ( n1716 , n299 );
    or g973 ( n3088 , n641 , n3573 );
    nor g974 ( n449 , n3330 , n3559 );
    nor g975 ( n128 , n3261 , n1775 );
    nor g976 ( n14 , n777 , n3576 );
    not g977 ( n1243 , n1265 );
    or g978 ( n1845 , n3693 , n1916 );
    not g979 ( n3475 , n1283 );
    or g980 ( n587 , n1059 , n288 );
    or g981 ( n2270 , n1934 , n876 );
    and g982 ( n2432 , n3231 , n3434 );
    or g983 ( n3100 , n325 , n3099 );
    or g984 ( n1643 , n2479 , n831 );
    not g985 ( n2760 , n2945 );
    and g986 ( n1196 , n3025 , n3726 );
    and g987 ( n2064 , n736 , n1609 );
    nor g988 ( n2732 , n1009 , n123 );
    or g989 ( n253 , n1255 , n3265 );
    or g990 ( n3238 , n2711 , n883 );
    nor g991 ( n3541 , n899 , n1921 );
    and g992 ( n2928 , n995 , n2813 );
    not g993 ( n1881 , n164 );
    not g994 ( n3196 , n2946 );
    or g995 ( n896 , n489 , n143 );
    and g996 ( n3538 , n817 , n2621 );
    and g997 ( n2692 , n412 , n2520 );
    and g998 ( n551 , n476 , n2480 );
    or g999 ( n3545 , n944 , n3709 );
    or g1000 ( n466 , n101 , n1188 );
    nor g1001 ( n3557 , n2685 , n2530 );
    and g1002 ( n2680 , n2625 , n1675 );
    nor g1003 ( n2377 , n1021 , n3508 );
    not g1004 ( n196 , n2475 );
    nor g1005 ( n2081 , n2123 , n2126 );
    and g1006 ( n603 , n217 , n3538 );
    or g1007 ( n3072 , n954 , n3449 );
    and g1008 ( n764 , n2994 , n2638 );
    or g1009 ( n1241 , n3024 , n97 );
    nor g1010 ( n1442 , n1676 , n1920 );
    and g1011 ( n2184 , n716 , n2568 );
    nor g1012 ( n1853 , n960 , n968 );
    or g1013 ( n3489 , n2353 , n2996 );
    not g1014 ( n2336 , n3345 );
    and g1015 ( n3544 , n1781 , n3213 );
    nor g1016 ( n1817 , n2720 , n1750 );
    and g1017 ( n1408 , n968 , n960 );
    or g1018 ( n1232 , n19 , n1911 );
    and g1019 ( n2832 , n1643 , n1550 );
    not g1020 ( n2216 , n103 );
    and g1021 ( n2492 , n1998 , n263 );
    or g1022 ( n3398 , n499 , n2020 );
    or g1023 ( n441 , n2220 , n1159 );
    not g1024 ( n2317 , n3379 );
    and g1025 ( n1415 , n713 , n2332 );
    or g1026 ( n3007 , n1731 , n1916 );
    and g1027 ( n2307 , n1939 , n240 );
    and g1028 ( n923 , n2679 , n3793 );
    and g1029 ( n1322 , n1595 , n3848 );
    and g1030 ( n569 , n3019 , n3056 );
    or g1031 ( n120 , n943 , n624 );
    or g1032 ( n927 , n845 , n1112 );
    or g1033 ( n2958 , n3549 , n2715 );
    nor g1034 ( n1650 , n1525 , n1284 );
    not g1035 ( n186 , n1341 );
    and g1036 ( n3436 , n1373 , n756 );
    or g1037 ( n1149 , n1861 , n1898 );
    not g1038 ( n1516 , n2579 );
    not g1039 ( n2034 , n675 );
    or g1040 ( n2633 , n2322 , n1169 );
    not g1041 ( n726 , n3631 );
    and g1042 ( n1713 , n2239 , n697 );
    or g1043 ( n278 , n3137 , n2607 );
    not g1044 ( n1493 , n1582 );
    and g1045 ( n81 , n3166 , n3138 );
    and g1046 ( n2024 , n1119 , n3752 );
    and g1047 ( n1412 , n3332 , n410 );
    and g1048 ( n268 , n3260 , n2111 );
    or g1049 ( n3291 , n3629 , n2763 );
    or g1050 ( n2650 , n3110 , n2553 );
    not g1051 ( n3735 , n1769 );
    and g1052 ( n624 , n1667 , n622 );
    and g1053 ( n2087 , n3381 , n2740 );
    or g1054 ( n3463 , n1287 , n1545 );
    not g1055 ( n1396 , n629 );
    or g1056 ( n2435 , n1140 , n731 );
    nor g1057 ( n1059 , n3843 , n1895 );
    or g1058 ( n126 , n1736 , n3903 );
    and g1059 ( n2647 , n1057 , n3819 );
    or g1060 ( n1391 , n3519 , n2607 );
    and g1061 ( n706 , n3409 , n1092 );
    not g1062 ( n3906 , n299 );
    or g1063 ( n2403 , n2026 , n3742 );
    or g1064 ( n2873 , n1738 , n724 );
    or g1065 ( n728 , n3631 , n1101 );
    and g1066 ( n173 , n1893 , n1043 );
    and g1067 ( n305 , n1388 , n189 );
    or g1068 ( n1951 , n907 , n1351 );
    and g1069 ( n2385 , n2625 , n386 );
    or g1070 ( n53 , n1622 , n2376 );
    nor g1071 ( n967 , n1822 , n2797 );
    not g1072 ( n798 , n3358 );
    nor g1073 ( n3830 , n3471 , n831 );
    and g1074 ( n2880 , n183 , n3895 );
    nor g1075 ( n3827 , n461 , n2349 );
    nor g1076 ( n68 , n3006 , n1893 );
    or g1077 ( n3622 , n1246 , n2824 );
    or g1078 ( n3891 , n1380 , n2114 );
    and g1079 ( n3364 , n437 , n1934 );
    not g1080 ( n2376 , n2538 );
    and g1081 ( n2751 , n3206 , n2758 );
    or g1082 ( n3884 , n3037 , n3425 );
    or g1083 ( n517 , n1966 , n571 );
    or g1084 ( n3503 , n1692 , n2031 );
    nor g1085 ( n2238 , n3544 , n621 );
    and g1086 ( n1777 , n3483 , n1008 );
    nor g1087 ( n1003 , n1532 , n1240 );
    not g1088 ( n613 , n1919 );
    nor g1089 ( n3851 , n649 , n2659 );
    not g1090 ( n1891 , n3682 );
    not g1091 ( n48 , n3547 );
    and g1092 ( n672 , n1608 , n1300 );
    or g1093 ( n2074 , n1944 , n2777 );
    and g1094 ( n45 , n2664 , n1039 );
    not g1095 ( n933 , n2398 );
    or g1096 ( n1617 , n435 , n3776 );
    or g1097 ( n3265 , n2509 , n2952 );
    nor g1098 ( n884 , n2445 , n3062 );
    nor g1099 ( n1539 , n3918 , n2408 );
    or g1100 ( n1310 , n2499 , n2225 );
    and g1101 ( n2382 , n3627 , n3402 );
    and g1102 ( n189 , n2098 , n3823 );
    not g1103 ( n1006 , n2436 );
    not g1104 ( n1929 , n2896 );
    or g1105 ( n992 , n2770 , n1529 );
    nor g1106 ( n5 , n3093 , n1227 );
    or g1107 ( n1912 , n2261 , n2001 );
    and g1108 ( n1690 , n3565 , n720 );
    nor g1109 ( n2394 , n830 , n835 );
    and g1110 ( n1748 , n1621 , n2887 );
    or g1111 ( n1616 , n232 , n1374 );
    or g1112 ( n2799 , n3481 , n2607 );
    nor g1113 ( n1737 , n2487 , n1554 );
    not g1114 ( n1131 , n3366 );
    and g1115 ( n1517 , n3129 , n583 );
    not g1116 ( n1562 , n373 );
    buf g1117 ( n3692 , n761 );
    and g1118 ( n2100 , n1810 , n2366 );
    or g1119 ( n2013 , n1421 , n3457 );
    or g1120 ( n2859 , n1602 , n3751 );
    or g1121 ( n1922 , n3231 , n3737 );
    not g1122 ( n1073 , n1514 );
    and g1123 ( n2519 , n2377 , n2481 );
    not g1124 ( n723 , n2736 );
    and g1125 ( n376 , n959 , n815 );
    nor g1126 ( n74 , n1298 , n918 );
    or g1127 ( n85 , n2294 , n1800 );
    not g1128 ( n2237 , n1114 );
    and g1129 ( n3069 , n1923 , n815 );
    or g1130 ( n175 , n1648 , n1898 );
    not g1131 ( n1169 , n282 );
    or g1132 ( n546 , n1506 , n2860 );
    not g1133 ( n2262 , n949 );
    nor g1134 ( n2357 , n471 , n2875 );
    or g1135 ( n1815 , n392 , n3628 );
    or g1136 ( n1619 , n3439 , n1207 );
    nor g1137 ( n159 , n579 , n1046 );
    or g1138 ( n2401 , n164 , n2607 );
    or g1139 ( n1316 , n1430 , n1441 );
    or g1140 ( n541 , n1842 , n1319 );
    or g1141 ( n2465 , n1580 , n1586 );
    not g1142 ( n2490 , n2473 );
    or g1143 ( n1553 , n285 , n3486 );
    not g1144 ( n1251 , n1852 );
    and g1145 ( n2215 , n1538 , n517 );
    nor g1146 ( n3162 , n1723 , n1675 );
    or g1147 ( n3639 , n2079 , n346 );
    or g1148 ( n243 , n3794 , n119 );
    nor g1149 ( n1659 , n1514 , n1881 );
    or g1150 ( n3136 , n2511 , n184 );
    and g1151 ( n3756 , n3500 , n165 );
    and g1152 ( n1112 , n1254 , n951 );
    not g1153 ( n2188 , n803 );
    or g1154 ( n1684 , n2424 , n509 );
    or g1155 ( n240 , n1693 , n3311 );
    and g1156 ( n525 , n2877 , n1967 );
    or g1157 ( n3761 , n606 , n1154 );
    nor g1158 ( n1449 , n250 , n1799 );
    not g1159 ( n1781 , n3224 );
    not g1160 ( n1545 , n2985 );
    or g1161 ( n1133 , n3434 , n509 );
    and g1162 ( n2668 , n3640 , n3914 );
    nor g1163 ( n1398 , n3373 , n1452 );
    not g1164 ( n1456 , n2856 );
    not g1165 ( n2891 , n604 );
    or g1166 ( n1598 , n1826 , n2739 );
    not g1167 ( n1575 , n2775 );
    not g1168 ( n3286 , n2946 );
    or g1169 ( n2603 , n1470 , n1188 );
    and g1170 ( n2325 , n2518 , n704 );
    nor g1171 ( n2787 , n2525 , n3040 );
    or g1172 ( n315 , n2281 , n2127 );
    or g1173 ( n3592 , n3082 , n1705 );
    nor g1174 ( n3140 , n1657 , n1928 );
    or g1175 ( n2185 , n2168 , n400 );
    and g1176 ( n2512 , n550 , n1492 );
    not g1177 ( n2636 , n2396 );
    or g1178 ( n58 , n3914 , n3692 );
    or g1179 ( n524 , n261 , n465 );
    and g1180 ( n2181 , n3019 , n1885 );
    nor g1181 ( n935 , n3590 , n2046 );
    or g1182 ( n791 , n3440 , n2778 );
    nor g1183 ( n3558 , n3043 , n386 );
    nor g1184 ( n3315 , n1130 , n1193 );
    and g1185 ( n108 , n1674 , n2775 );
    or g1186 ( n1682 , n487 , n880 );
    and g1187 ( n1985 , n1893 , n923 );
    and g1188 ( n151 , n3136 , n1480 );
    and g1189 ( n1803 , n3803 , n1216 );
    nor g1190 ( n1140 , n2051 , n2831 );
    buf g1191 ( n437 , n2625 );
    nor g1192 ( n3082 , n3682 , n853 );
    and g1193 ( n1934 , n2714 , n56 );
    or g1194 ( n3782 , n3331 , n1228 );
    not g1195 ( n2229 , n1195 );
    or g1196 ( n1405 , n1985 , n3834 );
    and g1197 ( n1501 , n1670 , n1838 );
    and g1198 ( n1247 , n1350 , n3441 );
    nor g1199 ( n3138 , n3610 , n207 );
    or g1200 ( n1863 , n3261 , n3742 );
    or g1201 ( n1204 , n1450 , n3096 );
    nor g1202 ( n1329 , n3011 , n602 );
    and g1203 ( n2664 , n1312 , n1292 );
    or g1204 ( n3728 , n1713 , n1579 );
    and g1205 ( n629 , n2789 , n2573 );
    not g1206 ( n2758 , n3294 );
    and g1207 ( n1789 , n2594 , n236 );
    or g1208 ( n2025 , n424 , n1414 );
    nor g1209 ( n3237 , n2656 , n1546 );
    not g1210 ( n1494 , n3763 );
    or g1211 ( n3157 , n2110 , n3120 );
    and g1212 ( n3487 , n2229 , n1316 );
    not g1213 ( n1272 , n3155 );
    nor g1214 ( n2361 , n1907 , n3527 );
    or g1215 ( n955 , n2077 , n2115 );
    and g1216 ( n1333 , n3483 , n3518 );
    and g1217 ( n443 , n2769 , n564 );
    or g1218 ( n2468 , n941 , n3692 );
    and g1219 ( n2875 , n3007 , n2433 );
    nor g1220 ( n2874 , n1751 , n2790 );
    and g1221 ( n750 , n230 , n364 );
    and g1222 ( n2767 , n3200 , n3726 );
    not g1223 ( n369 , n446 );
    or g1224 ( n2961 , n3122 , n1874 );
    and g1225 ( n2364 , n2871 , n2755 );
    not g1226 ( n1365 , n752 );
    and g1227 ( n1783 , n3040 , n2525 );
    or g1228 ( n2899 , n3338 , n3394 );
    and g1229 ( n3039 , n17 , n199 );
    and g1230 ( n2794 , n3818 , n896 );
    or g1231 ( n660 , n667 , n3118 );
    nor g1232 ( n106 , n2222 , n2903 );
    and g1233 ( n3450 , n844 , n2567 );
    and g1234 ( n3350 , n2152 , n3600 );
    or g1235 ( n1556 , n3484 , n2607 );
    or g1236 ( n3540 , n2986 , n3903 );
    and g1237 ( n344 , n3595 , n94 );
    or g1238 ( n1927 , n1086 , n2148 );
    and g1239 ( n2334 , n3517 , n3501 );
    or g1240 ( n2379 , n3537 , n239 );
    not g1241 ( n2120 , n3538 );
    not g1242 ( n109 , n1167 );
    nor g1243 ( n931 , n3213 , n769 );
    not g1244 ( n1752 , n1432 );
    and g1245 ( n3190 , n2039 , n1054 );
    nor g1246 ( n2500 , n795 , n3866 );
    or g1247 ( n553 , n2596 , n2559 );
    nor g1248 ( n1531 , n2290 , n972 );
    or g1249 ( n3587 , n2243 , n3903 );
    not g1250 ( n1784 , n3124 );
    or g1251 ( n1030 , n1274 , n3169 );
    not g1252 ( n3397 , n1285 );
    and g1253 ( n1074 , n1184 , n3036 );
    or g1254 ( n304 , n3314 , n2292 );
    or g1255 ( n368 , n2648 , n3466 );
    and g1256 ( n2702 , n1902 , n2742 );
    or g1257 ( n2566 , n1862 , n1916 );
    or g1258 ( n3482 , n1561 , n1410 );
    nor g1259 ( n1174 , n3308 , n3910 );
    and g1260 ( n651 , n300 , n1613 );
    or g1261 ( n1092 , n3574 , n1052 );
    or g1262 ( n1503 , n50 , n490 );
    and g1263 ( n3613 , n2678 , n3521 );
    not g1264 ( n11 , n2685 );
    or g1265 ( n1751 , n2593 , n925 );
    not g1266 ( n2716 , n3379 );
    and g1267 ( n1580 , n3010 , n2644 );
    or g1268 ( n2912 , n3048 , n1840 );
    and g1269 ( n242 , n141 , n3792 );
    or g1270 ( n1608 , n2505 , n2405 );
    nor g1271 ( n2588 , n2170 , n311 );
    not g1272 ( n115 , n33 );
    not g1273 ( n3429 , n3711 );
    and g1274 ( n1200 , n533 , n3654 );
    and g1275 ( n1939 , n3487 , n3668 );
    or g1276 ( n1836 , n2257 , n2469 );
    or g1277 ( n505 , n1831 , n2607 );
    nor g1278 ( n455 , n2964 , n3039 );
    and g1279 ( n229 , n1397 , n627 );
    not g1280 ( n562 , n1341 );
    and g1281 ( n2770 , n1871 , n1805 );
    not g1282 ( n721 , n1144 );
    and g1283 ( n3335 , n736 , n3799 );
    or g1284 ( n2138 , n2157 , n3169 );
    or g1285 ( n3059 , n1305 , n2956 );
    or g1286 ( n609 , n1306 , n1125 );
    buf g1287 ( n200 , n3548 );
    nor g1288 ( n2367 , n1719 , n722 );
    or g1289 ( n964 , n1626 , n2611 );
    nor g1290 ( n1270 , n2245 , n616 );
    or g1291 ( n2962 , n353 , n3396 );
    not g1292 ( n2103 , n2946 );
    and g1293 ( n1626 , n2086 , n1981 );
    and g1294 ( n34 , n2556 , n712 );
    not g1295 ( n3560 , n2986 );
    and g1296 ( n1066 , n3894 , n1590 );
    or g1297 ( n410 , n3553 , n3887 );
    or g1298 ( n3568 , n1347 , n1207 );
    and g1299 ( n86 , n3485 , n699 );
    or g1300 ( n1220 , n3876 , n1443 );
    nor g1301 ( n638 , n3825 , n3099 );
    and g1302 ( n1147 , n2343 , n1769 );
    nor g1303 ( n1351 , n1908 , n442 );
    nor g1304 ( n2923 , n1232 , n2845 );
    not g1305 ( n2016 , n495 );
    and g1306 ( n8 , n1456 , n1392 );
    and g1307 ( n3127 , n2071 , n3825 );
    and g1308 ( n3180 , n3205 , n3529 );
    or g1309 ( n1159 , n1002 , n3829 );
    and g1310 ( n3411 , n2701 , n2243 );
    and g1311 ( n3590 , n365 , n2986 );
    not g1312 ( n1223 , n954 );
    and g1313 ( n1042 , n1293 , n801 );
    and g1314 ( n3668 , n2717 , n270 );
    nor g1315 ( n1610 , n1195 , n2156 );
    and g1316 ( n2207 , n839 , n2066 );
    and g1317 ( n1168 , n2921 , n2979 );
    nor g1318 ( n3535 , n1841 , n1699 );
    or g1319 ( n3135 , n1527 , n698 );
    or g1320 ( n744 , n3708 , n571 );
    or g1321 ( n1577 , n2037 , n3903 );
    nor g1322 ( n2572 , n2794 , n811 );
    not g1323 ( n3892 , n2946 );
    or g1324 ( n879 , n1136 , n1188 );
    not g1325 ( n1199 , n2006 );
    and g1326 ( n3132 , n83 , n1311 );
    or g1327 ( n1371 , n2430 , n3692 );
    and g1328 ( n2862 , n1106 , n2850 );
    and g1329 ( n3534 , n3911 , n318 );
    and g1330 ( n1995 , n1498 , n3861 );
    nor g1331 ( n2203 , n1166 , n3207 );
    nor g1332 ( n821 , n1457 , n1477 );
    not g1333 ( n1069 , n3606 );
    and g1334 ( n1595 , n1681 , n27 );
    nor g1335 ( n1971 , n3613 , n2894 );
    and g1336 ( n2246 , n721 , n1576 );
    and g1337 ( n328 , n2983 , n3148 );
    and g1338 ( n1910 , n2325 , n3812 );
    or g1339 ( n1955 , n1012 , n994 );
    or g1340 ( n1217 , n2749 , n2452 );
    and g1341 ( n0 , n1899 , n798 );
    and g1342 ( n1275 , n1816 , n1407 );
    or g1343 ( n2296 , n3027 , n3449 );
    or g1344 ( n418 , n3215 , n3692 );
    nor g1345 ( n347 , n2859 , n2769 );
    and g1346 ( n3678 , n1257 , n398 );
    and g1347 ( n1463 , n3483 , n3869 );
    nor g1348 ( n2019 , n2361 , n871 );
    nor g1349 ( n2509 , n2289 , n1188 );
    and g1350 ( n3284 , n102 , n3116 );
    or g1351 ( n1424 , n2199 , n1965 );
    or g1352 ( n104 , n2744 , n3684 );
    and g1353 ( n3746 , n2447 , n2977 );
    nor g1354 ( n1798 , n15 , n1224 );
    nor g1355 ( n1447 , n33 , n978 );
    not g1356 ( n3246 , n1341 );
    and g1357 ( n2254 , n2543 , n2353 );
    not g1358 ( n3642 , n2702 );
    or g1359 ( n799 , n2002 , n1992 );
    and g1360 ( n733 , n2796 , n3472 );
    not g1361 ( n136 , n527 );
    and g1362 ( n2959 , n3700 , n3370 );
    buf g1363 ( n3483 , n2881 );
    and g1364 ( n3019 , n1264 , n2889 );
    or g1365 ( n3121 , n1827 , n48 );
    nor g1366 ( n2197 , n2173 , n2360 );
    not g1367 ( n67 , n3608 );
    and g1368 ( n1152 , n2769 , n3385 );
    or g1369 ( n2886 , n796 , n3466 );
    or g1370 ( n2764 , n1067 , n3425 );
    or g1371 ( n440 , n737 , n3395 );
    and g1372 ( n1733 , n1624 , n3553 );
    nor g1373 ( n2591 , n2210 , n2237 );
    and g1374 ( n1210 , n3271 , n3272 );
    nor g1375 ( n192 , n3490 , n2951 );
    not g1376 ( n3604 , n3379 );
    nor g1377 ( n2409 , n985 , n1424 );
    and g1378 ( n3344 , n1845 , n3657 );
    and g1379 ( n2718 , n2838 , n2578 );
    not g1380 ( n299 , n2263 );
    buf g1381 ( n3449 , n3900 );
    or g1382 ( n3067 , n1606 , n3636 );
    not g1383 ( n1994 , n1907 );
    or g1384 ( n1019 , n2968 , n3903 );
    or g1385 ( n1363 , n3310 , n3015 );
    nor g1386 ( n898 , n3265 , n3907 );
    or g1387 ( n2384 , n1406 , n3807 );
    not g1388 ( n1057 , n991 );
    and g1389 ( n3022 , n1823 , n373 );
    or g1390 ( n550 , n256 , n3466 );
    or g1391 ( n3064 , n3477 , n2713 );
    not g1392 ( n3164 , n3370 );
    and g1393 ( n871 , n511 , n3843 );
    not g1394 ( n3260 , n3833 );
    nor g1395 ( n3141 , n2606 , n2956 );
    and g1396 ( n1259 , n3797 , n1712 );
    and g1397 ( n2727 , n2965 , n2161 );
    and g1398 ( n3247 , n2963 , n3100 );
    not g1399 ( n1165 , n3686 );
    nor g1400 ( n2631 , n709 , n3902 );
    not g1401 ( n138 , n1163 );
    or g1402 ( n1851 , n3034 , n3466 );
    or g1403 ( n1385 , n2924 , n1129 );
    nor g1404 ( n2684 , n3106 , n3052 );
    and g1405 ( n2063 , n2834 , n3749 );
    and g1406 ( n801 , n372 , n3680 );
    nor g1407 ( n993 , n3326 , n59 );
    and g1408 ( n320 , n2360 , n1542 );
    and g1409 ( n3200 , n2055 , n938 );
    and g1410 ( n2617 , n1272 , n582 );
    and g1411 ( n2031 , n2216 , n2984 );
    and g1412 ( n548 , n3906 , n2006 );
    or g1413 ( n523 , n2703 , n1854 );
    and g1414 ( n3770 , n2917 , n3340 );
    or g1415 ( n3473 , n3071 , n2571 );
    and g1416 ( n2086 , n3514 , n2462 );
    or g1417 ( n3497 , n2075 , n2389 );
    or g1418 ( n2276 , n1807 , n1207 );
    nor g1419 ( n793 , n1136 , n279 );
    and g1420 ( n400 , n1293 , n2718 );
    and g1421 ( n3838 , n466 , n1927 );
    or g1422 ( n2557 , n1627 , n3128 );
    or g1423 ( n1078 , n2060 , n3865 );
    and g1424 ( n1079 , n1860 , n3781 );
    or g1425 ( n1361 , n651 , n2003 );
    and g1426 ( n448 , n2603 , n2104 );
    or g1427 ( n2908 , n2856 , n1188 );
    nor g1428 ( n961 , n2516 , n3647 );
    and g1429 ( n3869 , n656 , n673 );
    nor g1430 ( n973 , n1932 , n1768 );
    and g1431 ( n79 , n551 , n3004 );
    or g1432 ( n1855 , n3364 , n548 );
    buf g1433 ( n3466 , n665 );
    or g1434 ( n2271 , n3557 , n3346 );
    not g1435 ( n2950 , n102 );
    nor g1436 ( n3327 , n1181 , n2815 );
    and g1437 ( n829 , n87 , n519 );
    not g1438 ( n3360 , n3887 );
    or g1439 ( n1727 , n2188 , n3764 );
    not g1440 ( n2870 , n1761 );
    or g1441 ( n934 , n1027 , n3903 );
    nor g1442 ( n2362 , n3009 , n2489 );
    or g1443 ( n2313 , n3423 , n908 );
    not g1444 ( n2056 , n3379 );
    and g1445 ( n352 , n3385 , n3397 );
    or g1446 ( n3014 , n2286 , n1342 );
    and g1447 ( n2249 , n2284 , n3313 );
    nor g1448 ( n2442 , n1765 , n1554 );
    nor g1449 ( n3055 , n1163 , n3645 );
    not g1450 ( n1962 , n219 );
    not g1451 ( n968 , n1583 );
    and g1452 ( n1685 , n2546 , n3806 );
    and g1453 ( n684 , n2301 , n3555 );
    or g1454 ( n2299 , n3443 , n3433 );
    and g1455 ( n2611 , n2086 , n1515 );
    and g1456 ( n1812 , n2625 , n3180 );
    or g1457 ( n1300 , n3349 , n2632 );
    and g1458 ( n1697 , n3597 , n227 );
    and g1459 ( n1931 , n3761 , n3639 );
    not g1460 ( n1164 , n1836 );
    not g1461 ( n510 , n1585 );
    and g1462 ( n94 , n3147 , n595 );
    and g1463 ( n2672 , n1133 , n2375 );
    and g1464 ( n739 , n2630 , n646 );
    and g1465 ( n395 , n1433 , n3614 );
    and g1466 ( n1346 , n3507 , n3121 );
    not g1467 ( n1170 , n2363 );
    and g1468 ( n1977 , n2231 , n3464 );
    or g1469 ( n390 , n3790 , n246 );
    nor g1470 ( n1744 , n1742 , n3745 );
    not g1471 ( n1246 , n1766 );
    nor g1472 ( n3493 , n27 , n3848 );
    and g1473 ( n294 , n2625 , n3585 );
    and g1474 ( n1948 , n437 , n1194 );
    or g1475 ( n2977 , n3565 , n2091 );
    nor g1476 ( n3750 , n2928 , n2241 );
    not g1477 ( n3357 , n1861 );
    or g1478 ( n1635 , n3204 , n3770 );
    nor g1479 ( n3299 , n3238 , n2962 );
    nor g1480 ( n366 , n3481 , n2319 );
    or g1481 ( n1320 , n1321 , n1843 );
    or g1482 ( n3445 , n3084 , n3333 );
    or g1483 ( n3068 , n3713 , n478 );
    nor g1484 ( n3554 , n1496 , n689 );
    not g1485 ( n1382 , n325 );
    or g1486 ( n2375 , n580 , n571 );
    and g1487 ( n3911 , n3447 , n2634 );
    and g1488 ( n428 , n1490 , n2469 );
    and g1489 ( n2876 , n2741 , n1844 );
    or g1490 ( n3521 , n2615 , n908 );
    and g1491 ( n1877 , n3179 , n598 );
    or g1492 ( n1000 , n2288 , n2924 );
    or g1493 ( n508 , n1536 , n81 );
    and g1494 ( n948 , n2095 , n3301 );
    or g1495 ( n3783 , n2784 , n831 );
    or g1496 ( n1377 , n112 , n2770 );
    and g1497 ( n2 , n1498 , n362 );
    and g1498 ( n1652 , n3134 , n3918 );
    or g1499 ( n1902 , n2322 , n3169 );
    and g1500 ( n3456 , n2472 , n1547 );
    and g1501 ( n3636 , n639 , n913 );
    nor g1502 ( n2097 , n1372 , n2318 );
    nor g1503 ( n2922 , n3181 , n3817 );
    not g1504 ( n3102 , n256 );
    not g1505 ( n962 , n3060 );
    and g1506 ( n156 , n3759 , n1713 );
    or g1507 ( n1638 , n1338 , n3742 );
    and g1508 ( n21 , n3324 , n1338 );
    or g1509 ( n3850 , n2236 , n3910 );
    and g1510 ( n2342 , n3483 , n1412 );
    and g1511 ( n3320 , n3478 , n3585 );
    nor g1512 ( n1117 , n977 , n3432 );
    or g1513 ( n1303 , n3897 , n3015 );
    and g1514 ( n342 , n2497 , n1997 );
    or g1515 ( n656 , n676 , n3466 );
    nor g1516 ( n1047 , n3224 , n1554 );
    not g1517 ( n3804 , n2595 );
    or g1518 ( n1376 , n3033 , n881 );
    nor g1519 ( n3652 , n2120 , n1782 );
    and g1520 ( n2809 , n2007 , n2302 );
    not g1521 ( n1552 , n1071 );
    not g1522 ( n3593 , n2056 );
    nor g1523 ( n2004 , n2064 , n1526 );
    or g1524 ( n2889 , n1542 , n3741 );
    or g1525 ( n187 , n2395 , n1850 );
    and g1526 ( n743 , n2203 , n2521 );
    or g1527 ( n2801 , n173 , n3858 );
    and g1528 ( n975 , n2086 , n861 );
    or g1529 ( n3792 , n2703 , n3692 );
    not g1530 ( n2881 , n1341 );
    not g1531 ( n237 , n3379 );
    nor g1532 ( n1513 , n1615 , n3421 );
    or g1533 ( n1654 , n3777 , n2950 );
    not g1534 ( n1293 , n2946 );
    and g1535 ( n3257 , n2693 , n2682 );
    not g1536 ( n3879 , n1116 );
    nor g1537 ( n3026 , n199 , n17 );
    and g1538 ( n619 , n2783 , n3880 );
    buf g1539 ( n963 , n3548 );
    or g1540 ( n297 , n1760 , n1669 );
    or g1541 ( n3657 , n1499 , n2136 );
    nor g1542 ( n918 , n1746 , n3567 );
    nor g1543 ( n957 , n3658 , n1554 );
    and g1544 ( n3235 , n1989 , n3679 );
    or g1545 ( n785 , n417 , n3690 );
    or g1546 ( n3813 , n422 , n761 );
    or g1547 ( n3755 , n498 , n3692 );
    nor g1548 ( n392 , n3552 , n935 );
    or g1549 ( n846 , n3808 , n3903 );
    or g1550 ( n2752 , n3632 , n1416 );
    or g1551 ( n1001 , n2738 , n509 );
    and g1552 ( n2544 , n2139 , n474 );
    and g1553 ( n102 , n3322 , n2427 );
    and g1554 ( n2340 , n437 , n3854 );
    not g1555 ( n2551 , n1526 );
    nor g1556 ( n2555 , n2674 , n3499 );
    or g1557 ( n920 , n2984 , n509 );
    and g1558 ( n3108 , n3907 , n22 );
    not g1559 ( n681 , n3731 );
    nor g1560 ( n1901 , n1947 , n3479 );
    and g1561 ( n3618 , n1937 , n813 );
    and g1562 ( n264 , n3783 , n3017 );
    nor g1563 ( n3660 , n745 , n926 );
    or g1564 ( n1986 , n378 , n1007 );
    not g1565 ( n380 , n2176 );
    and g1566 ( n2225 , n614 , n2894 );
    nor g1567 ( n2151 , n3598 , n701 );
    nor g1568 ( n288 , n1907 , n1893 );
    and g1569 ( n3890 , n1768 , n1932 );
    not g1570 ( n866 , n3233 );
    and g1571 ( n2411 , n3102 , n886 );
    not g1572 ( n2400 , n419 );
    or g1573 ( n897 , n2791 , n3113 );
    or g1574 ( n1394 , n960 , n1207 );
    or g1575 ( n2749 , n377 , n1584 );
    or g1576 ( n3116 , n705 , n735 );
    nor g1577 ( n458 , n2252 , n2125 );
    and g1578 ( n1342 , n3483 , n1480 );
    or g1579 ( n3001 , n762 , n3348 );
    or g1580 ( n2098 , n1163 , n509 );
    and g1581 ( n3570 , n701 , n3598 );
    not g1582 ( n394 , n3484 );
    or g1583 ( n3036 , n803 , n982 );
    or g1584 ( n1458 , n1811 , n2692 );
    and g1585 ( n2941 , n2316 , n3871 );
    nor g1586 ( n171 , n174 , n2389 );
    not g1587 ( n3409 , n1641 );
    and g1588 ( n361 , n307 , n2008 );
    or g1589 ( n2309 , n770 , n2220 );
    or g1590 ( n2346 , n2328 , n1642 );
    nor g1591 ( n1709 , n1756 , n3163 );
    or g1592 ( n2398 , n198 , n3038 );
    nor g1593 ( n1800 , n1533 , n2345 );
    or g1594 ( n1903 , n381 , n86 );
    nor g1595 ( n2993 , n3255 , n1554 );
    or g1596 ( n2717 , n2718 , n1182 );
    or g1597 ( n3580 , n3630 , n758 );
    or g1598 ( n1173 , n2698 , n3697 );
    nor g1599 ( n3363 , n2964 , n3111 );
    or g1600 ( n664 , n922 , n2388 );
    buf g1601 ( n3742 , n908 );
    and g1602 ( n497 , n825 , n1762 );
    or g1603 ( n411 , n1892 , n3318 );
    not g1604 ( n1353 , n3787 );
    not g1605 ( n3184 , n3379 );
    or g1606 ( n1023 , n2116 , n1207 );
    or g1607 ( n3148 , n1947 , n3887 );
    buf g1608 ( n509 , n1050 );
    and g1609 ( n1226 , n1604 , n2487 );
    nor g1610 ( n1242 , n602 , n1249 );
    or g1611 ( n3338 , n2972 , n2186 );
    nor g1612 ( n649 , n1611 , n423 );
    and g1613 ( n1518 , n2717 , n240 );
    not g1614 ( n3578 , n467 );
    and g1615 ( n3437 , n389 , n276 );
    not g1616 ( n722 , n3379 );
    not g1617 ( n1806 , n1662 );
    and g1618 ( n797 , n1367 , n3177 );
    not g1619 ( n2148 , n3379 );
    or g1620 ( n3842 , n3268 , n271 );
    not g1621 ( n251 , n2622 );
    nor g1622 ( n2952 , n152 , n237 );
    and g1623 ( n2198 , n3435 , n557 );
    and g1624 ( n179 , n763 , n2249 );
    or g1625 ( n2429 , n3384 , n2503 );
    and g1626 ( n1675 , n2274 , n411 );
    and g1627 ( n3517 , n2645 , n878 );
    nor g1628 ( n296 , n3237 , n2926 );
    not g1629 ( n206 , n2638 );
    not g1630 ( n2902 , n23 );
    and g1631 ( n2416 , n1182 , n2718 );
    or g1632 ( n1182 , n3623 , n3073 );
    or g1633 ( n825 , n3852 , n1188 );
    not g1634 ( n856 , n2625 );
    or g1635 ( n3478 , n2524 , n1011 );
    or g1636 ( n3242 , n8 , n1409 );
    and g1637 ( n598 , n273 , n3130 );
    or g1638 ( n3394 , n1225 , n1317 );
    or g1639 ( n210 , n1903 , n3150 );
    nor g1640 ( n3448 , n2024 , n3886 );
    or g1641 ( n1349 , n1047 , n931 );
    not g1642 ( n3840 , n579 );
    and g1643 ( n919 , n553 , n3359 );
    and g1644 ( n1407 , n2296 , n1534 );
    and g1645 ( n1811 , n2769 , n903 );
    nor g1646 ( n1649 , n446 , n1554 );
    and g1647 ( n824 , n168 , n743 );
    not g1648 ( n1718 , n710 );
    not g1649 ( n2827 , n1731 );
    or g1650 ( n500 , n2668 , n3250 );
    or g1651 ( n1870 , n1871 , n1529 );
    not g1652 ( n688 , n3247 );
    not g1653 ( n2223 , n3862 );
    or g1654 ( n3717 , n3736 , n2058 );
    or g1655 ( n1348 , n3092 , n246 );
    not g1656 ( n3725 , n1341 );
    and g1657 ( n1780 , n2359 , n742 );
    or g1658 ( n641 , n1393 , n2515 );
    or g1659 ( n1525 , n2105 , n1543 );
    nor g1660 ( n1286 , n3460 , n1727 );
    nor g1661 ( n2137 , n1302 , n3769 );
    and g1662 ( n1417 , n688 , n694 );
    or g1663 ( n947 , n590 , n2341 );
    and g1664 ( n2199 , n3242 , n1987 );
    or g1665 ( n3806 , n1179 , n726 );
    nor g1666 ( n1289 , n3353 , n2804 );
    nor g1667 ( n1231 , n764 , n324 );
    and g1668 ( n2867 , n1281 , n2119 );
    and g1669 ( n1430 , n60 , n84 );
    nor g1670 ( n2080 , n1032 , n2409 );
    or g1671 ( n1084 , n779 , n797 );
    or g1672 ( n2191 , n2535 , n3175 );
    and g1673 ( n556 , n1732 , n148 );
    not g1674 ( n7 , n3462 );
    and g1675 ( n419 , n681 , n710 );
    or g1676 ( n3004 , n1315 , n522 );
    and g1677 ( n2251 , n1066 , n109 );
    not g1678 ( n995 , n3030 );
    or g1679 ( n3677 , n1113 , n571 );
    nor g1680 ( n2879 , n1802 , n1222 );
    or g1681 ( n3301 , n1991 , n2345 );
    not g1682 ( n1306 , n869 );
    or g1683 ( n236 , n3303 , n3742 );
    not g1684 ( n630 , n2862 );
    and g1685 ( n1177 , n1562 , n2991 );
    nor g1686 ( n1070 , n163 , n538 );
    or g1687 ( n3365 , n2283 , n3541 );
    not g1688 ( n3878 , n2102 );
    and g1689 ( n3737 , n3077 , n1139 );
    nor g1690 ( n2078 , n2200 , n2513 );
    nor g1691 ( n1454 , n1156 , n3140 );
    and g1692 ( n2387 , n2475 , n534 );
    or g1693 ( n146 , n1251 , n3294 );
    not g1694 ( n2466 , n3023 );
    and g1695 ( n802 , n1452 , n3373 );
    not g1696 ( n3321 , n3871 );
    and g1697 ( n3543 , n916 , n423 );
    and g1698 ( n1483 , n3288 , n2333 );
    or g1699 ( n2227 , n1838 , n1670 );
    or g1700 ( n620 , n2643 , n402 );
    or g1701 ( n1625 , n1812 , n3104 );
    or g1702 ( n1519 , n337 , n3742 );
    nor g1703 ( n3591 , n363 , n3578 );
    not g1704 ( n1033 , n3208 );
    and g1705 ( n1975 , n2818 , n2729 );
    and g1706 ( n3440 , n1978 , n1679 );
    nor g1707 ( n3103 , n1956 , n2184 );
    or g1708 ( n107 , n3874 , n2354 );
    or g1709 ( n3611 , n2500 , n2795 );
    or g1710 ( n1746 , n671 , n1745 );
    and g1711 ( n2461 , n3502 , n3656 );
    or g1712 ( n2539 , n1882 , n2458 );
    and g1713 ( n755 , n3047 , n3430 );
    nor g1714 ( n2172 , n521 , n1127 );
    or g1715 ( n1441 , n1174 , n2422 );
    and g1716 ( n1813 , n2090 , n1757 );
    or g1717 ( n2075 , n1045 , n1698 );
    and g1718 ( n959 , n2472 , n3524 );
    nor g1719 ( n190 , n2941 , n1326 );
    not g1720 ( n302 , n2336 );
    or g1721 ( n937 , n3429 , n1118 );
    or g1722 ( n2714 , n1366 , n1188 );
    and g1723 ( n70 , n2099 , n3664 );
    not g1724 ( n406 , n3399 );
    and g1725 ( n1125 , n2041 , n1215 );
    nor g1726 ( n2949 , n3581 , n1554 );
    nor g1727 ( n1450 , n1572 , n856 );
    nor g1728 ( n4 , n1862 , n2657 );
    or g1729 ( n917 , n1906 , n1188 );
    or g1730 ( n1605 , n3296 , n3015 );
    nor g1731 ( n1928 , n263 , n2884 );
    and g1732 ( n2111 , n2021 , n3259 );
    and g1733 ( n1860 , n316 , n118 );
    nor g1734 ( n1225 , n1938 , n333 );
    not g1735 ( n3659 , n2946 );
    not g1736 ( n2686 , n3869 );
    and g1737 ( n1772 , n740 , n3393 );
    or g1738 ( n3447 , n76 , n1188 );
    and g1739 ( n3216 , n2293 , n2144 );
    or g1740 ( n1089 , n2061 , n3910 );
    or g1741 ( n1094 , n1171 , n1777 );
    nor g1742 ( n2323 , n3621 , n3689 );
    and g1743 ( n3855 , n1853 , n2751 );
    and g1744 ( n1594 , n562 , n3340 );
    and g1745 ( n259 , n1029 , n1589 );
    not g1746 ( n576 , n986 );
    or g1747 ( n123 , n3154 , n2727 );
    not g1748 ( n1622 , n966 );
    not g1749 ( n2318 , n3634 );
    or g1750 ( n2558 , n3263 , n425 );
    not g1751 ( n2230 , n3217 );
    or g1752 ( n3886 , n2958 , n3665 );
    buf g1753 ( n1341 , n2393 );
    and g1754 ( n185 , n948 , n809 );
    not g1755 ( n2649 , n1229 );
    or g1756 ( n2776 , n1239 , n1714 );
    and g1757 ( n72 , n437 , n1432 );
    not g1758 ( n1121 , n2946 );
    and g1759 ( n2924 , n491 , n2236 );
    or g1760 ( n2624 , n3152 , n1207 );
    not g1761 ( n835 , n1194 );
    not g1762 ( n1864 , n2967 );
    and g1763 ( n1724 , n1655 , n2134 );
    nor g1764 ( n3685 , n2195 , n258 );
    not g1765 ( n978 , n3379 );
    or g1766 ( n1413 , n3739 , n3903 );
    and g1767 ( n1236 , n3095 , n2466 );
    and g1768 ( n549 , n663 , n694 );
    or g1769 ( n674 , n3029 , n3127 );
    and g1770 ( n2614 , n1223 , n2149 );
    nor g1771 ( n487 , n859 , n1243 );
    not g1772 ( n2737 , n1150 );
    or g1773 ( n1546 , n2610 , n3915 );
    not g1774 ( n217 , n467 );
    nor g1775 ( n2145 , n1190 , n3135 );
    or g1776 ( n209 , n1425 , n319 );
    or g1777 ( n3090 , n3234 , n1132 );
    and g1778 ( n2091 , n2267 , n720 );
    or g1779 ( n2036 , n3686 , n1916 );
    or g1780 ( n3800 , n2419 , n3185 );
    nor g1781 ( n1875 , n2982 , n202 );
    or g1782 ( n1786 , n3731 , n761 );
    and g1783 ( n820 , n1566 , n117 );
    and g1784 ( n2654 , n3612 , n2079 );
    or g1785 ( n3359 , n1830 , n2824 );
    nor g1786 ( n2663 , n226 , n2490 );
    and g1787 ( n2552 , n2597 , n3626 );
    not g1788 ( n1211 , n1963 );
    nor g1789 ( n2926 , n2748 , n1289 );
    and g1790 ( n2077 , n3539 , n2414 );
    or g1791 ( n2067 , n675 , n866 );
    and g1792 ( n2723 , n3013 , n631 );
    and g1793 ( n2728 , n1893 , n2107 );
    and g1794 ( n3628 , n2190 , n1630 );
    and g1795 ( n3351 , n2490 , n226 );
    not g1796 ( n3419 , n2946 );
    and g1797 ( n2659 , n1977 , n3896 );
    or g1798 ( n37 , n1959 , n2432 );
    or g1799 ( n1834 , n3602 , n1990 );
    and g1800 ( n861 , n3265 , n1255 );
    or g1801 ( n2901 , n3917 , n2092 );
    not g1802 ( n1673 , n3867 );
    nor g1803 ( n3673 , n775 , n2565 );
    not g1804 ( n3863 , n2852 );
    or g1805 ( n859 , n1649 , n2323 );
    not g1806 ( n3202 , n3379 );
    and g1807 ( n3204 , n613 , n77 );
    not g1808 ( n365 , n2848 );
    or g1809 ( n552 , n940 , n3304 );
    nor g1810 ( n1148 , n2794 , n1788 );
    or g1811 ( n457 , n1484 , n748 );
    or g1812 ( n2532 , n2885 , n2010 );
    not g1813 ( n2167 , n2424 );
    or g1814 ( n140 , n805 , n2863 );
    nor g1815 ( n2267 , n2065 , n1283 );
    nor g1816 ( n745 , n3819 , n1057 );
    or g1817 ( n2818 , n3444 , n638 );
    not g1818 ( n25 , n2181 );
    nor g1819 ( n671 , n1807 , n2050 );
    nor g1820 ( n168 , n1880 , n3334 );
    nor g1821 ( n3432 , n151 , n2019 );
    nor g1822 ( n157 , n3911 , n3446 );
    not g1823 ( n2773 , n2563 );
    or g1824 ( n113 , n530 , n2523 );
    or g1825 ( n3339 , n2680 , n3126 );
    nor g1826 ( n3849 , n2663 , n544 );
    or g1827 ( n1921 , n2309 , n1159 );
    not g1828 ( n132 , n3039 );
    nor g1829 ( n678 , n609 , n3038 );
    not g1830 ( n2258 , n2946 );
    and g1831 ( n2746 , n3218 , n3192 );
    not g1832 ( n3683 , n3379 );
    or g1833 ( n3192 , n43 , n2329 );
    not g1834 ( n2994 , n3747 );
    not g1835 ( n1327 , n3020 );
    or g1836 ( n127 , n2706 , n3887 );
    not g1837 ( n2907 , n2590 );
    not g1838 ( n1753 , n3885 );
    nor g1839 ( n2488 , n1814 , n1654 );
    and g1840 ( n1691 , n2565 , n775 );
    or g1841 ( n147 , n601 , n908 );
    and g1842 ( n3387 , n730 , n2504 );
    or g1843 ( n3032 , n1847 , n1146 );
    and g1844 ( n1802 , n115 , n2820 );
    and g1845 ( n2206 , n1327 , n924 );
    nor g1846 ( n3223 , n2049 , n1172 );
    and g1847 ( n2099 , n2226 , n3059 );
    or g1848 ( n291 , n1263 , n1973 );
    or g1849 ( n273 , n1827 , n3169 );
    and g1850 ( n1526 , n736 , n61 );
    and g1851 ( n650 , n2264 , n2890 );
    or g1852 ( n292 , n13 , n3197 );
    not g1853 ( n65 , n533 );
    not g1854 ( n2518 , n3552 );
    and g1855 ( n3290 , n2085 , n699 );
    and g1856 ( n2656 , n2883 , n1863 );
    nor g1857 ( n1756 , n694 , n688 );
    or g1858 ( n2675 , n1879 , n3910 );
    not g1859 ( n655 , n2946 );
    not g1860 ( n1620 , n44 );
    not g1861 ( n2917 , n2687 );
    or g1862 ( n2739 , n3146 , n2821 );
    or g1863 ( n2772 , n1211 , n341 );
    not g1864 ( n1312 , n225 );
    and g1865 ( n527 , n1391 , n657 );
    and g1866 ( n2725 , n543 , n2764 );
    nor g1867 ( n852 , n2251 , n1783 );
    or g1868 ( n1339 , n3391 , n3038 );
    and g1869 ( n753 , n1910 , n2449 );
    not g1870 ( n2187 , n3618 );
    or g1871 ( n415 , n2731 , n3318 );
    not g1872 ( n6 , n1364 );
    nor g1873 ( n3499 , n2033 , n2362 );
    and g1874 ( n241 , n2016 , n116 );
    nor g1875 ( n1443 , n2637 , n1155 );
    nor g1876 ( n536 , n2659 , n887 );
    not g1877 ( n3170 , n1807 );
    or g1878 ( n2245 , n3872 , n2338 );
    or g1879 ( n1389 , n979 , n3714 );
    and g1880 ( n632 , n1854 , n2703 );
    or g1881 ( n387 , n1581 , n2100 );
    or g1882 ( n1460 , n2088 , n1646 );
    and g1883 ( n2123 , n3835 , n998 );
    and g1884 ( n3675 , n888 , n2706 );
    and g1885 ( n125 , n210 , n535 );
    not g1886 ( n2583 , n1933 );
    not g1887 ( n1694 , n3887 );
    or g1888 ( n2803 , n1980 , n215 );
    or g1889 ( n1192 , n160 , n661 );
    not g1890 ( n1208 , n941 );
    or g1891 ( n1137 , n3836 , n3692 );
    and g1892 ( n855 , n3688 , n445 );
    not g1893 ( n3501 , n1412 );
    not g1894 ( n2774 , n3379 );
    and g1895 ( n714 , n2666 , n3186 );
    not g1896 ( n1998 , n503 );
    nor g1897 ( n3670 , n815 , n1816 );
    not g1898 ( n245 , n2333 );
    or g1899 ( n535 , n2619 , n1079 );
    or g1900 ( n1459 , n1995 , n1951 );
    or g1901 ( n1961 , n536 , n1687 );
    and g1902 ( n883 , n3199 , n298 );
    and g1903 ( n3250 , n3640 , n2653 );
    or g1904 ( n1894 , n2049 , n1207 );
    not g1905 ( n1895 , n2946 );
    or g1906 ( n3239 , n1282 , n3616 );
    or g1907 ( n60 , n953 , n1898 );
    nor g1908 ( n1359 , n3908 , n3448 );
    or g1909 ( n1254 , n2642 , n2155 );
    nor g1910 ( n1653 , n2596 , n3359 );
    or g1911 ( n2089 , n2119 , n1281 );
    and g1912 ( n585 , n768 , n3011 );
    and g1913 ( n666 , n3723 , n3540 );
    or g1914 ( n38 , n2030 , n1639 );
    and g1915 ( n2161 , n2618 , n1386 );
    and g1916 ( n3314 , n3692 , n1897 );
    or g1917 ( n2302 , n1068 , n740 );
    or g1918 ( n3579 , n359 , n1188 );
    and g1919 ( n3508 , n3421 , n1615 );
    and g1920 ( n1876 , n1716 , n739 );
    or g1921 ( n2531 , n1849 , n2892 );
    nor g1922 ( n2528 , n3430 , n2898 );
    not g1923 ( n3650 , n2938 );
    not g1924 ( n2418 , n2832 );
    or g1925 ( n3666 , n428 , n131 );
    or g1926 ( n1569 , n754 , n2898 );
    and g1927 ( n1782 , n3838 , n1396 );
    or g1928 ( n92 , n2157 , n881 );
    nor g1929 ( n1153 , n3545 , n906 );
    nor g1930 ( n3802 , n1879 , n1033 );
    and g1931 ( n3734 , n772 , n3323 );
    or g1932 ( n636 , n2627 , n2878 );
    or g1933 ( n1422 , n2414 , n3449 );
    not g1934 ( n3654 , n1008 );
    or g1935 ( n57 , n1168 , n2455 );
    or g1936 ( n421 , n106 , n987 );
    not g1937 ( n3134 , n2946 );
    not g1938 ( n3491 , n1481 );
    or g1939 ( n2038 , n2529 , n3742 );
    and g1940 ( n1839 , n12 , n2005 );
    or g1941 ( n2681 , n460 , n1791 );
    or g1942 ( n80 , n3264 , n1639 );
    or g1943 ( n3337 , n1779 , n3887 );
    nor g1944 ( n808 , n3342 , n1278 );
    or g1945 ( n1191 , n3208 , n3015 );
    or g1946 ( n2645 , n2587 , n1916 );
    and g1947 ( n2507 , n1353 , n2121 );
    not g1948 ( n3334 , n2615 );
    and g1949 ( n807 , n1834 , n2465 );
    and g1950 ( n2574 , n3839 , n2620 );
    or g1951 ( n2202 , n2250 , n989 );
    or g1952 ( n1085 , n2414 , n3539 );
    not g1953 ( n3801 , n623 );
    or g1954 ( n716 , n1104 , n1262 );
    and g1955 ( n3028 , n405 , n1062 );
    or g1956 ( n2015 , n3619 , n1478 );
    nor g1957 ( n2643 , n2896 , n988 );
    and g1958 ( n1195 , n584 , n630 );
    or g1959 ( n965 , n1150 , n761 );
    buf g1960 ( n2946 , n2393 );
    not g1961 ( n39 , n180 );
    or g1962 ( n1717 , n1403 , n1207 );
    and g1963 ( n1009 , n2230 , n818 );
    and g1964 ( n3040 , n2799 , n1553 );
    nor g1965 ( n3444 , n687 , n2607 );
    or g1966 ( n2586 , n286 , n2558 );
    nor g1967 ( n690 , n660 , n3052 );
    nor g1968 ( n2661 , n1473 , n508 );
    and g1969 ( n3219 , n2526 , n214 );
    and g1970 ( n752 , n3850 , n1303 );
    nor g1971 ( n3465 , n2487 , n2169 );
    or g1972 ( n784 , n2385 , n3531 );
    or g1973 ( n1283 , n3734 , n289 );
    not g1974 ( n870 , n2211 );
    nor g1975 ( n3736 , n1499 , n1334 );
    or g1976 ( n3722 , n915 , n867 );
    or g1977 ( n1970 , n169 , n2847 );
    or g1978 ( n1655 , n1360 , n2996 );
    or g1979 ( n3415 , n895 , n3015 );
    nor g1980 ( n845 , n325 , n414 );
    or g1981 ( n1427 , n3685 , n208 );
    not g1982 ( n2651 , n2056 );
    or g1983 ( n2673 , n464 , n1075 );
    not g1984 ( n414 , n1219 );
    or g1985 ( n727 , n96 , n509 );
    nor g1986 ( n2947 , n582 , n1272 );
    nor g1987 ( n3745 , n2900 , n1288 );
    or g1988 ( n2180 , n47 , n2661 );
    not g1989 ( n2288 , n889 );
    or g1990 ( n2460 , n293 , n3015 );
    or g1991 ( n3244 , n2781 , n447 );
    nor g1992 ( n2261 , n474 , n1989 );
    or g1993 ( n2452 , n3414 , n1148 );
    or g1994 ( n2578 , n3633 , n571 );
    not g1995 ( n3240 , n971 );
    and g1996 ( n1107 , n3012 , n2613 );
    or g1997 ( n2391 , n128 , n1739 );
    nor g1998 ( n2593 , n2358 , n53 );
    nor g1999 ( n3758 , n891 , n395 );
    or g2000 ( n1067 , n2527 , n3037 );
    or g2001 ( n813 , n1116 , n3903 );
    and g2002 ( n2306 , n879 , n1363 );
    or g2003 ( n2101 , n3178 , n196 );
    and g2004 ( n1708 , n1023 , n2721 );
    nor g2005 ( n2698 , n1481 , n2649 );
    and g2006 ( n3198 , n368 , n58 );
    or g2007 ( n1185 , n2702 , n323 );
    and g2008 ( n3625 , n1784 , n2788 );
    or g2009 ( n2201 , n3323 , n509 );
    or g2010 ( n583 , n1743 , n3184 );
    and g2011 ( n1698 , n23 , n356 );
    and g2012 ( n1448 , n3404 , n1724 );
    nor g2013 ( n2934 , n512 , n1153 );
    nor g2014 ( n2560 , n2894 , n2652 );
    and g2015 ( n900 , n437 , n3247 );
    or g2016 ( n375 , n3624 , n3742 );
    and g2017 ( n880 , n1243 , n2512 );
    or g2018 ( n2029 , n2560 , n1979 );
    or g2019 ( n3329 , n1933 , n3692 );
    nor g2020 ( n1825 , n1267 , n1231 );
    or g2021 ( n1957 , n2813 , n62 );
    not g2022 ( n1871 , n1736 );
    or g2023 ( n2577 , n644 , n3057 );
    or g2024 ( n1087 , n2189 , n1207 );
    or g2025 ( n3332 , n1829 , n1898 );
    not g2026 ( n2608 , n3051 );
    not g2027 ( n2831 , n2430 );
    and g2028 ( n3193 , n1165 , n3189 );
    and g2029 ( n3065 , n2138 , n375 );
    nor g2030 ( n3418 , n108 , n436 );
    or g2031 ( n3645 , n1806 , n836 );
    and g2032 ( n2017 , n3240 , n284 );
    or g2033 ( n1072 , n99 , n125 );
    not g2034 ( n2851 , n998 );
    or g2035 ( n1762 , n912 , n1101 );
    not g2036 ( n3626 , n3006 );
    or g2037 ( n1520 , n385 , n672 );
    and g2038 ( n2729 , n1149 , n846 );
    and g2039 ( n3788 , n3483 , n1713 );
    nor g2040 ( n590 , n915 , n1438 );
    nor g2041 ( n823 , n3530 , n1188 );
    and g2042 ( n843 , n3542 , n3322 );
    not g2043 ( n1367 , n1341 );
    or g2044 ( n3811 , n2628 , n1916 );
    or g2045 ( n575 , n990 , n347 );
    and g2046 ( n2472 , n1891 , n1587 );
    and g2047 ( n2298 , n451 , n789 );
    or g2048 ( n1402 , n2896 , n3692 );
    not g2049 ( n3018 , n2925 );
    or g2050 ( n191 , n582 , n509 );
    not g2051 ( n3111 , n1079 );
    not g2052 ( n1792 , n2564 );
    and g2053 ( n607 , n1427 , n2554 );
    nor g2054 ( n554 , n800 , n98 );
    and g2055 ( n581 , n384 , n3117 );
    and g2056 ( n3245 , n2154 , n2496 );
    nor g2057 ( n370 , n1770 , n3837 );
    not g2058 ( n2980 , n1341 );
    or g2059 ( n3446 , n318 , n981 );
    or g2060 ( n3768 , n3561 , n1567 );
    or g2061 ( n2989 , n2863 , n137 );
    and g2062 ( n158 , n467 , n254 );
    or g2063 ( n2247 , n2547 , n2384 );
    and g2064 ( n1375 , n2707 , n833 );
    and g2065 ( n3006 , n1945 , n3669 );
    not g2066 ( n130 , n3180 );
    or g2067 ( n2093 , n2131 , n806 );
    and g2068 ( n570 , n3899 , n1500 );
    or g2069 ( n1889 , n573 , n3428 );
    or g2070 ( n2301 , n18 , n1188 );
    and g2071 ( n476 , n2745 , n2299 );
    or g2072 ( n1790 , n1328 , n1263 );
    and g2073 ( n1570 , n2351 , n2043 );
    buf g2074 ( n1188 , n3666 );
    not g2075 ( n495 , n1664 );
    not g2076 ( n595 , n2279 );
    nor g2077 ( n3564 , n3216 , n2471 );
    not g2078 ( n2697 , n1899 );
    or g2079 ( n2846 , n139 , n1916 );
    and g2080 ( n944 , n420 , n2223 );
    nor g2081 ( n460 , n1700 , n3698 );
    and g2082 ( n1720 , n2625 , n2964 );
    and g2083 ( n2341 , n927 , n2912 );
    nor g2084 ( n2957 , n3081 , n296 );
    or g2085 ( n1127 , n1162 , n1471 );
    not g2086 ( n1978 , n617 );
    or g2087 ( n479 , n945 , n3449 );
    and g2088 ( n2824 , n1376 , n92 );
    and g2089 ( n3126 , n3483 , n3245 );
    and g2090 ( n2033 , n6 , n598 );
    or g2091 ( n1701 , n1335 , n1218 );
    not g2092 ( n3716 , n1233 );
    or g2093 ( n153 , n3474 , n3692 );
    or g2094 ( n1022 , n3693 , n3533 );
    nor g2095 ( n3234 , n760 , n70 );
    or g2096 ( n3555 , n2768 , n1101 );
    not g2097 ( n2273 , n1341 );
    or g2098 ( n3662 , n421 , n2961 );
    not g2099 ( n622 , n1358 );
    and g2100 ( n2853 , n3182 , n1605 );
    nor g2101 ( n2002 , n1831 , n1796 );
    or g2102 ( n2592 , n2057 , n3235 );
    not g2103 ( n3280 , n420 );
    nor g2104 ( n3056 , n564 , n2935 );
    and g2105 ( n3605 , n2903 , n2222 );
    and g2106 ( n698 , n1385 , n2514 );
    not g2107 ( n2130 , n854 );
    not g2108 ( n3647 , n3221 );
    and g2109 ( n3569 , n3091 , n3712 );
    or g2110 ( n3588 , n1233 , n908 );
    or g2111 ( n2963 , n1219 , n1916 );
    and g2112 ( n1982 , n437 , n2741 );
    nor g2113 ( n1968 , n1809 , n3070 );
    or g2114 ( n20 , n2438 , n3788 );
    not g2115 ( n1104 , n555 );
    and g2116 ( n1527 , n3638 , n3172 );
    or g2117 ( n787 , n2357 , n1941 );
    and g2118 ( n2265 , n791 , n2227 );
    nor g2119 ( n429 , n765 , n3194 );
    and g2120 ( n2124 , n3183 , n974 );
    and g2121 ( n3010 , n2671 , n1884 );
    or g2122 ( n2637 , n1357 , n1290 );
    not g2123 ( n2112 , n637 );
    not g2124 ( n1474 , n2587 );
    not g2125 ( n213 , n2595 );
    or g2126 ( n1172 , n177 , n3699 );
    nor g2127 ( n2900 , n116 , n3403 );
    or g2128 ( n1988 , n3233 , n3742 );
    nor g2129 ( n696 , n3222 , n1875 );
    nor g2130 ( n382 , n3492 , n95 );
    and g2131 ( n2523 , n1986 , n3532 );
    or g2132 ( n1952 , n3461 , n2854 );
    or g2133 ( n95 , n843 , n2809 );
    or g2134 ( n2154 , n1015 , n271 );
    not g2135 ( n2730 , n1821 );
    or g2136 ( n3130 , n3547 , n908 );
    and g2137 ( n270 , n1717 , n1638 );
    not g2138 ( n224 , n2935 );
    and g2139 ( n2421 , n1070 , n2118 );
    and g2140 ( n2108 , n2542 , n3065 );
    and g2141 ( n2541 , n3483 , n2166 );
    not g2142 ( n2981 , n3095 );
    nor g2143 ( n3201 , n2773 , n1712 );
    buf g2144 ( n1101 , n2062 );
    and g2145 ( n2719 , n1474 , n1924 );
    or g2146 ( n307 , n930 , n1603 );
    nor g2147 ( n2105 , n3051 , n831 );
    buf g2148 ( n2996 , n665 );
    or g2149 ( n996 , n182 , n1976 );
    or g2150 ( n1202 , n2373 , n2549 );
    and g2151 ( n3109 , n2769 , n1667 );
    or g2152 ( n2830 , n2576 , n1599 );
    or g2153 ( n1747 , n1805 , n3360 );
    and g2154 ( n2835 , n3717 , n3064 );
    or g2155 ( n646 , n1051 , n571 );
    or g2156 ( n2927 , n1514 , n2112 );
    not g2157 ( n3780 , n3511 );
    or g2158 ( n445 , n1434 , n908 );
    not g2159 ( n3316 , n1341 );
    and g2160 ( n3651 , n1597 , n1279 );
    or g2161 ( n788 , n3825 , n2071 );
    not g2162 ( n1146 , n2325 );
    and g2163 ( n50 , n2769 , n1528 );
    and g2164 ( n2781 , n2582 , n2228 );
    nor g2165 ( n1776 , n2902 , n1730 );
    and g2166 ( n2255 , n2607 , n1201 );
    nor g2167 ( n3146 , n1783 , n2042 );
    or g2168 ( n118 , n3340 , n2917 );
    or g2169 ( n1370 , n3729 , n3362 );
    not g2170 ( n3153 , n3379 );
    nor g2171 ( n2020 , n3749 , n2834 );
    or g2172 ( n1589 , n2448 , n1101 );
    and g2173 ( n2048 , n1494 , n304 );
    and g2174 ( n1295 , n3775 , n265 );
    and g2175 ( n869 , n1747 , n126 );
    and g2176 ( n3385 , n3811 , n2577 );
    and g2177 ( n3779 , n1893 , n3319 );
    or g2178 ( n3115 , n2602 , n1578 );
    or g2179 ( n2974 , n1210 , n2690 );
    and g2180 ( n3177 , n1573 , n3050 );
    or g2181 ( n1044 , n228 , n761 );
    and g2182 ( n77 , n260 , n1413 );
    nor g2183 ( n3694 , n3570 , n2278 );
    and g2184 ( n2390 , n406 , n1743 );
    and g2185 ( n1167 , n1087 , n418 );
    nor g2186 ( n3292 , n348 , n3450 );
    or g2187 ( n725 , n432 , n2704 );
    or g2188 ( n763 , n3253 , n1296 );
    or g2189 ( n2582 , n2719 , n167 );
    not g2190 ( n1818 , n2322 );
    not g2191 ( n1723 , n3245 );
    nor g2192 ( n621 , n3471 , n3188 );
    and g2193 ( n2407 , n3374 , n2547 );
    and g2194 ( n1742 , n3403 , n116 );
    or g2195 ( n2092 , n171 , n1955 );
    nor g2196 ( n1102 , n2061 , n3786 );
    or g2197 ( n1258 , n1838 , n3466 );
    or g2198 ( n121 , n2170 , n2317 );
    not g2199 ( n1214 , n2946 );
    and g2200 ( n420 , n1541 , n3251 );
    or g2201 ( n2704 , n794 , n750 );
    not g2202 ( n2828 , n1758 );
    nor g2203 ( n3166 , n2501 , n1767 );
    and g2204 ( n2135 , n1479 , n3437 );
    nor g2205 ( n3594 , n3383 , n3545 );
    nor g2206 ( n2641 , n1048 , n664 );
    and g2207 ( n2931 , n1508 , n1969 );
    not g2208 ( n1426 , n3754 );
    not g2209 ( n2204 , n2892 );
    or g2210 ( n3638 , n872 , n1389 );
    or g2211 ( n939 , n604 , n1101 );
    not g2212 ( n1989 , n467 );
    nor g2213 ( n3252 , n1375 , n541 );
    and g2214 ( n2921 , n1754 , n2272 );
    and g2215 ( n3380 , n1619 , n1158 );
    not g2216 ( n2536 , n3058 );
    nor g2217 ( n2422 , n2446 , n302 );
    not g2218 ( n3835 , n2723 );
    not g2219 ( n904 , n1269 );
    not g2220 ( n2819 , n3119 );
    nor g2221 ( n3488 , n183 , n3286 );
    and g2222 ( n1641 , n2891 , n810 );
    buf g2223 ( n2607 , n1188 );
    not g2224 ( n2745 , n2334 );
    nor g2225 ( n1842 , n644 , n1475 );
    nor g2226 ( n2857 , n3820 , n343 );
    and g2227 ( n3275 , n1555 , n3576 );
    or g2228 ( n1706 , n3335 , n93 );
    not g2229 ( n2350 , n757 );
    or g2230 ( n1558 , n192 , n493 );
    or g2231 ( n1699 , n3079 , n419 );
    and g2232 ( n3120 , n3566 , n2249 );
    and g2233 ( n2059 , n3334 , n1880 );
    nor g2234 ( n2122 , n352 , n3341 );
    or g2235 ( n3799 , n3162 , n3550 );
    nor g2236 ( n1340 , n3718 , n3575 );
    nor g2237 ( n3807 , n434 , n2148 );
    not g2238 ( n2090 , n3905 );
    or g2239 ( n201 , n2859 , n946 );
    not g2240 ( n3687 , n953 );
    or g2241 ( n2224 , n1958 , n3742 );
    not g2242 ( n3297 , n1491 );
    nor g2243 ( n2576 , n3233 , n2034 );
    not g2244 ( n3046 , n2625 );
    and g2245 ( n1593 , n2208 , n1804 );
    or g2246 ( n3793 , n2622 , n2136 );
    and g2247 ( n1591 , n560 , n2977 );
    or g2248 ( n3791 , n3030 , n1188 );
    nor g2249 ( n66 , n1844 , n2741 );
    not g2250 ( n1624 , n1829 );
    nor g2251 ( n1888 , n384 , n2273 );
    not g2252 ( n2129 , n1341 );
    and g2253 ( n731 , n594 , n1063 );
    or g2254 ( n2888 , n2137 , n654 );
    nor g2255 ( n1440 , n457 , n2901 );
    and g2256 ( n1187 , n2072 , n3030 );
    or g2257 ( n2850 , n2954 , n3887 );
    nor g2258 ( n2402 , n159 , n185 );
    and g2259 ( n765 , n850 , n3124 );
    not g2260 ( n195 , n644 );
    or g2261 ( n3515 , n1932 , n831 );
    nor g2262 ( n3331 , n423 , n2413 );
    or g2263 ( n1444 , n2017 , n1523 );
    not g2264 ( n2027 , n3815 );
    or g2265 ( n2789 , n691 , n3169 );
    not g2266 ( n1750 , n1341 );
    and g2267 ( n1560 , n2129 , n3117 );
    not g2268 ( n2235 , n492 );
    nor g2269 ( n453 , n3278 , n2382 );
    nor g2270 ( n3596 , n1415 , n3826 );
    not g2271 ( n295 , n3887 );
    and g2272 ( n1423 , n782 , n728 );
    and g2273 ( n3276 , n2273 , n1295 );
    and g2274 ( n1642 , n458 , n2013 );
    nor g2275 ( n1479 , n1940 , n2441 );
    and g2276 ( n628 , n2625 , n3912 );
    or g2277 ( n2406 , n3416 , n1207 );
    nor g2278 ( n1689 , n3266 , n3483 );
    nor g2279 ( n1020 , n1352 , n2022 );
    not g2280 ( n1284 , n2946 );
    and g2281 ( n3282 , n1575 , n3303 );
    nor g2282 ( n1799 , n2206 , n1825 );
    or g2283 ( n3112 , n2967 , n3449 );
    or g2284 ( n786 , n3055 , n3041 );
    nor g2285 ( n1508 , n2736 , n3561 );
    nor g2286 ( n1135 , n1663 , n1365 );
    or g2287 ( n938 , n2436 , n100 );
    and g2288 ( n1722 , n3725 , n830 );
    nor g2289 ( n990 , n3045 , n655 );
    or g2290 ( n1567 , n618 , n70 );
    and g2291 ( n605 , n2756 , n3217 );
    not g2292 ( n899 , n1253 );
    buf g2293 ( n3903 , n761 );
    and g2294 ( n1088 , n3744 , n3497 );
    or g2295 ( n3149 , n3608 , n2996 );
    or g2296 ( n1729 , n3245 , n24 );
    nor g2297 ( n2232 , n2144 , n2293 );
    or g2298 ( n3386 , n3101 , n3169 );
    or g2299 ( n316 , n77 , n613 );
    and g2300 ( n1313 , n3828 , n1765 );
    nor g2301 ( n1400 , n2459 , n2167 );
    and g2302 ( n254 , n505 , n3415 );
    and g2303 ( n1581 , n1037 , n1925 );
    or g2304 ( n2008 , n1688 , n1702 );
    or g2305 ( n1824 , n2955 , n1916 );
    and g2306 ( n780 , n514 , n1123 );
    nor g2307 ( n377 , n2683 , n693 );
    or g2308 ( n2534 , n928 , n2817 );
    or g2309 ( n2708 , n899 , n441 );
    nor g2310 ( n436 , n1557 , n2124 );
    nor g2311 ( n1920 , n2429 , n3454 );
    and g2312 ( n3729 , n962 , n2194 );
    not g2313 ( n2162 , n197 );
    and g2314 ( n3093 , n338 , n1285 );
    and g2315 ( n2964 , n2368 , n1866 );
    or g2316 ( n3894 , n263 , n1554 );
    and g2317 ( n1963 , n479 , n3877 );
    or g2318 ( n3050 , n3867 , n3903 );
    nor g2319 ( n2909 , n3467 , n2937 );
    or g2320 ( n2381 , n2767 , n3025 );
    or g2321 ( n3877 , n3279 , n3903 );
    or g2322 ( n828 , n2482 , n3887 );
    not g2323 ( n1604 , n2606 );
    or g2324 ( n1278 , n3424 , n2623 );
    and g2325 ( n1837 , n1718 , n3731 );
    or g2326 ( n372 , n15 , n3466 );
    or g2327 ( n2975 , n269 , n1463 );
    nor g2328 ( n166 , n3459 , n2402 );
    or g2329 ( n1984 , n2052 , n831 );
    and g2330 ( n3358 , n3489 , n2966 );
    or g2331 ( n1028 , n1563 , n2709 );
    not g2332 ( n2747 , n507 );
    or g2333 ( n3218 , n851 , n1346 );
    or g2334 ( n1323 , n1926 , n394 );
    or g2335 ( n3070 , n1006 , n2940 );
    or g2336 ( n2208 , n1814 , n1554 );
    not g2337 ( n1572 , n584 );
    nor g2338 ( n3470 , n3724 , n3377 );
    or g2339 ( n711 , n2195 , n3692 );
    and g2340 ( n1979 , n3286 , n3613 );
    or g2341 ( n2849 , n180 , n1101 );
    or g2342 ( n3325 , n1659 , n2495 );
    nor g2343 ( n2965 , n1568 , n2874 );
    or g2344 ( n357 , n3582 , n2673 );
    not g2345 ( n946 , n3045 );
    not g2346 ( n3707 , n3379 );
    and g2347 ( n3095 , n1344 , n2011 );
    nor g2348 ( n692 , n1917 , n2959 );
    buf g2349 ( n761 , n3887 );
    and g2350 ( n1162 , n2262 , n2470 );
    and g2351 ( n2405 , n2934 , n201 );
    and g2352 ( n1156 , n2319 , n3481 );
    or g2353 ( n3719 , n729 , n1232 );
    or g2354 ( n3551 , n317 , n3276 );
    and g2355 ( n3264 , n3164 , n3268 );
    not g2356 ( n1711 , n145 );
    and g2357 ( n1311 , n1502 , n1644 );
    not g2358 ( n1759 , n1113 );
    or g2359 ( n2173 , n952 , n781 );
    buf g2360 ( n2769 , n2625 );
    and g2361 ( n1755 , n2625 , n145 );
    and g2362 ( n3653 , n3281 , n3176 );
    not g2363 ( n3762 , n1046 );
    nor g2364 ( n1336 , n3763 , n3804 );
    and g2365 ( n3144 , n3455 , n2257 );
    not g2366 ( n1674 , n3303 );
    not g2367 ( n2537 , n3416 );
    or g2368 ( n3226 , n2949 , n2009 );
    or g2369 ( n563 , n3240 , n1523 );
    or g2370 ( n3710 , n1062 , n3272 );
    nor g2371 ( n3407 , n786 , n1361 );
    or g2372 ( n2790 , n1867 , n619 );
    or g2373 ( n1260 , n2841 , n305 );
    nor g2374 ( n3706 , n2667 , n1190 );
    not g2375 ( n3232 , n1778 );
    and g2376 ( n1478 , n496 , n1700 );
    not g2377 ( n2763 , n1862 );
    and g2378 ( n2744 , n1299 , n388 );
    nor g2379 ( n1477 , n3852 , n2793 );
    and g2380 ( n3874 , n2769 , n650 );
    not g2381 ( n2321 , n1470 );
    and g2382 ( n2646 , n3352 , n103 );
    nor g2383 ( n2754 , n1310 , n2913 );
    and g2384 ( n1658 , n1173 , n2805 );
    and g2385 ( n1704 , n3650 , n3809 );
    nor g2386 ( n2484 , n2919 , n3683 );
    and g2387 ( n3443 , n3072 , n1237 );
    and g2388 ( n876 , n1883 , n2187 );
    or g2389 ( n1245 , n847 , n1848 );
    and g2390 ( n353 , n161 , n2247 );
    or g2391 ( n670 , n1737 , n3141 );
    and g2392 ( n2825 , n2730 , n3708 );
    or g2393 ( n327 , n228 , n1864 );
    not g2394 ( n663 , n2297 );
    or g2395 ( n3709 , n1329 , n2797 );
    or g2396 ( n2356 , n2628 , n195 );
    or g2397 ( n1466 , n91 , n571 );
    or g2398 ( n1404 , n3016 , n509 );
    buf g2399 ( n3910 , n1026 );
    not g2400 ( n3057 , n3379 );
    and g2401 ( n2250 , n2387 , n71 );
    not g2402 ( n3664 , n739 );
    or g2403 ( n2554 , n676 , n2819 );
    nor g2404 ( n2110 , n3901 , n2542 );
    or g2405 ( n626 , n109 , n3058 );
    or g2406 ( n2153 , n799 , n3778 );
    and g2407 ( n3159 , n249 , n409 );
    nor g2408 ( n2035 , n2418 , n3906 );
    not g2409 ( n3520 , n1757 );
    or g2410 ( n1451 , n2920 , n2835 );
    nor g2411 ( n520 , n3538 , n670 );
    not g2412 ( n2944 , n1719 );
    or g2413 ( n1529 , n2113 , n3674 );
    nor g2414 ( n3632 , n229 , n3453 );
    or g2415 ( n205 , n1673 , n3674 );
    nor g2416 ( n1380 , n3658 , n2101 );
    not g2417 ( n1115 , n2210 );
    or g2418 ( n3021 , n1733 , n2614 );
    not g2419 ( n2062 , n3379 );
    not g2420 ( n513 , n556 );
    and g2421 ( n3094 , n110 , n1577 );
    or g2422 ( n1636 , n1392 , n3015 );
    not g2423 ( n3161 , n3713 );
    nor g2424 ( n1502 , n2507 , n1803 );
    and g2425 ( n2426 , n1058 , n1013 );
    and g2426 ( n3071 , n51 , n739 );
    or g2427 ( n262 , n3186 , n2836 );
    or g2428 ( n2483 , n45 , n367 );
    and g2429 ( n1528 , n2401 , n2927 );
    or g2430 ( n2953 , n1724 , n2178 );
    nor g2431 ( n2054 , n3402 , n3627 );
    or g2432 ( n1590 , n503 , n380 );
    and g2433 ( n2687 , n3579 , n3249 );
    and g2434 ( n1183 , n674 , n2074 );
    or g2435 ( n2634 , n2995 , n1620 );
    nor g2436 ( n667 , n3422 , n1554 );
    and g2437 ( n252 , n1525 , n2915 );
    and g2438 ( n748 , n3066 , n3065 );
    or g2439 ( n2526 , n1954 , n3449 );
    or g2440 ( n2315 , n3488 , n2454 );
    and g2441 ( n2547 , n741 , n828 );
    and g2442 ( n1055 , n2842 , n1700 );
    or g2443 ( n221 , n1435 , n1212 );
    not g2444 ( n502 , n3213 );
    and g2445 ( n98 , n1193 , n1130 );
    and g2446 ( n3037 , n2864 , n1015 );
    and g2447 ( n1046 , n3910 , n571 );
    not g2448 ( n2595 , n1865 );
    and g2449 ( n64 , n437 , n3653 );
    or g2450 ( n1297 , n905 , n2726 );
    not g2451 ( n271 , n3887 );
    and g2452 ( n1007 , n3325 , n1034 );
    or g2453 ( n3492 , n2488 , n1772 );
    or g2454 ( n3563 , n1017 , n2407 );
    or g2455 ( n2233 , n41 , n320 );
    or g2456 ( n265 , n1063 , n571 );
    nor g2457 ( n1600 , n304 , n2769 );
    and g2458 ( n1186 , n504 , n3354 );
    nor g2459 ( n13 , n1546 , n3404 );
    and g2460 ( n2612 , n1284 , n2087 );
    or g2461 ( n635 , n2282 , n2932 );
    not g2462 ( n1388 , n2946 );
    or g2463 ( n2496 , n1013 , n3692 );
    or g2464 ( n3845 , n2194 , n3689 );
    or g2465 ( n3646 , n690 , n662 );
    or g2466 ( n3498 , n1873 , n2996 );
    and g2467 ( n3005 , n3316 , n729 );
    and g2468 ( n280 , n3594 , n660 );
    nor g2469 ( n3798 , n3080 , n3371 );
    not g2470 ( n1644 , n1177 );
    or g2471 ( n55 , n1428 , n1898 );
    or g2472 ( n3251 , n373 , n2800 );
    nor g2473 ( n3163 , n1417 , n1909 );
    or g2474 ( n122 , n3048 , n831 );
    and g2475 ( n3912 , n3187 , n1230 );
    and g2476 ( n2915 , n911 , n1786 );
    nor g2477 ( n2999 , n2043 , n2351 );
    or g2478 ( n3173 , n64 , n599 );
    not g2479 ( n3599 , n3732 );
    and g2480 ( n2308 , n2107 , n904 );
    or g2481 ( n2159 , n2417 , n3098 );
    and g2482 ( n3278 , n3079 , n1841 );
    nor g2483 ( n3829 , n2731 , n1535 );
    not g2484 ( n1445 , n2289 );
    and g2485 ( n2855 , n3436 , n3226 );
    or g2486 ( n2169 , n1604 , n1431 );
    and g2487 ( n1700 , n3842 , n1797 );
    and g2488 ( n1176 , n547 , n757 );
    and g2489 ( n364 , n2689 , n2636 );
    not g2490 ( n943 , n3065 );
    and g2491 ( n456 , n3487 , n2416 );
    or g2492 ( n809 , n3840 , n3762 );
    not g2493 ( n471 , n2744 );
    or g2494 ( n782 , n1179 , n831 );
    not g2495 ( n3271 , n1062 );
    and g2496 ( n465 , n3483 , n3181 );
    and g2497 ( n2778 , n2830 , n3305 );
    buf g2498 ( n463 , n3548 );
    and g2499 ( n894 , n3483 , n1780 );
    and g2500 ( n3875 , n947 , n2089 );
    and g2501 ( n3000 , n1164 , n914 );
    nor g2502 ( n207 , n2157 , n1376 );
    or g2503 ( n1158 , n165 , n3742 );
    or g2504 ( n906 , n2303 , n717 );
    and g2505 ( n2417 , n1893 , n1899 );
    or g2506 ( n1540 , n1183 , n2802 );
    and g2507 ( n1171 , n437 , n533 );
    and g2508 ( n1181 , n2350 , n3860 );
    nor g2509 ( n1714 , n0 , n2140 );
    nor g2510 ( n2283 , n969 , n1159 );
    and g2511 ( n2571 , n427 , n848 );
    and g2512 ( n1410 , n3786 , n2061 );
    and g2513 ( n881 , n2737 , n3648 );
    and g2514 ( n2935 , n2306 , n1091 );
    or g2515 ( n2497 , n823 , n2528 );
    or g2516 ( n2598 , n837 , n3330 );
    not g2517 ( n3230 , n1873 );
    or g2518 ( n3305 , n1679 , n1978 );
    not g2519 ( n3583 , n462 );
    and g2520 ( n837 , n2907 , n2052 );
    not g2521 ( n3486 , n3379 );
    and g2522 ( n30 , n3483 , n1279 );
    or g2523 ( n3778 , n449 , n2172 );
    or g2524 ( n983 , n2193 , n30 );
    and g2525 ( n2878 , n3212 , n2710 );
    not g2526 ( n2992 , n804 );
    or g2527 ( n2264 , n2589 , n1188 );
    and g2528 ( n1769 , n1138 , n1988 );
    or g2529 ( n1122 , n746 , n2174 );
    and g2530 ( n708 , n2337 , n1269 );
    nor g2531 ( n1941 , n3857 , n1695 );
    or g2532 ( n3576 , n936 , n1523 );
    and g2533 ( n1997 , n1486 , n308 );
    and g2534 ( n3414 , n1446 , n3219 );
    or g2535 ( n2221 , n3400 , n3516 );
    or g2536 ( n1381 , n7 , n684 );
    nor g2537 ( n2171 , n3054 , n3637 );
    not g2538 ( n2343 , n3653 );
    and g2539 ( n1669 , n2413 , n3061 );
    and g2540 ( n3826 , n859 , n2512 );
    or g2541 ( n2682 , n2353 , n2543 );
    buf g2542 ( n571 , n3887 );
    not g2543 ( n3383 , n3376 );
    not g2544 ( n2816 , n3895 );
    or g2545 ( n2397 , n3828 , n2279 );
    or g2546 ( n512 , n566 , n374 );
    and g2547 ( n1285 , n1108 , n3495 );
    and g2548 ( n2823 , n3438 , n1332 );
    not g2549 ( n1993 , n703 );
    and g2550 ( n778 , n3419 , n3094 );
    not g2551 ( n2178 , n707 );
    nor g2552 ( n997 , n3614 , n1433 );
    not g2553 ( n258 , n3152 );
    or g2554 ( n3045 , n3889 , n2255 );
    nor g2555 ( n1788 , n1656 , n1706 );
    not g2556 ( n1854 , n2872 );
    not g2557 ( n3881 , n1773 );
    or g2558 ( n2635 , n1821 , n1898 );
    or g2559 ( n310 , n3236 , n3887 );
    or g2560 ( n3859 , n2938 , n1101 );
    nor g2561 ( n2735 , n1147 , n1401 );
    not g2562 ( n645 , n1977 );
    nor g2563 ( n3655 , n3221 , n222 );
    nor g2564 ( n2415 , n3882 , n611 );
    and g2565 ( n905 , n2625 , n752 );
    and g2566 ( n3256 , n2036 , n290 );
    nor g2567 ( n3211 , n1349 , n3317 );
    not g2568 ( n547 , n3860 );
    nor g2569 ( n2241 , n2784 , n814 );
    or g2570 ( n3841 , n473 , n1916 );
    or g2571 ( n3371 , n2897 , n3406 );
    nor g2572 ( n36 , n3890 , n1270 );
    and g2573 ( n2155 , n387 , n3463 );
    or g2574 ( n3615 , n1507 , n1302 );
    not g2575 ( n3715 , n1265 );
    not g2576 ( n715 , n2358 );
    and g2577 ( n3690 , n213 , n3287 );
    nor g2578 ( n2795 , n3888 , n1787 );
    not g2579 ( n2329 , n2529 );
    not g2580 ( n3143 , n2533 );
    or g2581 ( n3744 , n2786 , n2389 );
    and g2582 ( n250 , n892 , n3020 );
    or g2583 ( n2146 , n2899 , n3289 );
    and g2584 ( n2396 , n3321 , n2133 );
    or g2585 ( n2522 , n1454 , n220 );
    or g2586 ( n3267 , n2054 , n2826 );
    not g2587 ( n1090 , n1839 );
    or g2588 ( n1953 , n2866 , n603 );
    nor g2589 ( n3704 , n1552 , n3374 );
    or g2590 ( n3816 , n413 , n1916 );
    not g2591 ( n3505 , n3910 );
    nor g2592 ( n3222 , n3016 , n1510 );
    or g2593 ( n3464 , n10 , n3015 );
    or g2594 ( n2911 , n1018 , n3368 );
    and g2595 ( n1409 , n2798 , n2446 );
    and g2596 ( n3913 , n2129 , n3023 );
    nor g2597 ( n1705 , n2808 , n3299 );
    not g2598 ( n3348 , n3255 );
    nor g2599 ( n860 , n650 , n2772 );
    nor g2600 ( n2688 , n1442 , n1259 );
    not g2601 ( n1844 , n1789 );
    and g2602 ( n1885 , n224 , n2858 );
    not g2603 ( n405 , n3272 );
    and g2604 ( n3011 , n391 , n640 );
    not g2605 ( n1865 , n2625 );
    not g2606 ( n3490 , n3838 );
    and g2607 ( n2363 , n1208 , n3171 );
    and g2608 ( n1678 , n1916 , n2910 );
    nor g2609 ( n2450 , n1954 , n2065 );
    and g2610 ( n1745 , n1586 , n2644 );
    not g2611 ( n100 , n1809 );
    not g2612 ( n2683 , n801 );
    nor g2613 ( n2812 , n328 , n1752 );
    and g2614 ( n145 , n2517 , n2218 );
    or g2615 ( n1095 , n1145 , n3018 );
    and g2616 ( n561 , n2344 , n1323 );
    nor g2617 ( n3766 , n211 , n1975 );
    or g2618 ( n142 , n204 , n539 );
    and g2619 ( n1773 , n2201 , n934 );
    and g2620 ( n732 , n1302 , n1507 );
    or g2621 ( n1064 , n2784 , n1187 );
    not g2622 ( n1846 , n624 );
    and g2623 ( n683 , n725 , n1256 );
    not g2624 ( n2312 , n2672 );
    and g2625 ( n2006 , n702 , n857 );
    and g2626 ( n724 , n3179 , n2670 );
    or g2627 ( n404 , n1252 , n1493 );
    and g2628 ( n322 , n130 , n16 );
    not g2629 ( n1024 , n1576 );
    nor g2630 ( n737 , n1570 , n3849 );
    or g2631 ( n2021 , n1679 , n3466 );
    and g2632 ( n3701 , n1451 , n2843 );
    not g2633 ( n518 , n2706 );
    buf g2634 ( n1554 , n1026 );
    or g2635 ( n3748 , n854 , n3169 );
    nor g2636 ( n1355 , n3511 , n3853 );
    not g2637 ( n3533 , n1499 );
    and g2638 ( n1269 , n191 , n172 );
    or g2639 ( n907 , n3292 , n3191 );
    not g2640 ( n701 , n754 );
    and g2641 ( n2268 , n556 , n3042 );
    not g2642 ( n199 , n189 );
    or g2643 ( n2839 , n1720 , n1551 );
    nor g2644 ( n83 , n3422 , n1495 );
    or g2645 ( n2715 , n1419 , n3132 );
    and g2646 ( n3362 , n2817 , n928 );
    and g2647 ( n3392 , n3615 , n3226 );
    and g2648 ( n2570 , n2769 , n2666 );
    and g2649 ( n588 , n882 , n652 );
    nor g2650 ( n686 , n2048 , n1520 );
    and g2651 ( n1913 , n3780 , n2491 );
    and g2652 ( n1578 , n3483 , n869 );
    and g2653 ( n1999 , n645 , n2087 );
    not g2654 ( n2439 , n178 );
    and g2655 ( n176 , n1232 , n729 );
    nor g2656 ( n3073 , n2436 , n3505 );
    and g2657 ( n2671 , n266 , n345 );
    nor g2658 ( n853 , n890 , n3898 );
    and g2659 ( n2549 , n367 , n3901 );
    not g2660 ( n2817 , n359 );
    or g2661 ( n3281 , n1925 , n1916 );
    nor g2662 ( n560 , n2725 , n633 );
    or g2663 ( n1266 , n1982 , n134 );
    nor g2664 ( n689 , n1506 , n2370 );
    or g2665 ( n3205 , n924 , n1916 );
    or g2666 ( n1857 , n2355 , n2936 );
    or g2667 ( n1004 , n219 , n3505 );
    or g2668 ( n2190 , n3267 , n552 );
    or g2669 ( n2128 , n3634 , n2971 );
    not g2670 ( n2256 , n2569 );
    and g2671 ( n2892 , n2723 , n2851 );
    or g2672 ( n2990 , n2358 , n3169 );
    and g2673 ( n2882 , n2080 , n3437 );
    or g2674 ( n2192 , n1056 , n1591 );
    nor g2675 ( n131 , n3144 , n1744 );
    and g2676 ( n832 , n2540 , n1466 );
    not g2677 ( n1828 , n477 );
    or g2678 ( n2559 , n2372 , n2824 );
    nor g2679 ( n3003 , n762 , n2716 );
    or g2680 ( n1492 , n886 , n908 );
    and g2681 ( n289 , n1224 , n15 );
    or g2682 ( n3013 , n1332 , n3910 );
    or g2683 ( n2447 , n1691 , n822 );
    and g2684 ( n1687 , n2753 , n1681 );
    not g2685 ( n3786 , n293 );
    and g2686 ( n2310 , n1893 , n2687 );
    buf g2687 ( n1916 , n1188 );
    or g2688 ( n172 , n3155 , n3692 );
    or g2689 ( n811 , n2004 , n2421 );
    and g2690 ( n3428 , n1121 , n27 );
    nor g2691 ( n3882 , n2166 , n1390 );
    and g2692 ( n486 , n476 , n176 );
    or g2693 ( n1830 , n3258 , n2372 );
    or g2694 ( n135 , n2045 , n3108 );
    and g2695 ( n1532 , n3893 , n2463 );
    and g2696 ( n3457 , n1081 , n3772 );
    nor g2697 ( n427 , n1071 , n3768 );
    or g2698 ( n1550 , n1688 , n3015 );
    and g2699 ( n2515 , n403 , n2865 );
    not g2700 ( n183 , n448 );
    and g2701 ( n1203 , n2221 , n1423 );
    or g2702 ( n2132 , n2437 , n509 );
    and g2703 ( n2579 , n2018 , n1470 );
    buf g2704 ( n336 , n3548 );
    or g2705 ( n985 , n1968 , n1196 );
    not g2706 ( n3902 , n1434 );
    or g2707 ( n2104 , n2213 , n2016 );
    nor g2708 ( n2303 , n3376 , n660 );
    and g2709 ( n1358 , n3868 , n965 );
    nor g2710 ( n1097 , n1703 , n2905 );
    and g2711 ( n2454 , n287 , n3895 );
    or g2712 ( n1108 , n3634 , n1898 );
    nor g2713 ( n2156 , n2987 , n3361 );
    nor g2714 ( n2326 , n486 , n79 );
    or g2715 ( n1014 , n112 , n3466 );
    or g2716 ( n3283 , n975 , n3822 );
    and g2717 ( n97 , n3769 , n2744 );
    or g2718 ( n1209 , n1710 , n2180 );
    and g2719 ( n3395 , n1076 , n2161 );
    or g2720 ( n2840 , n72 , n783 );
    or g2721 ( n865 , n3171 , n3449 );
    and g2722 ( n3253 , n2276 , n3588 );
    not g2723 ( n608 , n29 );
    nor g2724 ( n2792 , n240 , n430 );
    nor g2725 ( n3209 , n450 , n2909 );
    and g2726 ( n417 , n437 , n3040 );
    or g2727 ( n148 , n2722 , n3687 );
    not g2728 ( n1384 , n2297 );
    nor g2729 ( n407 , n1109 , n2444 );
    or g2730 ( n2440 , n1731 , n3583 );
    and g2731 ( n1374 , n3483 , n3862 );
    or g2732 ( n3129 , n3399 , n2607 );
    and g2733 ( n2378 , n277 , n2467 );
    or g2734 ( n2567 , n2205 , n343 );
    nor g2735 ( n806 , n579 , n2769 );
    nor g2736 ( n3550 , n909 , n2461 );
    nor g2737 ( n184 , n2918 , n769 );
    and g2738 ( n1547 , n2182 , n3190 );
    not g2739 ( n1840 , n915 );
    or g2740 ( n2883 , n2705 , n3466 );
    and g2741 ( n3340 , n3112 , n1044 );
    nor g2742 ( n3485 , n2597 , n3626 );
    and g2743 ( n2150 , n390 , n1348 );
    or g2744 ( n290 , n3189 , n2844 );
    nor g2745 ( n3243 , n268 , n267 );
    or g2746 ( n819 , n277 , n3351 );
    or g2747 ( n567 , n3712 , n3887 );
    not g2748 ( n203 , n467 );
    or g2749 ( n3176 , n3426 , n3153 );
    or g2750 ( n3495 , n1372 , n908 );
    and g2751 ( n2065 , n2760 , n1703 );
    and g2752 ( n2096 , n3483 , n855 );
    not g2753 ( n1052 , n1728 );
    nor g2754 ( n2807 , n3871 , n62 );
    not g2755 ( n3907 , n2946 );
    or g2756 ( n1878 , n2907 , n2823 );
    nor g2757 ( n232 , n3280 , n3196 );
    and g2758 ( n2234 , n2060 , n18 );
    and g2759 ( n3376 , n2132 , n153 );
    or g2760 ( n2805 , n2955 , n433 );
    or g2761 ( n1596 , n2260 , n3611 );
    and g2762 ( n3413 , n980 , n1672 );
    and g2763 ( n2674 , n1364 , n1637 );
    or g2764 ( n2269 , n82 , n996 );
    nor g2765 ( n3509 , n855 , n3106 );
    nor g2766 ( n3195 , n1615 , n831 );
    or g2767 ( n2428 , n3629 , n2844 );
    nor g2768 ( n2140 , n485 , n1709 );
    buf g2769 ( n467 , n2625 );
    and g2770 ( n255 , n437 , n693 );
    and g2771 ( n1457 , n501 , n1395 );
    nor g2772 ( n397 , n3226 , n213 );
    not g2773 ( n249 , n796 );
    nor g2774 ( n1850 , n3458 , n3592 );
    or g2775 ( n2368 , n3203 , n3910 );
    not g2776 ( n3769 , n2946 );
    nor g2777 ( n2451 , n2788 , n1131 );
    or g2778 ( n812 , n2792 , n841 );
    nor g2779 ( n2662 , n2820 , n2607 );
    not g2780 ( n568 , n2263 );
    or g2781 ( n431 , n2766 , n2145 );
    nor g2782 ( n1749 , n3429 , n3088 );
    not g2783 ( n2971 , n1372 );
    and g2784 ( n841 , n663 , n270 );
    or g2785 ( n141 , n2872 , n2996 );
    and g2786 ( n2640 , n870 , n96 );
    and g2787 ( n695 , n727 , n1565 );
    not g2788 ( n3627 , n1549 );
    not g2789 ( n323 , n1528 );
    or g2790 ( n3584 , n3109 , n2219 );
    nor g2791 ( n396 , n1972 , n3605 );
    not g2792 ( n790 , n321 );
    and g2793 ( n804 , n1014 , n1019 );
    not g2794 ( n816 , n386 );
    or g2795 ( n1945 , n459 , n1898 );
    not g2796 ( n1438 , n3048 );
    and g2797 ( n2750 , n3892 , n2305 );
    and g2798 ( n3396 , n2078 , n2574 );
    not g2799 ( n1100 , n1664 );
    or g2800 ( n2030 , n1178 , n3264 );
    and g2801 ( n2305 , n3748 , n950 );
    nor g2802 ( n3273 , n820 , n793 );
    or g2803 ( n3705 , n3152 , n3536 );
    nor g2804 ( n3183 , n1400 , n2893 );
    and g2805 ( n783 , n496 , n328 );
    not g2806 ( n1050 , n3887 );
    not g2807 ( n1683 , n1780 );
    and g2808 ( n2597 , n2143 , n358 );
    nor g2809 ( n2689 , n1913 , n2380 );
    or g2810 ( n2228 , n1924 , n1474 );
    or g2811 ( n174 , n356 , n23 );
    or g2812 ( n1048 , n1053 , n21 );
    nor g2813 ( n2314 , n18 , n1078 );
    nor g2814 ( n3794 , n1395 , n501 );
    and g2815 ( n2335 , n2235 , n3227 );
    or g2816 ( n3355 , n3767 , n1483 );
    and g2817 ( n654 , n3404 , n1507 );
    or g2818 ( n932 , n3412 , n2612 );
    or g2819 ( n1 , n1336 , n1600 );
    not g2820 ( n1535 , n73 );
    not g2821 ( n333 , n3423 );
    not g2822 ( n1847 , n422 );
    or g2823 ( n2370 , n1759 , n1307 );
    nor g2824 ( n378 , n3815 , n612 );
    or g2825 ( n2248 , n2149 , n1223 );
    not g2826 ( n222 , n3379 );
    and g2827 ( n3367 , n3575 , n3718 );
    and g2828 ( n3822 , n2611 , n2173 );
    and g2829 ( n1883 , n2675 , n1191 );
    or g2830 ( n719 , n1291 , n1961 );
    not g2831 ( n2785 , n3261 );
    not g2832 ( n653 , n337 );
    nor g2833 ( n47 , n2640 , n3554 );
    not g2834 ( n2441 , n3382 );
    or g2835 ( n2053 , n413 , n979 );
    not g2836 ( n1446 , n3818 );
    and g2837 ( n447 , n1935 , n2869 );
    or g2838 ( n873 , n3591 , n2342 );
    not g2839 ( n2316 , n2133 );
    and g2840 ( n469 , n1887 , n3599 );
    nor g2841 ( n2118 , n678 , n1055 );
    nor g2842 ( n1325 , n1648 , n1647 );
    nor g2843 ( n3908 , n3752 , n1119 );
    not g2844 ( n1091 , n2670 );
    and g2845 ( n1439 , n3719 , n3004 );
    and g2846 ( n3667 , n2209 , n469 );
    and g2847 ( n1120 , n3483 , n77 );
    or g2848 ( n2285 , n73 , n1916 );
    and g2849 ( n2372 , n1246 , n2116 );
    not g2850 ( n3128 , n3319 );
    or g2851 ( n1038 , n4 , n2298 );
    and g2852 ( n1345 , n3483 , n1969 );
    or g2853 ( n1735 , n397 , n778 );
    not g2854 ( n2176 , n2774 );
    buf g2855 ( n334 , n3548 );
    and g2856 ( n1060 , n1024 , n1144 );
    nor g2857 ( n2815 , n1176 , n2390 );
    nor g2858 ( n450 , n2334 , n3620 );
    buf g2859 ( n3169 , n1694 );
    not g2860 ( n988 , n3034 );
    nor g2861 ( n3556 , n648 , n2320 );
    or g2862 ( n308 , n1049 , n3903 );
    or g2863 ( n3743 , n409 , n571 );
    or g2864 ( n3375 , n581 , n3827 );
    nor g2865 ( n3384 , n1063 , n594 );
    nor g2866 ( n2514 , n2911 , n2347 );
    or g2867 ( n2546 , n3730 , n2012 );
    and g2868 ( n3113 , n3246 , n362 );
    buf g2869 ( n1026 , n2607 );
    nor g2870 ( n2916 , n1539 , n3320 );
    and g2871 ( n3025 , n3200 , n1715 );
    or g2872 ( n3703 , n3780 , n2396 );
    or g2873 ( n482 , n2638 , n1916 );
    nor g2874 ( n3160 , n2026 , n67 );
    and g2875 ( n2338 , n3846 , n2613 );
    or g2876 ( n2359 , n703 , n3449 );
    or g2877 ( n3391 , n2992 , n90 );
    and g2878 ( n3009 , n1618 , n2686 );
    nor g2879 ( n3917 , n1088 , n3798 );
    nor g2880 ( n385 , n1331 , n635 );
    or g2881 ( n3042 , n3633 , n2548 );
    and g2882 ( n890 , n2418 , n1524 );
    and g2883 ( n987 , n2947 , n3757 );
    or g2884 ( n2284 , n1758 , n2996 );
    and g2885 ( n1043 , n124 , n2849 );
    nor g2886 ( n3424 , n623 , n3766 );
    or g2887 ( n3644 , n3754 , n1101 );
    and g2888 ( n3287 , n1614 , n1137 );
    and g2889 ( n3274 , n839 , n1792 );
    nor g2890 ( n2753 , n3493 , n3916 );
    and g2891 ( n1298 , n2747 , n1151 );
    nor g2892 ( n2082 , n3708 , n2730 );
    and g2893 ( n614 , n2696 , n3613 );
    and g2894 ( n3898 , n85 , n242 );
    or g2895 ( n3669 , n29 , n3887 );
    or g2896 ( n3295 , n3873 , n3015 );
    or g2897 ( n1767 , n162 , n3293 );
    or g2898 ( n416 , n885 , n942 );
    not g2899 ( n532 , n3215 );
    not g2900 ( n3896 , n2087 );
    and g2901 ( n3781 , n132 , n3198 );
    nor g2902 ( n3870 , n3119 , n3158 );
    nor g2903 ( n3194 , n1060 , n1795 );
    nor g2904 ( n3311 , n3726 , n32 );
    or g2905 ( n488 , n1229 , n831 );
    or g2906 ( n248 , n477 , n3887 );
    or g2907 ( n2838 , n1314 , n3466 );
    or g2908 ( n162 , n1571 , n1653 );
    nor g2909 ( n2444 , n34 , n3049 );
    not g2910 ( n318 , n1295 );
    nor g2911 ( n1401 , n1200 , n2957 );
    or g2912 ( n214 , n720 , n908 );
    or g2913 ( n1129 , n3398 , n2609 );
    or g2914 ( n3868 , n3648 , n3449 );
    or g2915 ( n481 , n1221 , n3365 );
    and g2916 ( n578 , n1753 , n774 );
    nor g2917 ( n522 , n2066 , n978 );
    not g2918 ( n1134 , n3219 );
    nor g2919 ( n2291 , n2492 , n1156 );
    or g2920 ( n2366 , n1925 , n1037 );
    and g2921 ( n78 , n3328 , n1933 );
    not g2922 ( n665 , n3887 );
    buf g2923 ( n3015 , n2062 );
    and g2924 ( n2070 , n1251 , n42 );
    and g2925 ( n3468 , n1261 , n1244 );
    not g2926 ( n1213 , n2461 );
    or g2927 ( n1294 , n1259 , n1970 );
    and g2928 ( n2508 , n3763 , n1665 );
    or g2929 ( n1712 , n1790 , n1973 );
    nor g2930 ( n847 , n282 , n1818 );
    or g2931 ( n2630 , n3600 , n2996 );
    not g2932 ( n3047 , n3530 );
    not g2933 ( n2810 , n3379 );
    not g2934 ( n2720 , n570 );
    and g2935 ( n2244 , n3483 , n3219 );
    and g2936 ( n597 , n2228 , n1095 );
    nor g2937 ( n2419 , n337 , n3297 );
    and g2938 ( n1542 , n2040 , n3074 );
    and g2939 ( n1471 , n2895 , n3750 );
    nor g2940 ( n2126 , n903 , n2531 );
    buf g2941 ( n3887 , n1601 );
    not g2942 ( n868 , n1086 );
    and g2943 ( n485 , n2697 , n3358 );
    and g2944 ( n2904 , n3715 , n3253 );
    nor g2945 ( n2854 , n3349 , n2769 );
    and g2946 ( n3697 , n113 , n529 );
    not g2947 ( n88 , n3253 );
    or g2948 ( n3899 , n2144 , n1188 );
    or g2949 ( n1523 , n1093 , n1181 );
    and g2950 ( n27 , n3753 , n2214 );
    not g2951 ( n2060 , n2768 );
    not g2952 ( n2521 , n2709 );
    and g2953 ( n740 , n3284 , n2695 );
    nor g2954 ( n202 , n3410 , n2605 );
    or g2955 ( n2344 , n2997 , n755 );
    nor g2956 ( n3525 , n3022 , n360 );
    not g2957 ( n3062 , n1548 );
    and g2958 ( n3858 , n856 , n2672 );
    and g2959 ( n2193 , n2769 , n3344 );
    or g2960 ( n384 , n2014 , n2451 );
    or g2961 ( n432 , n314 , n1858 );
    and g2962 ( n3080 , n3741 , n1542 );
    not g2963 ( n1974 , n568 );
    and g2964 ( n1267 , n206 , n3747 );
    and g2965 ( n1667 , n3791 , n1957 );
    or g2966 ( n3087 , n1888 , n1560 );
    not g2967 ( n2263 , n2625 );
    nor g2968 ( n760 , n2880 , n2931 );
    nor g2969 ( n314 , n3571 , n2280 );
    not g2970 ( n2530 , n2738 );
    and g2971 ( n3759 , n2620 , n1579 );
    and g2972 ( n3699 , n2831 , n2051 );
    nor g2973 ( n494 , n605 , n2732 );
    nor g2974 ( n589 , n858 , n3032 );
    nor g2975 ( n969 , n3678 , n1206 );
    or g2976 ( n163 , n776 , n416 );
    nor g2977 ( n1053 , n1314 , n444 );
    nor g2978 ( n1496 , n863 , n468 );
    and g2979 ( n41 , n437 , n2253 );
    and g2980 ( n23 , n3123 , n3805 );
    or g2981 ( n3603 , n628 , n3008 );
    nor g2982 ( n2395 , n848 , n1552 );
    or g2983 ( n616 , n361 , n683 );
    or g2984 ( n274 , n456 , n2307 );
    or g2985 ( n730 , n1178 , n3169 );
    or g2986 ( n110 , n3097 , n2996 );
    or g2987 ( n3442 , n1764 , n1677 );
    nor g2988 ( n324 , n2647 , n2275 );
    and g2989 ( n1399 , n3246 , n2215 );
    not g2990 ( n769 , n3379 );
    not g2991 ( n3139 , n2625 );
    or g2992 ( n3249 , n928 , n3015 );
    or g2993 ( n480 , n561 , n2581 );
    or g2994 ( n558 , n2825 , n2688 );
    nor g2995 ( n3369 , n3269 , n767 );
    or g2996 ( n137 , n335 , n884 );
    or g2997 ( n2969 , n3606 , n921 );
    and g2998 ( n1677 , n1189 , n743 );
    or g2999 ( n574 , n1930 , n2339 );
    and g3000 ( n1166 , n1563 , n1347 );
    nor g3001 ( n3214 , n2240 , n1192 );
    not g3002 ( n2601 , n2443 );
    nor g3003 ( n2009 , n71 , n2032 );
    and g3004 ( n1972 , n532 , n2189 );
    nor g3005 ( n2610 , n3477 , n1554 );
    or g3006 ( n3880 , n3569 , n355 );
    or g3007 ( n543 , n790 , n3884 );
    not g3008 ( n150 , n842 );
    or g3009 ( n2069 , n1253 , n1101 );
    and g3010 ( n3695 , n3288 , n695 );
    or g3011 ( n9 , n1126 , n1685 );
    not g3012 ( n2330 , n1618 );
    not g3013 ( n1058 , n1015 );
    nor g3014 ( n1657 , n1886 , n251 );
    or g3015 ( n2783 , n1904 , n2604 );
    or g3016 ( n3796 , n303 , n3887 );
    or g3017 ( n84 , n2722 , n908 );
    and g3018 ( n1695 , n2476 , n1914 );
    nor g3019 ( n3089 , n766 , n1973 );
    nor g3020 ( n1561 , n3873 , n3785 );
    or g3021 ( n3336 , n1650 , n212 );
    and g3022 ( n3356 , n454 , n2858 );
    and g3023 ( n1421 , n706 , n1180 );
    and g3024 ( n1307 , n468 , n863 );
    and g3025 ( n1530 , n3647 , n2516 );
    or g3026 ( n592 , n2262 , n521 );
    and g3027 ( n1725 , n3046 , n1524 );
    not g3028 ( n1637 , n598 );
    or g3029 ( n3696 , n1948 , n1722 );
    nor g3030 ( n2733 , n1426 , n833 );
    or g3031 ( n2707 , n1426 , n574 );
    not g3032 ( n2906 , n747 );
    nor g3033 ( n3857 , n3061 , n1387 );
    and g3034 ( n2348 , n2970 , n2868 );
    and g3035 ( n3312 , n1859 , n2672 );
    or g3036 ( n1029 , n1216 , n1916 );
    and g3037 ( n3834 , n3483 , n2868 );
    nor g3038 ( n3406 , n564 , n25 );
    not g3039 ( n1281 , n516 );
    or g3040 ( n3458 , n3456 , n376 );
    and g3041 ( n2639 , n502 , n3224 );
    not g3042 ( n2765 , n43 );
    and g3043 ( n3091 , n2538 , n1378 );
    nor g3044 ( n2423 , n1833 , n3888 );
    or g3045 ( n2259 , n3808 , n3357 );
    not g3046 ( n3053 , n2918 );
    or g3047 ( n1538 , n3258 , n1898 );
    and g3048 ( n212 , n600 , n2915 );
    not g3049 ( n3052 , n467 );
    or g3050 ( n1935 , n1308 , n3239 );
    and g3051 ( n3679 , n920 , n3285 );
    and g3052 ( n3306 , n3433 , n3443 );
    or g3053 ( n3452 , n2978 , n1748 );
    and g3054 ( n464 , n1421 , n3772 );
    nor g3055 ( n1419 , n1803 , n3525 );
    and g3056 ( n354 , n3483 , n242 );
    nor g3057 ( n1835 , n2818 , n3483 );
    and g3058 ( n1907 , n1422 , n2453 );
    nor g3059 ( n2420 , n322 , n1820 );
    buf g3060 ( n2625 , n2364 );
    or g3061 ( n1308 , n3315 , n1497 );
    or g3062 ( n2504 , n838 , n3692 );
    or g3063 ( n3277 , n1082 , n3442 );
    not g3064 ( n2127 , n495 );
    and g3065 ( n3096 , n3721 , n2862 );
    or g3066 ( n3154 , n2999 , n440 );
    buf g3067 ( n1268 , n3548 );
    or g3068 ( n3510 , n2658 , n509 );
    or g3069 ( n2988 , n1393 , n1916 );
    and g3070 ( n3199 , n2574 , n2710 );
    and g3071 ( n167 , n3018 , n1145 );
    or g3072 ( n1949 , n43 , n1207 );
    or g3073 ( n3044 , n1576 , n1188 );
    and g3074 ( n1969 , n1521 , n3408 );
    nor g3075 ( n1189 , n2059 , n3214 );
    or g3076 ( n3507 , n3870 , n607 );
    or g3077 ( n40 , n1485 , n194 );
    nor g3078 ( n2513 , n3283 , n2752 );
    or g3079 ( n124 , n3643 , n1188 );
    or g3080 ( n2887 , n1801 , n1350 );
    or g3081 ( n69 , n294 , n1652 );
    or g3082 ( n2677 , n3772 , n1101 );
    nor g3083 ( n994 , n1088 , n1220 );
    not g3084 ( n2018 , n2213 );
    nor g3085 ( n2553 , n3387 , n1893 );
    not g3086 ( n1386 , n3351 );
    or g3087 ( n3309 , n2194 , n962 );
    and g3088 ( n1602 , n3692 , n818 );
    or g3089 ( n2540 , n438 , n3169 );
    not g3090 ( n3738 , n858 );
    and g3091 ( n1414 , n2845 , n804 );
    or g3092 ( n2814 , n770 , n1554 );
    nor g3093 ( n2365 , n66 , n1469 );
    not g3094 ( n2371 , n2103 );
    or g3095 ( n2374 , n772 , n289 );
    nor g3096 ( n1227 , n2922 , n1203 );
    or g3097 ( n2568 , n565 , n3482 );
    or g3098 ( n1198 , n1114 , n1115 );
    or g3099 ( n2657 , n331 , n3863 );
    nor g3100 ( n1820 , n2876 , n2365 );
    and g3101 ( n2079 , n175 , n2224 );
    or g3102 ( n3172 , n2053 , n3714 );
    and g3103 ( n317 , n2625 , n3911 );
    not g3104 ( n1563 , n601 );
    nor g3105 ( n1819 , n2597 , n203 );
    or g3106 ( n272 , n589 , n1273 );
    nor g3107 ( n1584 , n1381 , n143 );
    not g3108 ( n1321 , n762 );
    and g3109 ( n3846 , n3012 , n3878 );
    and g3110 ( n3552 , n3560 , n2848 );
    and g3111 ( n2581 , n2269 , n57 );
    or g3112 ( n2913 , n1931 , n1175 );
    not g3113 ( n51 , n2099 );
    not g3114 ( n634 , n1623 );
    and g3115 ( n1250 , n3479 , n1947 );
    and g3116 ( n3649 , n369 , n3621 );
    not g3117 ( n3764 , n1184 );
    nor g3118 ( n618 , n1969 , n723 );
    not g3119 ( n3262 , n3366 );
    and g3120 ( n2349 , n3641 , n1707 );
    or g3121 ( n235 , n2684 , n2096 );
    nor g3122 ( n658 , n1296 , n3715 );
    and g3123 ( n1012 , n2177 , n2215 );
    or g3124 ( n1614 , n2222 , n3466 );
    not g3125 ( n2940 , n2055 );
    not g3126 ( n3672 , n844 );
    or g3127 ( n2721 , n1766 , n3742 );
    and g3128 ( n3181 , n3149 , n2403 );
    not g3129 ( n1566 , n3810 );
    and g3130 ( n2003 , n1209 , n500 );
    or g3131 ( n749 , n3586 , n1877 );
    or g3132 ( n2352 , n1242 , n2782 );
    or g3133 ( n1904 , n3388 , n3855 );
    and g3134 ( n3682 , n2832 , n3883 );
    or g3135 ( n1105 , n1835 , n1607 );
    not g3136 ( n3417 , n2946 );
    not g3137 ( n2939 , n2026 );
    nor g3138 ( n389 , n1226 , n3216 );
    or g3139 ( n1826 , n2787 , n3413 );
    nor g3140 ( n231 , n76 , n2600 );
    and g3141 ( n1431 , n868 , n101 );
    or g3142 ( n2561 , n443 , n3356 );
    and g3143 ( n2290 , n3062 , n2445 );
    not g3144 ( n331 , n3629 );
    or g3145 ( n3225 , n2035 , n1725 );
    or g3146 ( n1884 , n1233 , n3170 );
    and g3147 ( n2480 , n3719 , n22 );
    or g3148 ( n346 , n3195 , n3771 );
    or g3149 ( n531 , n1065 , n354 );
    and g3150 ( n989 , n2387 , n1537 );
    and g3151 ( n223 , n3274 , n2066 );
    or g3152 ( n2786 , n3854 , n1698 );
    or g3153 ( n266 , n3227 , n2235 );
    and g3154 ( n1515 , n253 , n2305 );
    and g3155 ( n1872 , n453 , n2400 );
    not g3156 ( n2525 , n3287 );
    and g3157 ( n3523 , n3280 , n3862 );
    and g3158 ( n1770 , n2321 , n2213 );
    nor g3159 ( n2627 , n298 , n412 );
    or g3160 ( n3617 , n1661 , n2112 );
    or g3161 ( n3789 , n1841 , n3449 );
    or g3162 ( n1660 , n2728 , n708 );
    or g3163 ( n3775 , n984 , n2996 );
    and g3164 ( n3609 , n1752 , n328 );
    not g3165 ( n3828 , n1559 );
    or g3166 ( n2134 , n775 , n571 );
    or g3167 ( n1555 , n777 , n1444 );
    and g3168 ( n367 , n2664 , n179 );
    or g3169 ( n2833 , n3494 , n2108 );
    or g3170 ( n188 , n3809 , n1916 );
    nor g3171 ( n2605 , n542 , n1856 );
    or g3172 ( n1476 , n3713 , n1207 );
    or g3173 ( n1261 , n2121 , n3910 );
    or g3174 ( n2871 , n3300 , n3254 );
    or g3175 ( n2843 , n3107 , n2295 );
    and g3176 ( n2868 , n865 , n2468 );
    nor g3177 ( n3254 , n2508 , n686 );
    or g3178 ( n2011 , n3819 , n1101 );
    nor g3179 ( n3206 , n2070 , n3350 );
    or g3180 ( n161 , n1248 , n156 );
    nor g3181 ( n2186 , n1805 , n1870 );
    not g3182 ( n2084 , n1179 );
    and g3183 ( n875 , n3317 , n3618 );
    or g3184 ( n950 , n2449 , n761 );
    and g3185 ( n2058 , n2771 , n1022 );
    nor g3186 ( n3844 , n1066 , n626 );
    or g3187 ( n1579 , n773 , n1355 );
    and g3188 ( n606 , n1349 , n3518 );
    or g3189 ( n1573 , n680 , n3449 );
    nor g3190 ( n1668 , n3420 , n137 );
    not g3191 ( n2072 , n2813 );
    nor g3192 ( n1909 , n1318 , n3243 );
    and g3193 ( n736 , n2327 , n2953 );
    or g3194 ( n1646 , n35 , n3252 );
    not g3195 ( n1025 , n1517 );
    and g3196 ( n2863 , n2583 , n2658 );
    or g3197 ( n2047 , n2473 , n761 );
    not g3198 ( n643 , n3474 );
    not g3199 ( n2413 , n2625 );
    nor g3200 ( n1795 , n2246 , n1449 );
    or g3201 ( n1041 , n2699 , n1188 );
    or g3202 ( n1288 , n1340 , n1077 );
    or g3203 ( n2700 , n170 , n3436 );
    nor g3204 ( n3263 , n3508 , n2238 );
    or g3205 ( n54 , n1353 , n1177 );
    or g3206 ( n1639 , n37 , n3737 );
    or g3207 ( n902 , n2893 , n3169 );
    and g3208 ( n2782 , n1730 , n3011 );
    and g3209 ( n848 , n1394 , n3727 );
    nor g3210 ( n335 , n165 , n3500 );
    or g3211 ( n3848 , n1330 , n2367 );
    and g3212 ( n593 , n2022 , n1352 );
    nor g3213 ( n2618 , n2378 , n1570 );
    and g3214 ( n3114 , n2852 , n3291 );
    and g3215 ( n3024 , n437 , n2875 );
    and g3216 ( n2388 , n3277 , n2811 );
    nor g3217 ( n360 , n2121 , n54 );
    or g3218 ( n340 , n2591 , n2575 );
    or g3219 ( n1083 , n2383 , n283 );
    nor g3220 ( n586 , n1145 , n3057 );
    and g3221 ( n3066 , n1846 , n2217 );
    or g3222 ( n559 , n1472 , n2743 );
    or g3223 ( n2573 , n712 , n571 );
    nor g3224 ( n182 , n802 , n3904 );
    nor g3225 ( n408 , n3350 , n1671 );
    not g3226 ( n2629 , n2906 );
    and g3227 ( n2575 , n840 , n1198 );
    and g3228 ( n3012 , n1612 , n3001 );
    nor g3229 ( n2841 , n2000 , n3892 );
    nor g3230 ( n1908 , n2 , n929 );
    and g3231 ( n584 , n2908 , n1636 );
    and g3232 ( n3104 , n3546 , n16 );
    not g3233 ( n2800 , n3593 );
    nor g3234 ( n3461 , n635 , n3419 );
    or g3235 ( n1473 , n1307 , n193 );
    or g3236 ( n2510 , n1926 , n3015 );
    or g3237 ( n2041 , n284 , n2607 );
    nor g3238 ( n2425 , n96 , n870 );
    nor g3239 ( n1425 , n692 , n1639 );
    and g3240 ( n1098 , n2472 , n3069 );
    or g3241 ( n345 , n886 , n3102 );
    nor g3242 ( n3549 , n1216 , n3803 );
    not g3243 ( n1665 , n304 );
    or g3244 ( n3106 , n3562 , n3145 );
    or g3245 ( n3567 , n528 , n807 );
    or g3246 ( n2327 , n1686 , n1213 );
    or g3247 ( n3075 , n3598 , n3910 );
    or g3248 ( n1797 , n3370 , n3692 );
    and g3249 ( n925 , n355 , n3712 );
    not g3250 ( n3700 , n3268 );
    or g3251 ( n2609 , n2184 , n1617 );
    not g3252 ( n312 , n2311 );
    or g3253 ( n3188 , n3773 , n2639 );
    not g3254 ( n454 , n1341 );
    or g3255 ( n3753 , n1151 , n3169 );
    and g3256 ( n2001 , n2258 , n470 );
    nor g3257 ( n1693 , n75 , n2607 );
    nor g3258 ( n3872 , n3255 , n1320 );
    and g3259 ( n795 , n570 , n1010 );
    or g3260 ( n1771 , n1964 , n2654 );
    nor g3261 ( n3085 , n2865 , n3635 );
    not g3262 ( n1495 , n31 );
    and g3263 ( n3459 , n2981 , n3023 );
    and g3264 ( n2046 , n3232 , n1049 );
    not g3265 ( n2109 , n3648 );
    nor g3266 ( n3676 , n1489 , n1121 );
    or g3267 ( n3270 , n2446 , n2798 );
    nor g3268 ( n1992 , n2470 , n592 );
    and g3269 ( n1524 , n2886 , n3743 );
    or g3270 ( n1054 , n803 , n571 );
    and g3271 ( n2997 , n394 , n1926 );
    not g3272 ( n2287 , n1309 );
    nor g3273 ( n940 , n2382 , n2914 );
    not g3274 ( n2929 , n44 );
    not g3275 ( n1462 , n3450 );
    nor g3276 ( n3776 , n357 , n2346 );
    or g3277 ( n2094 , n3405 , n2386 );
    or g3278 ( n3727 , n1583 , n571 );
    or g3279 ( n2604 , n408 , n1354 );
    and g3280 ( n1248 , n874 , n3679 );
    and g3281 ( n1618 , n488 , n1379 );
    and g3282 ( n306 , n3139 , n3476 );
    not g3283 ( n3741 , n2253 );
    not g3284 ( n2543 , n2477 );
    or g3285 ( n49 , n3670 , n1275 );
    and g3286 ( n17 , n2566 , n2428 );
    and g3287 ( n3054 , n2506 , n941 );
    or g3288 ( n3381 , n3402 , n3466 );
    nor g3289 ( n1081 , n2234 , n3865 );
    not g3290 ( n1452 , n10 );
    not g3291 ( n3366 , n3345 );
    not g3292 ( n637 , n747 );
    nor g3293 ( n633 , n2146 , n1633 );
    nor g3294 ( n2294 , n197 , n831 );
    and g3295 ( n402 , n2271 , n2478 );
    or g3296 ( n3433 , n3241 , n586 );
    nor g3297 ( n1142 , n3519 , n1000 );
    and g3298 ( n1435 , n917 , n2677 );
    not g3299 ( n3212 , n2625 );
    nor g3300 ( n515 , n2320 , n2081 );
    or g3301 ( n2584 , n2923 , n3005 );
    nor g3302 ( n2998 , n1651 , n3802 );
    and g3303 ( n2562 , n1893 , n1919 );
    not g3304 ( n363 , n3517 );
    not g3305 ( n735 , n1814 );
    nor g3306 ( n1436 , n2616 , n2601 );
    or g3307 ( n247 , n2705 , n2785 );
    and g3308 ( n758 , n2337 , n998 );
    nor g3309 ( n773 , n2491 , n831 );
    and g3310 ( n1255 , n2724 , n3813 );
    nor g3311 ( n2937 , n3473 , n3090 );
    and g3312 ( n1760 , n1893 , n1914 );
    nor g3313 ( n3821 , n272 , n1815 );
    or g3314 ( n3123 , n2865 , n1916 );
    and g3315 ( n329 , n2291 , n634 );
    and g3316 ( n1021 , n3773 , n3471 );
    or g3317 ( n12 , n2043 , n3169 );
    nor g3318 ( n2200 , n2710 , n298 );
    or g3319 ( n538 , n2415 , n2122 );
    or g3320 ( n2740 , n1549 , n761 );
    or g3321 ( n3818 , n221 , n143 );
    and g3322 ( n3531 , n2486 , n3380 );
    not g3323 ( n1334 , n3693 );
    and g3324 ( n470 , n3568 , n147 );
    and g3325 ( n528 , n3431 , n266 );
    nor g3326 ( n1946 , n723 , n3483 );
    and g3327 ( n3476 , n3720 , n3587 );
    not g3328 ( n2071 , n687 );
    and g3329 ( n1611 , n3789 , n301 );
    and g3330 ( n2982 , n1510 , n3016 );
    and g3331 ( n3732 , n2502 , n691 );
    not g3332 ( n3522 , n3066 );
    or g3333 ( n2050 , n3716 , n2147 );
    not g3334 ( n2506 , n3171 );
    and g3335 ( n2320 , n254 , n144 );
    and g3336 ( n2166 , n1511 , n2313 );
    not g3337 ( n2179 , n2664 );
    or g3338 ( n2182 , n2993 , n3003 );
    and g3339 ( n3681 , n3487 , n1518 );
    or g3340 ( n1031 , n3060 , n1916 );
    not g3341 ( n2486 , n2625 );
    not g3342 ( n1833 , n855 );
    and g3343 ( n3665 , n3369 , n1311 );
    or g3344 ( n1235 , n1817 , n2580 );
    nor g3345 ( n2895 , n3706 , n431 );
    and g3346 ( n1672 , n852 , n2536 );
    or g3347 ( n3125 , n805 , n509 );
    not g3348 ( n1664 , n3379 );
    or g3349 ( n3035 , n88 , n1593 );
    or g3350 ( n673 , n3119 , n761 );
    not g3351 ( n87 , n1897 );
    and g3352 ( n490 , n1249 , n2702 );
    or g3353 ( n1304 , n3553 , n1624 );
    or g3354 ( n1230 , n3574 , n3604 );
    or g3355 ( n999 , n1491 , n653 );
    not g3356 ( n1475 , n2628 );
    or g3357 ( n1036 , n974 , n761 );
    and g3358 ( n3861 , n1365 , n1663 );
    or g3359 ( n3469 , n1099 , n2420 );
    and g3360 ( n1905 , n1893 , n684 );
    and g3361 ( n1551 , n3804 , n3198 );
    and g3362 ( n2852 , n3309 , n2534 );
    and g3363 ( n2897 , n3019 , n1103 );
    and g3364 ( n362 , n1894 , n3755 );
    and g3365 ( n2743 , n1974 , n3190 );
    and g3366 ( n533 , n155 , n121 );
    nor g3367 ( n3122 , n3605 , n2171 );
    and g3368 ( n2219 , n3566 , n1358 );
    nor g3369 ( n887 , n252 , n3543 );
    nor g3370 ( n26 , n2497 , n1367 );
    and g3371 ( n2936 , n2585 , n1123 );
    or g3372 ( n332 , n227 , n3742 );
    or g3373 ( n483 , n3810 , n831 );
    nor g3374 ( n2014 , n3124 , n2607 );
    or g3375 ( n1487 , n2429 , n1294 );
    or g3376 ( n1726 , n1610 , n1453 );
    and g3377 ( n3674 , n333 , n1938 );
    not g3378 ( n412 , n2371 );
    and g3379 ( n3814 , n3490 , n629 );
    not g3380 ( n3438 , n652 );
    and g3381 ( n2220 , n2806 , n1061 );
    and g3382 ( n3410 , n3230 , n3236 );
    nor g3383 ( n1315 , n2564 , n1554 );
    and g3384 ( n3269 , n1495 , n3422 );
    or g3385 ( n3435 , n2867 , n3875 );
    not g3386 ( n2297 , n1214 );
    nor g3387 ( n1472 , n2182 , n3578 );
    or g3388 ( n1344 , n991 , n2607 );
    or g3389 ( n2139 , n3518 , n1349 );
    not g3390 ( n3266 , n733 );
    and g3391 ( n2837 , n2485 , n1708 );
    or g3392 ( n234 , n1666 , n1898 );
    and g3393 ( n2332 , n3589 , n154 );
    or g3394 ( n3150 , n515 , n3290 );
    and g3395 ( n2726 , n2652 , n1663 );
    or g3396 ( n300 , n3832 , n3671 );
    not g3397 ( n2844 , n1100 );
    not g3398 ( n1943 , n1827 );
    and g3399 ( n3513 , n186 , n1997 );
    and g3400 ( n694 , n1258 , n2163 );
    not g3401 ( n1224 , n1629 );
    and g3402 ( n530 , n3053 , n526 );
    or g3403 ( n1437 , n1286 , n1247 );
    and g3404 ( n3619 , n2625 , n497 );
    or g3405 ( n771 , n2945 , n908 );
    and g3406 ( n699 , n3556 , n2204 );
    and g3407 ( n599 , n3134 , n1769 );
    and g3408 ( n2012 , n3174 , n2440 );
    and g3409 ( n3353 , n3344 , n105 );
    or g3410 ( n2694 , n3002 , n3742 );
    and g3411 ( n3058 , n923 , n3909 );
    not g3412 ( n287 , n467 );
    nor g3413 ( n2511 , n526 , n1916 );
    not g3414 ( n713 , n3256 );
    or g3415 ( n2869 , n2207 , n3274 );
    and g3416 ( n2930 , n2151 , n329 );
    and g3417 ( n1651 , n3785 , n3873 );
    or g3418 ( n1161 , n3779 , n349 );
    nor g3419 ( n1592 , n1697 , n2426 );
    and g3420 ( n1512 , n3652 , n670 );
    nor g3421 ( n3293 , n919 , n3572 );
    and g3422 ( n1175 , n1785 , n2696 );
    or g3423 ( n1521 , n42 , n2996 );
    or g3424 ( n3307 , n997 , n780 );
    or g3425 ( n2550 , n2197 , n2750 );
    and g3426 ( n3029 , n2777 , n1944 );
    not g3427 ( n1119 , n1201 );
    or g3428 ( n3354 , n140 , n137 );
    not g3429 ( n3317 , n467 );
    and g3430 ( n929 , n1498 , n136 );
    not g3431 ( n2845 , n467 );
    nor g3432 ( n3378 , n713 , n3212 );
    or g3433 ( n3131 , n3378 , n452 );
    nor g3434 ( n3795 , n2287 , n3354 );
    or g3435 ( n3812 , n422 , n3738 );
    or g3436 ( n374 , n967 , n280 );
    and g3437 ( n1981 , n253 , n2173 );
    nor g3438 ( n348 , n3919 , n157 );
    not g3439 ( n872 , n1276 );
endmodule
