module top( n19 , n22 , n27 , n29 , n36 , n40 , n65 , n86 , n94 , 
n95 , n97 , n99 , n104 , n105 , n114 , n115 , n118 , n121 , n123 , 
n124 , n125 , n128 , n133 , n137 , n145 , n147 , n148 , n159 , n161 , 
n178 , n190 , n192 , n193 , n195 , n196 , n198 , n200 , n201 , n204 , 
n208 , n211 , n212 , n214 , n221 , n223 , n238 , n241 , n258 , n280 , 
n281 , n285 , n287 , n288 , n293 , n294 , n303 , n325 , n328 );
    input n22 , n27 , n36 , n65 , n94 , n99 , n104 , n105 , n114 , 
n115 , n118 , n123 , n125 , n128 , n145 , n147 , n190 , n196 , n200 , 
n201 , n208 , n211 , n221 , n223 , n238 , n258 , n281 , n287 , n288 , 
n294 , n303 , n325 , n328 ;
    output n19 , n29 , n40 , n86 , n95 , n97 , n121 , n124 , n133 , 
n137 , n148 , n159 , n161 , n178 , n192 , n193 , n195 , n198 , n204 , 
n212 , n214 , n241 , n280 , n285 , n293 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , 
n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , 
n20 , n21 , n23 , n24 , n25 , n26 , n28 , n30 , n31 , n32 , 
n33 , n34 , n35 , n37 , n38 , n39 , n41 , n42 , n43 , n44 , 
n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , 
n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , 
n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , 
n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , 
n87 , n88 , n89 , n90 , n91 , n92 , n93 , n96 , n98 , n100 , 
n101 , n102 , n103 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , 
n113 , n116 , n117 , n119 , n120 , n122 , n126 , n127 , n129 , n130 , 
n131 , n132 , n134 , n135 , n136 , n138 , n139 , n140 , n141 , n142 , 
n143 , n144 , n146 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , 
n156 , n157 , n158 , n160 , n162 , n163 , n164 , n165 , n166 , n167 , 
n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , 
n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , 
n189 , n191 , n194 , n197 , n199 , n202 , n203 , n205 , n206 , n207 , 
n209 , n210 , n213 , n215 , n216 , n217 , n218 , n219 , n220 , n222 , 
n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , 
n234 , n235 , n236 , n237 , n239 , n240 , n242 , n243 , n244 , n245 , 
n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , 
n256 , n257 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , 
n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , 
n277 , n278 , n279 , n282 , n283 , n284 , n286 , n289 , n290 , n291 , 
n292 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n304 , 
n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , 
n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , 
n326 , n327 , n329 , n330 , n331 , n332 , n333 , n334 ;
    or g0 ( n72 , n290 , n318 );
    nor g1 ( n76 , n294 , n49 );
    xnor g2 ( n285 , n278 , n328 );
    not g3 ( n129 , n200 );
    or g4 ( n171 , n224 , n23 );
    not g5 ( n17 , n324 );
    or g6 ( n53 , n219 , n211 );
    xnor g7 ( n97 , n227 , n99 );
    and g8 ( n249 , n295 , n4 );
    not g9 ( n320 , n199 );
    not g10 ( n120 , n257 );
    or g11 ( n78 , n72 , n237 );
    not g12 ( n314 , n174 );
    or g13 ( n10 , n28 , n249 );
    nor g14 ( n131 , n89 , n119 );
    xnor g15 ( n6 , n79 , n101 );
    xnor g16 ( n71 , n229 , n51 );
    or g17 ( n259 , n58 , n12 );
    xnor g18 ( n253 , n328 , n147 );
    xnor g19 ( n168 , n176 , n287 );
    nor g20 ( n59 , n205 , n170 );
    or g21 ( n286 , n177 , n170 );
    or g22 ( n77 , n252 , n9 );
    not g23 ( n33 , n22 );
    xnor g24 ( n236 , n221 , n94 );
    xnor g25 ( n256 , n84 , n46 );
    or g26 ( n226 , n47 , n186 );
    or g27 ( n9 , n102 , n186 );
    or g28 ( n315 , n205 , n284 );
    or g29 ( n12 , n183 , n275 );
    xnor g30 ( n84 , n232 , n166 );
    nor g31 ( n245 , n294 , n256 );
    or g32 ( n274 , n85 , n242 );
    or g33 ( n45 , n299 , n186 );
    or g34 ( n189 , n157 , n120 );
    xnor g35 ( n317 , n236 , n36 );
    and g36 ( n246 , n179 , n235 );
    xnor g37 ( n192 , n313 , n36 );
    nor g38 ( n88 , n205 , n231 );
    or g39 ( n284 , n42 , n320 );
    and g40 ( n183 , n325 , n210 );
    xnor g41 ( n46 , n196 , n94 );
    or g42 ( n133 , n117 , n112 );
    or g43 ( n186 , n72 , n12 );
    not g44 ( n74 , n34 );
    or g45 ( n34 , n87 , n93 );
    xnor g46 ( n275 , n279 , n65 );
    nor g47 ( n56 , n211 , n297 );
    nor g48 ( n220 , n144 , n78 );
    xnor g49 ( n291 , n265 , n55 );
    or g50 ( n103 , n251 , n108 );
    or g51 ( n144 , n298 , n168 );
    xnor g52 ( n160 , n291 , n53 );
    xnor g53 ( n193 , n139 , n94 );
    not g54 ( n224 , n208 );
    nor g55 ( n1 , n219 , n18 );
    nor g56 ( n148 , n43 , n262 );
    not g57 ( n80 , n321 );
    xnor g58 ( n241 , n301 , n196 );
    not g59 ( n82 , n128 );
    xnor g60 ( n178 , n164 , n288 );
    and g61 ( n92 , n156 , n23 );
    or g62 ( n11 , n231 , n237 );
    or g63 ( n112 , n109 , n307 );
    nor g64 ( n3 , n2 , n78 );
    and g65 ( n322 , n23 , n149 );
    not g66 ( n98 , n258 );
    xnor g67 ( n49 , n308 , n6 );
    or g68 ( n307 , n151 , n113 );
    nor g69 ( n167 , n205 , n299 );
    not g70 ( n306 , n309 );
    or g71 ( n248 , n177 , n126 );
    not g72 ( n244 , n201 );
    or g73 ( n0 , n102 , n186 );
    nor g74 ( n271 , n83 , n197 );
    or g75 ( n15 , n191 , n155 );
    xnor g76 ( n86 , n103 , n304 );
    xnor g77 ( n280 , n163 , n238 );
    xnor g78 ( n276 , n49 , n154 );
    or g79 ( n302 , n152 , n146 );
    xor g80 ( n332 , n30 , n223 );
    or g81 ( n106 , n257 , n169 );
    or g82 ( n209 , n286 , n58 );
    xor g83 ( n30 , n303 , n99 );
    not g84 ( n313 , n107 );
    nor g85 ( n235 , n2 , n259 );
    or g86 ( n62 , n57 , n282 );
    xnor g87 ( n304 , n140 , n106 );
    or g88 ( n252 , n127 , n170 );
    nor g89 ( n41 , n205 , n231 );
    or g90 ( n136 , n177 , n26 );
    and g91 ( n309 , n44 , n5 );
    or g92 ( n215 , n177 , n299 );
    nor g93 ( n247 , n2 , n186 );
    or g94 ( n87 , n127 , n284 );
    or g95 ( n135 , n174 , n255 );
    or g96 ( n47 , n298 , n194 );
    nor g97 ( n296 , n127 , n2 );
    xnor g98 ( n90 , n190 , n223 );
    or g99 ( n324 , n300 , n91 );
    xnor g100 ( n308 , n243 , n303 );
    or g101 ( n138 , n127 , n284 );
    nor g102 ( n95 , n43 , n260 );
    or g103 ( n67 , n23 , n189 );
    nor g104 ( n198 , n43 , n264 );
    xnor g105 ( n222 , n250 , n245 );
    not g106 ( n194 , n168 );
    xnor g107 ( n134 , n130 , n125 );
    nor g108 ( n57 , n184 , n153 );
    not g109 ( n96 , n105 );
    not g110 ( n110 , n246 );
    and g111 ( n43 , n211 , n82 );
    or g112 ( n210 , n244 , n294 );
    nor g113 ( n182 , n30 , n111 );
    and g114 ( n279 , n23 , n160 );
    xnor g115 ( n204 , n110 , n221 );
    nor g116 ( n214 , n43 , n276 );
    or g117 ( n217 , n311 , n306 );
    or g118 ( n184 , n299 , n231 );
    xnor g119 ( n185 , n333 , n330 );
    nor g120 ( n331 , n181 , n119 );
    and g121 ( n321 , n88 , n220 );
    nor g122 ( n66 , n170 , n186 );
    nor g123 ( n295 , n289 , n58 );
    or g124 ( n272 , n58 , n237 );
    or g125 ( n292 , n23 , n316 );
    and g126 ( n174 , n41 , n66 );
    xnor g127 ( n262 , n160 , n131 );
    and g128 ( n310 , n296 , n268 );
    xnor g129 ( n121 , n77 , n223 );
    xnor g130 ( n48 , n332 , n190 );
    and g131 ( n176 , n23 , n13 );
    xnor g132 ( n243 , n90 , n238 );
    or g133 ( n163 , n116 , n0 );
    or g134 ( n237 , n183 , n254 );
    or g135 ( n164 , n180 , n226 );
    nor g136 ( n4 , n284 , n237 );
    or g137 ( n68 , n98 , n123 );
    or g138 ( n267 , n62 , n20 );
    xnor g139 ( n38 , n70 , n175 );
    xor g140 ( n40 , n310 , n190 );
    nor g141 ( n140 , n211 , n309 );
    or g142 ( n270 , n75 , n269 );
    nor g143 ( n161 , n43 , n16 );
    nor g144 ( n165 , n205 , n47 );
    xnor g145 ( n264 , n149 , n239 );
    nor g146 ( n239 , n171 , n119 );
    xnor g147 ( n79 , n162 , n132 );
    xnor g148 ( n162 , n196 , n147 );
    xnor g149 ( n232 , n332 , n238 );
    xnor g150 ( n13 , n38 , n216 );
    or g151 ( n297 , n188 , n244 );
    nor g152 ( n5 , n135 , n150 );
    not g153 ( n156 , n123 );
    not g154 ( n172 , n287 );
    not g155 ( n188 , n325 );
    and g156 ( n81 , n211 , n18 );
    or g157 ( n316 , n250 , n119 );
    and g158 ( n107 , n230 , n31 );
    and g159 ( n157 , n201 , n123 );
    not g160 ( n24 , n210 );
    nor g161 ( n31 , n2 , n259 );
    or g162 ( n20 , n50 , n334 );
    not g163 ( n254 , n275 );
    and g164 ( n191 , n59 , n266 );
    or g165 ( n60 , n107 , n246 );
    xnor g166 ( n124 , n61 , n125 );
    or g167 ( n326 , n310 , n14 );
    xnor g168 ( n29 , n34 , n303 );
    or g169 ( n39 , n172 , n23 );
    or g170 ( n7 , n251 , n1 );
    nor g171 ( n151 , n233 , n272 );
    not g172 ( n119 , n217 );
    xnor g173 ( n54 , n288 , n190 );
    or g174 ( n261 , n23 , n327 );
    or g175 ( n83 , n215 , n58 );
    or g176 ( n319 , n81 , n182 );
    or g177 ( n58 , n290 , n141 );
    or g178 ( n206 , n231 , n237 );
    xnor g179 ( n298 , n218 , n22 );
    not g180 ( n228 , n92 );
    or g181 ( n173 , n299 , n231 );
    or g182 ( n139 , n158 , n323 );
    not g183 ( n213 , n115 );
    nor g184 ( n50 , n143 , n11 );
    not g185 ( n14 , n77 );
    or g186 ( n154 , n23 , n274 );
    nor g187 ( n212 , n43 , n122 );
    or g188 ( n2 , n222 , n199 );
    or g189 ( n301 , n315 , n45 );
    xnor g190 ( n70 , n145 , n147 );
    not g191 ( n203 , n311 );
    xnor g192 ( n333 , n253 , n225 );
    not g193 ( n278 , n155 );
    nor g194 ( n207 , n39 , n242 );
    xnor g195 ( n132 , n32 , n63 );
    or g196 ( n69 , n170 , n259 );
    not g197 ( n187 , n81 );
    or g198 ( n202 , n82 , n157 );
    xnor g199 ( n216 , n48 , n27 );
    or g200 ( n181 , n33 , n23 );
    xnor g201 ( n35 , n27 , n288 );
    or g202 ( n146 , n326 , n270 );
    or g203 ( n180 , n205 , n231 );
    nor g204 ( n266 , n2 , n78 );
    or g205 ( n311 , n60 , n302 );
    or g206 ( n91 , n102 , n78 );
    and g207 ( n257 , n211 , n21 );
    xnor g208 ( n277 , n238 , n221 );
    xnor g209 ( n16 , n13 , n207 );
    or g210 ( n158 , n127 , n299 );
    or g211 ( n289 , n177 , n299 );
    xnor g212 ( n234 , n111 , n63 );
    nor g213 ( n108 , n96 , n21 );
    nor g214 ( n229 , n211 , n203 );
    nor g215 ( n130 , n211 , n64 );
    or g216 ( n64 , n213 , n123 );
    xnor g217 ( n63 , n283 , n145 );
    and g218 ( n255 , n167 , n247 );
    and g219 ( n127 , n177 , n261 );
    or g220 ( n152 , n100 , n74 );
    or g221 ( n73 , n299 , n231 );
    and g222 ( n155 , n165 , n3 );
    and g223 ( n205 , n177 , n67 );
    xnor g224 ( n195 , n314 , n27 );
    or g225 ( n116 , n127 , n47 );
    not g226 ( n8 , n65 );
    nor g227 ( n109 , n73 , n136 );
    or g228 ( n300 , n205 , n299 );
    nor g229 ( n282 , n37 , n240 );
    nor g230 ( n142 , n211 , n68 );
    or g231 ( n197 , n2 , n237 );
    not g232 ( n21 , n281 );
    not g233 ( n23 , n294 );
    and g234 ( n263 , n30 , n111 );
    xnor g235 ( n137 , n329 , n145 );
    nor g236 ( n268 , n144 , n186 );
    xnor g237 ( n141 , n85 , n76 );
    or g238 ( n323 , n102 , n259 );
    not g239 ( n61 , n255 );
    xnor g240 ( n265 , n111 , n32 );
    xnor g241 ( n122 , n185 , n331 );
    not g242 ( n269 , n139 );
    not g243 ( n42 , n222 );
    or g244 ( n299 , n312 , n194 );
    or g245 ( n150 , n305 , n15 );
    or g246 ( n102 , n42 , n199 );
    not g247 ( n329 , n191 );
    or g248 ( n231 , n222 , n320 );
    or g249 ( n85 , n213 , n92 );
    or g250 ( n89 , n8 , n23 );
    or g251 ( n93 , n170 , n78 );
    not g252 ( n251 , n211 );
    xnor g253 ( n159 , n80 , n147 );
    or g254 ( n26 , n141 , n237 );
    or g255 ( n177 , n211 , n202 );
    and g256 ( n290 , n258 , n228 );
    or g257 ( n305 , n321 , n17 );
    or g258 ( n334 , n271 , n52 );
    nor g259 ( n52 , n209 , n206 );
    xnor g260 ( n175 , n142 , n36 );
    xnor g261 ( n166 , n56 , n104 );
    not g262 ( n242 , n217 );
    or g263 ( n117 , n10 , n267 );
    xnor g264 ( n260 , n256 , n292 );
    or g265 ( n273 , n177 , n47 );
    or g266 ( n233 , n299 , n231 );
    not g267 ( n318 , n141 );
    not g268 ( n219 , n114 );
    xnor g269 ( n32 , n35 , n125 );
    or g270 ( n101 , n96 , n211 );
    nor g271 ( n28 , n173 , n248 );
    not g272 ( n18 , n118 );
    not g273 ( n100 , n163 );
    or g274 ( n240 , n177 , n78 );
    or g275 ( n153 , n177 , n259 );
    or g276 ( n126 , n58 , n254 );
    not g277 ( n312 , n298 );
    or g278 ( n143 , n273 , n58 );
    xnor g279 ( n149 , n134 , n234 );
    xnor g280 ( n55 , n196 , n99 );
    and g281 ( n218 , n23 , n185 );
    or g282 ( n250 , n129 , n24 );
    not g283 ( n169 , n79 );
    xnor g284 ( n283 , n328 , n104 );
    or g285 ( n37 , n299 , n231 );
    nor g286 ( n179 , n127 , n47 );
    xnor g287 ( n293 , n7 , n71 );
    xnor g288 ( n330 , n54 , n277 );
    or g289 ( n170 , n312 , n168 );
    xnor g290 ( n111 , n243 , n317 );
    or g291 ( n51 , n263 , n319 );
    or g292 ( n227 , n138 , n69 );
    or g293 ( n25 , n129 , n244 );
    nor g294 ( n225 , n211 , n25 );
    nor g295 ( n230 , n127 , n170 );
    or g296 ( n113 , n211 , n217 );
    not g297 ( n75 , n227 );
    and g298 ( n44 , n164 , n301 );
    xnor g299 ( n199 , n322 , n208 );
    or g300 ( n327 , n157 , n187 );
    xnor g301 ( n19 , n324 , n104 );
endmodule
