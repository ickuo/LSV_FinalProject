// Benchmark "top" written by ABC on Sun Dec 21 18:08:54 2025

module top ( 
    n5, n13, n17, n20, n36, n37, n53, n75, n80, n86, n93, n105, n106, n111,
    n117, n139, n147, n157, n161, n182, n190, n198, n204, n208, n214, n217,
    n219, n224, n226, n229, n235, n244, n249, n281, n287, n289, n300, n303,
    n319, n346, n364, n365, n368, n384, n393, n403, n409, n410, n417, n439,
    n457, n465, n473, n477, n503, n506, n511, n518, n521, n532, n537, n587,
    n588, n593, n594, n595, n606, n642, n648, n656, n671, n680, n684, n690,
    n693, n699, n702, n706, n716, n741, n742, n743, n746, n777, n782, n788,
    n27, n62, n145, n175, n176, n225, n241, n256, n294, n345, n387, n389,
    n430, n442, n489, n491, n493, n515, n618, n630, n691, n703, n704, n753,
    n756, n765  );
  input  n5, n13, n17, n20, n36, n37, n53, n75, n80, n86, n93, n105,
    n106, n111, n117, n139, n147, n157, n161, n182, n190, n198, n204, n208,
    n214, n217, n219, n224, n226, n229, n235, n244, n249, n281, n287, n289,
    n300, n303, n319, n346, n364, n365, n368, n384, n393, n403, n409, n410,
    n417, n439, n457, n465, n473, n477, n503, n506, n511, n518, n521, n532,
    n537, n587, n588, n593, n594, n595, n606, n642, n648, n656, n671, n680,
    n684, n690, n693, n699, n702, n706, n716, n741, n742, n743, n746, n777,
    n782, n788;
  output n27, n62, n145, n175, n176, n225, n241, n256, n294, n345, n387, n389,
    n430, n442, n489, n491, n493, n515, n618, n630, n691, n703, n704, n753,
    n756, n765;
  wire new_n113, new_n114, new_n115, new_n116, new_n117_1, new_n118,
    new_n119, new_n120, new_n121, new_n122, new_n123, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139_1,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145_1, new_n146,
    new_n147_1, new_n148, new_n149, new_n150, new_n151, new_n152, new_n153,
    new_n154, new_n155, new_n156, new_n157_1, new_n158, new_n159, new_n160,
    new_n161_1, new_n162, new_n163, new_n164, new_n165, new_n166, new_n167,
    new_n168, new_n169, new_n170, new_n171, new_n172, new_n173, new_n174,
    new_n175_1, new_n176_1, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182_1, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190_1, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198_1, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204_1, new_n205, new_n206, new_n207,
    new_n208_1, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214_1, new_n215, new_n216, new_n217_1, new_n218, new_n219_1,
    new_n220, new_n221, new_n222, new_n223, new_n224_1, new_n225_1,
    new_n226_1, new_n227, new_n228, new_n229_1, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235_1, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241_1, new_n242, new_n243, new_n244_1,
    new_n245, new_n246, new_n247, new_n248, new_n249_1, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256_1, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281_1, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287_1, new_n288, new_n289_1, new_n290, new_n291, new_n292,
    new_n293, new_n294_1, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300_1, new_n301, new_n302, new_n303_1, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319_1,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345_1, new_n346_1,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n356, new_n357, new_n358, new_n359, new_n360,
    new_n361, new_n362, new_n363, new_n364_1, new_n365_1, new_n366,
    new_n367, new_n368_1, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384_1, new_n385, new_n386,
    new_n387_1, new_n388, new_n389_1, new_n390, new_n391, new_n392,
    new_n393_1, new_n394, new_n395, new_n396, new_n397, new_n398, new_n399,
    new_n400, new_n401, new_n402, new_n403_1, new_n404, new_n405, new_n406,
    new_n407, new_n408, new_n409_1, new_n410_1, new_n411, new_n412,
    new_n413, new_n414, new_n415, new_n416, new_n417_1, new_n418, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n430_1, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n439_1, new_n440,
    new_n441, new_n442_1, new_n443, new_n444, new_n445, new_n446, new_n447,
    new_n448, new_n449, new_n450, new_n451, new_n452, new_n453, new_n454,
    new_n455, new_n456, new_n457_1, new_n458, new_n459, new_n460, new_n461,
    new_n462, new_n463, new_n464, new_n465_1, new_n466, new_n467, new_n468,
    new_n469, new_n470, new_n471, new_n472, new_n473_1, new_n474, new_n475,
    new_n476, new_n477_1, new_n478, new_n479, new_n480, new_n481, new_n482,
    new_n483, new_n484, new_n485, new_n486, new_n487, new_n488, new_n489_1,
    new_n490, new_n491_1, new_n492, new_n493_1, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506_1, new_n507, new_n508, new_n509,
    new_n511_1, new_n512, new_n513, new_n514, new_n515_1, new_n516,
    new_n517, new_n518_1, new_n519, new_n521_1, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532_1,
    new_n533, new_n534, new_n535, new_n536, new_n537_1, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587_1, new_n588_1, new_n590, new_n591,
    new_n592, new_n593_1, new_n594_1, new_n595_1, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606_1,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618_1, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630_1, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642_1, new_n643, new_n645, new_n646,
    new_n648_1, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656_1, new_n657, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671_1,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684_1, new_n686, new_n687, new_n688,
    new_n689, new_n690_1, new_n692, new_n693_1, new_n694, new_n695,
    new_n697, new_n698, new_n699_1, new_n700;
  assign new_n113 = n217 & n690;
  assign new_n114 = n217 & n365;
  assign new_n115 = ~n690 & ~new_n114;
  assign new_n116 = ~new_n113 & ~new_n115;
  assign new_n117_1 = ~n503 & ~new_n116;
  assign new_n118 = n503 & new_n116;
  assign new_n119 = n217 & ~n365;
  assign new_n120 = n690 & ~new_n119;
  assign new_n121 = ~n690 & new_n119;
  assign new_n122 = ~new_n120 & ~new_n121;
  assign new_n123 = n503 & new_n122;
  assign new_n124 = ~n503 & ~new_n122;
  assign new_n125 = ~n217 & ~n365;
  assign new_n126 = ~new_n114 & ~new_n125;
  assign new_n127 = ~n680 & ~new_n126;
  assign new_n128 = n680 & new_n126;
  assign new_n129 = n5 & n365;
  assign new_n130 = ~new_n128 & ~new_n129;
  assign new_n131 = ~new_n127 & ~new_n130;
  assign new_n132 = ~new_n124 & ~new_n131;
  assign new_n133 = ~new_n123 & ~new_n132;
  assign new_n134 = ~new_n118 & ~new_n133;
  assign new_n135 = ~new_n117_1 & ~new_n134;
  assign new_n136 = new_n113 & new_n135;
  assign new_n137 = n393 & new_n136;
  assign new_n138 = ~n300 & ~n537;
  assign new_n139_1 = ~n403 & new_n138;
  assign new_n140 = ~n393 & new_n139_1;
  assign new_n141 = ~n106 & new_n140;
  assign new_n142 = n139 & new_n141;
  assign new_n143 = ~new_n137 & ~new_n142;
  assign new_n144 = ~n182 & ~n503;
  assign new_n145_1 = n182 & n503;
  assign new_n146 = ~n594 & ~n680;
  assign new_n147_1 = n594 & n680;
  assign new_n148 = n5 & n671;
  assign new_n149 = ~n5 & ~n671;
  assign new_n150 = n157 & n303;
  assign new_n151 = ~new_n149 & new_n150;
  assign new_n152 = ~new_n148 & ~new_n151;
  assign new_n153 = ~new_n147_1 & new_n152;
  assign new_n154 = ~new_n146 & ~new_n153;
  assign new_n155 = ~new_n145_1 & ~new_n154;
  assign new_n156 = ~new_n144 & ~new_n155;
  assign new_n157_1 = n777 & new_n156;
  assign new_n158 = n281 & new_n157_1;
  assign new_n159 = n699 & new_n158;
  assign new_n160 = ~n699 & ~new_n158;
  assign new_n161_1 = ~new_n159 & ~new_n160;
  assign new_n162 = n656 & ~new_n161_1;
  assign new_n163 = ~n518 & ~n656;
  assign new_n164 = ~new_n162 & ~new_n163;
  assign new_n165 = ~new_n143 & new_n164;
  assign new_n166 = new_n143 & ~new_n164;
  assign new_n167 = n319 & new_n141;
  assign new_n168 = ~new_n113 & ~new_n135;
  assign new_n169 = n393 & ~new_n136;
  assign new_n170 = ~new_n168 & new_n169;
  assign new_n171 = ~new_n167 & ~new_n170;
  assign new_n172 = ~n281 & ~new_n157_1;
  assign new_n173 = ~new_n158 & ~new_n172;
  assign new_n174 = n656 & ~new_n173;
  assign new_n175_1 = ~n219 & ~n656;
  assign new_n176_1 = ~new_n174 & ~new_n175_1;
  assign new_n177 = ~new_n171 & new_n176_1;
  assign new_n178 = new_n171 & ~new_n176_1;
  assign new_n179 = n5 & n157;
  assign new_n180 = n680 & new_n179;
  assign new_n181 = n503 & new_n180;
  assign new_n182_1 = n403 & new_n181;
  assign new_n183 = ~n106 & new_n139_1;
  assign new_n184 = n93 & new_n183;
  assign new_n185 = ~n393 & ~new_n184;
  assign new_n186 = ~new_n182_1 & new_n185;
  assign new_n187 = ~new_n117_1 & ~new_n118;
  assign new_n188 = new_n133 & ~new_n187;
  assign new_n189 = ~new_n133 & new_n187;
  assign new_n190_1 = n393 & ~new_n189;
  assign new_n191 = ~new_n188 & new_n190_1;
  assign new_n192 = ~new_n186 & ~new_n191;
  assign new_n193 = n346 & ~n656;
  assign new_n194 = ~n777 & ~new_n156;
  assign new_n195 = ~new_n157_1 & ~new_n194;
  assign new_n196 = n656 & new_n195;
  assign new_n197 = ~new_n193 & ~new_n196;
  assign new_n198_1 = new_n192 & ~new_n197;
  assign new_n199 = ~new_n192 & new_n197;
  assign new_n200 = n13 & n17;
  assign new_n201 = ~n13 & ~n17;
  assign new_n202 = ~n439 & ~n742;
  assign new_n203 = n439 & n742;
  assign new_n204_1 = n111 & n642;
  assign new_n205 = ~new_n203 & ~new_n204_1;
  assign new_n206 = ~new_n202 & ~new_n205;
  assign new_n207 = ~new_n201 & new_n206;
  assign new_n208_1 = n106 & ~new_n207;
  assign new_n209 = ~new_n200 & new_n208_1;
  assign new_n210 = ~n106 & ~n746;
  assign new_n211 = ~n300 & ~new_n210;
  assign new_n212 = ~new_n209 & new_n211;
  assign new_n213 = n17 & n782;
  assign new_n214_1 = ~n17 & ~n782;
  assign new_n215 = ~n117 & ~n439;
  assign new_n216 = n117 & n439;
  assign new_n217_1 = n606 & n642;
  assign new_n218 = ~new_n216 & ~new_n217_1;
  assign new_n219_1 = ~new_n215 & ~new_n218;
  assign new_n220 = ~new_n214_1 & new_n219_1;
  assign new_n221 = ~new_n213 & ~new_n220;
  assign new_n222 = n300 & ~new_n221;
  assign new_n223 = ~n537 & ~new_n222;
  assign new_n224_1 = ~new_n212 & new_n223;
  assign new_n225_1 = ~n17 & ~n693;
  assign new_n226_1 = ~n249 & ~n439;
  assign new_n227 = n249 & n439;
  assign new_n228 = n409 & n642;
  assign new_n229_1 = ~new_n227 & ~new_n228;
  assign new_n230 = ~new_n226_1 & ~new_n229_1;
  assign new_n231 = ~new_n225_1 & new_n230;
  assign new_n232 = n17 & n693;
  assign new_n233 = n537 & ~new_n232;
  assign new_n234 = ~new_n231 & new_n233;
  assign new_n235_1 = ~n403 & ~new_n234;
  assign new_n236 = ~new_n224_1 & new_n235_1;
  assign new_n237 = ~n503 & ~new_n180;
  assign new_n238 = n403 & ~new_n237;
  assign new_n239 = ~new_n181 & new_n238;
  assign new_n240 = ~n393 & ~new_n239;
  assign new_n241_1 = ~new_n236 & new_n240;
  assign new_n242 = ~new_n123 & ~new_n124;
  assign new_n243 = ~new_n131 & new_n242;
  assign new_n244_1 = new_n131 & ~new_n242;
  assign new_n245 = n393 & ~new_n244_1;
  assign new_n246 = ~new_n243 & new_n245;
  assign new_n247 = ~new_n241_1 & ~new_n246;
  assign new_n248 = ~n287 & ~n656;
  assign new_n249_1 = ~new_n144 & ~new_n145_1;
  assign new_n250 = new_n154 & ~new_n249_1;
  assign new_n251 = ~new_n154 & new_n249_1;
  assign new_n252 = ~new_n250 & ~new_n251;
  assign new_n253 = n656 & new_n252;
  assign new_n254 = ~new_n248 & ~new_n253;
  assign new_n255 = ~new_n247 & ~new_n254;
  assign new_n256_1 = ~new_n200 & ~new_n201;
  assign new_n257 = new_n206 & ~new_n256_1;
  assign new_n258 = ~new_n206 & new_n256_1;
  assign new_n259 = ~new_n257 & ~new_n258;
  assign new_n260 = n106 & ~new_n259;
  assign new_n261 = ~n106 & n473;
  assign new_n262 = ~n300 & ~new_n261;
  assign new_n263 = ~new_n260 & new_n262;
  assign new_n264 = ~new_n213 & ~new_n214_1;
  assign new_n265 = ~new_n219_1 & new_n264;
  assign new_n266 = new_n219_1 & ~new_n264;
  assign new_n267 = n300 & ~new_n266;
  assign new_n268 = ~new_n265 & new_n267;
  assign new_n269 = ~new_n263 & ~new_n268;
  assign new_n270 = ~n537 & ~new_n269;
  assign new_n271 = ~new_n225_1 & ~new_n232;
  assign new_n272 = ~new_n230 & new_n271;
  assign new_n273 = new_n230 & ~new_n271;
  assign new_n274 = n537 & ~new_n273;
  assign new_n275 = ~new_n272 & new_n274;
  assign new_n276 = ~n403 & ~new_n275;
  assign new_n277 = ~new_n270 & new_n276;
  assign new_n278 = ~n680 & ~new_n179;
  assign new_n279 = n403 & ~new_n278;
  assign new_n280 = ~new_n180 & new_n279;
  assign new_n281_1 = ~n393 & ~new_n280;
  assign new_n282 = ~new_n277 & new_n281_1;
  assign new_n283 = ~new_n127 & new_n130;
  assign new_n284 = ~new_n127 & ~new_n128;
  assign new_n285 = new_n129 & ~new_n284;
  assign new_n286 = n393 & ~new_n285;
  assign new_n287_1 = ~new_n283 & new_n286;
  assign new_n288 = ~new_n282 & ~new_n287_1;
  assign new_n289_1 = ~n656 & ~n706;
  assign new_n290 = ~new_n146 & ~new_n147_1;
  assign new_n291 = new_n152 & new_n290;
  assign new_n292 = ~new_n152 & ~new_n290;
  assign new_n293 = ~new_n291 & ~new_n292;
  assign new_n294_1 = n656 & new_n293;
  assign new_n295 = ~new_n289_1 & ~new_n294_1;
  assign new_n296 = ~new_n288 & ~new_n295;
  assign new_n297 = ~n5 & ~n365;
  assign new_n298 = ~new_n129 & ~new_n297;
  assign new_n299 = n393 & ~new_n298;
  assign new_n300_1 = ~n106 & ~n511;
  assign new_n301 = ~n300 & ~new_n300_1;
  assign new_n302 = ~new_n202 & ~new_n203;
  assign new_n303_1 = new_n204_1 & ~new_n302;
  assign new_n304 = ~new_n204_1 & new_n302;
  assign new_n305 = ~new_n303_1 & ~new_n304;
  assign new_n306 = n106 & new_n305;
  assign new_n307 = new_n301 & ~new_n306;
  assign new_n308 = ~new_n215 & ~new_n216;
  assign new_n309 = new_n217_1 & new_n308;
  assign new_n310 = ~new_n217_1 & ~new_n308;
  assign new_n311 = n300 & ~new_n310;
  assign new_n312 = ~new_n309 & new_n311;
  assign new_n313 = ~new_n307 & ~new_n312;
  assign new_n314 = ~n537 & ~new_n313;
  assign new_n315 = ~new_n226_1 & ~new_n227;
  assign new_n316 = ~new_n228 & ~new_n315;
  assign new_n317 = new_n228 & new_n315;
  assign new_n318 = ~new_n316 & ~new_n317;
  assign new_n319_1 = n537 & new_n318;
  assign new_n320 = ~new_n314 & ~new_n319_1;
  assign new_n321 = ~n403 & ~new_n320;
  assign new_n322 = ~n5 & ~n157;
  assign new_n323 = ~new_n179 & ~new_n322;
  assign new_n324 = n403 & new_n323;
  assign new_n325 = ~new_n321 & ~new_n324;
  assign new_n326 = ~n393 & new_n325;
  assign new_n327 = ~new_n299 & ~new_n326;
  assign new_n328 = ~n656 & n684;
  assign new_n329 = ~n157 & ~n303;
  assign new_n330 = n656 & ~new_n329;
  assign new_n331 = ~new_n150 & new_n330;
  assign new_n332 = ~new_n328 & ~new_n331;
  assign new_n333 = n157 & n393;
  assign new_n334 = ~n111 & ~n642;
  assign new_n335 = ~new_n204_1 & ~new_n334;
  assign new_n336 = n106 & ~new_n335;
  assign new_n337 = ~n106 & ~n289;
  assign new_n338 = ~n300 & ~new_n337;
  assign new_n339 = ~new_n336 & new_n338;
  assign new_n340 = ~n606 & ~n642;
  assign new_n341 = n300 & ~new_n217_1;
  assign new_n342 = ~new_n340 & new_n341;
  assign new_n343 = ~new_n339 & ~new_n342;
  assign new_n344 = ~n537 & ~new_n343;
  assign new_n345_1 = ~n409 & ~n642;
  assign new_n346_1 = n537 & ~new_n345_1;
  assign new_n347 = ~new_n228 & new_n346_1;
  assign new_n348 = ~n403 & ~new_n347;
  assign new_n349 = ~new_n344 & new_n348;
  assign new_n350 = n157 & n403;
  assign new_n351 = ~n393 & ~new_n350;
  assign new_n352 = ~new_n349 & new_n351;
  assign new_n353 = ~new_n333 & ~new_n352;
  assign new_n354 = ~new_n332 & ~new_n353;
  assign new_n355 = ~n593 & ~n656;
  assign new_n356 = ~new_n148 & ~new_n149;
  assign new_n357 = new_n150 & new_n356;
  assign new_n358 = ~new_n150 & ~new_n356;
  assign new_n359 = ~new_n357 & ~new_n358;
  assign new_n360 = n656 & ~new_n359;
  assign new_n361 = ~new_n355 & ~new_n360;
  assign new_n362 = new_n354 & new_n361;
  assign new_n363 = ~new_n327 & ~new_n362;
  assign new_n364_1 = ~new_n354 & ~new_n361;
  assign new_n365_1 = ~new_n363 & ~new_n364_1;
  assign new_n366 = new_n288 & new_n295;
  assign new_n367 = ~new_n365_1 & ~new_n366;
  assign new_n368_1 = ~new_n296 & ~new_n367;
  assign new_n369 = new_n247 & new_n254;
  assign new_n370 = ~new_n368_1 & ~new_n369;
  assign new_n371 = ~new_n255 & ~new_n370;
  assign new_n372 = ~new_n199 & new_n371;
  assign new_n373 = ~new_n198_1 & ~new_n372;
  assign new_n374 = ~new_n178 & ~new_n373;
  assign new_n375 = ~new_n177 & ~new_n374;
  assign new_n376 = ~new_n166 & ~new_n375;
  assign new_n377 = ~new_n165 & ~new_n376;
  assign new_n378 = n384 & new_n159;
  assign new_n379 = n457 & new_n378;
  assign new_n380 = n648 & new_n379;
  assign new_n381 = ~n648 & ~new_n379;
  assign new_n382 = ~new_n380 & ~new_n381;
  assign new_n383 = n656 & ~new_n382;
  assign new_n384_1 = ~n588 & ~n656;
  assign new_n385 = ~new_n383 & ~new_n384_1;
  assign new_n386 = ~n656 & n743;
  assign new_n387_1 = ~n384 & ~new_n159;
  assign new_n388 = ~new_n378 & ~new_n387_1;
  assign new_n389_1 = n656 & new_n388;
  assign new_n390 = ~new_n386 & ~new_n389_1;
  assign new_n391 = ~n457 & ~new_n378;
  assign new_n392 = ~new_n379 & ~new_n391;
  assign new_n393_1 = n656 & ~new_n392;
  assign new_n394 = ~n368 & ~n656;
  assign new_n395 = ~new_n393_1 & ~new_n394;
  assign new_n396 = ~new_n390 & new_n395;
  assign new_n397 = new_n385 & new_n396;
  assign new_n398 = n204 & new_n380;
  assign new_n399 = n417 & new_n398;
  assign new_n400 = ~n417 & ~new_n398;
  assign new_n401 = ~new_n399 & ~new_n400;
  assign new_n402 = n656 & ~new_n401;
  assign new_n403_1 = ~n465 & ~n656;
  assign new_n404 = ~new_n402 & ~new_n403_1;
  assign new_n405 = new_n397 & new_n404;
  assign new_n406 = n244 & ~n656;
  assign new_n407 = ~n204 & ~new_n380;
  assign new_n408 = ~new_n398 & ~new_n407;
  assign new_n409_1 = n656 & new_n408;
  assign new_n410_1 = ~new_n406 & ~new_n409_1;
  assign new_n411 = new_n405 & ~new_n410_1;
  assign new_n412 = ~new_n377 & new_n411;
  assign new_n413 = n587 & ~n656;
  assign new_n414 = n20 & new_n399;
  assign new_n415 = ~n20 & ~new_n399;
  assign new_n416 = n656 & ~new_n415;
  assign new_n417_1 = ~new_n414 & new_n416;
  assign new_n418 = ~new_n413 & ~new_n417_1;
  assign new_n419 = new_n412 & ~new_n418;
  assign new_n420 = n595 & ~n656;
  assign new_n421 = n36 & new_n414;
  assign new_n422 = ~n36 & ~new_n414;
  assign new_n423 = n656 & ~new_n422;
  assign new_n424 = ~new_n421 & new_n423;
  assign new_n425 = ~new_n420 & ~new_n424;
  assign new_n426 = new_n419 & ~new_n425;
  assign new_n427 = n788 & new_n421;
  assign new_n428 = ~n788 & ~new_n421;
  assign new_n429 = ~new_n427 & ~new_n428;
  assign new_n430_1 = n656 & ~new_n429;
  assign new_n431 = ~n364 & ~n656;
  assign new_n432 = ~new_n430_1 & ~new_n431;
  assign new_n433 = new_n426 & new_n432;
  assign new_n434 = n741 & new_n427;
  assign new_n435 = ~n741 & ~new_n427;
  assign new_n436 = ~new_n434 & ~new_n435;
  assign new_n437 = n656 & ~new_n436;
  assign new_n438 = ~n235 & ~n656;
  assign new_n439_1 = ~new_n437 & ~new_n438;
  assign new_n440 = new_n433 & new_n439_1;
  assign new_n441 = n161 & ~n656;
  assign new_n442_1 = n716 & new_n434;
  assign new_n443 = ~n716 & ~new_n434;
  assign new_n444 = n656 & ~new_n443;
  assign new_n445 = ~new_n442_1 & new_n444;
  assign new_n446 = ~new_n441 & ~new_n445;
  assign new_n447 = new_n440 & ~new_n446;
  assign new_n448 = n190 & new_n442_1;
  assign new_n449 = ~n190 & ~new_n442_1;
  assign new_n450 = n656 & ~new_n449;
  assign new_n451 = ~new_n448 & new_n450;
  assign new_n452 = n532 & ~n656;
  assign new_n453 = ~new_n451 & ~new_n452;
  assign new_n454 = new_n447 & ~new_n453;
  assign new_n455 = ~n656 & ~new_n454;
  assign new_n456 = new_n143 & new_n164;
  assign new_n457_1 = ~new_n143 & ~new_n164;
  assign new_n458 = new_n171 & new_n176_1;
  assign new_n459 = ~new_n171 & ~new_n176_1;
  assign new_n460 = ~new_n192 & ~new_n197;
  assign new_n461 = new_n192 & new_n197;
  assign new_n462 = ~new_n247 & new_n254;
  assign new_n463 = new_n247 & ~new_n254;
  assign new_n464 = ~new_n288 & new_n295;
  assign new_n465_1 = new_n288 & ~new_n295;
  assign new_n466 = ~new_n327 & new_n361;
  assign new_n467 = new_n327 & ~new_n361;
  assign new_n468 = ~new_n331 & ~new_n353;
  assign new_n469 = ~new_n328 & new_n468;
  assign new_n470 = ~new_n467 & ~new_n469;
  assign new_n471 = ~new_n466 & ~new_n470;
  assign new_n472 = ~new_n465_1 & ~new_n471;
  assign new_n473_1 = ~new_n464 & ~new_n472;
  assign new_n474 = ~new_n463 & ~new_n473_1;
  assign new_n475 = ~new_n462 & ~new_n474;
  assign new_n476 = ~new_n461 & ~new_n475;
  assign new_n477_1 = ~new_n460 & ~new_n476;
  assign new_n478 = ~new_n459 & ~new_n477_1;
  assign new_n479 = ~new_n458 & ~new_n478;
  assign new_n480 = ~new_n457_1 & ~new_n479;
  assign new_n481 = ~new_n456 & ~new_n480;
  assign new_n482 = ~new_n385 & ~new_n395;
  assign new_n483 = new_n410_1 & new_n482;
  assign new_n484 = new_n390 & new_n483;
  assign new_n485 = new_n481 & new_n484;
  assign new_n486 = ~new_n404 & new_n485;
  assign new_n487 = new_n418 & new_n425;
  assign new_n488 = ~new_n432 & new_n487;
  assign new_n489_1 = new_n486 & new_n488;
  assign new_n490 = ~new_n439_1 & new_n489_1;
  assign new_n491_1 = n656 & ~new_n490;
  assign new_n492 = ~new_n445 & ~new_n491_1;
  assign new_n493_1 = ~new_n451 & new_n492;
  assign new_n494 = ~new_n455 & new_n493_1;
  assign new_n495 = ~n147 & ~new_n448;
  assign new_n496 = n147 & new_n448;
  assign new_n497 = ~new_n495 & ~new_n496;
  assign new_n498 = n656 & ~new_n497;
  assign new_n499 = ~n229 & ~n656;
  assign new_n500 = ~new_n498 & ~new_n499;
  assign new_n501 = new_n494 & new_n500;
  assign new_n502 = ~new_n494 & ~new_n500;
  assign n27 = ~new_n501 & ~new_n502;
  assign new_n504 = ~n656 & new_n368_1;
  assign new_n505 = n656 & new_n473_1;
  assign new_n506_1 = ~new_n504 & ~new_n505;
  assign new_n507 = ~new_n462 & ~new_n463;
  assign new_n508 = new_n506_1 & new_n507;
  assign new_n509 = ~new_n506_1 & ~new_n507;
  assign n62 = ~new_n508 & ~new_n509;
  assign new_n511_1 = ~n656 & ~new_n377;
  assign new_n512 = new_n397 & new_n511_1;
  assign new_n513 = n656 & new_n481;
  assign new_n514 = ~new_n388 & new_n513;
  assign new_n515_1 = ~new_n395 & new_n514;
  assign new_n516 = ~new_n385 & new_n515_1;
  assign new_n517 = ~new_n512 & ~new_n516;
  assign new_n518_1 = ~new_n410_1 & ~new_n517;
  assign new_n519 = new_n410_1 & new_n517;
  assign n145 = ~new_n518_1 & ~new_n519;
  assign new_n521_1 = new_n332 & new_n353;
  assign n175 = ~new_n354 & ~new_n521_1;
  assign new_n523 = ~new_n198_1 & ~new_n199;
  assign new_n524 = ~n656 & new_n371;
  assign new_n525 = n656 & new_n475;
  assign new_n526 = ~new_n524 & ~new_n525;
  assign new_n527 = ~new_n523 & new_n526;
  assign new_n528 = new_n523 & ~new_n526;
  assign n176 = ~new_n527 & ~new_n528;
  assign new_n530 = new_n454 & new_n500;
  assign new_n531 = ~n656 & n702;
  assign new_n532_1 = n521 & new_n496;
  assign new_n533 = ~n521 & ~new_n496;
  assign new_n534 = n656 & ~new_n533;
  assign new_n535 = ~new_n532_1 & new_n534;
  assign new_n536 = ~new_n531 & ~new_n535;
  assign new_n537_1 = new_n530 & ~new_n536;
  assign new_n538 = ~n656 & ~new_n537_1;
  assign new_n539 = ~n80 & ~n656;
  assign new_n540 = new_n453 & ~new_n500;
  assign new_n541 = new_n446 & new_n540;
  assign new_n542 = new_n490 & new_n541;
  assign new_n543 = n506 & new_n532_1;
  assign new_n544 = ~n506 & ~new_n532_1;
  assign new_n545 = ~new_n543 & ~new_n544;
  assign new_n546 = n656 & ~new_n545;
  assign new_n547 = ~new_n539 & ~new_n546;
  assign new_n548 = new_n536 & ~new_n547;
  assign new_n549 = new_n542 & new_n548;
  assign new_n550 = n656 & ~new_n549;
  assign new_n551 = ~new_n539 & ~new_n550;
  assign new_n552 = ~new_n538 & new_n551;
  assign new_n553 = n86 & new_n543;
  assign new_n554 = ~n86 & ~new_n543;
  assign new_n555 = n656 & ~new_n554;
  assign new_n556 = ~new_n553 & new_n555;
  assign new_n557 = n224 & ~n656;
  assign new_n558 = ~new_n556 & ~new_n557;
  assign new_n559 = ~n656 & new_n558;
  assign new_n560 = ~new_n556 & ~new_n559;
  assign new_n561 = new_n552 & new_n560;
  assign new_n562 = n208 & new_n553;
  assign new_n563 = ~n208 & ~new_n553;
  assign new_n564 = n656 & ~new_n563;
  assign new_n565 = ~new_n562 & new_n564;
  assign new_n566 = n75 & ~n656;
  assign new_n567 = ~new_n565 & ~new_n566;
  assign new_n568 = new_n561 & new_n567;
  assign new_n569 = ~new_n561 & ~new_n567;
  assign n225 = new_n568 | new_n569;
  assign new_n571 = ~new_n485 & ~new_n512;
  assign new_n572 = ~n244 & ~n656;
  assign new_n573 = ~new_n571 & ~new_n572;
  assign new_n574 = new_n404 & new_n573;
  assign new_n575 = ~new_n404 & ~new_n573;
  assign n241 = ~new_n574 & ~new_n575;
  assign new_n577 = ~n656 & ~new_n447;
  assign new_n578 = new_n492 & ~new_n577;
  assign new_n579 = ~new_n453 & new_n578;
  assign new_n580 = new_n453 & ~new_n578;
  assign n256 = ~new_n579 & ~new_n580;
  assign new_n582 = n656 & ~new_n486;
  assign new_n583 = ~new_n417_1 & ~new_n582;
  assign new_n584 = ~n656 & ~new_n426;
  assign new_n585 = ~new_n424 & ~new_n584;
  assign new_n586 = new_n583 & new_n585;
  assign new_n587_1 = new_n432 & new_n586;
  assign new_n588_1 = ~new_n432 & ~new_n586;
  assign n294 = ~new_n587_1 & ~new_n588_1;
  assign new_n590 = ~n656 & ~new_n375;
  assign new_n591 = n656 & new_n479;
  assign new_n592 = ~new_n590 & ~new_n591;
  assign new_n593_1 = ~new_n165 & ~new_n166;
  assign new_n594_1 = new_n592 & ~new_n593_1;
  assign new_n595_1 = ~new_n592 & new_n593_1;
  assign n345 = ~new_n594_1 & ~new_n595_1;
  assign new_n597 = n656 & ~new_n489_1;
  assign new_n598 = ~new_n431 & ~new_n597;
  assign new_n599 = ~new_n584 & new_n598;
  assign new_n600 = new_n439_1 & new_n599;
  assign new_n601 = ~new_n439_1 & ~new_n599;
  assign n387 = ~new_n600 & ~new_n601;
  assign new_n603 = n743 & new_n511_1;
  assign new_n604 = ~new_n514 & ~new_n603;
  assign new_n605 = ~new_n395 & new_n604;
  assign new_n606_1 = new_n395 & ~new_n604;
  assign n389 = ~new_n605 & ~new_n606_1;
  assign new_n608 = n656 & ~new_n471;
  assign new_n609 = ~n656 & ~new_n365_1;
  assign new_n610 = ~new_n608 & ~new_n609;
  assign new_n611 = ~new_n464 & ~new_n465_1;
  assign new_n612 = new_n610 & ~new_n611;
  assign new_n613 = ~new_n610 & new_n611;
  assign n430 = ~new_n612 & ~new_n613;
  assign new_n615 = ~n214 & ~new_n562;
  assign new_n616 = n214 & new_n562;
  assign new_n617 = n656 & ~new_n616;
  assign new_n618_1 = ~new_n615 & new_n617;
  assign new_n619 = ~n656 & new_n567;
  assign new_n620 = new_n561 & ~new_n619;
  assign new_n621 = ~new_n565 & new_n620;
  assign new_n622 = ~n105 & ~n656;
  assign new_n623 = new_n621 & ~new_n622;
  assign new_n624 = ~new_n618_1 & new_n623;
  assign new_n625 = n53 & new_n616;
  assign new_n626 = ~n53 & ~new_n616;
  assign new_n627 = n656 & ~new_n626;
  assign new_n628 = ~new_n625 & new_n627;
  assign new_n629 = n410 & ~n656;
  assign new_n630_1 = ~new_n628 & ~new_n629;
  assign new_n631 = ~new_n624 & new_n630_1;
  assign new_n632 = new_n624 & ~new_n630_1;
  assign n442 = ~new_n631 & ~new_n632;
  assign new_n634 = n656 & ~new_n542;
  assign new_n635 = ~new_n535 & ~new_n634;
  assign new_n636 = ~new_n538 & new_n635;
  assign new_n637 = new_n547 & ~new_n636;
  assign new_n638 = ~new_n547 & new_n636;
  assign n489 = new_n637 | new_n638;
  assign new_n640 = new_n395 & new_n603;
  assign new_n641 = ~new_n515_1 & ~new_n640;
  assign new_n642_1 = new_n385 & ~new_n641;
  assign new_n643 = ~new_n385 & new_n641;
  assign n491 = ~new_n642_1 & ~new_n643;
  assign new_n645 = new_n552 & ~new_n558;
  assign new_n646 = ~new_n552 & new_n558;
  assign n493 = ~new_n645 & ~new_n646;
  assign new_n648_1 = ~new_n511_1 & ~new_n513;
  assign new_n649 = ~new_n390 & new_n648_1;
  assign new_n650 = new_n390 & ~new_n648_1;
  assign n515 = new_n649 | new_n650;
  assign new_n652 = ~new_n458 & ~new_n459;
  assign new_n653 = ~n656 & ~new_n373;
  assign new_n654 = n656 & new_n477_1;
  assign new_n655 = ~new_n653 & ~new_n654;
  assign new_n656_1 = ~new_n652 & new_n655;
  assign new_n657 = new_n652 & ~new_n655;
  assign n618 = new_n656_1 | new_n657;
  assign new_n659 = ~n656 & ~new_n419;
  assign new_n660 = new_n583 & ~new_n659;
  assign new_n661 = ~new_n425 & new_n660;
  assign new_n662 = new_n425 & ~new_n660;
  assign n630 = ~new_n661 & ~new_n662;
  assign new_n664 = ~n410 & ~n656;
  assign new_n665 = ~new_n628 & ~new_n664;
  assign new_n666 = new_n624 & new_n665;
  assign new_n667 = n37 & ~new_n625;
  assign new_n668 = ~n37 & new_n625;
  assign new_n669 = ~new_n667 & ~new_n668;
  assign new_n670 = n656 & ~new_n669;
  assign new_n671_1 = n226 & ~n656;
  assign new_n672 = ~new_n670 & ~new_n671_1;
  assign new_n673 = ~new_n666 & ~new_n672;
  assign new_n674 = new_n666 & new_n672;
  assign n691 = new_n673 | new_n674;
  assign new_n676 = ~n656 & ~new_n412;
  assign new_n677 = ~new_n582 & ~new_n676;
  assign new_n678 = ~new_n418 & new_n677;
  assign new_n679 = new_n418 & ~new_n677;
  assign n703 = ~new_n678 & ~new_n679;
  assign new_n681 = n105 & ~n656;
  assign new_n682 = ~new_n618_1 & ~new_n681;
  assign new_n683 = new_n621 & new_n682;
  assign new_n684_1 = ~new_n621 & ~new_n682;
  assign n704 = new_n683 | new_n684_1;
  assign new_n686 = ~new_n466 & ~new_n467;
  assign new_n687 = ~n656 & ~n684;
  assign new_n688 = new_n468 & ~new_n687;
  assign new_n689 = new_n686 & new_n688;
  assign new_n690_1 = ~new_n686 & ~new_n688;
  assign n753 = new_n689 | new_n690_1;
  assign new_n692 = ~n656 & ~new_n440;
  assign new_n693_1 = ~new_n491_1 & ~new_n692;
  assign new_n694 = ~new_n446 & new_n693_1;
  assign new_n695 = new_n446 & ~new_n693_1;
  assign n756 = ~new_n694 & ~new_n695;
  assign new_n697 = ~new_n499 & ~new_n634;
  assign new_n698 = ~new_n455 & new_n697;
  assign new_n699_1 = ~new_n536 & new_n698;
  assign new_n700 = new_n536 & ~new_n698;
  assign n765 = ~new_n699_1 & ~new_n700;
endmodule


