module top( n1 , n8 , n9 , n21 , n24 , n32 , n54 , n61 , n64 , 
n67 , n69 , n76 , n83 , n84 , n96 , n97 , n107 , n110 , n117 , 
n120 , n128 , n135 , n137 , n142 , n145 , n147 , n150 , n154 , n167 , 
n170 , n172 , n182 , n184 , n190 , n198 , n204 , n209 , n210 , n220 , 
n222 , n230 , n231 , n232 , n233 , n240 , n253 , n265 , n268 , n269 , 
n283 , n289 , n290 , n291 , n292 , n293 , n296 , n313 , n324 , n325 , 
n330 , n336 , n342 , n347 , n350 , n356 , n362 , n363 , n364 , n365 , 
n368 , n373 , n383 , n386 , n388 , n403 , n415 , n418 , n421 , n427 , 
n432 , n434 , n468 , n476 , n478 , n480 , n481 , n489 , n490 , n506 , 
n507 , n514 , n524 , n526 , n532 , n543 , n565 , n574 , n576 , n579 , 
n588 , n596 , n598 , n605 , n608 , n614 , n615 , n618 , n623 , n629 , 
n633 , n635 , n640 , n646 , n654 , n656 , n663 , n664 , n675 , n676 , 
n677 , n678 , n691 , n693 , n704 , n710 , n716 , n717 , n722 , n726 , 
n727 , n737 , n740 , n750 , n751 , n765 , n769 , n785 , n786 , n790 , 
n793 , n794 , n797 , n800 , n814 , n818 , n821 , n824 , n829 , n835 , 
n836 , n837 , n840 , n842 , n845 , n848 , n851 , n857 , n859 , n869 , 
n877 , n887 , n894 , n901 , n909 , n923 , n928 , n933 , n934 , n938 , 
n950 , n956 , n964 , n973 , n974 , n989 , n990 , n1013 , n1014 , n1019 , 
n1021 , n1023 , n1025 , n1026 , n1030 , n1032 , n1036 , n1039 , n1042 , n1043 , 
n1049 , n1052 , n1058 , n1065 , n1070 , n1091 , n1093 , n1098 , n1099 , n1108 , 
n1117 , n1121 , n1122 , n1131 , n1134 , n1138 , n1143 , n1146 , n1150 , n1151 , 
n1157 , n1160 , n1161 , n1162 , n1165 , n1170 , n1177 , n1184 , n1187 , n1189 , 
n1192 , n1194 , n1198 , n1223 , n1239 , n1240 , n1243 , n1251 , n1253 , n1255 , 
n1275 , n1276 , n1280 , n1303 , n1310 , n1311 , n1314 , n1331 , n1335 , n1339 , 
n1361 , n1366 , n1373 , n1375 , n1378 , n1389 , n1392 , n1396 , n1398 , n1407 , 
n1409 , n1411 , n1412 , n1413 , n1418 , n1422 , n1425 , n1438 , n1442 , n1454 , 
n1474 , n1475 , n1478 , n1479 , n1485 , n1508 , n1511 , n1512 , n1515 , n1518 , 
n1530 , n1531 , n1542 , n1545 , n1547 , n1549 , n1551 , n1552 , n1555 , n1556 , 
n1562 , n1574 , n1575 , n1580 , n1581 , n1589 , n1594 , n1596 , n1601 , n1604 , 
n1606 , n1620 , n1628 , n1629 , n1630 , n1631 , n1645 , n1648 , n1655 , n1665 , 
n1671 , n1676 );
    input n1 , n9 , n67 , n69 , n84 , n96 , n107 , n120 , n128 , 
n135 , n137 , n145 , n147 , n182 , n184 , n198 , n209 , n220 , n222 , 
n230 , n233 , n268 , n283 , n289 , n290 , n293 , n296 , n325 , n330 , 
n342 , n356 , n362 , n365 , n373 , n386 , n403 , n415 , n418 , n421 , 
n432 , n468 , n478 , n481 , n490 , n507 , n514 , n526 , n532 , n574 , 
n576 , n579 , n588 , n596 , n605 , n615 , n629 , n635 , n646 , n654 , 
n664 , n677 , n704 , n710 , n716 , n726 , n727 , n737 , n750 , n751 , 
n765 , n769 , n793 , n794 , n797 , n818 , n824 , n829 , n835 , n837 , 
n842 , n848 , n851 , n857 , n859 , n869 , n877 , n901 , n909 , n923 , 
n933 , n934 , n938 , n950 , n956 , n973 , n974 , n989 , n990 , n1013 , 
n1014 , n1025 , n1030 , n1042 , n1049 , n1052 , n1058 , n1065 , n1070 , n1091 , 
n1093 , n1098 , n1099 , n1108 , n1121 , n1131 , n1134 , n1143 , n1146 , n1150 , 
n1161 , n1162 , n1165 , n1170 , n1184 , n1187 , n1189 , n1223 , n1240 , n1243 , 
n1251 , n1253 , n1255 , n1276 , n1280 , n1303 , n1310 , n1311 , n1331 , n1335 , 
n1339 , n1361 , n1366 , n1373 , n1378 , n1389 , n1396 , n1398 , n1407 , n1409 , 
n1412 , n1413 , n1418 , n1422 , n1425 , n1438 , n1475 , n1479 , n1485 , n1508 , 
n1511 , n1515 , n1518 , n1530 , n1545 , n1549 , n1551 , n1555 , n1562 , n1575 , 
n1580 , n1581 , n1596 , n1606 , n1620 , n1630 , n1648 , n1655 , n1676 ;
    output n8 , n21 , n24 , n32 , n54 , n61 , n64 , n76 , n83 , 
n97 , n110 , n117 , n142 , n150 , n154 , n167 , n170 , n172 , n190 , 
n204 , n210 , n231 , n232 , n240 , n253 , n265 , n269 , n291 , n292 , 
n313 , n324 , n336 , n347 , n350 , n363 , n364 , n368 , n383 , n388 , 
n427 , n434 , n476 , n480 , n489 , n506 , n524 , n543 , n565 , n598 , 
n608 , n614 , n618 , n623 , n633 , n640 , n656 , n663 , n675 , n676 , 
n678 , n691 , n693 , n717 , n722 , n740 , n785 , n786 , n790 , n800 , 
n814 , n821 , n836 , n840 , n845 , n887 , n894 , n928 , n964 , n1019 , 
n1021 , n1023 , n1026 , n1032 , n1036 , n1039 , n1043 , n1117 , n1122 , n1138 , 
n1151 , n1157 , n1160 , n1177 , n1192 , n1194 , n1198 , n1239 , n1275 , n1314 , 
n1375 , n1392 , n1411 , n1442 , n1454 , n1474 , n1478 , n1512 , n1531 , n1542 , 
n1547 , n1552 , n1556 , n1574 , n1589 , n1594 , n1601 , n1604 , n1628 , n1629 , 
n1631 , n1645 , n1665 , n1671 ;
    wire n0 , n2 , n3 , n4 , n5 , n6 , n7 , n10 , n11 , 
n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n22 , 
n23 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n33 , n34 , 
n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , 
n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n55 , 
n56 , n57 , n58 , n59 , n60 , n62 , n63 , n65 , n66 , n68 , 
n70 , n71 , n72 , n73 , n74 , n75 , n77 , n78 , n79 , n80 , 
n81 , n82 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , 
n93 , n94 , n95 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , 
n105 , n106 , n108 , n109 , n111 , n112 , n113 , n114 , n115 , n116 , 
n118 , n119 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n129 , 
n130 , n131 , n132 , n133 , n134 , n136 , n138 , n139 , n140 , n141 , 
n143 , n144 , n146 , n148 , n149 , n151 , n152 , n153 , n155 , n156 , 
n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
n168 , n169 , n171 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
n180 , n181 , n183 , n185 , n186 , n187 , n188 , n189 , n191 , n192 , 
n193 , n194 , n195 , n196 , n197 , n199 , n200 , n201 , n202 , n203 , 
n205 , n206 , n207 , n208 , n211 , n212 , n213 , n214 , n215 , n216 , 
n217 , n218 , n219 , n221 , n223 , n224 , n225 , n226 , n227 , n228 , 
n229 , n234 , n235 , n236 , n237 , n238 , n239 , n241 , n242 , n243 , 
n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n254 , 
n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , 
n266 , n267 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , 
n278 , n279 , n280 , n281 , n282 , n284 , n285 , n286 , n287 , n288 , 
n294 , n295 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , 
n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n314 , n315 , 
n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n326 , n327 , 
n328 , n329 , n331 , n332 , n333 , n334 , n335 , n337 , n338 , n339 , 
n340 , n341 , n343 , n344 , n345 , n346 , n348 , n349 , n351 , n352 , 
n353 , n354 , n355 , n357 , n358 , n359 , n360 , n361 , n366 , n367 , 
n369 , n370 , n371 , n372 , n374 , n375 , n376 , n377 , n378 , n379 , 
n380 , n381 , n382 , n384 , n385 , n387 , n389 , n390 , n391 , n392 , 
n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , 
n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , 
n414 , n416 , n417 , n419 , n420 , n422 , n423 , n424 , n425 , n426 , 
n428 , n429 , n430 , n431 , n433 , n435 , n436 , n437 , n438 , n439 , 
n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n469 , n470 , 
n471 , n472 , n473 , n474 , n475 , n477 , n479 , n482 , n483 , n484 , 
n485 , n486 , n487 , n488 , n491 , n492 , n493 , n494 , n495 , n496 , 
n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n508 , 
n509 , n510 , n511 , n512 , n513 , n515 , n516 , n517 , n518 , n519 , 
n520 , n521 , n522 , n523 , n525 , n527 , n528 , n529 , n530 , n531 , 
n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , 
n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , 
n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , 
n564 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n575 , 
n577 , n578 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , 
n589 , n590 , n591 , n592 , n593 , n594 , n595 , n597 , n599 , n600 , 
n601 , n602 , n603 , n604 , n606 , n607 , n609 , n610 , n611 , n612 , 
n613 , n616 , n617 , n619 , n620 , n621 , n622 , n624 , n625 , n626 , 
n627 , n628 , n630 , n631 , n632 , n634 , n636 , n637 , n638 , n639 , 
n641 , n642 , n643 , n644 , n645 , n647 , n648 , n649 , n650 , n651 , 
n652 , n653 , n655 , n657 , n658 , n659 , n660 , n661 , n662 , n665 , 
n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n679 , 
n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
n690 , n692 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , 
n702 , n703 , n705 , n706 , n707 , n708 , n709 , n711 , n712 , n713 , 
n714 , n715 , n718 , n719 , n720 , n721 , n723 , n724 , n725 , n728 , 
n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n738 , n739 , 
n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n752 , 
n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , 
n763 , n764 , n766 , n767 , n768 , n770 , n771 , n772 , n773 , n774 , 
n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , 
n787 , n788 , n789 , n791 , n792 , n795 , n796 , n798 , n799 , n801 , 
n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , 
n812 , n813 , n815 , n816 , n817 , n819 , n820 , n822 , n823 , n825 , 
n826 , n827 , n828 , n830 , n831 , n832 , n833 , n834 , n838 , n839 , 
n841 , n843 , n844 , n846 , n847 , n849 , n850 , n852 , n853 , n854 , 
n855 , n856 , n858 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , 
n867 , n868 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n878 , 
n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n888 , n889 , 
n890 , n891 , n892 , n893 , n895 , n896 , n897 , n898 , n899 , n900 , 
n902 , n903 , n904 , n905 , n906 , n907 , n908 , n910 , n911 , n912 , 
n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , 
n924 , n925 , n926 , n927 , n929 , n930 , n931 , n932 , n935 , n936 , 
n937 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , 
n948 , n949 , n951 , n952 , n953 , n954 , n955 , n957 , n958 , n959 , 
n960 , n961 , n962 , n963 , n965 , n966 , n967 , n968 , n969 , n970 , 
n971 , n972 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , 
n983 , n984 , n985 , n986 , n987 , n988 , n991 , n992 , n993 , n994 , 
n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , 
n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1015 , n1016 , 
n1017 , n1018 , n1020 , n1022 , n1024 , n1027 , n1028 , n1029 , n1031 , n1033 , 
n1034 , n1035 , n1037 , n1038 , n1040 , n1041 , n1044 , n1045 , n1046 , n1047 , 
n1048 , n1050 , n1051 , n1053 , n1054 , n1055 , n1056 , n1057 , n1059 , n1060 , 
n1061 , n1062 , n1063 , n1064 , n1066 , n1067 , n1068 , n1069 , n1071 , n1072 , 
n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , 
n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1092 , n1094 , 
n1095 , n1096 , n1097 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , 
n1107 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1118 , 
n1119 , n1120 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , 
n1132 , n1133 , n1135 , n1136 , n1137 , n1139 , n1140 , n1141 , n1142 , n1144 , 
n1145 , n1147 , n1148 , n1149 , n1152 , n1153 , n1154 , n1155 , n1156 , n1158 , 
n1159 , n1163 , n1164 , n1166 , n1167 , n1168 , n1169 , n1171 , n1172 , n1173 , 
n1174 , n1175 , n1176 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1185 , 
n1186 , n1188 , n1190 , n1191 , n1193 , n1195 , n1196 , n1197 , n1199 , n1200 , 
n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , 
n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , 
n1221 , n1222 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , 
n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1241 , n1242 , n1244 , 
n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1252 , n1254 , n1256 , n1257 , 
n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , 
n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1277 , n1278 , n1279 , 
n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , 
n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , 
n1301 , n1302 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1312 , n1313 , 
n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , 
n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1332 , n1333 , n1334 , n1336 , 
n1337 , n1338 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , 
n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , 
n1358 , n1359 , n1360 , n1362 , n1363 , n1364 , n1365 , n1367 , n1368 , n1369 , 
n1370 , n1371 , n1372 , n1374 , n1376 , n1377 , n1379 , n1380 , n1381 , n1382 , 
n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1390 , n1391 , n1393 , n1394 , 
n1395 , n1397 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , 
n1408 , n1410 , n1414 , n1415 , n1416 , n1417 , n1419 , n1420 , n1421 , n1423 , 
n1424 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , 
n1435 , n1436 , n1437 , n1439 , n1440 , n1441 , n1443 , n1444 , n1445 , n1446 , 
n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1455 , n1456 , n1457 , 
n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , 
n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1476 , n1477 , n1480 , n1481 , 
n1482 , n1483 , n1484 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , 
n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , 
n1503 , n1504 , n1505 , n1506 , n1507 , n1509 , n1510 , n1513 , n1514 , n1516 , 
n1517 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , 
n1528 , n1529 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
n1540 , n1541 , n1543 , n1544 , n1546 , n1548 , n1550 , n1553 , n1554 , n1557 , 
n1558 , n1559 , n1560 , n1561 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , 
n1569 , n1570 , n1571 , n1572 , n1573 , n1576 , n1577 , n1578 , n1579 , n1582 , 
n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1590 , n1591 , n1592 , n1593 , 
n1595 , n1597 , n1598 , n1599 , n1600 , n1602 , n1603 , n1605 , n1607 , n1608 , 
n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , 
n1619 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1632 , n1633 , 
n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , 
n1644 , n1646 , n1647 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1656 , 
n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1666 , n1667 , 
n1668 , n1669 , n1670 , n1672 , n1673 , n1674 , n1675 , n1677 ;
    nor g0 ( n806 , n1255 , n1030 );
    nor g1 ( n1163 , n1422 , n148 );
    nor g2 ( n1015 , n1041 , n967 );
    not g3 ( n1516 , n47 );
    or g4 ( n394 , n413 , n513 );
    nor g5 ( n1359 , n198 , n1053 );
    nor g6 ( n360 , n1255 , n1251 );
    not g7 ( n1472 , n1408 );
    not g8 ( n936 , n51 );
    xnor g9 ( n1635 , n915 , n1554 );
    xnor g10 ( n1447 , n1127 , n742 );
    nor g11 ( n402 , n1255 , n209 );
    or g12 ( n1043 , n1629 , n1529 );
    nor g13 ( n1294 , n605 , n734 );
    xor g14 ( n1282 , n1295 , n71 );
    or g15 ( n191 , n641 , n539 );
    and g16 ( n1033 , n1348 , n1535 );
    and g17 ( n667 , n1491 , n632 );
    not g18 ( n518 , n1365 );
    or g19 ( n1007 , n713 , n519 );
    or g20 ( n890 , n1517 , n1139 );
    or g21 ( n1491 , n275 , n277 );
    and g22 ( n71 , n975 , n570 );
    nor g23 ( n28 , n272 , n1283 );
    or g24 ( n1085 , n944 , n774 );
    or g25 ( n524 , n1629 , n1089 );
    not g26 ( n60 , n218 );
    not g27 ( n434 , n1587 );
    or g28 ( n151 , n917 , n783 );
    nor g29 ( n822 , n1133 , n931 );
    xor g30 ( n1496 , n1242 , n1265 );
    and g31 ( n1010 , n954 , n938 );
    or g32 ( n610 , n1530 , n245 );
    not g33 ( n1229 , n729 );
    or g34 ( n720 , n940 , n841 );
    not g35 ( n1384 , n847 );
    nor g36 ( n1320 , n1311 , n1030 );
    not g37 ( n1190 , n770 );
    not g38 ( n1324 , n825 );
    or g39 ( n79 , n1495 , n1446 );
    or g40 ( n598 , n425 , n177 );
    xnor g41 ( n1619 , n116 , n1669 );
    or g42 ( n506 , n1629 , n323 );
    not g43 ( n504 , n1624 );
    and g44 ( n981 , n1143 , n325 );
    nor g45 ( n542 , n402 , n1027 );
    nor g46 ( n1272 , n1274 , n1518 );
    or g47 ( n1609 , n243 , n28 );
    xnor g48 ( n949 , n453 , n500 );
    nor g49 ( n985 , n300 , n1211 );
    or g50 ( n47 , n550 , n320 );
    or g51 ( n287 , n559 , n492 );
    nor g52 ( n206 , n289 , n62 );
    xnor g53 ( n163 , n1554 , n1599 );
    nor g54 ( n1344 , n10 , n1478 );
    nor g55 ( n862 , n403 , n789 );
    and g56 ( n1428 , n224 , n514 );
    not g57 ( n1269 , n397 );
    or g58 ( n427 , n449 , n168 );
    nor g59 ( n1593 , n960 , n654 );
    not g60 ( n66 , n1290 );
    and g61 ( n57 , n707 , n877 );
    not g62 ( n1199 , n1356 );
    nor g63 ( n1178 , n622 , n677 );
    not g64 ( n140 , n1378 );
    xnor g65 ( n339 , n1481 , n662 );
    not g66 ( n558 , n532 );
    not g67 ( n400 , n902 );
    nor g68 ( n32 , n1629 , n1323 );
    not g69 ( n1181 , n646 );
    and g70 ( n1368 , n1338 , n1354 );
    nor g71 ( n87 , n848 , n525 );
    not g72 ( n174 , n1435 );
    xnor g73 ( n260 , n763 , n1058 );
    or g74 ( n725 , n922 , n1420 );
    xnor g75 ( n550 , n1390 , n147 );
    nor g76 ( n728 , n615 , n1199 );
    not g77 ( n2 , n1108 );
    not g78 ( n761 , n1147 );
    and g79 ( n83 , n224 , n415 );
    not g80 ( n649 , n1384 );
    and g81 ( n1100 , n737 , n1243 );
    nor g82 ( n927 , n483 , n239 );
    not g83 ( n962 , n1235 );
    or g84 ( n1219 , n584 , n81 );
    nor g85 ( n45 , n135 , n385 );
    nor g86 ( n286 , n464 , n248 );
    xnor g87 ( n746 , n121 , n600 );
    and g88 ( n540 , n929 , n1339 );
    or g89 ( n41 , n102 , n404 );
    or g90 ( n185 , n242 , n371 );
    nor g91 ( n471 , n1676 , n1195 );
    nor g92 ( n1454 , n1099 , n1499 );
    not g93 ( n227 , n1193 );
    and g94 ( n106 , n969 , n403 );
    or g95 ( n808 , n1180 , n1528 );
    and g96 ( n1647 , n1268 , n726 );
    nor g97 ( n895 , n950 , n644 );
    or g98 ( n543 , n1629 , n890 );
    nor g99 ( n1626 , n238 , n1143 );
    not g100 ( n72 , n956 );
    or g101 ( n534 , n658 , n849 );
    and g102 ( n370 , n1302 , n1379 );
    not g103 ( n754 , n196 );
    or g104 ( n1275 , n165 , n326 );
    and g105 ( n23 , n1465 , n751 );
    and g106 ( n343 , n1011 , n181 );
    nor g107 ( n1371 , n527 , n962 );
    nor g108 ( n644 , n1504 , n1248 );
    not g109 ( n1211 , n1457 );
    not g110 ( n1244 , n220 );
    nor g111 ( n1246 , n6 , n1272 );
    nor g112 ( n1258 , n120 , n930 );
    or g113 ( n854 , n331 , n104 );
    not g114 ( n517 , n121 );
    nor g115 ( n1179 , n42 , n1283 );
    or g116 ( n1417 , n839 , n1371 );
    nor g117 ( n1322 , n848 , n424 );
    nor g118 ( n1060 , n960 , n859 );
    or g119 ( n1604 , n1629 , n444 );
    or g120 ( n811 , n319 , n1543 );
    not g121 ( n1547 , n842 );
    not g122 ( n964 , n1520 );
    not g123 ( n1477 , n902 );
    and g124 ( n25 , n647 , n1 );
    nor g125 ( n169 , n256 , n1645 );
    or g126 ( n954 , n1320 , n1330 );
    xnor g127 ( n1191 , n1524 , n1435 );
    not g128 ( n1153 , n877 );
    not g129 ( n187 , n297 );
    and g130 ( n695 , n401 , n1108 );
    or g131 ( n7 , n228 , n714 );
    not g132 ( n1419 , n1038 );
    not g133 ( n463 , n573 );
    or g134 ( n1476 , n1654 , n736 );
    nor g135 ( n1316 , n960 , n646 );
    xnor g136 ( n1617 , n112 , n125 );
    not g137 ( n398 , n372 );
    nor g138 ( n1250 , n561 , n752 );
    or g139 ( n815 , n442 , n7 );
    xnor g140 ( n961 , n454 , n594 );
    and g141 ( n1576 , n800 , n507 );
    and g142 ( n682 , n628 , n184 );
    not g143 ( n670 , n1336 );
    nor g144 ( n913 , n1255 , n1518 );
    or g145 ( n1046 , n540 , n1203 );
    nor g146 ( n529 , n1606 , n1181 );
    or g147 ( n1375 , n1629 , n1657 );
    and g148 ( n1416 , n1234 , n93 );
    and g149 ( n589 , n564 , n1378 );
    not g150 ( n270 , n514 );
    or g151 ( n1531 , n8 , n741 );
    or g152 ( n1657 , n82 , n1079 );
    not g153 ( n438 , n550 );
    or g154 ( n254 , n4 , n44 );
    not g155 ( n801 , n863 );
    xnor g156 ( n1140 , n419 , n1634 );
    and g157 ( n531 , n135 , n325 );
    or g158 ( n495 , n1046 , n787 );
    or g159 ( n1095 , n943 , n724 );
    or g160 ( n1570 , n1215 , n864 );
    xor g161 ( n688 , n1304 , n1564 );
    nor g162 ( n333 , n198 , n72 );
    not g163 ( n1307 , n393 );
    nor g164 ( n1443 , n1014 , n166 );
    not g165 ( n1631 , n523 );
    or g166 ( n1210 , n295 , n1185 );
    and g167 ( n839 , n1524 , n1479 );
    and g168 ( n747 , n1013 , n1606 );
    or g169 ( n836 , n984 , n1559 );
    nor g170 ( n789 , n772 , n1376 );
    or g171 ( n473 , n1334 , n169 );
    not g172 ( n1493 , n184 );
    nor g173 ( n907 , n694 , n590 );
    and g174 ( n880 , n1364 , n765 );
    or g175 ( n1437 , n68 , n1659 );
    and g176 ( n123 , n1140 , n632 );
    nor g177 ( n810 , n289 , n819 );
    nor g178 ( n73 , n1410 , n1404 );
    nor g179 ( n1301 , n198 , n1105 );
    not g180 ( n618 , n797 );
    not g181 ( n75 , n932 );
    or g182 ( n849 , n728 , n465 );
    nor g183 ( n19 , n706 , n1593 );
    not g184 ( n0 , n997 );
    or g185 ( n1397 , n433 , n1399 );
    nor g186 ( n1565 , n1367 , n261 );
    or g187 ( n1343 , n1335 , n162 );
    nor g188 ( n1497 , n1042 , n183 );
    nor g189 ( n1018 , n735 , n1039 );
    xnor g190 ( n1076 , n870 , n1496 );
    nor g191 ( n607 , n1398 , n1560 );
    nor g192 ( n805 , n256 , n621 );
    not g193 ( n1129 , n573 );
    or g194 ( n844 , n118 , n698 );
    nor g195 ( n872 , n468 , n670 );
    not g196 ( n130 , n1360 );
    or g197 ( n24 , n1629 , n639 );
    or g198 ( n952 , n1124 , n200 );
    nor g199 ( n65 , n342 , n757 );
    and g200 ( n1583 , n1243 , n1253 );
    nor g201 ( n733 , n1 , n1632 );
    or g202 ( n1050 , n856 , n100 );
    not g203 ( n1499 , n1412 );
    nor g204 ( n208 , n198 , n1526 );
    and g205 ( n1651 , n1596 , n1606 );
    nor g206 ( n1468 , n221 , n1302 );
    not g207 ( n416 , n280 );
    or g208 ( n1214 , n874 , n1449 );
    not g209 ( n1012 , n517 );
    xnor g210 ( n500 , n620 , n241 );
    or g211 ( n1313 , n1221 , n1625 );
    xnor g212 ( n1109 , n1335 , n629 );
    xnor g213 ( n1613 , n859 , n677 );
    nor g214 ( n1394 , n283 , n792 );
    not g215 ( n675 , n196 );
    nor g216 ( n515 , n1243 , n72 );
    or g217 ( n194 , n103 , n322 );
    not g218 ( n781 , n1587 );
    nor g219 ( n965 , n933 , n1156 );
    not g220 ( n112 , n975 );
    not g221 ( n1578 , n1405 );
    or g222 ( n1502 , n1140 , n318 );
    nor g223 ( n1567 , n615 , n1022 );
    nor g224 ( n1224 , n818 , n544 );
    xnor g225 ( n1257 , n268 , n209 );
    and g226 ( n972 , n746 , n632 );
    and g227 ( n219 , n616 , n765 );
    or g228 ( n297 , n747 , n886 );
    xor g229 ( n216 , n940 , n1329 );
    and g230 ( n1450 , n69 , n1243 );
    and g231 ( n327 , n156 , n145 );
    nor g232 ( n81 , n1227 , n291 );
    or g233 ( n387 , n1346 , n208 );
    nor g234 ( n1273 , n1511 , n959 );
    buf g235 ( n717 , n1134 );
    and g236 ( n1217 , n579 , n1243 );
    and g237 ( n617 , n956 , n325 );
    not g238 ( n1288 , n625 );
    nor g239 ( n226 , n236 , n1251 );
    xnor g240 ( n930 , n1308 , n835 );
    or g241 ( n1079 , n1238 , n5 );
    not g242 ( n1402 , n652 );
    not g243 ( n55 , n1251 );
    not g244 ( n1039 , n1440 );
    or g245 ( n846 , n1094 , n983 );
    xnor g246 ( n911 , n361 , n1165 );
    xnor g247 ( n121 , n1430 , n1389 );
    not g248 ( n1636 , n931 );
    or g249 ( n1466 , n267 , n1400 );
    nor g250 ( n1188 , n198 , n884 );
    and g251 ( n1020 , n407 , n632 );
    or g252 ( n1594 , n484 , n475 );
    xnor g253 ( n1632 , n1463 , n1434 );
    nor g254 ( n1287 , n198 , n935 );
    not g255 ( n94 , n115 );
    xor g256 ( n1107 , n1319 , n1264 );
    nor g257 ( n1399 , n735 , n964 );
    and g258 ( n1653 , n490 , n325 );
    nor g259 ( n876 , n843 , n1177 );
    and g260 ( n1369 , n1413 , n989 );
    xnor g261 ( n454 , n1572 , n1591 );
    not g262 ( n887 , n1247 );
    buf g263 ( n1629 , n1090 );
    xnor g264 ( n1434 , n372 , n613 );
    xnor g265 ( n116 , n161 , n625 );
    or g266 ( n401 , n1600 , n947 );
    not g267 ( n304 , n982 );
    not g268 ( n1204 , n306 );
    nor g269 ( n464 , n1255 , n135 );
    nor g270 ( n111 , n1398 , n665 );
    nor g271 ( n888 , n1425 , n999 );
    or g272 ( n1130 , n1481 , n1292 );
    or g273 ( n683 , n140 , n1416 );
    or g274 ( n1154 , n38 , n867 );
    xnor g275 ( n1483 , n1635 , n1298 );
    and g276 ( n597 , n149 , n796 );
    and g277 ( n50 , n416 , n570 );
    or g278 ( n199 , n759 , n1359 );
    nor g279 ( n1505 , n882 , n1256 );
    or g280 ( n1510 , n1293 , n548 );
    nor g281 ( n281 , n367 , n52 );
    or g282 ( n165 , n1000 , n307 );
    not g283 ( n1427 , n507 );
    nor g284 ( n1633 , n1091 , n665 );
    or g285 ( n894 , n1629 , n472 );
    and g286 ( n714 , n1067 , n1520 );
    nor g287 ( n1112 , n897 , n971 );
    and g288 ( n1644 , n1143 , n230 );
    and g289 ( n1220 , n351 , n869 );
    xnor g290 ( n443 , n738 , n1002 );
    not g291 ( n734 , n908 );
    not g292 ( n259 , n1615 );
    nor g293 ( n486 , n1667 , n686 );
    not g294 ( n1247 , n392 );
    buf g295 ( n232 , n480 );
    nor g296 ( n702 , n1606 , n800 );
    xnor g297 ( n419 , n625 , n403 );
    not g298 ( n1062 , n1432 );
    nor g299 ( n580 , n355 , n556 );
    and g300 ( n623 , n455 , n521 );
    not g301 ( n320 , n493 );
    or g302 ( n736 , n1007 , n1437 );
    and g303 ( n1135 , n997 , n1121 );
    and g304 ( n314 , n356 , n1243 );
    or g305 ( n467 , n1471 , n537 );
    and g306 ( n1618 , n481 , n1606 );
    nor g307 ( n447 , n451 , n316 );
    not g308 ( n1159 , n731 );
    and g309 ( n1507 , n1492 , n147 );
    nor g310 ( n703 , n882 , n394 );
    and g311 ( n445 , n176 , n950 );
    not g312 ( n1465 , n218 );
    not g313 ( n512 , n1409 );
    and g314 ( n560 , n1331 , n1243 );
    nor g315 ( n309 , n342 , n649 );
    and g316 ( n730 , n1470 , n1232 );
    nor g317 ( n175 , n304 , n863 );
    or g318 ( n698 , n681 , n131 );
    nor g319 ( n906 , n1311 , n135 );
    not g320 ( n1105 , n135 );
    or g321 ( n347 , n1629 , n1313 );
    xnor g322 ( n282 , n643 , n1047 );
    nor g323 ( n631 , n1108 , n1077 );
    nor g324 ( n759 , n1311 , n646 );
    not g325 ( n545 , n1166 );
    nor g326 ( n986 , n272 , n210 );
    and g327 ( n834 , n416 , n94 );
    nor g328 ( n1061 , n1184 , n1650 );
    and g329 ( n85 , n1152 , n490 );
    or g330 ( n203 , n23 , n430 );
    or g331 ( n181 , n1357 , n70 );
    not g332 ( n1333 , n57 );
    not g333 ( n1557 , n621 );
    not g334 ( n1432 , n1173 );
    xnor g335 ( n788 , n1047 , n1128 );
    or g336 ( n1540 , n1186 , n705 );
    and g337 ( n493 , n274 , n777 );
    or g338 ( n313 , n1629 , n1461 );
    buf g339 ( n786 , n478 );
    or g340 ( n1340 , n171 , n764 );
    or g341 ( n1083 , n349 , n1344 );
    or g342 ( n484 , n1607 , n900 );
    not g343 ( n861 , n1342 );
    and g344 ( n4 , n373 , n1243 );
    not g345 ( n385 , n365 );
    not g346 ( n902 , n138 );
    not g347 ( n882 , n1290 );
    xnor g348 ( n1084 , n1035 , n1619 );
    or g349 ( n99 , n1264 , n657 );
    or g350 ( n828 , n1289 , n978 );
    and g351 ( n275 , n968 , n1421 );
    nor g352 ( n1292 , n1242 , n600 );
    or g353 ( n168 , n1055 , n805 );
    or g354 ( n104 , n186 , n437 );
    and g355 ( n22 , n1382 , n1165 );
    or g356 ( n231 , n284 , n650 );
    or g357 ( n721 , n1226 , n1502 );
    or g358 ( n1654 , n749 , n538 );
    nor g359 ( n1215 , n1378 , n1527 );
    or g360 ( n966 , n271 , n216 );
    nor g361 ( n582 , n577 , n643 );
    not g362 ( n125 , n459 );
    nor g363 ( n511 , n1311 , n1518 );
    nor g364 ( n946 , n1146 , n130 );
    xnor g365 ( n141 , n1627 , n376 );
    not g366 ( n825 , n1137 );
    or g367 ( n117 , n811 , n1284 );
    or g368 ( n150 , n1629 , n1154 );
    and g369 ( n706 , n654 , n325 );
    not g370 ( n884 , n209 );
    or g371 ( n1577 , n375 , n795 );
    nor g372 ( n638 , n1605 , n824 );
    not g373 ( n43 , n283 );
    nor g374 ( n1185 , n1058 , n385 );
    not g375 ( n753 , n419 );
    xnor g376 ( n431 , n264 , n922 );
    xnor g377 ( n587 , n1637 , n1045 );
    or g378 ( n93 , n1181 , n700 );
    not g379 ( n34 , n1436 );
    and g380 ( n1193 , n488 , n1551 );
    nor g381 ( n382 , n1621 , n860 );
    not g382 ( n1022 , n1336 );
    or g383 ( n35 , n578 , n571 );
    not g384 ( n183 , n701 );
    or g385 ( n684 , n965 , n143 );
    not g386 ( n1342 , n66 );
    nor g387 ( n29 , n1064 , n124 );
    not g388 ( n1148 , n1170 );
    and g389 ( n1088 , n1545 , n230 );
    or g390 ( n1519 , n1658 , n1590 );
    or g391 ( n444 , n651 , n976 );
    and g392 ( n1525 , n107 , n1243 );
    nor g393 ( n396 , n1361 , n1480 );
    nor g394 ( n1347 , n1309 , n1256 );
    nor g395 ( n1453 , n909 , n1031 );
    nor g396 ( n1055 , n1162 , n1480 );
    nor g397 ( n1145 , n1152 , n1547 );
    and g398 ( n864 , n199 , n1378 );
    or g399 ( n592 , n824 , n385 );
    and g400 ( n685 , n647 , n1555 );
    or g401 ( n100 , n1202 , n555 );
    nor g402 ( n900 , n1374 , n545 );
    not g403 ( n611 , n1647 );
    xnor g404 ( n823 , n1430 , n361 );
    nor g405 ( n1424 , n605 , n959 );
    not g406 ( n352 , n824 );
    or g407 ( n255 , n1494 , n1048 );
    xnor g408 ( n261 , n141 , n949 );
    or g409 ( n1658 , n1032 , n523 );
    not g410 ( n466 , n1592 );
    and g411 ( n91 , n122 , n1005 );
    or g412 ( n621 , n203 , n202 );
    or g413 ( n1283 , n916 , n593 );
    not g414 ( n991 , n692 );
    or g415 ( n21 , n473 , n1174 );
    and g416 ( n858 , n677 , n325 );
    or g417 ( n1514 , n1278 , n1612 );
    and g418 ( n516 , n1472 , n438 );
    nor g419 ( n768 , n1002 , n48 );
    and g420 ( n161 , n1381 , n1606 );
    not g421 ( n671 , n1335 );
    not g422 ( n300 , n1365 );
    or g423 ( n475 , n567 , n1468 );
    or g424 ( n655 , n448 , n13 );
    and g425 ( n242 , n395 , n1580 );
    or g426 ( n520 , n18 , n1595 );
    and g427 ( n1296 , n956 , n230 );
    or g428 ( n204 , n197 , n712 );
    or g429 ( n657 , n1319 , n854 );
    or g430 ( n1661 , n1489 , n1576 );
    not g431 ( n1356 , n611 );
    or g432 ( n110 , n1127 , n59 );
    or g433 ( n449 , n745 , n541 );
    xnor g434 ( n921 , n927 , n672 );
    not g435 ( n1436 , n26 );
    and g436 ( n591 , n995 , n753 );
    nor g437 ( n739 , n1161 , n162 );
    nor g438 ( n1386 , n1255 , n956 );
    and g439 ( n277 , n577 , n1016 );
    or g440 ( n1524 , n39 , n515 );
    or g441 ( n54 , n1155 , n699 );
    or g442 ( n284 , n1443 , n382 );
    and g443 ( n331 , n1343 , n1315 );
    nor g444 ( n496 , n933 , n1544 );
    or g445 ( n748 , n467 , n1582 );
    nor g446 ( n672 , n1158 , n106 );
    or g447 ( n814 , n1214 , n666 );
    not g448 ( n1001 , n1173 );
    not g449 ( n791 , n962 );
    or g450 ( n250 , n1126 , n101 );
    nor g451 ( n487 , n1485 , n1560 );
    buf g452 ( n1026 , n740 );
    nor g453 ( n774 , n861 , n1120 );
    nor g454 ( n764 , n504 , n1601 );
    nor g455 ( n1248 , n1605 , n209 );
    nor g456 ( n1113 , n1427 , n1058 );
    nor g457 ( n126 , n1146 , n1031 );
    not g458 ( n1408 , n35 );
    or g459 ( n1435 , n1217 , n108 );
    and g460 ( n1073 , n1369 , n1515 );
    or g461 ( n499 , n511 , n305 );
    nor g462 ( n1103 , n1024 , n336 );
    nor g463 ( n18 , n934 , n734 );
    or g464 ( n1350 , n278 , n1266 );
    nor g465 ( n1500 , n1391 , n682 );
    or g466 ( n298 , n191 , n583 );
    nor g467 ( n172 , n1629 , n1643 );
    or g468 ( n600 , n685 , n1270 );
    or g469 ( n1256 , n1431 , n547 );
    xnor g470 ( n1072 , n582 , n788 );
    xnor g471 ( n408 , n1372 , n426 );
    nor g472 ( n1584 , n956 , n344 );
    or g473 ( n1634 , n77 , n398 );
    and g474 ( n278 , n361 , n1165 );
    and g475 ( n410 , n832 , n654 );
    buf g476 ( n1442 , n574 );
    or g477 ( n1364 , n1539 , n45 );
    not g478 ( n1535 , n1413 );
    not g479 ( n1090 , n1310 );
    not g480 ( n1537 , n899 );
    not g481 ( n1149 , n1243 );
    not g482 ( n461 , n31 );
    or g483 ( n850 , n1651 , n129 );
    and g484 ( n1387 , n251 , n576 );
    nor g485 ( n180 , n843 , n566 );
    nor g486 ( n953 , n152 , n754 );
    not g487 ( n910 , n1190 );
    not g488 ( n62 , n1403 );
    or g489 ( n779 , n71 , n50 );
    or g490 ( n146 , n1164 , n828 );
    or g491 ( n1492 , n601 , n508 );
    nor g492 ( n873 , n1016 , n1159 );
    nor g493 ( n1586 , n1511 , n1063 );
    and g494 ( n354 , n1368 , n1116 );
    not g495 ( n186 , n1372 );
    nor g496 ( n1662 , n1245 , n968 );
    not g497 ( n868 , n760 );
    nor g498 ( n178 , n1425 , n352 );
    and g499 ( n1489 , n629 , n325 );
    and g500 ( n1433 , n1647 , n1121 );
    or g501 ( n122 , n637 , n237 );
    nor g502 ( n745 , n9 , n227 );
    nor g503 ( n1202 , n1093 , n400 );
    and g504 ( n1169 , n1008 , n283 );
    not g505 ( n10 , n1033 );
    or g506 ( n636 , n708 , n1010 );
    xnor g507 ( n328 , n557 , n1484 );
    and g508 ( n1183 , n1007 , n1005 );
    not g509 ( n115 , n1663 );
    nor g510 ( n1132 , n1388 , n566 );
    and g511 ( n578 , n414 , n938 );
    xnor g512 ( n1484 , n554 , n1546 );
    not g513 ( n152 , n536 );
    not g514 ( n1031 , n1384 );
    or g515 ( n856 , n65 , n436 );
    or g516 ( n170 , n163 , n766 );
    or g517 ( n1319 , n626 , n1501 );
    or g518 ( n1315 , n671 , n832 );
    or g519 ( n1194 , n1629 , n1050 );
    or g520 ( n477 , n2 , n174 );
    or g521 ( n1209 , n1493 , n1419 );
    nor g522 ( n1041 , n1255 , n859 );
    buf g523 ( n154 , n478 );
    or g524 ( n442 , n206 , n88 );
    not g525 ( n915 , n1548 );
    nor g526 ( n963 , n851 , n34 );
    not g527 ( n509 , n1406 );
    or g528 ( n1235 , n1205 , n516 );
    not g529 ( n238 , n507 );
    or g530 ( n302 , n1497 , n17 );
    or g531 ( n1671 , n423 , n1397 );
    nor g532 ( n541 , n285 , n1157 );
    and g533 ( n652 , n877 , n182 );
    not g534 ( n1589 , n889 );
    xnor g535 ( n1009 , n1191 , n961 );
    nor g536 ( n1558 , n1309 , n1003 );
    and g537 ( n249 , n811 , n1005 );
    nor g538 ( n1623 , n222 , n218 );
    and g539 ( n1338 , n412 , n477 );
    xnor g540 ( n1411 , n1614 , n260 );
    and g541 ( n393 , n235 , n84 );
    nor g542 ( n809 , n1255 , n646 );
    and g543 ( n1133 , n1417 , n1420 );
    buf g544 ( n1192 , n1134 );
    not g545 ( n1554 , n366 );
    not g546 ( n1207 , n1534 );
    or g547 ( n1122 , n1510 , n1085 );
    and g548 ( n202 , n681 , n632 );
    nor g549 ( n1252 , n1451 , n1143 );
    buf g550 ( n1117 , n110 );
    nand g551 ( n1574 , n96 , n1150 );
    not g552 ( n994 , n1033 );
    nor g553 ( n755 , n1467 , n11 );
    and g554 ( n430 , n1654 , n1005 );
    and g555 ( n1097 , n1503 , n1655 );
    nor g556 ( n322 , n897 , n640 );
    not g557 ( n735 , n1097 );
    not g558 ( n494 , n1624 );
    xnor g559 ( n879 , n482 , n1257 );
    not g560 ( n1067 , n1448 );
    or g561 ( n680 , n327 , n338 );
    xnor g562 ( n1383 , n1350 , n1447 );
    buf g563 ( n1064 , n1573 );
    or g564 ( n1486 , n1267 , n29 );
    or g565 ( n863 , n1439 , n1325 );
    nor g566 ( n1249 , n765 , n286 );
    nor g567 ( n1048 , n329 , n535 );
    nor g568 ( n92 , n1274 , n135 );
    and g569 ( n892 , n1251 , n325 );
    nor g570 ( n246 , n1213 , n343 );
    not g571 ( n1317 , n1377 );
    and g572 ( n1628 , n167 , n794 );
    nor g573 ( n1080 , n1534 , n1636 );
    xnor g574 ( n738 , n113 , n784 );
    or g575 ( n1231 , n1305 , n791 );
    and g576 ( n1119 , n491 , n1005 );
    buf g577 ( n1023 , n1630 );
    or g578 ( n661 , n945 , n315 );
    and g579 ( n224 , n421 , n1412 );
    and g580 ( n1295 , n94 , n720 );
    nor g581 ( n1225 , n1523 , n1395 );
    nor g582 ( n228 , n1485 , n34 );
    or g583 ( n1314 , n1490 , n357 );
    or g584 ( n265 , n797 , n1244 );
    or g585 ( n1517 , n1273 , n1081 );
    xnor g586 ( n1008 , n1660 , n1483 );
    not g587 ( n1541 , n495 );
    or g588 ( n1490 , n1118 , n1112 );
    not g589 ( n1268 , n84 );
    not g590 ( n573 , n1448 );
    or g591 ( n472 , n1212 , n1340 );
    or g592 ( n766 , n431 , n844 );
    xnor g593 ( n271 , n113 , n16 );
    nor g594 ( n519 , n1108 , n1250 );
    not g595 ( n922 , n857 );
    nor g596 ( n1201 , n704 , n1269 );
    not g597 ( n458 , n859 );
    xnor g598 ( n1380 , n870 , n339 );
    nor g599 ( n1522 , n493 , n35 );
    or g600 ( n190 , n761 , n99 );
    or g601 ( n919 , n1677 , n1423 );
    nor g602 ( n335 , n1098 , n1269 );
    nor g603 ( n1068 , n147 , n865 );
    and g604 ( n48 , n1338 , n1540 );
    nor g605 ( n552 , n386 , n130 );
    and g606 ( n1670 , n585 , n683 );
    nor g607 ( n1494 , n418 , n649 );
    or g608 ( n741 , n335 , n460 );
    not g609 ( n1672 , n590 );
    nor g610 ( n425 , n1366 , n218 );
    nor g611 ( n58 , n435 , n812 );
    or g612 ( n1302 , n912 , n177 );
    and g613 ( n223 , n1251 , n230 );
    or g614 ( n423 , n1322 , n866 );
    not g615 ( n1608 , n905 );
    not g616 ( n1308 , n75 );
    not g617 ( n1285 , n218 );
    and g618 ( n886 , n1675 , n1161 );
    nor g619 ( n1334 , n526 , n668 );
    not g620 ( n1156 , n939 );
    not g621 ( n1230 , n1402 );
    not g622 ( n1245 , n1351 );
    or g623 ( n1395 , n846 , n86 );
    buf g624 ( n1005 , n1445 );
    and g625 ( n1488 , n68 , n1005 );
    nor g626 ( n143 , n1578 , n466 );
    and g627 ( n1357 , n517 , n30 );
    not g628 ( n109 , n1417 );
    and g629 ( n348 , n1551 , n1655 );
    or g630 ( n1421 , n1555 , n234 );
    or g631 ( n1546 , n560 , n1429 );
    nor g632 ( n80 , n1064 , n1652 );
    not g633 ( n762 , n1350 );
    or g634 ( n1506 , n487 , n266 );
    and g635 ( n1002 , n936 , n841 );
    not g636 ( n980 , n569 );
    not g637 ( n1242 , n225 );
    xnor g638 ( n479 , n443 , n299 );
    or g639 ( n1649 , n153 , n1018 );
    or g640 ( n1392 , n288 , n337 );
    nor g641 ( n390 , n1024 , n1532 );
    or g642 ( n993 , n158 , n294 );
    not g643 ( n1173 , n1445 );
    buf g644 ( n663 , n350 );
    buf g645 ( n218 , n1362 );
    or g646 ( n1461 , n173 , n687 );
    or g647 ( n1234 , n646 , n1102 );
    not g648 ( n525 , n57 );
    not g649 ( n406 , n910 );
    not g650 ( n321 , n1044 );
    not g651 ( n162 , n1311 );
    nor g652 ( n1600 , n1311 , n1143 );
    not g653 ( n105 , n1406 );
    not g654 ( n366 , n1564 );
    not g655 ( n674 , n950 );
    not g656 ( n622 , n507 );
    or g657 ( n1625 , n1294 , n755 );
    or g658 ( n1139 , n1353 , n1037 );
    not g659 ( n778 , n1141 );
    nor g660 ( n1643 , n78 , n813 );
    or g661 ( n1284 , n122 , n748 );
    and g662 ( n1385 , n387 , n1530 );
    nor g663 ( n1611 , n1394 , n1169 );
    not g664 ( n1337 , n970 );
    not g665 ( n996 , n661 );
    xnor g666 ( n376 , n811 , n1500 );
    or g667 ( n976 , n1567 , n447 );
    not g668 ( n441 , n750 );
    nor g669 ( n1426 , n238 , n956 );
    nor g670 ( n947 , n198 , n606 );
    nor g671 ( n367 , n769 , n1246 );
    not g672 ( n1568 , n138 );
    nor g673 ( n258 , n67 , n918 );
    not g674 ( n1605 , n507 );
    not g675 ( n1106 , n1300 );
    and g676 ( n480 , n132 , n742 );
    or g677 ( n1599 , n609 , n379 );
    nor g678 ( n551 , n1187 , n400 );
    or g679 ( n1512 , n194 , n257 );
    nor g680 ( n1329 , n51 , n768 );
    or g681 ( n139 , n1066 , n776 );
    not g682 ( n897 , n31 );
    xnor g683 ( n213 , n1611 , n891 );
    not g684 ( n1665 , n1610 );
    nor g685 ( n1464 , n1091 , n406 );
    or g686 ( n1638 , n943 , n420 );
    buf g687 ( n1552 , n478 );
    not g688 ( n1274 , n507 );
    nor g689 ( n1429 , n1243 , n352 );
    nor g690 ( n1236 , n631 , n695 );
    nor g691 ( n214 , n1676 , n1123 );
    nor g692 ( n332 , n198 , n977 );
    or g693 ( n523 , n512 , n405 );
    or g694 ( n1239 , n984 , n988 );
    xnor g695 ( n124 , n1306 , n926 );
    nor g696 ( n874 , n793 , n311 );
    buf g697 ( n565 , n1547 );
    and g698 ( n787 , n431 , n632 );
    nor g699 ( n1376 , n1425 , n935 );
    or g700 ( n318 , n746 , n312 );
    not g701 ( n306 , n1498 );
    not g702 ( n606 , n1143 );
    nor g703 ( n319 , n1240 , n709 );
    or g704 ( n59 , n932 , n1638 );
    not g705 ( n536 , n1307 );
    not g706 ( n134 , n251 );
    or g707 ( n351 , n1258 , n826 );
    xnor g708 ( n1656 , n659 , n1616 );
    nor g709 ( n630 , n1425 , n72 );
    or g710 ( n1138 , n1629 , n1553 );
    and g711 ( n144 , n824 , n325 );
    nor g712 ( n1197 , n300 , n345 );
    or g713 ( n926 , n14 , n1473 );
    xor g714 ( n20 , n661 , n1663 );
    nor g715 ( n40 , n1427 , n490 );
    or g716 ( n1011 , n70 , n600 );
    and g717 ( n1051 , n727 , n1606 );
    nor g718 ( n1228 , n913 , n888 );
    not g719 ( n1127 , n1297 );
    not g720 ( n1336 , n0 );
    xnor g721 ( n439 , n956 , n1143 );
    not g722 ( n1374 , n1405 );
    and g723 ( n77 , n995 , n1555 );
    nor g724 ( n1401 , n596 , n525 );
    not g725 ( n1615 , n1333 );
    or g726 ( n1400 , n1656 , n721 );
    not g727 ( n210 , n212 );
    and g728 ( n33 , n770 , n1515 );
    nor g729 ( n807 , n1311 , n654 );
    and g730 ( n56 , n163 , n632 );
    or g731 ( n521 , n391 , n193 );
    xnor g732 ( n98 , n1352 , n1370 );
    nor g733 ( n1118 , n1162 , n273 );
    nor g734 ( n1452 , n568 , n1507 );
    nor g735 ( n378 , n1621 , n722 );
    buf g736 ( n632 , n771 );
    or g737 ( n614 , n991 , n1622 );
    or g738 ( n982 , n1513 , n1034 );
    not g739 ( n1650 , n939 );
    nor g740 ( n1561 , n1311 , n677 );
    or g741 ( n522 , n1260 , n333 );
    not g742 ( n1227 , n1318 );
    or g743 ( n1382 , n1521 , n942 );
    or g744 ( n310 , n609 , n264 );
    or g745 ( n1142 , n852 , n718 );
    nor g746 ( n1167 , n152 , n1355 );
    and g747 ( n1459 , n1428 , n1549 );
    not g748 ( n640 , n1059 );
    nor g749 ( n200 , n1667 , n562 );
    not g750 ( n397 , n134 );
    or g751 ( n875 , n669 , n1068 );
    not g752 ( n1645 , n980 );
    or g753 ( n1212 , n817 , n58 );
    or g754 ( n1019 , n1104 , n146 );
    nor g755 ( n160 , n1042 , n1261 );
    xnor g756 ( n1028 , n1613 , n136 );
    not g757 ( n893 , n536 );
    nor g758 ( n1115 , n144 , n638 );
    or g759 ( n456 , n1487 , n411 );
    xnor g760 ( n719 , n439 , n879 );
    not g761 ( n847 , n1647 );
    or g762 ( n955 , n27 , n1263 );
    and g763 ( n1205 , n1390 , n147 );
    and g764 ( n1471 , n151 , n950 );
    not g765 ( n1003 , n980 );
    or g766 ( n782 , n309 , n986 );
    nor g767 ( n1328 , n596 , n1004 );
    nor g768 ( n1346 , n1311 , n824 );
    xnor g769 ( n1669 , n1144 , n1444 );
    or g770 ( n413 , n572 , n878 );
    not g771 ( n1175 , n229 );
    not g772 ( n1592 , n1029 );
    not g773 ( n303 , n262 );
    buf g774 ( n253 , n481 );
    not g775 ( n860 , n1610 );
    nor g776 ( n865 , n360 , n830 );
    or g777 ( n173 , n946 , n1132 );
    or g778 ( n625 , n1051 , n831 );
    or g779 ( n240 , n1629 , n723 );
    xnor g780 ( n613 , n659 , n1006 );
    not g781 ( n1172 , n1326 );
    not g782 ( n819 , n1377 );
    and g783 ( n503 , n610 , n79 );
    nor g784 ( n294 , n1102 , n1518 );
    and g785 ( n448 , n1455 , n664 );
    not g786 ( n374 , n652 );
    nor g787 ( n470 , n1456 , n725 );
    or g788 ( n590 , n655 , n80 );
    and g789 ( n6 , n1518 , n325 );
    buf g790 ( n324 , n293 );
    not g791 ( n742 , n932 );
    xnor g792 ( n1640 , n1441 , n1380 );
    not g793 ( n1601 , n1541 );
    or g794 ( n1372 , n799 , n739 );
    or g795 ( n1040 , n25 , n1270 );
    or g796 ( n37 , n458 , n700 );
    not g797 ( n694 , n1281 );
    not g798 ( n350 , n128 );
    or g799 ( n699 , n1491 , n1466 );
    not g800 ( n156 , n218 );
    not g801 ( n446 , n624 );
    not g802 ( n889 , n1355 );
    and g803 ( n1277 , n267 , n632 );
    or g804 ( n639 , n1609 , n520 );
    or g805 ( n1474 , n1629 , n1639 );
    not g806 ( n1610 , n345 );
    xnor g807 ( n407 , n48 , n112 );
    not g808 ( n485 , n503 );
    and g809 ( n1237 , n673 , n37 );
    xor g810 ( n870 , n30 , n1012 );
    or g811 ( n1641 , n223 , n226 );
    or g812 ( n650 , n1401 , n1505 );
    nor g813 ( n369 , n661 , n459 );
    nor g814 ( n103 , n1581 , n273 );
    and g815 ( n1504 , n209 , n325 );
    nor g816 ( n817 , n710 , n819 );
    or g817 ( n1571 , n552 , n308 );
    or g818 ( n821 , n1623 , n1486 );
    or g819 ( n1642 , n1453 , n876 );
    nor g820 ( n612 , n1056 , n1113 );
    or g821 ( n653 , n1526 , n700 );
    nor g822 ( n1449 , n1374 , n686 );
    not g823 ( n1034 , n597 );
    and g824 ( n775 , n1264 , n1005 );
    not g825 ( n958 , n730 );
    or g826 ( n666 , n214 , n937 );
    not g827 ( n420 , n647 );
    not g828 ( n1195 , n853 );
    and g829 ( n1668 , n251 , n1648 );
    nor g830 ( n708 , n938 , n188 );
    not g831 ( n1544 , n57 );
    not g832 ( n777 , n1563 );
    nor g833 ( n555 , n1129 , n392 );
    not g834 ( n1044 , n1333 );
    not g835 ( n999 , n1518 );
    nor g836 ( n1158 , n403 , n612 );
    buf g837 ( n678 , n623 );
    buf g838 ( n388 , n1013 );
    or g839 ( n392 , n36 , n56 );
    or g840 ( n114 , n807 , n410 );
    nor g841 ( n248 , n1425 , n1105 );
    not g842 ( n344 , n365 );
    xnor g843 ( n453 , n1236 , n580 );
    and g844 ( n52 , n499 , n769 );
    or g845 ( n452 , n1586 , n1167 );
    nor g846 ( n95 , n1165 , n1458 );
    and g847 ( n39 , n1407 , n1243 );
    not g848 ( n207 , n348 );
    not g849 ( n31 , n1172 );
    nor g850 ( n903 , n531 , n92 );
    nor g851 ( n795 , n1324 , n624 );
    and g852 ( n102 , n1030 , n230 );
    or g853 ( n409 , n157 , n966 );
    and g854 ( n559 , n1285 , n1508 );
    not g855 ( n1213 , n730 );
    nor g856 ( n1082 , n470 , n1472 );
    or g857 ( n1241 , n407 , n409 );
    or g858 ( n3 , n1328 , n1197 );
    nor g859 ( n603 , n120 , n1661 );
    nor g860 ( n831 , n1606 , n935 );
    or g861 ( n562 , n595 , n1486 );
    buf g862 ( n608 , n1596 );
    nor g863 ( n450 , n215 , n1060 );
    not g864 ( n1455 , n218 );
    not g865 ( n236 , n365 );
    or g866 ( n1096 , n979 , n1488 );
    not g867 ( n166 , n1230 );
    xnor g868 ( n1370 , n921 , n408 );
    or g869 ( n840 , n1629 , n534 );
    nor g870 ( n308 , n10 , n345 );
    nor g871 ( n428 , n1425 , n1053 );
    nor g872 ( n508 , n198 , n55 );
    and g873 ( n1290 , n1153 , n182 );
    or g874 ( n643 , n589 , n1662 );
    xnor g875 ( n252 , n1435 , n1108 );
    and g876 ( n1066 , n1460 , n1049 );
    not g877 ( n358 , n1001 );
    and g878 ( n983 , n796 , n589 );
    or g879 ( n1354 , n252 , n1171 );
    nor g880 ( n1458 , n1653 , n40 );
    and g881 ( n987 , n1223 , n1606 );
    not g882 ( n1004 , n868 );
    not g883 ( n1536 , n1432 );
    and g884 ( n838 , n1338 , n1663 );
    nor g885 ( n1607 , n1280 , n311 );
    not g886 ( n1520 , n394 );
    not g887 ( n604 , n509 );
    not g888 ( n707 , n182 );
    xnor g889 ( n241 , n1452 , n636 );
    nor g890 ( n1664 , n1425 , n1545 );
    not g891 ( n855 , n1545 );
    xnor g892 ( n1444 , n564 , n850 );
    xnor g893 ( n528 , n1569 , n175 );
    or g894 ( n383 , n1387 , n1222 );
    nor g895 ( n433 , n1581 , n1123 );
    not g896 ( n148 , n306 );
    nor g897 ( n830 , n1425 , n55 );
    not g898 ( n530 , n229 );
    nand g899 ( n790 , n1562 , n128 );
    nor g900 ( n539 , n769 , n1228 );
    xor g901 ( n1035 , n1447 , n823 );
    not g902 ( n1448 , n1379 );
    not g903 ( n760 , n1193 );
    or g904 ( n312 , n1229 , n970 );
    not g905 ( n42 , n1318 );
    and g906 ( n276 , n646 , n325 );
    or g907 ( n1588 , n452 , n1642 );
    or g908 ( n1174 , n1579 , n907 );
    or g909 ( n712 , n1069 , n377 );
    not g910 ( n1318 , n994 );
    nor g911 ( n263 , n622 , n1030 );
    or g912 ( n1196 , n1245 , n982 );
    and g913 ( n372 , n801 , n1196 );
    nor g914 ( n457 , n346 , n827 );
    or g915 ( n78 , n1433 , n1291 );
    not g916 ( n960 , n507 );
    nor g917 ( n465 , n604 , n316 );
    or g918 ( n1616 , n873 , n643 );
    not g919 ( n1456 , n274 );
    or g920 ( n363 , n808 , n1220 );
    not g921 ( n1286 , n1190 );
    or g922 ( n76 , n1629 , n1588 );
    and g923 ( n338 , n331 , n1005 );
    nor g924 ( n243 , n468 , n1317 );
    xor g925 ( n359 , n1101 , n438 );
    or g926 ( n1591 , n1583 , n599 );
    not g927 ( n336 , n446 );
    xnor g928 ( n1332 , n1617 , n20 );
    not g929 ( n1360 , n63 );
    nor g930 ( n944 , n1184 , n1544 );
    and g931 ( n553 , n271 , n632 );
    not g932 ( n391 , n1240 );
    xnor g933 ( n1420 , n1572 , n950 );
    nor g934 ( n1391 , n184 , n450 );
    or g935 ( n197 , n802 , n1312 );
    or g936 ( n1550 , n160 , n119 );
    xnor g937 ( n1006 , n1159 , n234 );
    not g938 ( n1087 , n293 );
    not g939 ( n951 , n446 );
    not g940 ( n462 , n252 );
    not g941 ( n435 , n105 );
    nor g942 ( n1124 , n923 , n374 );
    nor g943 ( n53 , n479 , n1368 );
    or g944 ( n414 , n314 , n211 );
    not g945 ( n1667 , n1300 );
    nor g946 ( n568 , n147 , n1136 );
    nor g947 ( n1263 , n494 , n887 );
    not g948 ( n1152 , n1606 );
    nor g949 ( n866 , n285 , n250 );
    nor g950 ( n164 , n617 , n1426 );
    xnor g951 ( n482 , n1030 , n1251 );
    nor g952 ( n584 , n710 , n1022 );
    xnor g953 ( n1321 , n654 , n490 );
    nor g954 ( n878 , n1062 , n503 );
    nor g955 ( n266 , n893 , n394 );
    nor g956 ( n411 , n1106 , n434 );
    nor g957 ( n334 , n329 , n1665 );
    nor g958 ( n90 , n1243 , n884 );
    or g959 ( n361 , n987 , n85 );
    not g960 ( n1451 , n365 );
    not g961 ( n179 , n705 );
    not g962 ( n280 , n48 );
    and g963 ( n1379 , n1535 , n989 );
    nor g964 ( n1306 , n733 , n1674 );
    nor g965 ( n802 , n362 , n321 );
    or g966 ( n257 , n87 , n703 );
    or g967 ( n74 , n744 , n1519 );
    nor g968 ( n1673 , n417 , n603 );
    not g969 ( n665 , n1568 );
    nor g970 ( n279 , n67 , n1004 );
    or g971 ( n323 , n1571 , n581 );
    and g972 ( n556 , n522 , n1479 );
    not g973 ( n992 , n149 );
    or g974 ( n269 , n456 , n767 );
    not g975 ( n127 , n1389 );
    or g976 ( n569 , n89 , n553 );
    not g977 ( n1024 , n1342 );
    and g978 ( n1585 , n1030 , n325 );
    nor g979 ( n498 , n290 , n1175 );
    not g980 ( n1513 , n1271 );
    nor g981 ( n239 , n198 , n855 );
    not g982 ( n1300 , n1172 );
    or g983 ( n633 , n3 , n1649 );
    nor g984 ( n709 , n858 , n1178 );
    nor g985 ( n355 , n1479 , n164 );
    not g986 ( n1467 , n393 );
    and g987 ( n833 , n1285 , n1131 );
    not g988 ( n1157 , n1233 );
    xnor g989 ( n1111 , n1575 , n1161 );
    xnor g990 ( n368 , n693 , n930 );
    nor g991 ( n537 , n950 , n542 );
    xor g992 ( n679 , n1661 , n331 );
    and g993 ( n1222 , n1428 , n1052 );
    not g994 ( n998 , n1030 );
    nor g995 ( n88 , n1227 , n250 );
    nor g996 ( n1533 , n504 , n624 );
    or g997 ( n1089 , n634 , n255 );
    xnor g998 ( n792 , n587 , n804 );
    or g999 ( n1029 , n139 , n317 );
    or g1000 ( n1566 , n1633 , n1558 );
    not g1001 ( n1102 , n365 );
    or g1002 ( n563 , n471 , n486 );
    not g1003 ( n1590 , n1411 );
    not g1004 ( n1086 , n1606 );
    nor g1005 ( n436 , n42 , n1345 );
    or g1006 ( n1216 , n1078 , n575 );
    not g1007 ( n235 , n726 );
    and g1008 ( n852 , n648 , n635 );
    nor g1009 ( n1206 , n1324 , n495 );
    nor g1010 ( n307 , n1578 , n781 );
    xnor g1011 ( n1144 , n743 , n234 );
    xor g1012 ( n155 , n51 , n738 );
    and g1013 ( n49 , n1025 , n1606 );
    or g1014 ( n1639 , n1566 , n1083 );
    nor g1015 ( n17 , n303 , n1355 );
    or g1016 ( n225 , n127 , n384 );
    nor g1017 ( n340 , n463 , n495 );
    not g1018 ( n1358 , n403 );
    and g1019 ( n1473 , n1040 , n1640 );
    nor g1020 ( n1092 , n1462 , n1385 );
    or g1021 ( n326 , n498 , n1666 );
    not g1022 ( n1646 , n770 );
    not g1023 ( n757 , n1360 );
    and g1024 ( n1114 , n929 , n1475 );
    xnor g1025 ( n975 , n554 , n765 );
    not g1026 ( n1289 , n676 );
    nor g1027 ( n237 , n938 , n440 );
    not g1028 ( n1603 , n1351 );
    nor g1029 ( n14 , n1299 , n1040 );
    not g1030 ( n984 , n1150 );
    or g1031 ( n1622 , n429 , n1207 );
    or g1032 ( n455 , n881 , n1349 );
    xnor g1033 ( n681 , n527 , n1231 );
    or g1034 ( n691 , n619 , n15 );
    or g1035 ( n743 , n798 , n1057 );
    and g1036 ( n885 , n1460 , n1189 );
    nor g1037 ( n502 , n463 , n951 );
    or g1038 ( n732 , n1644 , n1252 );
    not g1039 ( n570 , n996 );
    not g1040 ( n11 , n1440 );
    not g1041 ( n693 , n627 );
    or g1042 ( n812 , n871 , n1277 );
    or g1043 ( n1390 , n1450 , n1363 );
    nor g1044 ( n474 , n435 , n469 );
    not g1045 ( n959 , n1436 );
    nor g1046 ( n1462 , n1530 , n1115 );
    nor g1047 ( n548 , n461 , n244 );
    and g1048 ( n669 , n1641 , n147 );
    not g1049 ( n1164 , n1630 );
    nor g1050 ( n1293 , n1361 , n374 );
    xnor g1051 ( n136 , n135 , n824 );
    or g1052 ( n585 , n1378 , n1415 );
    not g1053 ( n1309 , n1379 );
    not g1054 ( n301 , n113 );
    nor g1055 ( n626 , n1389 , n19 );
    nor g1056 ( n377 , n461 , n590 );
    not g1057 ( n1675 , n1606 );
    or g1058 ( n1469 , n419 , n372 );
    and g1059 ( n941 , n1455 , n716 );
    not g1060 ( n1059 , n250 );
    and g1061 ( n914 , n60 , n1620 );
    xnor g1062 ( n1652 , n1308 , n246 );
    or g1063 ( n723 , n1182 , n1506 );
    and g1064 ( n979 , n395 , n233 );
    nor g1065 ( n1569 , n597 , n846 );
    not g1066 ( n1457 , n316 );
    and g1067 ( n776 , n191 , n1005 );
    nor g1068 ( n460 , n974 , n1204 );
    not g1069 ( n843 , n509 );
    nor g1070 ( n1415 , n809 , n428 );
    or g1071 ( n1171 , n43 , n217 );
    nor g1072 ( n129 , n1606 , n999 );
    or g1073 ( n978 , n74 , n1084 );
    not g1074 ( n1120 , n1541 );
    not g1075 ( n229 , n207 );
    not g1076 ( n1063 , n910 );
    nor g1077 ( n620 , n895 , n445 );
    and g1078 ( n1057 , n1086 , n1575 );
    or g1079 ( n581 , n1424 , n1347 );
    or g1080 ( n288 , n258 , n1103 );
    nor g1081 ( n1081 , n346 , n1589 );
    or g1082 ( n1659 , n485 , n778 );
    xnor g1083 ( n157 , n125 , n779 );
    not g1084 ( n648 , n218 );
    or g1085 ( n1232 , n1148 , n1675 );
    nor g1086 ( n341 , n1064 , n213 );
    xnor g1087 ( n896 , n1101 , n924 );
    nor g1088 ( n1077 , n981 , n1626 );
    or g1089 ( n705 , n922 , n1207 );
    xnor g1090 ( n113 , n254 , n1240 );
    or g1091 ( n1298 , n1133 , n1080 );
    or g1092 ( n554 , n1100 , n12 );
    or g1093 ( n827 , n1096 , n1020 );
    or g1094 ( n1126 , n833 , n775 );
    not g1095 ( n977 , n859 );
    nor g1096 ( n1075 , n1064 , n1337 );
    not g1097 ( n940 , n1110 );
    nor g1098 ( n1341 , n1070 , n1259 );
    not g1099 ( n744 , n785 );
    not g1100 ( n935 , n1058 );
    xnor g1101 ( n763 , n399 , n1111 );
    and g1102 ( n770 , n726 , n84 );
    xnor g1103 ( n557 , n1038 , n254 );
    and g1104 ( n645 , n216 , n632 );
    or g1105 ( n1553 , n782 , n955 );
    not g1106 ( n1621 , n1326 );
    not g1107 ( n133 , n812 );
    not g1108 ( n948 , n198 );
    not g1109 ( n1351 , n187 );
    not g1110 ( n908 , n1646 );
    and g1111 ( n1078 , n60 , n1418 );
    and g1112 ( n997 , n1348 , n1413 );
    and g1113 ( n1094 , n850 , n769 );
    nor g1114 ( n533 , n1608 , n827 );
    xnor g1115 ( n426 , n281 , n1570 );
    nor g1116 ( n1218 , n1274 , n1251 );
    not g1117 ( n1259 , n397 );
    not g1118 ( n832 , n198 );
    xor g1119 ( n149 , n564 , n1378 );
    or g1120 ( n217 , n915 , n47 );
    or g1121 ( n957 , n586 , n219 );
    and g1122 ( n251 , n1537 , n270 );
    or g1123 ( n767 , n1224 , n533 );
    not g1124 ( n379 , n725 );
    not g1125 ( n1377 , n611 );
    nor g1126 ( n153 , n1014 , n668 );
    xnor g1127 ( n594 , n414 , n1390 );
    and g1128 ( n1501 , n114 , n1389 );
    nor g1129 ( n567 , n923 , n530 );
    nor g1130 ( n5 , n1129 , n928 );
    not g1131 ( n1587 , n566 );
    not g1132 ( n1233 , n1283 );
    nor g1133 ( n159 , n1438 , n1204 );
    not g1134 ( n1381 , n574 );
    not g1135 ( n63 , n997 );
    nor g1136 ( n967 , n1425 , n458 );
    and g1137 ( n1141 , n389 , n1538 );
    or g1138 ( n429 , n881 , n720 );
    nor g1139 ( n752 , n1425 , n606 );
    or g1140 ( n1221 , n898 , n334 );
    not g1141 ( n697 , n1572 );
    not g1142 ( n1186 , n692 );
    and g1143 ( n799 , n1161 , n198 );
    not g1144 ( n920 , n1302 );
    not g1145 ( n311 , n1193 );
    nor g1146 ( n12 , n1243 , n1105 );
    and g1147 ( n1305 , n1516 , n857 );
    or g1148 ( n711 , n551 , n340 );
    and g1149 ( n205 , n1210 , n403 );
    not g1150 ( n46 , n1670 );
    nor g1151 ( n883 , n1386 , n630 );
    not g1152 ( n256 , n825 );
    not g1153 ( n1404 , n1247 );
    nor g1154 ( n492 , n358 , n1141 );
    or g1155 ( n177 , n1565 , n341 );
    or g1156 ( n616 , n906 , n1301 );
    and g1157 ( n641 , n993 , n769 );
    and g1158 ( n690 , n1268 , n235 );
    nor g1159 ( n1027 , n1425 , n884 );
    and g1160 ( n912 , n901 , n1065 );
    or g1161 ( n1021 , n476 , n1514 );
    xnor g1162 ( n1299 , n1383 , n1076 );
    and g1163 ( n1365 , n488 , n1503 );
    not g1164 ( n1074 , n1034 );
    not g1165 ( n167 , n899 );
    and g1166 ( n1254 , n696 , n393 );
    not g1167 ( n292 , n1134 );
    and g1168 ( n1539 , n135 , n230 );
    nor g1169 ( n171 , n1187 , n189 );
    xnor g1170 ( n399 , n646 , n1518 );
    or g1171 ( n658 , n501 , n1533 );
    and g1172 ( n1125 , n545 , n1033 );
    nor g1173 ( n601 , n1311 , n1251 );
    or g1174 ( n1431 , n1168 , n1183 );
    not g1175 ( n1367 , n1001 );
    not g1176 ( n1053 , n646 );
    xnor g1177 ( n1327 , n1522 , n359 );
    xnor g1178 ( n299 , n1617 , n1282 );
    not g1179 ( n1016 , n1555 );
    and g1180 ( n295 , n1058 , n230 );
    not g1181 ( n609 , n381 );
    and g1182 ( n44 , n1149 , n677 );
    not g1183 ( n1200 , n664 );
    and g1184 ( n1265 , n762 , n730 );
    xnor g1185 ( n1271 , n161 , n1545 );
    not g1186 ( n881 , n301 );
    not g1187 ( n26 , n1369 );
    not g1188 ( n796 , n659 );
    xnor g1189 ( n676 , n328 , n1009 );
    nor g1190 ( n1423 , n1410 , n696 );
    not g1191 ( n905 , n66 );
    or g1192 ( n583 , n549 , n46 );
    not g1193 ( n212 , n686 );
    or g1194 ( n89 , n1114 , n249 );
    not g1195 ( n272 , n105 );
    nor g1196 ( n510 , n1255 , n824 );
    nor g1197 ( n898 , n386 , n1199 );
    not g1198 ( n264 , n1563 );
    nor g1199 ( n561 , n1255 , n1143 );
    or g1200 ( n1470 , n1606 , n671 );
    nor g1201 ( n662 , n958 , n181 );
    or g1202 ( n82 , n872 , n1179 );
    or g1203 ( n1151 , n1577 , n803 );
    or g1204 ( n316 , n680 , n1075 );
    not g1205 ( n722 , n1457 );
    nor g1206 ( n1393 , n1608 , n1262 );
    and g1207 ( n195 , n648 , n1303 );
    xnor g1208 ( n1226 , n1271 , n1225 );
    or g1209 ( n1538 , n1493 , n1237 );
    not g1210 ( n497 , n994 );
    or g1211 ( n651 , n963 , n502 );
    not g1212 ( n929 , n218 );
    nor g1213 ( n1278 , n330 , n1259 );
    or g1214 ( n566 , n185 , n972 );
    and g1215 ( n1203 , n467 , n1005 );
    or g1216 ( n619 , n1061 , n247 );
    nor g1217 ( n349 , n418 , n62 );
    xnor g1218 ( n1627 , n1092 , n957 );
    nor g1219 ( n1267 , n1536 , n98 );
    or g1220 ( n689 , n1135 , n1125 );
    nor g1221 ( n101 , n1064 , n729 );
    not g1222 ( n424 , n868 );
    nor g1223 ( n108 , n1243 , n606 );
    xnor g1224 ( n729 , n911 , n1130 );
    not g1225 ( n221 , n262 );
    not g1226 ( n1137 , n1097 );
    not g1227 ( n1560 , n1286 );
    or g1228 ( n412 , n1186 , n109 );
    and g1229 ( n749 , n353 , n1479 );
    xnor g1230 ( n1660 , n1327 , n546 );
    or g1231 ( n628 , n1176 , n332 );
    nor g1232 ( n1579 , n362 , n227 );
    or g1233 ( n871 , n941 , n422 );
    or g1234 ( n624 , n287 , n645 );
    xnor g1235 ( n970 , n1213 , n343 );
    not g1236 ( n968 , n731 );
    not g1237 ( n800 , n629 );
    or g1238 ( n1559 , n1201 , n159 );
    and g1239 ( n942 , n948 , n490 );
    nor g1240 ( n27 , n1093 , n189 );
    not g1241 ( n70 , n762 );
    not g1242 ( n1503 , n1551 );
    and g1243 ( n371 , n1319 , n1005 );
    not g1244 ( n1345 , n212 );
    not g1245 ( n451 , n497 );
    or g1246 ( n68 , n880 , n1249 );
    not g1247 ( n138 , n1369 );
    and g1248 ( n417 , n1200 , n120 );
    not g1249 ( n1478 , n1672 );
    nor g1250 ( n1595 , n494 , n621 );
    or g1251 ( n687 , n111 , n457 );
    not g1252 ( n488 , n1655 );
    and g1253 ( n599 , n1149 , n268 );
    and g1254 ( n826 , n1652 , n120 );
    nor g1255 ( n1612 , n990 , n148 );
    not g1256 ( n1534 , n217 );
    and g1257 ( n1180 , n1276 , n1396 );
    nor g1258 ( n1353 , n909 , n670 );
    or g1259 ( n924 , n179 , n1417 );
    or g1260 ( n1264 , n95 , n22 );
    and g1261 ( n637 , n41 , n938 );
    xor g1262 ( n274 , n414 , n938 );
    xnor g1263 ( n1128 , n613 , n528 );
    not g1264 ( n1564 , n274 );
    or g1265 ( n357 , n1602 , n390 );
    and g1266 ( n647 , n591 , n1603 );
    not g1267 ( n773 , n652 );
    not g1268 ( n1410 , n905 );
    xnor g1269 ( n659 , n850 , n769 );
    nor g1270 ( n816 , n793 , n259 );
    xnor g1271 ( n527 , n1524 , n1479 );
    and g1272 ( n931 , n109 , n777 );
    nor g1273 ( n1260 , n1311 , n956 );
    or g1274 ( n1032 , n441 , n1087 );
    not g1275 ( n853 , n1402 );
    or g1276 ( n131 , n896 , n1241 );
    nor g1277 ( n571 , n381 , n1456 );
    not g1278 ( n1304 , n550 );
    buf g1279 ( n1556 , n829 );
    and g1280 ( n575 , n875 , n1005 );
    and g1281 ( n317 , n1656 , n632 );
    buf g1282 ( n234 , n297 );
    and g1283 ( n1291 , n562 , n690 );
    nor g1284 ( n188 , n1585 , n263 );
    or g1285 ( n867 , n607 , n953 );
    xnor g1286 ( n118 , n1304 , n1082 );
    nor g1287 ( n1330 , n198 , n998 );
    or g1288 ( n1038 , n1017 , n602 );
    not g1289 ( n1155 , n1652 );
    not g1290 ( n939 , n760 );
    not g1291 ( n1532 , n1557 );
    or g1292 ( n1430 , n49 , n904 );
    xnor g1293 ( n546 , n756 , n310 );
    or g1294 ( n51 , n1414 , n369 );
    nor g1295 ( n1527 , n276 , n1316 );
    not g1296 ( n692 , n252 );
    or g1297 ( n64 , n952 , n919 );
    xnor g1298 ( n1463 , n282 , n1597 );
    not g1299 ( n8 , n1150 );
    nor g1300 ( n1208 , n1311 , n1058 );
    and g1301 ( n1674 , n1072 , n1 );
    or g1302 ( n1182 , n810 , n474 );
    not g1303 ( n285 , n1281 );
    nor g1304 ( n440 , n806 , n1598 );
    not g1305 ( n899 , n224 );
    not g1306 ( n1406 , n690 );
    nor g1307 ( n937 , n221 , n392 );
    nor g1308 ( n501 , n851 , n406 );
    and g1309 ( n1414 , n1546 , n1530 );
    not g1310 ( n1348 , n989 );
    nor g1311 ( n247 , n694 , n812 );
    or g1312 ( n820 , n784 , n936 );
    nor g1313 ( n1323 , n689 , n505 );
    nor g1314 ( n538 , n1479 , n883 );
    not g1315 ( n627 , n1155 );
    or g1316 ( n1355 , n1216 , n201 );
    or g1317 ( n673 , n859 , n1451 );
    or g1318 ( n15 , n396 , n1206 );
    not g1319 ( n668 , n348 );
    not g1320 ( n1177 , n1592 );
    or g1321 ( n758 , n816 , n73 );
    not g1322 ( n346 , n1067 );
    nor g1323 ( n1677 , n1280 , n259 );
    and g1324 ( n1325 , n846 , n1271 );
    not g1325 ( n1403 , n63 );
    xnor g1326 ( n1352 , n679 , n1107 );
    buf g1327 ( n61 , n845 );
    and g1328 ( n1446 , n592 , n653 );
    not g1329 ( n544 , n1044 );
    not g1330 ( n273 , n853 );
    or g1331 ( n564 , n1618 , n529 );
    nor g1332 ( n602 , n1243 , n977 );
    and g1333 ( n547 , n896 , n632 );
    and g1334 ( n798 , n1606 , n588 );
    buf g1335 ( n489 , n350 );
    not g1336 ( n196 , n827 );
    not g1337 ( n1110 , n784 );
    and g1338 ( n642 , n549 , n1005 );
    xnor g1339 ( n784 , n1038 , n184 );
    xnor g1340 ( n1045 , n381 , n1235 );
    not g1341 ( n395 , n218 );
    or g1342 ( n813 , n33 , n1254 );
    not g1343 ( n1297 , n958 );
    not g1344 ( n1498 , n1428 );
    or g1345 ( n549 , n1088 , n1664 );
    not g1346 ( n1526 , n824 );
    not g1347 ( n30 , n911 );
    and g1348 ( n1326 , n707 , n1153 );
    or g1349 ( n337 , n1509 , n378 );
    xnor g1350 ( n785 , n1028 , n719 );
    or g1351 ( n505 , n1073 , n370 );
    nor g1352 ( n211 , n1243 , n998 );
    not g1353 ( n731 , n992 );
    nor g1354 ( n783 , n236 , n209 );
    or g1355 ( n780 , n1561 , n1279 );
    nor g1356 ( n1136 , n892 , n1218 );
    not g1357 ( n928 , n1557 );
    and g1358 ( n595 , n837 , n1065 );
    xnor g1359 ( n1047 , n1513 , n753 );
    not g1360 ( n384 , n1430 );
    and g1361 ( n1168 , n1465 , n432 );
    or g1362 ( n841 , n975 , n459 );
    xor g1363 ( n925 , n991 , n1548 );
    not g1364 ( n291 , n133 );
    or g1365 ( n353 , n1296 , n1584 );
    not g1366 ( n995 , n982 );
    nor g1367 ( n1509 , n1373 , n773 );
    and g1368 ( n513 , n157 , n632 );
    nor g1369 ( n1521 , n1311 , n490 );
    not g1370 ( n1460 , n218 );
    and g1371 ( n724 , n1469 , n1054 );
    or g1372 ( n686 , n1142 , n667 );
    and g1373 ( n158 , n1518 , n230 );
    nor g1374 ( n1000 , n818 , n1650 );
    not g1375 ( n1270 , n724 );
    nor g1376 ( n16 , n1295 , n834 );
    xnor g1377 ( n1597 , n1395 , n234 );
    not g1378 ( n315 , n554 );
    xnor g1379 ( n1637 , n35 , n925 );
    not g1380 ( n1388 , n497 );
    or g1381 ( n38 , n126 , n180 );
    and g1382 ( n1279 , n948 , n677 );
    and g1383 ( n215 , n859 , n325 );
    not g1384 ( n1495 , n1530 );
    xnor g1385 ( n459 , n1546 , n1530 );
    or g1386 ( n380 , n496 , n1393 );
    or g1387 ( n1054 , n1358 , n1288 );
    nor g1388 ( n660 , n1311 , n209 );
    nor g1389 ( n1666 , n303 , n675 );
    not g1390 ( n1104 , n829 );
    nor g1391 ( n1363 , n1243 , n55 );
    nor g1392 ( n305 , n198 , n999 );
    nor g1393 ( n1528 , n869 , n1673 );
    and g1394 ( n1523 , n1074 , n1555 );
    or g1395 ( n176 , n660 , n1188 );
    not g1396 ( n1101 , n462 );
    not g1397 ( n943 , n1357 );
    not g1398 ( n405 , n296 );
    and g1399 ( n577 , n149 , n1603 );
    and g1400 ( n904 , n1086 , n654 );
    not g1401 ( n1482 , n1420 );
    nor g1402 ( n404 , n1030 , n344 );
    nor g1403 ( n772 , n1255 , n1058 );
    nor g1404 ( n1312 , n861 , n569 );
    buf g1405 ( n1542 , n750 );
    not g1406 ( n845 , n128 );
    and g1407 ( n917 , n209 , n230 );
    not g1408 ( n945 , n765 );
    and g1409 ( n1543 , n780 , n1240 );
    xnor g1410 ( n1116 , n155 , n1332 );
    not g1411 ( n1563 , n1482 );
    xnor g1412 ( n1614 , n1109 , n1321 );
    not g1413 ( n535 , n1672 );
    nor g1414 ( n192 , n1467 , n569 );
    and g1415 ( n1056 , n1058 , n325 );
    not g1416 ( n1624 , n1307 );
    and g1417 ( n572 , n156 , n973 );
    buf g1418 ( n142 , n614 );
    nor g1419 ( n1266 , n225 , n911 );
    not g1420 ( n696 , n920 );
    or g1421 ( n969 , n1208 , n1287 );
    not g1422 ( n193 , n254 );
    not g1423 ( n656 , n1084 );
    not g1424 ( n918 , n1615 );
    or g1425 ( n36 , n195 , n91 );
    and g1426 ( n1017 , n137 , n1243 );
    nor g1427 ( n1598 , n1425 , n998 );
    or g1428 ( n916 , n642 , n885 );
    and g1429 ( n1445 , n1071 , n558 );
    or g1430 ( n932 , n1145 , n702 );
    nor g1431 ( n1176 , n1311 , n859 );
    not g1432 ( n1166 , n562 );
    or g1433 ( n1573 , n1065 , n558 );
    not g1434 ( n1071 , n1065 );
    not g1435 ( n1405 , n518 );
    not g1436 ( n469 , n1059 );
    or g1437 ( n1572 , n1525 , n90 );
    nor g1438 ( n1238 , n934 , n1477 );
    or g1439 ( n1349 , n1295 , n838 );
    or g1440 ( n1198 , n302 , n684 );
    or g1441 ( n345 , n715 , n123 );
    or g1442 ( n715 , n914 , n1119 );
    and g1443 ( n1481 , n1012 , n225 );
    or g1444 ( n1160 , n1629 , n815 );
    xnor g1445 ( n804 , n822 , n688 );
    xnor g1446 ( n1441 , n1447 , n181 );
    nor g1447 ( n756 , n1516 , n791 );
    nor g1448 ( n1069 , n526 , n773 );
    not g1449 ( n1147 , n1661 );
    or g1450 ( n1362 , n532 , n1071 );
    not g1451 ( n329 , n690 );
    and g1452 ( n86 , n597 , n234 );
    or g1453 ( n1582 , n875 , n1476 );
    nor g1454 ( n1602 , n9 , n544 );
    not g1455 ( n1281 , n518 );
    and g1456 ( n132 , n1095 , n1265 );
    xnor g1457 ( n267 , n234 , n1555 );
    and g1458 ( n593 , n1226 , n632 );
    not g1459 ( n771 , n1573 );
    not g1460 ( n1440 , n1256 );
    not g1461 ( n189 , n908 );
    not g1462 ( n262 , n1137 );
    or g1463 ( n740 , n1668 , n1459 );
    and g1464 ( n483 , n855 , n325 );
    or g1465 ( n491 , n205 , n862 );
    nor g1466 ( n586 , n765 , n903 );
    or g1467 ( n1036 , n563 , n758 );
    not g1468 ( n1261 , n1230 );
    not g1469 ( n244 , n133 );
    or g1470 ( n97 , n380 , n1550 );
    nor g1471 ( n375 , n1373 , n530 );
    and g1472 ( n1663 , n820 , n1209 );
    buf g1473 ( n364 , n842 );
    not g1474 ( n1548 , n527 );
    or g1475 ( n634 , n1464 , n192 );
    not g1476 ( n1480 , n701 );
    or g1477 ( n891 , n354 , n53 );
    and g1478 ( n13 , n761 , n1005 );
    and g1479 ( n713 , n732 , n1108 );
    nor g1480 ( n422 , n1536 , n1372 );
    nor g1481 ( n119 , n1106 , n1029 );
    not g1482 ( n1123 , n348 );
    or g1483 ( n389 , n184 , n1015 );
    or g1484 ( n803 , n279 , n985 );
    or g1485 ( n1529 , n1219 , n711 );
    not g1486 ( n476 , n1150 );
    not g1487 ( n971 , n1233 );
    nor g1488 ( n1037 , n1388 , n1029 );
    not g1489 ( n701 , n207 );
    nor g1490 ( n1439 , n855 , n161 );
    or g1491 ( n381 , n674 , n697 );
    or g1492 ( n988 , n1341 , n1163 );
    nor g1493 ( n718 , n1367 , n1670 );
    not g1494 ( n1262 , n889 );
    and g1495 ( n201 , n118 , n632 );
    nor g1496 ( n1487 , n290 , n166 );
    not g1497 ( n700 , n230 );
    or g1498 ( n437 , n491 , n298 );
    nor g1499 ( n245 , n510 , n178 );
endmodule
