module top( n4 , n37 , n44 , n56 , n66 , n84 , n88 , n132 , n181 , 
n185 , n196 , n220 , n274 , n308 , n335 , n422 , n493 , n504 , n523 , 
n530 , n642 , n670 , n705 , n722 , n770 , n772 , n794 , n824 , n829 , 
n835 , n850 , n866 , n872 , n873 , n891 , n927 , n928 , n935 , n940 , 
n944 , n955 , n1066 , n1103 , n1140 , n1156 , n1157 , n1202 , n1229 , n1234 , 
n1240 , n1273 , n1280 , n1361 , n1367 , n1387 , n1398 , n1404 , n1432 , n1507 , 
n1521 , n1540 , n1541 , n1638 , n1646 , n1761 , n1775 , n1793 , n1808 , n1820 , 
n1861 , n1874 , n1889 , n1938 , n2031 , n2050 , n2055 , n2073 , n2110 , n2112 , 
n2165 , n2195 , n2223 , n2252 , n2258 , n2313 , n2324 , n2371 , n2385 , n2402 , 
n2463 , n2490 , n2514 , n2523 , n2567 , n2572 , n2622 , n2640 , n2664 , n2724 , 
n2727 , n2744 , n2757 , n2760 , n2806 , n2830 , n2864 , n2886 , n2888 , n2912 , 
n3038 , n3092 , n3120 , n3209 , n3321 , n3340 , n3365 , n3384 , n3411 , n3444 , 
n3452 , n3465 , n3481 , n3506 , n3510 , n3536 , n3615 , n3631 , n3690 , n3742 , 
n3774 , n3800 , n3805 , n3806 , n3898 );
    input n4 , n44 , n56 , n66 , n88 , n181 , n185 , n196 , n220 , 
n274 , n308 , n335 , n422 , n493 , n504 , n523 , n530 , n642 , n670 , 
n705 , n722 , n770 , n772 , n794 , n824 , n829 , n835 , n866 , n873 , 
n891 , n927 , n928 , n935 , n940 , n944 , n955 , n1066 , n1103 , n1140 , 
n1156 , n1202 , n1234 , n1240 , n1273 , n1280 , n1361 , n1367 , n1387 , n1404 , 
n1432 , n1507 , n1521 , n1541 , n1638 , n1646 , n1761 , n1775 , n1793 , n1808 , 
n1820 , n1861 , n1874 , n1938 , n2031 , n2050 , n2055 , n2073 , n2110 , n2112 , 
n2165 , n2195 , n2223 , n2252 , n2258 , n2313 , n2324 , n2371 , n2402 , n2463 , 
n2514 , n2523 , n2567 , n2572 , n2640 , n2664 , n2724 , n2727 , n2744 , n2757 , 
n2760 , n2806 , n2830 , n2886 , n2888 , n2912 , n3038 , n3092 , n3120 , n3321 , 
n3340 , n3365 , n3384 , n3411 , n3444 , n3465 , n3481 , n3506 , n3510 , n3536 , 
n3615 , n3631 , n3690 , n3742 , n3774 , n3800 , n3805 , n3898 ;
    output n37 , n84 , n132 , n850 , n872 , n1157 , n1229 , n1398 , n1540 , 
n1889 , n2385 , n2490 , n2622 , n2864 , n3209 , n3452 , n3806 ;
    wire n0 , n1 , n2 , n3 , n5 , n6 , n7 , n8 , n9 , 
n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
n30 , n31 , n32 , n33 , n34 , n35 , n36 , n38 , n39 , n40 , 
n41 , n42 , n43 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , 
n52 , n53 , n54 , n55 , n57 , n58 , n59 , n60 , n61 , n62 , 
n63 , n64 , n65 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , 
n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , 
n85 , n86 , n87 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , 
n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , 
n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , 
n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , 
n126 , n127 , n128 , n129 , n130 , n131 , n133 , n134 , n135 , n136 , 
n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , 
n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , 
n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
n177 , n178 , n179 , n180 , n182 , n183 , n184 , n186 , n187 , n188 , 
n189 , n190 , n191 , n192 , n193 , n194 , n195 , n197 , n198 , n199 , 
n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
n271 , n272 , n273 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , 
n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , 
n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , 
n302 , n303 , n304 , n305 , n306 , n307 , n309 , n310 , n311 , n312 , 
n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , 
n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , 
n333 , n334 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , 
n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , 
n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , 
n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , 
n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , 
n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , 
n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , 
n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , 
n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n423 , n424 , 
n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , 
n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , 
n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , 
n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , 
n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , 
n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , 
n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n494 , n495 , 
n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n505 , n506 , 
n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , 
n517 , n518 , n519 , n520 , n521 , n522 , n524 , n525 , n526 , n527 , 
n528 , n529 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , 
n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , 
n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , 
n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , 
n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , 
n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , 
n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , 
n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , 
n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , 
n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , 
n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , 
n639 , n640 , n641 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , 
n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , 
n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , 
n701 , n702 , n703 , n704 , n706 , n707 , n708 , n709 , n710 , n711 , 
n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , 
n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , 
n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , 
n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , 
n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , 
n763 , n764 , n765 , n766 , n767 , n768 , n769 , n771 , n773 , n774 , 
n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , 
n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n795 , 
n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , 
n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , 
n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n825 , n826 , 
n827 , n828 , n830 , n831 , n832 , n833 , n834 , n836 , n837 , n838 , 
n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , 
n849 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
n860 , n861 , n862 , n863 , n864 , n865 , n867 , n868 , n869 , n870 , 
n871 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , 
n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n892 , n893 , 
n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , 
n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , 
n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , 
n924 , n925 , n926 , n929 , n930 , n931 , n932 , n933 , n934 , n936 , 
n937 , n938 , n939 , n941 , n942 , n943 , n945 , n946 , n947 , n948 , 
n949 , n950 , n951 , n952 , n953 , n954 , n956 , n957 , n958 , n959 , 
n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1067 , n1068 , n1069 , n1070 , 
n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , 
n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , 
n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , 
n1101 , n1102 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , 
n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , 
n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , 
n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1141 , n1142 , 
n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , 
n1153 , n1154 , n1155 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , 
n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , 
n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , 
n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , 
n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1203 , n1204 , n1205 , 
n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , 
n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , 
n1226 , n1227 , n1228 , n1230 , n1231 , n1232 , n1233 , n1235 , n1236 , n1237 , 
n1238 , n1239 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , 
n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , 
n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , 
n1269 , n1270 , n1271 , n1272 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , 
n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , 
n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , 
n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , 
n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , 
n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , 
n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , 
n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , 
n1362 , n1363 , n1364 , n1365 , n1366 , n1368 , n1369 , n1370 , n1371 , n1372 , 
n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , 
n1383 , n1384 , n1385 , n1386 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , 
n1394 , n1395 , n1396 , n1397 , n1399 , n1400 , n1401 , n1402 , n1403 , n1405 , 
n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , 
n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , 
n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1433 , n1434 , n1435 , n1436 , 
n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , 
n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , 
n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , 
n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , 
n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , 
n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , 
n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , 
n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , 
n1518 , n1519 , n1520 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , 
n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , 
n1539 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , 
n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , 
n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , 
n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , 
n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , 
n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , 
n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , 
n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , 
n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , 
n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1639 , n1640 , n1641 , 
n1642 , n1643 , n1644 , n1645 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , 
n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , 
n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , 
n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , 
n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , 
n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , 
n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , 
n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , 
n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , 
n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , 
n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , 
n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1762 , n1763 , 
n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , 
n1774 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , 
n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1794 , n1795 , 
n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , 
n1806 , n1807 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , 
n1817 , n1818 , n1819 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , 
n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , 
n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , 
n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , 
n1858 , n1859 , n1860 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , 
n1869 , n1870 , n1871 , n1872 , n1873 , n1875 , n1876 , n1877 , n1878 , n1879 , 
n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1890 , 
n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , 
n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , 
n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , 
n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , 
n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1939 , n1940 , n1941 , 
n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , 
n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , 
n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , 
n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , 
n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , 
n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , 
n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , 
n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , 
n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2032 , 
n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , 
n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2051 , n2052 , n2053 , 
n2054 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , 
n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2074 , n2075 , 
n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , 
n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , 
n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , 
n2106 , n2107 , n2108 , n2109 , n2111 , n2113 , n2114 , n2115 , n2116 , n2117 , 
n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , 
n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , 
n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , 
n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , 
n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2166 , n2167 , n2168 , 
n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , 
n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , 
n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2196 , n2197 , n2198 , n2199 , 
n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
n2220 , n2221 , n2222 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , 
n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , 
n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , 
n2251 , n2253 , n2254 , n2255 , n2256 , n2257 , n2259 , n2260 , n2261 , n2262 , 
n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , 
n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , 
n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , 
n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , 
n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , 
n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , 
n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , 
n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , 
n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , 
n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , 
n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2372 , n2373 , n2374 , n2375 , 
n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2386 , 
n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , 
n2397 , n2398 , n2399 , n2400 , n2401 , n2403 , n2404 , n2405 , n2406 , n2407 , 
n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , 
n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , 
n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , 
n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , 
n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , 
n2458 , n2459 , n2460 , n2461 , n2462 , n2464 , n2465 , n2466 , n2467 , n2468 , 
n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , 
n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , 
n2489 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
n2510 , n2511 , n2512 , n2513 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , 
n2521 , n2522 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , 
n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , 
n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , 
n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , 
n2562 , n2563 , n2564 , n2565 , n2566 , n2568 , n2569 , n2570 , n2571 , n2573 , 
n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , 
n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , 
n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , 
n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , 
n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2623 , n2624 , 
n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , 
n2635 , n2636 , n2637 , n2638 , n2639 , n2641 , n2642 , n2643 , n2644 , n2645 , 
n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , 
n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2665 , n2666 , 
n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , 
n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , 
n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , 
n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , 
n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , 
n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2725 , n2726 , n2728 , 
n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , 
n2739 , n2740 , n2741 , n2742 , n2743 , n2745 , n2746 , n2747 , n2748 , n2749 , 
n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2758 , n2759 , n2761 , 
n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , 
n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , 
n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , 
n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , 
n2802 , n2803 , n2804 , n2805 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , 
n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , 
n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2831 , n2832 , n2833 , 
n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , 
n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , 
n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , 
n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , 
n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , 
n2885 , n2887 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , 
n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , 
n2907 , n2908 , n2909 , n2910 , n2911 , n2913 , n2914 , n2915 , n2916 , n2917 , 
n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , 
n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , 
n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , 
n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , 
n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , 
n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , 
n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , 
n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , 
n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , 
n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , 
n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , 
n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , 
n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , 
n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , 
n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , 
n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , 
n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , 
n3089 , n3090 , n3091 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , 
n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , 
n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , 
n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , 
n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , 
n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , 
n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3210 , n3211 , 
n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , 
n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , 
n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , 
n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , 
n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , 
n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , 
n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , 
n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , 
n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , 
n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , 
n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3322 , 
n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , 
n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3341 , n3342 , n3343 , 
n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , 
n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , 
n3364 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , 
n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3385 , 
n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , 
n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , 
n3406 , n3407 , n3408 , n3409 , n3410 , n3412 , n3413 , n3414 , n3415 , n3416 , 
n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , 
n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , 
n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3445 , n3446 , n3447 , 
n3448 , n3449 , n3450 , n3451 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , 
n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3466 , n3467 , n3468 , n3469 , 
n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
n3480 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
n3501 , n3502 , n3503 , n3504 , n3505 , n3507 , n3508 , n3509 , n3511 , n3512 , 
n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , 
n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , 
n3533 , n3534 , n3535 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , 
n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , 
n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , 
n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , 
n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , 
n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , 
n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , 
n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , 
n3614 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , 
n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3632 , n3633 , n3634 , n3635 , 
n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , 
n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , 
n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , 
n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , 
n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , 
n3686 , n3687 , n3688 , n3689 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , 
n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , 
n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , 
n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , 
n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , 
n3737 , n3738 , n3739 , n3740 , n3741 , n3743 , n3744 , n3745 , n3746 , n3747 , 
n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , 
n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , 
n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3775 , n3776 , n3777 , n3778 , 
n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , 
n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , 
n3799 , n3801 , n3802 , n3803 , n3804 , n3807 , n3808 , n3809 , n3810 , n3811 , 
n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , 
n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , 
n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , 
n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , 
n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , 
n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , 
n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , 
n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , 
n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3899 , n3900 , n3901 , n3902 ;
    xnor g0 ( n381 , n2720 , n2736 );
    not g1 ( n1688 , n1656 );
    xnor g2 ( n1087 , n3601 , n3652 );
    and g3 ( n780 , n2333 , n2097 );
    not g4 ( n1584 , n2822 );
    xnor g5 ( n1575 , n2950 , n2954 );
    xnor g6 ( n3618 , n1271 , n3801 );
    and g7 ( n584 , n1833 , n3231 );
    not g8 ( n2951 , n2324 );
    and g9 ( n1679 , n2686 , n677 );
    or g10 ( n3699 , n1733 , n427 );
    xnor g11 ( n3825 , n787 , n2306 );
    xnor g12 ( n1490 , n2341 , n1218 );
    xnor g13 ( n3222 , n1907 , n502 );
    nor g14 ( n3248 , n487 , n277 );
    and g15 ( n120 , n1766 , n2156 );
    not g16 ( n2194 , n3742 );
    or g17 ( n2674 , n3839 , n1227 );
    and g18 ( n96 , n732 , n1027 );
    not g19 ( n655 , n789 );
    nor g20 ( n2020 , n853 , n1231 );
    xnor g21 ( n2768 , n275 , n1556 );
    nor g22 ( n129 , n3405 , n1755 );
    or g23 ( n724 , n3058 , n3210 );
    xnor g24 ( n3532 , n223 , n2131 );
    not g25 ( n2561 , n1735 );
    xnor g26 ( n2238 , n2083 , n1736 );
    or g27 ( n571 , n1678 , n1660 );
    and g28 ( n1560 , n877 , n1390 );
    or g29 ( n3766 , n310 , n3741 );
    xor g30 ( n77 , n1993 , n1759 );
    or g31 ( n807 , n2620 , n3394 );
    not g32 ( n3785 , n3649 );
    xnor g33 ( n1848 , n2986 , n966 );
    or g34 ( n3663 , n365 , n593 );
    or g35 ( n1582 , n2662 , n210 );
    and g36 ( n1311 , n730 , n331 );
    or g37 ( n1858 , n290 , n1987 );
    xnor g38 ( n656 , n1605 , n2665 );
    not g39 ( n1804 , n2209 );
    xnor g40 ( n3042 , n1095 , n3879 );
    and g41 ( n1401 , n1829 , n3237 );
    and g42 ( n2146 , n1271 , n2154 );
    xnor g43 ( n2088 , n49 , n1680 );
    not g44 ( n2124 , n2804 );
    xnor g45 ( n2288 , n3034 , n1618 );
    xnor g46 ( n631 , n540 , n1911 );
    or g47 ( n1226 , n431 , n2331 );
    or g48 ( n3417 , n3130 , n476 );
    or g49 ( n2774 , n605 , n1758 );
    or g50 ( n3706 , n2392 , n2790 );
    xnor g51 ( n684 , n1546 , n1977 );
    or g52 ( n1830 , n3324 , n3072 );
    xnor g53 ( n178 , n3691 , n2068 );
    and g54 ( n1873 , n3262 , n2962 );
    not g55 ( n2682 , n2567 );
    xnor g56 ( n1412 , n3363 , n2634 );
    xnor g57 ( n198 , n5 , n2443 );
    not g58 ( n754 , n3742 );
    xnor g59 ( n3477 , n3757 , n293 );
    xnor g60 ( n1670 , n2846 , n2057 );
    or g61 ( n1591 , n3622 , n2935 );
    not g62 ( n128 , n3360 );
    xnor g63 ( n288 , n1686 , n904 );
    and g64 ( n1846 , n1614 , n1778 );
    and g65 ( n1247 , n69 , n968 );
    not g66 ( n538 , n211 );
    and g67 ( n811 , n3608 , n1635 );
    not g68 ( n2859 , n3365 );
    or g69 ( n2186 , n1994 , n2922 );
    or g70 ( n820 , n1620 , n2243 );
    and g71 ( n1469 , n1543 , n2518 );
    or g72 ( n1120 , n1794 , n1431 );
    and g73 ( n1117 , n956 , n3216 );
    not g74 ( n1053 , n422 );
    not g75 ( n285 , n185 );
    or g76 ( n3653 , n1808 , n1434 );
    xnor g77 ( n3083 , n2673 , n2033 );
    or g78 ( n3639 , n1776 , n3483 );
    xnor g79 ( n2893 , n1100 , n3044 );
    and g80 ( n3421 , n2722 , n640 );
    and g81 ( n252 , n57 , n2699 );
    not g82 ( n3460 , n422 );
    or g83 ( n171 , n880 , n830 );
    and g84 ( n1397 , n2566 , n957 );
    xnor g85 ( n1305 , n2217 , n526 );
    and g86 ( n462 , n260 , n2389 );
    xnor g87 ( n1523 , n1537 , n2970 );
    and g88 ( n1918 , n3289 , n91 );
    xnor g89 ( n517 , n901 , n698 );
    xnor g90 ( n2046 , n2656 , n1305 );
    not g91 ( n2284 , n3340 );
    or g92 ( n2375 , n355 , n1821 );
    or g93 ( n1709 , n2412 , n3071 );
    or g94 ( n595 , n2081 , n1661 );
    and g95 ( n2015 , n3733 , n3211 );
    xnor g96 ( n52 , n1633 , n2214 );
    not g97 ( n2594 , n2912 );
    xnor g98 ( n3580 , n3487 , n2290 );
    xnor g99 ( n35 , n1423 , n1353 );
    and g100 ( n1878 , n327 , n980 );
    xnor g101 ( n23 , n3215 , n3116 );
    or g102 ( n1336 , n211 , n256 );
    or g103 ( n907 , n3815 , n3168 );
    not g104 ( n3584 , n2402 );
    xnor g105 ( n3635 , n2142 , n1663 );
    or g106 ( n1416 , n3565 , n1358 );
    not g107 ( n1381 , n2231 );
    and g108 ( n1452 , n750 , n3713 );
    xnor g109 ( n1781 , n2908 , n3016 );
    not g110 ( n1064 , n935 );
    or g111 ( n326 , n511 , n1993 );
    xnor g112 ( n2896 , n2462 , n2414 );
    xnor g113 ( n2866 , n2491 , n1586 );
    and g114 ( n1433 , n2144 , n209 );
    and g115 ( n1097 , n3122 , n2992 );
    or g116 ( n1827 , n3612 , n621 );
    and g117 ( n3673 , n2730 , n3443 );
    or g118 ( n3099 , n3051 , n2468 );
    not g119 ( n1505 , n3038 );
    or g120 ( n2019 , n2278 , n625 );
    xnor g121 ( n3106 , n3751 , n1159 );
    not g122 ( n727 , n3359 );
    or g123 ( n3077 , n2302 , n3157 );
    not g124 ( n2602 , n3383 );
    or g125 ( n957 , n3002 , n2965 );
    xnor g126 ( n399 , n3079 , n2916 );
    not g127 ( n72 , n2725 );
    and g128 ( n1050 , n994 , n3517 );
    or g129 ( n690 , n24 , n3083 );
    or g130 ( n3496 , n2959 , n3404 );
    xnor g131 ( n2399 , n1394 , n2155 );
    and g132 ( n404 , n1995 , n3661 );
    not g133 ( n997 , n3092 );
    xnor g134 ( n1633 , n1921 , n3846 );
    xnor g135 ( n3276 , n8 , n3357 );
    and g136 ( n962 , n608 , n2604 );
    or g137 ( n3789 , n2957 , n473 );
    and g138 ( n3274 , n827 , n1920 );
    or g139 ( n346 , n2789 , n627 );
    not g140 ( n187 , n1361 );
    xnor g141 ( n3193 , n648 , n1433 );
    not g142 ( n3348 , n3371 );
    and g143 ( n742 , n583 , n1238 );
    not g144 ( n3183 , n2450 );
    xnor g145 ( n208 , n2108 , n3583 );
    or g146 ( n1347 , n1734 , n3475 );
    xnor g147 ( n2236 , n2170 , n1701 );
    or g148 ( n739 , n3855 , n2949 );
    not g149 ( n3140 , n2982 );
    or g150 ( n2645 , n1610 , n2439 );
    or g151 ( n2147 , n3431 , n2533 );
    or g152 ( n887 , n2425 , n2492 );
    xnor g153 ( n1434 , n2216 , n2692 );
    and g154 ( n3252 , n3364 , n2047 );
    not g155 ( n2117 , n1682 );
    and g156 ( n3109 , n3407 , n1445 );
    not g157 ( n3887 , n873 );
    xnor g158 ( n3764 , n1564 , n1598 );
    xnor g159 ( n3683 , n2321 , n448 );
    not g160 ( n1489 , n2073 );
    xnor g161 ( n236 , n2166 , n2698 );
    or g162 ( n157 , n328 , n168 );
    and g163 ( n1268 , n2761 , n331 );
    and g164 ( n402 , n560 , n1786 );
    not g165 ( n2666 , n3724 );
    not g166 ( n2379 , n2514 );
    or g167 ( n3544 , n2005 , n1413 );
    or g168 ( n426 , n2758 , n1073 );
    not g169 ( n2234 , n1030 );
    or g170 ( n1559 , n1538 , n646 );
    and g171 ( n3311 , n943 , n374 );
    xnor g172 ( n1169 , n3326 , n3410 );
    not g173 ( n660 , n642 );
    or g174 ( n2801 , n235 , n2511 );
    not g175 ( n1191 , n2993 );
    xnor g176 ( n67 , n2871 , n2259 );
    or g177 ( n3094 , n2605 , n534 );
    nor g178 ( n3875 , n1459 , n2899 );
    not g179 ( n2938 , n2593 );
    or g180 ( n1669 , n1113 , n1626 );
    xnor g181 ( n64 , n3179 , n206 );
    or g182 ( n2298 , n2738 , n3367 );
    xnor g183 ( n369 , n3495 , n67 );
    not g184 ( n1399 , n3084 );
    xnor g185 ( n2207 , n605 , n1515 );
    not g186 ( n2537 , n335 );
    or g187 ( n1137 , n3835 , n620 );
    or g188 ( n3097 , n240 , n2092 );
    and g189 ( n2057 , n3441 , n832 );
    or g190 ( n1328 , n648 , n1433 );
    xnor g191 ( n119 , n3544 , n2255 );
    not g192 ( n2386 , n1804 );
    and g193 ( n1033 , n765 , n3902 );
    or g194 ( n2576 , n613 , n851 );
    not g195 ( n3817 , n1320 );
    or g196 ( n3533 , n469 , n2498 );
    and g197 ( n1001 , n933 , n2337 );
    or g198 ( n3022 , n2227 , n419 );
    and g199 ( n1357 , n1130 , n1753 );
    xnor g200 ( n3442 , n1445 , n452 );
    or g201 ( n3524 , n2477 , n1872 );
    xnor g202 ( n874 , n168 , n2980 );
    or g203 ( n1583 , n1708 , n3546 );
    or g204 ( n498 , n2027 , n2505 );
    or g205 ( n3852 , n2194 , n881 );
    or g206 ( n2028 , n2644 , n3732 );
    and g207 ( n3879 , n1908 , n139 );
    xnor g208 ( n3320 , n1105 , n3207 );
    xnor g209 ( n1828 , n3160 , n1651 );
    xnor g210 ( n3459 , n3178 , n2565 );
    or g211 ( n3391 , n1937 , n2365 );
    or g212 ( n2972 , n1461 , n3700 );
    not g213 ( n290 , n3742 );
    or g214 ( n1887 , n895 , n1871 );
    xnor g215 ( n857 , n917 , n951 );
    not g216 ( n2099 , n1938 );
    nor g217 ( n749 , n2262 , n2428 );
    xnor g218 ( n886 , n2999 , n1409 );
    nor g219 ( n1073 , n723 , n2369 );
    not g220 ( n2250 , n927 );
    or g221 ( n609 , n3288 , n920 );
    or g222 ( n2656 , n2894 , n2496 );
    or g223 ( n3069 , n430 , n2611 );
    not g224 ( n2706 , n3743 );
    and g225 ( n2804 , n77 , n2481 );
    and g226 ( n2828 , n2826 , n481 );
    or g227 ( n2981 , n963 , n2569 );
    and g228 ( n2149 , n1758 , n605 );
    or g229 ( n3237 , n1505 , n2592 );
    xnor g230 ( n3883 , n1331 , n3832 );
    xor g231 ( n3811 , n330 , n165 );
    xnor g232 ( n3822 , n1990 , n2978 );
    xnor g233 ( n580 , n2879 , n3689 );
    not g234 ( n1113 , n1432 );
    xnor g235 ( n3305 , n117 , n2890 );
    nor g236 ( n1046 , n1291 , n3891 );
    and g237 ( n1773 , n2083 , n735 );
    not g238 ( n926 , n1892 );
    not g239 ( n130 , n3120 );
    and g240 ( n3263 , n3056 , n869 );
    xnor g241 ( n3669 , n3889 , n2433 );
    nor g242 ( n2227 , n1320 , n2840 );
    not g243 ( n2012 , n1541 );
    or g244 ( n3113 , n643 , n3647 );
    and g245 ( n915 , n1091 , n99 );
    and g246 ( n1661 , n724 , n557 );
    xnor g247 ( n1147 , n3076 , n1612 );
    nor g248 ( n397 , n78 , n3156 );
    xnor g249 ( n1470 , n1104 , n1905 );
    or g250 ( n2923 , n1992 , n1868 );
    or g251 ( n3179 , n736 , n797 );
    or g252 ( n3812 , n808 , n1490 );
    and g253 ( n1948 , n3663 , n1923 );
    or g254 ( n3119 , n2448 , n1050 );
    and g255 ( n624 , n891 , n2888 );
    not g256 ( n2611 , n1761 );
    xor g257 ( n1337 , n3134 , n268 );
    and g258 ( n2013 , n2915 , n1415 );
    or g259 ( n3757 , n2808 , n2167 );
    and g260 ( n1192 , n1703 , n1009 );
    or g261 ( n3870 , n3697 , n896 );
    or g262 ( n1710 , n2660 , n1619 );
    not g263 ( n2548 , n2724 );
    or g264 ( n1730 , n1059 , n1647 );
    not g265 ( n2887 , n1938 );
    or g266 ( n505 , n919 , n1976 );
    not g267 ( n2287 , n927 );
    or g268 ( n1925 , n1884 , n2887 );
    or g269 ( n2254 , n1482 , n1069 );
    xnor g270 ( n1153 , n427 , n2456 );
    and g271 ( n3210 , n2228 , n3591 );
    or g272 ( n1460 , n1348 , n3555 );
    and g273 ( n930 , n703 , n3264 );
    and g274 ( n261 , n2892 , n3715 );
    or g275 ( n2665 , n1076 , n3164 );
    or g276 ( n3225 , n2677 , n1413 );
    or g277 ( n3287 , n1547 , n3049 );
    or g278 ( n3306 , n2923 , n2836 );
    and g279 ( n2181 , n3430 , n2740 );
    xnor g280 ( n3617 , n3161 , n2104 );
    or g281 ( n1519 , n1011 , n1868 );
    xnor g282 ( n2135 , n2380 , n755 );
    not g283 ( n1610 , n1874 );
    or g284 ( n3651 , n1744 , n1605 );
    xnor g285 ( n2961 , n2436 , n23 );
    not g286 ( n2010 , n3327 );
    or g287 ( n2821 , n3556 , n154 );
    not g288 ( n1249 , n39 );
    and g289 ( n587 , n1840 , n2735 );
    or g290 ( n2251 , n49 , n604 );
    or g291 ( n1966 , n581 , n2679 );
    or g292 ( n2623 , n3573 , n471 );
    and g293 ( n2822 , n2878 , n1444 );
    and g294 ( n3424 , n2001 , n2209 );
    or g295 ( n1644 , n0 , n1333 );
    xor g296 ( n1480 , n1920 , n12 );
    or g297 ( n2208 , n819 , n281 );
    or g298 ( n702 , n2858 , n2441 );
    or g299 ( n650 , n680 , n166 );
    and g300 ( n244 , n3339 , n1068 );
    xor g301 ( n2306 , n3027 , n1138 );
    not g302 ( n1262 , n722 );
    or g303 ( n3570 , n1462 , n2447 );
    xnor g304 ( n1832 , n2018 , n2669 );
    nor g305 ( n542 , n3160 , n1705 );
    and g306 ( n2750 , n1235 , n3586 );
    and g307 ( n1719 , n2514 , n1367 );
    and g308 ( n2473 , n2166 , n3011 );
    or g309 ( n1851 , n855 , n1292 );
    and g310 ( n3529 , n58 , n1901 );
    or g311 ( n267 , n975 , n500 );
    nor g312 ( n3447 , n2010 , n1331 );
    or g313 ( n876 , n1167 , n1514 );
    or g314 ( n2404 , n282 , n630 );
    xnor g315 ( n2275 , n503 , n64 );
    or g316 ( n170 , n3882 , n392 );
    xnor g317 ( n1196 , n2048 , n3462 );
    or g318 ( n1562 , n3764 , n3013 );
    and g319 ( n936 , n752 , n1423 );
    xnor g320 ( n3360 , n152 , n3693 );
    xnor g321 ( n2732 , n1930 , n3280 );
    xnor g322 ( n3373 , n3387 , n789 );
    and g323 ( n1812 , n1755 , n3405 );
    not g324 ( n1516 , n3387 );
    not g325 ( n1857 , n2468 );
    xor g326 ( n3499 , n1846 , n2996 );
    xnor g327 ( n1634 , n2961 , n2158 );
    and g328 ( n2038 , n1597 , n1461 );
    not g329 ( n388 , n1209 );
    nor g330 ( n3239 , n381 , n911 );
    xnor g331 ( n312 , n247 , n2937 );
    and g332 ( n2162 , n3187 , n2406 );
    and g333 ( n1293 , n3252 , n86 );
    or g334 ( n2712 , n1190 , n1627 );
    nor g335 ( n3730 , n822 , n2673 );
    xnor g336 ( n1465 , n2936 , n1254 );
    or g337 ( n665 , n2291 , n3271 );
    and g338 ( n864 , n3838 , n2298 );
    and g339 ( n2447 , n757 , n3079 );
    or g340 ( n3535 , n1391 , n3558 );
    xnor g341 ( n1172 , n623 , n2785 );
    or g342 ( n512 , n2052 , n3597 );
    xnor g343 ( n1574 , n2813 , n2897 );
    and g344 ( n2257 , n1350 , n1770 );
    xnor g345 ( n2440 , n288 , n885 );
    not g346 ( n3358 , n2889 );
    or g347 ( n3376 , n2473 , n2701 );
    or g348 ( n2044 , n198 , n2323 );
    not g349 ( n2705 , n2932 );
    or g350 ( n2532 , n2477 , n2809 );
    and g351 ( n1228 , n2715 , n611 );
    or g352 ( n2635 , n1533 , n1977 );
    and g353 ( n2204 , n3391 , n3676 );
    and g354 ( n1612 , n3818 , n2802 );
    xnor g355 ( n3693 , n1006 , n3271 );
    xnor g356 ( n1897 , n915 , n2952 );
    or g357 ( n202 , n3879 , n3296 );
    and g358 ( n1951 , n695 , n3825 );
    and g359 ( n2416 , n95 , n1328 );
    or g360 ( n2077 , n3896 , n1312 );
    not g361 ( n1482 , n1634 );
    or g362 ( n1021 , n2835 , n51 );
    or g363 ( n3445 , n1844 , n2526 );
    xnor g364 ( n1841 , n97 , n421 );
    or g365 ( n2542 , n1897 , n3420 );
    not g366 ( n2413 , n2258 );
    or g367 ( n1629 , n2831 , n1694 );
    and g368 ( n3579 , n3197 , n2119 );
    nor g369 ( n2369 , n1311 , n438 );
    or g370 ( n2226 , n3703 , n149 );
    and g371 ( n911 , n3744 , n595 );
    or g372 ( n3431 , n599 , n3830 );
    and g373 ( n3605 , n3159 , n2395 );
    not g374 ( n3301 , n1604 );
    not g375 ( n1694 , n1638 );
    and g376 ( n706 , n2767 , n1745 );
    or g377 ( n1984 , n1045 , n1135 );
    or g378 ( n2187 , n2436 , n1602 );
    or g379 ( n3327 , n3465 , n586 );
    or g380 ( n3241 , n1028 , n2164 );
    not g381 ( n296 , n2223 );
    or g382 ( n975 , n1083 , n947 );
    or g383 ( n3361 , n2491 , n1586 );
    and g384 ( n1916 , n2908 , n637 );
    and g385 ( n1317 , n1361 , n1234 );
    not g386 ( n320 , n1273 );
    nor g387 ( n1295 , n374 , n943 );
    xnor g388 ( n3219 , n3139 , n2583 );
    nor g389 ( n2281 , n2224 , n3342 );
    not g390 ( n3900 , n1446 );
    xnor g391 ( n1860 , n3872 , n1603 );
    xor g392 ( n1797 , n7 , n1182 );
    xnor g393 ( n3833 , n3304 , n444 );
    or g394 ( n3389 , n1031 , n1542 );
    or g395 ( n1561 , n1863 , n1394 );
    or g396 ( n10 , n1697 , n3266 );
    not g397 ( n3609 , n2486 );
    nor g398 ( n682 , n1341 , n2403 );
    and g399 ( n1200 , n424 , n2197 );
    or g400 ( n34 , n3479 , n1228 );
    or g401 ( n1814 , n563 , n2696 );
    and g402 ( n3415 , n1885 , n786 );
    xnor g403 ( n1603 , n1368 , n3634 );
    not g404 ( n1689 , n2624 );
    not g405 ( n3472 , n1204 );
    not g406 ( n3103 , n2532 );
    and g407 ( n2526 , n3496 , n1037 );
    or g408 ( n1168 , n6 , n3755 );
    not g409 ( n2512 , n3795 );
    not g410 ( n2973 , n824 );
    xnor g411 ( n2963 , n3166 , n2989 );
    xnor g412 ( n978 , n3176 , n684 );
    and g413 ( n3125 , n2820 , n2307 );
    and g414 ( n33 , n3124 , n3047 );
    or g415 ( n1555 , n2280 , n2474 );
    and g416 ( n1108 , n484 , n507 );
    xnor g417 ( n1763 , n2283 , n3565 );
    nor g418 ( n3439 , n12 , n1058 );
    and g419 ( n1015 , n756 , n2545 );
    and g420 ( n3634 , n2285 , n3261 );
    nor g421 ( n1904 , n3421 , n3308 );
    or g422 ( n1500 , n843 , n2880 );
    xnor g423 ( n2698 , n3011 , n2701 );
    or g424 ( n478 , n2906 , n2420 );
    or g425 ( n375 , n3252 , n86 );
    and g426 ( n1985 , n812 , n3406 );
    not g427 ( n3597 , n1234 );
    not g428 ( n2588 , n3690 );
    and g429 ( n1942 , n2210 , n3107 );
    not g430 ( n696 , n3408 );
    or g431 ( n1659 , n147 , n997 );
    and g432 ( n2059 , n1226 , n400 );
    not g433 ( n2998 , n3805 );
    not g434 ( n3104 , n705 );
    xnor g435 ( n951 , n3599 , n472 );
    or g436 ( n1671 , n2886 , n1558 );
    xnor g437 ( n2612 , n821 , n1725 );
    and g438 ( n3736 , n63 , n2960 );
    or g439 ( n1778 , n3327 , n1952 );
    or g440 ( n1508 , n147 , n2184 );
    and g441 ( n1477 , n1562 , n2451 );
    and g442 ( n3799 , n1426 , n3195 );
    and g443 ( n3323 , n876 , n1021 );
    xnor g444 ( n103 , n967 , n597 );
    not g445 ( n1389 , n1945 );
    nor g446 ( n2171 , n3547 , n2237 );
    nor g447 ( n2873 , n2112 , n1017 );
    not g448 ( n1034 , n2123 );
    and g449 ( n2871 , n3330 , n1717 );
    xnor g450 ( n279 , n3329 , n517 );
    and g451 ( n558 , n694 , n1859 );
    xnor g452 ( n28 , n1755 , n3669 );
    not g453 ( n590 , n2523 );
    xnor g454 ( n3657 , n1508 , n2222 );
    not g455 ( n3593 , n1305 );
    not g456 ( n2016 , n1202 );
    or g457 ( n2741 , n649 , n1108 );
    not g458 ( n1950 , n3686 );
    xnor g459 ( n2805 , n494 , n874 );
    xnor g460 ( n3185 , n419 , n354 );
    and g461 ( n1183 , n1740 , n1441 );
    or g462 ( n2102 , n321 , n1284 );
    and g463 ( n633 , n1721 , n1310 );
    not g464 ( n848 , n928 );
    or g465 ( n31 , n2233 , n3446 );
    not g466 ( n207 , n66 );
    not g467 ( n3074 , n196 );
    or g468 ( n2415 , n3127 , n1899 );
    and g469 ( n1212 , n133 , n1047 );
    and g470 ( n2133 , n815 , n941 );
    xnor g471 ( n663 , n1272 , n3747 );
    and g472 ( n2175 , n2629 , n26 );
    xnor g473 ( n568 , n3675 , n1285 );
    and g474 ( n1285 , n450 , n3854 );
    or g475 ( n3692 , n3301 , n3112 );
    not g476 ( n1868 , n3384 );
    xnor g477 ( n2520 , n426 , n3224 );
    and g478 ( n1390 , n378 , n2951 );
    xnor g479 ( n2433 , n3899 , n304 );
    and g480 ( n3032 , n1043 , n331 );
    and g481 ( n3563 , n2325 , n3295 );
    xnor g482 ( n1643 , n3158 , n1236 );
    or g483 ( n411 , n3725 , n3562 );
    or g484 ( n91 , n1720 , n411 );
    or g485 ( n846 , n2128 , n3563 );
    nor g486 ( n1590 , n878 , n1792 );
    and g487 ( n1055 , n1781 , n3675 );
    not g488 ( n3509 , n829 );
    and g489 ( n3063 , n2657 , n21 );
    xor g490 ( n2722 , n2015 , n2489 );
    or g491 ( n1931 , n3108 , n3850 );
    xnor g492 ( n440 , n2209 , n1004 );
    not g493 ( n2585 , n3465 );
    or g494 ( n3860 , n390 , n1172 );
    or g495 ( n3335 , n752 , n1423 );
    or g496 ( n3436 , n1629 , n2818 );
    xnor g497 ( n3007 , n1606 , n1658 );
    xnor g498 ( n1738 , n461 , n2070 );
    xnor g499 ( n3418 , n3784 , n760 );
    or g500 ( n3413 , n3 , n777 );
    and g501 ( n3619 , n2414 , n2462 );
    not g502 ( n3694 , n2643 );
    nor g503 ( n658 , n66 , n836 );
    xnor g504 ( n1221 , n3431 , n2704 );
    not g505 ( n764 , n3898 );
    not g506 ( n3561 , n3399 );
    or g507 ( n1747 , n2886 , n3580 );
    and g508 ( n1086 , n3334 , n3077 );
    or g509 ( n2001 , n1992 , n1262 );
    xnor g510 ( n651 , n411 , n3253 );
    or g511 ( n2667 , n124 , n2413 );
    or g512 ( n2837 , n2263 , n180 );
    or g513 ( n110 , n1127 , n3732 );
    and g514 ( n1739 , n3125 , n623 );
    or g515 ( n3201 , n3788 , n1552 );
    and g516 ( n653 , n1038 , n2763 );
    or g517 ( n2659 , n356 , n368 );
    or g518 ( n1571 , n609 , n3023 );
    and g519 ( n1734 , n787 , n3027 );
    and g520 ( n2689 , n1352 , n833 );
    and g521 ( n3451 , n2688 , n3484 );
    xnor g522 ( n1766 , n2781 , n2729 );
    or g523 ( n2309 , n2644 , n3830 );
    xnor g524 ( n1903 , n2224 , n3152 );
    or g525 ( n1599 , n3509 , n3460 );
    not g526 ( n2022 , n3139 );
    xnor g527 ( n3105 , n3056 , n3349 );
    and g528 ( n3207 , n1267 , n3523 );
    not g529 ( n1413 , n2463 );
    nor g530 ( n2037 , n773 , n92 );
    or g531 ( n2418 , n2152 , n1141 );
    or g532 ( n2011 , n1160 , n1870 );
    or g533 ( n3756 , n2974 , n1284 );
    nor g534 ( n1017 , n2292 , n3239 );
    not g535 ( n621 , n3615 );
    and g536 ( n2605 , n3053 , n2208 );
    not g537 ( n329 , n1361 );
    xnor g538 ( n1217 , n857 , n2059 );
    or g539 ( n3521 , n3643 , n1293 );
    nor g540 ( n1955 , n1030 , n3372 );
    nor g541 ( n638 , n3015 , n1309 );
    or g542 ( n2582 , n413 , n3169 );
    not g543 ( n1446 , n1463 );
    and g544 ( n3072 , n1032 , n1253 );
    and g545 ( n1069 , n1400 , n578 );
    xnor g546 ( n3743 , n1983 , n2943 );
    not g547 ( n2809 , n824 );
    and g548 ( n3494 , n193 , n2834 );
    or g549 ( n950 , n516 , n1437 );
    nor g550 ( n238 , n1177 , n1347 );
    and g551 ( n2206 , n2956 , n3097 );
    xnor g552 ( n2461 , n127 , n2636 );
    and g553 ( n2218 , n1100 , n2239 );
    not g554 ( n3330 , n2710 );
    or g555 ( n3519 , n1075 , n804 );
    or g556 ( n63 , n3004 , n1486 );
    or g557 ( n3648 , n5 , n871 );
    xnor g558 ( n1085 , n215 , n614 );
    or g559 ( n2222 , n2591 , n169 );
    nor g560 ( n496 , n3856 , n3347 );
    xnor g561 ( n2723 , n2312 , n2838 );
    or g562 ( n2853 , n1890 , n881 );
    not g563 ( n2098 , n455 );
    or g564 ( n3081 , n2796 , n3088 );
    or g565 ( n3159 , n2589 , n2739 );
    nor g566 ( n1707 , n1070 , n1341 );
    not g567 ( n3748 , n2214 );
    not g568 ( n2766 , n3092 );
    xnor g569 ( n3064 , n2269 , n119 );
    or g570 ( n2920 , n2440 , n303 );
    and g571 ( n1780 , n1639 , n137 );
    and g572 ( n1588 , n3502 , n525 );
    or g573 ( n3129 , n2452 , n3505 );
    xnor g574 ( n3209 , n900 , n2275 );
    nor g575 ( n2348 , n1797 , n3234 );
    or g576 ( n1026 , n1690 , n2273 );
    xor g577 ( n377 , n877 , n1787 );
    xnor g578 ( n3367 , n1542 , n902 );
    not g579 ( n3208 , n2252 );
    and g580 ( n890 , n650 , n3165 );
    not g581 ( n1297 , n490 );
    xnor g582 ( n2687 , n1150 , n243 );
    xnor g583 ( n125 , n487 , n3198 );
    xnor g584 ( n1145 , n2573 , n878 );
    not g585 ( n947 , n705 );
    or g586 ( n669 , n94 , n2499 );
    and g587 ( n2890 , n3466 , n3894 );
    not g588 ( n734 , n1616 );
    xnor g589 ( n2814 , n83 , n2317 );
    or g590 ( n3620 , n2994 , n782 );
    nor g591 ( n3181 , n1406 , n3671 );
    xnor g592 ( n3285 , n343 , n2343 );
    not g593 ( n2568 , n1882 );
    and g594 ( n1322 , n2151 , n2254 );
    or g595 ( n345 , n3795 , n3255 );
    xnor g596 ( n3548 , n3633 , n50 );
    xnor g597 ( n1686 , n1265 , n1659 );
    nor g598 ( n1866 , n1390 , n877 );
    or g599 ( n338 , n3585 , n1789 );
    and g600 ( n946 , n1329 , n1953 );
    not g601 ( n1706 , n3615 );
    or g602 ( n2299 , n988 , n1518 );
    xor g603 ( n378 , n1342 , n1134 );
    xnor g604 ( n2367 , n1669 , n3440 );
    not g605 ( n2633 , n4 );
    and g606 ( n2131 , n665 , n3769 );
    or g607 ( n2451 , n3162 , n1019 );
    and g608 ( n25 , n857 , n48 );
    or g609 ( n449 , n1913 , n3503 );
    and g610 ( n2481 , n1731 , n1588 );
    or g611 ( n137 , n2929 , n2238 );
    and g612 ( n1422 , n2695 , n3363 );
    or g613 ( n1132 , n3553 , n2780 );
    and g614 ( n3595 , n2914 , n2582 );
    or g615 ( n2154 , n182 , n2875 );
    xnor g616 ( n2205 , n1714 , n1534 );
    or g617 ( n2904 , n2174 , n280 );
    xnor g618 ( n2081 , n1350 , n1239 );
    and g619 ( n51 , n3737 , n1438 );
    and g620 ( n1359 , n2883 , n1762 );
    or g621 ( n444 , n2895 , n2498 );
    nor g622 ( n1765 , n3186 , n2206 );
    not g623 ( n11 , n1793 );
    and g624 ( n1568 , n2507 , n2251 );
    not g625 ( n1011 , n1432 );
    and g626 ( n2754 , n1225 , n3009 );
    xnor g627 ( n159 , n442 , n2927 );
    or g628 ( n3093 , n3723 , n3265 );
    xnor g629 ( n3770 , n53 , n519 );
    not g630 ( n150 , n3049 );
    or g631 ( n968 , n2000 , n3772 );
    or g632 ( n2716 , n716 , n3235 );
    xnor g633 ( n2349 , n2725 , n1395 );
    xnor g634 ( n2215 , n980 , n2718 );
    not g635 ( n2592 , n3481 );
    not g636 ( n2265 , n2371 );
    not g637 ( n1872 , n56 );
    not g638 ( n235 , n794 );
    not g639 ( n1723 , n1938 );
    and g640 ( n2454 , n1210 , n2470 );
    and g641 ( n1594 , n3293 , n2826 );
    and g642 ( n1494 , n1297 , n2276 );
    or g643 ( n2957 , n799 , n1440 );
    nor g644 ( n3432 , n2512 , n1760 );
    xnor g645 ( n2784 , n3547 , n2354 );
    xnor g646 ( n784 , n2792 , n3728 );
    not g647 ( n1662 , n955 );
    and g648 ( n2152 , n262 , n681 );
    or g649 ( n1373 , n3579 , n1197 );
    xnor g650 ( n885 , n619 , n2316 );
    xnor g651 ( n3053 , n923 , n2814 );
    or g652 ( n1896 , n3177 , n3842 );
    not g653 ( n3405 , n3889 );
    nor g654 ( n1728 , n2304 , n1551 );
    and g655 ( n1774 , n1057 , n2549 );
    not g656 ( n3788 , n220 );
    or g657 ( n554 , n1018 , n2001 );
    xnor g658 ( n3473 , n2835 , n1529 );
    not g659 ( n2826 , n1808 );
    and g660 ( n3608 , n505 , n497 );
    or g661 ( n407 , n1975 , n1308 );
    or g662 ( n1082 , n2831 , n3893 );
    xnor g663 ( n212 , n1870 , n1988 );
    not g664 ( n161 , n3384 );
    xnor g665 ( n3828 , n906 , n431 );
    not g666 ( n2271 , n3600 );
    or g667 ( n2948 , n1667 , n2348 );
    or g668 ( n1923 , n3294 , n468 );
    not g669 ( n3150 , n927 );
    xnor g670 ( n442 , n909 , n3532 );
    and g671 ( n167 , n866 , n1367 );
    and g672 ( n2758 , n438 , n1311 );
    and g673 ( n1462 , n3535 , n3067 );
    or g674 ( n562 , n2984 , n2529 );
    xnor g675 ( n392 , n3373 , n2180 );
    and g676 ( n1892 , n3615 , n1240 );
    or g677 ( n1179 , n2633 , n3596 );
    not g678 ( n3877 , n2828 );
    or g679 ( n3586 , n2557 , n2562 );
    xnor g680 ( n2909 , n2854 , n2319 );
    or g681 ( n3795 , n1808 , n2046 );
    and g682 ( n2442 , n1452 , n3064 );
    or g683 ( n685 , n216 , n1053 );
    xnor g684 ( n3146 , n1032 , n3324 );
    xnor g685 ( n418 , n2435 , n3390 );
    xor g686 ( n2199 , n600 , n1764 );
    not g687 ( n20 , n927 );
    or g688 ( n3131 , n3039 , n1567 );
    and g689 ( n2240 , n3541 , n823 );
    not g690 ( n405 , n2664 );
    or g691 ( n262 , n472 , n1545 );
    not g692 ( n2962 , n3465 );
    and g693 ( n3576 , n1368 , n3872 );
    xnor g694 ( n2557 , n3243 , n3592 );
    xnor g695 ( n798 , n1873 , n841 );
    or g696 ( n1288 , n1674 , n3076 );
    xor g697 ( n382 , n2885 , n377 );
    and g698 ( n2087 , n2115 , n2597 );
    not g699 ( n1762 , n1808 );
    or g700 ( n2176 , n1921 , n3846 );
    xnor g701 ( n3823 , n1363 , n1732 );
    not g702 ( n2527 , n3623 );
    not g703 ( n3449 , n1451 );
    and g704 ( n3855 , n2900 , n3667 );
    nor g705 ( n2762 , n2885 , n2948 );
    xnor g706 ( n2346 , n838 , n592 );
    and g707 ( n1382 , n3781 , n1090 );
    not g708 ( n1524 , n2186 );
    or g709 ( n566 , n2882 , n1700 );
    or g710 ( n2506 , n1727 , n3746 );
    or g711 ( n2148 , n1118 , n3225 );
    and g712 ( n3638 , n759 , n2911 );
    or g713 ( n821 , n1051 , n3164 );
    or g714 ( n2034 , n1584 , n3843 );
    and g715 ( n222 , n2965 , n3002 );
    or g716 ( n767 , n3183 , n1150 );
    or g717 ( n42 , n223 , n2131 );
    and g718 ( n556 , n839 , n2336 );
    and g719 ( n2501 , n562 , n2122 );
    or g720 ( n787 , n1164 , n1790 );
    not g721 ( n2955 , n772 );
    xnor g722 ( n2361 , n3282 , n635 );
    or g723 ( n1400 , n288 , n617 );
    or g724 ( n953 , n2537 , n2099 );
    and g725 ( n2421 , n3553 , n2780 );
    and g726 ( n1604 , n3185 , n640 );
    or g727 ( n94 , n3783 , n2766 );
    and g728 ( n2039 , n1007 , n3403 );
    or g729 ( n2042 , n3577 , n587 );
    or g730 ( n3740 , n1836 , n2189 );
    or g731 ( n420 , n550 , n654 );
    and g732 ( n214 , n1799 , n1561 );
    or g733 ( n1010 , n275 , n653 );
    or g734 ( n1772 , n2877 , n3456 );
    and g735 ( n123 , n3123 , n1290 );
    not g736 ( n2239 , n1268 );
    xnor g737 ( n1893 , n2559 , n2204 );
    not g738 ( n2477 , n1432 );
    and g739 ( n3479 , n987 , n791 );
    and g740 ( n359 , n403 , n3249 );
    xnor g741 ( n2574 , n111 , n3270 );
    xnor g742 ( n3232 , n1059 , n45 );
    or g743 ( n610 , n3853 , n2301 );
    not g744 ( n3401 , n2448 );
    not g745 ( n1119 , n670 );
    or g746 ( n1536 , n2623 , n3219 );
    or g747 ( n1301 , n321 , n818 );
    xnor g748 ( n3662 , n306 , n3552 );
    or g749 ( n1777 , n1065 , n2249 );
    xnor g750 ( n544 , n2884 , n3677 );
    or g751 ( n2781 , n3668 , n2856 );
    or g752 ( n2504 , n1165 , n1061 );
    or g753 ( n3282 , n3753 , n2030 );
    xnor g754 ( n2387 , n404 , n369 );
    xnor g755 ( n295 , n2400 , n2454 );
    or g756 ( n1768 , n589 , n1232 );
    and g757 ( n219 , n2178 , n357 );
    nor g758 ( n1242 , n1381 , n1891 );
    xnor g759 ( n3569 , n1137 , n1825 );
    and g760 ( n3841 , n1054 , n651 );
    not g761 ( n417 , n44 );
    xnor g762 ( n1206 , n2527 , n919 );
    xnor g763 ( n2810 , n970 , n3522 );
    or g764 ( n520 , n1861 , n571 );
    or g765 ( n2632 , n584 , n1630 );
    and g766 ( n2336 , n3578 , n1444 );
    or g767 ( n1271 , n3705 , n460 );
    or g768 ( n1067 , n661 , n3383 );
    or g769 ( n630 , n598 , n296 );
    and g770 ( n2096 , n1697 , n3266 );
    or g771 ( n3545 , n3887 , n2099 );
    or g772 ( n53 , n2668 , n1473 );
    or g773 ( n1881 , n1355 , n1232 );
    not g774 ( n1319 , n1944 );
    xnor g775 ( n2405 , n2446 , n1190 );
    xnor g776 ( n3425 , n3082 , n2730 );
    and g777 ( n112 , n2874 , n3784 );
    xnor g778 ( n2089 , n420 , n364 );
    not g779 ( n1393 , n2572 );
    or g780 ( n1922 , n221 , n38 );
    xnor g781 ( n1815 , n2517 , n979 );
    or g782 ( n2317 , n613 , n515 );
    or g783 ( n3711 , n189 , n1814 );
    nor g784 ( n17 , n1399 , n1616 );
    or g785 ( n3087 , n1445 , n3407 );
    or g786 ( n3070 , n1119 , n3356 );
    xnor g787 ( n337 , n1316 , n2599 );
    or g788 ( n774 , n1800 , n2663 );
    or g789 ( n2900 , n237 , n602 );
    not g790 ( n2652 , n3690 );
    or g791 ( n1752 , n3201 , n719 );
    not g792 ( n2644 , n829 );
    not g793 ( n2276 , n1248 );
    or g794 ( n1833 , n3655 , n485 );
    or g795 ( n522 , n3771 , n2856 );
    or g796 ( n2549 , n2700 , n3142 );
    nor g797 ( n2084 , n1554 , n2632 );
    or g798 ( n1520 , n2642 , n3402 );
    or g799 ( n3107 , n160 , n31 );
    not g800 ( n1727 , n3365 );
    and g801 ( n3678 , n3620 , n3624 );
    xnor g802 ( n398 , n1306 , n3411 );
    and g803 ( n961 , n2312 , n1098 );
    nor g804 ( n3555 , n1467 , n519 );
    or g805 ( n1744 , n1662 , n2023 );
    and g806 ( n487 , n1148 , n1081 );
    and g807 ( n2347 , n969 , n2876 );
    not g808 ( n351 , n1638 );
    not g809 ( n2432 , n944 );
    nor g810 ( n1369 , n2573 , n1544 );
    not g811 ( n1552 , n2252 );
    xor g812 ( n1558 , n1898 , n2750 );
    not g813 ( n3771 , n3805 );
    or g814 ( n2063 , n2 , n2901 );
    and g815 ( n3826 , n3241 , n702 );
    not g816 ( n2167 , n422 );
    and g817 ( n3498 , n1905 , n1591 );
    xnor g818 ( n3493 , n604 , n2088 );
    and g819 ( n2763 , n1862 , n1036 );
    not g820 ( n3566 , n1847 );
    nor g821 ( n2412 , n1071 , n687 );
    and g822 ( n3577 , n2560 , n1653 );
    or g823 ( n201 , n524 , n1504 );
    xnor g824 ( n195 , n3569 , n1008 );
    nor g825 ( n708 , n2770 , n828 );
    or g826 ( n1708 , n1890 , n3396 );
    or g827 ( n701 , n2551 , n710 );
    or g828 ( n2695 , n358 , n660 );
    xnor g829 ( n678 , n2330 , n3149 );
    xnor g830 ( n648 , n2161 , n1222 );
    or g831 ( n3195 , n1800 , n273 );
    or g832 ( n494 , n1900 , n1493 );
    xnor g833 ( n2319 , n2373 , n115 );
    or g834 ( n240 , n483 , n3834 );
    or g835 ( n2990 , n1754 , n1466 );
    xnor g836 ( n2765 , n1153 , n1287 );
    or g837 ( n993 , n214 , n399 );
    and g838 ( n55 , n821 , n854 );
    and g839 ( n3865 , n1824 , n3756 );
    and g840 ( n2004 , n3302 , n3228 );
    not g841 ( n3485 , n1212 );
    not g842 ( n816 , n1150 );
    or g843 ( n1338 , n3184 , n3304 );
    not g844 ( n3213 , n504 );
    and g845 ( n2224 , n3250 , n373 );
    or g846 ( n3462 , n1864 , n2335 );
    and g847 ( n1000 , n1669 , n875 );
    not g848 ( n3461 , n274 );
    or g849 ( n2625 , n2422 , n121 );
    not g850 ( n910 , n1294 );
    or g851 ( n474 , n29 , n460 );
    or g852 ( n3450 , n1307 , n675 );
    or g853 ( n3096 , n3726 , n2423 );
    and g854 ( n525 , n2757 , n935 );
    not g855 ( n1104 , n230 );
    xnor g856 ( n3317 , n3388 , n2841 );
    or g857 ( n1354 , n2986 , n1684 );
    and g858 ( n3379 , n2246 , n976 );
    and g859 ( n3565 , n2504 , n267 );
    or g860 ( n1464 , n3613 , n2267 );
    xor g861 ( n3767 , n2320 , n1566 );
    or g862 ( n3085 , n1685 , n1180 );
    and g863 ( n2583 , n2525 , n2198 );
    not g864 ( n2662 , n2727 );
    not g865 ( n1378 , n3775 );
    or g866 ( n1096 , n1039 , n3513 );
    or g867 ( n3624 , n1677 , n3259 );
    and g868 ( n364 , n2475 , n3031 );
    or g869 ( n277 , n2455 , n432 );
    not g870 ( n75 , n1991 );
    or g871 ( n58 , n1827 , n3115 );
    not g872 ( n882 , n991 );
    and g873 ( n1803 , n2213 , n1692 );
    xnor g874 ( n1712 , n260 , n3604 );
    and g875 ( n782 , n3259 , n1677 );
    and g876 ( n3300 , n1957 , n1332 );
    and g877 ( n2521 , n156 , n348 );
    or g878 ( n282 , n2548 , n2766 );
    not g879 ( n733 , n3007 );
    not g880 ( n2052 , n335 );
    not g881 ( n1488 , n2192 );
    or g882 ( n2735 , n3467 , n2881 );
    and g883 ( n2021 , n3431 , n2533 );
    not g884 ( n654 , n2055 );
    and g885 ( n2927 , n1600 , n2091 );
    or g886 ( n2802 , n2800 , n41 );
    xnor g887 ( n3182 , n2746 , n1933 );
    and g888 ( n3895 , n3473 , n3060 );
    not g889 ( n1809 , n1272 );
    xnor g890 ( n3116 , n1863 , n2399 );
    and g891 ( n1920 , n2236 , n1762 );
    or g892 ( n2437 , n110 , n2661 );
    and g893 ( n2085 , n3374 , n727 );
    not g894 ( n1077 , n928 );
    or g895 ( n3143 , n3875 , n1382 );
    and g896 ( n1928 , n953 , n3438 );
    xor g897 ( n964 , n1896 , n2921 );
    and g898 ( n3017 , n2666 , n3751 );
    or g899 ( n2363 , n931 , n353 );
    and g900 ( n561 , n3704 , n840 );
    and g901 ( n1998 , n479 , n2587 );
    and g902 ( n2601 , n2110 , n185 );
    or g903 ( n1570 , n1327 , n1771 );
    not g904 ( n1649 , n2349 );
    xnor g905 ( n1006 , n1881 , n3425 );
    or g906 ( n49 , n1355 , n2094 );
    xnor g907 ( n2715 , n1962 , n2120 );
    or g908 ( n768 , n1388 , n3775 );
    nor g909 ( n1935 , n2561 , n1111 );
    not g910 ( n581 , n770 );
    or g911 ( n385 , n208 , n2318 );
    or g912 ( n179 , n1082 , n384 );
    xnor g913 ( n477 , n3662 , n2574 );
    not g914 ( n1495 , n842 );
    or g915 ( n1909 , n3779 , n3584 );
    xnor g916 ( n177 , n1954 , n2788 );
    not g917 ( n1204 , n1461 );
    xnor g918 ( n1825 , n333 , n89 );
    or g919 ( n1927 , n2317 , n3492 );
    not g920 ( n1720 , n3401 );
    and g921 ( n844 , n985 , n3526 );
    and g922 ( n3647 , n2226 , n1984 );
    not g923 ( n2093 , n1874 );
    and g924 ( n1732 , n2002 , n201 );
    xnor g925 ( n1598 , n3488 , n2410 );
    nor g926 ( n2534 , n1947 , n2683 );
    and g927 ( n895 , n121 , n2422 );
    and g928 ( n3049 , n3598 , n2145 );
    or g929 ( n3010 , n2326 , n1473 );
    and g930 ( n1062 , n1820 , n1507 );
    or g931 ( n981 , n2886 , n3588 );
    xnor g932 ( n1609 , n3294 , n3645 );
    or g933 ( n2476 , n1363 , n1495 );
    and g934 ( n2940 , n1385 , n3626 );
    not g935 ( n331 , n66 );
    xnor g936 ( n2064 , n762 , n2225 );
    and g937 ( n852 , n2090 , n742 );
    xnor g938 ( n1254 , n512 , n580 );
    and g939 ( n2388 , n1579 , n233 );
    xnor g940 ( n3076 , n552 , n3727 );
    xnor g941 ( n1298 , n1042 , n706 );
    or g942 ( n2198 , n3803 , n1456 );
    or g943 ( n2624 , n1836 , n3200 );
    and g944 ( n1491 , n3434 , n3469 );
    not g945 ( n2922 , n866 );
    or g946 ( n317 , n2717 , n2101 );
    xnor g947 ( n2991 , n372 , n2711 );
    and g948 ( n3089 , n3119 , n1429 );
    or g949 ( n3453 , n299 , n845 );
    nor g950 ( n3048 , n1747 , n3640 );
    and g951 ( n1047 , n1103 , n1234 );
    and g952 ( n3497 , n3240 , n2137 );
    or g953 ( n2159 , n2115 , n2597 );
    xnor g954 ( n743 , n2780 , n3553 );
    xnor g955 ( n1314 , n3298 , n732 );
    and g956 ( n1769 , n3376 , n2032 );
    xnor g957 ( n2359 , n1453 , n508 );
    xnor g958 ( n3028 , n159 , n709 );
    or g959 ( n2445 , n2053 , n3863 );
    nor g960 ( n3842 , n1883 , n2409 );
    xnor g961 ( n1531 , n3724 , n3106 );
    or g962 ( n3299 , n3348 , n1214 );
    xnor g963 ( n850 , n2957 , n2595 );
    not g964 ( n1075 , n181 );
    and g965 ( n776 , n2118 , n938 );
    or g966 ( n1450 , n3835 , n1503 );
    and g967 ( n470 , n1541 , n1387 );
    or g968 ( n999 , n3767 , n3328 );
    or g969 ( n591 , n3382 , n2332 );
    not g970 ( n1836 , n1202 );
    not g971 ( n908 , n3506 );
    and g972 ( n3297 , n3161 , n173 );
    or g973 ( n2458 , n2548 , n1929 );
    xnor g974 ( n1648 , n886 , n3548 );
    xnor g975 ( n3086 , n3490 , n3456 );
    xnor g976 ( n1529 , n51 , n1514 );
    not g977 ( n245 , n2110 );
    or g978 ( n2151 , n3117 , n1201 );
    and g979 ( n2790 , n1478 , n527 );
    or g980 ( n2868 , n1880 , n898 );
    and g981 ( n1341 , n2601 , n803 );
    xnor g982 ( n2599 , n3012 , n565 );
    not g983 ( n2357 , n2371 );
    xnor g984 ( n93 , n1311 , n723 );
    or g985 ( n2688 , n2516 , n672 );
    or g986 ( n2142 , n2432 , n3233 );
    or g987 ( n1855 , n363 , n1175 );
    xnor g988 ( n280 , n2425 , n3892 );
    xnor g989 ( n1203 , n3640 , n3110 );
    not g990 ( n2947 , n1880 );
    and g991 ( n3726 , n3167 , n2813 );
    or g992 ( n2703 , n1186 , n3895 );
    not g993 ( n802 , n2139 );
    or g994 ( n3735 , n3490 , n1109 );
    or g995 ( n1799 , n2155 , n3665 );
    and g996 ( n2241 , n3738 , n2731 );
    and g997 ( n465 , n744 , n2678 );
    nor g998 ( n217 , n2886 , n897 );
    or g999 ( n2479 , n3246 , n2021 );
    or g1000 ( n979 , n0 , n2743 );
    or g1001 ( n2966 , n3485 , n618 );
    or g1002 ( n1587 , n929 , n545 );
    and g1003 ( n3027 , n177 , n611 );
    or g1004 ( n3331 , n2268 , n3030 );
    or g1005 ( n3399 , n3309 , n1269 );
    not g1006 ( n1365 , n1782 );
    or g1007 ( n905 , n1749 , n1474 );
    or g1008 ( n1022 , n1573 , n351 );
    nor g1009 ( n2546 , n1359 , n2524 );
    not g1010 ( n2541 , n2523 );
    xnor g1011 ( n1606 , n479 , n383 );
    not g1012 ( n2577 , n940 );
    nor g1013 ( n939 , n3231 , n1833 );
    or g1014 ( n3011 , n1051 , n3189 );
    or g1015 ( n1639 , n2431 , n3607 );
    and g1016 ( n3866 , n1522 , n2476 );
    or g1017 ( n2829 , n474 , n1476 );
    not g1018 ( n1012 , n15 );
    xnor g1019 ( n2071 , n1936 , n3564 );
    and g1020 ( n102 , n226 , n1873 );
    and g1021 ( n992 , n1316 , n3012 );
    xnor g1022 ( n1759 , n511 , n126 );
    and g1023 ( n3080 , n3840 , n2610 );
    xnor g1024 ( n553 , n3617 , n1803 );
    or g1025 ( n3567 , n2143 , n3524 );
    or g1026 ( n1188 , n1942 , n3196 );
    xnor g1027 ( n2915 , n651 , n1941 );
    and g1028 ( n1788 , n1644 , n3798 );
    not g1029 ( n2086 , n3718 );
    and g1030 ( n3336 , n741 , n1681 );
    and g1031 ( n2201 , n551 , n3299 );
    xnor g1032 ( n3832 , n2010 , n36 );
    xnor g1033 ( n3636 , n3395 , n2987 );
    xnor g1034 ( n73 , n104 , n2391 );
    or g1035 ( n1448 , n581 , n654 );
    xnor g1036 ( n132 , n972 , n398 );
    or g1037 ( n2414 , n116 , n1650 );
    not g1038 ( n3741 , n1938 );
    not g1039 ( n1782 , n145 );
    xor g1040 ( n3428 , n2710 , n1717 );
    not g1041 ( n3173 , n874 );
    not g1042 ( n3026 , n873 );
    and g1043 ( n3797 , n3633 , n886 );
    or g1044 ( n1645 , n1924 , n1838 );
    or g1045 ( n2614 , n1254 , n1281 );
    not g1046 ( n859 , n1280 );
    xnor g1047 ( n3169 , n3007 , n3014 );
    xnor g1048 ( n1133 , n500 , n975 );
    and g1049 ( n769 , n1830 , n40 );
    or g1050 ( n1235 , n2938 , n1263 );
    xnor g1051 ( n785 , n3478 , n2274 );
    xnor g1052 ( n1525 , n3419 , n3585 );
    or g1053 ( n970 , n3213 , n1269 );
    xnor g1054 ( n3408 , n1766 , n1377 );
    xnor g1055 ( n41 , n457 , n3029 );
    or g1056 ( n3295 , n769 , n3678 );
    xnor g1057 ( n3552 , n2643 , n197 );
    and g1058 ( n1852 , n517 , n3329 );
    or g1059 ( n211 , n2459 , n3493 );
    xnor g1060 ( n1398 , n1934 , n731 );
    xnor g1061 ( n480 , n3370 , n683 );
    not g1062 ( n2875 , n3092 );
    and g1063 ( n2295 , n2712 , n3762 );
    not g1064 ( n3572 , n2237 );
    xnor g1065 ( n2787 , n1112 , n2552 );
    xnor g1066 ( n509 , n2081 , n1661 );
    or g1067 ( n1125 , n2668 , n2030 );
    xor g1068 ( n1657 , n2804 , n3277 );
    not g1069 ( n983 , n519 );
    not g1070 ( n2657 , n2173 );
    or g1071 ( n3066 , n662 , n1960 );
    or g1072 ( n827 , n3205 , n1435 );
    not g1073 ( n2648 , n1181 );
    xnor g1074 ( n3016 , n637 , n16 );
    not g1075 ( n1503 , n2110 );
    and g1076 ( n3231 , n738 , n1193 );
    and g1077 ( n2628 , n114 , n2608 );
    and g1078 ( n468 , n2471 , n151 );
    or g1079 ( n2946 , n66 , n3450 );
    or g1080 ( n2647 , n1515 , n2149 );
    or g1081 ( n2488 , n2600 , n539 );
    and g1082 ( n1166 , n2108 , n1969 );
    and g1083 ( n2945 , n3269 , n570 );
    or g1084 ( n969 , n3048 , n1875 );
    or g1085 ( n3114 , n249 , n621 );
    or g1086 ( n3759 , n2886 , n2297 );
    xnor g1087 ( n2552 , n110 , n2661 );
    xnor g1088 ( n3186 , n2039 , n2639 );
    and g1089 ( n3271 , n1811 , n2457 );
    xnor g1090 ( n694 , n1428 , n199 );
    or g1091 ( n1350 , n577 , n2242 );
    or g1092 ( n1129 , n717 , n2867 );
    xnor g1093 ( n1148 , n3037 , n2376 );
    or g1094 ( n2228 , n2442 , n142 );
    or g1095 ( n1653 , n3606 , n366 );
    or g1096 ( n1225 , n1663 , n1509 );
    or g1097 ( n3221 , n543 , n561 );
    not g1098 ( n613 , n523 );
    xor g1099 ( n1229 , n2288 , n2694 );
    or g1100 ( n2137 , n3153 , n3741 );
    xnor g1101 ( n1894 , n3325 , n3697 );
    or g1102 ( n2006 , n465 , n252 );
    or g1103 ( n2002 , n707 , n3351 );
    and g1104 ( n2283 , n2564 , n2924 );
    or g1105 ( n1741 , n3387 , n2421 );
    or g1106 ( n3568 , n2824 , n3874 );
    xor g1107 ( n1123 , n607 , n1947 );
    not g1108 ( n368 , n3481 );
    xnor g1109 ( n2942 , n2932 , n539 );
    not g1110 ( n3573 , n44 );
    xor g1111 ( n1764 , n867 , n3804 );
    and g1112 ( n1895 , n3778 , n1531 );
    not g1113 ( n2770 , n1085 );
    xnor g1114 ( n1251 , n2676 , n657 );
    xnor g1115 ( n1750 , n499 , n3891 );
    not g1116 ( n3319 , n770 );
    xnor g1117 ( n1272 , n1187 , n19 );
    and g1118 ( n3435 , n3398 , n2975 );
    xnor g1119 ( n723 , n3369 , n3317 );
    not g1120 ( n2505 , n449 );
    or g1121 ( n3364 , n1278 , n558 );
    or g1122 ( n1478 , n116 , n3461 );
    not g1123 ( n3897 , n248 );
    or g1124 ( n695 , n1843 , n3508 );
    or g1125 ( n1244 , n2907 , n1262 );
    xnor g1126 ( n2671 , n672 , n3484 );
    and g1127 ( n713 , n2890 , n117 );
    or g1128 ( n3591 , n3064 , n1452 );
    or g1129 ( n1431 , n417 , n2379 );
    or g1130 ( n428 , n3543 , n3062 );
    not g1131 ( n704 , n493 );
    or g1132 ( n1031 , n3319 , n606 );
    or g1133 ( n2397 , n1691 , n3878 );
    or g1134 ( n333 , n2652 , n1694 );
    nor g1135 ( n3607 , n3063 , n3681 );
    xnor g1136 ( n1859 , n2910 , n1575 );
    or g1137 ( n3175 , n1241 , n1609 );
    or g1138 ( n2269 , n3827 , n441 );
    and g1139 ( n3679 , n2125 , n2075 );
    and g1140 ( n43 , n1373 , n200 );
    not g1141 ( n2293 , n2496 );
    or g1142 ( n703 , n2159 , n2788 );
    nor g1143 ( n3455 , n3816 , n749 );
    or g1144 ( n2738 , n1127 , n3659 );
    not g1145 ( n1379 , n922 );
    or g1146 ( n1110 , n3670 , n318 );
    xnor g1147 ( n1816 , n1241 , n1617 );
    not g1148 ( n1131 , n2726 );
    or g1149 ( n3864 , n570 , n3269 );
    nor g1150 ( n2292 , n2720 , n2736 );
    or g1151 ( n1310 , n821 , n854 );
    not g1152 ( n1402 , n2744 );
    not g1153 ( n3843 , n1914 );
    xnor g1154 ( n2466 , n2828 , n1628 );
    xnor g1155 ( n1693 , n808 , n2248 );
    and g1156 ( n545 , n3350 , n10 );
    nor g1157 ( n2272 , n2554 , n1578 );
    or g1158 ( n2116 , n2341 , n1599 );
    xnor g1159 ( n2908 , n2695 , n1412 );
    not g1160 ( n1007 , n433 );
    xnor g1161 ( n2967 , n1539 , n3218 );
    or g1162 ( n812 , n3800 , n3291 );
    or g1163 ( n1250 , n2417 , n664 );
    xnor g1164 ( n292 , n3646 , n1679 );
    not g1165 ( n3630 , n3536 );
    xnor g1166 ( n3262 , n991 , n2940 );
    or g1167 ( n2791 , n528 , n2575 );
    nor g1168 ( n2362 , n2051 , n507 );
    xnor g1169 ( n2104 , n173 , n359 );
    or g1170 ( n1796 , n2324 , n2168 );
    and g1171 ( n16 , n1416 , n3283 );
    not g1172 ( n1371 , n1280 );
    and g1173 ( n2150 , n2344 , n2411 );
    and g1174 ( n3341 , n1403 , n420 );
    not g1175 ( n998 , n1570 );
    nor g1176 ( n2051 , n1013 , n2390 );
    nor g1177 ( n1551 , n1117 , n3899 );
    and g1178 ( n3293 , n2894 , n3614 );
    xor g1179 ( n872 , n229 , n3180 );
    not g1180 ( n2684 , n3444 );
    or g1181 ( n524 , n1084 , n515 );
    or g1182 ( n3400 , n1256 , n2555 );
    and g1183 ( n2256 , n838 , n34 );
    or g1184 ( n1673 , n1594 , n1060 );
    or g1185 ( n421 , n1295 , n435 );
    xnor g1186 ( n1101 , n459 , n3069 );
    not g1187 ( n3443 , n2202 );
    not g1188 ( n3829 , n2112 );
    xnor g1189 ( n3357 , n3679 , n1831 );
    not g1190 ( n2539 , n1507 );
    and g1191 ( n3071 , n3338 , n1673 );
    xnor g1192 ( n427 , n121 , n513 );
    xnor g1193 ( n2443 , n2822 , n1914 );
    not g1194 ( n310 , n955 );
    and g1195 ( n231 , n1207 , n1508 );
    not g1196 ( n1440 , n28 );
    not g1197 ( n1270 , n1140 );
    not g1198 ( n1987 , n772 );
    not g1199 ( n514 , n1345 );
    xor g1200 ( n2261 , n1588 , n622 );
    xnor g1201 ( n2704 , n2533 , n3246 );
    and g1202 ( n537 , n3111 , n3511 );
    or g1203 ( n586 , n682 , n3511 );
    or g1204 ( n2356 , n249 , n3104 );
    not g1205 ( n965 , n3372 );
    or g1206 ( n2524 , n3052 , n3641 );
    or g1207 ( n1423 , n3509 , n1064 );
    not g1208 ( n748 , n220 );
    not g1209 ( n374 , n127 );
    and g1210 ( n472 , n3400 , n1756 );
    and g1211 ( n3215 , n3131 , n3812 );
    xnor g1212 ( n3310 , n1179 , n522 );
    and g1213 ( n534 , n2598 , n3651 );
    or g1214 ( n967 , n3622 , n3144 );
    and g1215 ( n3019 , n3792 , n188 );
    and g1216 ( n3587 , n2402 , n2727 );
    and g1217 ( n707 , n1504 , n524 );
    and g1218 ( n3244 , n626 , n2979 );
    xnor g1219 ( n3793 , n3252 , n86 );
    or g1220 ( n636 , n1477 , n1517 );
    or g1221 ( n2053 , n182 , n2679 );
    and g1222 ( n3707 , n62 , n3545 );
    not g1223 ( n332 , n162 );
    xor g1224 ( n106 , n3032 , n1853 );
    or g1225 ( n3304 , n3520 , n997 );
    not g1226 ( n210 , n3631 );
    or g1227 ( n2849 , n2014 , n924 );
    xnor g1228 ( n1255 , n178 , n995 );
    or g1229 ( n801 , n3771 , n2229 );
    xnor g1230 ( n1798 , n70 , n861 );
    and g1231 ( n1680 , n325 , n3073 );
    not g1232 ( n1499 , n2031 );
    not g1233 ( n1972 , n2112 );
    not g1234 ( n563 , n3805 );
    and g1235 ( n3846 , n2917 , n1842 );
    or g1236 ( n2525 , n3284 , n3722 );
    and g1237 ( n3149 , n1997 , n3099 );
    nor g1238 ( n458 , n2975 , n3398 );
    and g1239 ( n2056 , n3688 , n2011 );
    xor g1240 ( n3255 , n237 , n2619 );
    xnor g1241 ( n2785 , n3125 , n3736 );
    or g1242 ( n1122 , n1485 , n2769 );
    xnor g1243 ( n1409 , n1768 , n1819 );
    not g1244 ( n321 , n3506 );
    xnor g1245 ( n3259 , n1253 , n3146 );
    or g1246 ( n394 , n1633 , n3748 );
    not g1247 ( n2655 , n3365 );
    xnor g1248 ( n3710 , n2359 , n3542 );
    or g1249 ( n3123 , n1925 , n2175 );
    or g1250 ( n1847 , n2326 , n2311 );
    and g1251 ( n1276 , n2821 , n1323 );
    xnor g1252 ( n1236 , n3089 , n3702 );
    not g1253 ( n15 , n3077 );
    xor g1254 ( n1219 , n1359 , n2638 );
    nor g1255 ( n3844 , n3765 , n1436 );
    xnor g1256 ( n1173 , n2965 , n3616 );
    and g1257 ( n593 , n1746 , n1939 );
    xnor g1258 ( n884 , n41 , n1696 );
    and g1259 ( n3313 , n2909 , n2540 );
    and g1260 ( n1792 , n1544 , n2573 );
    and g1261 ( n1054 , n1687 , n3204 );
    and g1262 ( n3115 , n3453 , n3852 );
    xnor g1263 ( n1496 , n2041 , n3136 );
    or g1264 ( n2166 , n329 , n2887 );
    not g1265 ( n3574 , n1387 );
    or g1266 ( n3762 , n2446 , n3618 );
    not g1267 ( n1002 , n3589 );
    not g1268 ( n2615 , n852 );
    nor g1269 ( n24 , n1989 , n2086 );
    xnor g1270 ( n841 , n1326 , n3454 );
    or g1271 ( n3118 , n102 , n2753 );
    not g1272 ( n549 , n873 );
    or g1273 ( n839 , n458 , n3214 );
    not g1274 ( n826 , n1361 );
    xnor g1275 ( n3763 , n2486 , n1675 );
    nor g1276 ( n254 , n3134 , n268 );
    or g1277 ( n933 , n195 , n2681 );
    or g1278 ( n155 , n2201 , n3220 );
    not g1279 ( n3437 , n541 );
    xor g1280 ( n1383 , n1989 , n3083 );
    and g1281 ( n921 , n645 , n795 );
    xnor g1282 ( n1258 , n3767 , n3120 );
    or g1283 ( n1905 , n3810 , n2611 );
    or g1284 ( n2631 , n3632 , n901 );
    or g1285 ( n2941 , n2113 , n2485 );
    xnor g1286 ( n2370 , n217 , n2690 );
    and g1287 ( n2964 , n3510 , n2888 );
    not g1288 ( n249 , n3742 );
    or g1289 ( n218 , n3393 , n2846 );
    xnor g1290 ( n1885 , n3053 , n2434 );
    and g1291 ( n3483 , n3221 , n68 );
    and g1292 ( n2492 , n1958 , n2506 );
    not g1293 ( n2280 , n2888 );
    and g1294 ( n1891 , n1010 , n2188 );
    not g1295 ( n2974 , n3690 );
    xnor g1296 ( n3541 , n3374 , n2732 );
    nor g1297 ( n1197 , n2759 , n1379 );
    and g1298 ( n2338 , n2647 , n2774 );
    not g1299 ( n253 , n1209 );
    xnor g1300 ( n3349 , n869 , n1121 );
    and g1301 ( n3640 , n2282 , n793 );
    not g1302 ( n1711 , n1185 );
    or g1303 ( n1637 , n2357 , n960 );
    or g1304 ( n1608 , n2886 , n80 );
    xnor g1305 ( n3816 , n2772 , n1940 );
    or g1306 ( n889 , n2017 , n1978 );
    or g1307 ( n3337 , n3140 , n1211 );
    or g1308 ( n1501 , n550 , n1929 );
    or g1309 ( n1965 , n3468 , n2346 );
    xnor g1310 ( n1837 , n3162 , n1592 );
    or g1311 ( n1207 , n29 , n1246 );
    and g1312 ( n2374 , n673 , n579 );
    or g1313 ( n2911 , n2284 , n3460 );
    or g1314 ( n148 , n174 , n1706 );
    or g1315 ( n2944 , n2847 , n1611 );
    and g1316 ( n2982 , n2419 , n3561 );
    and g1317 ( n529 , n3479 , n1228 );
    and g1318 ( n2420 , n2315 , n3528 );
    nor g1319 ( n3238 , n190 , n1496 );
    not g1320 ( n1444 , n3465 );
    or g1321 ( n2121 , n2541 , n370 );
    not g1322 ( n746 , n1097 );
    not g1323 ( n3649 , n3703 );
    not g1324 ( n2591 , n2757 );
    xnor g1325 ( n1672 , n3143 , n2617 );
    not g1326 ( n577 , n4 );
    not g1327 ( n2302 , n44 );
    xnor g1328 ( n3015 , n1003 , n298 );
    and g1329 ( n2994 , n1188 , n3491 );
    xor g1330 ( n3434 , n1886 , n2388 );
    or g1331 ( n3538 , n3188 , n1374 );
    xnor g1332 ( n900 , n1817 , n788 );
    xor g1333 ( n2921 , n1491 , n2199 );
    or g1334 ( n1199 , n3668 , n2305 );
    or g1335 ( n691 , n2609 , n3003 );
    or g1336 ( n1138 , n2324 , n2787 );
    or g1337 ( n151 , n3240 , n2137 );
    or g1338 ( n3272 , n453 , n2078 );
    not g1339 ( n1065 , n3340 );
    or g1340 ( n1597 , n1967 , n2852 );
    not g1341 ( n3095 , n1202 );
    and g1342 ( n2530 , n2465 , n2707 );
    or g1343 ( n578 , n619 , n2316 );
    or g1344 ( n1346 , n1403 , n420 );
    and g1345 ( n2874 , n352 , n3346 );
    and g1346 ( n1364 , n1695 , n2792 );
    or g1347 ( n349 , n1301 , n2038 );
    or g1348 ( n1253 , n187 , n851 );
    or g1349 ( n1900 , n714 , n3275 );
    or g1350 ( n1901 , n3453 , n3852 );
    xnor g1351 ( n2571 , n2386 , n2836 );
    xnor g1352 ( n2179 , n2130 , n3305 );
    or g1353 ( n548 , n2970 , n3040 );
    not g1354 ( n1414 , n873 );
    or g1355 ( n1474 , n1443 , n2189 );
    or g1356 ( n1428 , n3637 , n441 );
    xnor g1357 ( n3256 , n3815 , n3168 );
    or g1358 ( n2589 , n356 , n2860 );
    or g1359 ( n246 , n3729 , n546 );
    not g1360 ( n3155 , n1494 );
    xnor g1361 ( n1115 , n1418 , n2185 );
    nor g1362 ( n1595 , n100 , n286 );
    or g1363 ( n413 , n533 , n532 );
    or g1364 ( n1195 , n3841 , n555 );
    or g1365 ( n677 , n2444 , n2821 );
    or g1366 ( n1682 , n2977 , n1771 );
    or g1367 ( n1463 , n3753 , n2311 );
    not g1368 ( n1930 , n3537 );
    xnor g1369 ( n121 , n2001 , n440 );
    or g1370 ( n2115 , n2966 , n2120 );
    xnor g1371 ( n489 , n3267 , n1942 );
    or g1372 ( n849 , n2295 , n3313 );
    xnor g1373 ( n3134 , n3857 , n2902 );
    xnor g1374 ( n3033 , n1909 , n3740 );
    and g1375 ( n143 , n2757 , n1273 );
    xnor g1376 ( n2127 , n2540 , n2295 );
    not g1377 ( n1964 , n835 );
    and g1378 ( n3468 , n3658 , n2536 );
    or g1379 ( n697 , n923 , n83 );
    not g1380 ( n606 , n1066 );
    xnor g1381 ( n257 , n3276 , n43 );
    not g1382 ( n3562 , n722 );
    nor g1383 ( n2243 , n958 , n2218 );
    and g1384 ( n1028 , n385 , n1932 );
    xnor g1385 ( n1189 , n1806 , n3230 );
    xnor g1386 ( n3124 , n1082 , n2007 );
    or g1387 ( n1286 , n2641 , n1389 );
    xor g1388 ( n2426 , n3193 , n3494 );
    or g1389 ( n3018 , n2432 , n2167 );
    or g1390 ( n3137 , n2259 , n451 );
    or g1391 ( n3008 , n3316 , n1617 );
    or g1392 ( n945 , n2581 , n3151 );
    not g1393 ( n373 , n2112 );
    not g1394 ( n3507 , n2513 );
    or g1395 ( n3528 , n1724 , n244 );
    or g1396 ( n1829 , n576 , n1270 );
    and g1397 ( n2026 , n392 , n3882 );
    or g1398 ( n3312 , n2928 , n3761 );
    xnor g1399 ( n773 , n3096 , n1867 );
    xnor g1400 ( n2180 , n2102 , n545 );
    or g1401 ( n652 , n576 , n1650 );
    and g1402 ( n3372 , n1748 , n1892 );
    or g1403 ( n3677 , n2280 , n1270 );
    or g1404 ( n2820 , n2616 , n175 );
    not g1405 ( n1943 , n167 );
    and g1406 ( n2301 , n2703 , n2203 );
    xnor g1407 ( n2925 , n74 , n1784 );
    and g1408 ( n1421 , n3901 , n3018 );
    or g1409 ( n3438 , n3026 , n3189 );
    and g1410 ( n3329 , n1220 , n733 );
    or g1411 ( n3540 , n1738 , n227 );
    or g1412 ( n854 , n1414 , n3098 );
    not g1413 ( n671 , n2733 );
    xnor g1414 ( n2642 , n90 , n1425 );
    xor g1415 ( n3075 , n3760 , n3811 );
    xnor g1416 ( n1699 , n1665 , n889 );
    and g1417 ( n729 , n691 , n3389 );
    xnor g1418 ( n2725 , n3471 , n2398 );
    or g1419 ( n683 , n2093 , n845 );
    xor g1420 ( n762 , n1854 , n2964 );
    xnor g1421 ( n2980 , n328 , n2220 );
    or g1422 ( n315 , n2345 , n3619 );
    xnor g1423 ( n919 , n1705 , n1828 );
    or g1424 ( n122 , n2389 , n260 );
    not g1425 ( n1232 , n308 );
    xnor g1426 ( n1218 , n1599 , n474 );
    not g1427 ( n679 , n2567 );
    and g1428 ( n1111 , n701 , n2868 );
    and g1429 ( n1627 , n2446 , n3618 );
    nor g1430 ( n1630 , n2967 , n939 );
    or g1431 ( n2411 , n3633 , n886 );
    and g1432 ( n2513 , n1300 , n2141 );
    and g1433 ( n2544 , n2279 , n3628 );
    and g1434 ( n191 , n971 , n157 );
    or g1435 ( n2767 , n2667 , n1401 );
    and g1436 ( n3112 , n2508 , n313 );
    xnor g1437 ( n2216 , n2811 , n2374 );
    xnor g1438 ( n1224 , n3166 , n3266 );
    not g1439 ( n960 , n3631 );
    or g1440 ( n251 , n1052 , n1860 );
    and g1441 ( n982 , n168 , n328 );
    not g1442 ( n1025 , n942 );
    nor g1443 ( n3043 , n1277 , n1279 );
    not g1444 ( n342 , n2724 );
    or g1445 ( n1256 , n1371 , n3412 );
    or g1446 ( n3480 , n1822 , n2287 );
    or g1447 ( n2515 , n2309 , n970 );
    and g1448 ( n1517 , n1860 , n1052 );
    xnor g1449 ( n1154 , n3477 , n1292 );
    and g1450 ( n2528 , n3393 , n2846 );
    xnor g1451 ( n12 , n277 , n125 );
    or g1452 ( n1472 , n706 , n2160 );
    xnor g1453 ( n2903 , n1695 , n784 );
    or g1454 ( n1865 , n306 , n3290 );
    not g1455 ( n387 , n148 );
    or g1456 ( n2307 , n1126 , n347 );
    or g1457 ( n3160 , n3465 , n785 );
    and g1458 ( n3878 , n1237 , n2713 );
    or g1459 ( n1802 , n66 , n2805 );
    and g1460 ( n3398 , n2542 , n498 );
    not g1461 ( n2840 , n3314 );
    or g1462 ( n2507 , n1680 , n232 );
    and g1463 ( n3672 , n1705 , n3160 );
    xnor g1464 ( n3056 , n1504 , n2558 );
    and g1465 ( n2499 , n3757 , n1448 );
    and g1466 ( n3888 , n228 , n1300 );
    nor g1467 ( n3695 , n2193 , n1326 );
    nor g1468 ( n3534 , n3359 , n39 );
    not g1469 ( n2253 , n1156 );
    xnor g1470 ( n454 , n2512 , n1760 );
    or g1471 ( n2598 , n2665 , n601 );
    xnor g1472 ( n2403 , n1516 , n743 );
    xor g1473 ( n693 , n1410 , n1099 );
    or g1474 ( n3133 , n3702 , n2872 );
    xnor g1475 ( n1912 , n3533 , n1518 );
    or g1476 ( n2389 , n2265 , n858 );
    xnor g1477 ( n3488 , n3237 , n3627 );
    and g1478 ( n2018 , n52 , n2962 );
    and g1479 ( n1345 , n225 , n1081 );
    xnor g1480 ( n1817 , n3332 , n2370 );
    xnor g1481 ( n3627 , n1829 , n2667 );
    nor g1482 ( n2423 , n2897 , n1102 );
    xor g1483 ( n393 , n509 , n3300 );
    or g1484 ( n69 , n628 , n1340 );
    nor g1485 ( n3423 , n2199 , n1078 );
    nor g1486 ( n3328 , n3120 , n1296 );
    or g1487 ( n9 , n2588 , n3527 );
    not g1488 ( n3065 , n3457 );
    xnor g1489 ( n3684 , n2441 , n1028 );
    not g1490 ( n182 , n829 );
    or g1491 ( n3325 , n3095 , n3584 );
    or g1492 ( n3381 , n2310 , n2393 );
    and g1493 ( n1977 , n1877 , n171 );
    not g1494 ( n3059 , n2748 );
    nor g1495 ( n602 , n949 , n3499 );
    xnor g1496 ( n2217 , n2353 , n544 );
    not g1497 ( n3671 , n672 );
    and g1498 ( n2983 , n2495 , n3813 );
    xnor g1499 ( n1592 , n1019 , n3764 );
    or g1500 ( n3848 , n1468 , n1879 );
    or g1501 ( n783 , n2854 , n3837 );
    not g1502 ( n410 , n1006 );
    or g1503 ( n3353 , n3900 , n652 );
    not g1504 ( n1162 , n523 );
    xnor g1505 ( n1926 , n204 , n3480 );
    not g1506 ( n573 , n3333 );
    and g1507 ( n3863 , n716 , n3235 );
    or g1508 ( n1326 , n1427 , n1375 );
    or g1509 ( n87 , n912 , n2852 );
    not g1510 ( n3216 , n66 );
    and g1511 ( n232 , n604 , n49 );
    or g1512 ( n311 , n3814 , n844 );
    xnor g1513 ( n1758 , n2246 , n3385 );
    xnor g1514 ( n1368 , n1922 , n1298 );
    or g1515 ( n1329 , n3297 , n359 );
    xnor g1516 ( n503 , n3093 , n1855 );
    or g1517 ( n805 , n954 , n2891 );
    not g1518 ( n674 , n3691 );
    not g1519 ( n903 , n1176 );
    xnor g1520 ( n842 , n2807 , n3807 );
    nor g1521 ( n2580 , n2830 , n1934 );
    and g1522 ( n2160 , n1042 , n1922 );
    nor g1523 ( n797 , n2638 , n2546 );
    xor g1524 ( n2329 , n2845 , n1001 );
    or g1525 ( n2341 , n2895 , n2061 );
    and g1526 ( n2867 , n259 , n2913 );
    or g1527 ( n937 , n3587 , n2985 );
    nor g1528 ( n1282 , n720 , n1709 );
    xnor g1529 ( n3652 , n250 , n2 );
    not g1530 ( n2929 , n3063 );
    or g1531 ( n491 , n679 , n2973 );
    not g1532 ( n2627 , n1387 );
    xnor g1533 ( n608 , n1451 , n2416 );
    xnor g1534 ( n2014 , n790 , n1912 );
    xnor g1535 ( n3881 , n3853 , n2301 );
    or g1536 ( n330 , n556 , n1595 );
    or g1537 ( n3704 , n1893 , n1322 );
    or g1538 ( n3715 , n1124 , n2501 );
    or g1539 ( n1290 , n2629 , n26 );
    and g1540 ( n2274 , n1351 , n1536 );
    xor g1541 ( n3578 , n195 , n2681 );
    and g1542 ( n1121 , n3094 , n2382 );
    or g1543 ( n2091 , n746 , n128 );
    and g1544 ( n635 , n3258 , n2819 );
    or g1545 ( n985 , n3243 , n283 );
    and g1546 ( n1602 , n3215 , n3116 );
    not g1547 ( n1716 , n414 );
    not g1548 ( n3625 , n316 );
    and g1549 ( n1266 , n2488 , n2200 );
    and g1550 ( n641 , n2008 , n1105 );
    not g1551 ( n162 , n3114 );
    xnor g1552 ( n1360 , n3647 , n3761 );
    xnor g1553 ( n1109 , n3867 , n2764 );
    not g1554 ( n3621 , n3465 );
    and g1555 ( n736 , n2524 , n1359 );
    not g1556 ( n532 , n3898 );
    xnor g1557 ( n755 , n3768 , n3210 );
    xnor g1558 ( n817 , n3186 , n2206 );
    or g1559 ( n1136 , n3202 , n2676 );
    xnor g1560 ( n3853 , n2332 , n1184 );
    xor g1561 ( n3882 , n1943 , n113 );
    and g1562 ( n2745 , n2402 , n181 );
    or g1563 ( n250 , n1662 , n2250 );
    and g1564 ( n2579 , n2987 , n3395 );
    or g1565 ( n2 , n1315 , n1723 );
    xnor g1566 ( n1726 , n477 , n3847 );
    xor g1567 ( n731 , n3222 , n2830 );
    and g1568 ( n2211 , n1576 , n415 );
    or g1569 ( n1037 , n2653 , n3070 );
    and g1570 ( n2193 , n3028 , n2536 );
    or g1571 ( n2584 , n253 , n3145 );
    not g1572 ( n2229 , n2031 );
    xnor g1573 ( n1456 , n1426 , n984 );
    xnor g1574 ( n2391 , n2429 , n1948 );
    or g1575 ( n3197 , n2059 , n25 );
    nor g1576 ( n2062 , n1430 , n1769 );
    xnor g1577 ( n1275 , n2745 , n3251 );
    not g1578 ( n1118 , n3610 );
    xnor g1579 ( n692 , n2367 , n3188 );
    or g1580 ( n3849 , n3232 , n3429 );
    or g1581 ( n1614 , n36 , n3447 );
    xnor g1582 ( n1090 , n2139 , n312 );
    xnor g1583 ( n1779 , n1144 , n3791 );
    or g1584 ( n1171 , n2792 , n1695 );
    or g1585 ( n2428 , n2850 , n3054 );
    xnor g1586 ( n105 , n2019 , n631 );
    xnor g1587 ( n2314 , n667 , n658 );
    not g1588 ( n154 , n3631 );
    and g1589 ( n758 , n2161 , n2162 );
    and g1590 ( n3685 , n3368 , n3469 );
    or g1591 ( n1807 , n3472 , n1597 );
    and g1592 ( n452 , n596 , n1354 );
    xor g1593 ( n3478 , n3333 , n1726 );
    nor g1594 ( n1971 , n2646 , n1857 );
    not g1595 ( n2856 , n196 );
    or g1596 ( n752 , n2253 , n320 );
    or g1597 ( n2219 , n3153 , n1981 );
    xnor g1598 ( n1941 , n1054 , n555 );
    not g1599 ( n2439 , n705 );
    or g1600 ( n501 , n3740 , n1909 );
    xnor g1601 ( n3041 , n1572 , n1568 );
    not g1602 ( n3873 , n709 );
    or g1603 ( n3090 , n635 , n1850 );
    xnor g1604 ( n2719 , n3756 , n688 );
    xnor g1605 ( n1911 , n3118 , n3366 );
    or g1606 ( n1063 , n3638 , n2480 );
    not g1607 ( n2889 , n2717 );
    and g1608 ( n1641 , n3899 , n1117 );
    xnor g1609 ( n3192 , n1814 , n189 );
    xnor g1610 ( n1211 , n2909 , n2127 );
    and g1611 ( n1538 , n2721 , n122 );
    or g1612 ( n3176 , n380 , n2095 );
    xnor g1613 ( n255 , n2137 , n1601 );
    and g1614 ( n3558 , n278 , n1966 );
    and g1615 ( n298 , n2635 , n2930 );
    or g1616 ( n2452 , n809 , n2875 );
    not g1617 ( n3520 , n2760 );
    and g1618 ( n1374 , n1643 , n2367 );
    or g1619 ( n1351 , n2190 , n2749 );
    not g1620 ( n1 , n722 );
    xnor g1621 ( n956 , n1255 , n2586 );
    not g1622 ( n3034 , n1247 );
    xnor g1623 ( n3158 , n2101 , n1980 );
    and g1624 ( n3324 , n2755 , n475 );
    or g1625 ( n1585 , n2723 , n3745 );
    or g1626 ( n3517 , n679 , n1872 );
    or g1627 ( n205 , n685 , n2544 );
    nor g1628 ( n2590 , n2433 , n129 );
    nor g1629 ( n1436 , n3888 , n7 );
    xnor g1630 ( n3452 , n3049 , n447 );
    and g1631 ( n863 , n2604 , n3024 );
    xnor g1632 ( n492 , n2738 , n2040 );
    or g1633 ( n1624 , n444 , n1550 );
    not g1634 ( n3814 , n2547 );
    not g1635 ( n3739 , n1854 );
    or g1636 ( n1862 , n1104 , n2579 );
    or g1637 ( n95 , n3193 , n3494 );
    and g1638 ( n113 , n2110 , n2572 );
    xnor g1639 ( n84 , n3406 , n2708 );
    or g1640 ( n3769 , n1006 , n3660 );
    and g1641 ( n528 , n849 , n2795 );
    or g1642 ( n883 , n3679 , n1831 );
    and g1643 ( n227 , n1250 , n1026 );
    and g1644 ( n2777 , n2972 , n179 );
    and g1645 ( n1613 , n2106 , n2550 );
    not g1646 ( n2793 , n2759 );
    nor g1647 ( n710 , n2947 , n239 );
    not g1648 ( n2743 , n2252 );
    or g1649 ( n457 , n1557 , n1259 );
    and g1650 ( n822 , n2362 , n373 );
    xnor g1651 ( n1840 , n888 , n1729 );
    and g1652 ( n3062 , n1468 , n1879 );
    or g1653 ( n1332 , n2135 , n946 );
    and g1654 ( n3837 , n115 , n2373 );
    nor g1655 ( n3402 , n1521 , n150 );
    and g1656 ( n2529 , n3025 , n2734 );
    or g1657 ( n2570 , n3590 , n2750 );
    or g1658 ( n1753 , n2179 , n1334 );
    and g1659 ( n3861 , n104 , n2429 );
    not g1660 ( n3835 , n493 );
    or g1661 ( n3869 , n3172 , n169 );
    and g1662 ( n1696 , n349 , n1807 );
    or g1663 ( n2711 , n1884 , n3055 );
    not g1664 ( n2430 , n1524 );
    or g1665 ( n3642 , n1350 , n1770 );
    or g1666 ( n596 , n633 , n3148 );
    or g1667 ( n3500 , n3006 , n3884 );
    or g1668 ( n1325 , n3796 , n3374 );
    or g1669 ( n2372 , n1636 , n2133 );
    or g1670 ( n200 , n2793 , n922 );
    or g1671 ( n1749 , n662 , n161 );
    or g1672 ( n877 , n3279 , n3844 );
    and g1673 ( n2646 , n3739 , n2964 );
    not g1674 ( n1870 , n1709 );
    nor g1675 ( n1974 , n1845 , n2293 );
    nor g1676 ( n2690 , n2324 , n397 );
    and g1677 ( n2331 , n103 , n906 );
    and g1678 ( n1956 , n1475 , n753 );
    or g1679 ( n3302 , n1637 , n1166 );
    or g1680 ( n2713 , n2230 , n890 );
    xnor g1681 ( n153 , n3060 , n1186 );
    not g1682 ( n2775 , n3038 );
    not g1683 ( n21 , n1526 );
    or g1684 ( n3268 , n512 , n2879 );
    or g1685 ( n3406 , n2247 , n2394 );
    or g1686 ( n875 , n848 , n1978 );
    xnor g1687 ( n1690 , n2915 , n3504 );
    and g1688 ( n2401 , n2751 , n907 );
    or g1689 ( n2344 , n50 , n3797 );
    or g1690 ( n778 , n145 , n1498 );
    or g1691 ( n516 , n3573 , n3412 );
    xnor g1692 ( n592 , n1228 , n3479 );
    xnor g1693 ( n70 , n2723 , n3745 );
    xnor g1694 ( n2797 , n3070 , n2653 );
    or g1695 ( n552 , n1967 , n2577 );
    or g1696 ( n1631 , n882 , n2940 );
    xnor g1697 ( n2182 , n2076 , n1555 );
    xnor g1698 ( n1142 , n3608 , n106 );
    not g1699 ( n3217 , n2728 );
    and g1700 ( n183 , n3173 , n675 );
    or g1701 ( n3067 , n1966 , n278 );
    nor g1702 ( n3355 , n760 , n112 );
    not g1703 ( n3088 , n1183 );
    or g1704 ( n2863 , n133 , n1047 );
    or g1705 ( n1936 , n3612 , n973 );
    or g1706 ( n3682 , n2222 , n231 );
    xor g1707 ( n2158 , n3790 , n1937 );
    or g1708 ( n2377 , n3215 , n3116 );
    xnor g1709 ( n2978 , n700 , n2378 );
    or g1710 ( n1160 , n1808 , n2630 );
    nor g1711 ( n1164 , n3751 , n2666 );
    and g1712 ( n172 , n2843 , n806 );
    and g1713 ( n2885 , n79 , n1972 );
    not g1714 ( n2438 , n3286 );
    or g1715 ( n2325 , n271 , n3273 );
    xnor g1716 ( n2996 , n3371 , n1672 );
    or g1717 ( n793 , n1652 , n3572 );
    and g1718 ( n2609 , n1542 , n1031 );
    not g1719 ( n2424 , n594 );
    or g1720 ( n2177 , n1489 , n1384 );
    or g1721 ( n753 , n2234 , n965 );
    xnor g1722 ( n2749 , n2623 , n3219 );
    nor g1723 ( n1128 , n2450 , n816 );
    xnor g1724 ( n2617 , n3468 , n2346 );
    and g1725 ( n856 , n1848 , n3822 );
    and g1726 ( n300 , n830 , n1682 );
    or g1727 ( n2697 , n1153 , n1287 );
    not g1728 ( n1856 , n642 );
    and g1729 ( n2747 , n1380 , n762 );
    xnor g1730 ( n3592 , n123 , n3866 );
    or g1731 ( n1353 , n809 , n2794 );
    and g1732 ( n1589 , n3858 , n388 );
    and g1733 ( n2140 , n3291 , n3800 );
    and g1734 ( n1544 , n3500 , n699 );
    xnor g1735 ( n3599 , n287 , n1470 );
    xnor g1736 ( n3110 , n1747 , n1796 );
    xnor g1737 ( n1161 , n3372 , n2234 );
    xnor g1738 ( n726 , n279 , n3595 );
    nor g1739 ( n1528 , n3760 , n820 );
    xnor g1740 ( n3141 , n3358 , n1474 );
    and g1741 ( n336 , n914 , n1801 );
    not g1742 ( n2693 , n3499 );
    or g1743 ( n3490 , n533 , n1626 );
    xnor g1744 ( n735 , n1858 , n480 );
    xnor g1745 ( n1308 , n2568 , n779 );
    xnor g1746 ( n47 , n3269 , n1839 );
    xnor g1747 ( n327 , n3900 , n2865 );
    xnor g1748 ( n513 , n2422 , n1871 );
    or g1749 ( n396 , n2568 , n1442 );
    or g1750 ( n994 , n1443 , n3200 );
    and g1751 ( n215 , n2449 , n3794 );
    not g1752 ( n248 , n3686 );
    not g1753 ( n2425 , n3566 );
    nor g1754 ( n625 , n1853 , n811 );
    not g1755 ( n446 , n230 );
    not g1756 ( n941 , n2245 );
    nor g1757 ( n355 , n537 , n3437 );
    xnor g1758 ( n3738 , n3644 , n1185 );
    and g1759 ( n2472 , n1308 , n1975 );
    and g1760 ( n725 , n1420 , n888 );
    not g1761 ( n1992 , n181 );
    and g1762 ( n1550 , n3184 , n3304 );
    not g1763 ( n2794 , n2744 );
    or g1764 ( n3525 , n343 , n2343 );
    xnor g1765 ( n2864 , n3343 , n1258 );
    and g1766 ( n2759 , n671 , n745 );
    and g1767 ( n1718 , n2612 , n834 );
    or g1768 ( n506 , n1714 , n1534 );
    xnor g1769 ( n604 , n3858 , n1702 );
    not g1770 ( n3632 , n190 );
    not g1771 ( n3098 , n2640 );
    not g1772 ( n1208 , n3321 );
    and g1773 ( n1141 , n1056 , n2482 );
    and g1774 ( n476 , n2458 , n2009 );
    or g1775 ( n2975 , n3465 , n1798 );
    not g1776 ( n1635 , n3032 );
    xnor g1777 ( n2906 , n1623 , n1780 );
    or g1778 ( n3047 , n1557 , n1783 );
    or g1779 ( n2008 , n2537 , n1392 );
    and g1780 ( n1231 , n574 , n1488 );
    not g1781 ( n1209 , n2910 );
    xnor g1782 ( n2246 , n926 , n1199 );
    or g1783 ( n2111 , n2481 , n77 );
    and g1784 ( n2702 , n3508 , n1843 );
    or g1785 ( n1267 , n629 , n1192 );
    or g1786 ( n3078 , n2013 , n3322 );
    and g1787 ( n763 , n2300 , n2497 );
    and g1788 ( n283 , n3866 , n123 );
    or g1789 ( n1906 , n1169 , n1537 );
    and g1790 ( n1640 , n999 , n1549 );
    xnor g1791 ( n2986 , n1703 , n258 );
    xnor g1792 ( n1056 , n717 , n1093 );
    not g1793 ( n3668 , n2912 );
    not g1794 ( n1384 , n2640 );
    not g1795 ( n380 , n3774 );
    or g1796 ( n2954 , n2650 , n845 );
    xnor g1797 ( n1420 , n1330 , n1525 );
    xnor g1798 ( n463 , n3344 , n198 );
    and g1799 ( n366 , n1170 , n1826 );
    nor g1800 ( n3290 , n1719 , n2643 );
    and g1801 ( n2739 , n831 , n1570 );
    or g1802 ( n2812 , n3817 , n3314 );
    xnor g1803 ( n1823 , n1841 , n2123 );
    and g1804 ( n1004 , n436 , n317 );
    not g1805 ( n3660 , n152 );
    or g1806 ( n716 , n1107 , n1402 );
    not g1807 ( n434 , n3631 );
    not g1808 ( n1081 , n66 );
    not g1809 ( n3755 , n940 );
    or g1810 ( n3266 , n1371 , n2379 );
    and g1811 ( n646 , n1606 , n1275 );
    xnor g1812 ( n2138 , n3613 , n3030 );
    or g1813 ( n1824 , n908 , n3755 );
    and g1814 ( n3698 , n1831 , n3679 );
    not g1815 ( n1044 , n1459 );
    and g1816 ( n2778 , n1900 , n937 );
    or g1817 ( n639 , n459 , n3069 );
    xnor g1818 ( n1439 , n1323 , n3516 );
    or g1819 ( n2192 , n3719 , n989 );
    not g1820 ( n2474 , n1820 );
    and g1821 ( n565 , n412 , n3712 );
    and g1822 ( n1008 , n3448 , n2109 );
    and g1823 ( n3030 , n2786 , n3777 );
    and g1824 ( n3202 , n2445 , n2716 );
    or g1825 ( n2382 , n2208 , n3053 );
    xnor g1826 ( n2621 , n31 , n2328 );
    not g1827 ( n2958 , n1191 );
    or g1828 ( n319 , n1693 , n3550 );
    xnor g1829 ( n1540 , n2466 , n2195 );
    not g1830 ( n3227 , n215 );
    xnor g1831 ( n3482 , n214 , n3896 );
    and g1832 ( n2169 , n160 , n31 );
    nor g1833 ( n918 , n981 , n1866 );
    or g1834 ( n3758 , n1669 , n875 );
    xor g1835 ( n869 , n3802 , n470 );
    or g1836 ( n141 , n3630 , n2918 );
    and g1837 ( n482 , n113 , n167 );
    xnor g1838 ( n1980 , n3358 , n2543 );
    not g1839 ( n2607 , n1387 );
    and g1840 ( n2673 , n2424 , n863 );
    or g1841 ( n3204 , n3066 , n1665 );
    not g1842 ( n1411 , n3321 );
    not g1843 ( n2005 , n1874 );
    xnor g1844 ( n1041 , n744 , n3046 );
    or g1845 ( n309 , n1417 , n1737 );
    or g1846 ( n437 , n466 , n1053 );
    xnor g1847 ( n2776 , n2009 , n3130 );
    or g1848 ( n2919 , n775 , n496 );
    nor g1849 ( n2487 , n3236 , n464 );
    xnor g1850 ( n3633 , n1165 , n1133 );
    or g1851 ( n766 , n1075 , n176 );
    or g1852 ( n2855 , n2112 , n2742 );
    and g1853 ( n1334 , n531 , n767 );
    not g1854 ( n2895 , n1156 );
    or g1855 ( n59 , n2768 , n2521 );
    or g1856 ( n3613 , n2284 , n777 );
    or g1857 ( n629 , n1535 , n2250 );
    and g1858 ( n540 , n3514 , n583 );
    nor g1859 ( n1790 , n1159 , n3017 );
    not g1860 ( n294 , n1701 );
    or g1861 ( n2129 , n3519 , n141 );
    not g1862 ( n1650 , n2252 );
    xor g1863 ( n163 , n257 , n2107 );
    and g1864 ( n3196 , n1512 , n3267 );
    or g1865 ( n3342 , n2702 , n1951 );
    or g1866 ( n2406 , n3701 , n3178 );
    or g1867 ( n3688 , n418 , n1282 );
    and g1868 ( n2232 , n393 , n3829 );
    xnor g1869 ( n3250 , n1085 , n828 );
    or g1870 ( n3307 , n380 , n370 );
    xnor g1871 ( n1651 , n3342 , n1903 );
    or g1872 ( n7 , n1260 , n3281 );
    or g1873 ( n2143 , n2907 , n161 );
    or g1874 ( n347 , n3831 , n3754 );
    or g1875 ( n1362 , n3872 , n1368 );
    xnor g1876 ( n3139 , n392 , n666 );
    xnor g1877 ( n3198 , n1645 , n1832 );
    or g1878 ( n1089 , n3380 , n1116 );
    or g1879 ( n750 , n2100 , n1174 );
    and g1880 ( n1437 , n3069 , n2993 );
    or g1881 ( n60 , n242 , n405 );
    or g1882 ( n1461 , n859 , n2922 );
    xnor g1883 ( n3385 , n976 , n3529 );
    and g1884 ( n1014 , n792 , n3268 );
    nor g1885 ( n1058 , n1920 , n827 );
    xnor g1886 ( n2332 , n3716 , n2072 );
    xnor g1887 ( n3277 , n3367 , n492 );
    or g1888 ( n868 , n2401 , n61 );
    not g1889 ( n2516 , n1406 );
    or g1890 ( n1406 , n3582 , n3507 );
    or g1891 ( n810 , n967 , n362 );
    not g1892 ( n589 , n1874 );
    xnor g1893 ( n888 , n2060 , n781 );
    xnor g1894 ( n2231 , n560 , n3611 );
    and g1895 ( n2296 , n1775 , n185 );
    xnor g1896 ( n3819 , n2903 , n1233 );
    xnor g1897 ( n3079 , n3399 , n572 );
    nor g1898 ( n339 , n3609 , n1675 );
    xnor g1899 ( n1396 , n2453 , n3310 );
    and g1900 ( n3896 , n2187 , n2377 );
    or g1901 ( n2378 , n1146 , n1964 );
    xnor g1902 ( n2230 , n271 , n2519 );
    xnor g1903 ( n954 , n48 , n1217 );
    not g1904 ( n1333 , n3510 );
    not g1905 ( n1372 , n1404 );
    not g1906 ( n197 , n1719 );
    xnor g1907 ( n1898 , n2547 , n844 );
    not g1908 ( n3121 , n998 );
    xnor g1909 ( n922 , n1056 , n2286 );
    or g1910 ( n972 , n2538 , n2466 );
    xnor g1911 ( n1729 , n1420 , n2530 );
    and g1912 ( n2244 , n2044 , n1122 );
    xor g1913 ( n738 , n261 , n3881 );
    or g1914 ( n531 , n3336 , n1128 );
    or g1915 ( n160 , n1414 , n405 );
    or g1916 ( n1130 , n3487 , n2290 );
    not g1917 ( n3537 , n727 );
    xor g1918 ( n991 , n2768 , n2521 );
    or g1919 ( n3820 , n2004 , n2240 );
    xnor g1920 ( n1566 , n1399 , n734 );
    xor g1921 ( n2554 , n1348 , n3770 );
    not g1922 ( n800 , n722 );
    not g1923 ( n1510 , n2583 );
    or g1924 ( n3430 , n1396 , n96 );
    or g1925 ( n3187 , n2565 , n3656 );
    or g1926 ( n2560 , n894 , n1487 );
    not g1927 ( n745 , n1168 );
    and g1928 ( n1578 , n1784 , n74 );
    and g1929 ( n1791 , n54 , n2296 );
    or g1930 ( n1029 , n3114 , n2853 );
    not g1931 ( n1392 , n1387 );
    xor g1932 ( n958 , n839 , n1049 );
    or g1933 ( n184 , n2717 , n3750 );
    or g1934 ( n792 , n3689 , n264 );
    not g1935 ( n2977 , n3774 );
    xnor g1936 ( n1975 , n1644 , n3654 );
    or g1937 ( n1005 , n1074 , n2945 );
    or g1938 ( n815 , n2594 , n3596 );
    or g1939 ( n2999 , n2998 , n1751 );
    or g1940 ( n699 , n1671 , n3557 );
    and g1941 ( n1983 , n1405 , n2351 );
    not g1942 ( n2351 , n3105 );
    and g1943 ( n3501 , n1565 , n170 );
    xnor g1944 ( n1853 , n226 , n798 );
    or g1945 ( n1009 , n549 , n2607 );
    and g1946 ( n127 , n2522 , n3602 );
    or g1947 ( n2710 , n2808 , n2926 );
    and g1948 ( n3068 , n2131 , n223 );
    and g1949 ( n1318 , n2951 , n143 );
    or g1950 ( n2910 , n235 , n621 );
    or g1951 ( n18 , n1016 , n2861 );
    xnor g1952 ( n241 , n212 , n1861 );
    and g1953 ( n3100 , n1555 , n2076 );
    and g1954 ( n3278 , n1712 , n766 );
    and g1955 ( n680 , n548 , n1906 );
    not g1956 ( n3650 , n891 );
    xnor g1957 ( n2225 , n1380 , n336 );
    and g1958 ( n1163 , n2639 , n2039 );
    not g1959 ( n3830 , n1273 );
    or g1960 ( n2755 , n3480 , n376 );
    not g1961 ( n3874 , n3495 );
    not g1962 ( n3236 , n2277 );
    not g1963 ( n3681 , n2238 );
    nor g1964 ( n2600 , n2932 , n852 );
    or g1965 ( n2156 , n1083 , n1499 );
    xor g1966 ( n2398 , n389 , n305 );
    or g1967 ( n3594 , n2170 , n294 );
    or g1968 ( n2197 , n786 , n1885 );
    or g1969 ( n2122 , n2734 , n3025 );
    or g1970 ( n700 , n138 , n1723 );
    xnor g1971 ( n657 , n3202 , n528 );
    and g1972 ( n133 , n1541 , n2664 );
    not g1973 ( n1626 , n3321 );
    or g1974 ( n1459 , n2112 , n2741 );
    or g1975 ( n1352 , n3861 , n1948 );
    or g1976 ( n1697 , n285 , n2861 );
    and g1977 ( n2694 , n1520 , n3287 );
    not g1978 ( n459 , n996 );
    xnor g1979 ( n1674 , n103 , n3828 );
    and g1980 ( n395 , n2329 , n54 );
    xnor g1981 ( n1512 , n60 , n32 );
    nor g1982 ( n1375 , n3152 , n2281 );
    xnor g1983 ( n2033 , n822 , n3397 );
    or g1984 ( n2751 , n18 , n371 );
    and g1985 ( n2300 , n879 , n1362 );
    and g1986 ( n988 , n790 , n3533 );
    and g1987 ( n1970 , n1564 , n3488 );
    or g1988 ( n2550 , n1453 , n508 );
    xor g1989 ( n2383 , n664 , n2417 );
    not g1990 ( n216 , n2760 );
    and g1991 ( n2562 , n202 , n847 );
    or g1992 ( n3369 , n1979 , n2037 );
    or g1993 ( n403 , n1916 , n16 );
    or g1994 ( n2467 , n337 , n289 );
    and g1995 ( n269 , n1956 , n3422 );
    or g1996 ( n2995 , n388 , n3858 );
    or g1997 ( n1879 , n2977 , n3650 );
    not g1998 ( n2789 , n3774 );
    xnor g1999 ( n3127 , n2064 , n495 );
    and g2000 ( n363 , n820 , n3760 );
    nor g2001 ( n3420 , n1020 , n449 );
    and g2002 ( n3279 , n7 , n3888 );
    or g2003 ( n1170 , n1439 , n3534 );
    and g2004 ( n2872 , n3089 , n3158 );
    not g2005 ( n1751 , n3615 );
    not g2006 ( n2861 , n88 );
    or g2007 ( n1863 , n3309 , n1246 );
    or g2008 ( n1786 , n1450 , n131 );
    nor g2009 ( n2393 , n2982 , n3512 );
    xnor g2010 ( n3856 , n2237 , n2784 );
    and g2011 ( n1072 , n2217 , n1125 );
    or g2012 ( n287 , n908 , n2663 );
    not g2013 ( n901 , n1496 );
    xnor g2014 ( n3616 , n2800 , n884 );
    nor g2015 ( n3234 , n2232 , n2266 );
    or g2016 ( n3235 , n3705 , n2766 );
    or g2017 ( n916 , n1686 , n780 );
    nor g2018 ( n1070 , n2601 , n803 );
    and g2019 ( n2355 , n3367 , n2738 );
    xnor g2020 ( n1513 , n2700 , n3142 );
    or g2021 ( n114 , n2327 , n3707 );
    and g2022 ( n588 , n2428 , n2262 );
    not g2023 ( n1388 , n183 );
    or g2024 ( n3804 , n2886 , n1189 );
    not g2025 ( n2752 , n2387 );
    not g2026 ( n1246 , n1273 );
    xor g2027 ( n605 , n2453 , n3122 );
    and g2028 ( n2681 , n3549 , n1585 );
    and g2029 ( n1518 , n2043 , n2404 );
    not g2030 ( n662 , n2371 );
    not g2031 ( n473 , n2595 );
    or g2032 ( n2282 , n2354 , n2171 );
    and g2033 ( n1100 , n2837 , n3786 );
    not g2034 ( n3005 , n1791 );
    or g2035 ( n1811 , n3379 , n3529 );
    xnor g2036 ( n3390 , n1484 , n3883 );
    and g2037 ( n3885 , n2372 , n932 );
    or g2038 ( n3712 , n888 , n1420 );
    not g2039 ( n2017 , n2567 );
    or g2040 ( n865 , n1812 , n2590 );
    and g2041 ( n1864 , n2948 , n2885 );
    and g2042 ( n134 , n1532 , n2626 );
    or g2043 ( n1035 , n148 , n3845 );
    or g2044 ( n2798 , n111 , n2756 );
    xnor g2045 ( n3559 , n3124 , n3603 );
    nor g2046 ( n3220 , n1319 , n1294 );
    nor g2047 ( n3780 , n3388 , n3369 );
    or g2048 ( n1403 , n3 , n3659 );
    and g2049 ( n2641 , n1289 , n2631 );
    or g2050 ( n145 , n2016 , n2973 );
    and g2051 ( n490 , n3170 , n3306 );
    or g2052 ( n3441 , n774 , n3080 );
    xnor g2053 ( n448 , n413 , n3169 );
    not g2054 ( n334 , n1066 );
    nor g2055 ( n78 , n1777 , n689 );
    and g2056 ( n555 , n2953 , n554 );
    or g2057 ( n3821 , n3158 , n3089 );
    xnor g2058 ( n2540 , n716 , n1704 );
    nor g2059 ( n3265 , n2368 , n2803 );
    or g2060 ( n1642 , n2056 , n3432 );
    xnor g2061 ( n1623 , n1781 , n568 );
    or g2062 ( n3790 , n1659 , n1265 );
    xnor g2063 ( n1886 , n2135 , n946 );
    not g2064 ( n2679 , n2223 );
    or g2065 ( n2692 , n1869 , n2825 );
    xnor g2066 ( n3487 , n2179 , n1334 );
    and g2067 ( n1913 , n3369 , n3388 );
    xnor g2068 ( n3709 , n1244 , n391 );
    or g2069 ( n1458 , n3229 , n19 );
    or g2070 ( n2097 , n1181 , n2079 );
    not g2071 ( n2345 , n998 );
    and g2072 ( n3292 , n1648 , n2578 );
    or g2073 ( n226 , n542 , n1813 );
    xnor g2074 ( n3604 , n2389 , n2933 );
    xnor g2075 ( n2352 , n3839 , n1116 );
    nor g2076 ( n3205 , n3653 , n2211 );
    not g2077 ( n2249 , n2223 );
    or g2078 ( n2795 , n2540 , n2909 );
    xnor g2079 ( n37 , n799 , n28 );
    xnor g2080 ( n2161 , n2578 , n1261 );
    xnor g2081 ( n361 , n455 , n98 );
    xnor g2082 ( n2685 , n236 , n2689 );
    or g2083 ( n2686 , n1519 , n1276 );
    and g2084 ( n1245 , n3312 , n3113 );
    not g2085 ( n460 , n2055 );
    xnor g2086 ( n164 , n1020 , n1897 );
    not g2087 ( n176 , n3898 );
    xnor g2088 ( n2058 , n366 , n894 );
    and g2089 ( n2408 , n3824 , n3474 );
    not g2090 ( n1748 , n1199 );
    and g2091 ( n3351 , n1927 , n697 );
    or g2092 ( n83 , n310 , n3446 );
    not g2093 ( n230 , n1591 );
    xnor g2094 ( n1702 , n2910 , n30 );
    xnor g2095 ( n194 , n2759 , n3579 );
    nor g2096 ( n1838 , n1818 , n1155 );
    not g2097 ( n90 , n3772 );
    or g2098 ( n3703 , n704 , n2935 );
    or g2099 ( n1740 , n1998 , n1668 );
    or g2100 ( n1024 , n107 , n1335 );
    or g2101 ( n2792 , n1742 , n1402 );
    and g2102 ( n929 , n3373 , n2102 );
    and g2103 ( n2869 , n1418 , n3518 );
    or g2104 ( n1565 , n921 , n2026 );
    xnor g2105 ( n3871 , n2731 , n3605 );
    or g2106 ( n384 , n1994 , n245 );
    not g2107 ( n2157 , n618 );
    not g2108 ( n2419 , n572 );
    or g2109 ( n1647 , n2017 , n3562 );
    not g2110 ( n777 , n2055 );
    or g2111 ( n3765 , n2324 , n2205 );
    or g2112 ( n2213 , n1285 , n1055 );
    xnor g2113 ( n622 , n1207 , n3657 );
    not g2114 ( n1083 , n794 );
    not g2115 ( n574 , n2219 );
    or g2116 ( n3345 , n3213 , n2249 );
    nor g2117 ( n2803 , n395 , n330 );
    xnor g2118 ( n984 , n3195 , n2777 );
    not g2119 ( n265 , n3411 );
    xnor g2120 ( n747 , n3259 , n2994 );
    or g2121 ( n3701 , n2594 , n2955 );
    xnor g2122 ( n1921 , n954 , n3285 );
    not g2123 ( n2350 , n835 );
    nor g2124 ( n3531 , n2648 , n1469 );
    not g2125 ( n356 , n2888 );
    or g2126 ( n2118 , n3736 , n1739 );
    or g2127 ( n3168 , n1573 , n2379 );
    and g2128 ( n2343 , n22 , n1288 );
    xnor g2129 ( n2469 , n2612 , n1014 );
    not g2130 ( n3023 , n322 );
    not g2131 ( n147 , n770 );
    or g2132 ( n2968 , n2400 , n2454 );
    or g2133 ( n209 , n389 , n3471 );
    xnor g2134 ( n1677 , n1087 , n1465 );
    not g2135 ( n3556 , n1202 );
    and g2136 ( n3629 , n282 , n630 );
    not g2137 ( n1300 , n2886 );
    xnor g2138 ( n1187 , n922 , n194 );
    not g2139 ( n996 , n2993 );
    or g2140 ( n741 , n1040 , n3244 );
    or g2141 ( n1596 , n191 , n3278 );
    or g2142 ( n3824 , n2685 , n219 );
    not g2143 ( n1269 , n935 );
    or g2144 ( n3154 , n3037 , n1915 );
    or g2145 ( n3894 , n3822 , n1848 );
    xnor g2146 ( n3243 , n1169 , n1523 );
    xor g2147 ( n2368 , n2948 , n382 );
    or g2148 ( n1973 , n3079 , n757 );
    and g2149 ( n3322 , n1887 , n2625 );
    and g2150 ( n3687 , n1993 , n511 );
    xnor g2151 ( n1257 , n1975 , n776 );
    xnor g2152 ( n1581 , n3004 , n1478 );
    nor g2153 ( n3303 , n183 , n1378 );
    or g2154 ( n535 , n1858 , n683 );
    xnor g2155 ( n2862 , n1176 , n3272 );
    xnor g2156 ( n2092 , n47 , n433 );
    nor g2157 ( n1664 , n1097 , n3360 );
    not g2158 ( n640 , n1808 );
    nor g2159 ( n1655 , n1094 , n2943 );
    or g2160 ( n2971 , n3883 , n1386 );
    and g2161 ( n987 , n2124 , n2111 );
    or g2162 ( n2566 , n3616 , n222 );
    xnor g2163 ( n808 , n1757 , n429 );
    not g2164 ( n1473 , n2258 );
    or g2165 ( n2429 , n826 , n2287 );
    or g2166 ( n2707 , n3709 , n3646 );
    or g2167 ( n139 , n869 , n3056 );
    and g2168 ( n3148 , n1684 , n2986 );
    nor g2169 ( n1078 , n1491 , n1896 );
    or g2170 ( n500 , n358 , n158 );
    nor g2171 ( n3199 , n1003 , n298 );
    xnor g2172 ( n304 , n1117 , n2304 );
    or g2173 ( n2924 , n1819 , n1768 );
    or g2174 ( n2190 , n1216 , n541 );
    and g2175 ( n149 , n1045 , n1135 );
    and g2176 ( n1979 , n566 , n2105 );
    or g2177 ( n68 , n2098 , n98 );
    or g2178 ( n3731 , n1944 , n910 );
    not g2179 ( n401 , n824 );
    or g2180 ( n709 , n1876 , n708 );
    not g2181 ( n2023 , n2664 );
    xnor g2182 ( n567 , n626 , n1040 );
    not g2183 ( n1967 , n185 );
    not g2184 ( n135 , n1095 );
    nor g2185 ( n3475 , n1138 , n2427 );
    xnor g2186 ( n1453 , n1857 , n1419 );
    or g2187 ( n2989 , n1371 , n2510 );
    xnor g2188 ( n391 , n1365 , n3734 );
    xnor g2189 ( n1572 , n1758 , n2207 );
    and g2190 ( n1737 , n423 , n883 );
    or g2191 ( n840 , n2559 , n2204 );
    and g2192 ( n1502 , n2101 , n536 );
    and g2193 ( n61 , n2867 , n717 );
    not g2194 ( n2831 , n185 );
    or g2195 ( n1605 , n1162 , n3597 );
    not g2196 ( n2189 , n56 );
    and g2197 ( n1190 , n3417 , n445 );
    xnor g2198 ( n3720 , n643 , n1360 );
    xnor g2199 ( n893 , n2238 , n2827 );
    xnor g2200 ( n2366 , n1044 , n1090 );
    xor g2201 ( n2815 , n1052 , n1477 );
    xnor g2202 ( n383 , n1969 , n1668 );
    not g2203 ( n2184 , n935 );
    and g2204 ( n3045 , n1244 , n2658 );
    and g2205 ( n1335 , n522 , n1179 );
    and g2206 ( n89 , n718 , n2649 );
    and g2207 ( n751 , n2332 , n3382 );
    and g2208 ( n3845 , n1858 , n683 );
    and g2209 ( n1880 , n2944 , n2129 );
    xnor g2210 ( n1628 , n742 , n3426 );
    or g2211 ( n1625 , n953 , n3438 );
    or g2212 ( n1755 , n3274 , n3439 );
    or g2213 ( n878 , n2886 , n1779 );
    or g2214 ( n737 , n748 , n38 );
    or g2215 ( n1330 , n2191 , n1960 );
    and g2216 ( n3554 , n3076 , n1674 );
    not g2217 ( n550 , n944 );
    and g2218 ( n3020 , n1990 , n700 );
    nor g2219 ( n1527 , n279 , n3595 );
    xor g2220 ( n2939 , n2232 , n1797 );
    xnor g2221 ( n3253 , n2654 , n712 );
    or g2222 ( n1471 , n2054 , n1961 );
    xnor g2223 ( n1114 , n2734 , n2984 );
    nor g2224 ( n92 , n2105 , n566 );
    nor g2225 ( n2949 , n1370 , n2602 );
    or g2226 ( n3283 , n1324 , n2283 );
    or g2227 ( n3260 , n2578 , n1648 );
    xnor g2228 ( n628 , n2531 , n1206 );
    or g2229 ( n2100 , n174 , n158 );
    xnor g2230 ( n76 , n1365 , n3524 );
    xnor g2231 ( n3224 , n1722 , n13 );
    or g2232 ( n344 , n1757 , n1501 );
    and g2233 ( n19 , n805 , n3525 );
    not g2234 ( n2242 , n772 );
    or g2235 ( n2144 , n305 , n1810 );
    and g2236 ( n1843 , n307 , n3829 );
    and g2237 ( n1999 , n1471 , n3685 );
    not g2238 ( n1622 , n1204 );
    not g2239 ( n2796 , n2773 );
    or g2240 ( n3171 , n115 , n2373 );
    not g2241 ( n2907 , n2727 );
    xnor g2242 ( n2434 , n2208 , n534 );
    xnor g2243 ( n1658 , n1275 , n1538 );
    xnor g2244 ( n3775 , n1712 , n3539 );
    nor g2245 ( n3884 , n2460 , n2772 );
    or g2246 ( n952 , n913 , n1856 );
    not g2247 ( n1995 , n864 );
    not g2248 ( n370 , n1820 );
    or g2249 ( n436 , n2543 , n1502 );
    or g2250 ( n681 , n3599 , n917 );
    or g2251 ( n1908 , n1121 , n3263 );
    xnor g2252 ( n152 , n2071 , n1161 );
    not g2253 ( n2604 , n2112 );
    or g2254 ( n2076 , n748 , n3834 );
    or g2255 ( n2047 , n694 , n1859 );
    not g2256 ( n2870 , n178 );
    xnor g2257 ( n2865 , n1442 , n3010 );
    and g2258 ( n1032 , n1710 , n1088 );
    and g2259 ( n2905 , n3639 , n1919 );
    or g2260 ( n443 , n2102 , n3373 );
    or g2261 ( n2285 , n2410 , n1970 );
    and g2262 ( n2455 , n2019 , n540 );
    and g2263 ( n672 , n3245 , n1300 );
    or g2264 ( n2717 , n3458 , n401 );
    and g2265 ( n2070 , n3078 , n1349 );
    and g2266 ( n619 , n669 , n3057 );
    or g2267 ( n2462 , n3674 , n627 );
    not g2268 ( n675 , n494 );
    or g2269 ( n1801 , n980 , n327 );
    or g2270 ( n3006 , n2324 , n2322 );
    and g2271 ( n268 , n945 , n3849 );
    or g2272 ( n2483 , n2257 , n2637 );
    not g2273 ( n2677 , n1240 );
    xnor g2274 ( n666 , n3882 , n921 );
    or g2275 ( n389 , n148 , n3782 );
    and g2276 ( n3502 , n770 , n1273 );
    not g2277 ( n1593 , n3891 );
    xnor g2278 ( n902 , n1031 , n3003 );
    not g2279 ( n3557 , n2772 );
    xnor g2280 ( n3029 , n1012 , n3334 );
    xnor g2281 ( n643 , n516 , n1101 );
    or g2282 ( n2556 , n1958 , n2506 );
    or g2283 ( n3084 , n1808 , n3022 );
    nor g2284 ( n1976 , n2527 , n2531 );
    xnor g2285 ( n728 , n1879 , n1468 );
    or g2286 ( n1112 , n2124 , n3277 );
    xnor g2287 ( n943 , n2554 , n2925 );
    xnor g2288 ( n256 , n801 , n3041 );
    or g2289 ( n2255 , n913 , n973 );
    xnor g2290 ( n2045 , n2484 , n1203 );
    not g2291 ( n2030 , n891 );
    not g2292 ( n2899 , n3708 );
    xnor g2293 ( n2559 , n399 , n3482 );
    or g2294 ( n400 , n906 , n103 );
    not g2295 ( n1071 , n1594 );
    and g2296 ( n406 , n2339 , n3766 );
    or g2297 ( n3623 , n66 , n726 );
    xnor g2298 ( n3606 , n2881 , n3467 );
    xnor g2299 ( n3407 , n2008 , n3320 );
    not g2300 ( n3189 , n835 );
    or g2301 ( n3543 , n590 , n486 );
    or g2302 ( n718 , n302 , n521 );
    xnor g2303 ( n2519 , n769 , n3678 );
    and g2304 ( n3178 , n2584 , n1457 );
    not g2305 ( n1934 , n1640 );
    xnor g2306 ( n32 , n3128 , n2660 );
    not g2307 ( n791 , n2324 );
    xnor g2308 ( n614 , n3360 , n360 );
    and g2309 ( n2670 , n1741 , n1132 );
    not g2310 ( n2233 , n1404 );
    and g2311 ( n1850 , n1041 , n3282 );
    not g2312 ( n934 , n1989 );
    xnor g2313 ( n192 , n3470 , n2356 );
    and g2314 ( n237 , n2971 , n1982 );
    or g2315 ( n1045 , n3810 , n3527 );
    not g2316 ( n3783 , n2757 );
    not g2317 ( n804 , n56 );
    not g2318 ( n3612 , n2912 );
    or g2319 ( n1681 , n2979 , n626 );
    and g2320 ( n860 , n2903 , n3428 );
    or g2321 ( n1687 , n889 , n1483 );
    not g2322 ( n118 , n1103 );
    and g2323 ( n3270 , n1587 , n443 );
    or g2324 ( n2517 , n2541 , n3356 );
    xnor g2325 ( n1454 , n1956 , n3254 );
    and g2326 ( n3745 , n350 , n2782 );
    or g2327 ( n1601 , n3091 , n3189 );
    and g2328 ( n136 , n3773 , n2848 );
    or g2329 ( n144 , n2936 , n1087 );
    or g2330 ( n2847 , n848 , n2672 );
    xnor g2331 ( n3603 , n3047 , n2670 );
    not g2332 ( n3719 , n2073 );
    xnor g2333 ( n2263 , n3398 , n1424 );
    xnor g2334 ( n1363 , n2629 , n603 );
    or g2335 ( n1576 , n1142 , n1339 );
    and g2336 ( n1586 , n1063 , n2606 );
    not g2337 ( n819 , n1541 );
    not g2338 ( n1094 , n1983 );
    and g2339 ( n2394 , n520 , n212 );
    xnor g2340 ( n3025 , n1308 , n1257 );
    or g2341 ( n3857 , n1968 , n1208 );
    or g2342 ( n2067 , n2087 , n1954 );
    xnor g2343 ( n2422 , n3066 , n1699 );
    not g2344 ( n3746 , n274 );
    not g2345 ( n221 , n1507 );
    xnor g2346 ( n974 , n3803 , n3284 );
    and g2347 ( n1698 , n3867 , n491 );
    nor g2348 ( n1607 , n1215 , n1588 );
    and g2349 ( n3122 , n308 , n794 );
    xnor g2350 ( n3691 , n1643 , n692 );
    or g2351 ( n1532 , n2003 , n2586 );
    and g2352 ( n3359 , n824 , n2371 );
    nor g2353 ( n3808 , n74 , n1784 );
    nor g2354 ( n1835 , n2876 , n969 );
    not g2355 ( n3527 , n940 );
    not g2356 ( n186 , n1027 );
    xnor g2357 ( n2558 , n524 , n3351 );
    or g2358 ( n661 , n66 , n1785 );
    xor g2359 ( n1883 , n969 , n2832 );
    and g2360 ( n3108 , n546 , n3729 );
    not g2361 ( n3315 , n1027 );
    not g2362 ( n6 , n1280 );
    xnor g2363 ( n717 , n774 , n1986 );
    nor g2364 ( n453 , n2260 , n369 );
    xnor g2365 ( n461 , n1109 , n3086 );
    or g2366 ( n1185 , n1327 , n3746 );
    or g2367 ( n1241 , n187 , n3574 );
    xnor g2368 ( n3514 , n2277 , n464 );
    or g2369 ( n3377 , n1928 , n2628 );
    xnor g2370 ( n1993 , n2309 , n2810 );
    nor g2371 ( n276 , n3857 , n2902 );
    not g2372 ( n3153 , n1404 );
    xnor g2373 ( n2360 , n2982 , n2310 );
    nor g2374 ( n836 , n276 , n254 );
    not g2375 ( n3644 , n2126 );
    or g2376 ( n340 , n1364 , n3728 );
    or g2377 ( n3713 , n3191 , n2801 );
    and g2378 ( n2680 , n887 , n2556 );
    or g2379 ( n1770 , n2005 , n1856 );
    nor g2380 ( n3347 , n962 , n3096 );
    nor g2381 ( n3581 , n1722 , n426 );
    xnor g2382 ( n2384 , n2105 , n773 );
    not g2383 ( n2852 , n1761 );
    and g2384 ( n3039 , n2479 , n2147 );
    xnor g2385 ( n2303 , n1859 , n1278 );
    xnor g2386 ( n1445 , n3240 , n255 );
    or g2387 ( n1701 , n3132 , n1563 );
    and g2388 ( n3344 , n3683 , n207 );
    not g2389 ( n2518 , n2065 );
    and g2390 ( n2932 , n2778 , n1081 );
    and g2391 ( n1476 , n2341 , n1599 );
    nor g2392 ( n2335 , n377 , n2762 );
    not g2393 ( n1084 , n955 );
    and g2394 ( n1134 , n506 , n2849 );
    and g2395 ( n3058 , n2380 , n3768 );
    not g2396 ( n1548 , n3272 );
    not g2397 ( n3637 , n2912 );
    or g2398 ( n1692 , n3675 , n1781 );
    xnor g2399 ( n2845 , n9 , n1015 );
    or g2400 ( n2543 , n3630 , n434 );
    xnor g2401 ( n3254 , n694 , n2303 );
    and g2402 ( n1831 , n2418 , n3036 );
    or g2403 ( n2772 , n892 , n3355 );
    and g2404 ( n2316 , n1851 , n1407 );
    xnor g2405 ( n1767 , n141 , n2847 );
    xnor g2406 ( n2916 , n757 , n1462 );
    and g2407 ( n1042 , n315 , n379 );
    xnor g2408 ( n3749 , n3729 , n3850 );
    not g2409 ( n2748 , n3077 );
    and g2410 ( n1619 , n60 , n3128 );
    xnor g2411 ( n759 , n3518 , n1115 );
    not g2412 ( n2132 , n2811 );
    xnor g2413 ( n547 , n2687 , n3563 );
    nor g2414 ( n1252 , n867 , n600 );
    and g2415 ( n1717 , n770 , n422 );
    or g2416 ( n439 , n1213 , n136 );
    or g2417 ( n475 , n2177 , n204 );
    or g2418 ( n189 , n2650 , n3104 );
    and g2419 ( n1668 , n778 , n3567 );
    not g2420 ( n1076 , n1541 );
    xnor g2421 ( n1988 , n720 , n418 );
    and g2422 ( n1281 , n1087 , n2936 );
    xnor g2423 ( n2267 , n282 , n518 );
    or g2424 ( n847 , n135 , n3625 );
    xnor g2425 ( n1342 , n1777 , n689 );
    or g2426 ( n1165 , n2194 , n3396 );
    xnor g2427 ( n1736 , n735 , n2150 );
    and g2428 ( n1278 , n1447 , n2148 );
    or g2429 ( n644 , n3410 , n3326 );
    or g2430 ( n2069 , n1809 , n3747 );
    and g2431 ( n2643 , n655 , n1516 );
    and g2432 ( n1933 , n1089 , n2674 );
    or g2433 ( n2328 , n138 , n3055 );
    xnor g2434 ( n2248 , n1490 , n3039 );
    xor g2435 ( n3392 , n3421 , n2520 );
    or g2436 ( n1932 , n2988 , n2060 );
    or g2437 ( n1526 , n2677 , n2511 );
    xnor g2438 ( n2120 , n2153 , n3194 );
    not g2439 ( n627 , n274 );
    and g2440 ( n3284 , n1366 , n3203 );
    xnor g2441 ( n2897 , n1544 , n1145 );
    or g2442 ( n2502 , n934 , n3718 );
    xnor g2443 ( n1986 , n2610 , n3840 );
    xnor g2444 ( n2060 , n2923 , n2571 );
    nor g2445 ( n101 , n1873 , n226 );
    or g2446 ( n408 , n1353 , n936 );
    xnor g2447 ( n3714 , n2113 , n2485 );
    or g2448 ( n830 , n2859 , n1552 );
    xnor g2449 ( n2490 , n1571 , n3457 );
    or g2450 ( n3676 , n3790 , n2961 );
    or g2451 ( n3167 , n588 , n3455 );
    or g2452 ( n923 , n3091 , n1981 );
    xor g2453 ( n1695 , n2065 , n1543 );
    xnor g2454 ( n3518 , n3413 , n3635 );
    and g2455 ( n50 , n1583 , n2844 );
    or g2456 ( n2833 , n1112 , n2552 );
    or g2457 ( n2048 , n1560 , n918 );
    and g2458 ( n481 , n891 , n1507 );
    xnor g2459 ( n1776 , n1251 , n575 );
    xnor g2460 ( n2083 , n1324 , n1763 );
    not g2461 ( n2095 , n3510 );
    or g2462 ( n765 , n1014 , n1718 );
    and g2463 ( n3511 , n2403 , n1341 );
    xnor g2464 ( n3383 , n2201 , n146 );
    or g2465 ( n1479 , n437 , n2028 );
    xor g2466 ( n2883 , n1309 , n3015 );
    or g2467 ( n2782 , n2746 , n3720 );
    or g2468 ( n1826 , n3796 , n1249 );
    not g2469 ( n1754 , n1103 );
    or g2470 ( n2103 , n3010 , n1963 );
    or g2471 ( n1152 , n336 , n2747 );
    and g2472 ( n1869 , n421 , n97 );
    nor g2473 ( n1386 , n1484 , n2435 );
    xnor g2474 ( n447 , n2642 , n1521 );
    not g2475 ( n1557 , n1367 );
    not g2476 ( n912 , n3690 );
    xnor g2477 ( n2464 , n719 , n3201 );
    xnor g2478 ( n3332 , n2873 , n3836 );
    or g2479 ( n467 , n2191 , n804 );
    or g2480 ( n938 , n623 , n3125 );
    not g2481 ( n1968 , n2567 );
    xor g2482 ( n1949 , n2735 , n3577 );
    or g2483 ( n3782 , n589 , n1499 );
    xnor g2484 ( n1391 , n2458 , n2776 );
    or g2485 ( n1665 , n1077 , n154 );
    not g2486 ( n2658 , n1782 );
    xnor g2487 ( n1184 , n3382 , n3323 );
    xnor g2488 ( n2841 , n2919 , n2045 );
    or g2489 ( n3697 , n1113 , n764 );
    or g2490 ( n879 , n3634 , n3576 );
    and g2491 ( n2877 , n1109 , n3490 );
    not g2492 ( n3834 , n891 );
    and g2493 ( n2636 , n1005 , n3864 );
    not g2494 ( n2672 , n3898 );
    xnor g2495 ( n3194 , n2990 , n2880 );
    or g2496 ( n2237 , n1369 , n1590 );
    xnor g2497 ( n1504 , n2192 , n2219 );
    xnor g2498 ( n3680 , n390 , n2620 );
    or g2499 ( n3744 , n509 , n3300 );
    not g2500 ( n483 , n670 );
    and g2501 ( n601 , n1744 , n1605 );
    or g2502 ( n760 , n2886 , n862 );
    or g2503 ( n2884 , n1198 , n370 );
    xnor g2504 ( n615 , n87 , n521 );
    not g2505 ( n818 , n88 );
    nor g2506 ( n1175 , n3811 , n1528 );
    or g2507 ( n3614 , n1062 , n624 );
    not g2508 ( n3862 , n2324 );
    xnor g2509 ( n632 , n3653 , n105 );
    xnor g2510 ( n1425 , n1321 , n628 );
    xnor g2511 ( n307 , n538 , n256 );
    not g2512 ( n2183 , n2656 );
    xnor g2513 ( n1356 , n3766 , n1158 );
    xnor g2514 ( n2970 , n1512 , n489 );
    or g2515 ( n357 , n73 , n559 );
    nor g2516 ( n2493 , n3199 , n638 );
    and g2517 ( n2933 , n1096 , n501 );
    or g2518 ( n3522 , n3319 , n2794 );
    and g2519 ( n2409 , n915 , n2855 );
    xnor g2520 ( n2773 , n3519 , n1767 );
    or g2521 ( n412 , n2530 , n725 );
    xnor g2522 ( n3218 , n1345 , n2263 );
    or g2523 ( n2553 , n2378 , n3020 );
    and g2524 ( n659 , n2211 , n3653 );
    nor g2525 ( n3666 , n540 , n2019 );
    nor g2526 ( n213 , n2134 , n2408 );
    not g2527 ( n1683 , n835 );
    or g2528 ( n2119 , n48 , n857 );
    or g2529 ( n3387 , n285 , n3157 );
    and g2530 ( n2634 , n1376 , n3711 );
    or g2531 ( n2221 , n197 , n3694 );
    not g2532 ( n2992 , n107 );
    not g2533 ( n2049 , n1808 );
    xnor g2534 ( n2482 , n1824 , n2719 );
    xor g2535 ( n730 , n134 , n2765 );
    not g2536 ( n3370 , n387 );
    or g2537 ( n2917 , n1397 , n402 );
    or g2538 ( n40 , n1253 , n1032 );
    xnor g2539 ( n414 , n3308 , n3392 );
    and g2540 ( n3700 , n1082 , n384 );
    and g2541 ( n318 , n3386 , n647 );
    not g2542 ( n1962 , n2966 );
    and g2543 ( n2320 , n1642 , n345 );
    and g2544 ( n2586 , n3154 , n2467 );
    xnor g2545 ( n3495 , n1991 , n1154 );
    or g2546 ( n2564 , n3082 , n1080 );
    and g2547 ( n3761 , n1274 , n218 );
    not g2548 ( n3446 , n1234 );
    and g2549 ( n2308 , n2800 , n41 );
    xnor g2550 ( n623 , n2959 , n2797 );
    and g2551 ( n1676 , n2309 , n970 );
    nor g2552 ( n3641 , n2893 , n2084 );
    and g2553 ( n3223 , n2923 , n2836 );
    xnor g2554 ( n1818 , n2428 , n65 );
    or g2555 ( n1059 , n1569 , n1208 );
    xnor g2556 ( n429 , n1501 , n3869 );
    or g2557 ( n2993 , n2652 , n2922 );
    not g2558 ( n2808 , n504 );
    and g2559 ( n1784 , n3135 , n1023 );
    or g2560 ( n1615 , n737 , n3489 );
    and g2561 ( n1320 , n3593 , n2183 );
    xor g2562 ( n813 , n1554 , n2893 );
    or g2563 ( n3363 , n563 , n947 );
    xnor g2564 ( n3314 , n1041 , n2361 );
    xnor g2565 ( n2619 , n949 , n2693 );
    or g2566 ( n832 , n1012 , n3840 );
    and g2567 ( n1167 , n51 , n2835 );
    xnor g2568 ( n541 , n1456 , n974 );
    and g2569 ( n3656 , n3178 , n3701 );
    xnor g2570 ( n2007 , n1622 , n384 );
    or g2571 ( n3491 , n1512 , n3267 );
    and g2572 ( n1201 , n2934 , n2920 );
    not g2573 ( n2668 , n3038 );
    and g2574 ( n2107 , n2069 , n1458 );
    not g2575 ( n2511 , n772 );
    and g2576 ( n2340 , n3677 , n2884 );
    not g2577 ( n1443 , n3536 );
    or g2578 ( n1805 , n1099 , n1410 );
    xnor g2579 ( n2676 , n546 , n3749 );
    nor g2580 ( n3876 , n925 , n842 );
    not g2581 ( n740 , n1323 );
    or g2582 ( n2475 , n3354 , n1421 );
    or g2583 ( n2563 , n3881 , n261 );
    and g2584 ( n3655 , n3308 , n3421 );
    xnor g2585 ( n3516 , n2821 , n1519 );
    or g2586 ( n3628 , n599 , n606 );
    or g2587 ( n234 , n3826 , n2675 );
    or g2588 ( n2136 , n229 , n3180 );
    and g2589 ( n2105 , n663 , n2585 );
    xor g2590 ( n165 , n395 , n2368 );
    or g2591 ( n3386 , n257 , n2107 );
    and g2592 ( n289 , n2042 , n425 );
    or g2593 ( n600 , n2347 , n3409 );
    and g2594 ( n353 , n427 , n1733 );
    xnor g2595 ( n2669 , n3167 , n1574 );
    or g2596 ( n688 , n430 , n818 );
    and g2597 ( n386 , n3521 , n375 );
    or g2598 ( n2843 , n159 , n3873 );
    xnor g2599 ( n1043 , n1506 , n3859 );
    and g2600 ( n1514 , n3445 , n3353 );
    not g2601 ( n2824 , n2871 );
    or g2602 ( n3784 , n2324 , n2862 );
    and g2603 ( n2555 , n3085 , n1943 );
    not g2604 ( n3661 , n3819 );
    or g2605 ( n203 , n1922 , n1042 );
    and g2606 ( n115 , n205 , n1834 );
    or g2607 ( n379 , n2414 , n2462 );
    xnor g2608 ( n1839 , n570 , n1074 );
    and g2609 ( n3675 , n1035 , n535 );
    or g2610 ( n2470 , n117 , n2890 );
    not g2611 ( n1546 , n1950 );
    and g2612 ( n3717 , n972 , n265 );
    and g2613 ( n1567 , n808 , n1490 );
    and g2614 ( n3551 , n3225 , n332 );
    nor g2615 ( n3503 , n2841 , n3780 );
    not g2616 ( n1216 , n537 );
    not g2617 ( n124 , n2523 );
    xnor g2618 ( n1380 , n280 , n3560 );
    and g2619 ( n2268 , n2267 , n3613 );
    and g2620 ( n2769 , n739 , n1067 );
    not g2621 ( n1691 , n547 );
    not g2622 ( n466 , n1156 );
    xnor g2623 ( n3422 , n3370 , n3782 );
    and g2624 ( n3665 , n1394 , n1863 );
    not g2625 ( n3827 , n3805 );
    or g2626 ( n1580 , n461 , n2070 );
    and g2627 ( n117 , n2553 , n2535 );
    not g2628 ( n3796 , n3359 );
    not g2629 ( n3590 , n1898 );
    and g2630 ( n2290 , n2397 , n846 );
    and g2631 ( n302 , n1022 , n87 );
    not g2632 ( n3622 , n2572 );
    xnor g2633 ( n2174 , n942 , n1815 );
    xnor g2634 ( n1424 , n2975 , n964 );
    or g2635 ( n795 , n3195 , n1426 );
    or g2636 ( n3382 , n483 , n1333 );
    or g2637 ( n1003 , n1727 , n2095 );
    and g2638 ( n3880 , n865 , n607 );
    or g2639 ( n3334 , n1455 , n3893 );
    and g2640 ( n1617 , n771 , n3087 );
    or g2641 ( n438 , n1641 , n1728 );
    not g2642 ( n1051 , n335 );
    and g2643 ( n1019 , n1460 , n3664 );
    and g2644 ( n1952 , n690 , n2502 );
    not g2645 ( n925 , n1363 );
    xnor g2646 ( n1143 , n2911 , n2480 );
    xnor g2647 ( n570 , n2121 , n109 );
    or g2648 ( n109 , n2775 , n3754 );
    not g2649 ( n3659 , n422 );
    xor g2650 ( n79 , n381 , n911 );
    or g2651 ( n3818 , n1696 , n2308 );
    or g2652 ( n2289 , n952 , n2645 );
    or g2653 ( n1530 , n3422 , n1956 );
    and g2654 ( n2880 , n2342 , n1139 );
    xor g2655 ( n1176 , n2440 , n303 );
    or g2656 ( n3598 , n3222 , n2580 );
    or g2657 ( n3886 , n729 , n860 );
    not g2658 ( n2094 , n2031 );
    and g2659 ( n1961 , n1965 , n3143 );
    or g2660 ( n2626 , n2870 , n995 );
    or g2661 ( n1415 , n1075 , n1411 );
    xnor g2662 ( n2153 , n1744 , n656 );
    or g2663 ( n2080 , n1428 , n3019 );
    or g2664 ( n3354 , n216 , n3732 );
    or g2665 ( n2009 , n598 , n2478 );
    xnor g2666 ( n3136 , n2773 , n1183 );
    xnor g2667 ( n2380 , n952 , n1343 );
    not g2668 ( n3589 , n491 );
    xnor g2669 ( n3696 , n1594 , n3338 );
    xor g2670 ( n1243 , n1513 , n2905 );
    not g2671 ( n1321 , n2000 );
    not g2672 ( n1484 , n2946 );
    not g2673 ( n2860 , n2258 );
    or g2674 ( n1158 , n1822 , n1683 );
    not g2675 ( n2569 , n1231 );
    xnor g2676 ( n899 , n3785 , n1135 );
    not g2677 ( n1783 , n1775 );
    or g2678 ( n1349 , n1415 , n2915 );
    xnor g2679 ( n834 , n2339 , n1356 );
    or g2680 ( n2032 , n2166 , n3011 );
    xnor g2681 ( n1144 , n2230 , n890 );
    not g2682 ( n441 , n642 );
    or g2683 ( n942 , n3788 , n368 );
    xnor g2684 ( n271 , n2979 , n567 );
    xor g2685 ( n2839 , n644 , n680 );
    or g2686 ( n1265 , n3783 , n296 );
    not g2687 ( n2709 , n2769 );
    xnor g2688 ( n1227 , n3393 , n1670 );
    xnor g2689 ( n1940 , n2460 , n3006 );
    or g2690 ( n1600 , n2338 , n1664 );
    and g2691 ( n3052 , n2632 , n1554 );
    xnor g2692 ( n1704 , n3235 , n2053 );
    nor g2693 ( n3132 , n2132 , n2374 );
    nor g2694 ( n3281 , n3804 , n1252 );
    or g2695 ( n2545 , n1137 , n333 );
    and g2696 ( n1427 , n3342 , n2224 );
    xnor g2697 ( n479 , n2624 , n1582 );
    and g2698 ( n1563 , n2692 , n2216 );
    or g2699 ( n3737 , n346 , n1788 );
    or g2700 ( n2649 , n1022 , n87 );
    or g2701 ( n612 , n1275 , n1606 );
    xor g2702 ( n2832 , n2876 , n1608 );
    xnor g2703 ( n1889 , n3288 , n2842 );
    nor g2704 ( n2291 , n410 , n152 );
    xnor g2705 ( n744 , n2345 , n2029 );
    or g2706 ( n2937 , n2324 , n2261 );
    not g2707 ( n3753 , n2523 );
    or g2708 ( n3718 , n3005 , n2271 );
    xnor g2709 ( n2858 , n1248 , n490 );
    and g2710 ( n3489 , n2485 , n3716 );
    and g2711 ( n2497 , n1472 , n203 );
    not g2712 ( n1370 , n661 );
    and g2713 ( n499 , n428 , n3848 );
    not g2714 ( n2128 , n2687 );
    or g2715 ( n3777 , n3518 , n1418 );
    and g2716 ( n3012 , n338 , n71 );
    not g2717 ( n2334 , n2830 );
    or g2718 ( n3463 , n3869 , n3102 );
    or g2719 ( n3130 , n3172 , n2926 );
    or g2720 ( n551 , n1846 , n27 );
    or g2721 ( n833 , n2429 , n104 );
    and g2722 ( n1611 , n3519 , n141 );
    not g2723 ( n169 , n2744 );
    or g2724 ( n1522 , n3876 , n1732 );
    nor g2725 ( n3368 , n2036 , n538 );
    and g2726 ( n843 , n2153 , n2990 );
    not g2727 ( n2061 , n1066 );
    xnor g2728 ( n1654 , n1181 , n1469 );
    or g2729 ( n2139 , n3181 , n3451 );
    and g2730 ( n376 , n2177 , n204 );
    xnor g2731 ( n2114 , n3105 , n1200 );
    nor g2732 ( n1620 , n2239 , n1100 );
    xnor g2733 ( n3454 , n2193 , n761 );
    xnor g2734 ( n1947 , n438 , n93 );
    not g2735 ( n2321 , n768 );
    not g2736 ( n1760 , n3255 );
    or g2737 ( n2746 , n3622 , n2577 );
    not g2738 ( n3051 , n2646 );
    not g2739 ( n920 , n2842 );
    not g2740 ( n1178 , n1446 );
    not g2741 ( n3810 , n1367 );
    xnor g2742 ( n80 , n295 , n1357 );
    or g2743 ( n229 , n2288 , n2694 );
    not g2744 ( n3117 , n2294 );
    or g2745 ( n3060 , n124 , n2095 );
    not g2746 ( n2478 , n2744 );
    or g2747 ( n2629 , n1162 , n2607 );
    xnor g2748 ( n1417 , n3720 , n3182 );
    not g2749 ( n3309 , n3340 );
    xnor g2750 ( n455 , n1211 , n2360 );
    not g2751 ( n1573 , n493 );
    not g2752 ( n1126 , n3566 );
    and g2753 ( n2736 , n2483 , n3642 );
    nor g2754 ( n451 , n2871 , n3495 );
    not g2755 ( n3575 , n2714 );
    and g2756 ( n1543 , n2760 , n1273 );
    not g2757 ( n599 , n944 );
    and g2758 ( n519 , n1711 , n2126 );
    and g2759 ( n1810 , n3471 , n389 );
    xnor g2760 ( n1806 , n73 , n559 );
    xor g2761 ( n3414 , n547 , n3878 );
    not g2762 ( n3893 , n2514 );
    xnor g2763 ( n904 , n780 , n1693 );
    xnor g2764 ( n2417 , n1690 , n2273 );
    or g2765 ( n2339 , n3719 , n20 );
    xnor g2766 ( n966 , n1684 , n633 );
    or g2767 ( n2065 , n466 , n1064 );
    and g2768 ( n1020 , n585 , n3621 );
    and g2769 ( n1174 , n2801 , n3298 );
    not g2770 ( n284 , n794 );
    and g2771 ( n3388 , n163 , n2962 );
    and g2772 ( n2318 , n2060 , n2988 );
    and g2773 ( n3546 , n2356 , n3470 );
    nor g2774 ( n1849 , n3730 , n3397 );
    xnor g2775 ( n2835 , n1847 , n1408 );
    and g2776 ( n1061 , n975 , n500 );
    and g2777 ( n867 , n3190 , n3862 );
    not g2778 ( n949 , n1802 );
    or g2779 ( n3275 , n2016 , n2672 );
    or g2780 ( n325 , n120 , n3885 );
    and g2781 ( n1260 , n600 , n867 );
    xnor g2782 ( n1945 , n2551 , n3101 );
    xnor g2783 ( n86 , n3701 , n3459 );
    and g2784 ( n1186 , n1313 , n407 );
    or g2785 ( n3242 , n3012 , n1316 );
    or g2786 ( n57 , n2353 , n2340 );
    and g2787 ( n433 , n3090 , n3530 );
    xnor g2788 ( n3294 , n62 , n3021 );
    xnor g2789 ( n2330 , n3025 , n1114 );
    xnor g2790 ( n1150 , n1848 , n2816 );
    and g2791 ( n3061 , n426 , n1722 );
    xnor g2792 ( n2764 , n491 , n1918 );
    not g2793 ( n3356 , n274 );
    xnor g2794 ( n3267 , n2177 , n1926 );
    not g2795 ( n3226 , n1582 );
    and g2796 ( n2637 , n2503 , n2289 );
    or g2797 ( n2471 , n1601 , n3497 );
    and g2798 ( n2173 , n1024 , n510 );
    xor g2799 ( n1182 , n3888 , n3765 );
    or g2800 ( n1296 , n2140 , n1985 );
    xnor g2801 ( n146 , n1294 , n1319 );
    and g2802 ( n2733 , n810 , n1120 );
    xnor g2803 ( n1632 , n3852 , n3453 );
    xnor g2804 ( n539 , n3718 , n1383 );
    not g2805 ( n1731 , n622 );
    xnor g2806 ( n1099 , n978 , n416 );
    nor g2807 ( n3378 , n1212 , n2157 );
    nor g2808 ( n2036 , n1577 , n1910 );
    or g2809 ( n976 , n290 , n3074 );
    and g2810 ( n803 , n1775 , n1280 );
    or g2811 ( n2731 , n1198 , n2783 );
    not g2812 ( n1794 , n3649 );
    not g2813 ( n2191 , n2727 );
    not g2814 ( n1220 , n3014 );
    and g2815 ( n575 , n3381 , n3337 );
    not g2816 ( n1259 , n88 );
    or g2817 ( n1068 , n2162 , n2161 );
    not g2818 ( n3200 , n3384 );
    not g2819 ( n515 , n3444 );
    or g2820 ( n1834 , n2279 , n3628 );
    xnor g2821 ( n322 , n2632 , n813 );
    not g2822 ( n3716 , n2117 );
    or g2823 ( n2043 , n3629 , n2754 );
    or g2824 ( n831 , n3674 , n488 );
    or g2825 ( n1376 , n1959 , n2651 );
    not g2826 ( n3458 , n181 );
    not g2827 ( n2311 , n3481 );
    nor g2828 ( n1660 , n3717 , n1306 );
    or g2829 ( n3308 , n3880 , n2534 );
    or g2830 ( n1407 , n3477 , n75 );
    and g2831 ( n3456 , n1195 , n2779 );
    not g2832 ( n291 , n111 );
    xor g2833 ( n3044 , n1268 , n958 );
    and g2834 ( n715 , n3201 , n719 );
    or g2835 ( n3050 , n3345 , n2146 );
    or g2836 ( n3549 , n70 , n861 );
    or g2837 ( n2848 , n2066 , n3867 );
    xnor g2838 ( n3839 , n1045 , n899 );
    and g2839 ( n775 , n3096 , n962 );
    or g2840 ( n3840 , n1393 , n1180 );
    and g2841 ( n1309 , n1805 , n1304 );
    and g2842 ( n1074 , n2006 , n1713 );
    or g2843 ( n2333 , n1221 , n3531 );
    or g2844 ( n790 , n1107 , n3233 );
    not g2845 ( n1466 , n2640 );
    or g2846 ( n3228 , n2587 , n2108 );
    not g2847 ( n469 , n2724 );
    xnor g2848 ( n2581 , n3232 , n3429 );
    or g2849 ( n3664 , n53 , n983 );
    or g2850 ( n3626 , n573 , n1726 );
    not g2851 ( n273 , n2110 );
    and g2852 ( n2155 , n3463 , n344 );
    and g2853 ( n416 , n3318 , n591 );
    and g2854 ( n2450 , n3217 , n1317 );
    not g2855 ( n1355 , n1793 );
    and g2856 ( n861 , n1110 , n309 );
    and g2857 ( n1537 , n1946 , n2981 );
    not g2858 ( n2610 , n2748 );
    or g2859 ( n3523 , n1703 , n1009 );
    nor g2860 ( n2364 , n291 , n3662 );
    or g2861 ( n1438 , n3897 , n1644 );
    or g2862 ( n3258 , n1072 , n2983 );
    not g2863 ( n3582 , n1318 );
    or g2864 ( n1442 , n3809 , n488 );
    xnor g2865 ( n823 , n994 , n1344 );
    or g2866 ( n870 , n2255 , n3544 );
    not g2867 ( n3298 , n3315 );
    or g2868 ( n3686 , n2859 , n2592 );
    not g2869 ( n3596 , n308 );
    and g2870 ( n931 , n3538 , n2500 );
    not g2871 ( n3396 , n642 );
    xnor g2872 ( n2381 , n3438 , n2628 );
    xnor g2873 ( n2742 , n553 , n1553 );
    xnor g2874 ( n2468 , n1172 , n3680 );
    not g2875 ( n2126 , n2659 );
    or g2876 ( n3264 , n1299 , n2114 );
    or g2877 ( n3467 , n1077 , n2918 );
    not g2878 ( n1331 , n1952 );
    xnor g2879 ( n2041 , n1439 , n3868 );
    not g2880 ( n2260 , n404 );
    xnor g2881 ( n2622 , n571 , n241 );
    or g2882 ( n224 , n3059 , n3334 );
    and g2883 ( n995 , n2969 , n3242 );
    or g2884 ( n557 , n3768 , n2380 );
    not g2885 ( n527 , n1025 );
    nor g2886 ( n2078 , n2752 , n1917 );
    xnor g2887 ( n2708 , n3291 , n3800 );
    or g2888 ( n2730 , n577 , n2229 );
    xor g2889 ( n100 , n2266 , n2939 );
    xnor g2890 ( n1419 , n2646 , n1743 );
    xnor g2891 ( n3174 , n1677 , n747 );
    not g2892 ( n3809 , n3774 );
    not g2893 ( n3 , n2724 );
    xnor g2894 ( n1343 , n2645 , n3787 );
    not g2895 ( n3055 , n3444 );
    not g2896 ( n598 , n944 );
    xnor g2897 ( n761 , n2874 , n3418 );
    and g2898 ( n3040 , n1537 , n1169 );
    and g2899 ( n1656 , n1823 , n1193 );
    not g2900 ( n2459 , n1577 );
    and g2901 ( n3723 , n330 , n395 );
    xnor g2902 ( n97 , n1837 , n1750 );
    xnor g2903 ( n3847 , n482 , n3501 );
    not g2904 ( n3674 , n220 );
    xnor g2905 ( n618 , n2576 , n2991 );
    and g2906 ( n3752 , n2673 , n822 );
    xnor g2907 ( n788 , n2314 , n1196 );
    xnor g2908 ( n2842 , n1833 , n686 );
    not g2909 ( n2027 , n1020 );
    or g2910 ( n2354 , n2324 , n2857 );
    xnor g2911 ( n3426 , n1791 , n3600 );
    not g2912 ( n2696 , n2463 );
    xnor g2913 ( n484 , n815 , n2603 );
    not g2914 ( n2003 , n1255 );
    or g2915 ( n2108 , n3095 , n800 );
    or g2916 ( n1939 , n2008 , n1105 );
    xnor g2917 ( n1511 , n2709 , n463 );
    or g2918 ( n3135 , n2241 , n3605 );
    or g2919 ( n1919 , n1251 , n575 );
    and g2920 ( n1845 , n1062 , n624 );
    or g2921 ( n3867 , n3163 , n1 );
    and g2922 ( n3492 , n923 , n83 );
    and g2923 ( n3722 , n1456 , n3803 );
    or g2924 ( n990 , n2064 , n763 );
    xnor g2925 ( n2446 , n2279 , n2035 );
    and g2926 ( n3013 , n1019 , n3162 );
    and g2927 ( n3014 , n1596 , n3352 );
    not g2928 ( n1960 , n3321 );
    nor g2929 ( n3156 , n1342 , n1134 );
    or g2930 ( n1441 , n3575 , n479 );
    and g2931 ( n1080 , n1819 , n1768 );
    or g2932 ( n634 , n3254 , n269 );
    xnor g2933 ( n3101 , n1880 , n239 );
    or g2934 ( n3288 , n3789 , n1716 );
    or g2935 ( n3601 , n1489 , n1392 );
    not g2936 ( n430 , n493 );
    and g2937 ( n30 , n837 , n1029 );
    not g2938 ( n2202 , n2999 );
    nor g2939 ( n1875 , n1796 , n3212 );
    xnor g2940 ( n597 , n3785 , n1431 );
    and g2941 ( n2984 , n807 , n3860 );
    or g2942 ( n2315 , n3449 , n2416 );
    and g2943 ( n986 , n2163 , n1752 );
    not g2944 ( n1685 , n3506 );
    or g2945 ( n1549 , n130 , n3343 );
    not g2946 ( n3257 , n1628 );
    or g2947 ( n1877 , n300 , n2680 );
    or g2948 ( n914 , n2718 , n1878 );
    or g2949 ( n3891 , n3808 , n2272 );
    xnor g2950 ( n1222 , n2162 , n386 );
    xor g2951 ( n2761 , n2581 , n3151 );
    and g2952 ( n2484 , n1449 , n2536 );
    xnor g2953 ( n1618 , n1656 , n1142 );
    or g2954 ( n771 , n3109 , n452 );
    or g2955 ( n204 , n1084 , n2627 );
    or g2956 ( n1539 , n3061 , n2976 );
    or g2957 ( n786 , n1754 , n2627 );
    xnor g2958 ( n3721 , n1370 , n2602 );
    or g2959 ( n2987 , n2302 , n1503 );
    and g2960 ( n3000 , n3720 , n2746 );
    not g2961 ( n1194 , n1347 );
    or g2962 ( n1944 , n3465 , n2375 );
    or g2963 ( n3416 , n1506 , n2931 );
    and g2964 ( n3273 , n3678 , n769 );
    or g2965 ( n2721 , n462 , n2933 );
    xnor g2966 ( n3397 , n1406 , n2671 );
    and g2967 ( n1116 , n868 , n1129 );
    not g2968 ( n3144 , n88 );
    xnor g2969 ( n3021 , n3545 , n2327 );
    and g2970 ( n3333 , n1510 , n2022 );
    and g2971 ( n1213 , n1059 , n1647 );
    xnor g2972 ( n977 , n1843 , n3825 );
    not g2973 ( n1039 , n740 );
    or g2974 ( n980 , n2655 , n2474 );
    xnor g2975 ( n2788 , n1299 , n2114 );
    not g2976 ( n3166 , n1524 );
    or g2977 ( n3147 , n2339 , n3766 );
    or g2978 ( n2630 , n1974 , n2183 );
    and g2979 ( n2728 , n2063 , n3851 );
    and g2980 ( n1509 , n3413 , n2142 );
    xnor g2981 ( n111 , n1591 , n3636 );
    xnor g2982 ( n2068 , n1494 , n3826 );
    or g2983 ( n2123 , n1163 , n1765 );
    and g2984 ( n1487 , n366 , n3606 );
    or g2985 ( n579 , n499 , n1593 );
    xnor g2986 ( n3588 , n2134 , n2408 );
    not g2987 ( n1193 , n1808 );
    or g2988 ( n1481 , n2269 , n2613 );
    or g2989 ( n1447 , n1936 , n3551 );
    or g2990 ( n497 , n3623 , n2244 );
    not g2991 ( n3798 , n248 );
    and g2992 ( n1395 , n569 , n42 );
    not g2993 ( n138 , n2073 );
    not g2994 ( n1455 , n2572 );
    not g2995 ( n1742 , n829 );
    or g2996 ( n2279 , n469 , n169 );
    or g2997 ( n2892 , n2489 , n2015 );
    and g2998 ( n1483 , n3066 , n1665 );
    xnor g2999 ( n3583 , n2532 , n1637 );
    or g3000 ( n1842 , n1786 , n560 );
    nor g3001 ( n1279 , n2845 , n1001 );
    xor g3002 ( n1506 , n1945 , n2641 );
    or g3003 ( n2196 , n3341 , n364 );
    or g3004 ( n2495 , n266 , n3100 );
    and g3005 ( n1292 , n340 , n1171 );
    xnor g3006 ( n108 , n3541 , n2004 );
    xnor g3007 ( n360 , n1097 , n2338 );
    and g3008 ( n3429 , n1772 , n3735 );
    and g3009 ( n5 , n155 , n3731 );
    not g3010 ( n2066 , n3589 );
    xnor g3011 ( n603 , n26 , n1925 );
    or g3012 ( n1888 , n1207 , n1508 );
    or g3013 ( n206 , n1571 , n3065 );
    or g3014 ( n2879 , n3887 , n2684 );
    not g3015 ( n973 , n705 );
    and g3016 ( n3371 , n2212 , n54 );
    and g3017 ( n1095 , n1492 , n470 );
    or g3018 ( n3724 , n529 , n2256 );
    or g3019 ( n3318 , n751 , n3323 );
    and g3020 ( n3251 , n56 , n2371 );
    and g3021 ( n2928 , n3647 , n643 );
    and g3022 ( n3316 , n1609 , n1241 );
    nor g3023 ( n2494 , n2773 , n1183 );
    or g3024 ( n173 , n11 , n2242 );
    not g3025 ( n1485 , n3344 );
    or g3026 ( n2163 , n2659 , n715 );
    not g3027 ( n3082 , n2202 );
    and g3028 ( n2220 , n3870 , n1795 );
    or g3029 ( n712 , n2682 , n210 );
    not g3030 ( n2783 , n2258 );
    xnor g3031 ( n65 , n2262 , n3816 );
    xnor g3032 ( n1666 , n1893 , n1322 );
    and g3033 ( n2850 , n1326 , n2193 );
    or g3034 ( n3261 , n1564 , n3488 );
    and g3035 ( n2040 , n3375 , n326 );
    or g3036 ( n3530 , n3282 , n1041 );
    or g3037 ( n3667 , n1802 , n2693 );
    and g3038 ( n2358 , n1896 , n1491 );
    not g3039 ( n1954 , n2159 );
    not g3040 ( n85 , n477 );
    or g3041 ( n906 , n912 , n273 );
    or g3042 ( n1088 , n60 , n3128 );
    nor g3043 ( n3177 , n2855 , n915 );
    nor g3044 ( n2675 , n1494 , n674 );
    and g3045 ( n2565 , n2080 , n959 );
    and g3046 ( n2701 , n3377 , n1625 );
    not g3047 ( n2390 , n1827 );
    xnor g3048 ( n2898 , n3018 , n3354 );
    and g3049 ( n98 , n2077 , n993 );
    xnor g3050 ( n1556 , n2763 , n1038 );
    xnor g3051 ( n781 , n2988 , n208 );
    xnor g3052 ( n2718 , n3644 , n2464 );
    or g3053 ( n1313 , n776 , n2472 );
    or g3054 ( n3773 , n1698 , n1918 );
    not g3055 ( n2453 , n2992 );
    and g3056 ( n1705 , n3648 , n2034 );
    and g3057 ( n1287 , n234 , n409 );
    or g3058 ( n247 , n2886 , n2596 );
    xnor g3059 ( n3892 , n347 , n2616 );
    xnor g3060 ( n3471 , n3643 , n3793 );
    xnor g3061 ( n894 , n3709 , n292 );
    or g3062 ( n270 , n790 , n3533 );
    or g3063 ( n350 , n1933 , n3000 );
    not g3064 ( n3343 , n1296 );
    xnor g3065 ( n2827 , n3063 , n2431 );
    or g3066 ( n372 , n1076 , n989 );
    or g3067 ( n3859 , n1852 , n1527 );
    and g3068 ( n896 , n467 , n3325 );
    and g3069 ( n39 , n3226 , n1689 );
    or g3070 ( n1457 , n2954 , n2950 );
    not g3071 ( n3831 , n3365 );
    or g3072 ( n2327 , n2233 , n2350 );
    nor g3073 ( n432 , n1911 , n3666 );
    not g3074 ( n948 , n1775 );
    not g3075 ( n2536 , n2112 );
    not g3076 ( n1569 , n928 );
    and g3077 ( n2734 , n1615 , n2941 );
    or g3078 ( n1703 , n2052 , n1466 );
    not g3079 ( n2510 , n1761 );
    and g3080 ( n1498 , n2143 , n3524 );
    not g3081 ( n2926 , n1066 );
    not g3082 ( n3732 , n2055 );
    and g3083 ( n2185 , n2196 , n1346 );
    or g3084 ( n22 , n1612 , n3554 );
    xnor g3085 ( n263 , n2997 , n3085 );
    nor g3086 ( n2323 , n3344 , n2709 );
    or g3087 ( n2465 , n3433 , n1679 );
    or g3088 ( n2082 , n1271 , n2154 );
    nor g3089 ( n1678 , n265 , n972 );
    xnor g3090 ( n2661 , n3819 , n864 );
    xnor g3091 ( n2597 , n1885 , n668 );
    not g3092 ( n38 , n3510 );
    or g3093 ( n3902 , n2612 , n834 );
    xnor g3094 ( n1991 , n1221 , n1654 );
    or g3095 ( n2500 , n2367 , n1643 );
    xnor g3096 ( n3286 , n827 , n1480 );
    xnor g3097 ( n495 , n2497 , n2300 );
    and g3098 ( n362 , n1431 , n3703 );
    not g3099 ( n1180 , n1761 );
    and g3100 ( n1486 , n979 , n2517 );
    and g3101 ( n2902 , n439 , n1730 );
    and g3102 ( n1013 , n2031 , n1240 );
    and g3103 ( n616 , n802 , n247 );
    or g3104 ( n711 , n1655 , n2817 );
    nor g3105 ( n286 , n2336 , n839 );
    or g3106 ( n1946 , n2807 , n2020 );
    or g3107 ( n450 , n2150 , n1773 );
    or g3108 ( n2699 , n3677 , n2884 );
    xnor g3109 ( n2551 , n3606 , n2058 );
    and g3110 ( n508 , n990 , n2024 );
    and g3111 ( n1743 , n1152 , n324 );
    and g3112 ( n3787 , n1481 , n870 );
    or g3113 ( n1289 , n3206 , n3238 );
    and g3114 ( n1092 , n952 , n2645 );
    and g3115 ( n3404 , n2653 , n3070 );
    not g3116 ( n536 , n2889 );
    or g3117 ( n3346 , n3759 , n1194 );
    and g3118 ( n2164 , n2441 , n2858 );
    or g3119 ( n3165 , n644 , n3174 );
    nor g3120 ( n1048 , n2484 , n2919 );
    or g3121 ( n2376 , n1935 , n2487 );
    xnor g3122 ( n668 , n786 , n2025 );
    xnor g3123 ( n2854 , n3901 , n2898 );
    or g3124 ( n3036 , n2482 , n1056 );
    or g3125 ( n3792 , n299 , n2439 );
    not g3126 ( n1492 , n3802 );
    or g3127 ( n796 , n457 , n1086 );
    or g3128 ( n423 , n8 , n3698 );
    not g3129 ( n1315 , n523 );
    nor g3130 ( n2753 , n841 , n101 );
    not g3131 ( n583 , n66 );
    not g3132 ( n3725 , n3536 );
    and g3133 ( n1554 , n693 , n2049 );
    and g3134 ( n2273 , n2363 , n3699 );
    or g3135 ( n2210 , n2328 , n2169 );
    and g3136 ( n126 , n3682 , n1888 );
    or g3137 ( n2395 , n3121 , n831 );
    and g3138 ( n3772 , n81 , n3692 );
    or g3139 ( n1079 , n2364 , n3270 );
    and g3140 ( n190 , n3251 , n2745 );
    or g3141 ( n2653 , n590 , n3208 );
    not g3142 ( n3157 , n866 );
    xnor g3143 ( n3457 , n2524 , n1219 );
    and g3144 ( n3585 , n140 , n676 );
    or g3145 ( n963 , n1146 , n281 );
    not g3146 ( n1884 , n1103 );
    and g3147 ( n2410 , n3706 , n1205 );
    xnor g3148 ( n278 , n437 , n3247 );
    and g3149 ( n1030 , n196 , n794 );
    or g3150 ( n3374 , n1011 , n800 );
    xnor g3151 ( n2286 , n2482 , n2152 );
    or g3152 ( n1982 , n2946 , n1266 );
    xnor g3153 ( n199 , n188 , n3792 );
    not g3154 ( n419 , n2812 );
    not g3155 ( n611 , n2886 );
    xnor g3156 ( n2491 , n2267 , n2138 );
    or g3157 ( n2616 , n2789 , n2783 );
    xnor g3158 ( n168 , n1039 , n3033 );
    nor g3159 ( n2825 , n1841 , n1034 );
    and g3160 ( n1358 , n2283 , n1324 );
    or g3161 ( n1366 , n33 , n2670 );
    xnor g3162 ( n518 , n630 , n2754 );
    and g3163 ( n1307 , n1493 , n1900 );
    or g3164 ( n1957 , n1886 , n2388 );
    xnor g3165 ( n260 , n2143 , n76 );
    or g3166 ( n837 , n2781 , n2799 );
    not g3167 ( n2997 , n167 );
    or g3168 ( n3464 , n986 , n1715 );
    xnor g3169 ( n2456 , n1733 , n931 );
    not g3170 ( n3233 , n3092 );
    xnor g3171 ( n2304 , n566 , n2384 );
    and g3172 ( n1312 , n399 , n214 );
    not g3173 ( n272 , n482 );
    and g3174 ( n2882 , n1645 , n2018 );
    and g3175 ( n2262 , n3427 , n3469 );
    or g3176 ( n1713 , n2678 , n744 );
    or g3177 ( n2101 , n2265 , n1 );
    or g3178 ( n1135 , n2588 , n3144 );
    and g3179 ( n2620 , n3464 , n2904 );
    or g3180 ( n3289 , n712 , n1996 );
    not g3181 ( n2305 , n2463 );
    or g3182 ( n1579 , n553 , n1553 );
    xnor g3183 ( n3600 , n863 , n594 );
    or g3184 ( n2075 , n1824 , n3756 );
    and g3185 ( n3542 , n3594 , n2415 );
    not g3186 ( n989 , n1234 );
    or g3187 ( n2485 , n3831 , n2413 );
    or g3188 ( n2913 , n446 , n1905 );
    not g3189 ( n1547 , n1521 );
    xnor g3190 ( n1714 , n2014 , n924 );
    and g3191 ( n2247 , n571 , n1861 );
    not g3192 ( n2090 , n3426 );
    xnor g3193 ( n3670 , n1417 , n1737 );
    or g3194 ( n62 , n242 , n2287 );
    and g3195 ( n1418 , n1624 , n1338 );
    xnor g3196 ( n2385 , n2136 , n3286 );
    or g3197 ( n3508 , n1999 , n1895 );
    or g3198 ( n140 , n3734 , n3045 );
    and g3199 ( n1667 , n2266 , n2232 );
    xnor g3200 ( n3247 , n2028 , n2452 );
    xnor g3201 ( n1239 , n1770 , n2637 );
    xnor g3202 ( n3504 , n1415 , n3322 );
    xor g3203 ( n585 , n318 , n3670 );
    not g3204 ( n3512 , n1211 );
    and g3205 ( n1789 , n3419 , n1330 );
    nor g3206 ( n667 , n1808 , n2493 );
    or g3207 ( n1745 , n1131 , n1829 );
    not g3208 ( n714 , n3587 );
    or g3209 ( n14 , n2990 , n2153 );
    xnor g3210 ( n2212 , n3511 , n3559 );
    not g3211 ( n1018 , n1804 );
    and g3212 ( n175 , n347 , n1847 );
    nor g3213 ( n2823 , n2018 , n1645 );
    or g3214 ( n2106 , n2359 , n3542 );
    nor g3215 ( n435 , n3311 , n2636 );
    or g3216 ( n193 , n1649 , n172 );
    or g3217 ( n188 , n754 , n2696 );
    xor g3218 ( n2857 , n361 , n561 );
    not g3219 ( n809 , n504 );
    xnor g3220 ( n1124 , n3473 , n153 );
    or g3221 ( n3851 , n3601 , n250 );
    not g3222 ( n1467 , n53 );
    xnor g3223 ( n1093 , n2867 , n2401 );
    or g3224 ( n1795 , n467 , n3325 );
    or g3225 ( n1205 , n942 , n1478 );
    xnor g3226 ( n1493 , n467 , n1894 );
    and g3227 ( n1394 , n2829 , n2116 );
    and g3228 ( n1684 , n2691 , n3147 );
    not g3229 ( n1821 , n2190 );
    or g3230 ( n1475 , n2071 , n1955 );
    and g3231 ( n689 , n2299 , n270 );
    not g3232 ( n858 , n2402 );
    or g3233 ( n2235 , n295 , n1357 );
    and g3234 ( n3760 , n1337 , n207 );
    or g3235 ( n424 , n2025 , n3415 );
    xor g3236 ( n456 , n2387 , n1917 );
    nor g3237 ( n180 , n1345 , n1539 );
    not g3238 ( n3469 , n2112 );
    not g3239 ( n1981 , n2664 );
    or g3240 ( n1303 , n2324 , n456 );
    not g3241 ( n1060 , n687 );
    or g3242 ( n3778 , n3685 , n1471 );
    and g3243 ( n1553 , n478 , n1106 );
    or g3244 ( n2503 , n1092 , n3787 );
    not g3245 ( n2498 , n2223 );
    or g3246 ( n3890 , n2655 , n3650 );
    xnor g3247 ( n3037 , n337 , n289 );
    xnor g3248 ( n2294 , n1634 , n1069 );
    xnor g3249 ( n2168 , n1776 , n3483 );
    xnor g3250 ( n2603 , n1892 , n1636 );
    xnor g3251 ( n2952 , n2855 , n1883 );
    or g3252 ( n2988 , n2682 , n858 );
    not g3253 ( n54 , n3465 );
    not g3254 ( n3486 , n2484 );
    xnor g3255 ( n2700 , n759 , n1143 );
    not g3256 ( n2531 , n2244 );
    not g3257 ( n3172 , n2760 );
    or g3258 ( n3326 , n118 , n1964 );
    xnor g3259 ( n2639 , n943 , n2461 );
    xnor g3260 ( n909 , n3422 , n1454 );
    or g3261 ( n2606 , n2911 , n759 );
    or g3262 ( n2109 , n1098 , n2312 );
    or g3263 ( n3362 , n1002 , n1000 );
    and g3264 ( n617 , n2316 , n619 );
    not g3265 ( n3001 , n3610 );
    and g3266 ( n2373 , n3050 , n2082 );
    or g3267 ( n2618 , n2866 , n1774 );
    or g3268 ( n2024 , n2497 , n2300 );
    or g3269 ( n2266 , n2358 , n3423 );
    not g3270 ( n2079 , n1469 );
    not g3271 ( n299 , n1240 );
    xnor g3272 ( n3152 , n1347 , n3515 );
    or g3273 ( n1636 , n754 , n2094 );
    xor g3274 ( n2297 , n3743 , n930 );
    or g3275 ( n1959 , n284 , n660 );
    and g3276 ( n3212 , n3640 , n1747 );
    or g3277 ( n1023 , n2731 , n3738 );
    and g3278 ( n301 , n1902 , n552 );
    nor g3279 ( n649 , n507 , n484 );
    and g3280 ( n3484 , n1607 , n3862 );
    and g3281 ( n924 , n3331 , n1464 );
    or g3282 ( n1990 , n329 , n515 );
    xnor g3283 ( n1324 , n1959 , n3192 );
    xnor g3284 ( n2807 , n160 , n2621 );
    or g3285 ( n2337 , n3569 , n1008 );
    or g3286 ( n838 , n2509 , n2771 );
    and g3287 ( n507 , n2390 , n1013 );
    nor g3288 ( n1264 , n3198 , n3248 );
    not g3289 ( n1929 , n935 );
    or g3290 ( n1323 , n2662 , n401 );
    xor g3291 ( n3291 , n2056 , n454 );
    not g3292 ( n3163 , n928 );
    or g3293 ( n2737 , n2765 , n134 );
    and g3294 ( n2891 , n2343 , n343 );
    and g3295 ( n3206 , n1559 , n612 );
    not g3296 ( n1127 , n2757 );
    not g3297 ( n1214 , n1672 );
    or g3298 ( n2596 , n3378 , n1962 );
    nor g3299 ( n367 , n1604 , n1907 );
    or g3300 ( n1430 , n187 , n1683 );
    xnor g3301 ( n3643 , n1396 , n1314 );
    or g3302 ( n2881 , n1968 , n764 );
    nor g3303 ( n3214 , n964 , n3435 );
    not g3304 ( n2270 , n1682 );
    xor g3305 ( n1616 , n3855 , n3721 );
    not g3306 ( n1910 , n3493 );
    or g3307 ( n2953 , n3424 , n1004 );
    or g3308 ( n2396 , n801 , n3041 );
    or g3309 ( n3009 , n3413 , n2142 );
    or g3310 ( n687 , n3877 , n3257 );
    xnor g3311 ( n3046 , n2678 , n252 );
    xnor g3312 ( n1348 , n2392 , n1581 );
    not g3313 ( n3754 , n1140 );
    xnor g3314 ( n1233 , n3428 , n729 );
    xor g3315 ( n2322 , n2294 , n1201 );
    or g3316 ( n3170 , n2386 , n3223 );
    or g3317 ( n1429 , n994 , n3517 );
    not g3318 ( n2894 , n1845 );
    or g3319 ( n2836 , n3163 , n1872 );
    not g3320 ( n488 , n1140 );
    and g3321 ( n1899 , n636 , n251 );
    and g3322 ( n1937 , n319 , n916 );
    xnor g3323 ( n546 , n1403 , n2089 );
    not g3324 ( n0 , n3038 );
    or g3325 ( n2178 , n1806 , n3230 );
    not g3326 ( n3403 , n47 );
    or g3327 ( n2535 , n1990 , n700 );
    or g3328 ( n582 , n2181 , n3292 );
    or g3329 ( n719 , n2775 , n3461 );
    or g3330 ( n3246 , n2253 , n2478 );
    or g3331 ( n3474 , n236 , n2689 );
    xnor g3332 ( n1377 , n2156 , n3885 );
    xnor g3333 ( n293 , n1448 , n94 );
    xnor g3334 ( n917 , n18 , n3256 );
    or g3335 ( n266 , n2539 , n486 );
    or g3336 ( n81 , n1511 , n367 );
    xor g3337 ( n2979 , n2728 , n1317 );
    and g3338 ( n305 , n634 , n1530 );
    not g3339 ( n1263 , n711 );
    or g3340 ( n2608 , n62 , n3545 );
    xnor g3341 ( n2134 , n1430 , n1769 );
    not g3342 ( n3164 , n3444 );
    or g3343 ( n324 , n762 , n1380 );
    or g3344 ( n2691 , n1158 , n406 );
    and g3345 ( n1871 , n3133 , n3821 );
    and g3346 ( n303 , n3137 , n3568 );
    not g3347 ( n358 , n1793 );
    nor g3348 ( n1238 , n532 , n2907 );
    or g3349 ( n348 , n272 , n85 );
    not g3350 ( n881 , n308 );
    or g3351 ( n3854 , n735 , n2083 );
    and g3352 ( n2310 , n3570 , n1973 );
    not g3353 ( n1177 , n3759 );
    and g3354 ( n3702 , n814 , n1325 );
    and g3355 ( n2818 , n2989 , n2186 );
    and g3356 ( n3230 , n2235 , n2968 );
    xor g3357 ( n2638 , n820 , n3075 );
    and g3358 ( n464 , n3416 , n1286 );
    or g3359 ( n1248 , n3556 , n1411 );
    not g3360 ( n720 , n1160 );
    xnor g3361 ( n2029 , n831 , n2589 );
    or g3362 ( n3031 , n3901 , n3018 );
    or g3363 ( n3768 , n2998 , n1987 );
    not g3364 ( n3412 , n1638 );
    or g3365 ( n3901 , n342 , n334 );
    or g3366 ( n1274 , n2528 , n2057 );
    or g3367 ( n415 , n1688 , n1247 );
    xnor g3368 ( n3515 , n1177 , n1303 );
    not g3369 ( n1284 , n2514 );
    not g3370 ( n2935 , n866 );
    and g3371 ( n1533 , n3176 , n3686 );
    xnor g3372 ( n316 , n842 , n3823 );
    not g3373 ( n2326 , n670 );
    or g3374 ( n259 , n287 , n3498 );
    xnor g3375 ( n698 , n190 , n3206 );
    or g3376 ( n425 , n2735 , n1840 );
    or g3377 ( n2960 , n979 , n2517 );
    not g3378 ( n1915 , n2376 );
    or g3379 ( n2200 , n2705 , n2615 );
    and g3380 ( n1675 , n1631 , n59 );
    xnor g3381 ( n3646 , n1749 , n3141 );
    xnor g3382 ( n3858 , n1827 , n1632 );
    and g3383 ( n2651 , n189 , n1814 );
    or g3384 ( n3138 , n30 , n1589 );
    not g3385 ( n2714 , n2532 );
    not g3386 ( n3111 , n3559 );
    xnor g3387 ( n1451 , n893 , n244 );
    or g3388 ( n2720 , n1610 , n2955 );
    xnor g3389 ( n3162 , n3890 , n3307 );
    or g3390 ( n2145 , n2334 , n1640 );
    or g3391 ( n3375 , n3687 , n126 );
    not g3392 ( n1890 , n1240 );
    and g3393 ( n3419 , n184 , n905 );
    or g3394 ( n3751 , n2886 , n2067 );
    and g3395 ( n1924 , n3118 , n721 );
    not g3396 ( n1016 , n44 );
    or g3397 ( n3781 , n1044 , n3708 );
    or g3398 ( n2203 , n3060 , n3473 );
    or g3399 ( n2264 , n2999 , n2730 );
    or g3400 ( n2000 , n1808 , n817 );
    and g3401 ( n2074 , n796 , n224 );
    or g3402 ( n3448 , n961 , n1245 );
    xnor g3403 ( n2595 , n865 , n1123 );
    xnor g3404 ( n1914 , n3508 , n977 );
    or g3405 ( n1721 , n1621 , n55 );
    or g3406 ( n1091 , n1203 , n1048 );
    xor g3407 ( n1049 , n2336 , n100 );
    nor g3408 ( n1215 , n3502 , n525 );
    and g3409 ( n3245 , n3485 , n2863 );
    xnor g3410 ( n3002 , n131 , n1450 );
    xnor g3411 ( n2486 , n2231 , n1891 );
    or g3412 ( n3802 , n1315 , n3098 );
    and g3413 ( n1040 , n2614 , n144 );
    or g3414 ( n1181 , n1742 , n2061 );
    xnor g3415 ( n1157 , n3789 , n414 );
    xor g3416 ( n1787 , n1390 , n981 );
    or g3417 ( n3466 , n1033 , n856 );
    nor g3418 ( n485 , n2520 , n1904 );
    not g3419 ( n281 , n2640 );
    xnor g3420 ( n2035 , n3628 , n685 );
    not g3421 ( n1822 , n523 );
    or g3422 ( n3803 , n1455 , n471 );
    nor g3423 ( n825 , n482 , n477 );
    or g3424 ( n3280 , n3458 , n960 );
    not g3425 ( n174 , n4 );
    xnor g3426 ( n74 , n3543 , n728 );
    or g3427 ( n647 , n3276 , n43 );
    nor g3428 ( n892 , n3784 , n2874 );
    or g3429 ( n2844 , n2356 , n3470 );
    or g3430 ( n107 , n11 , n1706 );
    xnor g3431 ( n2436 , n278 , n1302 );
    xnor g3432 ( n275 , n3002 , n1173 );
    and g3433 ( n1902 , n3436 , n2172 );
    or g3434 ( n3035 , n3428 , n2903 );
    and g3435 ( n2025 , n1500 , n14 );
    not g3436 ( n2538 , n2195 );
    or g3437 ( n1757 , n342 , n320 );
    not g3438 ( n2435 , n1266 );
    nor g3439 ( n897 , n2062 , n213 );
    xnor g3440 ( n13 , n449 , n164 );
    and g3441 ( n2901 , n3601 , n250 );
    or g3442 ( n1953 , n173 , n3161 );
    or g3443 ( n313 , n3084 , n734 );
    xnor g3444 ( n2400 , n1609 , n1816 );
    or g3445 ( n645 , n3799 , n2777 );
    and g3446 ( n1577 , n696 , n1108 );
    or g3447 ( n3350 , n2186 , n2096 );
    xnor g3448 ( n2312 , n1022 , n615 );
    not g3449 ( n1327 , n1507 );
    or g3450 ( n1106 , n1623 , n1780 );
    not g3451 ( n486 , n1140 );
    not g3452 ( n1771 , n3481 );
    not g3453 ( n2650 , n1793 );
    not g3454 ( n314 , n1539 );
    xnor g3455 ( n2816 , n3822 , n1033 );
    not g3456 ( n533 , n3536 );
    and g3457 ( n2054 , n2346 , n3468 );
    or g3458 ( n3813 , n1555 , n2076 );
    or g3459 ( n3057 , n3757 , n1448 );
    or g3460 ( n3470 , n284 , n2305 );
    and g3461 ( n1996 , n411 , n2448 );
    and g3462 ( n2365 , n2961 , n3790 );
    and g3463 ( n2965 , n1865 , n2221 );
    or g3464 ( n1652 , n2886 , n3414 );
    not g3465 ( n3091 , n2073 );
    or g3466 ( n1210 , n2130 , n713 );
    xor g3467 ( n3190 , n2866 , n1774 );
    or g3468 ( n789 , n859 , n1259 );
    and g3469 ( n2613 , n2255 , n3544 );
    nor g3470 ( n2817 , n2706 , n930 );
    or g3471 ( n1997 , n1743 , n1971 );
    not g3472 ( n2522 , n109 );
    nor g3473 ( n1876 , n3227 , n614 );
    xnor g3474 ( n2578 , n1526 , n2173 );
    or g3475 ( n2779 , n651 , n1054 );
    nor g3476 ( n1102 , n2813 , n3167 );
    xnor g3477 ( n1426 , n1697 , n1224 );
    nor g3478 ( n3296 , n1095 , n316 );
    xnor g3479 ( n2277 , n1735 , n1111 );
    xnor g3480 ( n3269 , n3738 , n3871 );
    not g3481 ( n158 , n2463 );
    not g3482 ( n845 , n196 );
    or g3483 ( n799 , n2136 , n2438 );
    and g3484 ( n3747 , n394 , n2176 );
    and g3485 ( n1844 , n652 , n1178 );
    or g3486 ( n1958 , n3809 , n3208 );
    or g3487 ( n1098 , n417 , n620 );
    or g3488 ( n3352 , n766 , n1712 );
    xnor g3489 ( n390 , n737 , n3714 );
    or g3490 ( n2956 , n2812 , n354 );
    not g3491 ( n620 , n940 );
    xnor g3492 ( n2729 , n332 , n2853 );
    not g3493 ( n576 , n670 );
    or g3494 ( n564 , n2695 , n3363 );
    and g3495 ( n664 , n2737 , n2697 );
    or g3496 ( n1139 , n2576 , n372 );
    xnor g3497 ( n46 , n3685 , n1531 );
    not g3498 ( n1994 , n3506 );
    not g3499 ( n3191 , n186 );
    xnor g3500 ( n3564 , n1118 , n3225 );
    not g3501 ( n1907 , n3112 );
    or g3502 ( n673 , n1837 , n1046 );
    and g3503 ( n2480 , n1931 , n246 );
    or g3504 ( n1299 , n118 , n3150 );
    or g3505 ( n156 , n3501 , n825 );
    xnor g3506 ( n2072 , n830 , n2680 );
    xnor g3507 ( n1261 , n1648 , n2181 );
    xnor g3508 ( n431 , n1256 , n263 );
    and g3509 ( n3505 , n437 , n2028 );
    or g3510 ( n932 , n941 , n815 );
    or g3511 ( n3395 , n704 , n948 );
    and g3512 ( n2876 , n1243 , n791 );
    xnor g3513 ( n594 , n1318 , n2513 );
    or g3514 ( n2209 , n3725 , n401 );
    or g3515 ( n2533 , n216 , n2184 );
    or g3516 ( n3073 , n2156 , n1766 );
    not g3517 ( n341 , n2919 );
    and g3518 ( n2799 , n2853 , n3001 );
    not g3519 ( n2587 , n2714 );
    nor g3520 ( n3836 , n3465 , n3043 );
    xnor g3521 ( n1230 , n1452 , n142 );
    xnor g3522 ( n3440 , n1002 , n875 );
    and g3523 ( n343 , n297 , n323 );
    nor g3524 ( n2427 , n3027 , n787 );
    or g3525 ( n3476 , n3522 , n1676 );
    and g3526 ( n1722 , n2383 , n3216 );
    and g3527 ( n2813 , n2426 , n1972 );
    not g3528 ( n853 , n963 );
    not g3529 ( n3602 , n2121 );
    and g3530 ( n1989 , n1707 , n3621 );
    xnor g3531 ( n637 , n2801 , n3126 );
    not g3532 ( n3004 , n1025 );
    xnor g3533 ( n45 , n1647 , n136 );
    and g3534 ( n855 , n75 , n3477 );
    xnor g3535 ( n48 , n1168 , n2733 );
    nor g3536 ( n27 , n3371 , n1672 );
    and g3537 ( n572 , n3129 , n1479 );
    or g3538 ( n1385 , n3478 , n2274 );
    xnor g3539 ( n36 , n2899 , n2366 );
    or g3540 ( n131 , n2974 , n948 );
    and g3541 ( n3188 , n3820 , n2407 );
    or g3542 ( n1057 , n1513 , n2905 );
    not g3543 ( n1535 , n1404 );
    and g3544 ( n828 , n1336 , n2396 );
    or g3545 ( n3128 , n549 , n989 );
    xnor g3546 ( n2496 , n266 , n2182 );
    xnor g3547 ( n862 , n2593 , n711 );
    nor g3548 ( n2771 , n2937 , n616 );
    not g3549 ( n1969 , n3103 );
    or g3550 ( n1237 , n1144 , n3791 );
    and g3551 ( n3433 , n3709 , n3646 );
    or g3552 ( n2819 , n1125 , n2217 );
    not g3553 ( n1405 , n1200 );
    not g3554 ( n880 , n2270 );
    nor g3555 ( n1339 , n1656 , n3034 );
    or g3556 ( n2392 , n221 , n2743 );
    or g3557 ( n2846 , n1016 , n2510 );
    or g3558 ( n2172 , n2430 , n2989 );
    xnor g3559 ( n1294 , n1471 , n46 );
    or g3560 ( n3249 , n637 , n2908 );
    xnor g3561 ( n1867 , n962 , n3856 );
    and g3562 ( n3142 , n2791 , n1136 );
    xnor g3563 ( n2878 , n1821 , n2749 );
    xnor g3564 ( n560 , n1674 , n1147 );
    or g3565 ( n2950 , n3827 , n1232 );
    xnor g3566 ( n104 , n953 , n2381 );
    nor g3567 ( n3054 , n761 , n3695 );
    not g3568 ( n2113 , n2270 );
    xnor g3569 ( n2547 , n3174 , n2839 );
    and g3570 ( n3380 , n1227 , n3839 );
    or g3571 ( n2678 , n1505 , n3571 );
    xnor g3572 ( n8 , n1227 , n2352 );
    or g3573 ( n3203 , n3047 , n3124 );
    xnor g3574 ( n2800 , n1629 , n2963 );
    not g3575 ( n471 , n1775 );
    and g3576 ( n371 , n3168 , n2958 );
    and g3577 ( n3394 , n1172 , n390 );
    and g3578 ( n1854 , n2103 , n396 );
    not g3579 ( n543 , n361 );
    not g3580 ( n3815 , n1191 );
    or g3581 ( n569 , n909 , n3068 );
    not g3582 ( n2444 , n740 );
    xnor g3583 ( n3806 , n609 , n322 );
    and g3584 ( n2851 , n2576 , n372 );
    or g3585 ( n2457 , n976 , n2246 );
    or g3586 ( n1756 , n2997 , n3085 );
    or g3587 ( n239 , n2494 , n3776 );
    and g3588 ( n3151 , n3540 , n1580 );
    nor g3589 ( n3024 , n1499 , n3637 );
    and g3590 ( n3791 , n2570 , n311 );
    not g3591 ( n1978 , n3384 );
    xnor g3592 ( n1564 , n1570 , n2896 );
    or g3593 ( n3410 , n2012 , n1723 );
    or g3594 ( n233 , n3617 , n1803 );
    not g3595 ( n1800 , n1367 );
    or g3596 ( n1027 , n2093 , n1751 );
    xnor g3597 ( n354 , n240 , n2092 );
    and g3598 ( n166 , n3174 , n644 );
    xnor g3599 ( n3658 , n1108 , n3408 );
    nor g3600 ( n1340 , n1321 , n90 );
    nor g3601 ( n1700 , n2669 , n2823 );
    xnor g3602 ( n3729 , n3184 , n3833 );
    or g3603 ( n2125 , n688 , n3865 );
    or g3604 ( n2780 , n1685 , n1783 );
    nor g3605 ( n1155 , n721 , n3118 );
    and g3606 ( n3003 , n3476 , n2515 );
    not g3607 ( n2245 , n926 );
    or g3608 ( n99 , n3486 , n341 );
    xor g3609 ( n1449 , n2420 , n2906 );
    and g3610 ( n521 , n950 , n639 );
    xor g3611 ( n686 , n3231 , n2967 );
    xnor g3612 ( n1344 , n2654 , n3517 );
    nor g3613 ( n2976 , n13 , n3581 );
    xor g3614 ( n228 , n2685 , n219 );
    and g3615 ( n607 , n1223 , n2049 );
    xnor g3616 ( n526 , n1125 , n2983 );
    xnor g3617 ( n3427 , n2349 , n172 );
    xnor g3618 ( n1408 , n2506 , n1958 );
    nor g3619 ( n1277 , n9 , n1015 );
    and g3620 ( n1715 , n2174 , n280 );
    not g3621 ( n851 , n2664 );
    or g3622 ( n1304 , n978 , n416 );
    or g3623 ( n297 , n2074 , n301 );
    nor g3624 ( n2278 , n1635 , n3608 );
    and g3625 ( n721 , n3763 , n2585 );
    or g3626 ( n1746 , n641 , n3207 );
    nor g3627 ( n2509 , n247 , n802 );
    or g3628 ( n1468 , n1119 , n3571 );
    or g3629 ( n806 , n442 , n2927 );
    xnor g3630 ( n502 , n1604 , n1511 );
    xnor g3631 ( n3161 , n3064 , n1230 );
    or g3632 ( n2407 , n3541 , n823 );
    and g3633 ( n1283 , n277 , n487 );
    and g3634 ( n1038 , n1079 , n2798 );
    nor g3635 ( n1435 , n105 , n659 );
    and g3636 ( n3728 , n408 , n3335 );
    or g3637 ( n510 , n522 , n1179 );
    xnor g3638 ( n1151 , n1622 , n1301 );
    not g3639 ( n3705 , n1156 );
    or g3640 ( n323 , n552 , n1902 );
    and g3641 ( n3145 , n2954 , n2950 );
    or g3642 ( n2448 , n1569 , n2809 );
    or g3643 ( n445 , n2458 , n2009 );
    and g3644 ( n3750 , n1749 , n1474 );
    nor g3645 ( n3409 , n1608 , n1835 );
    xnor g3646 ( n757 , n3618 , n2405 );
    xnor g3647 ( n3872 , n327 , n2215 );
    or g3648 ( n2936 , n2012 , n2350 );
    or g3649 ( n2914 , n768 , n448 );
    not g3650 ( n1198 , n220 );
    or g3651 ( n1052 , n3307 , n3890 );
    or g3652 ( n3838 , n2040 , n2355 );
    and g3653 ( n2575 , n2676 , n3202 );
    or g3654 ( n1036 , n2987 , n3395 );
    or g3655 ( n676 , n145 , n1244 );
    or g3656 ( n814 , n3280 , n2085 );
    xnor g3657 ( n1542 , n752 , n35 );
    not g3658 ( n3794 , n1572 );
    xor g3659 ( n2593 , n2557 , n2562 );
    and g3660 ( n3776 , n3081 , n2041 );
    or g3661 ( n1663 , n3520 , n2679 );
    and g3662 ( n1545 , n3599 , n917 );
    xor g3663 ( n3126 , n3315 , n2100 );
    not g3664 ( n1291 , n499 );
    xnor g3665 ( n243 , n2450 , n3336 );
    or g3666 ( n1819 , n2633 , n3074 );
    or g3667 ( n3689 , n1535 , n281 );
    and g3668 ( n223 , n1149 , n2264 );
    and g3669 ( n1917 , n2833 , n2437 );
    or g3670 ( n3889 , n1808 , n3710 );
    not g3671 ( n3571 , n1820 );
    or g3672 ( n3339 , n386 , n758 );
    not g3673 ( n116 , n2888 );
    or g3674 ( n2573 , n2324 , n1666 );
    and g3675 ( n559 , n3008 , n3175 );
    xnor g3676 ( n306 , n1597 , n1151 );
    or g3677 ( n2353 , n2539 , n2860 );
    xnor g3678 ( n3645 , n468 , n593 );
    and g3679 ( n264 , n512 , n2879 );
    xnor g3680 ( n258 , n1009 , n629 );
    xnor g3681 ( n3654 , n3897 , n346 );
    not g3682 ( n1146 , n955 );
    not g3683 ( n2654 , n3401 );
    or g3684 ( n971 , n982 , n2220 );
    or g3685 ( n3526 , n123 , n3866 );
    and g3686 ( n3850 , n783 , n3171 );
    or g3687 ( n2508 , n2320 , n17 );
    not g3688 ( n2449 , n1568 );
    or g3689 ( n3393 , n1393 , n351 );
    and g3690 ( n3550 , n780 , n1686 );
    or g3691 ( n1105 , n3026 , n3150 );
    xnor g3692 ( n2838 , n1098 , n1245 );
    nor g3693 ( n2141 , n1884 , n2023 );
    or g3694 ( n3553 , n6 , n245 );
    not g3695 ( n1882 , n1463 );
    xnor g3696 ( n1302 , n1966 , n1391 );
    not g3697 ( n1107 , n3340 );
    or g3698 ( n2188 , n2763 , n1038 );
    xnor g3699 ( n2943 , n316 , n3042 );
    xnor g3700 ( n1306 , n687 , n3696 );
    not g3701 ( n242 , n335 );
    xnor g3702 ( n2170 , n3127 , n1899 );
    nor g3703 ( n2683 , n607 , n865 );
    xnor g3704 ( n3801 , n2154 , n3345 );
    xor g3705 ( n225 , n227 , n1738 );
    or g3706 ( n71 , n1330 , n3419 );
    xor g3707 ( n1223 , n1613 , n678 );
    or g3708 ( n1785 , n3303 , n2321 );
    or g3709 ( n3211 , n2330 , n3149 );
    and g3710 ( n3513 , n3740 , n1909 );
    or g3711 ( n2214 , n1242 , n339 );
    xnor g3712 ( n3807 , n963 , n1231 );
    xnor g3713 ( n2489 , n1124 , n2501 );
    xor g3714 ( n3611 , n1786 , n1397 );
    or g3715 ( n2834 , n72 , n1395 );
    and g3716 ( n2431 , n582 , n3260 );
    xnor g3717 ( n2441 , n823 , n108 );
    or g3718 ( n1149 , n1881 , n3673 );
    xnor g3719 ( n3338 , n2615 , n2942 );
    or g3720 ( n1621 , n1372 , n3574 );
    or g3721 ( n3708 , n3752 , n1849 );
    or g3722 ( n3733 , n678 , n1613 );
    not g3723 ( n29 , n504 );
    or g3724 ( n3786 , n514 , n314 );
    xnor g3725 ( n3560 , n2174 , n986 );
    not g3726 ( n2663 , n1638 );
    not g3727 ( n898 , n239 );
    xnor g3728 ( n626 , n834 , n2469 );
    nor g3729 ( n1813 , n1651 , n3672 );
    or g3730 ( n3899 , n1283 , n1264 );
    or g3731 ( n2934 , n903 , n1548 );
    not g3732 ( n1724 , n893 );
    not g3733 ( n3229 , n1187 );
    xnor g3734 ( n1735 , n1840 , n1949 );
    xnor g3735 ( n3366 , n721 , n1818 );
    and g3736 ( n1534 , n2618 , n3361 );
    or g3737 ( n2660 , n1372 , n2684 );
    xnor g3738 ( n1316 , n2858 , n3684 );
    not g3739 ( n3779 , n1432 );
    or g3740 ( n2969 , n565 , n992 );
    and g3741 ( n365 , n468 , n3294 );
    not g3742 ( n2460 , n1671 );
    not g3743 ( n2918 , n2402 );
    and g3744 ( n1515 , n3138 , n2995 );
    and g3745 ( n1410 , n2563 , n610 );
    not g3746 ( n2931 , n3859 );
    not g3747 ( n913 , n4 );
    not g3748 ( n3610 , n3114 );
    or g3749 ( n2342 , n2711 , n2851 );
    xnor g3750 ( n732 , n1708 , n192 );
    or g3751 ( n3184 , n1065 , n606 );
    xnor g3752 ( n2811 , n1860 , n2815 );
    or g3753 ( n352 , n1303 , n238 );
    xnor g3754 ( n3727 , n1902 , n2074 );
    not g3755 ( n2756 , n3662 );
    and g3756 ( n3102 , n1757 , n1501 );
    or g3757 ( n2740 , n3191 , n732 );
    or g3758 ( n26 , n819 , n20 );
    not g3759 ( n2726 , n3237 );
    xnor g3760 ( n3180 , n2211 , n632 );
    and g3761 ( n2259 , n3886 , n3035 );
    or g3762 ( n2786 , n2869 , n2185 );
    xnor g3763 ( n3539 , n766 , n191 );
    not g3764 ( n3547 , n1652 );
    xnor g3765 ( n779 , n652 , n2526 );
    or g3766 ( n511 , n2591 , n334 );
    xnor g3767 ( n1725 , n854 , n1621 );
    or g3768 ( n3734 , n3779 , n434 );
    xnor g3769 ( n3868 , n1930 , n39 );
    or g3770 ( n3240 , n826 , n1384 );
    and g3771 ( n142 , n1497 , n564 );
    and g3772 ( n1733 , n3362 , n3758 );
    or g3773 ( n2930 , n1546 , n3176 );
    and g3774 ( n1963 , n1442 , n1463 );
    and g3775 ( n82 , n1137 , n333 );
    or g3776 ( n1497 , n1422 , n2634 );
    or g3777 ( n409 , n3155 , n3691 );
    or g3778 ( n959 , n3792 , n188 );
    or g3779 ( n756 , n82 , n89 );
    or g3780 ( n328 , n2357 , n176 );
    xnor g3781 ( n2130 , n3407 , n3442 );
    nor g3782 ( n871 , n2822 , n1914 );
    or g3783 ( n1159 , n2324 , n1657 );
    not g3784 ( n2959 , n2726 );
    not g3785 ( n2985 , n3275 );
endmodule
