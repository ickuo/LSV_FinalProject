module top( n2 , n5 , n6 , n7 , n8 , n15 , n27 , n31 , n33 , 
n37 , n40 , n45 , n49 , n58 , n78 , n79 , n83 , n87 , n88 , 
n92 , n98 , n113 , n121 , n123 , n129 , n135 , n143 , n144 , n145 , 
n165 , n168 , n173 , n177 , n181 , n185 , n188 , n196 , n200 , n201 , 
n202 , n204 , n205 , n212 , n213 , n220 , n222 , n226 , n230 , n231 , 
n232 , n245 , n246 , n250 , n251 , n255 , n257 , n258 , n281 , n287 , 
n302 , n324 , n331 , n344 , n349 , n350 , n351 , n354 , n357 , n365 , 
n368 , n369 , n371 , n373 , n378 , n380 , n381 , n382 , n396 , n400 , 
n404 , n415 , n426 , n428 , n429 , n432 , n433 , n439 , n451 , n467 , 
n469 , n474 , n487 , n490 , n494 , n499 , n500 , n502 , n513 , n517 , 
n521 , n523 , n524 , n533 , n539 , n540 , n543 );
    input n2 , n5 , n6 , n8 , n31 , n33 , n40 , n49 , n58 , 
n78 , n79 , n98 , n123 , n129 , n145 , n177 , n181 , n188 , n200 , 
n201 , n202 , n204 , n205 , n213 , n220 , n222 , n230 , n245 , n251 , 
n257 , n287 , n302 , n324 , n331 , n344 , n349 , n351 , n354 , n357 , 
n380 , n396 , n400 , n415 , n428 , n432 , n433 , n451 , n467 , n474 , 
n494 , n500 , n502 , n517 , n521 , n523 , n524 , n533 , n540 , n543 ;
    output n7 , n15 , n27 , n37 , n45 , n83 , n87 , n88 , n92 , 
n113 , n121 , n135 , n143 , n144 , n165 , n168 , n173 , n185 , n196 , 
n212 , n226 , n231 , n232 , n246 , n250 , n255 , n258 , n281 , n350 , 
n365 , n368 , n369 , n371 , n373 , n378 , n381 , n382 , n404 , n426 , 
n429 , n439 , n469 , n487 , n490 , n499 , n513 , n539 ;
    wire n0 , n1 , n3 , n4 , n9 , n10 , n11 , n12 , n13 , 
n14 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , 
n25 , n26 , n28 , n29 , n30 , n32 , n34 , n35 , n36 , n38 , 
n39 , n41 , n42 , n43 , n44 , n46 , n47 , n48 , n50 , n51 , 
n52 , n53 , n54 , n55 , n56 , n57 , n59 , n60 , n61 , n62 , 
n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , 
n73 , n74 , n75 , n76 , n77 , n80 , n81 , n82 , n84 , n85 , 
n86 , n89 , n90 , n91 , n93 , n94 , n95 , n96 , n97 , n99 , 
n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
n110 , n111 , n112 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
n122 , n124 , n125 , n126 , n127 , n128 , n130 , n131 , n132 , n133 , 
n134 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n146 , n147 , 
n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , 
n158 , n159 , n160 , n161 , n162 , n163 , n164 , n166 , n167 , n169 , 
n170 , n171 , n172 , n174 , n175 , n176 , n178 , n179 , n180 , n182 , 
n183 , n184 , n186 , n187 , n189 , n190 , n191 , n192 , n193 , n194 , 
n195 , n197 , n198 , n199 , n203 , n206 , n207 , n208 , n209 , n210 , 
n211 , n214 , n215 , n216 , n217 , n218 , n219 , n221 , n223 , n224 , 
n225 , n227 , n228 , n229 , n233 , n234 , n235 , n236 , n237 , n238 , 
n239 , n240 , n241 , n242 , n243 , n244 , n247 , n248 , n249 , n252 , 
n253 , n254 , n256 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , 
n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , 
n276 , n277 , n278 , n279 , n280 , n282 , n283 , n284 , n285 , n286 , 
n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , 
n298 , n299 , n300 , n301 , n303 , n304 , n305 , n306 , n307 , n308 , 
n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , 
n319 , n320 , n321 , n322 , n323 , n325 , n326 , n327 , n328 , n329 , 
n330 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , 
n341 , n342 , n343 , n345 , n346 , n347 , n348 , n352 , n353 , n355 , 
n356 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n366 , n367 , 
n370 , n372 , n374 , n375 , n376 , n377 , n379 , n383 , n384 , n385 , 
n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , 
n397 , n398 , n399 , n401 , n402 , n403 , n405 , n406 , n407 , n408 , 
n409 , n410 , n411 , n412 , n413 , n414 , n416 , n417 , n418 , n419 , 
n420 , n421 , n422 , n423 , n424 , n425 , n427 , n430 , n431 , n434 , 
n435 , n436 , n437 , n438 , n440 , n441 , n442 , n443 , n444 , n445 , 
n446 , n447 , n448 , n449 , n450 , n452 , n453 , n454 , n455 , n456 , 
n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , 
n468 , n470 , n471 , n472 , n473 , n475 , n476 , n477 , n478 , n479 , 
n480 , n481 , n482 , n483 , n484 , n485 , n486 , n488 , n489 , n491 , 
n492 , n493 , n495 , n496 , n497 , n498 , n501 , n503 , n504 , n505 , 
n506 , n507 , n508 , n509 , n510 , n511 , n512 , n514 , n515 , n516 , 
n518 , n519 , n520 , n522 , n525 , n526 , n527 , n528 , n529 , n530 , 
n531 , n532 , n534 , n535 , n536 , n537 , n538 , n541 , n542 , n544 , 
n545 , n546 ;
    nor g0 ( n272 , n540 , n58 );
    and g1 ( n353 , n215 , n59 );
    buf g2 ( n526 , n116 );
    nor g3 ( n227 , n188 , n95 );
    xnor g4 ( n240 , n231 , n108 );
    and g5 ( n55 , n228 , n483 );
    xnor g6 ( n113 , n76 , n320 );
    or g7 ( n194 , n217 , n480 );
    and g8 ( n450 , n271 , n263 );
    nor g9 ( n424 , n433 , n488 );
    or g10 ( n108 , n51 , n436 );
    and g11 ( n341 , n103 , n458 );
    and g12 ( n484 , n468 , n180 );
    and g13 ( n274 , n401 , n62 );
    xnor g14 ( n369 , n421 , n466 );
    and g15 ( n159 , n213 , n241 );
    or g16 ( n329 , n478 , n104 );
    nor g17 ( n170 , n202 , n291 );
    not g18 ( n491 , n188 );
    xnor g19 ( n234 , n127 , n526 );
    and g20 ( n280 , n307 , n292 );
    or g21 ( n218 , n450 , n544 );
    or g22 ( n335 , n306 , n391 );
    and g23 ( n464 , n481 , n48 );
    xnor g24 ( n496 , n300 , n32 );
    or g25 ( n401 , n468 , n387 );
    nor g26 ( n465 , n437 , n388 );
    xnor g27 ( n348 , n245 , n344 );
    xnor g28 ( n486 , n218 , n125 );
    xnor g29 ( n121 , n96 , n482 );
    or g30 ( n46 , n311 , n261 );
    nor g31 ( n541 , n202 , n79 );
    nor g32 ( n293 , n202 , n336 );
    not g33 ( n294 , n423 );
    or g34 ( n308 , n73 , n4 );
    not g35 ( n326 , n539 );
    not g36 ( n21 , n180 );
    nor g37 ( n391 , n314 , n81 );
    not g38 ( n534 , n286 );
    not g39 ( n193 , n146 );
    xnor g40 ( n221 , n219 , n66 );
    and g41 ( n480 , n406 , n190 );
    or g42 ( n448 , n219 , n59 );
    xnor g43 ( n239 , n83 , n461 );
    and g44 ( n346 , n430 , n229 );
    and g45 ( n325 , n386 , n198 );
    not g46 ( n345 , n248 );
    not g47 ( n153 , n507 );
    not g48 ( n368 , n478 );
    or g49 ( n20 , n536 , n337 );
    or g50 ( n87 , n519 , n298 );
    and g51 ( n65 , n33 , n507 );
    and g52 ( n191 , n390 , n152 );
    xnor g53 ( n296 , n144 , n188 );
    and g54 ( n214 , n209 , n279 );
    xnor g55 ( n144 , n498 , n90 );
    nor g56 ( n407 , n200 , n34 );
    or g57 ( n419 , n202 , n288 );
    nor g58 ( n260 , n197 , n254 );
    and g59 ( n69 , n375 , n238 );
    and g60 ( n342 , n343 , n509 );
    not g61 ( n416 , n98 );
    or g62 ( n100 , n252 , n206 );
    or g63 ( n483 , n73 , n538 );
    not g64 ( n66 , n59 );
    not g65 ( n212 , n524 );
    not g66 ( n477 , n220 );
    not g67 ( n25 , n410 );
    or g68 ( n77 , n236 , n438 );
    xnor g69 ( n429 , n480 , n234 );
    nor g70 ( n93 , n202 , n527 );
    nor g71 ( n1 , n441 , n303 );
    and g72 ( n312 , n83 , n461 );
    not g73 ( n426 , n79 );
    or g74 ( n24 , n403 , n530 );
    xnor g75 ( n478 , n155 , n220 );
    and g76 ( n146 , n134 , n225 );
    and g77 ( n299 , n263 , n376 );
    xor g78 ( n531 , n539 , n126 );
    nor g79 ( n510 , n354 , n415 );
    xnor g80 ( n226 , n319 , n240 );
    xnor g81 ( n281 , n426 , n348 );
    or g82 ( n189 , n425 , n414 );
    xnor g83 ( n488 , n100 , n98 );
    not g84 ( n84 , n543 );
    nor g85 ( n497 , n197 , n221 );
    not g86 ( n88 , n475 );
    and g87 ( n392 , n140 , n94 );
    and g88 ( n243 , n521 , n202 );
    or g89 ( n457 , n491 , n29 );
    nor g90 ( n437 , n433 , n177 );
    and g91 ( n515 , n433 , n177 );
    or g92 ( n210 , n290 , n46 );
    or g93 ( n62 , n147 , n210 );
    nor g94 ( n112 , n202 , n299 );
    or g95 ( n439 , n431 , n420 );
    and g96 ( n270 , n474 , n202 );
    or g97 ( n340 , n14 , n503 );
    and g98 ( n75 , n354 , n415 );
    not g99 ( n505 , n8 );
    xnor g100 ( n262 , n123 , n230 );
    nor g101 ( n362 , n202 , n39 );
    nor g102 ( n101 , n347 , n9 );
    not g103 ( n110 , n62 );
    and g104 ( n249 , n85 , n189 );
    nor g105 ( n135 , n340 , n53 );
    not g106 ( n119 , n245 );
    or g107 ( n365 , n289 , n393 );
    nor g108 ( n157 , n222 , n8 );
    nor g109 ( n17 , n338 , n472 );
    xnor g110 ( n514 , n375 , n182 );
    and g111 ( n479 , n506 , n89 );
    and g112 ( n167 , n171 , n170 );
    nor g113 ( n278 , n0 , n542 );
    and g114 ( n208 , n500 , n131 );
    or g115 ( n161 , n471 , n479 );
    not g116 ( n360 , n438 );
    and g117 ( n252 , n302 , n5 );
    or g118 ( n459 , n243 , n214 );
    xnor g119 ( n128 , n341 , n376 );
    not g120 ( n436 , n513 );
    nor g121 ( n393 , n242 , n233 );
    and g122 ( n206 , n301 , n498 );
    xnor g123 ( n338 , n540 , n58 );
    or g124 ( n136 , n271 , n178 );
    xnor g125 ( n162 , n15 , n368 );
    not g126 ( n288 , n77 );
    not g127 ( n469 , n116 );
    and g128 ( n277 , n331 , n202 );
    not g129 ( n15 , n39 );
    or g130 ( n319 , n312 , n203 );
    and g131 ( n130 , n478 , n104 );
    or g132 ( n92 , n156 , n93 );
    or g133 ( n535 , n341 , n101 );
    and g134 ( n336 , n398 , n209 );
    or g135 ( n297 , n202 , n427 );
    xnor g136 ( n39 , n524 , n79 );
    or g137 ( n219 , n473 , n18 );
    and g138 ( n447 , n64 , n153 );
    and g139 ( n38 , n41 , n327 );
    and g140 ( n163 , n144 , n283 );
    not g141 ( n107 , n487 );
    and g142 ( n473 , n349 , n202 );
    or g143 ( n307 , n150 , n197 );
    nor g144 ( n504 , n484 , n183 );
    not g145 ( n425 , n200 );
    and g146 ( n384 , n526 , n280 );
    or g147 ( n499 , n10 , n379 );
    or g148 ( n103 , n366 , n541 );
    nor g149 ( n154 , n191 , n192 );
    nor g150 ( n532 , n197 , n456 );
    not g151 ( n41 , n129 );
    and g152 ( n179 , n489 , n317 );
    and g153 ( n172 , n326 , n30 );
    or g154 ( n321 , n277 , n422 );
    and g155 ( n472 , n457 , n20 );
    or g156 ( n461 , n51 , n107 );
    not g157 ( n546 , n344 );
    xnor g158 ( n14 , n0 , n324 );
    or g159 ( n283 , n491 , n328 );
    and g160 ( n385 , n78 , n202 );
    not g161 ( n126 , n335 );
    and g162 ( n111 , n153 , n399 );
    and g163 ( n388 , n454 , n334 );
    or g164 ( n423 , n477 , n195 );
    or g165 ( n406 , n79 , n39 );
    or g166 ( n246 , n91 , n542 );
    xnor g167 ( n320 , n231 , n354 );
    or g168 ( n511 , n363 , n361 );
    not g169 ( n152 , n105 );
    xnor g170 ( n54 , n433 , n177 );
    not g171 ( n313 , n500 );
    and g172 ( n374 , n426 , n529 );
    xnor g173 ( n356 , n188 , n31 );
    nor g174 ( n82 , n171 , n345 );
    not g175 ( n458 , n94 );
    not g176 ( n137 , n97 );
    nor g177 ( n379 , n61 , n43 );
    not g178 ( n403 , n161 );
    xnor g179 ( n165 , n325 , n148 );
    not g180 ( n133 , n432 );
    xnor g181 ( n284 , n56 , n265 );
    nor g182 ( n16 , n197 , n514 );
    not g183 ( n267 , n396 );
    not g184 ( n518 , n540 );
    and g185 ( n314 , n358 , n445 );
    and g186 ( n187 , n136 , n535 );
    or g187 ( n371 , n497 , n13 );
    nor g188 ( n259 , n202 , n447 );
    xnor g189 ( n265 , n324 , n517 );
    or g190 ( n225 , n28 , n244 );
    nor g191 ( n536 , n188 , n31 );
    nor g192 ( n364 , n216 , n389 );
    xnor g193 ( n207 , n388 , n54 );
    not g194 ( n323 , n222 );
    or g195 ( n115 , n202 , n105 );
    not g196 ( n47 , n100 );
    or g197 ( n233 , n202 , n359 );
    or g198 ( n53 , n224 , n512 );
    or g199 ( n34 , n75 , n268 );
    nor g200 ( n408 , n197 , n132 );
    not g201 ( n29 , n31 );
    or g202 ( n489 , n309 , n449 );
    or g203 ( n60 , n44 , n124 );
    nor g204 ( n23 , n515 , n465 );
    or g205 ( n386 , n39 , n176 );
    xnor g206 ( n173 , n95 , n296 );
    or g207 ( n215 , n126 , n442 );
    nor g208 ( n363 , n467 , n65 );
    nor g209 ( n217 , n127 , n469 );
    or g210 ( n196 , n260 , n102 );
    and g211 ( n263 , n103 , n94 );
    or g212 ( n253 , n416 , n47 );
    and g213 ( n74 , n356 , n337 );
    or g214 ( n405 , n146 , n187 );
    buf g215 ( n37 , n426 );
    xor g216 ( n382 , n441 , n262 );
    and g217 ( n12 , n164 , n293 );
    not g218 ( n235 , n281 );
    and g219 ( n72 , n540 , n58 );
    and g220 ( n412 , n428 , n202 );
    or g221 ( n180 , n228 , n483 );
    or g222 ( n32 , n97 , n62 );
    xnor g223 ( n513 , n52 , n237 );
    and g224 ( n507 , n129 , n208 );
    and g225 ( n71 , n330 , n411 );
    not g226 ( n516 , n257 );
    or g227 ( n383 , n269 , n452 );
    or g228 ( n509 , n51 , n35 );
    nor g229 ( n160 , n272 , n472 );
    and g230 ( n30 , n151 , n19 );
    or g231 ( n169 , n323 , n382 );
    and g232 ( n105 , n321 , n359 );
    or g233 ( n7 , n539 , n455 );
    not g234 ( n4 , n261 );
    and g235 ( n142 , n145 , n202 );
    and g236 ( n422 , n333 , n501 );
    not g237 ( n174 , n46 );
    and g238 ( n359 , n161 , n288 );
    or g239 ( n151 , n526 , n280 );
    and g240 ( n397 , n144 , n96 );
    or g241 ( n192 , n202 , n57 );
    or g242 ( n68 , n478 , n526 );
    or g243 ( n304 , n202 , n229 );
    or g244 ( n330 , n531 , n30 );
    or g245 ( n290 , n270 , n372 );
    not g246 ( n83 , n488 );
    or g247 ( n454 , n84 , n522 );
    xnor g248 ( n45 , n528 , n162 );
    and g249 ( n442 , n280 , n534 );
    not g250 ( n434 , n433 );
    or g251 ( n56 , n119 , n546 );
    or g252 ( n185 , n408 , n106 );
    xnor g253 ( n318 , n469 , n207 );
    nor g254 ( n268 , n510 , n48 );
    not g255 ( n506 , n149 );
    and g256 ( n242 , n403 , n77 );
    nor g257 ( n417 , n202 , n407 );
    xnor g258 ( n237 , n99 , n60 );
    nor g259 ( n86 , n324 , n517 );
    and g260 ( n300 , n122 , n511 );
    xnor g261 ( n316 , n543 , n351 );
    xor g262 ( n402 , n15 , n284 );
    not g263 ( n275 , n189 );
    nor g264 ( n462 , n144 , n96 );
    or g265 ( n343 , n382 , n273 );
    and g266 ( n366 , n202 , n205 );
    not g267 ( n95 , n328 );
    not g268 ( n127 , n478 );
    and g269 ( n372 , n327 , n276 );
    xor g270 ( n503 , n144 , n543 );
    not g271 ( n209 , n159 );
    xnor g272 ( n255 , n475 , n451 );
    or g273 ( n334 , n141 , n179 );
    xor g274 ( n26 , n382 , n509 );
    and g275 ( n476 , n332 , n112 );
    buf g276 ( n250 , 1'b0 );
    not g277 ( n158 , n483 );
    xor g278 ( n482 , n144 , n36 );
    or g279 ( n421 , n227 , n163 );
    nor g280 ( n184 , n197 , n274 );
    not g281 ( n375 , n321 );
    or g282 ( n370 , n202 , n21 );
    not g283 ( n64 , n33 );
    and g284 ( n427 , n338 , n472 );
    or g285 ( n441 , n267 , n133 );
    and g286 ( n155 , n524 , n79 );
    nor g287 ( n76 , n114 , n264 );
    and g288 ( n138 , n389 , n259 );
    not g289 ( n80 , n442 );
    xnor g290 ( n104 , n179 , n316 );
    or g291 ( n339 , n51 , n235 );
    and g292 ( n131 , n380 , n159 );
    xnor g293 ( n27 , n352 , n440 );
    and g294 ( n61 , n73 , n538 );
    nor g295 ( n13 , n435 , n419 );
    not g296 ( n508 , n213 );
    nor g297 ( n446 , n202 , n82 );
    or g298 ( n19 , n384 , n413 );
    nor g299 ( n495 , n430 , n229 );
    not g300 ( n315 , n494 );
    and g301 ( n306 , n6 , n202 );
    not g302 ( n414 , n34 );
    not g303 ( n347 , n271 );
    xnor g304 ( n376 , n9 , n347 );
    and g305 ( n525 , n531 , n30 );
    and g306 ( n11 , n137 , n410 );
    not g307 ( n238 , n182 );
    or g308 ( n97 , n412 , n138 );
    not g309 ( n178 , n9 );
    not g310 ( n228 , n290 );
    xnor g311 ( n444 , n469 , n280 );
    not g312 ( n390 , n459 );
    xor g313 ( n452 , n231 , n40 );
    or g314 ( n286 , n193 , n537 );
    not g315 ( n389 , n65 );
    and g316 ( n18 , n189 , n417 );
    or g317 ( n171 , n285 , n516 );
    not g318 ( n285 , n451 );
    nor g319 ( n10 , n197 , n485 );
    or g320 ( n492 , n518 , n421 );
    nor g321 ( n156 , n197 , n377 );
    and g322 ( n229 , n97 , n25 );
    or g323 ( n394 , n323 , n505 );
    not g324 ( n387 , n210 );
    and g325 ( n539 , n502 , n294 );
    or g326 ( n440 , n539 , n469 );
    or g327 ( n261 , n459 , n117 );
    nor g328 ( n124 , n207 , n493 );
    not g329 ( n327 , n208 );
    xnor g330 ( n248 , n323 , n8 );
    and g331 ( n453 , n508 , n333 );
    nor g332 ( n3 , n15 , n374 );
    and g333 ( n485 , n308 , n46 );
    nor g334 ( n141 , n543 , n351 );
    not g335 ( n195 , n155 );
    nor g336 ( n298 , n55 , n370 );
    xnor g337 ( n166 , n0 , n222 );
    xnor g338 ( n475 , n396 , n432 );
    xnor g339 ( n125 , n368 , n146 );
    or g340 ( n232 , n367 , n71 );
    and g341 ( n542 , n475 , n199 );
    not g342 ( n449 , n517 );
    or g343 ( n147 , n142 , n111 );
    not g344 ( n0 , n382 );
    and g345 ( n256 , n375 , n120 );
    nor g346 ( n269 , n434 , n83 );
    and g347 ( n352 , n68 , n194 );
    not g348 ( n413 , n211 );
    and g349 ( n63 , n202 , n204 );
    or g350 ( n282 , n368 , n193 );
    or g351 ( n445 , n72 , n160 );
    and g352 ( n114 , n518 , n421 );
    xnor g353 ( n377 , n280 , n286 );
    and g354 ( n203 , n109 , n42 );
    not g355 ( n216 , n467 );
    and g356 ( n544 , n9 , n22 );
    and g357 ( n149 , n357 , n275 );
    not g358 ( n468 , n147 );
    and g359 ( n266 , n123 , n230 );
    nor g360 ( n305 , n222 , n0 );
    xnor g361 ( n254 , n97 , n110 );
    not g362 ( n247 , n400 );
    or g363 ( n332 , n263 , n376 );
    and g364 ( n409 , n313 , n164 );
    xnor g365 ( n90 , n302 , n5 );
    and g366 ( n132 , n405 , n286 );
    or g367 ( n183 , n202 , n25 );
    and g368 ( n264 , n83 , n492 );
    nor g369 ( n276 , n202 , n409 );
    nor g370 ( n279 , n202 , n453 );
    nor g371 ( n102 , n11 , n304 );
    and g372 ( n36 , n201 , n165 );
    nor g373 ( n106 , n202 , n486 );
    nor g374 ( n411 , n202 , n525 );
    and g375 ( n545 , n49 , n202 );
    or g376 ( n373 , n184 , n504 );
    or g377 ( n70 , n186 , n248 );
    not g378 ( n430 , n300 );
    not g379 ( n150 , n251 );
    or g380 ( n168 , n16 , n139 );
    not g381 ( n273 , n542 );
    xnor g382 ( n481 , n354 , n415 );
    and g383 ( n355 , n127 , n193 );
    not g384 ( n120 , n359 );
    not g385 ( n176 , n374 );
    xnor g386 ( n99 , n40 , n181 );
    or g387 ( n498 , n266 , n1 );
    or g388 ( n59 , n335 , n80 );
    nor g389 ( n399 , n202 , n38 );
    and g390 ( n67 , n70 , n446 );
    and g391 ( n460 , n24 , n182 );
    or g392 ( n94 , n463 , n167 );
    not g393 ( n48 , n445 );
    xnor g394 ( n143 , n295 , n166 );
    or g395 ( n109 , n83 , n461 );
    not g396 ( n529 , n348 );
    or g397 ( n96 , n278 , n342 );
    not g398 ( n530 , n448 );
    or g399 ( n198 , n3 , n284 );
    nor g400 ( n223 , n197 , n128 );
    or g401 ( n295 , n285 , n88 );
    and g402 ( n241 , n400 , n149 );
    xnor g403 ( n52 , n326 , n23 );
    not g404 ( n418 , n2 );
    or g405 ( n182 , n161 , n448 );
    xnor g406 ( n527 , n211 , n444 );
    not g407 ( n35 , n381 );
    or g408 ( n292 , n17 , n297 );
    xnor g409 ( n466 , n83 , n518 );
    not g410 ( n164 , n131 );
    and g411 ( n337 , n394 , n470 );
    nor g412 ( n310 , n462 , n36 );
    or g413 ( n311 , n545 , n12 );
    and g414 ( n471 , n287 , n202 );
    or g415 ( n271 , n63 , n362 );
    nor g416 ( n28 , n356 , n337 );
    or g417 ( n438 , n126 , n172 );
    not g418 ( n537 , n187 );
    nor g419 ( n367 , n197 , n353 );
    xor g420 ( n116 , n423 , n502 );
    not g421 ( n57 , n538 );
    or g422 ( n190 , n39 , n478 );
    not g423 ( n186 , n171 );
    not g424 ( n522 , n351 );
    or g425 ( n361 , n202 , n364 );
    or g426 ( n378 , n476 , n223 );
    xnor g427 ( n404 , n542 , n26 );
    or g428 ( n410 , n468 , n180 );
    xor g429 ( n456 , n390 , n69 );
    nor g430 ( n431 , n197 , n496 );
    or g431 ( n538 , n390 , n152 );
    not g432 ( n117 , n69 );
    or g433 ( n350 , n532 , n154 );
    not g434 ( n528 , n406 );
    xnor g435 ( n231 , n253 , n523 );
    and g436 ( n493 , n526 , n520 );
    nor g437 ( n291 , n451 , n257 );
    xnor g438 ( n381 , n374 , n402 );
    or g439 ( n322 , n202 , n495 );
    not g440 ( n51 , n201 );
    or g441 ( n512 , n424 , n383 );
    not g442 ( n199 , n339 );
    xnor g443 ( n224 , n475 , n245 );
    and g444 ( n443 , n295 , n169 );
    or g445 ( n244 , n202 , n74 );
    nor g446 ( n420 , n346 , n322 );
    or g447 ( n328 , n305 , n443 );
    or g448 ( n42 , n397 , n310 );
    and g449 ( n520 , n329 , n118 );
    not g450 ( n73 , n311 );
    or g451 ( n81 , n202 , n464 );
    not g452 ( n309 , n324 );
    nor g453 ( n435 , n219 , n360 );
    xor g454 ( n50 , n228 , n174 );
    xnor g455 ( n148 , n127 , n104 );
    or g456 ( n118 , n130 , n325 );
    nor g457 ( n519 , n197 , n50 );
    or g458 ( n122 , n315 , n197 );
    not g459 ( n333 , n241 );
    not g460 ( n140 , n103 );
    or g461 ( n134 , n418 , n197 );
    nor g462 ( n501 , n202 , n175 );
    not g463 ( n236 , n219 );
    nor g464 ( n44 , n526 , n520 );
    xnor g465 ( n490 , n42 , n239 );
    or g466 ( n43 , n202 , n158 );
    nor g467 ( n289 , n197 , n460 );
    nor g468 ( n455 , n526 , n352 );
    xnor g469 ( n487 , n520 , n318 );
    not g470 ( n358 , n481 );
    and g471 ( n91 , n88 , n339 );
    not g472 ( n197 , n202 );
    or g473 ( n258 , n392 , n341 );
    nor g474 ( n139 , n256 , n115 );
    not g475 ( n85 , n357 );
    nor g476 ( n89 , n202 , n249 );
    and g477 ( n395 , n282 , n218 );
    or g478 ( n317 , n56 , n86 );
    or g479 ( n470 , n171 , n157 );
    or g480 ( n211 , n355 , n395 );
    nor g481 ( n303 , n123 , n230 );
    not g482 ( n398 , n380 );
    and g483 ( n175 , n247 , n506 );
    or g484 ( n301 , n302 , n5 );
    or g485 ( n22 , n271 , n263 );
    and g486 ( n463 , n533 , n202 );
    or g487 ( n9 , n385 , n67 );
endmodule
