module top( n11 , n21 , n22 , n23 , n27 , n29 , n30 , n40 , n45 , 
n50 , n52 , n54 , n56 , n58 , n71 , n77 , n82 , n85 , n86 , 
n87 , n94 , n107 , n112 , n117 , n126 , n130 , n138 , n143 , n153 , 
n155 , n156 , n159 , n161 , n164 , n173 , n181 , n184 , n200 , n216 , 
n219 , n220 , n222 , n223 , n230 , n233 , n243 , n244 , n246 , n247 , 
n251 , n254 , n262 , n268 , n273 , n275 , n284 , n288 , n292 , n293 , 
n299 , n300 , n301 , n304 , n307 , n310 , n312 , n314 , n315 , n318 , 
n337 , n341 , n344 , n346 , n352 , n362 , n364 , n370 , n374 , n376 , 
n378 , n380 , n391 , n392 , n396 , n399 , n408 , n409 , n416 , n417 , 
n420 , n428 , n430 , n453 , n457 , n460 , n477 , n478 , n487 , n489 , 
n497 , n498 , n501 , n502 , n506 , n507 , n509 , n510 , n516 , n517 , 
n534 , n545 , n553 , n559 , n560 , n561 , n567 , n574 , n581 , n582 , 
n585 , n589 , n593 , n595 , n597 , n598 , n600 , n607 , n608 , n609 , 
n625 , n626 , n638 , n640 , n641 , n645 , n663 , n669 , n671 , n676 , 
n690 , n693 , n695 , n701 , n710 , n714 , n719 , n726 , n727 , n729 , 
n734 , n742 , n743 , n755 , n769 , n773 , n775 , n778 , n779 , n782 , 
n787 , n790 , n794 , n821 , n823 , n831 , n832 , n839 , n842 , n849 , 
n879 , n882 , n885 , n894 , n905 , n916 , n918 , n920 , n936 , n947 , 
n952 , n953 , n961 , n969 , n980 , n984 , n986 , n990 , n992 , n997 , 
n1006 , n1017 , n1023 , n1040 , n1042 , n1044 , n1050 , n1051 , n1054 , n1058 , 
n1060 , n1061 , n1063 , n1065 , n1071 , n1095 , n1103 , n1114 , n1121 , n1138 , 
n1152 , n1154 , n1156 , n1164 , n1172 , n1175 , n1177 , n1186 , n1187 , n1191 , 
n1193 , n1195 , n1205 , n1209 , n1211 , n1225 , n1227 , n1231 , n1234 , n1239 , 
n1246 , n1250 , n1253 , n1263 , n1278 , n1281 , n1283 , n1285 , n1286 , n1288 , 
n1289 , n1292 , n1296 , n1299 , n1301 , n1302 , n1305 , n1306 , n1320 , n1322 , 
n1337 , n1345 , n1346 , n1350 , n1359 , n1361 , n1368 , n1375 , n1386 , n1387 , 
n1389 , n1391 , n1393 , n1401 , n1411 , n1415 , n1418 , n1420 , n1421 , n1427 , 
n1428 , n1435 , n1438 , n1443 , n1446 , n1448 , n1463 , n1470 , n1474 , n1476 , 
n1500 , n1502 , n1506 , n1516 , n1520 , n1521 , n1523 , n1527 , n1534 , n1536 , 
n1547 , n1548 , n1566 , n1569 , n1576 , n1586 , n1588 , n1592 , n1594 , n1609 , 
n1613 , n1616 , n1626 , n1627 , n1632 , n1639 , n1644 , n1645 , n1647 , n1656 , 
n1687 , n1729 , n1738 , n1750 , n1752 , n1753 );
    input n11 , n21 , n29 , n40 , n45 , n50 , n52 , n54 , n56 , 
n58 , n71 , n77 , n82 , n86 , n87 , n94 , n107 , n117 , n138 , 
n143 , n153 , n155 , n156 , n159 , n200 , n219 , n220 , n222 , n223 , 
n243 , n244 , n246 , n251 , n254 , n262 , n268 , n273 , n284 , n288 , 
n293 , n299 , n300 , n307 , n310 , n312 , n314 , n315 , n318 , n341 , 
n344 , n346 , n374 , n376 , n380 , n391 , n392 , n399 , n408 , n409 , 
n416 , n420 , n430 , n477 , n478 , n487 , n489 , n502 , n506 , n507 , 
n510 , n545 , n559 , n560 , n561 , n567 , n574 , n581 , n582 , n589 , 
n593 , n598 , n600 , n607 , n608 , n609 , n626 , n641 , n645 , n663 , 
n671 , n676 , n690 , n695 , n701 , n710 , n727 , n729 , n734 , n742 , 
n743 , n755 , n769 , n775 , n778 , n779 , n787 , n790 , n823 , n831 , 
n832 , n839 , n849 , n879 , n882 , n885 , n905 , n920 , n936 , n947 , 
n953 , n961 , n969 , n980 , n984 , n986 , n992 , n997 , n1023 , n1040 , 
n1044 , n1054 , n1061 , n1071 , n1095 , n1103 , n1114 , n1121 , n1138 , n1152 , 
n1154 , n1156 , n1164 , n1172 , n1175 , n1187 , n1191 , n1193 , n1205 , n1225 , 
n1227 , n1239 , n1246 , n1250 , n1263 , n1278 , n1281 , n1283 , n1286 , n1289 , 
n1299 , n1301 , n1305 , n1345 , n1346 , n1350 , n1361 , n1386 , n1387 , n1389 , 
n1393 , n1401 , n1411 , n1415 , n1418 , n1428 , n1435 , n1438 , n1443 , n1446 , 
n1448 , n1463 , n1470 , n1474 , n1476 , n1500 , n1502 , n1506 , n1516 , n1520 , 
n1521 , n1523 , n1536 , n1566 , n1569 , n1576 , n1586 , n1592 , n1609 , n1613 , 
n1616 , n1626 , n1627 , n1644 , n1647 , n1656 , n1750 , n1753 ;
    output n22 , n23 , n27 , n30 , n85 , n112 , n126 , n130 , n161 , 
n164 , n173 , n181 , n184 , n216 , n230 , n233 , n247 , n275 , n292 , 
n301 , n304 , n337 , n352 , n362 , n364 , n370 , n378 , n396 , n417 , 
n428 , n453 , n457 , n460 , n497 , n498 , n501 , n509 , n516 , n517 , 
n534 , n553 , n585 , n595 , n597 , n625 , n638 , n640 , n669 , n693 , 
n714 , n719 , n726 , n773 , n782 , n794 , n821 , n842 , n894 , n916 , 
n918 , n952 , n990 , n1006 , n1017 , n1042 , n1050 , n1051 , n1058 , n1060 , 
n1063 , n1065 , n1177 , n1186 , n1195 , n1209 , n1211 , n1231 , n1234 , n1253 , 
n1285 , n1288 , n1292 , n1296 , n1302 , n1306 , n1320 , n1322 , n1337 , n1359 , 
n1368 , n1375 , n1391 , n1420 , n1421 , n1427 , n1527 , n1534 , n1547 , n1548 , 
n1588 , n1594 , n1632 , n1639 , n1645 , n1687 , n1729 , n1738 , n1752 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , 
n9 , n10 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
n20 , n24 , n25 , n26 , n28 , n31 , n32 , n33 , n34 , n35 , 
n36 , n37 , n38 , n39 , n41 , n42 , n43 , n44 , n46 , n47 , 
n48 , n49 , n51 , n53 , n55 , n57 , n59 , n60 , n61 , n62 , 
n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n72 , n73 , 
n74 , n75 , n76 , n78 , n79 , n80 , n81 , n83 , n84 , n88 , 
n89 , n90 , n91 , n92 , n93 , n95 , n96 , n97 , n98 , n99 , 
n100 , n101 , n102 , n103 , n104 , n105 , n106 , n108 , n109 , n110 , 
n111 , n113 , n114 , n115 , n116 , n118 , n119 , n120 , n121 , n122 , 
n123 , n124 , n125 , n127 , n128 , n129 , n131 , n132 , n133 , n134 , 
n135 , n136 , n137 , n139 , n140 , n141 , n142 , n144 , n145 , n146 , 
n147 , n148 , n149 , n150 , n151 , n152 , n154 , n157 , n158 , n160 , 
n162 , n163 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , 
n174 , n175 , n176 , n177 , n178 , n179 , n180 , n182 , n183 , n185 , 
n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , 
n196 , n197 , n198 , n199 , n201 , n202 , n203 , n204 , n205 , n206 , 
n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n217 , 
n218 , n221 , n224 , n225 , n226 , n227 , n228 , n229 , n231 , n232 , 
n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n245 , 
n248 , n249 , n250 , n252 , n253 , n255 , n256 , n257 , n258 , n259 , 
n260 , n261 , n263 , n264 , n265 , n266 , n267 , n269 , n270 , n271 , 
n272 , n274 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , 
n285 , n286 , n287 , n289 , n290 , n291 , n294 , n295 , n296 , n297 , 
n298 , n302 , n303 , n305 , n306 , n308 , n309 , n311 , n313 , n316 , 
n317 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , 
n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n338 , 
n339 , n340 , n342 , n343 , n345 , n347 , n348 , n349 , n350 , n351 , 
n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n363 , 
n365 , n366 , n367 , n368 , n369 , n371 , n372 , n373 , n375 , n377 , 
n379 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
n390 , n393 , n394 , n395 , n397 , n398 , n400 , n401 , n402 , n403 , 
n404 , n405 , n406 , n407 , n410 , n411 , n412 , n413 , n414 , n415 , 
n418 , n419 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n429 , 
n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , 
n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , 
n451 , n452 , n454 , n455 , n456 , n458 , n459 , n461 , n462 , n463 , 
n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , 
n474 , n475 , n476 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , 
n486 , n488 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n499 , 
n500 , n503 , n504 , n505 , n508 , n511 , n512 , n513 , n514 , n515 , 
n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , 
n528 , n529 , n530 , n531 , n532 , n533 , n535 , n536 , n537 , n538 , 
n539 , n540 , n541 , n542 , n543 , n544 , n546 , n547 , n548 , n549 , 
n550 , n551 , n552 , n554 , n555 , n556 , n557 , n558 , n562 , n563 , 
n564 , n565 , n566 , n568 , n569 , n570 , n571 , n572 , n573 , n575 , 
n576 , n577 , n578 , n579 , n580 , n583 , n584 , n586 , n587 , n588 , 
n590 , n591 , n592 , n594 , n596 , n599 , n601 , n602 , n603 , n604 , 
n605 , n606 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , 
n618 , n619 , n620 , n621 , n622 , n623 , n624 , n627 , n628 , n629 , 
n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n639 , n642 , 
n643 , n644 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , 
n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n664 , 
n665 , n666 , n667 , n668 , n670 , n672 , n673 , n674 , n675 , n677 , 
n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , 
n688 , n689 , n691 , n692 , n694 , n696 , n697 , n698 , n699 , n700 , 
n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n711 , n712 , 
n713 , n715 , n716 , n717 , n718 , n720 , n721 , n722 , n723 , n724 , 
n725 , n728 , n730 , n731 , n732 , n733 , n735 , n736 , n737 , n738 , 
n739 , n740 , n741 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , 
n751 , n752 , n753 , n754 , n756 , n757 , n758 , n759 , n760 , n761 , 
n762 , n763 , n764 , n765 , n766 , n767 , n768 , n770 , n771 , n772 , 
n774 , n776 , n777 , n780 , n781 , n783 , n784 , n785 , n786 , n788 , 
n789 , n791 , n792 , n793 , n795 , n796 , n797 , n798 , n799 , n800 , 
n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , 
n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , 
n822 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n833 , n834 , 
n835 , n836 , n837 , n838 , n840 , n841 , n843 , n844 , n845 , n846 , 
n847 , n848 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , 
n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , 
n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , 
n878 , n880 , n881 , n883 , n884 , n886 , n887 , n888 , n889 , n890 , 
n891 , n892 , n893 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , 
n902 , n903 , n904 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , 
n913 , n914 , n915 , n917 , n919 , n921 , n922 , n923 , n924 , n925 , 
n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , 
n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , 
n948 , n949 , n950 , n951 , n954 , n955 , n956 , n957 , n958 , n959 , 
n960 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n970 , n971 , 
n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n981 , n982 , 
n983 , n985 , n987 , n988 , n989 , n991 , n993 , n994 , n995 , n996 , 
n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1007 , n1008 , 
n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1018 , n1019 , 
n1020 , n1021 , n1022 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , 
n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1041 , 
n1043 , n1045 , n1046 , n1047 , n1048 , n1049 , n1052 , n1053 , n1055 , n1056 , 
n1057 , n1059 , n1062 , n1064 , n1066 , n1067 , n1068 , n1069 , n1070 , n1072 , 
n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , 
n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , 
n1093 , n1094 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1104 , 
n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1115 , 
n1116 , n1117 , n1118 , n1119 , n1120 , n1122 , n1123 , n1124 , n1125 , n1126 , 
n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , 
n1137 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , 
n1148 , n1149 , n1150 , n1151 , n1153 , n1155 , n1157 , n1158 , n1159 , n1160 , 
n1161 , n1162 , n1163 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , 
n1173 , n1174 , n1176 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , 
n1185 , n1188 , n1189 , n1190 , n1192 , n1194 , n1196 , n1197 , n1198 , n1199 , 
n1200 , n1201 , n1202 , n1203 , n1204 , n1206 , n1207 , n1208 , n1210 , n1212 , 
n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , 
n1223 , n1224 , n1226 , n1228 , n1229 , n1230 , n1232 , n1233 , n1235 , n1236 , 
n1237 , n1238 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1247 , n1248 , 
n1249 , n1251 , n1252 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , 
n1261 , n1262 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , 
n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1279 , n1280 , n1282 , n1284 , 
n1287 , n1290 , n1291 , n1293 , n1294 , n1295 , n1297 , n1298 , n1300 , n1303 , 
n1304 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , 
n1316 , n1317 , n1318 , n1319 , n1321 , n1323 , n1324 , n1325 , n1326 , n1327 , 
n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1338 , 
n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1347 , n1348 , n1349 , n1351 , 
n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1360 , n1362 , n1363 , 
n1364 , n1365 , n1366 , n1367 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , 
n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , 
n1388 , n1390 , n1392 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , 
n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1412 , 
n1413 , n1414 , n1416 , n1417 , n1419 , n1422 , n1423 , n1424 , n1425 , n1426 , 
n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1436 , n1437 , n1439 , n1440 , 
n1441 , n1442 , n1444 , n1445 , n1447 , n1449 , n1450 , n1451 , n1452 , n1453 , 
n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1464 , 
n1465 , n1466 , n1467 , n1468 , n1469 , n1471 , n1472 , n1473 , n1475 , n1477 , 
n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , 
n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , 
n1498 , n1499 , n1501 , n1503 , n1504 , n1505 , n1507 , n1508 , n1509 , n1510 , 
n1511 , n1512 , n1513 , n1514 , n1515 , n1517 , n1518 , n1519 , n1522 , n1524 , 
n1525 , n1526 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1535 , n1537 , 
n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1549 , 
n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1567 , n1568 , n1570 , n1571 , 
n1572 , n1573 , n1574 , n1575 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , 
n1583 , n1584 , n1585 , n1587 , n1589 , n1590 , n1591 , n1593 , n1595 , n1596 , 
n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , 
n1607 , n1608 , n1610 , n1611 , n1612 , n1614 , n1615 , n1617 , n1618 , n1619 , 
n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1628 , n1629 , n1630 , n1631 , 
n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1640 , n1641 , n1642 , n1643 , 
n1646 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1657 , 
n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , 
n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , 
n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1688 , 
n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , 
n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , 
n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , 
n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , 
n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1739 , n1740 , 
n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1751 , 
n1754 , n1755 , n1756 ;
    or g0 ( n426 , n422 , n1543 );
    or g1 ( n1664 , n889 , n1101 );
    xnor g2 ( n1637 , n456 , n1142 );
    xnor g3 ( n1067 , n1402 , n145 );
    xnor g4 ( n993 , n780 , n1263 );
    xor g5 ( n1517 , n206 , n1725 );
    or g6 ( n1735 , n1116 , n1429 );
    and g7 ( n1539 , n1683 , n1276 );
    not g8 ( n154 , n1002 );
    nor g9 ( n1347 , n142 , n1105 );
    not g10 ( n1537 , n1540 );
    xnor g11 ( n1608 , n1573 , n866 );
    not g12 ( n960 , n1377 );
    and g13 ( n476 , n768 , n1126 );
    or g14 ( n805 , n1485 , n192 );
    xnor g15 ( n752 , n88 , n540 );
    not g16 ( n1048 , n654 );
    nor g17 ( n1698 , n1343 , n109 );
    nor g18 ( n1326 , n289 , n1230 );
    not g19 ( n721 , n728 );
    not g20 ( n1555 , n886 );
    or g21 ( n1578 , n1194 , n25 );
    or g22 ( n1383 , n802 , n218 );
    buf g23 ( n821 , n374 );
    not g24 ( n802 , n837 );
    or g25 ( n103 , n1706 , n1557 );
    or g26 ( n175 , n717 , n943 );
    not g27 ( n468 , n1419 );
    xnor g28 ( n38 , n1207 , n557 );
    or g29 ( n1585 , n1115 , n238 );
    or g30 ( n1105 , n1416 , n467 );
    or g31 ( n1648 , n935 , n266 );
    not g32 ( n165 , n1664 );
    or g33 ( n212 , n1721 , n500 );
    and g34 ( n624 , n885 , n197 );
    and g35 ( n1218 , n986 , n0 );
    or g36 ( n1002 , n228 , n1551 );
    or g37 ( n256 , n1357 , n1533 );
    or g38 ( n102 , n1531 , n686 );
    xnor g39 ( n1617 , n1373 , n1417 );
    xnor g40 ( n123 , n1512 , n1355 );
    and g41 ( n272 , n1100 , n177 );
    or g42 ( n305 , n1481 , n272 );
    nor g43 ( n104 , n721 , n1401 );
    or g44 ( n973 , n1408 , n379 );
    not g45 ( n70 , n923 );
    not g46 ( n1365 , n1506 );
    xnor g47 ( n1316 , n632 , n1595 );
    and g48 ( n1015 , n376 , n1168 );
    xnor g49 ( n1302 , n837 , n933 );
    and g50 ( n1480 , n779 , n721 );
    and g51 ( n1719 , n251 , n1555 );
    or g52 ( n1188 , n1268 , n1458 );
    nor g53 ( n148 , n721 , n1138 );
    xnor g54 ( n436 , n777 , n194 );
    xnor g55 ( n1247 , n1037 , n72 );
    not g56 ( n747 , n1708 );
    not g57 ( n579 , n1293 );
    xnor g58 ( n1556 , n723 , n518 );
    and g59 ( n471 , n1558 , n1312 );
    not g60 ( n327 , n843 );
    not g61 ( n846 , n324 );
    xnor g62 ( n1488 , n623 , n1382 );
    nand g63 ( n1237 , n380 , n701 );
    and g64 ( n785 , n63 , n807 );
    and g65 ( n1370 , n559 , n491 );
    not g66 ( n388 , n1559 );
    or g67 ( n658 , n1696 , n835 );
    not g68 ( n914 , n1387 );
    xnor g69 ( n331 , n1107 , n1707 );
    xnor g70 ( n1212 , n999 , n24 );
    not g71 ( n1623 , n891 );
    nor g72 ( n488 , n1535 , n1628 );
    and g73 ( n681 , n1172 , n602 );
    buf g74 ( n1017 , n1476 );
    not g75 ( n298 , n1521 );
    and g76 ( n923 , n1692 , n474 );
    not g77 ( n670 , n626 );
    and g78 ( n554 , n134 , n1400 );
    not g79 ( n1515 , n1008 );
    or g80 ( n1325 , n1579 , n423 );
    or g81 ( n1201 , n1623 , n1511 );
    nor g82 ( n549 , n63 , n32 );
    or g83 ( n1158 , n1241 , n1354 );
    not g84 ( n197 , n1314 );
    or g85 ( n861 , n64 , n1244 );
    nor g86 ( n801 , n1615 , n1336 );
    and g87 ( n151 , n312 , n1458 );
    buf g88 ( n516 , n1187 );
    and g89 ( n1075 , n124 , n1482 );
    or g90 ( n946 , n568 , n999 );
    xnor g91 ( n1525 , n1339 , n615 );
    nor g92 ( n587 , n1734 , n772 );
    not g93 ( n1179 , n545 );
    nor g94 ( n686 , n1178 , n175 );
    or g95 ( n1465 , n1254 , n1167 );
    and g96 ( n1477 , n89 , n495 );
    or g97 ( n1687 , n523 , n73 );
    or g98 ( n1538 , n1013 , n444 );
    not g99 ( n1355 , n188 );
    or g100 ( n1736 , n687 , n979 );
    nor g101 ( n1119 , n257 , n200 );
    not g102 ( n26 , n778 );
    xnor g103 ( n1714 , n1445 , n1084 );
    or g104 ( n1658 , n1261 , n10 );
    and g105 ( n1596 , n1393 , n530 );
    not g106 ( n1673 , n993 );
    or g107 ( n1743 , n359 , n434 );
    nor g108 ( n1335 , n1686 , n1073 );
    nor g109 ( n1612 , n721 , n56 );
    not g110 ( n1458 , n808 );
    and g111 ( n182 , n1346 , n602 );
    xnor g112 ( n1468 , n1597 , n980 );
    and g113 ( n195 , n1251 , n1598 );
    xnor g114 ( n1307 , n1273 , n427 );
    xnor g115 ( n324 , n1721 , n732 );
    or g116 ( n828 , n1752 , n493 );
    and g117 ( n958 , n1673 , n798 );
    buf g118 ( n301 , n318 );
    not g119 ( n316 , n1201 );
    xnor g120 ( n174 , n1597 , n923 );
    not g121 ( n119 , n567 );
    and g122 ( n124 , n395 , n1034 );
    buf g123 ( n460 , n21 );
    xnor g124 ( n1496 , n1049 , n630 );
    not g125 ( n1214 , n339 );
    xnor g126 ( n504 , n49 , n1406 );
    xnor g127 ( n1107 , n83 , n724 );
    not g128 ( n811 , n1475 );
    and g129 ( n1189 , n2 , n323 );
    not g130 ( n17 , n865 );
    or g131 ( n474 , n803 , n905 );
    xnor g132 ( n1084 , n1648 , n1018 );
    xnor g133 ( n1287 , n261 , n1727 );
    nor g134 ( n252 , n522 , n132 );
    and g135 ( n760 , n1230 , n873 );
    or g136 ( n1497 , n721 , n346 );
    xnor g137 ( n606 , n1537 , n60 );
    or g138 ( n481 , n1182 , n1238 );
    or g139 ( n306 , n1577 , n1203 );
    xnor g140 ( n99 , n1535 , n1442 );
    or g141 ( n35 , n636 , n1620 );
    not g142 ( n1394 , n1681 );
    or g143 ( n1099 , n1489 , n806 );
    or g144 ( n1306 , n1204 , n1619 );
    xnor g145 ( n302 , n1173 , n608 );
    xnor g146 ( n1600 , n32 , n1473 );
    not g147 ( n308 , n1239 );
    xnor g148 ( n611 , n1166 , n1699 );
    xnor g149 ( n1058 , n1667 , n810 );
    not g150 ( n687 , n1711 );
    not g151 ( n1430 , n307 );
    nor g152 ( n414 , n1470 , n910 );
    not g153 ( n1511 , n907 );
    and g154 ( n340 , n613 , n698 );
    and g155 ( n1621 , n934 , n1697 );
    nor g156 ( n1532 , n1667 , n840 );
    xor g157 ( n1404 , n133 , n375 );
    and g158 ( n921 , n1644 , n1136 );
    not g159 ( n835 , n413 );
    not g160 ( n1395 , n738 );
    xnor g161 ( n1072 , n899 , n938 );
    nor g162 ( n492 , n900 , n86 );
    and g163 ( n637 , n1672 , n1475 );
    xor g164 ( n213 , n142 , n1083 );
    nor g165 ( n1269 , n999 , n703 );
    not g166 ( n999 , n1419 );
    xnor g167 ( n373 , n740 , n407 );
    or g168 ( n1170 , n903 , n694 );
    and g169 ( n271 , n1750 , n238 );
    nor g170 ( n177 , n1230 , n1335 );
    xnor g171 ( n1689 , n1200 , n707 );
    or g172 ( n1282 , n454 , n639 );
    or g173 ( n1235 , n1722 , n649 );
    not g174 ( n900 , n413 );
    or g175 ( n1747 , n1102 , n75 );
    or g176 ( n1148 , n798 , n1390 );
    or g177 ( n96 , n687 , n1139 );
    and g178 ( n140 , n651 , n248 );
    nor g179 ( n1194 , n1099 , n189 );
    or g180 ( n635 , n1668 , n197 );
    and g181 ( n137 , n1415 , n530 );
    and g182 ( n1018 , n479 , n840 );
    not g183 ( n530 , n808 );
    and g184 ( n1085 , n899 , n1264 );
    or g185 ( n1162 , n803 , n1191 );
    nor g186 ( n357 , n367 , n158 );
    or g187 ( n91 , n985 , n443 );
    or g188 ( n1083 , n1015 , n804 );
    xnor g189 ( n1091 , n876 , n33 );
    and g190 ( n367 , n1360 , n575 );
    or g191 ( n1274 , n1698 , n1075 );
    or g192 ( n379 , n964 , n717 );
    xnor g193 ( n1229 , n922 , n1651 );
    not g194 ( n1126 , n852 );
    not g195 ( n1197 , n179 );
    xnor g196 ( n962 , n1686 , n1498 );
    and g197 ( n47 , n1083 , n1492 );
    not g198 ( n1113 , n1188 );
    xnor g199 ( n1457 , n206 , n1343 );
    or g200 ( n1155 , n1405 , n567 );
    xnor g201 ( n866 , n654 , n1629 );
    or g202 ( n1353 , n204 , n577 );
    or g203 ( n537 , n1291 , n1098 );
    or g204 ( n1618 , n761 , n465 );
    and g205 ( n1397 , n219 , n1168 );
    not g206 ( n758 , n565 );
    xnor g207 ( n1582 , n1641 , n1476 );
    nor g208 ( n1272 , n146 , n481 );
    or g209 ( n592 , n760 , n1327 );
    and g210 ( n1226 , n1585 , n569 );
    or g211 ( n1642 , n1561 , n250 );
    xnor g212 ( n1380 , n1573 , n1133 );
    nor g213 ( n1132 , n324 , n241 );
    not g214 ( n1135 , n888 );
    or g215 ( n746 , n1493 , n503 );
    buf g216 ( n1320 , n1263 );
    nor g217 ( n100 , n354 , n1137 );
    xnor g218 ( n1009 , n1340 , n1636 );
    not g219 ( n259 , n908 );
    or g220 ( n719 , n1361 , n1225 );
    nor g221 ( n245 , n803 , n769 );
    or g222 ( n486 , n614 , n1012 );
    nor g223 ( n1604 , n572 , n1682 );
    xnor g224 ( n525 , n1673 , n1148 );
    xnor g225 ( n1056 , n555 , n730 );
    not g226 ( n9 , n1284 );
    buf g227 ( n1738 , n45 );
    or g228 ( n718 , n629 , n636 );
    or g229 ( n266 , n1552 , n1222 );
    or g230 ( n120 , n1288 , n1322 );
    or g231 ( n807 , n1136 , n1435 );
    not g232 ( n1565 , n1747 );
    xor g233 ( n812 , n1623 , n907 );
    nor g234 ( n874 , n1535 , n1695 );
    or g235 ( n1190 , n695 , n653 );
    nor g236 ( n646 , n852 , n1436 );
    or g237 ( n1133 , n883 , n1048 );
    or g238 ( n229 , n793 , n59 );
    xnor g239 ( n383 , n948 , n1148 );
    and g240 ( n1709 , n849 , n776 );
    or g241 ( n1358 , n1700 , n212 );
    nor g242 ( n1215 , n1601 , n998 );
    not g243 ( n348 , n1307 );
    not g244 ( n731 , n1694 );
    or g245 ( n1716 , n1304 , n333 );
    and g246 ( n798 , n249 , n1129 );
    not g247 ( n1381 , n1043 );
    not g248 ( n1493 , n225 );
    not g249 ( n180 , n1386 );
    and g250 ( n1399 , n930 , n655 );
    or g251 ( n1740 , n824 , n618 );
    or g252 ( n777 , n137 , n207 );
    or g253 ( n1315 , n1328 , n900 );
    nor g254 ( n1513 , n1405 , n823 );
    or g255 ( n199 , n915 , n257 );
    and g256 ( n1267 , n416 , n444 );
    not g257 ( n239 , n50 );
    xnor g258 ( n48 , n613 , n405 );
    nor g259 ( n800 , n318 , n781 );
    or g260 ( n1033 , n514 , n989 );
    or g261 ( n738 , n682 , n668 );
    and g262 ( n536 , n790 , n240 );
    not g263 ( n551 , n1007 );
    xnor g264 ( n93 , n899 , n960 );
    or g265 ( n639 , n1657 , n403 );
    xnor g266 ( n1037 , n469 , n1055 );
    and g267 ( n511 , n637 , n1078 );
    or g268 ( n326 , n1333 , n1150 );
    not g269 ( n1297 , n1077 );
    or g270 ( n1741 , n1141 , n1731 );
    not g271 ( n80 , n938 );
    or g272 ( n1243 , n47 , n1022 );
    or g273 ( n1624 , n838 , n983 );
    not g274 ( n240 , n808 );
    or g275 ( n483 , n238 , n839 );
    or g276 ( n1718 , n5 , n1722 );
    and g277 ( n303 , n691 , n639 );
    not g278 ( n134 , n1261 );
    and g279 ( n1016 , n755 , n721 );
    not g280 ( n1150 , n668 );
    xnor g281 ( n422 , n675 , n1398 );
    nor g282 ( n817 , n736 , n1422 );
    or g283 ( n88 , n20 , n864 );
    or g284 ( n1482 , n170 , n1545 );
    not g285 ( n1599 , n887 );
    or g286 ( n963 , n1461 , n444 );
    and g287 ( n1106 , n119 , n1002 );
    buf g288 ( n230 , n831 );
    nor g289 ( n1526 , n630 , n1355 );
    and g290 ( n1570 , n1673 , n1390 );
    xnor g291 ( n1661 , n99 , n129 );
    xnor g292 ( n242 , n1637 , n606 );
    not g293 ( n1324 , n1396 );
    or g294 ( n1043 , n1724 , n386 );
    buf g295 ( n509 , n769 );
    or g296 ( n1614 , n1298 , n1394 );
    not g297 ( n249 , n1116 );
    or g298 ( n1437 , n1542 , n875 );
    xnor g299 ( n378 , n224 , n211 );
    nor g300 ( n1087 , n721 , n1502 );
    nand g301 ( n1221 , n1438 , n1536 );
    xnor g302 ( n437 , n1220 , n394 );
    or g303 ( n1427 , n1407 , n1562 );
    or g304 ( n235 , n1377 , n1756 );
    xnor g305 ( n570 , n708 , n948 );
    or g306 ( n1375 , n229 , n770 );
    and g307 ( n1455 , n1004 , n1044 );
    xnor g308 ( n90 , n265 , n24 );
    not g309 ( n1486 , n1635 );
    or g310 ( n227 , n150 , n1290 );
    and g311 ( n1094 , n1319 , n205 );
    or g312 ( n1384 , n309 , n444 );
    not g313 ( n749 , n419 );
    xnor g314 ( n1417 , n1303 , n1641 );
    not g315 ( n883 , n1629 );
    xnor g316 ( n1045 , n43 , n33 );
    or g317 ( n387 , n217 , n877 );
    not g318 ( n820 , n203 );
    not g319 ( n1314 , n263 );
    not g320 ( n1144 , n212 );
    or g321 ( n466 , n441 , n636 );
    and g322 ( n950 , n1692 , n483 );
    or g323 ( n655 , n971 , n530 );
    xnor g324 ( n112 , n42 , n907 );
    xnor g325 ( n794 , n225 , n1208 );
    or g326 ( n167 , n238 , n222 );
    or g327 ( n1251 , n1293 , n708 );
    or g328 ( n1019 , n651 , n527 );
    and g329 ( n1396 , n100 , n1666 );
    and g330 ( n660 , n676 , n197 );
    and g331 ( n1078 , n248 , n527 );
    not g332 ( n135 , n1073 );
    xnor g333 ( n1051 , n689 , n168 );
    and g334 ( n496 , n564 , n473 );
    xnor g335 ( n1339 , n66 , n336 );
    or g336 ( n1629 , n2 , n684 );
    buf g337 ( n1177 , n487 );
    xnor g338 ( n1639 , n302 , n801 );
    and g339 ( n465 , n1152 , n491 );
    nand g340 ( n433 , n315 , n997 );
    or g341 ( n677 , n1648 , n1232 );
    or g342 ( n1011 , n1513 , n1426 );
    or g343 ( n740 , n1309 , n1742 );
    not g344 ( n1321 , n691 );
    xnor g345 ( n534 , n248 , n472 );
    or g346 ( n515 , n579 , n706 );
    not g347 ( n386 , n1174 );
    xnor g348 ( n1459 , n321 , n1507 );
    or g349 ( n490 , n1029 , n748 );
    and g350 ( n519 , n1682 , n994 );
    or g351 ( n1060 , n762 , n1702 );
    not g352 ( n850 , n1061 );
    not g353 ( n803 , n413 );
    not g354 ( n14 , n1279 );
    or g355 ( n1151 , n868 , n212 );
    or g356 ( n1501 , n1140 , n148 );
    not g357 ( n429 , n1629 );
    not g358 ( n1700 , n1582 );
    and g359 ( n231 , n565 , n1150 );
    or g360 ( n463 , n836 , n240 );
    or g361 ( n32 , n884 , n745 );
    xnor g362 ( n1527 , n311 , n1706 );
    and g363 ( n768 , n214 , n981 );
    not g364 ( n1219 , n561 );
    or g365 ( n406 , n845 , n1070 );
    or g366 ( n662 , n282 , n496 );
    or g367 ( n943 , n1491 , n1722 );
    and g368 ( n1035 , n732 , n340 );
    or g369 ( n451 , n979 , n647 );
    nor g370 ( n1454 , n1742 , n1035 );
    or g371 ( n1349 , n1630 , n1405 );
    and g372 ( n228 , n268 , n1168 );
    or g373 ( n926 , n1413 , n356 );
    and g374 ( n991 , n1059 , n946 );
    nor g375 ( n928 , n1089 , n787 );
    or g376 ( n1216 , n1057 , n226 );
    and g377 ( n1597 , n1692 , n1509 );
    and g378 ( n1522 , n1103 , n491 );
    buf g379 ( n292 , n408 );
    xnor g380 ( n1462 , n1572 , n769 );
    nor g381 ( n858 , n490 , n1229 );
    or g382 ( n359 , n1216 , n932 );
    or g383 ( n419 , n591 , n530 );
    not g384 ( n221 , n605 );
    and g385 ( n867 , n1555 , n117 );
    xnor g386 ( n442 , n1515 , n1487 );
    or g387 ( n765 , n774 , n982 );
    or g388 ( n533 , n1367 , n149 );
    xnor g389 ( n1142 , n371 , n1665 );
    not g390 ( n784 , n1648 );
    and g391 ( n1020 , n906 , n1371 );
    or g392 ( n1607 , n679 , n389 );
    or g393 ( n41 , n721 , n223 );
    nor g394 ( n1117 , n408 , n704 );
    and g395 ( n1602 , n63 , n1374 );
    and g396 ( n1007 , n1349 , n1077 );
    xnor g397 ( n717 , n1402 , n895 );
    or g398 ( n1086 , n1479 , n738 );
    and g399 ( n1228 , n84 , n777 );
    or g400 ( n289 , n811 , n1432 );
    or g401 ( n1708 , n529 , n1555 );
    not g402 ( n1715 , n1064 );
    or g403 ( n697 , n1493 , n677 );
    xnor g404 ( n121 , n1623 , n739 );
    xnor g405 ( n1694 , n841 , n1470 );
    nor g406 ( n1080 , n994 , n242 );
    or g407 ( n1467 , n1655 , n1119 );
    or g408 ( n69 , n1049 , n368 );
    and g409 ( n1655 , n589 , n835 );
    nor g410 ( n989 , n1399 , n452 );
    xnor g411 ( n1734 , n1232 , n225 );
    nor g412 ( n809 , n1493 , n435 );
    nor g413 ( n588 , n18 , n1726 );
    not g414 ( n1076 , n1250 );
    xnor g415 ( n1169 , n321 , n1336 );
    not g416 ( n1357 , n1432 );
    nor g417 ( n1434 , n1535 , n659 );
    and g418 ( n653 , n1528 , n1703 );
    nor g419 ( n25 , n144 , n306 );
    nor g420 ( n956 , n1364 , n901 );
    or g421 ( n930 , n238 , n1071 );
    and g422 ( n1323 , n40 , n257 );
    or g423 ( n364 , n1477 , n1508 );
    and g424 ( n1407 , n1212 , n1650 );
    xnor g425 ( n1279 , n1530 , n138 );
    nor g426 ( n183 , n741 , n891 );
    or g427 ( n1484 , n467 , n363 );
    xnor g428 ( n1483 , n1159 , n610 );
    and g429 ( n682 , n545 , n758 );
    not g430 ( n564 , n479 );
    not g431 ( n139 , n78 );
    xnor g432 ( n187 , n38 , n1009 );
    and g433 ( n142 , n735 , n887 );
    xnor g434 ( n772 , n859 , n825 );
    nor g435 ( n661 , n803 , n94 );
    or g436 ( n1028 , n921 , n1541 );
    or g437 ( n126 , n1449 , n566 );
    xnor g438 ( n12 , n236 , n1496 );
    or g439 ( n869 , n1127 , n197 );
    xnor g440 ( n1543 , n1659 , n111 );
    or g441 ( n1332 , n1379 , n578 );
    xnor g442 ( n1340 , n874 , n1635 );
    or g443 ( n735 , n524 , n257 );
    or g444 ( n1173 , n1553 , n198 );
    nor g445 ( n443 , n1575 , n402 );
    or g446 ( n913 , n1106 , n1559 );
    xor g447 ( n1727 , n949 , n857 );
    not g448 ( n896 , n1734 );
    not g449 ( n269 , n750 );
    nor g450 ( n253 , n1537 , n1307 );
    and g451 ( n1240 , n689 , n576 );
    or g452 ( n1545 , n169 , n1728 );
    xor g453 ( n1196 , n1021 , n1301 );
    nor g454 ( n659 , n1405 , n1389 );
    not g455 ( n484 , n1202 );
    and g456 ( n250 , n1193 , n491 );
    xnor g457 ( n427 , n470 , n157 );
    and g458 ( n819 , n159 , n835 );
    nor g459 ( n390 , n1026 , n340 );
    not g460 ( n190 , n1627 );
    buf g461 ( n1253 , n1050 );
    xnor g462 ( n369 , n66 , n172 );
    or g463 ( n1293 , n980 , n358 );
    xnor g464 ( n1166 , n1249 , n957 );
    and g465 ( n683 , n1126 , n1204 );
    and g466 ( n333 , n1121 , n491 );
    xnor g467 ( n89 , n249 , n327 );
    and g468 ( n1184 , n1672 , n1634 );
    or g469 ( n448 , n98 , n1383 );
    or g470 ( n505 , n976 , n1705 );
    nor g471 ( n774 , n205 , n1390 );
    xnor g472 ( n542 , n654 , n1380 );
    xnor g473 ( n754 , n752 , n851 );
    not g474 ( n602 , n413 );
    or g475 ( n1590 , n1483 , n1030 );
    not g476 ( n461 , n302 );
    xnor g477 ( n753 , n543 , n1716 );
    and g478 ( n1414 , n446 , n476 );
    or g479 ( n0 , n627 , n1341 );
    or g480 ( n750 , n1210 , n747 );
    xnor g481 ( n1273 , n1604 , n505 );
    or g482 ( n1392 , n1275 , n1046 );
    nor g483 ( n1128 , n896 , n783 );
    or g484 ( n211 , n1080 , n1621 );
    or g485 ( n815 , n1649 , n1088 );
    nor g486 ( n1693 , n1217 , n911 );
    and g487 ( n1571 , n879 , n900 );
    or g488 ( n573 , n1007 , n145 );
    and g489 ( n1717 , n1200 , n1664 );
    not g490 ( n1079 , n538 );
    not g491 ( n906 , n1733 );
    xnor g492 ( n181 , n1468 , n1505 );
    and g493 ( n804 , n262 , n602 );
    not g494 ( n42 , n1743 );
    or g495 ( n512 , n369 , n1271 );
    and g496 ( n20 , n1419 , n237 );
    or g497 ( n1490 , n1518 , n1053 );
    xnor g498 ( n1171 , n1260 , n1725 );
    and g499 ( n1070 , n409 , n1136 );
    xnor g500 ( n557 , n1530 , n841 );
    or g501 ( n698 , n1324 , n61 );
    or g502 ( n377 , n1414 , n583 );
    xnor g503 ( n1507 , n302 , n473 );
    not g504 ( n1622 , n941 );
    nor g505 ( n1460 , n811 , n1079 );
    buf g506 ( n23 , n346 );
    or g507 ( n863 , n835 , n1500 );
    xor g508 ( n957 , n653 , n972 );
    or g509 ( n97 , n1189 , n449 );
    buf g510 ( n1534 , n920 );
    or g511 ( n616 , n687 , n979 );
    xnor g512 ( n418 , n471 , n332 );
    xnor g513 ( n893 , n1700 , n339 );
    or g514 ( n1676 , n1660 , n681 );
    not g515 ( n1568 , n1476 );
    or g516 ( n1050 , n1361 , n1237 );
    or g517 ( n771 , n1144 , n1579 );
    and g518 ( n651 , n287 , n1382 );
    not g519 ( n1352 , n972 );
    xnor g520 ( n129 , n1434 , n488 );
    nor g521 ( n432 , n1135 , n265 );
    and g522 ( n618 , n87 , n602 );
    or g523 ( n709 , n110 , n377 );
    or g524 ( n908 , n1739 , n1116 );
    nor g525 ( n813 , n721 , n775 );
    not g526 ( n578 , n635 );
    or g527 ( n1236 , n531 , n1701 );
    or g528 ( n736 , n1190 , n1493 );
    and g529 ( n49 , n1180 , n163 );
    xnor g530 ( n1359 , n654 , n901 );
    or g531 ( n1270 , n313 , n105 );
    and g532 ( n877 , n1276 , n757 );
    nor g533 ( n1160 , n570 , n1505 );
    and g534 ( n1318 , n668 , n754 );
    xnor g535 ( n363 , n1416 , n142 );
    nor g536 ( n1531 , n573 , n759 );
    and g537 ( n1681 , n1560 , n1025 );
    xnor g538 ( n940 , n579 , n756 );
    not g539 ( n886 , n728 );
    nor g540 ( n1124 , n257 , n1616 );
    buf g541 ( n85 , n153 );
    xnor g542 ( n1207 , n1317 , n1572 );
    nor g543 ( n1542 , n644 , n1484 );
    xnor g544 ( n1475 , n1392 , n1592 );
    and g545 ( n619 , n107 , n1206 );
    nor g546 ( n711 , n1574 , n1650 );
    or g547 ( n1248 , n1321 , n1217 );
    and g548 ( n295 , n1396 , n326 );
    xnor g549 ( n766 , n1019 , n203 );
    or g550 ( n53 , n1591 , n1478 );
    buf g551 ( n173 , n823 );
    xnor g552 ( n384 , n471 , n68 );
    and g553 ( n36 , n1681 , n1539 );
    not g554 ( n263 , n308 );
    xnor g555 ( n907 , n750 , n293 );
    or g556 ( n297 , n345 , n384 );
    not g557 ( n558 , n977 );
    not g558 ( n844 , n1468 );
    or g559 ( n909 , n26 , n238 );
    or g560 ( n873 , n858 , n978 );
    or g561 ( n517 , n398 , n1198 );
    xnor g562 ( n751 , n1021 , n725 );
    buf g563 ( n453 , n1359 );
    not g564 ( n925 , n248 );
    or g565 ( n623 , n258 , n1113 );
    or g566 ( n1487 , n271 , n51 );
    or g567 ( n1029 , n1184 , n1153 );
    nand g568 ( n208 , n478 , n1095 );
    and g569 ( n672 , n468 , n322 );
    xnor g570 ( n767 , n580 , n1043 );
    or g571 ( n1518 , n361 , n1272 );
    or g572 ( n1654 , n19 , n1098 );
    and g573 ( n1529 , n199 , n1451 );
    xnor g574 ( n72 , n929 , n650 );
    or g575 ( n713 , n36 , n387 );
    xnor g576 ( n636 , n133 , n857 );
    nor g577 ( n464 , n868 , n829 );
    xnor g578 ( n19 , n353 , n1291 );
    xnor g579 ( n237 , n722 , n222 );
    not g580 ( n1046 , n1310 );
    not g581 ( n351 , n613 );
    xnor g582 ( n825 , n8 , n1262 );
    and g583 ( n1704 , n902 , n1650 );
    and g584 ( n68 , n909 , n1703 );
    or g585 ( n1595 , n1447 , n819 );
    or g586 ( n1588 , n956 , n1334 );
    not g587 ( n783 , n772 );
    not g588 ( n1453 , n441 );
    nor g589 ( n786 , n7 , n911 );
    or g590 ( n366 , n776 , n608 );
    and g591 ( n878 , n1041 , n899 );
    and g592 ( n1669 , n1713 , n1269 );
    not g593 ( n1294 , n1251 );
    or g594 ( n1062 , n900 , n727 );
    or g595 ( n1178 , n614 , n649 );
    or g596 ( n1258 , n1378 , n1348 );
    or g597 ( n1678 , n988 , n1743 );
    or g598 ( n945 , n508 , n1460 );
    and g599 ( n1304 , n1222 , n314 );
    not g600 ( n797 , n33 );
    and g601 ( n270 , n837 , n519 );
    nor g602 ( n1697 , n911 , n253 );
    or g603 ( n1587 , n1375 , n120 );
    not g604 ( n1112 , n945 );
    and g605 ( n583 , n446 , n646 );
    xnor g606 ( n44 , n1583 , n856 );
    nor g607 ( n1649 , n721 , n399 );
    nor g608 ( n1643 , n636 , n1409 );
    and g609 ( n604 , n977 , n1756 );
    nor g610 ( n995 , n201 , n1395 );
    or g611 ( n8 , n784 , n321 );
    not g612 ( n792 , n1572 );
    or g613 ( n81 , n1120 , n994 );
    or g614 ( n1322 , n1590 , n426 );
    not g615 ( n446 , n28 );
    not g616 ( n205 , n993 );
    buf g617 ( n428 , n1588 );
    nor g618 ( n1755 , n602 , n45 );
    or g619 ( n555 , n1331 , n1601 );
    not g620 ( n74 , n1226 );
    and g621 ( n1466 , n254 , n491 );
    and g622 ( n1561 , n1289 , n197 );
    buf g623 ( n1632 , n1186 );
    and g624 ( n133 , n853 , n959 );
    and g625 ( n1254 , n673 , n1224 );
    or g626 ( n1422 , n461 , n1667 );
    or g627 ( n1611 , n1199 , n325 );
    nor g628 ( n1424 , n603 , n715 );
    not g629 ( n1111 , n489 );
    or g630 ( n854 , n1720 , n39 );
    or g631 ( n657 , n669 , n126 );
    buf g632 ( n1042 , n1566 );
    or g633 ( n360 , n672 , n1395 );
    or g634 ( n493 , n1594 , n1587 );
    xnor g635 ( n540 , n888 , n134 );
    or g636 ( n22 , n1027 , n1549 );
    nand g637 ( n255 , n1054 , n1040 );
    and g638 ( n322 , n568 , n703 );
    and g639 ( n1514 , n598 , n444 );
    xnor g640 ( n216 , n1462 , n1746 );
    not g641 ( n708 , n706 );
    or g642 ( n757 , n462 , n1 );
    xnor g643 ( n902 , n1311 , n991 );
    or g644 ( n725 , n660 , n1599 );
    not g645 ( n1089 , n1388 );
    and g646 ( n1598 , n515 , n495 );
    xnor g647 ( n1082 , n611 , n1109 );
    not g648 ( n935 , n612 );
    buf g649 ( n1729 , n138 );
    and g650 ( n1153 , n140 , n637 );
    or g651 ( n43 , n624 , n250 );
    and g652 ( n576 , n311 , n789 );
    buf g653 ( n726 , n1296 );
    and g654 ( n903 , n1652 , n1708 );
    xnor g655 ( n1410 , n613 , n968 );
    not g656 ( n1505 , n982 );
    xnor g657 ( n92 , n513 , n90 );
    nor g658 ( n1580 , n587 , n1554 );
    xor g659 ( n723 , n1579 , n1026 );
    buf g660 ( n1285 , n1401 );
    nor g661 ( n440 , n846 , n1610 );
    not g662 ( n1102 , n984 );
    nor g663 ( n884 , n602 , n1656 );
    nor g664 ( n1653 , n1135 , n1125 );
    buf g665 ( n585 , n553 );
    not g666 ( n281 , n295 );
    nand g667 ( n319 , n593 , n1286 );
    and g668 ( n445 , n1523 , n900 );
    buf g669 ( n501 , n200 );
    or g670 ( n1257 , n1656 , n1486 );
    or g671 ( n450 , n1047 , n528 );
    xnor g672 ( n1665 , n1694 , n1279 );
    nor g673 ( n1141 , n1196 , n342 );
    nor g674 ( n356 , n49 , n1718 );
    nor g675 ( n528 , n1248 , n320 );
    or g676 ( n186 , n19 , n1199 );
    and g677 ( n834 , n302 , n496 );
    xor g678 ( n818 , n172 , n1456 );
    nor g679 ( n330 , n14 , n1284 );
    nor g680 ( n122 , n1640 , n718 );
    not g681 ( n791 , n998 );
    or g682 ( n28 , n1235 , n486 );
    not g683 ( n1450 , n742 );
    xnor g684 ( n597 , n1179 , n321 );
    buf g685 ( n1337 , n1138 );
    or g686 ( n402 , n1499 , n466 );
    or g687 ( n1031 , n34 , n1168 );
    nor g688 ( n875 , n974 , n1170 );
    or g689 ( n1010 , n303 , n160 );
    or g690 ( n656 , n190 , n1168 );
    not g691 ( n1110 , n323 );
    not g692 ( n495 , n982 );
    xnor g693 ( n1130 , n79 , n535 );
    or g694 ( n1385 , n1596 , n1466 );
    or g695 ( n146 , n632 , n763 );
    nor g696 ( n1198 , n1072 , n42 );
    xnor g697 ( n1261 , n154 , n567 );
    not g698 ( n1104 , n138 );
    or g699 ( n1485 , n1163 , n826 );
    or g700 ( n210 , n926 , n252 );
    xnor g701 ( n888 , n1740 , n374 );
    nor g702 ( n1619 , n28 , n1754 );
    xor g703 ( n898 , n68 , n406 );
    not g704 ( n796 , n243 );
    not g705 ( n1165 , n950 );
    not g706 ( n780 , n880 );
    not g707 ( n24 , n568 );
    or g708 ( n1147 , n1550 , n629 );
    not g709 ( n704 , n1303 );
    or g710 ( n1489 , n1535 , n928 );
    nor g711 ( n1367 , n769 , n792 );
    buf g712 ( n497 , n1656 );
    and g713 ( n1351 , n1694 , n39 );
    and g714 ( n841 , n63 , n382 );
    and g715 ( n1402 , n1680 , n656 );
    xnor g716 ( n1711 , n74 , n1344 );
    and g717 ( n904 , n558 , n960 );
    or g718 ( n584 , n471 , n647 );
    or g719 ( n1579 , n870 , n601 );
    not g720 ( n890 , n671 );
    xnor g721 ( n793 , n1287 , n1661 );
    nor g722 ( n168 , n1228 , n576 );
    or g723 ( n538 , n140 , n1078 );
    not g724 ( n1266 , n1616 );
    not g725 ( n62 , n506 );
    xnor g726 ( n795 , n385 , n92 );
    nor g727 ( n688 , n545 , n264 );
    and g728 ( n531 , n562 , n1356 );
    xnor g729 ( n277 , n1577 , n815 );
    xnor g730 ( n629 , n949 , n375 );
    not g731 ( n1328 , n1114 );
    not g732 ( n1115 , n392 );
    not g733 ( n1341 , n487 );
    and g734 ( n1720 , n1104 , n1530 );
    and g735 ( n304 , n420 , n832 );
    not g736 ( n543 , n1529 );
    not g737 ( n1131 , n1717 );
    not g738 ( n1309 , n500 );
    xnor g739 ( n164 , n1672 , n482 );
    and g740 ( n739 , n37 , n1511 );
    or g741 ( n1161 , n1136 , n980 );
    and g742 ( n876 , n1093 , n1384 );
    and g743 ( n527 , n1228 , n689 );
    xnor g744 ( n264 , n1714 , n954 );
    not g745 ( n1074 , n1283 );
    or g746 ( n901 , n639 , n1693 );
    xor g747 ( n513 , n237 , n468 );
    or g748 ( n548 , n847 , n1222 );
    nor g749 ( n983 , n335 , n1663 );
    nor g750 ( n523 , n276 , n1134 );
    nor g751 ( n762 , n183 , n1678 );
    xnor g752 ( n467 , n1083 , n1492 );
    and g753 ( n1635 , n1692 , n1372 );
    or g754 ( n565 , n1422 , n746 );
    and g755 ( n1343 , n658 , n869 );
    xnor g756 ( n1090 , n1291 , n1165 );
    not g757 ( n191 , n604 );
    not g758 ( n703 , n237 );
    and g759 ( n149 , n586 , n1462 );
    or g760 ( n569 , n193 , n1222 );
    xnor g761 ( n613 , n543 , n1401 );
    not g762 ( n401 , n589 );
    xnor g763 ( n675 , n1546 , n1091 );
    not g764 ( n413 , n308 );
    and g765 ( n978 , n490 , n158 );
    or g766 ( n1097 , n1377 , n1201 );
    not g767 ( n345 , n101 );
    and g768 ( n415 , n958 , n490 );
    or g769 ( n1680 , n1089 , n153 );
    xnor g770 ( n1737 , n785 , n1392 );
    xnor g771 ( n1030 , n285 , n215 );
    and g772 ( n1731 , n899 , n499 );
    or g773 ( n1260 , n1605 , n618 );
    or g774 ( n918 , n657 , n828 );
    or g775 ( n700 , n1223 , n279 );
    xnor g776 ( n1159 , n1404 , n1233 );
    nor g777 ( n127 , n1733 , n1000 );
    xnor g778 ( n518 , n1742 , n893 );
    not g779 ( n939 , n1018 );
    not g780 ( n2 , n986 );
    xnor g781 ( n837 , n1317 , n626 );
    not g782 ( n673 , n698 );
    not g783 ( n1388 , n1314 );
    not g784 ( n911 , n994 );
    xnor g785 ( n625 , n1236 , n1465 );
    and g786 ( n1176 , n1260 , n1725 );
    and g787 ( n870 , n1631 , n580 );
    xnor g788 ( n16 , n322 , n1270 );
    or g789 ( n508 , n296 , n1634 );
    nor g790 ( n720 , n996 , n1284 );
    not g791 ( n836 , n1156 );
    or g792 ( n605 , n291 , n530 );
    xnor g793 ( n1671 , n1385 , n722 );
    nor g794 ( n761 , n257 , n408 );
    not g795 ( n521 , n1451 );
    or g796 ( n1329 , n979 , n647 );
    nor g797 ( n816 , n688 , n1580 );
    nor g798 ( n354 , n374 , n1646 );
    or g799 ( n1638 , n627 , n559 );
    or g800 ( n1705 , n533 , n9 );
    or g801 ( n196 , n835 , n1566 );
    or g802 ( n724 , n425 , n333 );
    not g803 ( n1503 , n347 );
    and g804 ( n1426 , n882 , n1405 );
    nor g805 ( n472 , n1019 , n1240 );
    xnor g806 ( n1232 , n653 , n695 );
    or g807 ( n325 , n1118 , n404 );
    or g808 ( n381 , n267 , n705 );
    not g809 ( n1510 , n321 );
    and g810 ( n1577 , n1161 , n1538 );
    xnor g811 ( n1391 , n14 , n833 );
    nor g812 ( n696 , n899 , n1264 );
    nor g813 ( n398 , n1085 , n830 );
    not g814 ( n1650 , n738 );
    or g815 ( n1100 , n1039 , n135 );
    not g816 ( n404 , n1593 );
    or g817 ( n1262 , n1677 , n939 );
    and g818 ( n666 , n607 , n1004 );
    not g819 ( n1723 , n502 );
    buf g820 ( n782 , n222 );
    not g821 ( n630 , n1295 );
    or g822 ( n347 , n1614 , n295 );
    or g823 ( n830 , n696 , n1743 );
    not g824 ( n1003 , n227 );
    and g825 ( n1724 , n1576 , n1458 );
    or g826 ( n462 , n594 , n1741 );
    or g827 ( n1284 , n98 , n1064 );
    nor g828 ( n294 , n1263 , n780 );
    xnor g829 ( n648 , n311 , n820 );
    or g830 ( n938 , n1584 , n1264 );
    not g831 ( n336 , n631 );
    or g832 ( n57 , n116 , n1405 );
    or g833 ( n1200 , n666 , n207 );
    and g834 ( n1362 , n1020 , n583 );
    buf g835 ( n1421 , n695 );
    not g836 ( n892 , n507 );
    or g837 ( n1049 , n1535 , n661 );
    not g838 ( n1564 , n1385 );
    or g839 ( n612 , n1369 , n530 );
    nor g840 ( n1 , n1245 , n1444 );
    or g841 ( n759 , n1722 , n614 );
    buf g842 ( n27 , n947 );
    not g843 ( n1001 , n622 );
    xnor g844 ( n1116 , n278 , n346 );
    or g845 ( n83 , n1259 , n521 );
    nor g846 ( n1423 , n1145 , n1318 );
    and g847 ( n840 , n736 , n697 );
    or g848 ( n912 , n187 , n1130 );
    or g849 ( n1211 , n1241 , n897 );
    not g850 ( n342 , n904 );
    nor g851 ( n61 , n1333 , n1395 );
    not g852 ( n1535 , n1747 );
    xnor g853 ( n1651 , n1123 , n940 );
    nor g854 ( n1185 , n721 , n1301 );
    not g855 ( n238 , n413 );
    nor g856 ( n715 , n680 , n622 );
    not g857 ( n1127 , n600 );
    xnor g858 ( n339 , n1303 , n408 );
    not g859 ( n1601 , n266 );
    or g860 ( n37 , n293 , n269 );
    or g861 ( n827 , n127 , n1158 );
    or g862 ( n1575 , n629 , n1620 );
    and g863 ( n1280 , n1020 , n1414 );
    and g864 ( n1431 , n248 , n1240 );
    nor g865 ( n355 , n721 , n374 );
    or g866 ( n343 , n1453 , n1499 );
    xnor g867 ( n1620 , n1494 , n664 );
    and g868 ( n5 , n57 , n605 );
    nor g869 ( n634 , n1581 , n1606 );
    or g870 ( n31 , n721 , n1592 );
    or g871 ( n714 , n1036 , n995 );
    xor g872 ( n1055 , n1412 , n74 );
    and g873 ( n296 , n1342 , n1392 );
    or g874 ( n7 , n14 , n448 );
    not g875 ( n108 , n722 );
    xnor g876 ( n891 , n1642 , n920 );
    nor g877 ( n226 , n1149 , n868 );
    and g878 ( n1412 , n1732 , n635 );
    not g879 ( n1390 , n756 );
    buf g880 ( n352 , n1463 );
    not g881 ( n1630 , n77 );
    nor g882 ( n1192 , n547 , n942 );
    buf g883 ( n417 , n399 );
    or g884 ( n1732 , n890 , n257 );
    not g885 ( n1242 , n601 );
    and g886 ( n1319 , n125 , n1602 );
    nor g887 ( n942 , n1181 , n599 );
    or g888 ( n494 , n1607 , n122 );
    nor g889 ( n328 , n900 , n831 );
    and g890 ( n603 , n680 , n274 );
    not g891 ( n915 , n82 );
    or g892 ( n1032 , n1376 , n238 );
    or g893 ( n965 , n1755 , n1709 );
    xnor g894 ( n321 , n266 , n612 );
    buf g895 ( n130 , n1592 );
    or g896 ( n553 , n450 , n1010 );
    xnor g897 ( n1498 , n311 , n945 );
    or g898 ( n1068 , n1722 , n614 );
    not g899 ( n1296 , n992 );
    and g900 ( n1615 , n545 , n283 );
    or g901 ( n1583 , n1129 , n843 );
    not g902 ( n1667 , n473 );
    or g903 ( n1581 , n494 , n91 );
    not g904 ( n1252 , n1569 );
    xnor g905 ( n1540 , n98 , n837 );
    nor g906 ( n562 , n698 , n1108 );
    nor g907 ( n55 , n628 , n1469 );
    or g908 ( n1186 , n1047 , n872 );
    and g909 ( n716 , n231 , n795 );
    and g910 ( n1101 , n969 , n1206 );
    or g911 ( n457 , n827 , n1452 );
    xnor g912 ( n1063 , n613 , n136 );
    or g913 ( n1356 , n1444 , n1001 );
    and g914 ( n1331 , n1222 , n1411 );
    or g915 ( n1238 , n1171 , n1457 );
    or g916 ( n405 , n1353 , n290 );
    and g917 ( n756 , n141 , n1688 );
    or g918 ( n1069 , n257 , n220 );
    and g919 ( n1683 , n1669 , n682 );
    or g920 ( n1093 , n257 , n293 );
    not g921 ( n1004 , n1314 );
    or g922 ( n642 , n1450 , n530 );
    or g923 ( n217 , n550 , n415 );
    or g924 ( n160 , n485 , n563 );
    not g925 ( n1136 , n413 );
    xnor g926 ( n1373 , n753 , n767 );
    or g927 ( n403 , n1351 , n720 );
    xnor g928 ( n763 , n179 , n1595 );
    or g929 ( n1077 , n298 , n1458 );
    or g930 ( n730 , n1455 , n1348 );
    xnor g931 ( n1065 , n592 , n305 );
    xnor g932 ( n1419 , n1385 , n1463 );
    not g933 ( n678 , n1595 );
    not g934 ( n491 , n413 );
    not g935 ( n1000 , n1581 );
    xnor g936 ( n954 , n896 , n1169 );
    or g937 ( n833 , n1705 , n480 );
    not g938 ( n198 , n569 );
    not g939 ( n776 , n1388 );
    or g940 ( n1657 , n414 , n329 );
    not g941 ( n162 , n1428 );
    or g942 ( n1471 , n316 , n191 );
    or g943 ( n951 , n19 , n1098 );
    not g944 ( n475 , n1149 );
    or g945 ( n1554 , n1179 , n1128 );
    not g946 ( n193 , n54 );
    nor g947 ( n1330 , n1165 , n970 );
    or g948 ( n110 , n1567 , n683 );
    and g949 ( n948 , n1293 , n844 );
    nor g950 ( n1744 , n55 , n911 );
    buf g951 ( n1547 , n420 );
    nor g952 ( n897 , n1733 , n634 );
    not g953 ( n1405 , n728 );
    nor g954 ( n1726 , n1206 , n1205 );
    nor g955 ( n712 , n1041 , n904 );
    not g956 ( n1491 , n964 );
    xor g957 ( n1377 , n725 , n1566 );
    buf g958 ( n498 , n293 );
    xnor g959 ( n1672 , n785 , n318 );
    or g960 ( n1433 , n95 , n332 );
    and g961 ( n1157 , n712 , n235 );
    nor g962 ( n1591 , n1512 , n69 );
    and g963 ( n1605 , n1753 , n1222 );
    or g964 ( n194 , n867 , n1522 );
    not g965 ( n1552 , n510 );
    or g966 ( n224 , n699 , n1744 );
    and g967 ( n407 , n1358 , n178 );
    or g968 ( n1473 , n182 , n328 );
    xnor g969 ( n649 , n551 , n1011 );
    or g970 ( n1139 , n101 , n384 );
    nor g971 ( n141 , n1319 , n259 );
    xnor g972 ( n421 , n652 , n1467 );
    and g973 ( n826 , n282 , n302 );
    or g974 ( n1464 , n784 , n1544 );
    nor g975 ( n1574 , n134 , n88 );
    xnor g976 ( n1610 , n431 , n411 );
    not g977 ( n591 , n1647 );
    xnor g978 ( n1546 , n1416 , n115 );
    not g979 ( n1551 , n869 );
    not g980 ( n1013 , n71 );
    xor g981 ( n456 , n1705 , n572 );
    nor g982 ( n1038 , n283 , n1336 );
    or g983 ( n1181 , n1179 , n716 );
    xnor g984 ( n1682 , n1635 , n1656 );
    not g985 ( n1066 , n1059 );
    nand g986 ( n566 , n1520 , n1613 );
    or g987 ( n1012 , n973 , n17 );
    and g988 ( n1557 , n367 , n1229 );
    and g989 ( n919 , n1658 , n711 );
    or g990 ( n852 , n1654 , n1611 );
    not g991 ( n1436 , n1490 );
    or g992 ( n974 , n876 , n1045 );
    or g993 ( n972 , n1397 , n1070 );
    or g994 ( n722 , n151 , n484 );
    not g995 ( n1369 , n1205 );
    or g996 ( n131 , n1117 , n106 );
    or g997 ( n934 , n1540 , n348 );
    or g998 ( n1451 , n850 , n1555 );
    buf g999 ( n275 , n1296 );
    xnor g1000 ( n917 , n846 , n48 );
    or g1001 ( n1118 , n232 , n67 );
    not g1002 ( n444 , n808 );
    or g1003 ( n1203 , n368 , n1014 );
    or g1004 ( n479 , n45 , n1352 );
    xnor g1005 ( n60 , n1682 , n941 );
    not g1006 ( n218 , n1682 );
    and g1007 ( n459 , n300 , n835 );
    not g1008 ( n1206 , n413 );
    not g1009 ( n1298 , n1276 );
    nor g1010 ( n1005 , n467 , n363 );
    not g1011 ( n1544 , n571 );
    nor g1012 ( n1666 , n338 , n1653 );
    xnor g1013 ( n439 , n814 , n256 );
    xnor g1014 ( n215 , n1439 , n1525 );
    or g1015 ( n1008 , n104 , n15 );
    or g1016 ( n1652 , n239 , n1405 );
    or g1017 ( n1452 , n1280 , n1362 );
    xnor g1018 ( n225 , n972 , n45 );
    xnor g1019 ( n449 , n1638 , n986 );
    or g1020 ( n1195 , n1704 , n919 );
    or g1021 ( n764 , n1674 , n1143 );
    xnor g1022 ( n368 , n1295 , n188 );
    not g1023 ( n499 , n235 );
    or g1024 ( n526 , n294 , n1094 );
    xnor g1025 ( n1685 , n876 , n903 );
    and g1026 ( n1413 , n1676 , n1618 );
    or g1027 ( n982 , n490 , n937 );
    or g1028 ( n1690 , n975 , n139 );
    not g1029 ( n532 , n1573 );
    not g1030 ( n1686 , n1039 );
    or g1031 ( n1492 , n1185 , n1480 );
    nor g1032 ( n334 , n405 , n855 );
    xnor g1033 ( n6 , n1489 , n806 );
    and g1034 ( n106 , n204 , n339 );
    xnor g1035 ( n931 , n1123 , n383 );
    or g1036 ( n105 , n913 , n554 );
    buf g1037 ( n773 , n980 );
    or g1038 ( n1174 , n1074 , n1555 );
    nor g1039 ( n628 , n1608 , n1282 );
    nor g1040 ( n1702 , n121 , n42 );
    nor g1041 ( n814 , n1228 , n311 );
    and g1042 ( n1241 , n986 , n737 );
    or g1043 ( n1567 , n1578 , n286 );
    not g1044 ( n397 , n664 );
    and g1045 ( n679 , n949 , n375 );
    xnor g1046 ( n111 , n438 , n410 );
    and g1047 ( n353 , n31 , n1031 );
    or g1048 ( n1308 , n1111 , n1555 );
    or g1049 ( n1312 , n1723 , n444 );
    xnor g1050 ( n1679 , n962 , n860 );
    or g1051 ( n317 , n834 , n817 );
    xnor g1052 ( n247 , n1700 , n1325 );
    buf g1053 ( n640 , n1345 );
    not g1054 ( n1376 , n953 );
    nor g1055 ( n855 , n1358 , n673 );
    nor g1056 ( n1027 , n1570 , n765 );
    nor g1057 ( n1223 , n993 , n908 );
    or g1058 ( n349 , n1624 , n861 );
    not g1059 ( n309 , n1448 );
    nor g1060 ( n985 , n1147 , n1096 );
    or g1061 ( n868 , n1214 , n1700 );
    not g1062 ( n1026 , n267 );
    or g1063 ( n617 , n685 , n336 );
    xnor g1064 ( n535 , n174 , n674 );
    or g1065 ( n853 , n1206 , n138 );
    not g1066 ( n971 , n341 );
    not g1067 ( n1631 , n823 );
    and g1068 ( n1208 , n78 , n435 );
    xnor g1069 ( n370 , n339 , n334 );
    xnor g1070 ( n59 , n546 , n12 );
    xnor g1071 ( n851 , n513 , n16 );
    or g1072 ( n541 , n162 , n238 );
    nor g1073 ( n889 , n257 , n1345 );
    xnor g1074 ( n203 , n811 , n1672 );
    xnor g1075 ( n158 , n44 , n931 );
    or g1076 ( n748 , n1684 , n511 );
    not g1077 ( n95 , n406 );
    nor g1078 ( n395 , n1171 , n1457 );
    xnor g1079 ( n201 , n888 , n1270 );
    nor g1080 ( n937 , n1360 , n1230 );
    and g1081 ( n18 , n729 , n900 );
    not g1082 ( n575 , n490 );
    buf g1083 ( n842 , n1205 );
    nor g1084 ( n1628 , n257 , n246 );
    or g1085 ( n144 , n1751 , n6 );
    or g1086 ( n998 , n197 , n18 );
    or g1087 ( n994 , n1503 , n713 );
    not g1088 ( n529 , n641 );
    not g1089 ( n1721 , n539 );
    nor g1090 ( n1562 , n1748 , n360 );
    not g1091 ( n741 , n37 );
    nor g1092 ( n1549 , n525 , n495 );
    nor g1093 ( n3 , n1206 , n487 );
    not g1094 ( n684 , n1092 );
    xnor g1095 ( n234 , n93 , n1471 );
    or g1096 ( n789 , n757 , n944 );
    not g1097 ( n1429 , n1583 );
    and g1098 ( n685 , n692 , n1188 );
    or g1099 ( n371 , n586 , n1715 );
    or g1100 ( n996 , n731 , n14 );
    and g1101 ( n280 , n1418 , n257 );
    not g1102 ( n241 , n1610 );
    xnor g1103 ( n881 , n166 , n520 );
    xnor g1104 ( n1006 , n237 , n1395 );
    nor g1105 ( n361 , n702 , n147 );
    and g1106 ( n1081 , n865 , n621 );
    xnor g1107 ( n615 , n165 , n1028 );
    nor g1108 ( n65 , n368 , n1014 );
    not g1109 ( n988 , n1756 );
    xnor g1110 ( n622 , n1441 , n234 );
    xnor g1111 ( n860 , n1256 , n766 );
    xnor g1112 ( n1024 , n812 , n1662 );
    or g1113 ( n594 , n1603 , n878 );
    and g1114 ( n632 , n167 , n1730 );
    and g1115 ( n848 , n1516 , n1222 );
    or g1116 ( n1096 , n924 , n35 );
    xnor g1117 ( n455 , n648 , n881 );
    and g1118 ( n1508 , n1735 , n1710 );
    or g1119 ( n101 , n266 , n791 );
    xnor g1120 ( n922 , n843 , n856 );
    and g1121 ( n283 , n473 , n1677 );
    xnor g1122 ( n236 , n1489 , n1751 );
    or g1123 ( n737 , n1638 , n1110 );
    and g1124 ( n1379 , n310 , n240 );
    and g1125 ( n172 , n541 , n419 );
    xnor g1126 ( n1699 , n1173 , n1332 );
    or g1127 ( n707 , n400 , n1522 );
    and g1128 ( n880 , n63 , n1069 );
    nor g1129 ( n1728 , n451 , n96 );
    or g1130 ( n1288 , n912 , n128 );
    or g1131 ( n1047 , n1218 , n429 );
    or g1132 ( n1703 , n1076 , n1004 );
    not g1133 ( n788 , n1282 );
    and g1134 ( n520 , n289 , n1112 );
    and g1135 ( n1137 , n1106 , n888 );
    not g1136 ( n976 , n448 );
    xnor g1137 ( n1039 , n689 , n925 );
    xnor g1138 ( n1233 , n924 , n1494 );
    and g1139 ( n214 , n690 , n1711 );
    and g1140 ( n1122 , n542 , n639 );
    and g1141 ( n1593 , n65 , n365 );
    and g1142 ( n643 , n637 , n1357 );
    nor g1143 ( n1408 , n83 , n1008 );
    nor g1144 ( n1363 , n1045 , n1685 );
    or g1145 ( n1752 , n118 , n208 );
    not g1146 ( n358 , n1597 );
    or g1147 ( n1742 , n1472 , n1633 );
    and g1148 ( n1371 , n590 , n1643 );
    or g1149 ( n932 , n131 , n464 );
    and g1150 ( n480 , n1462 , n270 );
    and g1151 ( n680 , n1151 , n1444 );
    not g1152 ( n424 , n1071 );
    nor g1153 ( n176 , n1683 , n281 );
    or g1154 ( n114 , n1533 , n1431 );
    or g1155 ( n1053 , n1176 , n1274 );
    and g1156 ( n1559 , n1066 , n1311 );
    xor g1157 ( n1589 , n154 , n1740 );
    or g1158 ( n1528 , n1252 , n1136 );
    or g1159 ( n702 , n1197 , n678 );
    and g1160 ( n15 , n1227 , n602 );
    nor g1161 ( n169 , n1433 , n616 );
    xor g1162 ( n1707 , n895 , n551 );
    not g1163 ( n862 , n36 );
    not g1164 ( n84 , n1345 );
    xnor g1165 ( n1249 , n871 , n1258 );
    not g1166 ( n150 , n689 );
    not g1167 ( n705 , n732 );
    nor g1168 ( n1603 , n1301 , n1675 );
    xnor g1169 ( n1670 , n93 , n604 );
    or g1170 ( n1245 , n1196 , n1097 );
    xnor g1171 ( n610 , n1600 , n421 );
    and g1172 ( n1378 , n240 , n1281 );
    or g1173 ( n857 , n1535 , n492 );
    buf g1174 ( n1368 , n420 );
    or g1175 ( n1021 , n733 , n804 );
    nor g1176 ( n434 , n1151 , n673 );
    xnor g1177 ( n1445 , n78 , n1507 );
    nor g1178 ( n1469 , n542 , n788 );
    not g1179 ( n454 , n1217 );
    or g1180 ( n692 , n1749 , n835 );
    and g1181 ( n824 , n645 , n1555 );
    and g1182 ( n400 , n240 , n1023 );
    or g1183 ( n1641 , n848 , n221 );
    or g1184 ( n571 , n1179 , n1510 );
    and g1185 ( n964 , n83 , n1008 );
    xnor g1186 ( n1398 , n504 , n1265 );
    or g1187 ( n941 , n330 , n854 );
    and g1188 ( n1572 , n63 , n393 );
    xnor g1189 ( n952 , n539 , n1454 );
    not g1190 ( n1584 , n1097 );
    or g1191 ( n1684 , n800 , n1425 );
    not g1192 ( n627 , n156 );
    and g1193 ( n1606 , n1371 , n709 );
    nor g1194 ( n1754 , n768 , n1490 );
    not g1195 ( n1333 , n1669 );
    not g1196 ( n1696 , n288 );
    not g1197 ( n291 , n710 );
    and g1198 ( n39 , n1279 , n533 );
    xnor g1199 ( n706 , n923 , n399 );
    xnor g1200 ( n1277 , n1038 , n1690 );
    not g1201 ( n968 , n893 );
    xnor g1202 ( n157 , n1519 , n1300 );
    or g1203 ( n1550 , n1535 , n1087 );
    xnor g1204 ( n411 , n1410 , n373 );
    or g1205 ( n147 , n1171 , n1457 );
    or g1206 ( n621 , n210 , n102 );
    not g1207 ( n1633 , n381 );
    or g1208 ( n1725 , n355 , n1016 );
    nand g1209 ( n118 , n581 , n743 );
    not g1210 ( n1677 , n746 );
    xnor g1211 ( n1220 , n331 , n556 );
    or g1212 ( n1271 , n1131 , n1098 );
    and g1213 ( n1478 , n1593 , n349 );
    not g1214 ( n1264 , n1157 );
    nor g1215 ( n1213 , n249 , n1583 );
    nor g1216 ( n547 , n545 , n1423 );
    or g1217 ( n669 , n1221 , n433 );
    xnor g1218 ( n1014 , n1512 , n1049 );
    not g1219 ( n1311 , n1261 );
    or g1220 ( n375 , n1146 , n459 );
    and g1221 ( n1553 , n1609 , n1555 );
    nor g1222 ( n966 , n721 , n1263 );
    and g1223 ( n577 , n870 , n1582 );
    and g1224 ( n1634 , n987 , n1475 );
    or g1225 ( n1640 , n397 , n260 );
    or g1226 ( n620 , n153 , n1381 );
    not g1227 ( n320 , n387 );
    or g1228 ( n76 , n1136 , n626 );
    buf g1229 ( n1733 , n97 );
    or g1230 ( n1134 , n1712 , n1743 );
    or g1231 ( n163 , n180 , n1168 );
    not g1232 ( n1342 , n1592 );
    or g1233 ( n500 , n705 , n351 );
    xnor g1234 ( n596 , n667 , n751 );
    buf g1235 ( n595 , n1301 );
    or g1236 ( n1303 , n1719 , n681 );
    not g1237 ( n1143 , n124 );
    not g1238 ( n665 , n829 );
    buf g1239 ( n1209 , n1071 );
    xnor g1240 ( n394 , n458 , n213 );
    or g1241 ( n887 , n1625 , n1458 );
    and g1242 ( n1057 , n339 , n577 );
    not g1243 ( n125 , n346 );
    and g1244 ( n66 , n1440 , n463 );
    or g1245 ( n1509 , n835 , n1278 );
    xnor g1246 ( n654 , n1092 , n986 );
    buf g1247 ( n638 , n420 );
    not g1248 ( n278 , n1602 );
    xnor g1249 ( n539 , n580 , n823 );
    not g1250 ( n552 , n1739 );
    xnor g1251 ( n674 , n1602 , n880 );
    or g1252 ( n843 , n552 , n1294 );
    xnor g1253 ( n438 , n1399 , n1344 );
    and g1254 ( n745 , n663 , n1136 );
    xnor g1255 ( n799 , n436 , n1488 );
    xor g1256 ( n1123 , n708 , n1468 );
    not g1257 ( n1125 , n554 );
    or g1258 ( n644 , n1052 , n797 );
    not g1259 ( n145 , n1011 );
    xnor g1260 ( n1439 , n353 , n970 );
    not g1261 ( n1691 , n1173 );
    nor g1262 ( n599 , n231 , n754 );
    xor g1263 ( n650 , n1343 , n1260 );
    buf g1264 ( n1292 , n1616 );
    or g1265 ( n544 , n673 , n440 );
    not g1266 ( n116 , n1586 );
    or g1267 ( n550 , n526 , n700 );
    xnor g1268 ( n1224 , n917 , n1556 );
    not g1269 ( n1230 , n789 );
    xnor g1270 ( n1073 , n439 , n455 );
    and g1271 ( n1530 , n1692 , n863 );
    xnor g1272 ( n894 , n811 , n114 );
    xnor g1273 ( n1745 , n1617 , n596 );
    or g1274 ( n1374 , n900 , n391 );
    or g1275 ( n977 , n920 , n1504 );
    not g1276 ( n1668 , n1175 );
    or g1277 ( n452 , n1412 , n687 );
    and g1278 ( n1425 , n296 , n1672 );
    not g1279 ( n1268 , n1443 );
    nor g1280 ( n838 , n617 , n1313 );
    or g1281 ( n335 , n66 , n1199 );
    buf g1282 ( n1548 , n567 );
    or g1283 ( n441 , n1535 , n209 );
    not g1284 ( n847 , n936 );
    nor g1285 ( n51 , n721 , n947 );
    and g1286 ( n206 , n1155 , n548 );
    or g1287 ( n189 , n368 , n1014 );
    or g1288 ( n435 , n571 , n1232 );
    nor g1289 ( n232 , n1200 , n1664 );
    buf g1290 ( n161 , n457 );
    or g1291 ( n568 , n222 , n108 );
    xnor g1292 ( n1265 , n1067 , n442 );
    and g1293 ( n425 , n1222 , n560 );
    xnor g1294 ( n1499 , n924 , n1550 );
    xnor g1295 ( n469 , n1056 , n898 );
    and g1296 ( n1291 , n1032 , n1310 );
    nor g1297 ( n412 , n941 , n786 );
    and g1298 ( n276 , n960 , n191 );
    not g1299 ( n1025 , n1151 );
    or g1300 ( n113 , n892 , n1458 );
    xnor g1301 ( n856 , n205 , n249 );
    not g1302 ( n808 , n263 );
    xor g1303 ( n1256 , n1228 , n1533 );
    nor g1304 ( n1701 , n136 , n1424 );
    not g1305 ( n1646 , n1740 );
    xnor g1306 ( n689 , n1382 , n1446 );
    not g1307 ( n46 , n1566 );
    xnor g1308 ( n152 , n960 , n1471 );
    or g1309 ( n1558 , n803 , n695 );
    nor g1310 ( n372 , n353 , n537 );
    or g1311 ( n1730 , n796 , n1168 );
    and g1312 ( n1259 , n344 , n197 );
    xnor g1313 ( n546 , n1366 , n1090 );
    xnor g1314 ( n1441 , n812 , n13 );
    nor g1315 ( n1713 , n1135 , n1261 );
    or g1316 ( n128 , n1745 , n1082 );
    or g1317 ( n1674 , n1215 , n297 );
    and g1318 ( n423 , n539 , n1035 );
    or g1319 ( n694 , n467 , n363 );
    or g1320 ( n1533 , n987 , n538 );
    or g1321 ( n1751 , n1535 , n350 );
    nor g1322 ( n1746 , n371 , n270 );
    or g1323 ( n179 , n1267 , n1466 );
    nor g1324 ( n927 , n257 , n920 );
    and g1325 ( n1041 , n46 , n725 );
    nor g1326 ( n652 , n1370 , n3 );
    not g1327 ( n899 , n1196 );
    or g1328 ( n580 , n536 , n1297 );
    nor g1329 ( n389 , n133 , n1495 );
    or g1330 ( n1059 , n1463 , n1564 );
    xnor g1331 ( n1659 , n1517 , n1316 );
    not g1332 ( n115 , n1492 );
    and g1333 ( n949 , n63 , n41 );
    xor g1334 ( n458 , n903 , n43 );
    xnor g1335 ( n274 , n1670 , n1024 );
    and g1336 ( n987 , n1266 , n623 );
    xnor g1337 ( n967 , n1577 , n1751 );
    nor g1338 ( n1145 , n668 , n795 );
    and g1339 ( n258 , n58 , n240 );
    and g1340 ( n1354 , n1020 , n110 );
    and g1341 ( n313 , n134 , n20 );
    or g1342 ( n601 , n475 , n665 );
    and g1343 ( n845 , n29 , n1004 );
    nand g1344 ( n1449 , n284 , n574 );
    or g1345 ( n1519 , n1403 , n371 );
    nor g1346 ( n1442 , n1535 , n1612 );
    or g1347 ( n1494 , n245 , n1571 );
    not g1348 ( n1749 , n52 );
    xnor g1349 ( n1199 , n1456 , n631 );
    and g1350 ( n279 , n205 , n1183 );
    not g1351 ( n1406 , n1618 );
    and g1352 ( n207 , n1246 , n491 );
    xnor g1353 ( n1366 , n1689 , n818 );
    and g1354 ( n924 , n76 , n963 );
    nor g1355 ( n482 , n945 , n1326 );
    not g1356 ( n1400 , n946 );
    xnor g1357 ( n13 , n739 , n80 );
    not g1358 ( n10 , n88 );
    nor g1359 ( n1036 , n432 , n1086 );
    nor g1360 ( n1108 , n359 , n274 );
    or g1361 ( n1204 , n1437 , n1243 );
    or g1362 ( n188 , n966 , n1323 );
    or g1363 ( n1594 , n255 , n319 );
    nor g1364 ( n73 , n152 , n42 );
    nor g1365 ( n1146 , n1405 , n1470 );
    or g1366 ( n1180 , n1405 , n1476 );
    nor g1367 ( n1710 , n1213 , n495 );
    xnor g1368 ( n1098 , n950 , n633 );
    and g1369 ( n1120 , n1608 , n744 );
    or g1370 ( n1663 , n172 , n951 );
    nor g1371 ( n202 , n1026 , n613 );
    not g1372 ( n1688 , n1183 );
    not g1373 ( n209 , n32 );
    and g1374 ( n171 , n1458 , n961 );
    not g1375 ( n136 , n698 );
    not g1376 ( n975 , n503 );
    or g1377 ( n396 , n195 , n1160 );
    not g1378 ( n34 , n1305 );
    not g1379 ( n1472 , n620 );
    nor g1380 ( n1244 , n186 , n512 );
    not g1381 ( n1625 , n1154 );
    not g1382 ( n257 , n728 );
    and g1383 ( n1348 , n299 , n491 );
    not g1384 ( n781 , n785 );
    nor g1385 ( n944 , n1394 , n176 );
    or g1386 ( n4 , n1136 , n1299 );
    xnor g1387 ( n1722 , n1676 , n1618 );
    nor g1388 ( n1034 , n763 , n185 );
    or g1389 ( n1313 , n19 , n1098 );
    not g1390 ( n1560 , n1245 );
    not g1391 ( n1675 , n1021 );
    xnor g1392 ( n431 , n202 , n771 );
    or g1393 ( n1310 , n1365 , n1458 );
    or g1394 ( n871 , n171 , n1601 );
    or g1395 ( n633 , n447 , n445 );
    nor g1396 ( n338 , n1135 , n388 );
    not g1397 ( n1222 , n886 );
    xnor g1398 ( n285 , n123 , n277 );
    and g1399 ( n1129 , n706 , n1468 );
    or g1400 ( n1255 , n62 , n1206 );
    not g1401 ( n910 , n841 );
    not g1402 ( n260 , n1494 );
    and g1403 ( n1275 , n1474 , n1168 );
    and g1404 ( n1512 , n1497 , n1308 );
    xnor g1405 ( n1364 , n1573 , n1629 );
    and g1406 ( n1088 , n1164 , n257 );
    xnor g1407 ( n859 , n1459 , n1277 );
    not g1408 ( n332 , n965 );
    and g1409 ( n1416 , n196 , n113 );
    not g1410 ( n572 , n1257 );
    xnor g1411 ( n647 , n406 , n965 );
    xnor g1412 ( n916 , n1682 , n911 );
    and g1413 ( n1660 , n734 , n240 );
    not g1414 ( n1563 , n200 );
    not g1415 ( n524 , n273 );
    xor g1416 ( n556 , n5 , n1676 );
    or g1417 ( n1756 , n37 , n1623 );
    nor g1418 ( n1327 , n357 , n103 );
    or g1419 ( n166 , n1003 , n1019 );
    not g1420 ( n1168 , n1314 );
    xnor g1421 ( n732 , n1043 , n153 );
    or g1422 ( n362 , n914 , n1361 );
    not g1423 ( n1461 , n143 );
    not g1424 ( n265 , n105 );
    or g1425 ( n1432 , n925 , n227 );
    and g1426 ( n282 , n424 , n1332 );
    and g1427 ( n204 , n1568 , n1641 );
    or g1428 ( n810 , n809 , n939 );
    or g1429 ( n1440 , n1206 , n1446 );
    xnor g1430 ( n1573 , n0 , n986 );
    not g1431 ( n970 , n633 );
    xor g1432 ( n929 , n1182 , n179 );
    nor g1433 ( n822 , n584 , n1524 );
    not g1434 ( n1456 , n685 );
    and g1435 ( n1276 , n958 , n643 );
    or g1436 ( n1092 , n627 , n1563 );
    and g1437 ( n1479 , n1135 , n265 );
    nor g1438 ( n192 , n1422 , n697 );
    nor g1439 ( n981 , n1329 , n764 );
    and g1440 ( n1210 , n244 , n197 );
    xnor g1441 ( n614 , n49 , n5 );
    or g1442 ( n1217 , n996 , n448 );
    and g1443 ( n329 , n1720 , n1694 );
    or g1444 ( n959 , n1219 , n444 );
    and g1445 ( n1334 , n1380 , n901 );
    xnor g1446 ( n955 , n588 , n1501 );
    and g1447 ( n586 , n670 , n1317 );
    or g1448 ( n770 , n437 , n1247 );
    xnor g1449 ( n1662 , n741 , n1157 );
    xnor g1450 ( n79 , n799 , n1737 );
    buf g1451 ( n1234 , n608 );
    not g1452 ( n1692 , n1565 );
    xnor g1453 ( n473 , n1332 , n1071 );
    or g1454 ( n1739 , n399 , n70 );
    nor g1455 ( n1338 , n1535 , n813 );
    nor g1456 ( n590 , n629 , n1620 );
    buf g1457 ( n184 , n420 );
    xnor g1458 ( n1420 , n1232 , n1464 );
    nor g1459 ( n1712 , n960 , n191 );
    and g1460 ( n1300 , n7 , n1622 );
    xnor g1461 ( n311 , n777 , n1345 );
    xnor g1462 ( n979 , n1399 , n1412 );
    or g1463 ( n631 , n1124 , n280 );
    not g1464 ( n1444 , n359 );
    not g1465 ( n1706 , n789 );
    or g1466 ( n1202 , n1430 , n240 );
    not g1467 ( n1290 , n311 );
    and g1468 ( n664 , n63 , n4 );
    buf g1469 ( n30 , n362 );
    and g1470 ( n78 , n1190 , n677 );
    not g1471 ( n287 , n1446 );
    buf g1472 ( n337 , n626 );
    and g1473 ( n733 , n1350 , n530 );
    and g1474 ( n323 , n156 , n401 );
    nor g1475 ( n1447 , n1405 , n1463 );
    or g1476 ( n1372 , n803 , n430 );
    xnor g1477 ( n667 , n1642 , n750 );
    or g1478 ( n1524 , n68 , n1736 );
    or g1479 ( n1064 , n1257 , n802 );
    xnor g1480 ( n990 , n1694 , n412 );
    nor g1481 ( n563 , n1248 , n347 );
    not g1482 ( n1403 , n1383 );
    and g1483 ( n1295 , n1692 , n1062 );
    or g1484 ( n267 , n1401 , n1529 );
    or g1485 ( n1382 , n1514 , n749 );
    and g1486 ( n895 , n1315 , n1174 );
    or g1487 ( n1149 , n620 , n1721 );
    xnor g1488 ( n261 , n1550 , n397 );
    and g1489 ( n1183 , n249 , n1294 );
    or g1490 ( n1495 , n857 , n629 );
    xnor g1491 ( n248 , n623 , n1616 );
    xnor g1492 ( n185 , n632 , n1182 );
    not g1493 ( n806 , n815 );
    or g1494 ( n393 , n602 , n477 );
    or g1495 ( n382 , n1206 , n582 );
    nor g1496 ( n447 , n803 , n318 );
    xnor g1497 ( n1636 , n1535 , n1338 );
    or g1498 ( n64 , n1330 , n372 );
    and g1499 ( n1317 , n1692 , n1162 );
    xnor g1500 ( n233 , n1192 , n816 );
    and g1501 ( n691 , n532 , n1048 );
    nor g1502 ( n1163 , n608 , n1691 );
    or g1503 ( n33 , n927 , n619 );
    nor g1504 ( n365 , n6 , n967 );
    not g1505 ( n744 , n639 );
    or g1506 ( n286 , n1526 , n53 );
    xnor g1507 ( n410 , n418 , n955 );
    or g1508 ( n1409 , n549 , n343 );
    nor g1509 ( n1748 , n999 , n322 );
    and g1510 ( n865 , n1005 , n1363 );
    and g1511 ( n1344 , n366 , n642 );
    not g1512 ( n1052 , n43 );
    and g1513 ( n1481 , n1706 , n1679 );
    xnor g1514 ( n470 , n1682 , n1665 );
    and g1515 ( n1182 , n1255 , n1202 );
    nor g1516 ( n290 , n1700 , n1242 );
    not g1517 ( n1504 , n1642 );
    or g1518 ( n132 , n895 , n1068 );
    nor g1519 ( n350 , n257 , n609 );
    not g1520 ( n178 , n405 );
    or g1521 ( n109 , n206 , n1171 );
    or g1522 ( n1336 , n662 , n1532 );
    not g1523 ( n98 , n1462 );
    nor g1524 ( n699 , n1122 , n81 );
    or g1525 ( n668 , n317 , n805 );
    xnor g1526 ( n1109 , n1671 , n1589 );
    xnor g1527 ( n693 , n732 , n390 );
    xnor g1528 ( n385 , n864 , n540 );
    buf g1529 ( n1645 , n1446 );
    or g1530 ( n829 , n1721 , n381 );
    not g1531 ( n75 , n11 );
    or g1532 ( n170 , n1033 , n822 );
    or g1533 ( n503 , n1510 , n1232 );
    and g1534 ( n1140 , n155 , n803 );
    not g1535 ( n1360 , n643 );
    buf g1536 ( n1231 , n1470 );
    not g1537 ( n63 , n1565 );
    not g1538 ( n728 , n308 );
    not g1539 ( n864 , n991 );
    nor g1540 ( n1695 , n257 , n1626 );
    nor g1541 ( n1167 , n1132 , n544 );
    or g1542 ( n522 , n1402 , n649 );
    or g1543 ( n1022 , n1347 , n1081 );
    nor g1544 ( n485 , n1248 , n862 );
    or g1545 ( n67 , n1717 , n369 );
    and g1546 ( n872 , n691 , n901 );
    nor g1547 ( n514 , n1226 , n1344 );
    nor g1548 ( n933 , n572 , n519 );
    nor g1549 ( n1541 , n721 , n21 );
endmodule
