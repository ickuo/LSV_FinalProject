module top( n0 , n21 , n29 , n34 , n36 , n38 , n45 , n49 , n60 , 
n77 , n81 , n82 , n88 , n90 , n91 , n95 , n98 , n104 , n107 , 
n108 , n112 , n116 , n122 , n127 , n128 , n129 , n130 , n135 , n138 , 
n150 , n153 , n159 , n167 , n168 , n175 , n185 , n190 , n192 , n193 , 
n196 , n200 , n204 , n206 , n207 , n208 , n218 , n221 , n223 , n227 , 
n228 , n229 , n231 , n236 , n240 , n244 , n245 , n246 , n252 , n258 , 
n260 , n262 , n267 , n268 , n275 , n281 , n284 , n288 , n299 , n301 , 
n305 , n307 , n310 , n319 , n323 , n324 , n332 , n336 , n342 , n347 , 
n359 , n360 , n364 , n366 , n374 , n381 , n383 , n384 , n389 , n393 , 
n398 , n408 , n409 , n410 , n415 , n421 , n423 , n431 , n432 , n433 , 
n438 , n439 , n441 , n444 , n448 , n449 , n452 , n456 , n475 , n491 , 
n492 , n500 , n505 , n507 , n510 , n516 , n519 , n532 , n536 , n540 , 
n554 , n571 , n577 , n580 , n589 , n592 , n598 , n599 , n607 , n608 , 
n610 , n613 , n617 , n621 , n623 , n627 , n631 , n635 , n638 , n640 , 
n644 , n650 , n651 , n653 , n657 , n662 , n667 , n679 , n683 , n685 , 
n688 , n695 , n707 , n710 , n714 , n716 , n718 , n723 , n733 , n734 , 
n741 , n745 , n747 , n749 , n766 , n767 , n771 , n774 , n779 , n785 , 
n787 , n801 , n802 , n804 , n806 , n807 , n808 , n817 , n818 , n819 , 
n823 , n825 , n826 , n833 , n835 , n839 , n841 , n842 , n845 , n851 , 
n853 , n854 , n857 , n862 , n863 , n866 , n870 , n877 , n879 , n893 , 
n896 , n901 , n905 , n908 , n927 , n928 , n929 , n936 , n944 , n952 , 
n955 , n961 , n962 , n966 , n973 , n975 , n976 , n986 , n997 , n999 , 
n1005 , n1022 , n1023 , n1027 , n1029 , n1035 , n1036 , n1041 , n1044 , n1045 , 
n1048 , n1057 , n1059 , n1061 , n1064 , n1067 , n1069 , n1072 , n1073 , n1077 , 
n1080 , n1081 , n1085 , n1089 , n1091 , n1097 , n1098 , n1099 , n1120 , n1131 , 
n1132 , n1140 , n1141 , n1143 , n1146 , n1150 , n1151 , n1153 , n1163 , n1164 , 
n1178 , n1180 , n1184 , n1191 , n1194 , n1198 , n1202 , n1206 , n1219 , n1226 , 
n1229 , n1231 , n1232 , n1236 , n1239 , n1257 , n1259 , n1264 , n1269 , n1273 , 
n1277 , n1279 , n1288 , n1298 , n1301 , n1308 , n1311 , n1321 , n1326 , n1342 , 
n1344 , n1352 );
    input n0 , n21 , n36 , n38 , n45 , n49 , n77 , n95 , n98 , 
n104 , n107 , n108 , n116 , n122 , n127 , n128 , n138 , n153 , n192 , 
n196 , n200 , n208 , n221 , n231 , n236 , n244 , n245 , n246 , n252 , 
n258 , n260 , n262 , n267 , n268 , n281 , n284 , n288 , n301 , n305 , 
n310 , n319 , n323 , n324 , n332 , n336 , n359 , n360 , n364 , n366 , 
n381 , n384 , n393 , n398 , n421 , n423 , n431 , n433 , n438 , n439 , 
n441 , n444 , n448 , n449 , n475 , n491 , n500 , n505 , n507 , n510 , 
n519 , n532 , n536 , n540 , n571 , n577 , n589 , n599 , n610 , n631 , 
n635 , n640 , n644 , n650 , n657 , n667 , n685 , n688 , n695 , n714 , 
n716 , n741 , n745 , n749 , n766 , n767 , n771 , n774 , n787 , n802 , 
n804 , n806 , n818 , n819 , n823 , n825 , n826 , n833 , n839 , n841 , 
n845 , n851 , n857 , n862 , n863 , n866 , n870 , n879 , n893 , n896 , 
n901 , n928 , n929 , n936 , n944 , n952 , n955 , n961 , n975 , n976 , 
n986 , n997 , n1005 , n1022 , n1029 , n1035 , n1036 , n1041 , n1044 , n1045 , 
n1048 , n1064 , n1067 , n1069 , n1072 , n1073 , n1077 , n1080 , n1081 , n1089 , 
n1091 , n1097 , n1098 , n1120 , n1131 , n1132 , n1140 , n1141 , n1143 , n1146 , 
n1151 , n1163 , n1164 , n1180 , n1191 , n1198 , n1219 , n1226 , n1229 , n1231 , 
n1236 , n1257 , n1269 , n1273 , n1277 , n1279 , n1298 , n1308 , n1311 , n1321 , 
n1326 , n1342 , n1344 , n1352 ;
    output n29 , n34 , n60 , n81 , n82 , n88 , n90 , n91 , n112 , 
n129 , n130 , n135 , n150 , n159 , n167 , n168 , n175 , n185 , n190 , 
n193 , n204 , n206 , n207 , n218 , n223 , n227 , n228 , n229 , n240 , 
n275 , n299 , n307 , n342 , n347 , n374 , n383 , n389 , n408 , n409 , 
n410 , n415 , n432 , n452 , n456 , n492 , n516 , n554 , n580 , n592 , 
n598 , n607 , n608 , n613 , n617 , n621 , n623 , n627 , n638 , n651 , 
n653 , n662 , n679 , n683 , n707 , n710 , n718 , n723 , n733 , n734 , 
n747 , n779 , n785 , n801 , n807 , n808 , n817 , n835 , n842 , n853 , 
n854 , n877 , n905 , n908 , n927 , n962 , n966 , n973 , n999 , n1023 , 
n1027 , n1057 , n1059 , n1061 , n1085 , n1099 , n1150 , n1153 , n1178 , n1184 , 
n1194 , n1202 , n1206 , n1232 , n1239 , n1259 , n1264 , n1288 , n1301 ;
    wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
n20 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n30 , n31 , 
n32 , n33 , n35 , n37 , n39 , n40 , n41 , n42 , n43 , n44 , 
n46 , n47 , n48 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , 
n57 , n58 , n59 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , 
n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n78 , 
n79 , n80 , n83 , n84 , n85 , n86 , n87 , n89 , n92 , n93 , 
n94 , n96 , n97 , n99 , n100 , n101 , n102 , n103 , n105 , n106 , 
n109 , n110 , n111 , n113 , n114 , n115 , n117 , n118 , n119 , n120 , 
n121 , n123 , n124 , n125 , n126 , n131 , n132 , n133 , n134 , n136 , 
n137 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , 
n148 , n149 , n151 , n152 , n154 , n155 , n156 , n157 , n158 , n160 , 
n161 , n162 , n163 , n164 , n165 , n166 , n169 , n170 , n171 , n172 , 
n173 , n174 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , 
n184 , n186 , n187 , n188 , n189 , n191 , n194 , n195 , n197 , n198 , 
n199 , n201 , n202 , n203 , n205 , n209 , n210 , n211 , n212 , n213 , 
n214 , n215 , n216 , n217 , n219 , n220 , n222 , n224 , n225 , n226 , 
n230 , n232 , n233 , n234 , n235 , n237 , n238 , n239 , n241 , n242 , 
n243 , n247 , n248 , n249 , n250 , n251 , n253 , n254 , n255 , n256 , 
n257 , n259 , n261 , n263 , n264 , n265 , n266 , n269 , n270 , n271 , 
n272 , n273 , n274 , n276 , n277 , n278 , n279 , n280 , n282 , n283 , 
n285 , n286 , n287 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , 
n296 , n297 , n298 , n300 , n302 , n303 , n304 , n306 , n308 , n309 , 
n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n320 , n321 , 
n322 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n333 , n334 , 
n335 , n337 , n338 , n339 , n340 , n341 , n343 , n344 , n345 , n346 , 
n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , 
n358 , n361 , n362 , n363 , n365 , n367 , n368 , n369 , n370 , n371 , 
n372 , n373 , n375 , n376 , n377 , n378 , n379 , n380 , n382 , n385 , 
n386 , n387 , n388 , n390 , n391 , n392 , n394 , n395 , n396 , n397 , 
n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n411 , 
n412 , n413 , n414 , n416 , n417 , n418 , n419 , n420 , n422 , n424 , 
n425 , n426 , n427 , n428 , n429 , n430 , n434 , n435 , n436 , n437 , 
n440 , n442 , n443 , n445 , n446 , n447 , n450 , n451 , n453 , n454 , 
n455 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , 
n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n476 , 
n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , 
n487 , n488 , n489 , n490 , n493 , n494 , n495 , n496 , n497 , n498 , 
n499 , n501 , n502 , n503 , n504 , n506 , n508 , n509 , n511 , n512 , 
n513 , n514 , n515 , n517 , n518 , n520 , n521 , n522 , n523 , n524 , 
n525 , n526 , n527 , n528 , n529 , n530 , n531 , n533 , n534 , n535 , 
n537 , n538 , n539 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , 
n548 , n549 , n550 , n551 , n552 , n553 , n555 , n556 , n557 , n558 , 
n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , 
n569 , n570 , n572 , n573 , n574 , n575 , n576 , n578 , n579 , n581 , 
n582 , n583 , n584 , n585 , n586 , n587 , n588 , n590 , n591 , n593 , 
n594 , n595 , n596 , n597 , n600 , n601 , n602 , n603 , n604 , n605 , 
n606 , n609 , n611 , n612 , n614 , n615 , n616 , n618 , n619 , n620 , 
n622 , n624 , n625 , n626 , n628 , n629 , n630 , n632 , n633 , n634 , 
n636 , n637 , n639 , n641 , n642 , n643 , n645 , n646 , n647 , n648 , 
n649 , n652 , n654 , n655 , n656 , n658 , n659 , n660 , n661 , n663 , 
n664 , n665 , n666 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , 
n675 , n676 , n677 , n678 , n680 , n681 , n682 , n684 , n686 , n687 , 
n689 , n690 , n691 , n692 , n693 , n694 , n696 , n697 , n698 , n699 , 
n700 , n701 , n702 , n703 , n704 , n705 , n706 , n708 , n709 , n711 , 
n712 , n713 , n715 , n717 , n719 , n720 , n721 , n722 , n724 , n725 , 
n726 , n727 , n728 , n729 , n730 , n731 , n732 , n735 , n736 , n737 , 
n738 , n739 , n740 , n742 , n743 , n744 , n746 , n748 , n750 , n751 , 
n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , 
n762 , n763 , n764 , n765 , n768 , n769 , n770 , n772 , n773 , n775 , 
n776 , n777 , n778 , n780 , n781 , n782 , n783 , n784 , n786 , n788 , 
n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , 
n799 , n800 , n803 , n805 , n809 , n810 , n811 , n812 , n813 , n814 , 
n815 , n816 , n820 , n821 , n822 , n824 , n827 , n828 , n829 , n830 , 
n831 , n832 , n834 , n836 , n837 , n838 , n840 , n843 , n844 , n846 , 
n847 , n848 , n849 , n850 , n852 , n855 , n856 , n858 , n859 , n860 , 
n861 , n864 , n865 , n867 , n868 , n869 , n871 , n872 , n873 , n874 , 
n875 , n876 , n878 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , 
n887 , n888 , n889 , n890 , n891 , n892 , n894 , n895 , n897 , n898 , 
n899 , n900 , n902 , n903 , n904 , n906 , n907 , n909 , n910 , n911 , 
n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , 
n922 , n923 , n924 , n925 , n926 , n930 , n931 , n932 , n933 , n934 , 
n935 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n945 , n946 , 
n947 , n948 , n949 , n950 , n951 , n953 , n954 , n956 , n957 , n958 , 
n959 , n960 , n963 , n964 , n965 , n967 , n968 , n969 , n970 , n971 , 
n972 , n974 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , 
n985 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , 
n996 , n998 , n1000 , n1001 , n1002 , n1003 , n1004 , n1006 , n1007 , n1008 , 
n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , 
n1019 , n1020 , n1021 , n1024 , n1025 , n1026 , n1028 , n1030 , n1031 , n1032 , 
n1033 , n1034 , n1037 , n1038 , n1039 , n1040 , n1042 , n1043 , n1046 , n1047 , 
n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1058 , n1060 , 
n1062 , n1063 , n1065 , n1066 , n1068 , n1070 , n1071 , n1074 , n1075 , n1076 , 
n1078 , n1079 , n1082 , n1083 , n1084 , n1086 , n1087 , n1088 , n1090 , n1092 , 
n1093 , n1094 , n1095 , n1096 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , 
n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , 
n1116 , n1117 , n1118 , n1119 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , 
n1127 , n1128 , n1129 , n1130 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , 
n1139 , n1142 , n1144 , n1145 , n1147 , n1148 , n1149 , n1152 , n1154 , n1155 , 
n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1165 , n1166 , n1167 , 
n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , 
n1179 , n1181 , n1182 , n1183 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , 
n1192 , n1193 , n1195 , n1196 , n1197 , n1199 , n1200 , n1201 , n1203 , n1204 , 
n1205 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , 
n1216 , n1217 , n1218 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1227 , 
n1228 , n1230 , n1233 , n1234 , n1235 , n1237 , n1238 , n1240 , n1241 , n1242 , 
n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , 
n1253 , n1254 , n1255 , n1256 , n1258 , n1260 , n1261 , n1262 , n1263 , n1265 , 
n1266 , n1267 , n1268 , n1270 , n1271 , n1272 , n1274 , n1275 , n1276 , n1278 , 
n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1289 , n1290 , 
n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1299 , n1300 , n1302 , 
n1303 , n1304 , n1305 , n1306 , n1307 , n1309 , n1310 , n1312 , n1313 , n1314 , 
n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1322 , n1323 , n1324 , n1325 , 
n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , 
n1337 , n1338 , n1339 , n1340 , n1341 , n1343 , n1345 , n1346 , n1347 , n1348 , 
n1349 , n1350 , n1351 , n1353 ;
    or g0 ( n55 , n1004 , n1113 );
    or g1 ( n1107 , n1214 , n636 );
    not g2 ( n487 , n942 );
    and g3 ( n682 , n1332 , n147 );
    xor g4 ( n1004 , n1158 , n974 );
    xnor g5 ( n744 , n89 , n393 );
    not g6 ( n502 , n375 );
    nor g7 ( n471 , n643 , n52 );
    xnor g8 ( n1240 , n152 , n499 );
    and g9 ( n1303 , n846 , n153 );
    xnor g10 ( n1168 , n78 , n1156 );
    or g11 ( n894 , n449 , n497 );
    nor g12 ( n472 , n838 , n727 );
    buf g13 ( n638 , n1311 );
    not g14 ( n313 , n634 );
    or g15 ( n216 , n579 , n1320 );
    and g16 ( n854 , n243 , n647 );
    not g17 ( n1052 , n505 );
    and g18 ( n584 , n525 , n1324 );
    xnor g19 ( n721 , n920 , n501 );
    or g20 ( n356 , n1093 , n435 );
    buf g21 ( n683 , n381 );
    not g22 ( n756 , n514 );
    not g23 ( n217 , n951 );
    nor g24 ( n827 , n440 , n522 );
    nor g25 ( n42 , n301 , n1312 );
    or g26 ( n652 , n1198 , n403 );
    nor g27 ( n1100 , n1224 , n317 );
    and g28 ( n563 , n987 , n269 );
    nor g29 ( n1253 , n1225 , n697 );
    or g30 ( n996 , n205 , n541 );
    and g31 ( n732 , n985 , n528 );
    and g32 ( n1109 , n1076 , n687 );
    nor g33 ( n478 , n703 , n189 );
    or g34 ( n509 , n1300 , n981 );
    and g35 ( n840 , n692 , n238 );
    buf g36 ( n60 , n1081 );
    or g37 ( n184 , n1216 , n1275 );
    xnor g38 ( n254 , n955 , n851 );
    and g39 ( n932 , n456 , n574 );
    nor g40 ( n1315 , n571 , n1047 );
    not g41 ( n836 , n796 );
    not g42 ( n490 , n631 );
    nor g43 ( n1245 , n1081 , n1205 );
    or g44 ( n1082 , n496 , n670 );
    xor g45 ( n1332 , n1038 , n1311 );
    buf g46 ( n227 , 1'b0 );
    not g47 ( n469 , n601 );
    not g48 ( n220 , n1091 );
    buf g49 ( n415 , n997 );
    nor g50 ( n964 , n805 , n550 );
    xnor g51 ( n1150 , n1015 , n1350 );
    xnor g52 ( n765 , n1130 , n957 );
    not g53 ( n27 , n239 );
    xnor g54 ( n956 , n1290 , n889 );
    and g55 ( n671 , n1236 , n319 );
    not g56 ( n871 , n656 );
    xor g57 ( n941 , n1213 , n1081 );
    nor g58 ( n1290 , n254 , n815 );
    or g59 ( n377 , n1198 , n520 );
    nor g60 ( n719 , n1126 , n1313 );
    or g61 ( n1139 , n36 , n1317 );
    and g62 ( n459 , n1273 , n688 );
    xnor g63 ( n1006 , n472 , n765 );
    and g64 ( n152 , n502 , n591 );
    not g65 ( n51 , n52 );
    or g66 ( n690 , n1351 , n214 );
    or g67 ( n161 , n941 , n416 );
    xnor g68 ( n969 , n188 , n1095 );
    and g69 ( n279 , n871 , n1345 );
    not g70 ( n1280 , n330 );
    not g71 ( n443 , n177 );
    or g72 ( n1086 , n53 , n602 );
    or g73 ( n1026 , n584 , n1248 );
    buf g74 ( n29 , n1259 );
    xnor g75 ( n733 , n1108 , n744 );
    nor g76 ( n211 , n777 , n1313 );
    and g77 ( n698 , n471 , n995 );
    and g78 ( n382 , n1116 , n1307 );
    and g79 ( n653 , n717 , n939 );
    nor g80 ( n890 , n524 , n261 );
    or g81 ( n145 , n332 , n970 );
    not g82 ( n1250 , n688 );
    and g83 ( n614 , n1062 , n831 );
    xnor g84 ( n429 , n1123 , n535 );
    xor g85 ( n183 , n1222 , n47 );
    and g86 ( n927 , n824 , n1027 );
    or g87 ( n80 , n688 , n759 );
    or g88 ( n552 , n371 , n405 );
    buf g89 ( n229 , n785 );
    not g90 ( n1104 , n3 );
    xnor g91 ( n991 , n1349 , n138 );
    not g92 ( n1042 , n630 );
    and g93 ( n253 , n485 , n264 );
    buf g94 ( n1057 , n332 );
    not g95 ( n177 , n257 );
    xnor g96 ( n1106 , n821 , n440 );
    or g97 ( n568 , n716 , n891 );
    nor g98 ( n762 , n885 , n143 );
    or g99 ( n1203 , n40 , n660 );
    or g100 ( n125 , n663 , n1049 );
    or g101 ( n461 , n272 , n583 );
    and g102 ( n753 , n403 , n695 );
    xnor g103 ( n1142 , n508 , n1034 );
    or g104 ( n895 , n219 , n1157 );
    not g105 ( n701 , n585 );
    and g106 ( n861 , n269 , n446 );
    xnor g107 ( n998 , n1011 , n641 );
    xnor g108 ( n659 , n1248 , n20 );
    and g109 ( n1058 , n198 , n131 );
    xnor g110 ( n24 , n799 , n1200 );
    buf g111 ( n1049 , n680 );
    nor g112 ( n792 , n559 , n457 );
    xnor g113 ( n249 , n775 , n259 );
    and g114 ( n62 , n1337 , n9 );
    xnor g115 ( n570 , n292 , n1142 );
    nor g116 ( n830 , n757 , n813 );
    not g117 ( n118 , n418 );
    xnor g118 ( n704 , n1262 , n1211 );
    or g119 ( n1338 , n1020 , n1299 );
    xor g120 ( n66 , n438 , n1048 );
    and g121 ( n1305 , n1098 , n688 );
    and g122 ( n643 , n1109 , n474 );
    or g123 ( n1285 , n688 , n100 );
    and g124 ( n1216 , n947 , n928 );
    not g125 ( n1007 , n991 );
    and g126 ( n1254 , n1018 , n585 );
    or g127 ( n198 , n688 , n1092 );
    or g128 ( n696 , n811 , n16 );
    or g129 ( n1155 , n350 , n743 );
    nor g130 ( n921 , n1321 , n1205 );
    and g131 ( n75 , n1316 , n958 );
    and g132 ( n731 , n1050 , n1056 );
    and g133 ( n357 , n1049 , n863 );
    not g134 ( n117 , n1332 );
    xnor g135 ( n847 , n604 , n1238 );
    xnor g136 ( n700 , n341 , n396 );
    not g137 ( n210 , n297 );
    xnor g138 ( n1255 , n296 , n96 );
    xnor g139 ( n348 , n1189 , n1030 );
    nor g140 ( n1260 , n1186 , n725 );
    not g141 ( n176 , n208 );
    nor g142 ( n1137 , n909 , n75 );
    and g143 ( n224 , n846 , n1164 );
    xnor g144 ( n865 , n1323 , n270 );
    xnor g145 ( n634 , n1190 , n36 );
    buf g146 ( n492 , 1'b0 );
    xnor g147 ( n286 , n25 , n1340 );
    or g148 ( n561 , n427 , n968 );
    nor g149 ( n978 , n1319 , n1192 );
    and g150 ( n971 , n1171 , n1207 );
    nor g151 ( n590 , n788 , n14 );
    xnor g152 ( n1293 , n1349 , n1213 );
    not g153 ( n770 , n330 );
    or g154 ( n626 , n1271 , n798 );
    xnor g155 ( n1186 , n609 , n573 );
    nor g156 ( n764 , n1123 , n457 );
    not g157 ( n121 , n1326 );
    and g158 ( n628 , n814 , n281 );
    not g159 ( n680 , n688 );
    and g160 ( n1208 , n1171 , n552 );
    and g161 ( n602 , n1205 , n1269 );
    xnor g162 ( n306 , n247 , n948 );
    or g163 ( n946 , n1315 , n387 );
    xnor g164 ( n1178 , n634 , n840 );
    and g165 ( n9 , n690 , n28 );
    nor g166 ( n1112 , n900 , n392 );
    not g167 ( n1284 , n1325 );
    or g168 ( n593 , n688 , n19 );
    or g169 ( n1084 , n706 , n357 );
    xnor g170 ( n609 , n466 , n1117 );
    and g171 ( n195 , n1049 , n818 );
    buf g172 ( n973 , n819 );
    nor g173 ( n565 , n982 , n195 );
    not g174 ( n178 , n310 );
    not g175 ( n604 , n586 );
    not g176 ( n776 , n796 );
    nor g177 ( n1015 , n792 , n912 );
    or g178 ( n206 , n732 , n118 );
    not g179 ( n1018 , n47 );
    not g180 ( n19 , n245 );
    not g181 ( n815 , n1330 );
    and g182 ( n670 , n1254 , n1222 );
    xnor g183 ( n167 , n1280 , n394 );
    or g184 ( n1259 , n691 , n1183 );
    or g185 ( n1145 , n31 , n646 );
    not g186 ( n684 , n528 );
    and g187 ( n518 , n766 , n635 );
    buf g188 ( n608 , 1'b0 );
    buf g189 ( n307 , n1308 );
    not g190 ( n158 , n1069 );
    xnor g191 ( n1258 , n953 , n1155 );
    not g192 ( n1094 , n744 );
    or g193 ( n529 , n688 , n1212 );
    nor g194 ( n703 , n241 , n907 );
    not g195 ( n1317 , n1190 );
    or g196 ( n967 , n1270 , n253 );
    or g197 ( n859 , n688 , n1229 );
    not g198 ( n344 , n75 );
    xnor g199 ( n1016 , n974 , n659 );
    or g200 ( n951 , n178 , n403 );
    and g201 ( n1287 , n1176 , n975 );
    or g202 ( n465 , n772 , n693 );
    or g203 ( n648 , n888 , n614 );
    and g204 ( n112 , n116 , n1257 );
    not g205 ( n1021 , n1313 );
    not g206 ( n881 , n1058 );
    or g207 ( n988 , n1282 , n742 );
    xnor g208 ( n736 , n291 , n79 );
    xnor g209 ( n915 , n770 , n261 );
    and g210 ( n385 , n118 , n1147 );
    not g211 ( n910 , n75 );
    and g212 ( n715 , n417 , n139 );
    xnor g213 ( n511 , n566 , n589 );
    xnor g214 ( n523 , n443 , n231 );
    or g215 ( n460 , n45 , n846 );
    nor g216 ( n506 , n153 , n688 );
    or g217 ( n738 , n661 , n812 );
    not g218 ( n1012 , n965 );
    nor g219 ( n812 , n997 , n1049 );
    nor g220 ( n1159 , n1094 , n367 );
    xor g221 ( n1099 , n1325 , n515 );
    and g222 ( n168 , n597 , n453 );
    and g223 ( n397 , n52 , n1332 );
    or g224 ( n32 , n419 , n1166 );
    not g225 ( n583 , n214 );
    or g226 ( n30 , n1246 , n295 );
    and g227 ( n1087 , n688 , n1163 );
    not g228 ( n64 , n1073 );
    buf g229 ( n383 , n1321 );
    xnor g230 ( n783 , n1055 , n216 );
    and g231 ( n282 , n293 , n1139 );
    or g232 ( n450 , n447 , n636 );
    and g233 ( n878 , n300 , n1207 );
    and g234 ( n22 , n1140 , n688 );
    not g235 ( n191 , n0 );
    and g236 ( n1172 , n846 , n233 );
    not g237 ( n1271 , n1249 );
    or g238 ( n189 , n139 , n979 );
    not g239 ( n706 , n125 );
    or g240 ( n109 , n217 , n102 );
    or g241 ( n256 , n421 , n1205 );
    not g242 ( n520 , n354 );
    xnor g243 ( n1302 , n458 , n820 );
    and g244 ( n404 , n403 , n221 );
    not g245 ( n566 , n165 );
    or g246 ( n201 , n618 , n977 );
    xnor g247 ( n180 , n576 , n461 );
    and g248 ( n661 , n846 , n774 );
    or g249 ( n1050 , n945 , n464 );
    xnor g250 ( n654 , n84 , n564 );
    buf g251 ( n613 , n592 );
    xor g252 ( n1301 , n71 , n133 );
    and g253 ( n513 , n846 , n267 );
    buf g254 ( n185 , n571 );
    not g255 ( n788 , n393 );
    not g256 ( n624 , n1110 );
    nor g257 ( n902 , n1011 , n1079 );
    or g258 ( n615 , n17 , n935 );
    or g259 ( n334 , n850 , n1275 );
    or g260 ( n123 , n436 , n187 );
    nor g261 ( n1068 , n757 , n1278 );
    or g262 ( n501 , n65 , n911 );
    and g263 ( n737 , n901 , n688 );
    or g264 ( n361 , n1136 , n789 );
    and g265 ( n585 , n965 , n7 );
    not g266 ( n1312 , n895 );
    nor g267 ( n203 , n455 , n3 );
    not g268 ( n1328 , n833 );
    xor g269 ( n557 , n109 , n332 );
    or g270 ( n480 , n1347 , n182 );
    xnor g271 ( n413 , n923 , n763 );
    xnor g272 ( n687 , n56 , n571 );
    nor g273 ( n50 , n738 , n44 );
    and g274 ( n464 , n550 , n1101 );
    not g275 ( n126 , n67 );
    or g276 ( n1292 , n688 , n220 );
    and g277 ( n219 , n1045 , n688 );
    or g278 ( n1165 , n521 , n878 );
    or g279 ( n691 , n1002 , n1032 );
    or g280 ( n147 , n1311 , n83 );
    xnor g281 ( n270 , n174 , n678 );
    xnor g282 ( n1274 , n995 , n31 );
    xnor g283 ( n1218 , n41 , n735 );
    nor g284 ( n63 , n1019 , n696 );
    xnor g285 ( n170 , n938 , n1293 );
    not g286 ( n67 , n1031 );
    nor g287 ( n1060 , n1022 , n839 );
    xnor g288 ( n129 , n378 , n352 );
    not g289 ( n209 , n1084 );
    not g290 ( n549 , n761 );
    not g291 ( n498 , n117 );
    not g292 ( n1333 , n731 );
    or g293 ( n402 , n274 , n1245 );
    or g294 ( n131 , n191 , n1049 );
    not g295 ( n238 , n600 );
    or g296 ( n297 , n688 , n1179 );
    nor g297 ( n897 , n1035 , n846 );
    buf g298 ( n347 , n1342 );
    not g299 ( n805 , n1201 );
    xnor g300 ( n595 , n1310 , n1152 );
    not g301 ( n272 , n212 );
    nor g302 ( n406 , n138 , n1049 );
    and g303 ( n371 , n1205 , n423 );
    or g304 ( n171 , n271 , n921 );
    nor g305 ( n855 , n682 , n764 );
    nor g306 ( n1116 , n57 , n772 );
    or g307 ( n1000 , n1286 , n1275 );
    and g308 ( n1296 , n1051 , n1205 );
    not g309 ( n427 , n532 );
    or g310 ( n1028 , n571 , n403 );
    or g311 ( n1322 , n173 , n76 );
    or g312 ( n632 , n688 , n278 );
    not g313 ( n495 , n1270 );
    not g314 ( n100 , n893 );
    and g315 ( n1222 , n708 , n70 );
    nor g316 ( n748 , n1004 , n1026 );
    buf g317 ( n130 , n716 );
    not g318 ( n239 , n731 );
    and g319 ( n1353 , n431 , n688 );
    xnor g320 ( n391 , n114 , n860 );
    and g321 ( n533 , n263 , n339 );
    not g322 ( n37 , n445 );
    and g323 ( n809 , n1108 , n1159 );
    not g324 ( n587 , n1270 );
    or g325 ( n686 , n786 , n340 );
    not g326 ( n1329 , n1330 );
    and g327 ( n139 , n837 , n1055 );
    buf g328 ( n554 , n360 );
    nor g329 ( n1154 , n433 , n403 );
    nor g330 ( n816 , n589 , n165 );
    and g331 ( n586 , n125 , n1285 );
    xor g332 ( n1133 , n553 , n1335 );
    xnor g333 ( n1061 , n712 , n1145 );
    nor g334 ( n1010 , n890 , n382 );
    xnor g335 ( n1243 , n517 , n1261 );
    and g336 ( n999 , n484 , n518 );
    xnor g337 ( n477 , n39 , n1274 );
    buf g338 ( n82 , n104 );
    or g339 ( n87 , n1105 , n276 );
    or g340 ( n417 , n729 , n110 );
    and g341 ( n993 , n364 , n688 );
    or g342 ( n938 , n232 , n404 );
    nor g343 ( n1 , n467 , n315 );
    not g344 ( n666 , n686 );
    or g345 ( n115 , n1322 , n395 );
    or g346 ( n837 , n222 , n588 );
    xnor g347 ( n1030 , n1158 , n1065 );
    or g348 ( n1055 , n539 , n512 );
    xnor g349 ( n1235 , n575 , n1122 );
    xnor g350 ( n909 , n180 , n1240 );
    not g351 ( n1252 , n849 );
    nor g352 ( n26 , n152 , n1054 );
    xnor g353 ( n1090 , n876 , n420 );
    not g354 ( n673 , n694 );
    not g355 ( n205 , n645 );
    and g356 ( n810 , n610 , n688 );
    xnor g357 ( n1126 , n622 , n298 );
    not g358 ( n390 , n317 );
    xnor g359 ( n775 , n37 , n287 );
    or g360 ( n25 , n746 , n210 );
    and g361 ( n134 , n213 , n1294 );
    xnor g362 ( n1281 , n601 , n881 );
    and g363 ( n1105 , n1204 , n501 );
    or g364 ( n488 , n454 , n282 );
    and g365 ( n900 , n1172 , n1020 );
    or g366 ( n1083 , n45 , n829 );
    and g367 ( n1276 , n836 , n749 );
    or g368 ( n47 , n358 , n285 );
    xnor g369 ( n90 , n442 , n375 );
    xnor g370 ( n889 , n343 , n639 );
    nor g371 ( n422 , n439 , n1329 );
    or g372 ( n1350 , n1187 , n1137 );
    xnor g373 ( n1319 , n1134 , n637 );
    xnor g374 ( n149 , n895 , n793 );
    and g375 ( n1175 , n988 , n953 );
    not g376 ( n326 , n71 );
    or g377 ( n280 , n1311 , n846 );
    xnor g378 ( n1211 , n294 , n904 );
    or g379 ( n70 , n567 , n796 );
    or g380 ( n1066 , n800 , n403 );
    not g381 ( n761 , n313 );
    not g382 ( n790 , n95 );
    and g383 ( n1283 , n280 , n632 );
    or g384 ( n755 , n1228 , n6 );
    and g385 ( n556 , n336 , n384 );
    nor g386 ( n17 , n339 , n263 );
    not g387 ( n462 , n612 );
    nor g388 ( n1334 , n37 , n141 );
    xor g389 ( n1223 , n583 , n576 );
    nor g390 ( n697 , n212 , n345 );
    and g391 ( n1088 , n688 , n252 );
    and g392 ( n954 , n124 , n168 );
    or g393 ( n317 , n1195 , n437 );
    or g394 ( n234 , n944 , n596 );
    or g395 ( n907 , n867 , n762 );
    and g396 ( n752 , n444 , n688 );
    not g397 ( n187 , n1242 );
    not g398 ( n213 , n304 );
    or g399 ( n821 , n993 , n404 );
    not g400 ( n309 , n685 );
    or g401 ( n7 , n1052 , n796 );
    not g402 ( n822 , n944 );
    not g403 ( n940 , n268 );
    not g404 ( n656 , n946 );
    nor g405 ( n15 , n136 , n1071 );
    or g406 ( n779 , n494 , n33 );
    not g407 ( n18 , n511 );
    not g408 ( n832 , n416 );
    not g409 ( n1185 , n482 );
    nor g410 ( n980 , n1109 , n946 );
    not g411 ( n784 , n761 );
    xnor g412 ( n906 , n376 , n120 );
    not g413 ( n481 , n1158 );
    and g414 ( n1201 , n1205 , n328 );
    or g415 ( n645 , n22 , n1268 );
    and g416 ( n1286 , n776 , n217 );
    and g417 ( n1074 , n403 , n741 );
    or g418 ( n674 , n289 , n30 );
    or g419 ( n367 , n1166 , n144 );
    or g420 ( n1056 , n997 , n209 );
    or g421 ( n54 , n58 , n414 );
    nor g422 ( n709 , n589 , n846 );
    or g423 ( n926 , n688 , n616 );
    or g424 ( n1196 , n688 , n176 );
    not g425 ( n257 , n1000 );
    xor g426 ( n1247 , n587 , n1040 );
    not g427 ( n1336 , n196 );
    not g428 ( n965 , n1148 );
    and g429 ( n850 , n814 , n507 );
    and g430 ( n639 , n1330 , n66 );
    or g431 ( n750 , n132 , n514 );
    and g432 ( n232 , n1191 , n688 );
    or g433 ( n199 , n557 , n473 );
    and g434 ( n350 , n403 , n540 );
    xnor g435 ( n672 , n682 , n980 );
    or g436 ( n186 , n688 , n1336 );
    or g437 ( n785 , n385 , n99 );
    not g438 ( n1267 , n620 );
    xnor g439 ( n658 , n291 , n619 );
    not g440 ( n970 , n109 );
    not g441 ( n1031 , n724 );
    or g442 ( n1129 , n701 , n711 );
    and g443 ( n1187 , n1121 , n2 );
    or g444 ( n76 , n873 , n478 );
    buf g445 ( n207 , n1198 );
    not g446 ( n913 , n3 );
    not g447 ( n1349 , n412 );
    or g448 ( n295 , n542 , n1181 );
    buf g449 ( n580 , n449 );
    and g450 ( n739 , n476 , n996 );
    xnor g451 ( n1059 , n553 , n302 );
    buf g452 ( n223 , 1'b0 );
    xnor g453 ( n607 , n1039 , n1253 );
    xnor g454 ( n375 , n601 , n104 );
    not g455 ( n553 , n875 );
    and g456 ( n1054 , n1121 , n591 );
    not g457 ( n503 , n510 );
    xnor g458 ( n303 , n626 , n780 );
    or g459 ( n1266 , n234 , n751 );
    not g460 ( n89 , n527 );
    or g461 ( n525 , n688 , n1125 );
    buf g462 ( n91 , n1259 );
    xnor g463 ( n948 , n1144 , n998 );
    nor g464 ( n1209 , n475 , n846 );
    and g465 ( n271 , n1205 , n1279 );
    xor g466 ( n942 , n356 , n1321 );
    not g467 ( n1130 , n313 );
    buf g468 ( n846 , n680 );
    buf g469 ( n853 , n589 );
    nor g470 ( n84 , n688 , n726 );
    or g471 ( n56 , n963 , n843 );
    xnor g472 ( n780 , n1124 , n794 );
    xnor g473 ( n793 , n356 , n105 );
    not g474 ( n1037 , n562 );
    not g475 ( n315 , n157 );
    or g476 ( n485 , n514 , n894 );
    xnor g477 ( n1239 , n1043 , n855 );
    xnor g478 ( n120 , n831 , n339 );
    xnor g479 ( n803 , n1118 , n837 );
    or g480 ( n136 , n1017 , n11 );
    not g481 ( n197 , n451 );
    not g482 ( n1121 , n344 );
    xnor g483 ( n1202 , n511 , n62 );
    not g484 ( n179 , n480 );
    and g485 ( n538 , n1129 , n47 );
    not g486 ( n1108 , n913 );
    and g487 ( n1246 , n1001 , n920 );
    nor g488 ( n53 , n381 , n846 );
    not g489 ( n947 , n796 );
    or g490 ( n340 , n1185 , n582 );
    xnor g491 ( n372 , n720 , n321 );
    and g492 ( n572 , n629 , n501 );
    not g493 ( n798 , n630 );
    xnor g494 ( n799 , n79 , n426 );
    or g495 ( n174 , n166 , n1303 );
    buf g496 ( n175 , n138 );
    and g497 ( n773 , n1205 , n77 );
    or g498 ( n354 , n119 , n430 );
    xor g499 ( n97 , n655 , n915 );
    and g500 ( n515 , n1267 , n670 );
    and g501 ( n867 , n369 , n1167 );
    and g502 ( n582 , n142 , n1094 );
    nor g503 ( n1002 , n1233 , n250 );
    or g504 ( n578 , n1008 , n13 );
    not g505 ( n437 , n322 );
    or g506 ( n751 , n454 , n784 );
    xnor g507 ( n882 , n72 , n795 );
    not g508 ( n106 , n1333 );
    not g509 ( n418 , n730 );
    or g510 ( n1278 , n611 , n164 );
    xnor g511 ( n1085 , n694 , n464 );
    and g512 ( n689 , n142 , n1114 );
    buf g513 ( n374 , 1'b0 );
    or g514 ( n786 , n581 , n285 );
    not g515 ( n534 , n720 );
    xor g516 ( n1189 , n1167 , n1309 );
    or g517 ( n376 , n43 , n984 );
    or g518 ( n3 , n917 , n887 );
    not g519 ( n1212 , n1077 );
    not g520 ( n442 , n910 );
    not g521 ( n600 , n234 );
    nor g522 ( n717 , n308 , n54 );
    or g523 ( n1340 , n983 , n753 );
    xor g524 ( n1169 , n881 , n360 );
    and g525 ( n222 , n846 , n441 );
    not g526 ( n304 , n834 );
    not g527 ( n497 , n361 );
    xnor g528 ( n71 , n462 , n38 );
    not g529 ( n33 , n711 );
    or g530 ( n226 , n1081 , n73 );
    not g531 ( n265 , n365 );
    xnor g532 ( n923 , n391 , n722 );
    and g533 ( n241 , n101 , n171 );
    not g534 ( n290 , n796 );
    xnor g535 ( n1162 , n946 , n429 );
    or g536 ( n992 , n644 , n1205 );
    and g537 ( n172 , n544 , n1217 );
    nor g538 ( n758 , n1100 , n79 );
    not g539 ( n1033 , n796 );
    and g540 ( n486 , n1205 , n857 );
    not g541 ( n1310 , n326 );
    xnor g542 ( n289 , n94 , n1155 );
    buf g543 ( n1153 , n231 );
    not g544 ( n1251 , n557 );
    or g545 ( n1177 , n1087 , n316 );
    not g546 ( n454 , n71 );
    and g547 ( n1020 , n1205 , n790 );
    buf g548 ( n1264 , n116 );
    xnor g549 ( n702 , n265 , n1010 );
    not g550 ( n655 , n1014 );
    nor g551 ( n1265 , n360 , n1049 );
    and g552 ( n746 , n745 , n688 );
    or g553 ( n1197 , n943 , n1205 );
    or g554 ( n52 , n42 , n279 );
    and g555 ( n165 , n322 , n728 );
    or g556 ( n1316 , n942 , n1348 );
    or g557 ( n740 , n1078 , n630 );
    xnor g558 ( n58 , n407 , n700 );
    and g559 ( n248 , n1263 , n1309 );
    or g560 ( n934 , n950 , n897 );
    nor g561 ( n242 , n303 , n731 );
    not g562 ( n1123 , n147 );
    or g563 ( n341 , n1136 , n753 );
    not g564 ( n188 , n255 );
    not g565 ( n829 , n938 );
    and g566 ( n1327 , n1097 , n688 );
    and g567 ( n924 , n315 , n1109 );
    and g568 ( n983 , n1044 , n688 );
    and g569 ( n85 , n408 , n817 );
    or g570 ( n591 , n104 , n469 );
    not g571 ( n849 , n1169 );
    or g572 ( n218 , n545 , n538 );
    not g573 ( n368 , n67 );
    xnor g574 ( n1345 , n895 , n301 );
    nor g575 ( n163 , n268 , n403 );
    nor g576 ( n235 , n1209 , n160 );
    or g577 ( n1192 , n24 , n1295 );
    not g578 ( n1092 , n1132 );
    xor g579 ( n111 , n151 , n1248 );
    or g580 ( n445 , n1025 , n1275 );
    and g581 ( n6 , n830 , n333 );
    not g582 ( n1125 , n323 );
    not g583 ( n164 , n1155 );
    not g584 ( n151 , n584 );
    nor g585 ( n318 , n1147 , n349 );
    xnor g586 ( n575 , n504 , n672 );
    or g587 ( n1188 , n1351 , n212 );
    buf g588 ( n842 , n1184 );
    and g589 ( n243 , n448 , n870 );
    not g590 ( n74 , n1079 );
    or g591 ( n333 , n338 , n1256 );
    xor g592 ( n483 , n754 , n991 );
    nor g593 ( n337 , n919 , n590 );
    and g594 ( n269 , n740 , n1083 );
    xnor g595 ( n1103 , n154 , n834 );
    and g596 ( n824 , n954 , n854 );
    and g597 ( n1119 , n1110 , n1307 );
    and g598 ( n4 , n827 , n821 );
    xnor g599 ( n576 , n1039 , n511 );
    not g600 ( n1233 , n1352 );
    not g601 ( n642 , n340 );
    and g602 ( n1330 , n708 , n947 );
    xnor g603 ( n325 , n380 , n400 );
    xnor g604 ( n5 , n1019 , n304 );
    nor g605 ( n388 , n132 , n509 );
    xnor g606 ( n931 , n777 , n194 );
    xnor g607 ( n20 , n1283 , n903 );
    not g608 ( n995 , n498 );
    and g609 ( n1289 , n543 , n971 );
    or g610 ( n293 , n549 , n692 );
    nor g611 ( n352 , n1215 , n428 );
    nand g612 ( n1176 , n1022 , n839 );
    and g613 ( n1306 , n290 , n936 );
    and g614 ( n99 , n299 , n349 );
    and g615 ( n1299 , n1287 , n1233 );
    nor g616 ( n496 , n701 , n1254 );
    not g617 ( n943 , n650 );
    nor g618 ( n266 , n874 , n876 );
    not g619 ( n1268 , n1285 );
    xnor g620 ( n1323 , n1190 , n462 );
    xnor g621 ( n251 , n922 , n286 );
    not g622 ( n754 , n782 );
    buf g623 ( n1275 , n1148 );
    not g624 ( n162 , n582 );
    not g625 ( n772 , n261 );
    xnor g626 ( n396 , n775 , n933 );
    buf g627 ( n403 , n1250 );
    or g628 ( n1001 , n1314 , n406 );
    nor g629 ( n778 , n689 , n531 );
    or g630 ( n1224 , n773 , n709 );
    or g631 ( n1166 , n1000 , n445 );
    not g632 ( n114 , n187 );
    and g633 ( n1076 , n669 , n255 );
    or g634 ( n541 , n664 , n50 );
    not g635 ( n31 , n51 );
    xnor g636 ( n757 , n953 , n988 );
    nor g637 ( n463 , n1115 , n113 );
    buf g638 ( n1205 , n1250 );
    not g639 ( n14 , n1104 );
    nor g640 ( n409 , n633 , n318 );
    and g641 ( n1237 , n110 , n216 );
    or g642 ( n1337 , n994 , n442 );
    xor g643 ( n562 , n361 , n449 );
    not g644 ( n782 , n941 );
    xnor g645 ( n641 , n660 , n1046 );
    not g646 ( n72 , n832 );
    not g647 ( n569 , n172 );
    and g648 ( n629 , n1106 , n555 );
    or g649 ( n299 , n1352 , n730 );
    xor g650 ( n194 , n557 , n523 );
    or g651 ( n1034 , n1272 , n242 );
    nor g652 ( n379 , n1289 , n300 );
    or g653 ( n601 , n459 , n512 );
    and g654 ( n887 , n465 , n468 );
    and g655 ( n618 , n436 , n368 );
    not g656 ( n1291 , n390 );
    not g657 ( n1213 , n73 );
    xnor g658 ( n559 , n1162 , n1173 );
    and g659 ( n228 , n238 , n883 );
    xnor g660 ( n308 , n372 , n149 );
    xnor g661 ( n1173 , n188 , n477 );
    not g662 ( n1307 , n655 );
    xnor g663 ( n573 , n645 , n181 );
    and g664 ( n581 , n776 , n1298 );
    or g665 ( n1038 , n737 , n675 );
    and g666 ( n1256 , n561 , n857 );
    xnor g667 ( n1039 , n720 , n107 );
    xnor g668 ( n1117 , n821 , n721 );
    buf g669 ( n342 , n299 );
    and g670 ( n10 , n424 , n86 );
    buf g671 ( n596 , n1201 );
    or g672 ( n953 , n224 , n46 );
    and g673 ( n864 , n846 , n246 );
    not g674 ( n886 , n648 );
    xnor g675 ( n292 , n480 , n1035 );
    xnor g676 ( n296 , n425 , n546 );
    xnor g677 ( n504 , n1009 , n353 );
    and g678 ( n1160 , n1161 , n677 );
    xnor g679 ( n922 , n1207 , n949 );
    or g680 ( n230 , n688 , n121 );
    and g681 ( n918 , n1242 , n1266 );
    xnor g682 ( n694 , n1084 , n997 );
    and g683 ( n888 , n294 , n376 );
    not g684 ( n985 , n1241 );
    buf g685 ( n516 , n301 );
    nor g686 ( n405 , n449 , n403 );
    or g687 ( n322 , n688 , n490 );
    nor g688 ( n373 , n1124 , n8 );
    and g689 ( n791 , n305 , n688 );
    not g690 ( n1078 , n508 );
    or g691 ( n456 , n215 , n115 );
    and g692 ( n789 , n846 , n841 );
    not g693 ( n977 , n681 );
    nor g694 ( n369 , n603 , n248 );
    not g695 ( n435 , n146 );
    or g696 ( n1228 , n1341 , n1127 );
    and g697 ( n489 , n1219 , n688 );
    or g698 ( n1217 , n1035 , n179 );
    or g699 ( n225 , n63 , n1165 );
    and g700 ( n950 , n846 , n929 );
    not g701 ( n378 , n365 );
    not g702 ( n436 , n751 );
    xnor g703 ( n1171 , n1340 , n660 );
    or g704 ( n1325 , n848 , n285 );
    or g705 ( n1127 , n4 , n87 );
    and g706 ( n214 , n872 , n61 );
    and g707 ( n419 , n937 , n788 );
    and g708 ( n1314 , n1049 , n1120 );
    and g709 ( n844 , n403 , n1229 );
    or g710 ( n676 , n346 , n715 );
    and g711 ( n1204 , n629 , n402 );
    or g712 ( n544 , n1331 , n563 );
    and g713 ( n440 , n460 , n363 );
    or g714 ( n302 , n871 , n924 );
    and g715 ( n560 , n1013 , n392 );
    nor g716 ( n588 , n104 , n403 );
    xnor g717 ( n904 , n184 , n1135 );
    xnor g718 ( n1046 , n565 , n552 );
    not g719 ( n669 , n498 );
    xor g720 ( n820 , n402 , n1001 );
    or g721 ( n335 , n107 , n1049 );
    not g722 ( n1149 , n1076 );
    or g723 ( n291 , n1305 , n844 );
    or g724 ( n276 , n35 , n769 );
    or g725 ( n446 , n1078 , n1249 );
    not g726 ( n1215 , n473 );
    or g727 ( n416 , n138 , n412 );
    buf g728 ( n617 , n598 );
    and g729 ( n1309 , n146 , n1197 );
    xnor g730 ( n637 , n664 , n1090 );
    or g731 ( n528 , n1276 , n1275 );
    or g732 ( n781 , n1308 , n1049 );
    and g733 ( n817 , n1260 , n493 );
    nor g734 ( n215 , n1160 , n451 );
    and g735 ( n1027 , n671 , n1221 );
    and g736 ( n974 , n1028 , n926 );
    not g737 ( n742 , n529 );
    not g738 ( n712 , n487 );
    and g739 ( n660 , n992 , n230 );
    nor g740 ( n370 , n1249 , n27 );
    not g741 ( n699 , n1345 );
    not g742 ( n1148 , n237 );
    xor g743 ( n858 , n126 , n282 );
    and g744 ( n545 , n1267 , n1254 );
    or g745 ( n868 , n38 , n612 );
    not g746 ( n59 , n1041 );
    and g747 ( n412 , n125 , n80 );
    not g748 ( n1110 , n1021 );
    not g749 ( n524 , n1346 );
    xnor g750 ( n81 , n495 , n351 );
    and g751 ( n994 , n9 , n1188 );
    or g752 ( n451 , n1283 , n55 );
    or g753 ( n883 , n822 , n805 );
    not g754 ( n801 , n385 );
    and g755 ( n1241 , n515 , n1284 );
    buf g756 ( n159 , 1'b0 );
    not g757 ( n558 , n687 );
    xnor g758 ( n508 , n938 , n45 );
    and g759 ( n182 , n403 , n1072 );
    xnor g760 ( n726 , n1022 , n839 );
    not g761 ( n287 , n786 );
    xnor g762 ( n298 , n587 , n97 );
    xnor g763 ( n808 , n106 , n991 );
    buf g764 ( n285 , n1296 );
    or g765 ( n979 , n140 , n914 );
    buf g766 ( n877 , n679 );
    not g767 ( n1263 , n171 );
    and g768 ( n166 , n688 , n128 );
    xor g769 ( n1156 , n422 , n41 );
    nor g770 ( n1071 , n1175 , n1068 );
    and g771 ( n1221 , n1029 , n952 );
    not g772 ( n551 , n239 );
    not g773 ( n875 , n1095 );
    buf g774 ( n410 , 1'b0 );
    nor g775 ( n1318 , n234 , n549 );
    xnor g776 ( n627 , n524 , n624 );
    xnor g777 ( n144 , n775 , n393 );
    xnor g778 ( n1096 , n1130 , n596 );
    or g779 ( n872 , n1252 , n380 );
    and g780 ( n720 , n256 , n859 );
    xnor g781 ( n96 , n770 , n702 );
    and g782 ( n1242 , n488 , n868 );
    nor g783 ( n574 , n560 , n379 );
    or g784 ( n1324 , n537 , n1049 );
    and g785 ( n358 , n836 , n398 );
    xnor g786 ( n311 , n960 , n1086 );
    or g787 ( n813 , n136 , n674 );
    not g788 ( n620 , n33 );
    xnor g789 ( n722 , n673 , n858 );
    and g790 ( n860 , n968 , n940 );
    nor g791 ( n960 , n163 , n486 );
    nor g792 ( n92 , n481 , n974 );
    and g793 ( n1282 , n1080 , n688 );
    not g794 ( n1348 , n1145 );
    and g795 ( n110 , n12 , n797 );
    xor g796 ( n259 , n1185 , n419 );
    nor g797 ( n1008 , n247 , n137 );
    xnor g798 ( n1261 , n94 , n988 );
    xnor g799 ( n420 , n311 , n1258 );
    and g800 ( n79 , n335 , n1196 );
    and g801 ( n1070 , n985 , n1218 );
    and g802 ( n1009 , n1335 , n1149 );
    xnor g803 ( n962 , n941 , n373 );
    and g804 ( n1195 , n823 , n688 );
    or g805 ( n1032 , n1112 , n605 );
    xnor g806 ( n707 , n523 , n465 );
    not g807 ( n1075 , n591 );
    and g808 ( n729 , n12 , n216 );
    nor g809 ( n48 , n434 , n273 );
    xor g810 ( n939 , n1174 , n847 );
    xor g811 ( n1304 , n1252 , n375 );
    or g812 ( n61 , n360 , n1058 );
    or g813 ( n531 , n809 , n203 );
    xnor g814 ( n78 , n528 , n1325 );
    buf g815 ( n193 , n644 );
    and g816 ( n647 , n324 , n577 );
    and g817 ( n597 , n1344 , n802 );
    nor g818 ( n912 , n1235 , n172 );
    or g819 ( n351 , n1040 , n211 );
    nor g820 ( n425 , n388 , n1343 );
    or g821 ( n432 , n976 , n127 );
    not g822 ( n69 , n1005 );
    not g823 ( n233 , n866 );
    or g824 ( n1313 , n816 , n1210 );
    or g825 ( n903 , n169 , n513 );
    not g826 ( n914 , n417 );
    nor g827 ( n386 , n376 , n294 );
    xnor g828 ( n795 , n269 , n483 );
    xnor g829 ( n835 , n687 , n990 );
    not g830 ( n711 , n666 );
    xnor g831 ( n1065 , n151 , n1297 );
    not g832 ( n1346 , n1014 );
    not g833 ( n616 , n1131 );
    not g834 ( n981 , n473 );
    nor g835 ( n86 , n386 , n760 );
    not g836 ( n675 , n1161 );
    xnor g837 ( n1230 , n1019 , n811 );
    xnor g838 ( n2 , n1223 , n325 );
    xnor g839 ( n493 , n658 , n348 );
    not g840 ( n1014 , n562 );
    xnor g841 ( n530 , n603 , n1016 );
    and g842 ( n1093 , n826 , n688 );
    xnor g843 ( n362 , n101 , n171 );
    and g844 ( n880 , n846 , n309 );
    and g845 ( n395 , n705 , n755 );
    nor g846 ( n892 , n1160 , n55 );
    or g847 ( n327 , n1308 , n586 );
    not g848 ( n1181 , n713 );
    not g849 ( n1351 , n1039 );
    or g850 ( n294 , n628 , n1275 );
    and g851 ( n1019 , n186 , n470 );
    nor g852 ( n394 , n989 , n1119 );
    or g853 ( n314 , n301 , n1049 );
    not g854 ( n103 , n262 );
    xnor g855 ( n499 , n1304 , n994 );
    not g856 ( n154 , n869 );
    and g857 ( n1157 , n1049 , n879 );
    not g858 ( n278 , n258 );
    not g859 ( n1184 , n862 );
    buf g860 ( n623 , 1'b0 );
    not g861 ( n919 , n177 );
    and g862 ( n664 , n781 , n1102 );
    xnor g863 ( n621 , n126 , n918 );
    not g864 ( n989 , n894 );
    or g865 ( n1170 , n724 , n114 );
    not g866 ( n625 , n80 );
    xor g867 ( n41 , n1227 , n183 );
    not g868 ( n665 , n1224 );
    not g869 ( n567 , n986 );
    xnor g870 ( n1238 , n1084 , n865 );
    xnor g871 ( n622 , n899 , n931 );
    not g872 ( n283 , n108 );
    xnor g873 ( n564 , n1172 , n235 );
    buf g874 ( n796 , n556 );
    or g875 ( n1190 , n752 , n1074 );
    not g876 ( n157 , n569 );
    or g877 ( n1193 , n1111 , n719 );
    xnor g878 ( n546 , n468 , n1247 );
    or g879 ( n339 , n688 , n804 );
    buf g880 ( n807 , n45 );
    xor g881 ( n1270 , n407 , n716 );
    nor g882 ( n273 , n944 , n93 );
    and g883 ( n1335 , n649 , n377 );
    or g884 ( n13 , n648 , n925 );
    or g885 ( n1102 , n688 , n1328 );
    not g886 ( n550 , n977 );
    buf g887 ( n710 , n36 );
    or g888 ( n713 , n572 , n1204 );
    not g889 ( n937 , n527 );
    not g890 ( n39 , n558 );
    and g891 ( n1183 , n932 , n155 );
    or g892 ( n401 , n688 , n69 );
    nor g893 ( n916 , n533 , n578 );
    or g894 ( n677 , n64 , n1049 );
    and g895 ( n155 , n10 , n886 );
    not g896 ( n547 , n1180 );
    xnor g897 ( n105 , n23 , n856 );
    and g898 ( n681 , n1170 , n327 );
    and g899 ( n428 , n1119 , n1300 );
    and g900 ( n1011 , n331 , n593 );
    nor g901 ( n1115 , n596 , n784 );
    buf g902 ( n1232 , n268 );
    not g903 ( n312 , n341 );
    nor g904 ( n760 , n831 , n1062 );
    or g905 ( n470 , n972 , n846 );
    and g906 ( n473 , n967 , n568 );
    and g907 ( n843 , n1205 , n200 );
    or g908 ( n204 , n337 , n141 );
    or g909 ( n728 , n547 , n1049 );
    not g910 ( n458 , n934 );
    and g911 ( n646 , n924 , n474 );
    xnor g912 ( n414 , n334 , n1168 );
    and g913 ( n543 , n74 , n479 );
    and g914 ( n930 , n85 , n653 );
    and g915 ( n1300 , n1280 , n495 );
    or g916 ( n831 , n688 , n519 );
    and g917 ( n1138 , n846 , n260 );
    and g918 ( n963 , n1036 , n688 );
    or g919 ( n202 , n111 , n189 );
    or g920 ( n263 , n1306 , n1275 );
    xnor g921 ( n619 , n1291 , n783 );
    not g922 ( n40 , n1340 );
    nor g923 ( n982 , n819 , n846 );
    and g924 ( n848 , n1033 , n896 );
    nor g925 ( n542 , n920 , n1001 );
    or g926 ( n1167 , n668 , n1157 );
    xnor g927 ( n1297 , n1160 , n1107 );
    not g928 ( n876 , n738 );
    and g929 ( n141 , n162 , n937 );
    buf g930 ( n1194 , n116 );
    not g931 ( n349 , n730 );
    not g932 ( n814 , n796 );
    xnor g933 ( n662 , n508 , n277 );
    and g934 ( n73 , n548 , n1066 );
    or g935 ( n1161 , n688 , n1024 );
    and g936 ( n453 , n288 , n359 );
    and g937 ( n1025 , n290 , n599 );
    xnor g938 ( n1295 , n906 , n306 );
    not g939 ( n611 , n94 );
    xor g940 ( n11 , n874 , n738 );
    not g941 ( n468 , n523 );
    or g942 ( n150 , n642 , n1334 );
    and g943 ( n579 , n657 , n688 );
    xnor g944 ( n747 , n1169 , n26 );
    not g945 ( n972 , n806 );
    or g946 ( n1062 , n329 , n285 );
    or g947 ( n331 , n716 , n403 );
    nor g948 ( n1210 , n18 , n62 );
    xnor g949 ( n320 , n798 , n882 );
    not g950 ( n759 , n845 );
    xnor g951 ( n455 , n89 , n249 );
    or g952 ( n958 , n1321 , n594 );
    nor g953 ( n16 , n1294 , n213 );
    and g954 ( n261 , n199 , n145 );
    not g955 ( n1320 , n198 );
    or g956 ( n363 , n688 , n503 );
    and g957 ( n539 , n1064 , n688 );
    xnor g958 ( n763 , n681 , n1199 );
    xnor g959 ( n181 , n44 , n1243 );
    xor g960 ( n1128 , n1167 , n603 );
    and g961 ( n12 , n736 , n1234 );
    not g962 ( n1047 , n56 );
    nor g963 ( n838 , n596 , n123 );
    not g964 ( n355 , n1151 );
    and g965 ( n484 , n21 , n1226 );
    nor g966 ( n1220 , n397 , n698 );
    and g967 ( n1343 , n899 , n562 );
    not g968 ( n83 , n1038 );
    xor g969 ( n400 , n9 , n1304 );
    and g970 ( n668 , n366 , n688 );
    and g971 ( n408 , n978 , n654 );
    nor g972 ( n743 , n36 , n1205 );
    and g973 ( n316 , n1049 , n1143 );
    or g974 ( n1294 , n864 , n884 );
    not g975 ( n237 , n1296 );
    not g976 ( n537 , n98 );
    and g977 ( n274 , n403 , n1141 );
    and g978 ( n346 , n1291 , n1224 );
    or g979 ( n1003 , n332 , n846 );
    or g980 ( n735 , n1082 , n686 );
    and g981 ( n160 , n1205 , n1231 );
    or g982 ( n389 , n515 , n68 );
    and g983 ( n693 , n428 , n265 );
    and g984 ( n1053 , n1033 , n771 );
    and g985 ( n447 , n688 , n767 );
    not g986 ( n692 , n860 );
    xnor g987 ( n135 , n669 , n172 );
    or g988 ( n28 , n107 , n534 );
    or g989 ( n94 , n1353 , n1074 );
    nor g990 ( n411 , n1203 , n1063 );
    xnor g991 ( n1199 , n1310 , n1096 );
    buf g992 ( n908 , n801 );
    not g993 ( n527 , n257 );
    xor g994 ( n1234 , n317 , n1118 );
    xnor g995 ( n1200 , n1263 , n530 );
    nor g996 ( n68 , n1222 , n545 );
    and g997 ( n512 , n1205 , n536 );
    not g998 ( n1051 , n796 );
    and g999 ( n8 , n106 , n416 );
    xnor g1000 ( n1134 , n440 , n1302 );
    or g1001 ( n212 , n502 , n1169 );
    not g1002 ( n1063 , n543 );
    nor g1003 ( n885 , n92 , n748 );
    xnor g1004 ( n1017 , n205 , n664 );
    nor g1005 ( n343 , n768 , n815 );
    xnor g1006 ( n1174 , n480 , n170 );
    not g1007 ( n365 , n1251 );
    not g1008 ( n594 , n356 );
    nor g1009 ( n35 , n399 , n458 );
    nor g1010 ( n1111 , n1255 , n624 );
    not g1011 ( n457 , n157 );
    buf g1012 ( n452 , n393 );
    and g1013 ( n1182 , n902 , n25 );
    nor g1014 ( n338 , n532 , n880 );
    or g1015 ( n173 , n1237 , n676 );
    nor g1016 ( n476 , n266 , n15 );
    or g1017 ( n143 , n1128 , n362 );
    and g1018 ( n156 , n1146 , n688 );
    not g1019 ( n1179 , n825 );
    xnor g1020 ( n633 , n78 , n1070 );
    buf g1021 ( n1288 , n1035 );
    and g1022 ( n727 , n391 , n596 );
    not g1023 ( n137 , n184 );
    not g1024 ( n869 , n1294 );
    not g1025 ( n113 , n282 );
    not g1026 ( n102 , n186 );
    nor g1027 ( n917 , n231 , n443 );
    or g1028 ( n725 , n956 , n704 );
    xor g1029 ( n935 , n247 , n184 );
    or g1030 ( n598 , n127 , n606 );
    nor g1031 ( n140 , n1055 , n837 );
    xnor g1032 ( n957 , n368 , n526 );
    not g1033 ( n142 , n1104 );
    and g1034 ( n329 , n1051 , n284 );
    xor g1035 ( n353 , n558 , n942 );
    and g1036 ( n65 , n714 , n688 );
    and g1037 ( n43 , n403 , n640 );
    or g1038 ( n1101 , n724 , n1266 );
    and g1039 ( n603 , n314 , n401 );
    buf g1040 ( n1206 , 1'b0 );
    and g1041 ( n1124 , n72 , n1007 );
    xnor g1042 ( n240 , n48 , n570 );
    or g1043 ( n1207 , n810 , n789 );
    xnor g1044 ( n535 , n712 , n1133 );
    nor g1045 ( n46 , n38 , n1049 );
    not g1046 ( n1147 , n1352 );
    nor g1047 ( n1214 , n1067 , n403 );
    xor g1048 ( n514 , n341 , n644 );
    xnor g1049 ( n1152 , n673 , n463 );
    not g1050 ( n777 , n253 );
    nor g1051 ( n1244 , n596 , n201 );
    xnor g1052 ( n856 , n354 , n56 );
    not g1053 ( n1095 , n1345 );
    nand g1054 ( n606 , n787 , n491 );
    buf g1055 ( n34 , n116 );
    xnor g1056 ( n555 , n399 , n934 );
    and g1057 ( n968 , n1049 , n685 );
    not g1058 ( n399 , n466 );
    or g1059 ( n920 , n791 , n625 );
    buf g1060 ( n275 , n1277 );
    and g1061 ( n387 , n467 , n39 );
    and g1062 ( n769 , n713 , n1246 );
    or g1063 ( n649 , n147 , n1043 );
    not g1064 ( n1331 , n292 );
    buf g1065 ( n88 , 1'b0 );
    not g1066 ( n1227 , n585 );
    not g1067 ( n874 , n44 );
    not g1068 ( n1339 , n667 );
    xnor g1069 ( n23 , n1038 , n450 );
    or g1070 ( n987 , n861 , n551 );
    xor g1071 ( n899 , n981 , n989 );
    and g1072 ( n612 , n529 , n148 );
    xnor g1073 ( n905 , n1227 , n686 );
    nor g1074 ( n424 , n533 , n615 );
    xnor g1075 ( n321 , n566 , n1281 );
    nor g1076 ( n605 , n560 , n916 );
    and g1077 ( n124 , n930 , n999 );
    and g1078 ( n891 , n951 , n297 );
    nor g1079 ( n526 , n964 , n1244 );
    or g1080 ( n146 , n688 , n158 );
    or g1081 ( n1158 , n1327 , n843 );
    buf g1082 ( n1023 , n38 );
    and g1083 ( n250 , n1060 , n975 );
    and g1084 ( n630 , n161 , n226 );
    or g1085 ( n548 , n688 , n355 );
    xnor g1086 ( n1122 , n1220 , n969 );
    xnor g1087 ( n828 , n361 , n1177 );
    xnor g1088 ( n898 , n109 , n828 );
    xnor g1089 ( n479 , n25 , n1011 );
    not g1090 ( n1136 , n951 );
    nor g1091 ( n169 , n1342 , n1205 );
    not g1092 ( n945 , n694 );
    or g1093 ( n1013 , n1172 , n1338 );
    xnor g1094 ( n517 , n880 , n506 );
    not g1095 ( n800 , n961 );
    or g1096 ( n1249 , n754 , n1007 );
    not g1097 ( n380 , n1075 );
    not g1098 ( n679 , n385 );
    and g1099 ( n730 , n1241 , n684 );
    and g1100 ( n873 , n758 , n291 );
    not g1101 ( n1118 , n665 );
    xor g1102 ( n724 , n604 , n1308 );
    xnor g1103 ( n794 , n483 , n861 );
    xnor g1104 ( n723 , n292 , n563 );
    or g1105 ( n133 , n1318 , n113 );
    not g1106 ( n101 , n1309 );
    or g1107 ( n521 , n134 , n1182 );
    not g1108 ( n430 , n525 );
    xnor g1109 ( n190 , n778 , n1193 );
    not g1110 ( n330 , n756 );
    or g1111 ( n990 , n1009 , n1 );
    not g1112 ( n663 , n122 );
    xor g1113 ( n1144 , n154 , n811 );
    and g1114 ( n119 , n236 , n688 );
    or g1115 ( n1079 , n1230 , n1103 );
    and g1116 ( n247 , n1205 , n1339 );
    not g1117 ( n132 , n1037 );
    or g1118 ( n705 , n892 , n197 );
    or g1119 ( n797 , n1138 , n1265 );
    buf g1120 ( n651 , n1184 );
    or g1121 ( n148 , n283 , n1049 );
    xnor g1122 ( n1135 , n1062 , n263 );
    and g1123 ( n300 , n543 , n1208 );
    and g1124 ( n1272 , n551 , n320 );
    and g1125 ( n434 , n413 , n944 );
    or g1126 ( n392 , n796 , n1299 );
    not g1127 ( n911 , n548 );
    not g1128 ( n345 , n344 );
    xnor g1129 ( n93 , n595 , n1006 );
    and g1130 ( n1040 , n253 , n750 );
    xor g1131 ( n768 , n49 , n244 );
    nor g1132 ( n884 , n231 , n1205 );
    xnor g1133 ( n426 , n797 , n803 );
    or g1134 ( n592 , n127 , n59 );
    xnor g1135 ( n255 , n354 , n1198 );
    not g1136 ( n1225 , n214 );
    or g1137 ( n949 , n1154 , n316 );
    xor g1138 ( n933 , n919 , n898 );
    xnor g1139 ( n328 , n940 , n685 );
    nor g1140 ( n984 , n393 , n1049 );
    buf g1141 ( n718 , n116 );
    buf g1142 ( n734 , n475 );
    or g1143 ( n834 , n1053 , n1275 );
    or g1144 ( n1113 , n143 , n202 );
    xnor g1145 ( n1262 , n251 , n5 );
    or g1146 ( n466 , n489 , n182 );
    not g1147 ( n482 , n1166 );
    and g1148 ( n1347 , n1089 , n688 );
    not g1149 ( n708 , n1012 );
    or g1150 ( n44 , n156 , n357 );
    not g1151 ( n1024 , n500 );
    not g1152 ( n474 , n699 );
    and g1153 ( n1114 , n32 , n144 );
    nor g1154 ( n277 , n1042 , n370 );
    not g1155 ( n407 , n891 );
    nor g1156 ( n494 , n287 , n642 );
    and g1157 ( n636 , n403 , n192 );
    or g1158 ( n264 , n644 , n312 );
    or g1159 ( n678 , n1088 , n968 );
    not g1160 ( n1043 , n255 );
    nor g1161 ( n522 , n934 , n466 );
    nor g1162 ( n1341 , n739 , n30 );
    or g1163 ( n852 , n688 , n103 );
    and g1164 ( n1248 , n652 , n852 );
    or g1165 ( n959 , n411 , n225 );
    and g1166 ( n57 , n1300 , n378 );
    and g1167 ( n925 , n959 , n155 );
    buf g1168 ( n966 , n107 );
    not g1169 ( n467 , n1335 );
    and g1170 ( n811 , n1003 , n1292 );
endmodule
