module top( n1 , n2 , n3 , n5 , n6 , n9 , n11 , n14 , n16 , 
n18 , n20 , n26 , n27 , n29 , n38 , n40 , n42 , n44 , n48 , 
n54 , n56 , n59 , n60 , n64 , n67 , n71 , n72 , n74 , n76 , 
n81 , n82 , n85 , n86 , n92 , n93 , n94 , n96 , n101 , n102 , 
n103 , n108 , n109 , n111 , n113 , n114 , n115 , n116 , n120 , n123 , 
n125 , n129 , n131 , n132 , n133 , n134 , n137 , n138 , n139 , n140 , 
n143 , n144 , n145 , n147 , n150 , n153 , n154 , n156 , n157 , n158 , 
n161 , n162 , n163 , n164 , n166 , n171 , n174 , n176 , n178 , n179 , 
n182 , n183 , n187 , n188 , n192 , n193 , n195 , n196 , n200 , n202 , 
n203 , n204 , n206 , n207 , n209 , n210 , n213 , n215 , n217 , n219 , 
n220 , n224 , n225 , n226 , n233 , n234 , n237 , n239 , n242 , n245 , 
n247 , n248 , n251 , n252 , n254 , n256 , n257 , n263 , n268 , n274 , 
n278 , n279 , n281 , n282 , n284 , n286 , n288 , n290 , n291 , n294 , 
n295 , n299 , n300 , n304 , n313 , n314 , n317 , n326 , n329 , n330 , 
n336 , n340 , n342 , n343 , n344 , n345 , n346 , n348 , n349 , n357 , 
n358 , n359 , n360 , n363 , n365 , n368 , n370 , n371 , n375 , n378 , 
n383 , n385 , n387 , n388 , n393 , n394 , n395 , n398 , n399 , n403 , 
n404 , n406 , n407 , n409 , n410 , n411 , n416 , n426 , n429 , n432 , 
n437 , n438 , n440 , n443 , n444 , n446 , n448 , n449 , n452 , n453 , 
n454 , n456 , n459 , n460 , n461 , n462 , n463 , n464 , n470 , n474 , 
n475 , n477 , n479 , n481 , n482 , n484 , n486 , n488 , n491 , n492 , 
n499 , n500 , n502 , n506 , n507 , n509 , n511 , n512 , n516 , n517 , 
n522 , n525 , n526 , n530 , n533 , n534 , n535 , n536 , n537 , n542 , 
n544 , n552 , n553 , n554 , n555 , n556 , n560 , n564 , n565 , n570 , 
n573 , n577 , n578 , n580 , n585 , n587 , n590 , n591 , n593 , n594 , 
n595 , n597 , n598 , n608 , n611 , n613 , n615 , n619 , n622 , n623 , 
n625 , n626 , n631 , n633 , n636 , n637 , n639 , n640 , n644 , n645 , 
n647 , n651 , n652 , n657 , n658 , n659 , n660 , n661 , n662 , n665 , 
n667 , n679 , n680 , n682 , n687 , n688 , n705 , n707 , n711 , n713 , 
n716 , n717 , n718 , n722 , n726 , n727 , n728 , n729 , n731 , n735 , 
n739 , n746 , n750 , n751 , n755 , n758 , n759 , n760 , n766 , n767 , 
n770 , n771 , n772 , n773 , n774 , n778 , n779 , n780 , n783 , n784 , 
n786 , n787 , n788 , n789 , n790 , n791 , n794 , n795 , n796 , n797 , 
n798 , n800 , n805 , n807 , n812 , n813 , n815 , n817 , n821 , n826 , 
n827 , n828 , n829 , n832 , n834 , n835 , n836 , n839 , n840 , n844 , 
n845 , n850 , n851 , n852 , n853 , n855 , n856 , n861 , n864 , n866 , 
n867 , n868 , n870 , n875 , n885 , n887 , n888 , n890 , n892 , n893 , 
n894 , n895 , n898 , n900 );
    input n1 , n2 , n3 , n9 , n14 , n18 , n20 , n27 , n29 , 
n38 , n40 , n42 , n44 , n48 , n59 , n60 , n64 , n71 , n72 , 
n81 , n85 , n86 , n93 , n96 , n103 , n111 , n114 , n115 , n123 , 
n129 , n131 , n132 , n133 , n137 , n138 , n139 , n143 , n144 , n145 , 
n147 , n154 , n156 , n157 , n158 , n162 , n163 , n164 , n166 , n171 , 
n174 , n178 , n179 , n182 , n183 , n187 , n188 , n192 , n202 , n203 , 
n206 , n209 , n210 , n215 , n224 , n225 , n237 , n242 , n247 , n248 , 
n251 , n252 , n263 , n274 , n278 , n284 , n286 , n290 , n291 , n294 , 
n295 , n299 , n304 , n313 , n317 , n326 , n330 , n342 , n343 , n345 , 
n348 , n357 , n358 , n359 , n360 , n365 , n368 , n370 , n371 , n375 , 
n378 , n383 , n387 , n388 , n393 , n395 , n398 , n399 , n403 , n404 , 
n409 , n410 , n411 , n429 , n438 , n440 , n443 , n444 , n446 , n448 , 
n449 , n454 , n456 , n459 , n460 , n461 , n463 , n464 , n474 , n477 , 
n482 , n486 , n488 , n491 , n500 , n507 , n516 , n522 , n525 , n526 , 
n535 , n542 , n544 , n552 , n553 , n554 , n555 , n556 , n564 , n585 , 
n587 , n591 , n594 , n595 , n597 , n598 , n608 , n611 , n613 , n622 , 
n623 , n625 , n626 , n631 , n633 , n636 , n639 , n645 , n651 , n652 , 
n657 , n658 , n659 , n660 , n661 , n665 , n667 , n680 , n682 , n687 , 
n688 , n707 , n713 , n722 , n727 , n728 , n729 , n731 , n739 , n759 , 
n766 , n767 , n770 , n771 , n774 , n778 , n780 , n783 , n784 , n786 , 
n787 , n789 , n791 , n794 , n796 , n797 , n798 , n807 , n812 , n813 , 
n817 , n821 , n826 , n827 , n828 , n832 , n834 , n840 , n844 , n852 , 
n855 , n856 , n864 , n866 , n867 , n868 , n870 , n875 , n887 , n888 , 
n890 , n892 , n894 , n900 ;
    output n5 , n6 , n11 , n16 , n26 , n54 , n56 , n67 , n74 , 
n76 , n82 , n92 , n94 , n101 , n102 , n108 , n109 , n113 , n116 , 
n120 , n125 , n134 , n140 , n150 , n153 , n161 , n176 , n193 , n195 , 
n196 , n200 , n204 , n207 , n213 , n217 , n219 , n220 , n226 , n233 , 
n234 , n239 , n245 , n254 , n256 , n257 , n268 , n279 , n281 , n282 , 
n288 , n300 , n314 , n329 , n336 , n340 , n344 , n346 , n349 , n363 , 
n385 , n394 , n406 , n407 , n416 , n426 , n432 , n437 , n452 , n453 , 
n462 , n470 , n475 , n479 , n481 , n484 , n492 , n499 , n502 , n506 , 
n509 , n511 , n512 , n517 , n530 , n533 , n534 , n536 , n537 , n560 , 
n565 , n570 , n573 , n577 , n578 , n580 , n590 , n593 , n615 , n619 , 
n637 , n640 , n644 , n647 , n662 , n679 , n705 , n711 , n716 , n717 , 
n718 , n726 , n735 , n746 , n750 , n751 , n755 , n758 , n760 , n772 , 
n773 , n779 , n788 , n790 , n795 , n800 , n805 , n815 , n829 , n835 , 
n836 , n839 , n845 , n850 , n851 , n853 , n861 , n885 , n893 , n895 , 
n898 ;
    wire n0 , n4 , n7 , n8 , n10 , n12 , n13 , n15 , n17 , 
n19 , n21 , n22 , n23 , n24 , n25 , n28 , n30 , n31 , n32 , 
n33 , n34 , n35 , n36 , n37 , n39 , n41 , n43 , n45 , n46 , 
n47 , n49 , n50 , n51 , n52 , n53 , n55 , n57 , n58 , n61 , 
n62 , n63 , n65 , n66 , n68 , n69 , n70 , n73 , n75 , n77 , 
n78 , n79 , n80 , n83 , n84 , n87 , n88 , n89 , n90 , n91 , 
n95 , n97 , n98 , n99 , n100 , n104 , n105 , n106 , n107 , n110 , 
n112 , n117 , n118 , n119 , n121 , n122 , n124 , n126 , n127 , n128 , 
n130 , n135 , n136 , n141 , n142 , n146 , n148 , n149 , n151 , n152 , 
n155 , n159 , n160 , n165 , n167 , n168 , n169 , n170 , n172 , n173 , 
n175 , n177 , n180 , n181 , n184 , n185 , n186 , n189 , n190 , n191 , 
n194 , n197 , n198 , n199 , n201 , n205 , n208 , n211 , n212 , n214 , 
n216 , n218 , n221 , n222 , n223 , n227 , n228 , n229 , n230 , n231 , 
n232 , n235 , n236 , n238 , n240 , n241 , n243 , n244 , n246 , n249 , 
n250 , n253 , n255 , n258 , n259 , n260 , n261 , n262 , n264 , n265 , 
n266 , n267 , n269 , n270 , n271 , n272 , n273 , n275 , n276 , n277 , 
n280 , n283 , n285 , n287 , n289 , n292 , n293 , n296 , n297 , n298 , 
n301 , n302 , n303 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , 
n312 , n315 , n316 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , 
n325 , n327 , n328 , n331 , n332 , n333 , n334 , n335 , n337 , n338 , 
n339 , n341 , n347 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , 
n361 , n362 , n364 , n366 , n367 , n369 , n372 , n373 , n374 , n376 , 
n377 , n379 , n380 , n381 , n382 , n384 , n386 , n389 , n390 , n391 , 
n392 , n396 , n397 , n400 , n401 , n402 , n405 , n408 , n412 , n413 , 
n414 , n415 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , 
n425 , n427 , n428 , n430 , n431 , n433 , n434 , n435 , n436 , n439 , 
n441 , n442 , n445 , n447 , n450 , n451 , n455 , n457 , n458 , n465 , 
n466 , n467 , n468 , n469 , n471 , n472 , n473 , n476 , n478 , n480 , 
n483 , n485 , n487 , n489 , n490 , n493 , n494 , n495 , n496 , n497 , 
n498 , n501 , n503 , n504 , n505 , n508 , n510 , n513 , n514 , n515 , 
n518 , n519 , n520 , n521 , n523 , n524 , n527 , n528 , n529 , n531 , 
n532 , n538 , n539 , n540 , n541 , n543 , n545 , n546 , n547 , n548 , 
n549 , n550 , n551 , n557 , n558 , n559 , n561 , n562 , n563 , n566 , 
n567 , n568 , n569 , n571 , n572 , n574 , n575 , n576 , n579 , n581 , 
n582 , n583 , n584 , n586 , n588 , n589 , n592 , n596 , n599 , n600 , 
n601 , n602 , n603 , n604 , n605 , n606 , n607 , n609 , n610 , n612 , 
n614 , n616 , n617 , n618 , n620 , n621 , n624 , n627 , n628 , n629 , 
n630 , n632 , n634 , n635 , n638 , n641 , n642 , n643 , n646 , n648 , 
n649 , n650 , n653 , n654 , n655 , n656 , n663 , n664 , n666 , n668 , 
n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , 
n681 , n683 , n684 , n685 , n686 , n689 , n690 , n691 , n692 , n693 , 
n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , 
n704 , n706 , n708 , n709 , n710 , n712 , n714 , n715 , n719 , n720 , 
n721 , n723 , n724 , n725 , n730 , n732 , n733 , n734 , n736 , n737 , 
n738 , n740 , n741 , n742 , n743 , n744 , n745 , n747 , n748 , n749 , 
n752 , n753 , n754 , n756 , n757 , n761 , n762 , n763 , n764 , n765 , 
n768 , n769 , n775 , n776 , n777 , n781 , n782 , n785 , n792 , n793 , 
n799 , n801 , n802 , n803 , n804 , n806 , n808 , n809 , n810 , n811 , 
n814 , n816 , n818 , n819 , n820 , n822 , n823 , n824 , n825 , n830 , 
n831 , n833 , n837 , n838 , n841 , n842 , n843 , n846 , n847 , n848 , 
n849 , n854 , n857 , n858 , n859 , n860 , n862 , n863 , n865 , n869 , 
n871 , n872 , n873 , n874 , n876 , n877 , n878 , n879 , n880 , n881 , 
n882 , n883 , n884 , n886 , n889 , n891 , n896 , n897 , n899 , n901 , 
n902 , n903 ;
    or g0 ( n630 , n892 , n540 );
    buf g1 ( n573 , n665 );
    or g2 ( n405 , n610 , n417 );
    or g3 ( n605 , n862 , n354 );
    not g4 ( n830 , n105 );
    buf g5 ( n340 , n533 );
    buf g6 ( n394 , n252 );
    buf g7 ( n850 , n48 );
    and g8 ( n271 , n263 , n209 );
    not g9 ( n420 , n896 );
    or g10 ( n689 , n778 , n420 );
    nor g11 ( n649 , n203 , n287 );
    or g12 ( n549 , n287 , n650 );
    xnor g13 ( n308 , n546 , n880 );
    not g14 ( n571 , n701 );
    or g15 ( n124 , n556 , n141 );
    nor g16 ( n246 , n465 , n264 );
    nor g17 ( n376 , n645 , n663 );
    or g18 ( n140 , n841 , n232 );
    not g19 ( n353 , n681 );
    or g20 ( n301 , n307 , n26 );
    not g21 ( n110 , n673 );
    or g22 ( n884 , n883 , n769 );
    and g23 ( n312 , n186 , n642 );
    and g24 ( n668 , n373 , n606 );
    or g25 ( n471 , n876 , n604 );
    nor g26 ( n341 , n2 , n579 );
    and g27 ( n505 , n710 , n553 );
    and g28 ( n10 , n138 , n892 );
    nor g29 ( n841 , n639 , n236 );
    nor g30 ( n208 , n71 , n75 );
    buf g31 ( n895 , n81 );
    nor g32 ( n819 , n597 , n155 );
    buf g33 ( n204 , n360 );
    xnor g34 ( n331 , n285 , n32 );
    or g35 ( n168 , n238 , n241 );
    nor g36 ( n238 , n278 , n88 );
    nor g37 ( n442 , n415 , n762 );
    and g38 ( n829 , n401 , n879 );
    xnor g39 ( n377 , n614 , n330 );
    nor g40 ( n824 , n727 , n392 );
    and g41 ( n666 , n755 , n309 );
    nor g42 ( n401 , n328 , n276 );
    not g43 ( n802 , n379 );
    and g44 ( n414 , n818 , n731 );
    nor g45 ( n351 , n749 , n47 );
    not g46 ( n540 , n730 );
    or g47 ( n106 , n843 , n77 );
    not g48 ( n790 , n343 );
    buf g49 ( n861 , n375 );
    not g50 ( n142 , n188 );
    xnor g51 ( n592 , n620 , n369 );
    not g52 ( n122 , n601 );
    not g53 ( n673 , n271 );
    nor g54 ( n352 , n561 , n858 );
    not g55 ( n476 , n56 );
    not g56 ( n296 , n100 );
    and g57 ( n696 , n689 , n531 );
    buf g58 ( n288 , n342 );
    nor g59 ( n741 , n203 , n220 );
    buf g60 ( n492 , n474 );
    and g61 ( n776 , n357 , n892 );
    nor g62 ( n52 , n359 , n541 );
    buf g63 ( n74 , n739 );
    or g64 ( n699 , n483 , n521 );
    nor g65 ( n223 , n135 , n361 );
    nor g66 ( n754 , n624 , n70 );
    xnor g67 ( n185 , n724 , n731 );
    xnor g68 ( n177 , n842 , n794 );
    or g69 ( n434 , n809 , n686 );
    or g70 ( n160 , n167 , n367 );
    buf g71 ( n735 , n502 );
    not g72 ( n654 , n255 );
    nor g73 ( n519 , n553 , n119 );
    and g74 ( n581 , n422 , n569 );
    not g75 ( n26 , n696 );
    not g76 ( n569 , n263 );
    and g77 ( n799 , n398 , n892 );
    not g78 ( n857 , n35 );
    and g79 ( n677 , n444 , n203 );
    nor g80 ( n136 , n115 , n199 );
    nor g81 ( n761 , n687 , n99 );
    buf g82 ( n101 , n866 );
    not g83 ( n382 , n534 );
    buf g84 ( n407 , n174 );
    xnor g85 ( n275 , n603 , n17 );
    or g86 ( n337 , n664 , n222 );
    xnor g87 ( n806 , n765 , n600 );
    nor g88 ( n431 , n410 , n364 );
    or g89 ( n79 , n404 , n145 );
    not g90 ( n697 , n731 );
    nor g91 ( n781 , n892 , n748 );
    buf g92 ( n716 , n123 );
    buf g93 ( n795 , n274 );
    xnor g94 ( n333 , n12 , n34 );
    xnor g95 ( n632 , n236 , n572 );
    not g96 ( n572 , n191 );
    not g97 ( n269 , n586 );
    buf g98 ( n679 , n158 );
    buf g99 ( n314 , n564 );
    and g100 ( n702 , n51 , n373 );
    not g101 ( n426 , n491 );
    buf g102 ( n537 , n187 );
    nor g103 ( n265 , n383 , n802 );
    nor g104 ( n897 , n230 , n323 );
    nor g105 ( n465 , n157 , n654 );
    not g106 ( n374 , n779 );
    or g107 ( n435 , n602 , n8 );
    nor g108 ( n457 , n61 , n311 );
    or g109 ( n836 , n699 , n43 );
    xnor g110 ( n212 , n553 , n114 );
    or g111 ( n533 , n690 , n53 );
    buf g112 ( n11 , n544 );
    nor g113 ( n588 , n744 , n435 );
    and g114 ( n39 , n756 , n764 );
    or g115 ( n126 , n667 , n823 );
    and g116 ( n63 , n240 , n639 );
    buf g117 ( n213 , n680 );
    xnor g118 ( n903 , n89 , n889 );
    not g119 ( n97 , n151 );
    nor g120 ( n367 , n313 , n244 );
    and g121 ( n683 , n836 , n822 );
    or g122 ( n229 , n504 , n152 );
    buf g123 ( n746 , n284 );
    nor g124 ( n306 , n443 , n388 );
    not g125 ( n748 , n808 );
    and g126 ( n493 , n607 , n794 );
    not g127 ( n321 , n567 );
    not g128 ( n530 , n829 );
    and g129 ( n871 , n672 , n513 );
    not g130 ( n503 , n737 );
    and g131 ( n437 , n433 , n104 );
    xor g132 ( n788 , n315 , n33 );
    not g133 ( n176 , n667 );
    xor g134 ( n578 , n742 , n592 );
    nor g135 ( n814 , n111 , n280 );
    nor g136 ( n551 , n657 , n121 );
    or g137 ( n231 , n761 , n871 );
    xnor g138 ( n380 , n145 , n330 );
    nor g139 ( n642 , n260 , n596 );
    buf g140 ( n835 , n680 );
    or g141 ( n319 , n824 , n265 );
    nor g142 ( n527 , n289 , n159 );
    and g143 ( n876 , n36 , n334 );
    not g144 ( n4 , n446 );
    and g145 ( n362 , n532 , n701 );
    xnor g146 ( n600 , n701 , n315 );
    and g147 ( n8 , n362 , n131 );
    xnor g148 ( n78 , n836 , n19 );
    nor g149 ( n452 , n162 , n472 );
    not g150 ( n627 , n424 );
    xnor g151 ( n529 , n691 , n852 );
    and g152 ( n50 , n215 , n892 );
    not g153 ( n822 , n203 );
    nor g154 ( n628 , n41 , n427 );
    nor g155 ( n700 , n831 , n464 );
    buf g156 ( n195 , n395 );
    xnor g157 ( n12 , n131 , n652 );
    not g158 ( n845 , n460 );
    not g159 ( n214 , n849 );
    and g160 ( n386 , n332 , n423 );
    or g161 ( n896 , n832 , n126 );
    not g162 ( n753 , n356 );
    nor g163 ( n417 , n247 , n235 );
    buf g164 ( n193 , n237 );
    or g165 ( n769 , n377 , n562 );
    nor g166 ( n297 , n709 , n186 );
    buf g167 ( n200 , n844 );
    and g168 ( n751 , n877 , n294 );
    buf g169 ( n760 , n680 );
    or g170 ( n643 , n757 , n384 );
    and g171 ( n22 , n84 , n330 );
    not g172 ( n747 , n127 );
    xnor g173 ( n736 , n489 , n846 );
    or g174 ( n672 , n229 , n458 );
    or g175 ( n515 , n469 , n873 );
    nor g176 ( n629 , n639 , n498 );
    xnor g177 ( n32 , n608 , n783 );
    or g178 ( n57 , n160 , n768 );
    xnor g179 ( n130 , n621 , n854 );
    nor g180 ( n617 , n864 , n467 );
    buf g181 ( n207 , n85 );
    or g182 ( n704 , n782 , n261 );
    xnor g183 ( n328 , n262 , n145 );
    or g184 ( n170 , n777 , n118 );
    not g185 ( n273 , n737 );
    and g186 ( n390 , n897 , n31 );
    or g187 ( n882 , n343 , n347 );
    not g188 ( n88 , n732 );
    xnor g189 ( n228 , n806 , n736 );
    xnor g190 ( n877 , n19 , n713 );
    or g191 ( n472 , n368 , n42 );
    nor g192 ( n860 , n591 , n296 );
    buf g193 ( n580 , n153 );
    or g194 ( n577 , n868 , n123 );
    or g195 ( n153 , n352 , n576 );
    or g196 ( n849 , n460 , n882 );
    and g197 ( n734 , n425 , n99 );
    buf g198 ( n134 , n890 );
    or g199 ( n466 , n350 , n298 );
    or g200 ( n279 , n275 , n535 );
    or g201 ( n128 , n142 , n173 );
    or g202 ( n534 , n184 , n405 );
    and g203 ( n54 , n165 , n745 );
    nor g204 ( n118 , n44 , n738 );
    not g205 ( n67 , n64 );
    xnor g206 ( n369 , n380 , n514 );
    or g207 ( n5 , n896 , n849 );
    nor g208 ( n842 , n528 , n683 );
    buf g209 ( n109 , n729 );
    not g210 ( n743 , n386 );
    nor g211 ( n508 , n817 , n266 );
    not g212 ( n520 , n543 );
    and g213 ( n413 , n869 , n540 );
    or g214 ( n675 , n436 , n366 );
    nor g215 ( n872 , n887 , n235 );
    nor g216 ( n838 , n771 , n541 );
    and g217 ( n837 , n135 , n468 );
    not g218 ( n885 , n672 );
    nor g219 ( n412 , n295 , n663 );
    or g220 ( n175 , n177 , n719 );
    or g221 ( n793 , n221 , n98 );
    not g222 ( n494 , n269 );
    buf g223 ( n619 , n526 );
    nor g224 ( n230 , n791 , n538 );
    or g225 ( n141 , n421 , n117 );
    xnor g226 ( n89 , n489 , n600 );
    xnor g227 ( n249 , n438 , n525 );
    not g228 ( n820 , n801 );
    nor g229 ( n809 , n678 , n515 );
    xnor g230 ( n87 , n390 , n382 );
    nor g231 ( n485 , n203 , n704 );
    nor g232 ( n323 , n129 , n510 );
    nor g233 ( n152 , n286 , n372 );
    or g234 ( n648 , n870 , n831 );
    buf g235 ( n481 , n786 );
    buf g236 ( n678 , n586 );
    and g237 ( n847 , n84 , n404 );
    nor g238 ( n698 , n651 , n258 );
    nor g239 ( n47 , n892 , n484 );
    buf g240 ( n416 , n409 );
    nor g241 ( n690 , n561 , n315 );
    nor g242 ( n528 , n894 , n146 );
    not g243 ( n709 , n260 );
    not g244 ( n467 , n271 );
    or g245 ( n899 , n400 , n471 );
    not g246 ( n372 , n545 );
    xnor g247 ( n620 , n166 , n404 );
    buf g248 ( n256 , n636 );
    not g249 ( n732 , n743 );
    nor g250 ( n148 , n613 , n820 );
    buf g251 ( n281 , n454 );
    buf g252 ( n94 , n290 );
    nor g253 ( n670 , n789 , n902 );
    nor g254 ( n400 , n498 , n638 );
    buf g255 ( n84 , n39 );
    buf g256 ( n239 , n461 );
    nor g257 ( n609 , n326 , n753 );
    xnor g258 ( n546 , n605 , n78 );
    and g259 ( n686 , n671 , n211 );
    not g260 ( n765 , n621 );
    nor g261 ( n31 , n617 , n376 );
    or g262 ( n307 , n797 , n162 );
    nor g263 ( n221 , n387 , n180 );
    or g264 ( n706 , n557 , n723 );
    nor g265 ( n243 , n96 , n802 );
    or g266 ( n334 , n335 , n734 );
    not g267 ( n506 , n18 );
    and g268 ( n574 , n666 , n512 );
    nor g269 ( n264 , n659 , n75 );
    buf g270 ( n102 , n812 );
    not g271 ( n45 , n722 );
    buf g272 ( n726 , n248 );
    buf g273 ( n815 , n595 );
    xnor g274 ( n68 , n854 , n632 );
    or g275 ( n261 , n860 , n609 );
    buf g276 ( n839 , n459 );
    or g277 ( n584 , n58 , n485 );
    not g278 ( n441 , n35 );
    not g279 ( n66 , n581 );
    nor g280 ( n624 , n145 , n353 );
    and g281 ( n320 , n453 , n578 );
    not g282 ( n583 , n250 );
    xnor g283 ( n514 , n611 , n794 );
    nor g284 ( n496 , n93 , n90 );
    nor g285 ( n289 , n758 , n878 );
    xnor g286 ( n655 , n311 , n704 );
    or g287 ( n37 , n508 , n698 );
    not g288 ( n419 , n672 );
    not g289 ( n356 , n902 );
    or g290 ( n531 , n796 , n214 );
    not g291 ( n62 , n100 );
    or g292 ( n458 , n148 , n539 );
    not g293 ( n575 , n225 );
    xnor g294 ( n846 , n854 , n87 );
    not g295 ( n402 , n250 );
    not g296 ( n258 , n583 );
    nor g297 ( n691 , n700 , n792 );
    nor g298 ( n568 , n144 , n62 );
    xnor g299 ( n883 , n584 , n404 );
    nor g300 ( n656 , n428 , n869 );
    not g301 ( n257 , n5 );
    or g302 ( n763 , n185 , n292 );
    buf g303 ( n565 , n20 );
    and g304 ( n602 , n702 , n652 );
    not g305 ( n25 , n166 );
    nor g306 ( n302 , n40 , n467 );
    not g307 ( n468 , n318 );
    buf g308 ( n718 , n403 );
    or g309 ( n385 , n223 , n216 );
    nor g310 ( n792 , n892 , n885 );
    buf g311 ( n499 , n826 );
    or g312 ( n604 , n253 , n804 );
    nor g313 ( n65 , n291 , n146 );
    not g314 ( n874 , n543 );
    buf g315 ( n346 , n1 );
    or g316 ( n311 , n793 , n338 );
    not g317 ( n379 , n66 );
    not g318 ( n800 , n397 );
    not g319 ( n601 , n901 );
    buf g320 ( n536 , n147 );
    not g321 ( n711 , n127 );
    not g322 ( n599 , n163 );
    buf g323 ( n217 , n29 );
    buf g324 ( n511 , n767 );
    not g325 ( n287 , n643 );
    buf g326 ( n336 , n123 );
    not g327 ( n708 , n871 );
    not g328 ( n424 , n99 );
    not g329 ( n146 , n203 );
    not g330 ( n681 , n408 );
    or g331 ( n755 , n4 , n903 );
    buf g332 ( n161 , n707 );
    not g333 ( n61 , n166 );
    or g334 ( n205 , n676 , n194 );
    or g335 ( n354 , n838 , n670 );
    buf g336 ( n570 , n807 );
    buf g337 ( n479 , n156 );
    xnor g338 ( n752 , n212 , n775 );
    xor g339 ( n603 , n112 , n331 );
    not g340 ( n250 , n712 );
    buf g341 ( n590 , n594 );
    not g342 ( n524 , n478 );
    not g343 ( n90 , n381 );
    and g344 ( n100 , n317 , n821 );
    not g345 ( n397 , n390 );
    nor g346 ( n717 , n171 , n301 );
    not g347 ( n859 , n373 );
    and g348 ( n99 , n628 , n703 );
    buf g349 ( n196 , n393 );
    buf g350 ( n662 , n507 );
    not g351 ( n439 , n382 );
    nor g352 ( n891 , n429 , n66 );
    and g353 ( n46 , n36 , n143 );
    not g354 ( n30 , n13 );
    not g355 ( n638 , n159 );
    and g356 ( n159 , n49 , n754 );
    nor g357 ( n300 , n330 , n803 );
    not g358 ( n582 , n892 );
    not g359 ( n738 , n712 );
    not g360 ( n105 , n69 );
    and g361 ( n135 , n136 , n476 );
    buf g362 ( n893 , n304 );
    and g363 ( n73 , n692 , n80 );
    nor g364 ( n723 , n626 , n579 );
    or g365 ( n858 , n810 , n15 );
    not g366 ( n579 , n391 );
    not g367 ( n650 , n684 );
    or g368 ( n184 , n523 , n169 );
    nor g369 ( n550 , n203 , n19 );
    buf g370 ( n120 , n154 );
    and g371 ( n253 , n73 , n676 );
    or g372 ( n782 , n322 , n814 );
    nor g373 ( n0 , n875 , n244 );
    or g374 ( n478 , n596 , n297 );
    xnor g375 ( n715 , n714 , n752 );
    nor g376 ( n218 , n828 , n703 );
    not g377 ( n423 , n317 );
    and g378 ( n51 , n848 , n473 );
    buf g379 ( n705 , n688 );
    buf g380 ( n772 , n371 );
    buf g381 ( n108 , n900 );
    and g382 ( n901 , n332 , n317 );
    and g383 ( n674 , n837 , n61 );
    or g384 ( n91 , n652 , n635 );
    nor g385 ( n504 , n399 , n547 );
    or g386 ( n384 , n490 , n190 );
    or g387 ( n186 , n493 , n46 );
    xnor g388 ( n285 , n348 , n660 );
    buf g389 ( n6 , n140 );
    not g390 ( n469 , n808 );
    buf g391 ( n329 , n224 );
    and g392 ( n36 , n710 , n45 );
    xnor g393 ( n112 , n225 , n840 );
    xnor g394 ( n863 , n476 , n57 );
    xnor g395 ( n880 , n863 , n495 );
    nor g396 ( n455 , n449 , n90 );
    buf g397 ( n853 , n542 );
    nor g398 ( n523 , n867 , n392 );
    not g399 ( n235 , n712 );
    nor g400 ( n694 , n463 , n97 );
    not g401 ( n277 , n571 );
    not g402 ( n902 , n543 );
    not g403 ( n545 , n310 );
    nor g404 ( n389 , n682 , n24 );
    or g405 ( n725 , n172 , n527 );
    or g406 ( n450 , n616 , n668 );
    or g407 ( n719 , n197 , n124 );
    not g408 ( n634 , n54 );
    and g409 ( n548 , n277 , n189 );
    or g410 ( n445 , n23 , n303 );
    nor g411 ( n733 , n776 , n781 );
    xnor g412 ( n201 , n633 , n179 );
    not g413 ( n104 , n494 );
    not g414 ( n303 , n361 );
    buf g415 ( n254 , n440 );
    and g416 ( n309 , n279 , n320 );
    or g417 ( n77 , n325 , n337 );
    xnor g418 ( n17 , n201 , n249 );
    not g419 ( n318 , n311 );
    and g420 ( n366 , n119 , n553 );
    nor g421 ( n646 , n25 , n7 );
    nor g422 ( n576 , n639 , n621 );
    not g423 ( n831 , n892 );
    not g424 ( n392 , n110 );
    not g425 ( n24 , n386 );
    or g426 ( n292 , n480 , n149 );
    and g427 ( n559 , n30 , n840 );
    not g428 ( n155 , n583 );
    or g429 ( n95 , n799 , n518 );
    not g430 ( n428 , n397 );
    nor g431 ( n181 , n299 , n180 );
    and g432 ( n232 , n800 , n639 );
    or g433 ( n804 , n312 , n721 );
    and g434 ( n712 , n569 , n209 );
    and g435 ( n49 , n524 , n205 );
    not g436 ( n475 , n770 );
    or g437 ( n823 , n64 , n491 );
    xnor g438 ( n489 , n644 , n419 );
    buf g439 ( n92 , 1'b1 );
    nor g440 ( n518 , n892 , n572 );
    buf g441 ( n851 , n488 );
    nor g442 ( n825 , n411 , n582 );
    nor g443 ( n430 , n263 , n370 );
    nor g444 ( n226 , n306 , n301 );
    not g445 ( n422 , n209 );
    and g446 ( n119 , n630 , n648 );
    or g447 ( n502 , n629 , n63 );
    not g448 ( n538 , n737 );
    or g449 ( n671 , n240 , n324 );
    not g450 ( n13 , n408 );
    nor g451 ( n198 , n65 , n487 );
    not g452 ( n497 , n391 );
    or g453 ( n621 , n599 , n678 );
    nor g454 ( n756 , n115 , n128 );
    and g455 ( n779 , n283 , n107 );
    nor g456 ( n762 , n892 , n805 );
    not g457 ( n21 , n598 );
    nor g458 ( n169 , n139 , n121 );
    not g459 ( n541 , n105 );
    not g460 ( n28 , n135 );
    nor g461 ( n557 , n178 , n97 );
    or g462 ( n55 , n575 , n84 );
    not g463 ( n391 , n520 );
    nor g464 ( n98 , n780 , n364 );
    or g465 ( n315 , n466 , n37 );
    xnor g466 ( n886 , n450 , n652 );
    or g467 ( n589 , n10 , n548 );
    or g468 ( n194 , n722 , n80 );
    and g469 ( n361 , n899 , n532 );
    not g470 ( n808 , n858 );
    buf g471 ( n219 , n456 );
    nor g472 ( n172 , n413 , n434 );
    not g473 ( n878 , n49 );
    not g474 ( n127 , n236 );
    not g475 ( n758 , n779 );
    or g476 ( n869 , n847 , n505 );
    not g477 ( n280 , n122 );
    nor g478 ( n305 , n455 , n243 );
    and g479 ( n432 , n574 , n696 );
    or g480 ( n810 , n302 , n551 );
    not g481 ( n180 , n255 );
    not g482 ( n710 , n13 );
    nor g483 ( n418 , n14 , n62 );
    or g484 ( n15 , n259 , n872 );
    xnor g485 ( n436 , n558 , n840 );
    nor g486 ( n721 , n656 , n725 );
    not g487 ( n676 , n747 );
    or g488 ( n586 , n319 , n881 );
    nor g489 ( n521 , n728 , n280 );
    or g490 ( n316 , n91 , n28 );
    or g491 ( n236 , n566 , n170 );
    xnor g492 ( n34 , n365 , n731 );
    not g493 ( n151 , n296 );
    not g494 ( n730 , n390 );
    buf g495 ( n82 , n813 );
    buf g496 ( n233 , n477 );
    buf g497 ( n125 , n103 );
    nor g498 ( n641 , n451 , n865 );
    and g499 ( n58 , n38 , n203 );
    buf g500 ( n615 , n486 );
    nor g501 ( n327 , n500 , n503 );
    xor g502 ( n267 , n635 , n643 );
    or g503 ( n80 , n22 , n785 );
    not g504 ( n165 , n162 );
    or g505 ( n19 , n563 , n501 );
    buf g506 ( n462 , n182 );
    not g507 ( n703 , n402 );
    buf g508 ( n245 , n27 );
    nor g509 ( n614 , n833 , n740 );
    or g510 ( n757 , n181 , n431 );
    xnor g511 ( n843 , n293 , n687 );
    and g512 ( n532 , n51 , n316 );
    not g513 ( n513 , n852 );
    xnor g514 ( n854 , n469 , n678 );
    nor g515 ( n53 , n639 , n228 );
    buf g516 ( n344 , n345 );
    or g517 ( n562 , n106 , n763 );
    nor g518 ( n339 , n164 , n497 );
    nor g519 ( n107 , n496 , n891 );
    buf g520 ( n363 , n103 );
    nor g521 ( n693 , n892 , n104 );
    nor g522 ( n16 , n598 , n858 );
    or g523 ( n293 , n50 , n618 );
    and g524 ( n487 , n468 , n146 );
    not g525 ( n517 , n432 );
    and g526 ( n701 , n695 , n305 );
    not g527 ( n567 , n901 );
    nor g528 ( n539 , n516 , n738 );
    nor g529 ( n406 , n796 , n634 );
    and g530 ( n335 , n419 , n852 );
    and g531 ( n425 , n708 , n687 );
    xnor g532 ( n421 , n575 , n733 );
    not g533 ( n121 , n581 );
    or g534 ( n862 , n816 , n0 );
    or g535 ( n197 , n811 , n550 );
    not g536 ( n76 , n832 );
    not g537 ( n764 , n56 );
    and g538 ( n618 , n627 , n582 );
    not g539 ( n7 , n681 );
    nor g540 ( n558 , n825 , n693 );
    and g541 ( n785 , n30 , n759 );
    not g542 ( n408 , n39 );
    or g543 ( n768 , n418 , n83 );
    or g544 ( n276 , n175 , n884 );
    nor g545 ( n720 , n787 , n396 );
    nor g546 ( n724 , n653 , n649 );
    buf g547 ( n150 , n855 );
    xnor g548 ( n325 , n442 , n143 );
    nor g549 ( n415 , n189 , n827 );
    and g550 ( n596 , n36 , n231 );
    not g551 ( n381 , n396 );
    nor g552 ( n270 , n9 , n422 );
    or g553 ( n744 , n457 , n414 );
    nor g554 ( n241 , n132 , n601 );
    not g555 ( n220 , n173 );
    not g556 ( n606 , n203 );
    nor g557 ( n607 , n353 , n722 );
    buf g558 ( n637 , n251 );
    or g559 ( n473 , n731 , n549 );
    buf g560 ( n640 , n888 );
    not g561 ( n240 , n494 );
    or g562 ( n355 , n697 , n7 );
    not g563 ( n268 , n571 );
    buf g564 ( n234 , n766 );
    nor g565 ( n740 , n203 , n764 );
    buf g566 ( n898 , n552 );
    or g567 ( n56 , n168 , n706 );
    not g568 ( n484 , n747 );
    xnor g569 ( n480 , n589 , n131 );
    nor g570 ( n70 , n114 , n84 );
    not g571 ( n364 , n321 );
    and g572 ( n543 , n423 , n821 );
    and g573 ( n873 , n355 , n55 );
    and g574 ( n373 , n246 , n641 );
    or g575 ( n262 , n677 , n741 );
    nor g576 ( n593 , n778 , n634 );
    or g577 ( n338 , n52 , n685 );
    or g578 ( n881 , n327 , n218 );
    xnor g579 ( n664 , n351 , n759 );
    nor g580 ( n83 , n587 , n874 );
    and g581 ( n260 , n534 , n45 );
    or g582 ( n347 , n18 , n770 );
    nor g583 ( n695 , n669 , n819 );
    or g584 ( n211 , n646 , n559 );
    buf g585 ( n773 , n59 );
    nor g586 ( n483 , n242 , n88 );
    not g587 ( n310 , n581 );
    nor g588 ( n749 , n658 , n582 );
    or g589 ( n272 , n268 , n650 );
    not g590 ( n663 , n545 );
    nor g591 ( n818 , n643 , n674 );
    not g592 ( n396 , n271 );
    xnor g593 ( n879 , n25 , n198 );
    nor g594 ( n669 , n3 , n503 );
    xnor g595 ( n775 , n687 , n852 );
    not g596 ( n199 , n128 );
    or g597 ( n803 , n794 , n79 );
    xnor g598 ( n222 , n95 , n114 );
    not g599 ( n75 , n321 );
    nor g600 ( n167 , n631 , n654 );
    nor g601 ( n259 , n86 , n857 );
    not g602 ( n805 , n439 );
    not g603 ( n227 , n386 );
    not g604 ( n173 , n57 );
    or g605 ( n43 , n694 , n339 );
    not g606 ( n848 , n674 );
    not g607 ( n644 , n424 );
    not g608 ( n255 , n227 );
    xnor g609 ( n495 , n655 , n267 );
    buf g610 ( n282 , n123 );
    nor g611 ( n350 , n202 , n547 );
    not g612 ( n561 , n639 );
    not g613 ( n547 , n110 );
    or g614 ( n512 , n4 , n308 );
    xor g615 ( n453 , n333 , n715 );
    and g616 ( n811 , n623 , n203 );
    not g617 ( n35 , n273 );
    not g618 ( n332 , n821 );
    buf g619 ( n470 , n123 );
    xnor g620 ( n889 , n87 , n68 );
    nor g621 ( n612 , n137 , n258 );
    xnor g622 ( n714 , n759 , n143 );
    buf g623 ( n509 , n798 );
    buf g624 ( n116 , n192 );
    not g625 ( n635 , n859 );
    nor g626 ( n298 , n210 , n372 );
    nor g627 ( n865 , n784 , n753 );
    nor g628 ( n447 , n834 , n820 );
    nor g629 ( n653 , n822 , n622 );
    or g630 ( n149 , n529 , n886 );
    nor g631 ( n490 , n183 , n830 );
    buf g632 ( n113 , n358 );
    not g633 ( n266 , n801 );
    nor g634 ( n610 , n554 , n538 );
    not g635 ( n191 , n374 );
    or g636 ( n433 , n21 , n765 );
    nor g637 ( n283 , n447 , n612 );
    and g638 ( n216 , n445 , n588 );
    not g639 ( n684 , n28 );
    or g640 ( n33 , n21 , n130 );
    buf g641 ( n750 , n133 );
    not g642 ( n189 , n892 );
    nor g643 ( n816 , n482 , n24 );
    not g644 ( n801 , n273 );
    nor g645 ( n23 , n131 , n272 );
    not g646 ( n69 , n100 );
    buf g647 ( n647 , n60 );
    nor g648 ( n692 , n478 , n722 );
    nor g649 ( n833 , n606 , n661 );
    nor g650 ( n322 , n625 , n743 );
    buf g651 ( n349 , n206 );
    nor g652 ( n777 , n585 , n441 );
    nor g653 ( n427 , n856 , n857 );
    or g654 ( n41 , n430 , n270 );
    or g655 ( n563 , n389 , n208 );
    xnor g656 ( n742 , n294 , n713 );
    buf g657 ( n560 , n555 );
    or g658 ( n566 , n720 , n412 );
    not g659 ( n324 , n515 );
    or g660 ( n501 , n568 , n341 );
    and g661 ( n616 , n522 , n203 );
    nor g662 ( n685 , n448 , n874 );
    nor g663 ( n451 , n72 , n830 );
    not g664 ( n244 , n901 );
    and g665 ( n737 , n422 , n263 );
    nor g666 ( n190 , n378 , n497 );
    or g667 ( n117 , n519 , n675 );
    not g668 ( n498 , n191 );
    not g669 ( n510 , n402 );
    not g670 ( n745 , n774 );
endmodule
