module top( n3 , n8 , n26 , n40 , n41 , n44 , n46 , n54 , n67 , 
n71 , n81 , n93 , n97 , n103 , n109 , n121 , n123 , n130 , n132 , 
n134 , n146 , n153 , n154 , n161 , n167 , n168 , n169 , n173 , n176 , 
n177 , n178 , n183 , n186 , n187 , n197 , n198 , n201 , n208 , n217 , 
n219 , n221 , n229 , n235 , n236 , n246 , n248 , n256 , n260 , n261 , 
n275 , n278 , n280 , n298 , n301 , n311 , n317 , n325 , n328 , n333 , 
n336 , n345 , n349 , n361 , n362 , n368 , n386 , n388 , n395 , n400 , 
n404 , n405 , n419 , n426 , n430 , n432 , n433 , n441 , n455 , n462 , 
n466 , n467 , n474 , n479 , n502 , n505 , n506 , n511 , n519 , n521 , 
n523 , n525 , n531 , n542 , n546 , n557 , n558 , n560 , n561 , n571 , 
n574 , n577 , n578 , n582 , n584 , n585 , n600 , n607 , n608 , n615 , 
n620 , n627 , n629 , n631 , n649 , n652 , n664 , n667 , n678 , n683 , 
n685 , n688 , n694 , n698 , n711 , n712 , n732 , n751 , n753 , n757 , 
n758 , n773 , n778 , n780 , n804 , n809 , n820 , n823 , n827 , n829 , 
n836 , n837 , n838 , n840 , n841 , n848 , n850 , n866 , n873 , n878 , 
n879 , n888 , n892 , n903 , n904 , n909 , n910 , n915 , n917 , n927 , 
n930 , n931 , n932 , n940 , n947 , n957 , n958 , n964 , n966 , n981 , 
n985 , n990 , n994 , n995 , n1002 , n1004 , n1015 , n1025 , n1043 , n1045 , 
n1049 , n1051 , n1067 , n1068 , n1071 , n1074 , n1075 , n1090 , n1099 , n1108 , 
n1118 , n1132 , n1138 , n1139 , n1141 , n1165 , n1170 , n1172 , n1177 , n1187 , 
n1200 , n1211 , n1217 , n1220 , n1222 , n1232 , n1239 , n1250 , n1254 , n1256 , 
n1259 , n1268 , n1272 , n1276 , n1281 , n1284 , n1285 , n1298 , n1305 , n1306 , 
n1307 , n1310 , n1314 , n1315 , n1320 , n1322 , n1324 , n1351 , n1366 , n1371 , 
n1376 , n1378 , n1382 , n1392 , n1393 , n1394 , n1395 , n1397 , n1399 , n1409 , 
n1420 , n1427 , n1432 , n1433 , n1448 , n1449 , n1451 , n1454 , n1467 , n1471 , 
n1474 , n1483 , n1490 , n1495 , n1504 , n1524 , n1529 , n1534 , n1543 , n1549 , 
n1550 , n1559 , n1565 , n1574 , n1575 , n1578 , n1580 , n1582 , n1584 , n1589 , 
n1596 , n1601 , n1605 , n1615 , n1622 , n1623 , n1624 , n1627 , n1629 , n1631 , 
n1633 , n1640 , n1645 , n1654 , n1669 , n1679 , n1680 , n1682 , n1686 , n1690 , 
n1691 , n1692 , n1700 , n1701 , n1702 , n1708 , n1718 , n1720 , n1726 , n1731 , 
n1736 , n1738 , n1751 , n1764 , n1775 , n1785 , n1787 , n1800 , n1804 , n1805 , 
n1806 , n1815 , n1817 , n1819 , n1822 , n1834 , n1842 , n1855 , n1863 , n1867 , 
n1873 , n1877 , n1884 , n1903 , n1904 , n1916 , n1920 , n1926 , n1936 , n1938 , 
n1941 , n1945 , n1947 , n1950 , n1962 , n1965 , n1975 , n1982 , n1999 , n2002 , 
n2004 , n2014 , n2017 , n2021 , n2027 , n2033 , n2034 , n2040 , n2043 , n2052 , 
n2065 , n2068 , n2076 , n2079 , n2087 , n2090 , n2095 , n2096 , n2097 , n2112 , 
n2118 , n2119 , n2121 , n2124 , n2140 , n2146 , n2151 , n2183 , n2185 , n2187 , 
n2188 , n2206 , n2216 , n2236 , n2242 , n2253 , n2255 , n2263 , n2273 , n2283 , 
n2286 , n2289 , n2293 , n2296 , n2297 , n2303 , n2307 , n2311 , n2312 , n2321 , 
n2325 , n2328 , n2330 , n2339 , n2344 , n2360 , n2378 , n2390 , n2393 , n2394 , 
n2397 , n2398 , n2405 , n2407 , n2417 , n2422 , n2431 , n2433 , n2437 , n2439 , 
n2440 , n2444 , n2445 , n2449 , n2474 , n2478 , n2484 , n2488 , n2493 , n2501 , 
n2502 , n2507 , n2520 , n2521 , n2543 , n2544 , n2547 , n2550 , n2553 , n2559 , 
n2572 , n2577 , n2578 , n2590 , n2609 , n2611 , n2621 , n2635 , n2636 , n2644 , 
n2647 , n2649 , n2651 , n2661 , n2662 , n2668 , n2671 , n2676 , n2693 , n2694 , 
n2705 , n2707 , n2711 , n2712 , n2721 , n2726 , n2731 , n2732 , n2734 , n2736 , 
n2745 , n2751 , n2752 , n2758 , n2761 , n2767 , n2773 , n2775 , n2787 , n2788 , 
n2800 , n2806 , n2812 , n2833 , n2843 , n2853 , n2855 , n2862 , n2865 , n2880 , 
n2883 , n2889 , n2890 , n2893 , n2895 , n2896 , n2912 , n2915 , n2928 , n2929 , 
n2932 , n2950 , n2954 , n2962 , n2971 , n2974 , n2975 , n2979 , n2990 , n2991 , 
n3001 , n3007 , n3013 , n3017 , n3021 , n3024 , n3025 , n3026 , n3035 , n3039 , 
n3044 , n3045 , n3050 , n3052 , n3054 , n3060 , n3068 , n3083 , n3092 , n3106 , 
n3114 , n3125 , n3133 , n3143 , n3145 , n3154 , n3156 , n3157 , n3158 , n3168 , 
n3186 , n3188 , n3199 , n3203 , n3206 , n3210 , n3214 , n3218 , n3245 , n3247 , 
n3248 , n3250 , n3266 , n3269 , n3278 , n3287 , n3288 , n3291 , n3299 , n3308 , 
n3314 , n3318 , n3323 , n3325 , n3327 , n3330 , n3335 , n3336 , n3359 , n3367 , 
n3373 , n3377 , n3381 , n3385 , n3387 , n3401 , n3415 , n3417 , n3418 , n3432 , 
n3436 , n3475 , n3487 , n3498 , n3502 , n3504 , n3511 , n3522 , n3525 , n3532 , 
n3539 , n3541 , n3543 , n3544 , n3552 , n3570 , n3573 , n3576 , n3582 , n3585 , 
n3586 , n3590 , n3607 , n3617 , n3626 , n3637 , n3639 , n3641 , n3642 , n3645 , 
n3646 , n3656 , n3672 , n3673 , n3676 , n3682 , n3684 , n3693 , n3696 , n3697 , 
n3698 , n3700 , n3702 , n3712 , n3714 , n3718 , n3721 , n3725 , n3732 , n3754 , 
n3755 , n3756 , n3758 , n3762 , n3776 , n3778 , n3784 , n3785 , n3786 , n3801 , 
n3807 , n3808 , n3809 , n3814 , n3819 , n3820 , n3822 , n3826 , n3827 , n3837 , 
n3843 , n3848 , n3854 );
    input n3 , n26 , n40 , n44 , n46 , n54 , n81 , n93 , n97 , 
n103 , n109 , n121 , n123 , n130 , n132 , n134 , n146 , n161 , n167 , 
n169 , n173 , n176 , n177 , n178 , n183 , n186 , n187 , n197 , n198 , 
n208 , n217 , n221 , n229 , n235 , n236 , n246 , n248 , n256 , n260 , 
n261 , n275 , n278 , n298 , n301 , n311 , n317 , n328 , n333 , n336 , 
n345 , n349 , n361 , n362 , n368 , n386 , n388 , n395 , n400 , n404 , 
n405 , n430 , n432 , n433 , n441 , n455 , n462 , n466 , n467 , n474 , 
n479 , n502 , n506 , n511 , n519 , n521 , n523 , n525 , n531 , n542 , 
n546 , n557 , n558 , n560 , n561 , n571 , n574 , n577 , n578 , n582 , 
n584 , n585 , n607 , n608 , n615 , n620 , n627 , n631 , n649 , n652 , 
n667 , n678 , n683 , n685 , n688 , n694 , n698 , n711 , n712 , n732 , 
n751 , n753 , n773 , n780 , n804 , n809 , n820 , n827 , n836 , n837 , 
n838 , n841 , n848 , n850 , n866 , n873 , n878 , n903 , n904 , n927 , 
n930 , n931 , n932 , n947 , n958 , n964 , n966 , n981 , n990 , n994 , 
n995 , n1002 , n1015 , n1043 , n1045 , n1049 , n1051 , n1068 , n1071 , n1074 , 
n1075 , n1099 , n1108 , n1118 , n1132 , n1139 , n1141 , n1170 , n1172 , n1187 , 
n1200 , n1211 , n1217 , n1220 , n1222 , n1232 , n1250 , n1254 , n1259 , n1268 , 
n1276 , n1281 , n1285 , n1298 , n1305 , n1314 , n1315 , n1322 , n1324 , n1351 , 
n1371 , n1376 , n1382 , n1392 , n1393 , n1395 , n1397 , n1420 , n1427 , n1433 , 
n1448 , n1449 , n1451 , n1454 , n1467 , n1471 , n1474 , n1483 , n1490 , n1495 , 
n1504 , n1524 , n1529 , n1534 , n1549 , n1550 , n1559 , n1574 , n1575 , n1578 , 
n1580 , n1582 , n1584 , n1589 , n1596 , n1601 , n1605 , n1615 , n1622 , n1623 , 
n1624 , n1627 , n1631 , n1640 , n1645 , n1654 , n1669 , n1680 , n1682 , n1686 , 
n1691 , n1692 , n1700 , n1701 , n1702 , n1708 , n1720 , n1726 , n1731 , n1736 , 
n1738 , n1764 , n1775 , n1785 , n1787 , n1800 , n1804 , n1805 , n1806 , n1817 , 
n1819 , n1822 , n1834 , n1842 , n1855 , n1873 , n1877 , n1884 , n1904 , n1916 , 
n1926 , n1938 , n1941 , n1947 , n1950 , n1962 , n1965 , n1975 , n1982 , n1999 , 
n2002 , n2004 , n2014 , n2017 , n2027 , n2034 , n2043 , n2052 , n2068 , n2076 , 
n2079 , n2090 , n2096 , n2097 , n2112 , n2118 , n2121 , n2124 , n2140 , n2146 , 
n2151 , n2183 , n2185 , n2187 , n2188 , n2216 , n2236 , n2242 , n2253 , n2255 , 
n2263 , n2283 , n2289 , n2296 , n2297 , n2303 , n2311 , n2312 , n2321 , n2325 , 
n2328 , n2330 , n2339 , n2378 , n2390 , n2393 , n2397 , n2405 , n2407 , n2417 , 
n2422 , n2431 , n2433 , n2437 , n2439 , n2444 , n2445 , n2449 , n2474 , n2478 , 
n2484 , n2488 , n2493 , n2507 , n2520 , n2521 , n2543 , n2544 , n2547 , n2550 , 
n2553 , n2559 , n2572 , n2577 , n2578 , n2590 , n2609 , n2611 , n2635 , n2636 , 
n2644 , n2647 , n2649 , n2651 , n2661 , n2662 , n2668 , n2671 , n2676 , n2693 , 
n2705 , n2711 , n2712 , n2721 , n2726 , n2731 , n2732 , n2736 , n2745 , n2752 , 
n2758 , n2761 , n2767 , n2773 , n2775 , n2787 , n2806 , n2812 , n2843 , n2853 , 
n2855 , n2862 , n2865 , n2883 , n2889 , n2890 , n2893 , n2896 , n2915 , n2928 , 
n2929 , n2932 , n2950 , n2962 , n2971 , n2975 , n2990 , n3001 , n3007 , n3013 , 
n3021 , n3024 , n3025 , n3026 , n3035 , n3044 , n3050 , n3052 , n3054 , n3060 , 
n3092 , n3106 , n3114 , n3125 , n3133 , n3143 , n3145 , n3154 , n3156 , n3157 , 
n3168 , n3186 , n3188 , n3199 , n3203 , n3210 , n3214 , n3218 , n3245 , n3248 , 
n3250 , n3266 , n3269 , n3278 , n3287 , n3288 , n3291 , n3299 , n3308 , n3314 , 
n3318 , n3323 , n3325 , n3335 , n3336 , n3367 , n3373 , n3377 , n3381 , n3385 , 
n3401 , n3415 , n3417 , n3418 , n3432 , n3436 , n3475 , n3487 , n3498 , n3502 , 
n3504 , n3522 , n3525 , n3539 , n3541 , n3544 , n3552 , n3570 , n3573 , n3576 , 
n3582 , n3585 , n3586 , n3590 , n3607 , n3626 , n3637 , n3639 , n3641 , n3646 , 
n3656 , n3672 , n3673 , n3682 , n3684 , n3693 , n3697 , n3698 , n3700 , n3702 , 
n3718 , n3721 , n3725 , n3732 , n3754 , n3755 , n3756 , n3758 , n3776 , n3784 , 
n3785 , n3786 , n3801 , n3807 , n3808 , n3819 , n3820 , n3822 , n3826 , n3827 , 
n3843 , n3848 , n3854 ;
    output n8 , n41 , n67 , n71 , n153 , n154 , n168 , n201 , n219 , 
n280 , n325 , n419 , n426 , n505 , n600 , n629 , n664 , n757 , n758 , 
n778 , n823 , n829 , n840 , n879 , n888 , n892 , n909 , n910 , n915 , 
n917 , n940 , n957 , n985 , n1004 , n1025 , n1067 , n1090 , n1138 , n1165 , 
n1177 , n1239 , n1256 , n1272 , n1284 , n1306 , n1307 , n1310 , n1320 , n1366 , 
n1378 , n1394 , n1399 , n1409 , n1432 , n1543 , n1565 , n1629 , n1633 , n1679 , 
n1690 , n1718 , n1751 , n1815 , n1863 , n1867 , n1903 , n1920 , n1936 , n1945 , 
n2021 , n2033 , n2040 , n2065 , n2087 , n2095 , n2119 , n2206 , n2273 , n2286 , 
n2293 , n2307 , n2344 , n2360 , n2394 , n2398 , n2440 , n2501 , n2502 , n2621 , 
n2694 , n2707 , n2734 , n2751 , n2788 , n2800 , n2833 , n2880 , n2895 , n2912 , 
n2954 , n2974 , n2979 , n2991 , n3017 , n3039 , n3045 , n3068 , n3083 , n3158 , 
n3206 , n3247 , n3327 , n3330 , n3359 , n3387 , n3511 , n3532 , n3543 , n3617 , 
n3642 , n3645 , n3676 , n3696 , n3712 , n3714 , n3762 , n3778 , n3809 , n3814 , 
n3837 ;
    wire n0 , n1 , n2 , n4 , n5 , n6 , n7 , n9 , n10 , 
n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
n21 , n22 , n23 , n24 , n25 , n27 , n28 , n29 , n30 , n31 , 
n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n42 , n43 , 
n45 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n55 , n56 , 
n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , 
n68 , n69 , n70 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , 
n79 , n80 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
n90 , n91 , n92 , n94 , n95 , n96 , n98 , n99 , n100 , n101 , 
n102 , n104 , n105 , n106 , n107 , n108 , n110 , n111 , n112 , n113 , 
n114 , n115 , n116 , n117 , n118 , n119 , n120 , n122 , n124 , n125 , 
n126 , n127 , n128 , n129 , n131 , n133 , n135 , n136 , n137 , n138 , 
n139 , n140 , n141 , n142 , n143 , n144 , n145 , n147 , n148 , n149 , 
n150 , n151 , n152 , n155 , n156 , n157 , n158 , n159 , n160 , n162 , 
n163 , n164 , n165 , n166 , n170 , n171 , n172 , n174 , n175 , n179 , 
n180 , n181 , n182 , n184 , n185 , n188 , n189 , n190 , n191 , n192 , 
n193 , n194 , n195 , n196 , n199 , n200 , n202 , n203 , n204 , n205 , 
n206 , n207 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , 
n218 , n220 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n230 , 
n231 , n232 , n233 , n234 , n237 , n238 , n239 , n240 , n241 , n242 , 
n243 , n244 , n245 , n247 , n249 , n250 , n251 , n252 , n253 , n254 , 
n255 , n257 , n258 , n259 , n262 , n263 , n264 , n265 , n266 , n267 , 
n268 , n269 , n270 , n271 , n272 , n273 , n274 , n276 , n277 , n279 , 
n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , 
n291 , n292 , n293 , n294 , n295 , n296 , n297 , n299 , n300 , n302 , 
n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n312 , n313 , 
n314 , n315 , n316 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , 
n326 , n327 , n329 , n330 , n331 , n332 , n334 , n335 , n337 , n338 , 
n339 , n340 , n341 , n342 , n343 , n344 , n346 , n347 , n348 , n350 , 
n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , 
n363 , n364 , n365 , n366 , n367 , n369 , n370 , n371 , n372 , n373 , 
n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , 
n384 , n385 , n387 , n389 , n390 , n391 , n392 , n393 , n394 , n396 , 
n397 , n398 , n399 , n401 , n402 , n403 , n406 , n407 , n408 , n409 , 
n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n420 , 
n421 , n422 , n423 , n424 , n425 , n427 , n428 , n429 , n431 , n434 , 
n435 , n436 , n437 , n438 , n439 , n440 , n442 , n443 , n444 , n445 , 
n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n456 , 
n457 , n458 , n459 , n460 , n461 , n463 , n464 , n465 , n468 , n469 , 
n470 , n471 , n472 , n473 , n475 , n476 , n477 , n478 , n480 , n481 , 
n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , 
n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , 
n503 , n504 , n507 , n508 , n509 , n510 , n512 , n513 , n514 , n515 , 
n516 , n517 , n518 , n520 , n522 , n524 , n526 , n527 , n528 , n529 , 
n530 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , 
n541 , n543 , n544 , n545 , n547 , n548 , n549 , n550 , n551 , n552 , 
n553 , n554 , n555 , n556 , n559 , n562 , n563 , n564 , n565 , n566 , 
n567 , n568 , n569 , n570 , n572 , n573 , n575 , n576 , n579 , n580 , 
n581 , n583 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , 
n594 , n595 , n596 , n597 , n598 , n599 , n601 , n602 , n603 , n604 , 
n605 , n606 , n609 , n610 , n611 , n612 , n613 , n614 , n616 , n617 , 
n618 , n619 , n621 , n622 , n623 , n624 , n625 , n626 , n628 , n630 , 
n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , 
n642 , n643 , n644 , n645 , n646 , n647 , n648 , n650 , n651 , n653 , 
n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , 
n665 , n666 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , 
n676 , n677 , n679 , n680 , n681 , n682 , n684 , n686 , n687 , n689 , 
n690 , n691 , n692 , n693 , n695 , n696 , n697 , n699 , n700 , n701 , 
n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n713 , 
n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , 
n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n733 , n734 , 
n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , 
n745 , n746 , n747 , n748 , n749 , n750 , n752 , n754 , n755 , n756 , 
n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , 
n769 , n770 , n771 , n772 , n774 , n775 , n776 , n777 , n779 , n781 , 
n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , 
n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , 
n802 , n803 , n805 , n806 , n807 , n808 , n810 , n811 , n812 , n813 , 
n814 , n815 , n816 , n817 , n818 , n819 , n821 , n822 , n824 , n825 , 
n826 , n828 , n830 , n831 , n832 , n833 , n834 , n835 , n839 , n842 , 
n843 , n844 , n845 , n846 , n847 , n849 , n851 , n852 , n853 , n854 , 
n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , 
n865 , n867 , n868 , n869 , n870 , n871 , n872 , n874 , n875 , n876 , 
n877 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n889 , 
n890 , n891 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , 
n901 , n902 , n905 , n906 , n907 , n908 , n911 , n912 , n913 , n914 , 
n916 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , 
n928 , n929 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n941 , 
n942 , n943 , n944 , n945 , n946 , n948 , n949 , n950 , n951 , n952 , 
n953 , n954 , n955 , n956 , n959 , n960 , n961 , n962 , n963 , n965 , 
n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , 
n977 , n978 , n979 , n980 , n982 , n983 , n984 , n986 , n987 , n988 , 
n989 , n991 , n992 , n993 , n996 , n997 , n998 , n999 , n1000 , n1001 , 
n1003 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , 
n1014 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , 
n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , 
n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1044 , n1046 , n1047 , 
n1048 , n1050 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1069 , n1070 , n1072 , 
n1073 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , 
n1085 , n1086 , n1087 , n1088 , n1089 , n1091 , n1092 , n1093 , n1094 , n1095 , 
n1096 , n1097 , n1098 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , 
n1107 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , 
n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , 
n1129 , n1130 , n1131 , n1133 , n1134 , n1135 , n1136 , n1137 , n1140 , n1142 , 
n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , 
n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , 
n1163 , n1164 , n1166 , n1167 , n1168 , n1169 , n1171 , n1173 , n1174 , n1175 , 
n1176 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , 
n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , 
n1198 , n1199 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , 
n1209 , n1210 , n1212 , n1213 , n1214 , n1215 , n1216 , n1218 , n1219 , n1221 , 
n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1233 , 
n1234 , n1235 , n1236 , n1237 , n1238 , n1240 , n1241 , n1242 , n1243 , n1244 , 
n1245 , n1246 , n1247 , n1248 , n1249 , n1251 , n1252 , n1253 , n1255 , n1257 , 
n1258 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1269 , 
n1270 , n1271 , n1273 , n1274 , n1275 , n1277 , n1278 , n1279 , n1280 , n1282 , 
n1283 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , 
n1295 , n1296 , n1297 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1308 , 
n1309 , n1311 , n1312 , n1313 , n1316 , n1317 , n1318 , n1319 , n1321 , n1323 , 
n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , 
n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , 
n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1352 , n1353 , n1354 , n1355 , 
n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , 
n1367 , n1368 , n1369 , n1370 , n1372 , n1373 , n1374 , n1375 , n1377 , n1379 , 
n1380 , n1381 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , 
n1391 , n1396 , n1398 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , 
n1407 , n1408 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , 
n1418 , n1419 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1428 , n1429 , 
n1430 , n1431 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , 
n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1450 , n1452 , n1453 , n1455 , 
n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , 
n1466 , n1468 , n1469 , n1470 , n1472 , n1473 , n1475 , n1476 , n1477 , n1478 , 
n1479 , n1480 , n1481 , n1482 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
n1491 , n1492 , n1493 , n1494 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , 
n1502 , n1503 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , 
n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , 
n1523 , n1525 , n1526 , n1527 , n1528 , n1530 , n1531 , n1532 , n1533 , n1535 , 
n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1544 , n1545 , n1546 , 
n1547 , n1548 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , 
n1560 , n1561 , n1562 , n1563 , n1564 , n1566 , n1567 , n1568 , n1569 , n1570 , 
n1571 , n1572 , n1573 , n1576 , n1577 , n1579 , n1581 , n1583 , n1585 , n1586 , 
n1587 , n1588 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1597 , n1598 , 
n1599 , n1600 , n1602 , n1603 , n1604 , n1606 , n1607 , n1608 , n1609 , n1610 , 
n1611 , n1612 , n1613 , n1614 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , 
n1625 , n1626 , n1628 , n1630 , n1632 , n1634 , n1635 , n1636 , n1637 , n1638 , 
n1639 , n1641 , n1642 , n1643 , n1644 , n1646 , n1647 , n1648 , n1649 , n1650 , 
n1651 , n1652 , n1653 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , 
n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1670 , n1671 , n1672 , 
n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1681 , n1683 , n1684 , n1685 , 
n1687 , n1688 , n1689 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
n1703 , n1704 , n1705 , n1706 , n1707 , n1709 , n1710 , n1711 , n1712 , n1713 , 
n1714 , n1715 , n1716 , n1717 , n1719 , n1721 , n1722 , n1723 , n1724 , n1725 , 
n1727 , n1728 , n1729 , n1730 , n1732 , n1733 , n1734 , n1735 , n1737 , n1739 , 
n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
n1750 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , 
n1761 , n1762 , n1763 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , 
n1772 , n1773 , n1774 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , 
n1783 , n1784 , n1786 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , 
n1795 , n1796 , n1797 , n1798 , n1799 , n1801 , n1802 , n1803 , n1807 , n1808 , 
n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1816 , n1818 , n1820 , n1821 , 
n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , 
n1833 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1843 , n1844 , 
n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , 
n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1864 , n1865 , n1866 , 
n1868 , n1869 , n1870 , n1871 , n1872 , n1874 , n1875 , n1876 , n1878 , n1879 , 
n1880 , n1881 , n1882 , n1883 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , 
n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , 
n1901 , n1902 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , 
n1913 , n1914 , n1915 , n1917 , n1918 , n1919 , n1921 , n1922 , n1923 , n1924 , 
n1925 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , 
n1937 , n1939 , n1940 , n1942 , n1943 , n1944 , n1946 , n1948 , n1949 , n1951 , 
n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , 
n1963 , n1964 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , 
n1974 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1983 , n1984 , n1985 , 
n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , 
n1996 , n1997 , n1998 , n2000 , n2001 , n2003 , n2005 , n2006 , n2007 , n2008 , 
n2009 , n2010 , n2011 , n2012 , n2013 , n2015 , n2016 , n2018 , n2019 , n2020 , 
n2022 , n2023 , n2024 , n2025 , n2026 , n2028 , n2029 , n2030 , n2031 , n2032 , 
n2035 , n2036 , n2037 , n2038 , n2039 , n2041 , n2042 , n2044 , n2045 , n2046 , 
n2047 , n2048 , n2049 , n2050 , n2051 , n2053 , n2054 , n2055 , n2056 , n2057 , 
n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2066 , n2067 , n2069 , 
n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2077 , n2078 , n2080 , n2081 , 
n2082 , n2083 , n2084 , n2085 , n2086 , n2088 , n2089 , n2091 , n2092 , n2093 , 
n2094 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , 
n2107 , n2108 , n2109 , n2110 , n2111 , n2113 , n2114 , n2115 , n2116 , n2117 , 
n2120 , n2122 , n2123 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , 
n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2141 , n2142 , 
n2143 , n2144 , n2145 , n2147 , n2148 , n2149 , n2150 , n2152 , n2153 , n2154 , 
n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , 
n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , 
n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2184 , n2186 , 
n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , 
n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2207 , n2208 , n2209 , 
n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2217 , n2218 , n2219 , n2220 , 
n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , 
n2231 , n2232 , n2233 , n2234 , n2235 , n2237 , n2238 , n2239 , n2240 , n2241 , 
n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , 
n2254 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2264 , n2265 , 
n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2274 , n2275 , n2276 , 
n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2284 , n2285 , n2287 , n2288 , 
n2290 , n2291 , n2292 , n2294 , n2295 , n2298 , n2299 , n2300 , n2301 , n2302 , 
n2304 , n2305 , n2306 , n2308 , n2309 , n2310 , n2313 , n2314 , n2315 , n2316 , 
n2317 , n2318 , n2319 , n2320 , n2322 , n2323 , n2324 , n2326 , n2327 , n2329 , 
n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2340 , n2341 , 
n2342 , n2343 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , 
n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2361 , n2362 , n2363 , 
n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , 
n2374 , n2375 , n2376 , n2377 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , 
n2385 , n2386 , n2387 , n2388 , n2389 , n2391 , n2392 , n2395 , n2396 , n2399 , 
n2400 , n2401 , n2402 , n2403 , n2404 , n2406 , n2408 , n2409 , n2410 , n2411 , 
n2412 , n2413 , n2414 , n2415 , n2416 , n2418 , n2419 , n2420 , n2421 , n2423 , 
n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2432 , n2434 , n2435 , 
n2436 , n2438 , n2441 , n2442 , n2443 , n2446 , n2447 , n2448 , n2450 , n2451 , 
n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , 
n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , 
n2472 , n2473 , n2475 , n2476 , n2477 , n2479 , n2480 , n2481 , n2482 , n2483 , 
n2485 , n2486 , n2487 , n2489 , n2490 , n2491 , n2492 , n2494 , n2495 , n2496 , 
n2497 , n2498 , n2499 , n2500 , n2503 , n2504 , n2505 , n2506 , n2508 , n2509 , 
n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , 
n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , 
n2542 , n2545 , n2546 , n2548 , n2549 , n2551 , n2552 , n2554 , n2555 , n2556 , 
n2557 , n2558 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , 
n2568 , n2569 , n2570 , n2571 , n2573 , n2574 , n2575 , n2576 , n2579 , n2580 , 
n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2591 , 
n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , 
n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2610 , n2612 , n2613 , 
n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2622 , n2623 , n2624 , 
n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , 
n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2645 , n2646 , n2648 , 
n2650 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
n2663 , n2664 , n2665 , n2666 , n2667 , n2669 , n2670 , n2672 , n2673 , n2674 , 
n2675 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , 
n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2695 , n2696 , n2697 , 
n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2706 , n2708 , n2709 , 
n2710 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2722 , 
n2723 , n2724 , n2725 , n2727 , n2728 , n2729 , n2730 , n2733 , n2735 , n2737 , 
n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2746 , n2747 , n2748 , 
n2749 , n2750 , n2753 , n2754 , n2755 , n2756 , n2757 , n2759 , n2760 , n2762 , 
n2763 , n2764 , n2765 , n2766 , n2768 , n2769 , n2770 , n2771 , n2772 , n2774 , 
n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , 
n2786 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , 
n2798 , n2799 , n2801 , n2802 , n2803 , n2804 , n2805 , n2807 , n2808 , n2809 , 
n2810 , n2811 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , 
n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , 
n2831 , n2832 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , 
n2842 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , 
n2854 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2863 , n2864 , n2866 , 
n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , 
n2877 , n2878 , n2879 , n2881 , n2882 , n2884 , n2885 , n2886 , n2887 , n2888 , 
n2891 , n2892 , n2894 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , 
n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2913 , n2914 , 
n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , 
n2926 , n2927 , n2930 , n2931 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , 
n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , 
n2949 , n2951 , n2952 , n2953 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , 
n2961 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2972 , 
n2973 , n2976 , n2977 , n2978 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , 
n2986 , n2987 , n2988 , n2989 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , 
n2998 , n2999 , n3000 , n3002 , n3003 , n3004 , n3005 , n3006 , n3008 , n3009 , 
n3010 , n3011 , n3012 , n3014 , n3015 , n3016 , n3018 , n3019 , n3020 , n3022 , 
n3023 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3036 , 
n3037 , n3038 , n3040 , n3041 , n3042 , n3043 , n3046 , n3047 , n3048 , n3049 , 
n3051 , n3053 , n3055 , n3056 , n3057 , n3058 , n3059 , n3061 , n3062 , n3063 , 
n3064 , n3065 , n3066 , n3067 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , 
n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3084 , n3085 , 
n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3093 , n3094 , n3095 , n3096 , 
n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3107 , 
n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3115 , n3116 , n3117 , n3118 , 
n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3126 , n3127 , n3128 , n3129 , 
n3130 , n3131 , n3132 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
n3141 , n3142 , n3144 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , 
n3153 , n3155 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , 
n3167 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , 
n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3187 , n3189 , 
n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3200 , 
n3201 , n3202 , n3204 , n3205 , n3207 , n3208 , n3209 , n3211 , n3212 , n3213 , 
n3215 , n3216 , n3217 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , 
n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , 
n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3246 , 
n3249 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3267 , n3268 , n3270 , n3271 , 
n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3279 , n3280 , n3281 , n3282 , 
n3283 , n3284 , n3285 , n3286 , n3289 , n3290 , n3292 , n3293 , n3294 , n3295 , 
n3296 , n3297 , n3298 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , 
n3307 , n3309 , n3310 , n3311 , n3312 , n3313 , n3315 , n3316 , n3317 , n3319 , 
n3320 , n3321 , n3322 , n3324 , n3326 , n3328 , n3329 , n3331 , n3332 , n3333 , 
n3334 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , 
n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , 
n3356 , n3357 , n3358 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , 
n3368 , n3369 , n3370 , n3371 , n3372 , n3374 , n3375 , n3376 , n3378 , n3379 , 
n3380 , n3382 , n3383 , n3384 , n3386 , n3388 , n3389 , n3390 , n3391 , n3392 , 
n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3402 , n3403 , 
n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , 
n3414 , n3416 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , 
n3427 , n3428 , n3429 , n3430 , n3431 , n3433 , n3434 , n3435 , n3437 , n3438 , 
n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , 
n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , 
n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , 
n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3476 , n3477 , n3478 , n3479 , 
n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3488 , n3489 , n3490 , 
n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3499 , n3500 , n3501 , 
n3503 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3512 , n3513 , n3514 , 
n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3523 , n3524 , n3526 , 
n3527 , n3528 , n3529 , n3530 , n3531 , n3533 , n3534 , n3535 , n3536 , n3537 , 
n3538 , n3540 , n3542 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , 
n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , 
n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3571 , n3572 , n3574 , 
n3575 , n3577 , n3578 , n3579 , n3580 , n3581 , n3583 , n3584 , n3587 , n3588 , 
n3589 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3608 , n3609 , n3610 , 
n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3618 , n3619 , n3620 , n3621 , 
n3622 , n3623 , n3624 , n3625 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , 
n3633 , n3634 , n3635 , n3636 , n3638 , n3640 , n3643 , n3644 , n3647 , n3648 , 
n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3657 , n3658 , n3659 , 
n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , 
n3670 , n3671 , n3674 , n3675 , n3677 , n3678 , n3679 , n3680 , n3681 , n3683 , 
n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3694 , n3695 , 
n3699 , n3701 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , 
n3711 , n3713 , n3715 , n3716 , n3717 , n3719 , n3720 , n3722 , n3723 , n3724 , 
n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3733 , n3734 , n3735 , n3736 , 
n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , 
n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3757 , n3759 , n3760 , 
n3761 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , 
n3772 , n3773 , n3774 , n3775 , n3777 , n3779 , n3780 , n3781 , n3782 , n3783 , 
n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , 
n3797 , n3798 , n3799 , n3800 , n3802 , n3803 , n3804 , n3805 , n3806 , n3810 , 
n3811 , n3812 , n3813 , n3815 , n3816 , n3817 , n3818 , n3821 , n3823 , n3824 , 
n3825 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , 
n3838 , n3839 , n3840 , n3841 , n3842 , n3844 , n3845 , n3846 , n3847 , n3849 , 
n3850 , n3851 , n3852 , n3853 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , 
n3861 , n3862 , n3863 ;
    nor g0 ( n1931 , n3561 , n2114 );
    not g1 ( n3069 , n3374 );
    or g2 ( n1111 , n3723 , n2902 );
    and g3 ( n3110 , n3037 , n3559 );
    or g4 ( n224 , n1754 , n832 );
    and g5 ( n3192 , n2978 , n3662 );
    nor g6 ( n651 , n1413 , n3747 );
    nor g7 ( n3113 , n1355 , n1999 );
    or g8 ( n1544 , n820 , n3665 );
    and g9 ( n2935 , n941 , n3553 );
    and g10 ( n978 , n1251 , n2071 );
    and g11 ( n989 , n1350 , n946 );
    or g12 ( n1989 , n346 , n3258 );
    and g13 ( n3527 , n2562 , n2597 );
    nor g14 ( n747 , n788 , n2030 );
    nor g15 ( n2320 , n2154 , n1021 );
    or g16 ( n647 , n2640 , n1332 );
    or g17 ( n2583 , n3025 , n1291 );
    nor g18 ( n3414 , n1573 , n3170 );
    nor g19 ( n2207 , n1086 , n1124 );
    and g20 ( n567 , n2371 , n3858 );
    nor g21 ( n2202 , n409 , n2447 );
    and g22 ( n210 , n944 , n971 );
    nor g23 ( n2083 , n3094 , n343 );
    and g24 ( n2850 , n267 , n1928 );
    nor g25 ( n632 , n1739 , n197 );
    or g26 ( n2822 , n902 , n1480 );
    nor g27 ( n2639 , n2780 , n1530 );
    not g28 ( n1767 , n3754 );
    nor g29 ( n2579 , n130 , n2725 );
    nor g30 ( n442 , n1216 , n3013 );
    and g31 ( n2229 , n289 , n978 );
    and g32 ( n1089 , n3013 , n1216 );
    and g33 ( n3193 , n2626 , n1848 );
    and g34 ( n3640 , n3426 , n2199 );
    nor g35 ( n392 , n2697 , n1444 );
    or g36 ( n1104 , n1471 , n2687 );
    or g37 ( n2252 , n3748 , n202 );
    and g38 ( n1362 , n3061 , n1598 );
    or g39 ( n3176 , n473 , n1939 );
    and g40 ( n2220 , n3771 , n3803 );
    nor g41 ( n3800 , n1258 , n3702 );
    nor g42 ( n3094 , n1346 , n286 );
    or g43 ( n3796 , n3582 , n3241 );
    nor g44 ( n283 , n3782 , n3021 );
    or g45 ( n2899 , n2224 , n3166 );
    and g46 ( n2984 , n2304 , n2381 );
    and g47 ( n3249 , n2334 , n2051 );
    not g48 ( n1145 , n2865 );
    not g49 ( n603 , n558 );
    not g50 ( n1032 , n2543 );
    nor g51 ( n2066 , n3678 , n3759 );
    and g52 ( n2826 , n102 , n3764 );
    nor g53 ( n2039 , n2909 , n3803 );
    nor g54 ( n1337 , n3839 , n3484 );
    nor g55 ( n1902 , n759 , n3250 );
    not g56 ( n2708 , n3592 );
    and g57 ( n2035 , n396 , n772 );
    or g58 ( n2172 , n2654 , n1368 );
    not g59 ( n3077 , n2985 );
    not g60 ( n1978 , n229 );
    or g61 ( n1501 , n3371 , n2849 );
    nor g62 ( n3507 , n723 , n3168 );
    not g63 ( n2877 , n1254 );
    or g64 ( n1883 , n1460 , n3053 );
    or g65 ( n3140 , n1438 , n2735 );
    or g66 ( n1158 , n2937 , n1879 );
    and g67 ( n2262 , n2651 , n66 );
    or g68 ( n1440 , n3757 , n3235 );
    not g69 ( n314 , n820 );
    nor g70 ( n1277 , n870 , n3829 );
    not g71 ( n1048 , n584 );
    or g72 ( n1239 , n3469 , n2089 );
    not g73 ( n3765 , n3625 );
    nor g74 ( n769 , n3260 , n761 );
    nor g75 ( n313 , n3552 , n1072 );
    not g76 ( n2763 , n3785 );
    nor g77 ( n653 , n3725 , n2708 );
    nor g78 ( n1131 , n1170 , n3185 );
    not g79 ( n3217 , n2049 );
    nor g80 ( n3766 , n1685 , n3806 );
    nor g81 ( n2055 , n1371 , n1899 );
    and g82 ( n1173 , n1608 , n365 );
    nor g83 ( n3587 , n3519 , n3477 );
    nor g84 ( n1946 , n272 , n3571 );
    nor g85 ( n830 , n2411 , n54 );
    not g86 ( n1603 , n3372 );
    nor g87 ( n3100 , n2448 , n3553 );
    or g88 ( n1814 , n2405 , n2200 );
    nor g89 ( n2695 , n3257 , n1890 );
    and g90 ( n192 , n3781 , n2066 );
    or g91 ( n756 , n2292 , n2139 );
    or g92 ( n332 , n721 , n3707 );
    not g93 ( n37 , n3576 );
    nor g94 ( n1193 , n1535 , n691 );
    nor g95 ( n3792 , n907 , n2883 );
    or g96 ( n2501 , n899 , n3236 );
    or g97 ( n1249 , n2578 , n1554 );
    nor g98 ( n2593 , n2461 , n2826 );
    or g99 ( n2000 , n81 , n1985 );
    or g100 ( n727 , n146 , n3746 );
    and g101 ( n2689 , n3343 , n1114 );
    nor g102 ( n1956 , n2645 , n345 );
    nor g103 ( n1869 , n1347 , n253 );
    and g104 ( n3261 , n2353 , n1199 );
    and g105 ( n1257 , n2226 , n1388 );
    and g106 ( n1588 , n1452 , n2152 );
    nor g107 ( n3458 , n3473 , n2392 );
    and g108 ( n810 , n2131 , n1721 );
    nor g109 ( n3334 , n2520 , n896 );
    not g110 ( n1484 , n3049 );
    nor g111 ( n1338 , n2540 , n837 );
    not g112 ( n3294 , n2169 );
    or g113 ( n1903 , n3240 , n1821 );
    nor g114 ( n717 , n830 , n287 );
    or g115 ( n3426 , n1068 , n1554 );
    or g116 ( n3599 , n2590 , n1878 );
    not g117 ( n1598 , n2776 );
    not g118 ( n1034 , n3418 );
    and g119 ( n1162 , n3126 , n3616 );
    or g120 ( n1644 , n567 , n1492 );
    or g121 ( n145 , n75 , n1774 );
    and g122 ( n3581 , n2166 , n596 );
    and g123 ( n1784 , n2333 , n31 );
    nor g124 ( n89 , n2427 , n3223 );
    not g125 ( n3803 , n2776 );
    or g126 ( n154 , n80 , n3010 );
    or g127 ( n1591 , n2359 , n3287 );
    nor g128 ( n746 , n2299 , n3631 );
    or g129 ( n1019 , n3487 , n1798 );
    or g130 ( n3295 , n702 , n1784 );
    or g131 ( n714 , n3188 , n789 );
    or g132 ( n1025 , n3149 , n3182 );
    or g133 ( n2400 , n1990 , n1729 );
    nor g134 ( n319 , n2865 , n95 );
    and g135 ( n2224 , n3373 , n2324 );
    or g136 ( n330 , n2236 , n3765 );
    or g137 ( n2502 , n3100 , n2205 );
    not g138 ( n1925 , n208 );
    and g139 ( n3282 , n1435 , n2829 );
    or g140 ( n1514 , n60 , n843 );
    or g141 ( n1343 , n30 , n2345 );
    or g142 ( n2660 , n2460 , n3309 );
    nor g143 ( n5 , n2907 , n1279 );
    nor g144 ( n650 , n1980 , n3664 );
    not g145 ( n1739 , n2962 );
    or g146 ( n1079 , n3129 , n3507 );
    not g147 ( n344 , n3035 );
    nor g148 ( n2749 , n2511 , n858 );
    not g149 ( n1140 , n2616 );
    or g150 ( n757 , n3572 , n2009 );
    nor g151 ( n494 , n1855 , n3598 );
    or g152 ( n846 , n1035 , n3026 );
    nor g153 ( n3602 , n3417 , n1539 );
    not g154 ( n3729 , n3570 );
    or g155 ( n3014 , n3031 , n2553 );
    and g156 ( n905 , n727 , n1520 );
    or g157 ( n12 , n3415 , n1235 );
    nor g158 ( n3562 , n3628 , n3553 );
    nor g159 ( n3326 , n3653 , n397 );
    nor g160 ( n2395 , n744 , n2887 );
    nor g161 ( n3204 , n627 , n2354 );
    not g162 ( n1675 , n2151 );
    or g163 ( n2694 , n1862 , n1377 );
    and g164 ( n2574 , n1602 , n2740 );
    nor g165 ( n2828 , n2242 , n341 );
    not g166 ( n3012 , n248 );
    or g167 ( n3683 , n2059 , n1210 );
    or g168 ( n2494 , n3331 , n3347 );
    or g169 ( n763 , n1017 , n1208 );
    nor g170 ( n2008 , n889 , n2660 );
    not g171 ( n1546 , n3188 );
    or g172 ( n444 , n267 , n1928 );
    and g173 ( n148 , n1806 , n3397 );
    or g174 ( n3039 , n9 , n3720 );
    not g175 ( n3333 , n2693 );
    and g176 ( n1476 , n2469 , n2061 );
    nor g177 ( n200 , n10 , n2526 );
    and g178 ( n731 , n1599 , n929 );
    nor g179 ( n48 , n1182 , n2467 );
    nor g180 ( n3384 , n3405 , n2634 );
    and g181 ( n1763 , n1075 , n509 );
    nor g182 ( n2672 , n3697 , n3090 );
    or g183 ( n3737 , n23 , n3237 );
    nor g184 ( n245 , n2268 , n691 );
    nor g185 ( n2210 , n2016 , n1701 );
    and g186 ( n238 , n804 , n427 );
    nor g187 ( n412 , n3525 , n1673 );
    or g188 ( n1799 , n3319 , n905 );
    nor g189 ( n1124 , n2271 , n105 );
    and g190 ( n3237 , n3322 , n251 );
    and g191 ( n2364 , n1786 , n3569 );
    nor g192 ( n1560 , n2397 , n2298 );
    not g193 ( n2737 , n3801 );
    or g194 ( n2150 , n138 , n1901 );
    nor g195 ( n3500 , n2962 , n2799 );
    not g196 ( n3743 , n700 );
    and g197 ( n1292 , n1954 , n1628 );
    nor g198 ( n2568 , n1812 , n3430 );
    nor g199 ( n3520 , n2183 , n3623 );
    or g200 ( n1651 , n841 , n3665 );
    nor g201 ( n19 , n1001 , n2046 );
    nor g202 ( n3716 , n1125 , n2339 );
    or g203 ( n1912 , n1314 , n1126 );
    nor g204 ( n355 , n881 , n2670 );
    and g205 ( n2276 , n2555 , n358 );
    nor g206 ( n1321 , n1734 , n914 );
    or g207 ( n1273 , n3114 , n3601 );
    or g208 ( n2064 , n3686 , n2901 );
    or g209 ( n3177 , n2572 , n1929 );
    nor g210 ( n346 , n2662 , n1137 );
    not g211 ( n2604 , n1785 );
    nor g212 ( n206 , n197 , n2026 );
    and g213 ( n1988 , n3014 , n1013 );
    not g214 ( n736 , n2668 );
    or g215 ( n341 , n3772 , n2744 );
    or g216 ( n2596 , n1682 , n1235 );
    and g217 ( n1489 , n1684 , n2382 );
    not g218 ( n1673 , n3592 );
    nor g219 ( n2807 , n246 , n611 );
    or g220 ( n3649 , n494 , n1725 );
    or g221 ( n2154 , n2011 , n2081 );
    nor g222 ( n2993 , n3266 , n2243 );
    nor g223 ( n1567 , n3142 , n2232 );
    nor g224 ( n938 , n1061 , n1012 );
    and g225 ( n3027 , n1273 , n2265 );
    nor g226 ( n3392 , n1524 , n43 );
    nor g227 ( n1050 , n1298 , n95 );
    or g228 ( n2012 , n764 , n956 );
    nor g229 ( n575 , n3415 , n2450 );
    nor g230 ( n869 , n2779 , n3244 );
    or g231 ( n1151 , n3308 , n3840 );
    not g232 ( n3397 , n40 );
    and g233 ( n1154 , n1170 , n3012 );
    or g234 ( n2309 , n1416 , n3184 );
    or g235 ( n2538 , n1811 , n2284 );
    nor g236 ( n3123 , n2742 , n1736 );
    or g237 ( n1178 , n2003 , n799 );
    not g238 ( n2924 , n848 );
    and g239 ( n3859 , n3850 , n1600 );
    or g240 ( n437 , n1139 , n2532 );
    or g241 ( n3071 , n1476 , n1668 );
    nor g242 ( n367 , n949 , n3047 );
    nor g243 ( n1487 , n1970 , n2612 );
    and g244 ( n997 , n1884 , n3440 );
    or g245 ( n1036 , n1106 , n1843 );
    or g246 ( n3663 , n349 , n1385 );
    nor g247 ( n2610 , n1634 , n323 );
    nor g248 ( n795 , n1806 , n1219 );
    and g249 ( n1888 , n275 , n543 );
    nor g250 ( n1959 , n200 , n2395 );
    nor g251 ( n2581 , n1654 , n3598 );
    or g252 ( n2788 , n394 , n3298 );
    nor g253 ( n3149 , n3730 , n3805 );
    and g254 ( n1517 , n1782 , n1891 );
    nor g255 ( n2506 , n1917 , n2893 );
    or g256 ( n1148 , n239 , n3406 );
    not g257 ( n3191 , n2253 );
    and g258 ( n2208 , n272 , n3571 );
    and g259 ( n3612 , n989 , n3553 );
    nor g260 ( n1693 , n2275 , n2784 );
    nor g261 ( n3342 , n979 , n2386 );
    or g262 ( n2995 , n2782 , n626 );
    not g263 ( n3259 , n3168 );
    nor g264 ( n463 , n2766 , n1603 );
    or g265 ( n1452 , n1044 , n3582 );
    and g266 ( n347 , n3858 , n1598 );
    or g267 ( n1744 , n3528 , n3282 );
    or g268 ( n1633 , n1885 , n1914 );
    not g269 ( n2748 , n2297 );
    nor g270 ( n473 , n3341 , n3819 );
    nor g271 ( n777 , n3413 , n1014 );
    or g272 ( n3793 , n2216 , n2026 );
    and g273 ( n17 , n2283 , n974 );
    or g274 ( n16 , n853 , n410 );
    or g275 ( n1887 , n11 , n3202 );
    or g276 ( n1409 , n2480 , n2504 );
    or g277 ( n114 , n1036 , n220 );
    nor g278 ( n1761 , n1215 , n3452 );
    and g279 ( n874 , n235 , n993 );
    and g280 ( n2952 , n514 , n2964 );
    or g281 ( n2465 , n3316 , n1417 );
    and g282 ( n876 , n1553 , n2231 );
    and g283 ( n3242 , n2848 , n3297 );
    or g284 ( n564 , n1570 , n2516 );
    and g285 ( n3227 , n336 , n2710 );
    or g286 ( n3330 , n375 , n2028 );
    or g287 ( n3614 , n3269 , n738 );
    and g288 ( n190 , n1287 , n2381 );
    nor g289 ( n3674 , n1119 , n2074 );
    or g290 ( n1425 , n1851 , n3846 );
    nor g291 ( n3108 , n2996 , n3641 );
    nor g292 ( n324 , n2280 , n1132 );
    nor g293 ( n2770 , n1346 , n2595 );
    nor g294 ( n3205 , n1709 , n2438 );
    nor g295 ( n659 , n3255 , n760 );
    nor g296 ( n1349 , n3621 , n3154 );
    and g297 ( n1808 , n669 , n2824 );
    and g298 ( n3230 , n3833 , n64 );
    or g299 ( n1745 , n290 , n581 );
    and g300 ( n3151 , n1974 , n2114 );
    nor g301 ( n2011 , n2405 , n2509 );
    or g302 ( n282 , n1316 , n3273 );
    not g303 ( n936 , n726 );
    nor g304 ( n3564 , n3480 , n3130 );
    and g305 ( n3853 , n1552 , n300 );
    not g306 ( n2888 , n1139 );
    nor g307 ( n3093 , n3534 , n2545 );
    or g308 ( n1378 , n950 , n1839 );
    and g309 ( n1810 , n875 , n2597 );
    and g310 ( n3146 , n3027 , n64 );
    and g311 ( n2555 , n284 , n2722 );
    or g312 ( n2728 , n176 , n2168 );
    and g313 ( n3545 , n3319 , n905 );
    and g314 ( n3111 , n2586 , n2667 );
    nor g315 ( n2063 , n1069 , n524 );
    or g316 ( n3515 , n3422 , n1142 );
    or g317 ( n917 , n617 , n2903 );
    or g318 ( n1488 , n377 , n3656 );
    nor g319 ( n2050 , n2134 , n2610 );
    nor g320 ( n760 , n740 , n3028 );
    not g321 ( n2087 , n3743 );
    or g322 ( n801 , n1451 , n3346 );
    not g323 ( n1977 , n3578 );
    not g324 ( n1385 , n2665 );
    nor g325 ( n3329 , n44 , n1072 );
    or g326 ( n302 , n417 , n1220 );
    nor g327 ( n2077 , n965 , n1114 );
    or g328 ( n3468 , n3073 , n1154 );
    not g329 ( n68 , n2248 );
    or g330 ( n1614 , n1079 , n2567 );
    nor g331 ( n2144 , n1498 , n3315 );
    or g332 ( n3115 , n1510 , n2625 );
    nor g333 ( n2566 , n2642 , n1301 );
    nor g334 ( n1278 , n1221 , n3852 );
    not g335 ( n1724 , n1474 );
    or g336 ( n2427 , n3613 , n305 );
    nor g337 ( n1441 , n3 , n2633 );
    nor g338 ( n3354 , n409 , n3833 );
    or g339 ( n2179 , n1995 , n2658 );
    or g340 ( n3483 , n1846 , n949 );
    nor g341 ( n517 , n1626 , n952 );
    nor g342 ( n3074 , n610 , n2932 );
    and g343 ( n1336 , n3480 , n3130 );
    nor g344 ( n3118 , n768 , n3857 );
    and g345 ( n1267 , n876 , n2757 );
    or g346 ( n2354 , n2888 , n2681 );
    not g347 ( n1668 , n3037 );
    nor g348 ( n2943 , n1358 , n2296 );
    not g349 ( n2254 , n1834 );
    nor g350 ( n2784 , n453 , n2264 );
    or g351 ( n3068 , n522 , n3612 );
    or g352 ( n2342 , n3312 , n1465 );
    not g353 ( n2757 , n2985 );
    nor g354 ( n2102 , n1456 , n3120 );
    and g355 ( n75 , n1876 , n1445 );
    nor g356 ( n2785 , n580 , n3644 );
    and g357 ( n960 , n3358 , n1292 );
    not g358 ( n3523 , n97 );
    not g359 ( n1212 , n1324 );
    and g360 ( n3355 , n3243 , n739 );
    and g361 ( n3120 , n461 , n3830 );
    nor g362 ( n1105 , n955 , n1525 );
    nor g363 ( n828 , n2390 , n2539 );
    or g364 ( n2143 , n2133 , n447 );
    nor g365 ( n2655 , n236 , n2026 );
    nor g366 ( n3303 , n2361 , n1986 );
    and g367 ( n3277 , n2906 , n2249 );
    and g368 ( n1755 , n196 , n1897 );
    nor g369 ( n3775 , n3338 , n1571 );
    and g370 ( n3343 , n2005 , n2970 );
    and g371 ( n1552 , n1303 , n2947 );
    and g372 ( n213 , n1986 , n64 );
    nor g373 ( n3357 , n1684 , n3803 );
    nor g374 ( n1670 , n3444 , n926 );
    and g375 ( n2700 , n227 , n3595 );
    or g376 ( n3393 , n3008 , n452 );
    and g377 ( n954 , n127 , n484 );
    not g378 ( n1190 , n700 );
    nor g379 ( n3296 , n3585 , n3598 );
    or g380 ( n2873 , n1203 , n2839 );
    nor g381 ( n834 , n1275 , n1887 );
    nor g382 ( n293 , n1028 , n1576 );
    not g383 ( n984 , n2255 );
    not g384 ( n1563 , n3718 );
    or g385 ( n965 , n2481 , n1400 );
    or g386 ( n431 , n3259 , n523 );
    and g387 ( n1980 , n198 , n3265 );
    or g388 ( n2391 , n1871 , n1269 );
    or g389 ( n3768 , n3085 , n3425 );
    nor g390 ( n1898 , n608 , n157 );
    or g391 ( n414 , n2541 , n1343 );
    and g392 ( n2624 , n1721 , n772 );
    nor g393 ( n2356 , n2448 , n141 );
    nor g394 ( n82 , n3839 , n1598 );
    and g395 ( n250 , n286 , n2087 );
    or g396 ( n1403 , n2779 , n2513 );
    or g397 ( n2820 , n2371 , n3858 );
    and g398 ( n901 , n2382 , n3032 );
    and g399 ( n3223 , n2290 , n1073 );
    nor g400 ( n2136 , n1379 , n3441 );
    and g401 ( n1123 , n1926 , n1642 );
    nor g402 ( n3699 , n1989 , n3032 );
    or g403 ( n1868 , n1264 , n51 );
    nor g404 ( n2965 , n2079 , n1037 );
    not g405 ( n2053 , n2185 );
    nor g406 ( n2306 , n2479 , n3494 );
    not g407 ( n1870 , n2263 );
    nor g408 ( n2322 , n3254 , n3615 );
    or g409 ( n2498 , n928 , n1562 );
    not g410 ( n150 , n1190 );
    nor g411 ( n576 , n3563 , n2228 );
    or g412 ( n1981 , n708 , n2076 );
    nor g413 ( n3431 , n3216 , n1819 );
    and g414 ( n672 , n809 , n655 );
    nor g415 ( n2887 , n1098 , n1991 );
    and g416 ( n2805 , n1397 , n2604 );
    and g417 ( n1464 , n2135 , n2757 );
    nor g418 ( n2480 , n2309 , n150 );
    nor g419 ( n350 , n3274 , n64 );
    nor g420 ( n3102 , n1797 , n1761 );
    not g421 ( n3526 , n3525 );
    nor g422 ( n478 , n1327 , n3278 );
    and g423 ( n1818 , n3436 , n497 );
    and g424 ( n2504 , n3481 , n322 );
    or g425 ( n982 , n2883 , n1484 );
    and g426 ( n2042 , n1300 , n143 );
    or g427 ( n719 , n2861 , n2341 );
    and g428 ( n1472 , n2882 , n2527 );
    or g429 ( n88 , n3058 , n2577 );
    nor g430 ( n3167 , n1849 , n2914 );
    and g431 ( n2669 , n1449 , n195 );
    not g432 ( n2114 , n726 );
    or g433 ( n299 , n3687 , n108 );
    or g434 ( n457 , n2573 , n1274 );
    or g435 ( n2361 , n3500 , n206 );
    and g436 ( n549 , n3167 , n116 );
    or g437 ( n2755 , n336 , n1484 );
    not g438 ( n993 , n1068 );
    nor g439 ( n249 , n1587 , n2442 );
    and g440 ( n2227 , n838 , n500 );
    nor g441 ( n21 , n904 , n611 );
    nor g442 ( n3631 , n2641 , n2267 );
    nor g443 ( n91 , n3734 , n923 );
    not g444 ( n3578 , n2352 );
    not g445 ( n3547 , n2644 );
    and g446 ( n3196 , n2883 , n907 );
    not g447 ( n43 , n790 );
    nor g448 ( n2861 , n893 , n2550 );
    nor g449 ( n2982 , n344 , n2668 );
    nor g450 ( n2548 , n1713 , n1265 );
    or g451 ( n3410 , n2677 , n3159 );
    and g452 ( n2681 , n1999 , n1355 );
    not g453 ( n3861 , n667 );
    and g454 ( n1227 , n802 , n705 );
    and g455 ( n396 , n2082 , n1747 );
    nor g456 ( n794 , n1521 , n247 );
    nor g457 ( n963 , n3250 , n3593 );
    nor g458 ( n1316 , n475 , n93 );
    and g459 ( n1157 , n2527 , n3553 );
    not g460 ( n1985 , n1140 );
    not g461 ( n480 , n796 );
    and g462 ( n1480 , n2787 , n1905 );
    nor g463 ( n2516 , n1650 , n1536 );
    or g464 ( n3327 , n2771 , n1464 );
    nor g465 ( n2294 , n2960 , n795 );
    or g466 ( n2173 , n3333 , n2731 );
    not g467 ( n2029 , n2550 );
    or g468 ( n2141 , n605 , n1592 );
    or g469 ( n2729 , n2843 , n3746 );
    not g470 ( n1114 , n2776 );
    nor g471 ( n2931 , n2 , n2773 );
    or g472 ( n707 , n468 , n1376 );
    not g473 ( n3081 , n3060 );
    nor g474 ( n1793 , n984 , n1631 );
    or g475 ( n854 , n2990 , n1235 );
    or g476 ( n3433 , n1546 , n176 );
    and g477 ( n2181 , n2180 , n669 );
    nor g478 ( n3535 , n1599 , n3217 );
    or g479 ( n602 , n1439 , n2187 );
    or g480 ( n1366 , n1716 , n3363 );
    not g481 ( n500 , n3848 );
    and g482 ( n3548 , n2491 , n3770 );
    and g483 ( n716 , n3336 , n595 );
    nor g484 ( n2497 , n3191 , n873 );
    and g485 ( n1169 , n3066 , n2925 );
    or g486 ( n2954 , n3713 , n504 );
    nor g487 ( n1826 , n3807 , n2708 );
    not g488 ( n3625 , n2616 );
    or g489 ( n1608 , n1179 , n1682 );
    not g490 ( n3220 , n433 );
    and g491 ( n13 , n44 , n1109 );
    not g492 ( n294 , n2896 );
    or g493 ( n512 , n2415 , n659 );
    nor g494 ( n3239 , n132 , n1698 );
    nor g495 ( n31 , n1056 , n2487 );
    and g496 ( n70 , n1289 , n1041 );
    not g497 ( n3316 , n3843 );
    nor g498 ( n3424 , n2477 , n1828 );
    nor g499 ( n3429 , n2449 , n896 );
    nor g500 ( n1174 , n2371 , n3829 );
    or g501 ( n1146 , n2323 , n313 );
    nor g502 ( n2092 , n971 , n924 );
    nor g503 ( n1431 , n998 , n3335 );
    nor g504 ( n2968 , n2613 , n1357 );
    nor g505 ( n2225 , n124 , n3630 );
    nor g506 ( n1507 , n3460 , n407 );
    or g507 ( n2319 , n3801 , n1985 );
    or g508 ( n3560 , n3755 , n2105 );
    or g509 ( n1867 , n2015 , n2454 );
    or g510 ( n2588 , n1160 , n2762 );
    or g511 ( n831 , n1805 , n3665 );
    or g512 ( n2197 , n2255 , n859 );
    or g513 ( n826 , n1859 , n2255 );
    not g514 ( n1864 , n3025 );
    and g515 ( n2203 , n541 , n111 );
    and g516 ( n1502 , n1720 , n3533 );
    nor g517 ( n2175 , n1884 , n3069 );
    nor g518 ( n2264 , n2412 , n1506 );
    nor g519 ( n3835 , n3708 , n2889 );
    or g520 ( n1553 , n1232 , n2532 );
    and g521 ( n3085 , n3314 , n2897 );
    nor g522 ( n3159 , n1675 , n2328 );
    and g523 ( n3546 , n3109 , n1614 );
    nor g524 ( n403 , n1582 , n2243 );
    nor g525 ( n1772 , n2235 , n1612 );
    not g526 ( n3032 , n1190 );
    or g527 ( n1908 , n2614 , n3485 );
    nor g528 ( n1510 , n3729 , n1708 );
    not g529 ( n2698 , n2726 );
    or g530 ( n3694 , n1122 , n1655 );
    or g531 ( n3198 , n1926 , n2168 );
    or g532 ( n3696 , n2056 , n3155 );
    or g533 ( n1060 , n752 , n3836 );
    and g534 ( n498 , n1667 , n2873 );
    nor g535 ( n1215 , n545 , n3465 );
    not g536 ( n2221 , n2572 );
    or g537 ( n1058 , n3701 , n3789 );
    and g538 ( n1705 , n1788 , n2391 );
    nor g539 ( n2658 , n130 , n814 );
    and g540 ( n460 , n2863 , n906 );
    nor g541 ( n566 , n804 , n1539 );
    nor g542 ( n824 , n1748 , n226 );
    or g543 ( n1009 , n3145 , n3148 );
    nor g544 ( n1717 , n1266 , n756 );
    and g545 ( n2009 , n2813 , n3077 );
    and g546 ( n144 , n2156 , n1598 );
    or g547 ( n783 , n3107 , n270 );
    and g548 ( n863 , n1434 , n2562 );
    or g549 ( n3178 , n3854 , n3148 );
    not g550 ( n592 , n2433 );
    or g551 ( n2621 , n3324 , n2793 );
    nor g552 ( n2659 , n2911 , n3210 );
    or g553 ( n1920 , n3173 , n1084 );
    nor g554 ( n2282 , n3323 , n2799 );
    or g555 ( n2277 , n3296 , n1470 );
    nor g556 ( n787 , n3636 , n1601 );
    or g557 ( n1396 , n2076 , n3765 );
    nor g558 ( n3015 , n3457 , n2060 );
    nor g559 ( n1976 , n1804 , n3583 );
    not g560 ( n543 , n3203 );
    nor g561 ( n3019 , n1746 , n3272 );
    nor g562 ( n230 , n406 , n2990 );
    and g563 ( n3774 , n1691 , n318 );
    nor g564 ( n2571 , n1495 , n1072 );
    and g565 ( n1924 , n2339 , n1125 );
    and g566 ( n2666 , n2736 , n2698 );
    and g567 ( n2836 , n409 , n3833 );
    nor g568 ( n1513 , n2711 , n896 );
    or g569 ( n3671 , n3421 , n2452 );
    nor g570 ( n112 , n2054 , n1750 );
    nor g571 ( n507 , n528 , n143 );
    nor g572 ( n2192 , n1149 , n697 );
    nor g573 ( n147 , n3186 , n3842 );
    or g574 ( n2848 , n3150 , n3219 );
    or g575 ( n1657 , n1782 , n1891 );
    nor g576 ( n3813 , n2149 , n2590 );
    or g577 ( n2226 , n1384 , n3556 );
    nor g578 ( n1069 , n2410 , n3525 );
    nor g579 ( n3209 , n3283 , n3384 );
    not g580 ( n3281 , n1451 );
    or g581 ( n408 , n2186 , n2638 );
    not g582 ( n2458 , n1045 );
    nor g583 ( n421 , n3590 , n1537 );
    nor g584 ( n3678 , n818 , n1250 );
    and g585 ( n120 , n1775 , n3316 );
    and g586 ( n1191 , n1405 , n3540 );
    or g587 ( n2209 , n627 , n3765 );
    or g588 ( n1857 , n1774 , n2783 );
    and g589 ( n700 , n1331 , n1940 );
    and g590 ( n504 , n3640 , n2757 );
    nor g591 ( n1811 , n1121 , n1162 );
    nor g592 ( n2249 , n180 , n666 );
    not g593 ( n1156 , n1605 );
    nor g594 ( n484 , n2419 , n3520 );
    or g595 ( n2448 , n566 , n337 );
    or g596 ( n550 , n1631 , n2921 );
    and g597 ( n2986 , n891 , n2135 );
    nor g598 ( n1714 , n2018 , n1650 );
    not g599 ( n1878 , n972 );
    nor g600 ( n3439 , n521 , n640 );
    not g601 ( n618 , n1420 );
    not g602 ( n32 , n2484 );
    and g603 ( n556 , n2503 , n2518 );
    or g604 ( n3554 , n569 , n1858 );
    and g605 ( n807 , n2526 , n2595 );
    and g606 ( n2530 , n1611 , n1951 );
    nor g607 ( n559 , n3393 , n1603 );
    or g608 ( n1556 , n3574 , n1955 );
    or g609 ( n973 , n2185 , n2921 );
    or g610 ( n1339 , n3311 , n2027 );
    nor g611 ( n3064 , n338 , n3815 );
    or g612 ( n690 , n1063 , n3591 );
    nor g613 ( n565 , n3365 , n1018 );
    nor g614 ( n622 , n887 , n2083 );
    and g615 ( n1721 , n992 , n2319 );
    nor g616 ( n1011 , n2791 , n2068 );
    nor g617 ( n39 , n1523 , n3229 );
    and g618 ( n3271 , n1129 , n3077 );
    nor g619 ( n3065 , n1260 , n2041 );
    or g620 ( n1650 , n1128 , n986 );
    nor g621 ( n1335 , n492 , n2835 );
    or g622 ( n689 , n2959 , n613 );
    and g623 ( n3067 , n545 , n3465 );
    nor g624 ( n1837 , n3087 , n3684 );
    or g625 ( n1046 , n2178 , n422 );
    nor g626 ( n656 , n873 , n640 );
    or g627 ( n533 , n2897 , n635 );
    and g628 ( n3619 , n2729 , n1511 );
    and g629 ( n3770 , n1342 , n295 );
    and g630 ( n2369 , n1029 , n1107 );
    or g631 ( n983 , n2029 , n298 );
    or g632 ( n3279 , n2805 , n1123 );
    and g633 ( n2435 , n1591 , n1919 );
    nor g634 ( n1133 , n837 , n665 );
    and g635 ( n1223 , n2325 , n3558 );
    or g636 ( n1150 , n574 , n3346 );
    nor g637 ( n3779 , n1602 , n226 );
    or g638 ( n3174 , n1002 , n1263 );
    or g639 ( n1919 , n3677 , n2388 );
    nor g640 ( n1400 , n1118 , n2298 );
    or g641 ( n1933 , n2619 , n158 );
    and g642 ( n635 , n2890 , n3362 );
    and g643 ( n1469 , n2260 , n271 );
    not g644 ( n529 , n3266 );
    and g645 ( n1783 , n3278 , n1327 );
    and g646 ( n1948 , n1463 , n1290 );
    nor g647 ( n935 , n2879 , n3051 );
    nor g648 ( n2585 , n1728 , n2715 );
    nor g649 ( n939 , n2453 , n1824 );
    nor g650 ( n3292 , n2380 , n661 );
    and g651 ( n1612 , n1561 , n2351 );
    not g652 ( n1905 , n2611 );
    or g653 ( n1727 , n3446 , n402 );
    or g654 ( n2991 , n1367 , n3110 );
    nor g655 ( n258 , n217 , n3583 );
    nor g656 ( n2959 , n2607 , n400 );
    nor g657 ( n290 , n1695 , n782 );
    nor g658 ( n2137 , n2955 , n2778 );
    and g659 ( n1839 , n3193 , n2597 );
    or g660 ( n604 , n3081 , n2297 );
    and g661 ( n1809 , n3052 , n2795 );
    or g662 ( n1910 , n467 , n2168 );
    nor g663 ( n1195 , n2488 , n1539 );
    or g664 ( n1737 , n1319 , n812 );
    and g665 ( n547 , n302 , n306 );
    or g666 ( n486 , n1999 , n1798 );
    or g667 ( n3255 , n3189 , n264 );
    nor g668 ( n2573 , n1015 , n1977 );
    or g669 ( n2373 , n2774 , n1369 );
    nor g670 ( n1402 , n2698 , n2736 );
    not g671 ( n1179 , n3335 );
    nor g672 ( n1264 , n947 , n1539 );
    or g673 ( n3404 , n1882 , n1077 );
    nor g674 ( n1786 , n1632 , n332 );
    or g675 ( n2318 , n3076 , n3306 );
    or g676 ( n713 , n3376 , n3647 );
    nor g677 ( n3225 , n2361 , n3553 );
    not g678 ( n2685 , n3288 );
    nor g679 ( n1053 , n2491 , n64 );
    nor g680 ( n3825 , n3013 , n3583 );
    nor g681 ( n34 , n1259 , n2708 );
    or g682 ( n3747 , n1016 , n459 );
    or g683 ( n1983 , n3001 , n789 );
    and g684 ( n3508 , n2194 , n3056 );
    nor g685 ( n3466 , n728 , n2392 );
    not g686 ( n3558 , n2661 );
    or g687 ( n2244 , n1402 , n1757 );
    and g688 ( n1269 , n2643 , n890 );
    and g689 ( n3309 , n2390 , n1816 );
    not g690 ( n998 , n1682 );
    not g691 ( n1327 , n947 );
    nor g692 ( n133 , n2147 , n2595 );
    not g693 ( n3374 , n1389 );
    not g694 ( n1125 , n1200 );
    nor g695 ( n734 , n2052 , n1037 );
    nor g696 ( n3509 , n2048 , n2124 );
    nor g697 ( n1283 , n3133 , n1698 );
    not g698 ( n1044 , n1471 );
    and g699 ( n2123 , n224 , n1974 );
    and g700 ( n3446 , n931 , n3550 );
    not g701 ( n2375 , n2971 );
    and g702 ( n42 , n1841 , n2223 );
    nor g703 ( n3162 , n2550 , n1537 );
    nor g704 ( n92 , n3023 , n2566 );
    nor g705 ( n3723 , n631 , n1673 );
    nor g706 ( n335 , n868 , n1259 );
    nor g707 ( n2232 , n1328 , n864 );
    nor g708 ( n1384 , n1222 , n2708 );
    and g709 ( n2987 , n1504 , n2794 );
    nor g710 ( n1921 , n3006 , n3211 );
    or g711 ( n514 , n1217 , n2921 );
    nor g712 ( n84 , n1779 , n3011 );
    or g713 ( n3680 , n97 , n1484 );
    nor g714 ( n2386 , n2495 , n1325 );
    or g715 ( n553 , n2363 , n2086 );
    or g716 ( n1194 , n523 , n3840 );
    and g717 ( n447 , n2378 , n2019 );
    and g718 ( n1930 , n2536 , n3042 );
    or g719 ( n1664 , n1674 , n2101 );
    nor g720 ( n894 , n1624 , n3593 );
    nor g721 ( n3234 , n3726 , n1958 );
    or g722 ( n1896 , n1116 , n1096 );
    and g723 ( n2592 , n74 , n1552 );
    or g724 ( n1967 , n400 , n3148 );
    and g725 ( n119 , n2316 , n425 );
    not g726 ( n2470 , n261 );
    or g727 ( n284 , n2928 , n2921 );
    and g728 ( n212 , n207 , n1585 );
    and g729 ( n364 , n2427 , n3223 );
    not g730 ( n2423 , n1305 );
    nor g731 ( n3477 , n2378 , n3824 );
    and g732 ( n244 , n1292 , n1357 );
    nor g733 ( n1963 , n2458 , n1451 );
    or g734 ( n681 , n1020 , n2468 );
    or g735 ( n1610 , n258 , n1133 );
    or g736 ( n262 , n1974 , n733 );
    and g737 ( n1655 , n2671 , n3744 );
    and g738 ( n2223 , n699 , n12 );
    nor g739 ( n1828 , n3632 , n3487 );
    not g740 ( n665 , n3374 );
    or g741 ( n2138 , n3392 , n1898 );
    nor g742 ( n3810 , n2507 , n3069 );
    or g743 ( n587 , n1454 , n2366 );
    and g744 ( n1262 , n3541 , n3831 );
    or g745 ( n2819 , n2787 , n1985 );
    nor g746 ( n1862 , n1031 , n358 );
    or g747 ( n2680 , n2620 , n2637 );
    not g748 ( n353 , n994 );
    or g749 ( n3307 , n202 , n2088 );
    nor g750 ( n476 , n3065 , n2961 );
    or g751 ( n2463 , n3634 , n2404 );
    nor g752 ( n1526 , n808 , n1550 );
    not g753 ( n1846 , n930 );
    or g754 ( n1792 , n2936 , n1874 );
    or g755 ( n3652 , n2613 , n3619 );
    nor g756 ( n3447 , n1904 , n3090 );
    nor g757 ( n2690 , n2604 , n1397 );
    or g758 ( n2467 , n312 , n3175 );
    or g759 ( n2180 , n1513 , n2259 );
    or g760 ( n1709 , n1892 , n2192 );
    and g761 ( n1360 , n3619 , n64 );
    nor g762 ( n2374 , n2967 , n1873 );
    not g763 ( n968 , n311 );
    or g764 ( n3232 , n2489 , n1639 );
    nor g765 ( n1414 , n503 , n3295 );
    nor g766 ( n1106 , n1759 , n2928 );
    nor g767 ( n2657 , n3074 , n908 );
    nor g768 ( n532 , n903 , n1977 );
    not g769 ( n387 , n1376 );
    or g770 ( n3000 , n850 , n1291 );
    and g771 ( n1265 , n2930 , n3580 );
    or g772 ( n3849 , n160 , n2102 );
    nor g773 ( n2919 , n3609 , n2870 );
    nor g774 ( n2257 , n388 , n2026 );
    or g775 ( n3664 , n1198 , n1768 );
    and g776 ( n2916 , n1275 , n11 );
    nor g777 ( n1093 , n298 , n611 );
    and g778 ( n1519 , n2370 , n322 );
    or g779 ( n596 , n2523 , n2347 );
    nor g780 ( n3324 , n457 , n3217 );
    nor g781 ( n2481 , n3573 , n3598 );
    or g782 ( n3194 , n519 , n2921 );
    and g783 ( n3470 , n1753 , n772 );
    or g784 ( n946 , n3827 , n1085 );
    nor g785 ( n2603 , n2731 , n2243 );
    nor g786 ( n1410 , n621 , n340 );
    nor g787 ( n2122 , n2422 , n3090 );
    nor g788 ( n2291 , n3818 , n936 );
    and g789 ( n923 , n170 , n2376 );
    nor g790 ( n3795 , n3564 , n953 );
    or g791 ( n2383 , n849 , n3411 );
    nor g792 ( n411 , n187 , n3221 );
    not g793 ( n358 , n2482 );
    or g794 ( n758 , n1931 , n2689 );
    nor g795 ( n1911 , n1434 , n2562 );
    or g796 ( n3062 , n3202 , n2099 );
    nor g797 ( n1103 , n2980 , n3808 );
    or g798 ( n3083 , n1193 , n1242 );
    or g799 ( n1802 , n1230 , n1888 );
    nor g800 ( n2387 , n3007 , n2190 );
    or g801 ( n1411 , n398 , n28 );
    nor g802 ( n2674 , n3255 , n3209 );
    or g803 ( n3454 , n3647 , n2430 );
    not g804 ( n1604 , n3508 );
    nor g805 ( n3524 , n2982 , n3618 );
    nor g806 ( n3407 , n878 , n1698 );
    not g807 ( n3669 , n3697 );
    and g808 ( n843 , n3724 , n2674 );
    and g809 ( n3438 , n1923 , n1932 );
    and g810 ( n1600 , n2515 , n2496 );
    not g811 ( n535 , n3743 );
    and g812 ( n453 , n671 , n2813 );
    or g813 ( n1021 , n3108 , n1948 );
    nor g814 ( n158 , n3768 , n369 );
    not g815 ( n2765 , n2166 );
    nor g816 ( n1927 , n2277 , n1598 );
    or g817 ( n2440 , n2528 , n117 );
    not g818 ( n1587 , n3715 );
    and g819 ( n3703 , n1790 , n2373 );
    or g820 ( n2315 , n1453 , n1705 );
    or g821 ( n1345 , n3082 , n2272 );
    not g822 ( n896 , n1295 );
    not g823 ( n818 , n711 );
    nor g824 ( n2084 , n2288 , n1946 );
    nor g825 ( n2963 , n545 , n143 );
    and g826 ( n3306 , n920 , n3692 );
    nor g827 ( n3018 , n658 , n884 );
    or g828 ( n1007 , n1095 , n3043 );
    or g829 ( n160 , n3462 , n156 );
    not g830 ( n1917 , n2330 );
    not g831 ( n1112 , n1298 );
    and g832 ( n644 , n2519 , n1169 );
    not g833 ( n322 , n919 );
    not g834 ( n723 , n523 );
    not g835 ( n902 , n3786 );
    or g836 ( n3274 , n2010 , n2196 );
    and g837 ( n2702 , n826 , n3140 );
    or g838 ( n729 , n2797 , n2574 );
    nor g839 ( n593 , n1770 , n2238 );
    nor g840 ( n96 , n2950 , n2799 );
    nor g841 ( n434 , n2431 , n665 );
    or g842 ( n1512 , n2303 , n1385 );
    and g843 ( n3833 , n3740 , n590 );
    or g844 ( n765 , n3301 , n2683 );
    nor g845 ( n1116 , n2953 , n2547 );
    nor g846 ( n3563 , n314 , n1549 );
    or g847 ( n1078 , n2329 , n1305 );
    nor g848 ( n1095 , n1486 , n1799 );
    and g849 ( n1548 , n2889 , n3708 );
    nor g850 ( n2115 , n3826 , n2190 );
    and g851 ( n1874 , n873 , n3191 );
    or g852 ( n2456 , n3106 , n3765 );
    not g853 ( n3829 , n2482 );
    nor g854 ( n1958 , n2651 , n385 );
    or g855 ( n2722 , n3700 , n738 );
    nor g856 ( n85 , n1211 , n3090 );
    not g857 ( n1137 , n3578 );
    or g858 ( n99 , n3847 , n2175 );
    nor g859 ( n3267 , n304 , n2342 );
    not g860 ( n1094 , n2311 );
    and g861 ( n3061 , n2466 , n1224 );
    nor g862 ( n1207 , n2006 , n132 );
    nor g863 ( n1206 , n1308 , n300 );
    or g864 ( n3004 , n96 , n3078 );
    nor g865 ( n1671 , n2464 , n405 );
    or g866 ( n215 , n1195 , n3029 );
    or g867 ( n1794 , n3165 , n1128 );
    or g868 ( n706 , n2181 , n14 );
    or g869 ( n803 , n2608 , n2261 );
    and g870 ( n1184 , n1981 , n2315 );
    nor g871 ( n1683 , n1627 , n1792 );
    not g872 ( n710 , n615 );
    nor g873 ( n3830 , n1734 , n539 );
    or g874 ( n204 , n1170 , n859 );
    or g875 ( n1815 , n3119 , n1519 );
    or g876 ( n3816 , n3226 , n135 );
    nor g877 ( n1062 , n10 , n1603 );
    nor g878 ( n3382 , n1708 , n157 );
    nor g879 ( n825 , n809 , n1137 );
    nor g880 ( n3862 , n98 , n2498 );
    or g881 ( n1064 , n2161 , n222 );
    nor g882 ( n3794 , n920 , n3692 );
    nor g883 ( n2937 , n3502 , n3124 );
    not g884 ( n2614 , n1442 );
    or g885 ( n2710 , n724 , n480 );
    and g886 ( n642 , n3531 , n2322 );
    and g887 ( n1054 , n2521 , n1846 );
    nor g888 ( n2772 , n3695 , n3443 );
    or g889 ( n833 , n319 , n2409 );
    nor g890 ( n555 , n694 , n157 );
    nor g891 ( n786 , n3761 , n1533 );
    nor g892 ( n1286 , n2893 , n2190 );
    nor g893 ( n3851 , n553 , n281 );
    or g894 ( n2139 , n3551 , n1271 );
    nor g895 ( n2525 , n3604 , n1149 );
    or g896 ( n2627 , n3204 , n2332 );
    nor g897 ( n1730 , n2716 , n225 );
    or g898 ( n951 , n1584 , n1126 );
    nor g899 ( n3752 , n728 , n2132 );
    and g900 ( n2652 , n1778 , n3217 );
    nor g901 ( n397 , n3517 , n991 );
    and g902 ( n2215 , n2803 , n3077 );
    nor g903 ( n1119 , n3393 , n1597 );
    nor g904 ( n623 , n2025 , n1624 );
    nor g905 ( n832 , n3504 , n157 );
    and g906 ( n2211 , n3484 , n2597 );
    nor g907 ( n3273 , n3136 , n2408 );
    and g908 ( n3130 , n3685 , n720 );
    and g909 ( n1442 , n983 , n1581 );
    not g910 ( n357 , n546 );
    nor g911 ( n1998 , n3351 , n2933 );
    or g912 ( n2334 , n2542 , n3382 );
    not g913 ( n3280 , n186 );
    not g914 ( n1357 , n3743 );
    not g915 ( n2472 , n753 );
    not g916 ( n1707 , n1584 );
    or g917 ( n891 , n2122 , n2655 );
    and g918 ( n423 , n3088 , n2278 );
    nor g919 ( n1183 , n618 , n2758 );
    and g920 ( n2239 , n3274 , n396 );
    or g921 ( n339 , n1333 , n443 );
    and g922 ( n3286 , n506 , n3190 );
    nor g923 ( n2998 , n121 , n1226 );
    or g924 ( n881 , n925 , n935 );
    nor g925 ( n2646 , n1558 , n114 );
    nor g926 ( n2518 , n1996 , n233 );
    nor g927 ( n1012 , n282 , n1507 );
    or g928 ( n2625 , n351 , n3353 );
    nor g929 ( n3403 , n3544 , n2298 );
    nor g930 ( n2868 , n3427 , n3524 );
    nor g931 ( n2358 , n1043 , n1662 );
    or g932 ( n1348 , n874 , n3703 );
    and g933 ( n1203 , n2017 , n3280 );
    and g934 ( n2300 , n1390 , n693 );
    or g935 ( n2979 , n675 , n530 );
    nor g936 ( n2938 , n1712 , n2629 );
    or g937 ( n2371 , n3264 , n185 );
    nor g938 ( n722 , n616 , n3018 );
    or g939 ( n1742 , n3147 , n3086 );
    nor g940 ( n3493 , n2179 , n300 );
    or g941 ( n1188 , n3245 , n3346 );
    or g942 ( n2780 , n2836 , n3249 );
    nor g943 ( n1493 , n1861 , n558 );
    or g944 ( n3781 , n3228 , n2151 );
    or g945 ( n2475 , n1938 , n2366 );
    not g946 ( n263 , n511 );
    and g947 ( n465 , n1043 , n1185 );
    nor g948 ( n570 , n927 , n3090 );
    not g949 ( n1895 , n1140 );
    nor g950 ( n925 , n3488 , n260 );
    and g951 ( n242 , n880 , n1814 );
    or g952 ( n3163 , n3179 , n2262 );
    or g953 ( n976 , n2368 , n2188 );
    and g954 ( n2517 , n1807 , n2421 );
    nor g955 ( n548 , n2131 , n64 );
    not g956 ( n977 , n519 );
    nor g957 ( n2556 , n3473 , n159 );
    or g958 ( n774 , n3366 , n3101 );
    nor g959 ( n3046 , n2764 , n2775 );
    nor g960 ( n2981 , n332 , n1370 );
    or g961 ( n1171 , n2437 , n738 );
    or g962 ( n2093 , n2445 , n1126 );
    and g963 ( n2557 , n956 , n226 );
    nor g964 ( n569 , n2825 , n173 );
    or g965 ( n1932 , n386 , n1085 );
    not g966 ( n3070 , n2647 );
    nor g967 ( n695 , n673 , n2044 );
    nor g968 ( n1935 , n3684 , n640 );
    not g969 ( n3805 , n2776 );
    or g970 ( n1293 , n2672 , n2310 );
    or g971 ( n2307 , n2798 , n2830 );
    and g972 ( n2560 , n2789 , n3445 );
    nor g973 ( n1621 , n442 , n1880 );
    or g974 ( n1323 , n3557 , n1915 );
    nor g975 ( n2856 , n2676 , n3598 );
    and g976 ( n3542 , n561 , n3634 );
    nor g977 ( n2302 , n3207 , n620 );
    nor g978 ( n1181 , n3214 , n814 );
    nor g979 ( n3264 , n1622 , n68 );
    nor g980 ( n315 , n2251 , n5 );
    or g981 ( n3769 , n2644 , n2532 );
    or g982 ( n2107 , n2522 , n1214 );
    not g983 ( n1741 , n130 );
    not g984 ( n3632 , n1393 );
    nor g985 ( n2406 , n732 , n2822 );
    nor g986 ( n3764 , n1076 , n2241 );
    and g987 ( n988 , n2675 , n1987 );
    nor g988 ( n1528 , n2987 , n2868 );
    or g989 ( n1039 , n1549 , n1895 );
    and g990 ( n3720 , n1246 , n300 );
    not g991 ( n1238 , n1622 );
    or g992 ( n1876 , n430 , n1929 );
    nor g993 ( n1533 , n2814 , n3797 );
    or g994 ( n1332 , n1480 , n1079 );
    or g995 ( n1422 , n1982 , n3749 );
    nor g996 ( n2892 , n1893 , n261 );
    or g997 ( n3195 , n2003 , n777 );
    or g998 ( n2496 , n3218 , n859 );
    or g999 ( n2814 , n1502 , n2653 );
    and g1000 ( n1164 , n3451 , n2537 );
    and g1001 ( n445 , n1982 , n2459 );
    nor g1002 ( n1328 , n2309 , n3481 );
    nor g1003 ( n3519 , n2957 , n3721 );
    and g1004 ( n3197 , n3692 , n535 );
    or g1005 ( n715 , n2146 , n1263 );
    not g1006 ( n1175 , n1842 );
    and g1007 ( n316 , n2493 , n2992 );
    or g1008 ( n1233 , n1427 , n1263 );
    or g1009 ( n2353 , n3024 , n3746 );
    or g1010 ( n900 , n745 , n1365 );
    not g1011 ( n3370 , n3186 );
    nor g1012 ( n3107 , n3607 , n68 );
    nor g1013 ( n100 , n1437 , n1446 );
    and g1014 ( n2966 , n1989 , n172 );
    not g1015 ( n2841 , n2758 );
    nor g1016 ( n2906 , n687 , n3468 );
    or g1017 ( n1561 , n3547 , n1474 );
    not g1018 ( n2532 , n959 );
    and g1019 ( n402 , n2183 , n2663 );
    or g1020 ( n3109 , n2335 , n2303 );
    nor g1021 ( n3857 , n1257 , n1730 );
    not g1022 ( n1859 , n1631 );
    or g1023 ( n2561 , n1364 , n2349 );
    or g1024 ( n1735 , n2187 , n859 );
    not g1025 ( n2881 , n1916 );
    nor g1026 ( n273 , n3495 , n975 );
    or g1027 ( n1748 , n2709 , n2007 );
    nor g1028 ( n2476 , n2084 , n1644 );
    and g1029 ( n297 , n88 , n371 );
    or g1030 ( n2069 , n1532 , n3133 );
    or g1031 ( n1922 , n997 , n48 );
    or g1032 ( n3048 , n2766 , n1038 );
    nor g1033 ( n658 , n1212 , n2676 );
    not g1034 ( n1355 , n652 );
    not g1035 ( n3746 , n1374 );
    and g1036 ( n3408 , n3571 , n2114 );
    nor g1037 ( n2007 , n2151 , n1537 );
    not g1038 ( n1478 , n3820 );
    nor g1039 ( n3666 , n123 , n713 );
    not g1040 ( n101 , n93 );
    or g1041 ( n2753 , n1789 , n2500 );
    or g1042 ( n2605 , n1955 , n1443 );
    or g1043 ( n2337 , n2118 , n2168 );
    or g1044 ( n2082 , n1916 , n3148 );
    nor g1045 ( n3745 , n856 , n3233 );
    not g1046 ( n318 , n827 );
    or g1047 ( n2692 , n3113 , n642 );
    nor g1048 ( n2237 , n1158 , n2117 );
    nor g1049 ( n3675 , n3819 , n68 );
    not g1050 ( n3144 , n1764 );
    and g1051 ( n15 , n2777 , n2148 );
    or g1052 ( n1952 , n1669 , n1878 );
    nor g1053 ( n1918 , n2459 , n1982 );
    not g1054 ( n417 , n3143 );
    and g1055 ( n613 , n602 , n586 );
    and g1056 ( n2403 , n161 , n2274 );
    or g1057 ( n27 , n1741 , n607 );
    not g1058 ( n2324 , n2950 );
    nor g1059 ( n2902 , n3576 , n3069 );
    nor g1060 ( n429 , n1913 , n3193 );
    or g1061 ( n1447 , n2752 , n1291 );
    and g1062 ( n3479 , n764 , n956 );
    not g1063 ( n3855 , n3586 );
    or g1064 ( n3511 , n1375 , n2313 );
    not g1065 ( n2280 , n2853 );
    and g1066 ( n819 , n2455 , n772 );
    not g1067 ( n1696 , n3585 );
    or g1068 ( n962 , n2570 , n301 );
    or g1069 ( n3243 , n3381 , n2687 );
    or g1070 ( n3322 , n2924 , n3288 );
    and g1071 ( n1503 , n54 , n2411 );
    and g1072 ( n184 , n2222 , n989 );
    nor g1073 ( n2436 , n557 , n1539 );
    or g1074 ( n505 , n862 , n3146 );
    and g1075 ( n1955 , n1382 , n3041 );
    or g1076 ( n3023 , n3046 , n3633 );
    and g1077 ( n1001 , n3522 , n3293 );
    or g1078 ( n2442 , n1391 , n3037 );
    and g1079 ( n3841 , n1549 , n314 );
    or g1080 ( n861 , n1783 , n465 );
    nor g1081 ( n583 , n303 , n786 );
    and g1082 ( n2815 , n1505 , n1852 );
    not g1083 ( n3533 , n1805 );
    or g1084 ( n1204 , n2666 , n689 );
    nor g1085 ( n3388 , n428 , n836 );
    nor g1086 ( n799 , n2305 , n326 );
    nor g1087 ( n3097 , n1081 , n1482 );
    nor g1088 ( n740 , n2400 , n1287 );
    not g1089 ( n1185 , n466 );
    or g1090 ( n643 , n331 , n2244 );
    or g1091 ( n2891 , n1312 , n2548 );
    or g1092 ( n648 , n455 , n43 );
    or g1093 ( n2350 , n492 , n3205 );
    nor g1094 ( n393 , n2577 , n3842 );
    nor g1095 ( n228 , n3424 , n291 );
    nor g1096 ( n122 , n2609 , n2633 );
    nor g1097 ( n1372 , n990 , n2601 );
    nor g1098 ( n1674 , n2759 , n1300 );
    or g1099 ( n2426 , n3505 , n793 );
    or g1100 ( n3201 , n1941 , n1878 );
    or g1101 ( n1241 , n1607 , n1184 );
    or g1102 ( n1398 , n2806 , n2200 );
    nor g1103 ( n617 , n2951 , n2114 );
    nor g1104 ( n285 , n2158 , n886 );
    or g1105 ( n1224 , n208 , n1798 );
    nor g1106 ( n129 , n3314 , n533 );
    nor g1107 ( n3603 , n2809 , n1392 );
    and g1108 ( n2308 , n1873 , n2967 );
    or g1109 ( n3066 , n3060 , n2532 );
    nor g1110 ( n1271 , n1363 , n2575 );
    or g1111 ( n3164 , n2796 , n3246 );
    or g1112 ( n864 , n429 , n794 );
    nor g1113 ( n398 , n46 , n95 );
    or g1114 ( n113 , n256 , n2532 );
    nor g1115 ( n2416 , n3401 , n1673 );
    or g1116 ( n1166 , n3288 , n1126 );
    and g1117 ( n2923 , n3361 , n3559 );
    nor g1118 ( n2650 , n3410 , n192 );
    nor g1119 ( n2130 , n3561 , n3343 );
    or g1120 ( n3158 , n2866 , n2418 );
    nor g1121 ( n3152 , n1551 , n2520 );
    not g1122 ( n3749 , n1140 );
    or g1123 ( n2939 , n1924 , n2524 );
    nor g1124 ( n3753 , n1020 , n143 );
    and g1125 ( n3738 , n3026 , n1035 );
    nor g1126 ( n3258 , n1627 , n1537 );
    not g1127 ( n2911 , n2393 );
    nor g1128 ( n2528 , n2138 , n300 );
    and g1129 ( n3202 , n2355 , n87 );
    or g1130 ( n3181 , n965 , n1778 );
    or g1131 ( n241 , n502 , n3840 );
    nor g1132 ( n1280 , n3377 , n1137 );
    and g1133 ( n1527 , n2020 , n1494 );
    or g1134 ( n1031 , n149 , n1022 );
    and g1135 ( n1593 , n1191 , n2597 );
    and g1136 ( n399 , n2623 , n982 );
    not g1137 ( n1473 , n43 );
    or g1138 ( n528 , n2436 , n3239 );
    not g1139 ( n3717 , n1232 );
    nor g1140 ( n2389 , n1979 , n3266 );
    or g1141 ( n1863 , n2039 , n363 );
    or g1142 ( n3472 , n1048 , n2669 );
    or g1143 ( n597 , n249 , n1717 );
    nor g1144 ( n3078 , n3373 , n1537 );
    nor g1145 ( n118 , n2763 , n1281 );
    or g1146 ( n612 , n3586 , n1985 );
    or g1147 ( n563 , n797 , n2981 );
    nor g1148 ( n2910 , n579 , n2063 );
    or g1149 ( n2148 , n1963 , n3773 );
    nor g1150 ( n634 , n2536 , n2392 );
    and g1151 ( n3395 , n321 , n1241 );
    and g1152 ( n1377 , n1155 , n3805 );
    nor g1153 ( n1319 , n2858 , n246 );
    nor g1154 ( n418 , n1426 , n1564 );
    or g1155 ( n1004 , n3449 , n1810 );
    or g1156 ( n1182 , n3132 , n1407 );
    nor g1157 ( n1325 , n568 , n703 );
    or g1158 ( n1699 , n3639 , n1263 );
    and g1159 ( n3604 , n1051 , n3499 );
    or g1160 ( n471 , n320 , n3395 );
    or g1161 ( n1434 , n85 , n2257 );
    or g1162 ( n1648 , n16 , n2181 );
    or g1163 ( n1466 , n36 , n3827 );
    and g1164 ( n1246 , n2583 , n1130 );
    or g1165 ( n3644 , n3812 , n142 );
    and g1166 ( n3647 , n1589 , n1545 );
    nor g1167 ( n3686 , n863 , n444 );
    or g1168 ( n379 , n2325 , n1895 );
    nor g1169 ( n3399 , n3480 , n136 );
    nor g1170 ( n255 , n2882 , n358 );
    nor g1171 ( n2818 , n3035 , n2633 );
    nor g1172 ( n3175 , n366 , n2150 );
    and g1173 ( n3428 , n1388 , n2757 );
    and g1174 ( n1663 , n2136 , n1594 );
    not g1175 ( n1798 , n2665 );
    nor g1176 ( n1136 , n2795 , n3052 );
    nor g1177 ( n80 , n1437 , n936 );
    or g1178 ( n2539 , n1816 , n2460 );
    not g1179 ( n2212 , n1454 );
    or g1180 ( n693 , n1196 , n834 );
    or g1181 ( n2367 , n2080 , n547 );
    nor g1182 ( n2267 , n3345 , n2505 );
    and g1183 ( n1147 , n3130 , n2757 );
    or g1184 ( n3256 , n2547 , n1484 );
    or g1185 ( n2119 , n3458 , n3497 );
    not g1186 ( n509 , n2578 );
    or g1187 ( n996 , n2432 , n1818 );
    nor g1188 ( n1571 , n2719 , n1528 );
    or g1189 ( n2882 , n1280 , n1935 );
    not g1190 ( n789 , n1722 );
    nor g1191 ( n2679 , n3504 , n1556 );
    nor g1192 ( n2284 , n1343 , n1225 );
    not g1193 ( n2059 , n146 );
    nor g1194 ( n1463 , n2551 , n692 );
    not g1195 ( n1515 , n1211 );
    and g1196 ( n3022 , n45 , n2746 );
    nor g1197 ( n1688 , n2191 , n136 );
    and g1198 ( n1252 , n1038 , n3803 );
    and g1199 ( n3600 , n528 , n639 );
    or g1200 ( n3272 , n354 , n2808 );
    nor g1201 ( n3788 , n427 , n804 );
    nor g1202 ( n1047 , n966 , n1537 );
    or g1203 ( n1617 , n3848 , n3148 );
    or g1204 ( n3662 , n62 , n3276 );
    not g1205 ( n2099 , n1390 );
    not g1206 ( n3372 , n700 );
    or g1207 ( n1897 , n260 , n1798 );
    or g1208 ( n334 , n1074 , n859 );
    or g1209 ( n425 , n1027 , n3639 );
    or g1210 ( n470 , n1911 , n106 );
    nor g1211 ( n1100 , n3541 , n665 );
    not g1212 ( n2794 , n103 );
    or g1213 ( n1107 , n1702 , n3749 );
    nor g1214 ( n797 , n3784 , n718 );
    nor g1215 ( n3413 , n3861 , n878 );
    or g1216 ( n3089 , n1947 , n3346 );
    nor g1217 ( n3008 , n3021 , n1977 );
    or g1218 ( n3473 , n216 , n3512 );
    nor g1219 ( n1509 , n3153 , n2649 );
    or g1220 ( n1329 , n1847 , n970 );
    or g1221 ( n3017 , n491 , n2127 );
    and g1222 ( n2468 , n1638 , n1457 );
    nor g1223 ( n3615 , n800 , n2646 );
    or g1224 ( n2290 , n2745 , n1554 );
    or g1225 ( n1436 , n1146 , n3002 );
    or g1226 ( n1599 , n912 , n3482 );
    nor g1227 ( n1304 , n2541 , n1838 );
    not g1228 ( n2248 , n390 );
    and g1229 ( n513 , n2781 , n1500 );
    or g1230 ( n2715 , n2840 , n948 );
    or g1231 ( n1082 , n1835 , n1035 );
    nor g1232 ( n3589 , n1403 , n516 );
    not g1233 ( n674 , n3732 );
    or g1234 ( n2157 , n3738 , n3095 );
    not g1235 ( n1537 , n2656 );
    and g1236 ( n2631 , n2369 , n150 );
    or g1237 ( n2925 , n2297 , n3765 );
    nor g1238 ( n2072 , n2180 , n669 );
    nor g1239 ( n3147 , n383 , n2474 );
    nor g1240 ( n1607 , n104 , n850 );
    nor g1241 ( n2885 , n1338 , n324 );
    nor g1242 ( n461 , n3435 , n3859 );
    or g1243 ( n1758 , n3669 , n3812 );
    or g1244 ( n3172 , n990 , n3749 );
    nor g1245 ( n1995 , n607 , n2708 );
    not g1246 ( n1979 , n1877 );
    not g1247 ( n1235 , n2665 );
    not g1248 ( n3376 , n1574 );
    nor g1249 ( n3638 , n773 , n3583 );
    and g1250 ( n281 , n2266 , n3234 );
    and g1251 ( n1128 , n2547 , n2953 );
    or g1252 ( n1906 , n595 , n3134 );
    or g1253 ( n3824 , n2019 , n2133 );
    or g1254 ( n1386 , n553 , n2443 );
    or g1255 ( n3319 , n734 , n3403 );
    nor g1256 ( n3620 , n2753 , n2940 );
    not g1257 ( n2953 , n169 );
    nor g1258 ( n2258 , n1926 , n3368 );
    not g1259 ( n3379 , n2843 );
    or g1260 ( n890 , n3596 , n2435 );
    and g1261 ( n1242 , n2489 , n2087 );
    and g1262 ( n1771 , n3442 , n1176 );
    nor g1263 ( n108 , n2104 , n308 );
    not g1264 ( n2663 , n958 );
    or g1265 ( n718 , n3529 , n721 );
    nor g1266 ( n420 , n3319 , n2824 );
    or g1267 ( n3584 , n215 , n139 );
    not g1268 ( n3741 , n1654 );
    nor g1269 ( n2164 , n495 , n2772 );
    or g1270 ( n725 , n3754 , n3665 );
    nor g1271 ( n657 , n3794 , n100 );
    nor g1272 ( n3173 , n783 , n691 );
    nor g1273 ( n2080 , n2973 , n3143 );
    and g1274 ( n980 , n2676 , n1212 );
    or g1275 ( n3623 , n2663 , n3446 );
    nor g1276 ( n3492 , n2096 , n2298 );
    or g1277 ( n1543 , n1706 , n527 );
    nor g1278 ( n3030 , n1141 , n1037 );
    not g1279 ( n2817 , n1817 );
    not g1280 ( n911 , n3656 );
    nor g1281 ( n877 , n3850 , n3829 );
    and g1282 ( n2051 , n3383 , n1151 );
    or g1283 ( n1424 , n3744 , n1122 );
    nor g1284 ( n1752 , n2701 , n3666 );
    or g1285 ( n1462 , n551 , n2782 );
    not g1286 ( n3486 , n1601 );
    nor g1287 ( n3104 , n1559 , n2190 );
    nor g1288 ( n2010 , n221 , n2799 );
    nor g1289 ( n2706 , n1281 , n1977 );
    nor g1290 ( n970 , n900 , n1261 );
    and g1291 ( n986 , n2118 , n3165 );
    and g1292 ( n240 , n3438 , n322 );
    nor g1293 ( n107 , n1737 , n1527 );
    not g1294 ( n76 , n1281 );
    nor g1295 ( n1538 , n729 , n749 );
    nor g1296 ( n3467 , n667 , n1302 );
    and g1297 ( n2404 , n1250 , n818 );
    nor g1298 ( n1665 , n1600 , n2606 );
    and g1299 ( n1778 , n1150 , n2535 );
    nor g1300 ( n2901 , n1312 , n3169 );
    or g1301 ( n1401 , n3281 , n1045 );
    or g1302 ( n1347 , n2744 , n3434 );
    not g1303 ( n1545 , n1686 );
    or g1304 ( n2964 , n2929 , n1484 );
    nor g1305 ( n3184 , n2544 , n1537 );
    or g1306 ( n629 , n2770 , n250 );
    and g1307 ( n792 , n3691 , n772 );
    and g1308 ( n2038 , n2740 , n2381 );
    or g1309 ( n3809 , n2684 , n2935 );
    nor g1310 ( n451 , n2915 , n611 );
    or g1311 ( n3608 , n3328 , n163 );
    nor g1312 ( n697 , n1207 , n1113 );
    and g1313 ( n2567 , n431 , n3390 );
    nor g1314 ( n1379 , n2430 , n1752 );
    nor g1315 ( n2637 , n1364 , n3521 );
    nor g1316 ( n115 , n1874 , n92 );
    nor g1317 ( n1380 , n578 , n1673 );
    nor g1318 ( n1583 , n698 , n1758 );
    and g1319 ( n1891 , n817 , n612 );
    nor g1320 ( n2125 , n1032 , n1395 );
    or g1321 ( n3224 , n2153 , n3192 );
    and g1322 ( n3481 , n1468 , n334 );
    and g1323 ( n2878 , n1748 , n3438 );
    or g1324 ( n1656 , n3287 , n1235 );
    or g1325 ( n3252 , n1185 , n1783 );
    not g1326 ( n195 , n932 );
    and g1327 ( n3142 , n2309 , n3481 );
    not g1328 ( n3505 , n1738 );
    or g1329 ( n2623 , n3291 , n2687 );
    or g1330 ( n168 , n2202 , n3230 );
    or g1331 ( n488 , n1229 , n2067 );
    nor g1332 ( n1779 , n2909 , n1635 );
    not g1333 ( n497 , n3381 );
    not g1334 ( n2482 , n700 );
    not g1335 ( n663 , n1825 );
    or g1336 ( n1149 , n1809 , n2403 );
    and g1337 ( n1928 , n1237 , n1000 );
    not g1338 ( n1659 , n3626 );
    or g1339 ( n537 , n3067 , n1797 );
    and g1340 ( n906 , n3195 , n3055 );
    and g1341 ( n949 , n3299 , n3220 );
    nor g1342 ( n3270 , n362 , n2633 );
    or g1343 ( n600 , n3225 , n213 );
    and g1344 ( n2127 , n923 , n3559 );
    nor g1345 ( n1406 , n2330 , n2799 );
    nor g1346 ( n1757 , n2140 , n813 );
    or g1347 ( n1117 , n3196 , n3528 );
    or g1348 ( n835 , n1441 , n3020 );
    and g1349 ( n793 , n836 , n428 );
    nor g1350 ( n2529 , n3718 , n157 );
    and g1351 ( n1635 , n550 , n2197 );
    or g1352 ( n1718 , n824 , n240 );
    or g1353 ( n2065 , n82 , n2211 );
    or g1354 ( n2575 , n2639 , n520 );
    and g1355 ( n2454 , n1018 , n2421 );
    and g1356 ( n1084 , n2032 , n691 );
    and g1357 ( n3497 , n159 , n936 );
    nor g1358 ( n3448 , n2563 , n273 );
    not g1359 ( n1161 , n1524 );
    or g1360 ( n2703 , n309 , n660 );
    or g1361 ( n401 , n3335 , n1929 );
    nor g1362 ( n2852 , n2680 , n2108 );
    nor g1363 ( n3427 , n736 , n3035 );
    nor g1364 ( n2074 , n2530 , n2704 );
    and g1365 ( n203 , n1308 , n3771 );
    or g1366 ( n385 , n66 , n3179 );
    nor g1367 ( n1023 , n1933 , n774 );
    or g1368 ( n3532 , n2854 , n3408 );
    or g1369 ( n3658 , n1474 , n2168 );
    and g1370 ( n1881 , n3730 , n3116 );
    and g1371 ( n1092 , n2031 , n1129 );
    not g1372 ( n383 , n2090 );
    nor g1373 ( n737 , n485 , n3024 );
    or g1374 ( n915 , n350 , n2035 );
    nor g1375 ( n2230 , n1563 , n3417 );
    nor g1376 ( n2247 , n2712 , n1302 );
    and g1377 ( n1352 , n3007 , n493 );
    or g1378 ( n2768 , n2992 , n3344 );
    nor g1379 ( n1576 , n1024 , n722 );
    nor g1380 ( n2409 , n577 , n3593 );
    and g1381 ( n2287 , n3637 , n3627 );
    nor g1382 ( n3098 , n474 , n2708 );
    nor g1383 ( n1516 , n2401 , n1186 );
    and g1384 ( n2988 , n525 , n3741 );
    nor g1385 ( n775 , n2848 , n3217 );
    and g1386 ( n472 , n1247 , n2802 );
    nor g1387 ( n3580 , n1681 , n2094 );
    nor g1388 ( n2500 , n2142 , n3742 );
    and g1389 ( n3298 , n782 , n3032 );
    not g1390 ( n679 , n349 );
    and g1391 ( n3605 , n70 , n1603 );
    or g1392 ( n3016 , n83 , n3679 );
    and g1393 ( n58 , n3681 , n136 );
    not g1394 ( n1539 , n1295 );
    not g1395 ( n2699 , n2321 );
    or g1396 ( n3734 , n1050 , n147 );
    nor g1397 ( n3369 , n3332 , n221 );
    not g1398 ( n3087 , n3377 );
    or g1399 ( n2376 , n2027 , n1235 );
    nor g1400 ( n2534 , n3004 , n300 );
    nor g1401 ( n2213 , n694 , n1462 );
    not g1402 ( n1258 , n3808 );
    not g1403 ( n2413 , n2169 );
    nor g1404 ( n3420 , n2491 , n3770 );
    or g1405 ( n2796 , n3549 , n2892 );
    and g1406 ( n1030 , n1111 , n3111 );
    and g1407 ( n1446 , n2165 , n3251 );
    not g1408 ( n2809 , n1315 );
    nor g1409 ( n1063 , n3831 , n3541 );
    and g1410 ( n3790 , n1169 , n3032 );
    not g1411 ( n595 , n964 );
    and g1412 ( n3155 , n2223 , n2597 );
    not g1413 ( n3553 , n726 );
    nor g1414 ( n1087 , n203 , n3118 );
    nor g1415 ( n3099 , n2022 , n2471 );
    and g1416 ( n2441 , n2838 , n2370 );
    nor g1417 ( n59 , n3730 , n3116 );
    and g1418 ( n2018 , n3698 , n3379 );
    and g1419 ( n1689 , n1653 , n1019 );
    nor g1420 ( n3750 , n2400 , n3032 );
    or g1421 ( n448 , n2761 , n1985 );
    nor g1422 ( n233 , n3688 , n1577 );
    nor g1423 ( n225 , n589 , n1693 );
    nor g1424 ( n1880 , n1089 , n3661 );
    or g1425 ( n3561 , n1093 , n3162 );
    not g1426 ( n2696 , n3432 );
    or g1427 ( n3657 , n86 , n2462 );
    nor g1428 ( n2271 , n3079 , n183 );
    nor g1429 ( n23 , n2685 , n848 );
    or g1430 ( n3457 , n638 , n2399 );
    not g1431 ( n614 , n1002 );
    not g1432 ( n1722 , n2413 );
    or g1433 ( n3778 , n1277 , n2276 );
    not g1434 ( n2359 , n3755 );
    or g1435 ( n1127 , n1255 , n2896 );
    not g1436 ( n2019 , n430 );
    or g1437 ( n3055 , n1323 , n1178 );
    or g1438 ( n784 , n1557 , n3752 );
    not g1439 ( n3148 , n1722 );
    or g1440 ( n1297 , n825 , n1560 );
    and g1441 ( n2338 , n1715 , n583 );
    not g1442 ( n2747 , n1276 );
    nor g1443 ( n979 , n483 , n866 );
    and g1444 ( n2653 , n3269 , n292 );
    not g1445 ( n2595 , n3372 );
    not g1446 ( n3461 , n3758 );
    or g1447 ( n3383 , n1700 , n3601 );
    not g1448 ( n2786 , n1825 );
    nor g1449 ( n2380 , n529 , n1877 );
    or g1450 ( n469 , n3385 , n1126 );
    or g1451 ( n892 , n1927 , n3402 );
    or g1452 ( n2612 , n2842 , n3490 );
    not g1453 ( n3079 , n1680 );
    or g1454 ( n2541 , n2969 , n1930 );
    not g1455 ( n3207 , n260 );
    nor g1456 ( n1506 , n961 , n84 );
    nor g1457 ( n2134 , n1112 , n3186 );
    or g1458 ( n1134 , n2130 , n2128 );
    and g1459 ( n1061 , n132 , n2006 );
    nor g1460 ( n356 , n2355 , n936 );
    not g1461 ( n2996 , n2745 );
    not g1462 ( n2607 , n2187 );
    or g1463 ( n3715 , n916 , n701 );
    nor g1464 ( n3618 , n283 , n1423 );
    nor g1465 ( n987 , n2817 , n229 );
    not g1466 ( n3634 , n927 );
    or g1467 ( n1426 , n1010 , n3851 );
    nor g1468 ( n320 , n2599 , n1669 );
    or g1469 ( n3860 , n632 , n1335 );
    or g1470 ( n1165 , n2193 , n3527 );
    or g1471 ( n170 , n395 , n2105 );
    and g1472 ( n3051 , n3722 , n717 );
    and g1473 ( n875 , n2195 , n2093 );
    and g1474 ( n310 , n2785 , n898 );
    or g1475 ( n439 , n652 , n2921 );
    or g1476 ( n3212 , n751 , n3665 );
    nor g1477 ( n1892 , n161 , n730 );
    and g1478 ( n2418 , n1755 , n2087 );
    and g1479 ( n2918 , n1865 , n3224 );
    and g1480 ( n2688 , n588 , n1781 );
    nor g1481 ( n3400 , n3649 , n3640 );
    or g1482 ( n2438 , n1136 , n3838 );
    and g1483 ( n669 , n3736 , n241 );
    or g1484 ( n2863 , n2483 , n1483 );
    not g1485 ( n3241 , n3625 );
    not g1486 ( n2366 , n972 );
    and g1487 ( n14 , n16 , n3567 );
    and g1488 ( n3571 , n562 , n166 );
    and g1489 ( n2629 , n477 , n2618 );
    or g1490 ( n2664 , n2875 , n3275 );
    and g1491 ( n1086 , n183 , n3079 );
    nor g1492 ( n2487 , n408 , n3267 );
    nor g1493 ( n1274 , n3052 , n814 );
    nor g1494 ( n3371 , n783 , n2032 );
    not g1495 ( n2274 , n2079 );
    not g1496 ( n1710 , n1322 );
    nor g1497 ( n2485 , n1103 , n852 );
    and g1498 ( n735 , n1559 , n2877 );
    nor g1499 ( n2288 , n2172 , n399 );
    or g1500 ( n308 , n3811 , n556 );
    and g1501 ( n2562 , n895 , n2116 );
    nor g1502 ( n1225 , n2225 , n1304 );
    not g1503 ( n3138 , n2752 );
    nor g1504 ( n2241 , n597 , n867 );
    or g1505 ( n2345 , n1472 , n776 );
    not g1506 ( n1216 , n1099 );
    or g1507 ( n1284 , n3391 , n1711 );
    nor g1508 ( n2037 , n1145 , n577 );
    or g1509 ( n2344 , n3562 , n205 );
    and g1510 ( n2062 , n966 , n2875 );
    not g1511 ( n342 , n362 );
    nor g1512 ( n1882 , n558 , n95 );
    nor g1513 ( n2250 , n2221 , n2004 );
    and g1514 ( n1711 , n1162 , n2824 );
    or g1515 ( n464 , n229 , n1085 );
    and g1516 ( n721 , n1392 , n2809 );
    or g1517 ( n291 , n1481 , n2942 );
    and g1518 ( n2219 , n3552 , n1646 );
    nor g1519 ( n3121 , n2268 , n1753 );
    not g1520 ( n2936 , n2662 );
    nor g1521 ( n2045 , n3033 , n3448 );
    nor g1522 ( n2295 , n90 , n1134 );
    nor g1523 ( n1208 , n3808 , n1662 );
    or g1524 ( n1511 , n3698 , n1085 );
    and g1525 ( n956 , n188 , n1910 );
    or g1526 ( n2450 , n1317 , n1548 );
    nor g1527 ( n768 , n1308 , n3771 );
    and g1528 ( n1845 , n126 , n2713 );
    not g1529 ( n3583 , n1295 );
    nor g1530 ( n3208 , n3420 , n1340 );
    nor g1531 ( n2917 , n2453 , n2595 );
    or g1532 ( n2023 , n1703 , n1049 );
    and g1533 ( n3034 , n639 , n2114 );
    nor g1534 ( n624 , n2254 , n1975 );
    nor g1535 ( n3798 , n1254 , n2799 );
    and g1536 ( n3254 , n167 , n2053 );
    and g1537 ( n1914 , n242 , n1114 );
    or g1538 ( n1364 , n193 , n1572 );
    nor g1539 ( n898 , n13 , n2377 );
    not g1540 ( n636 , n990 );
    nor g1541 ( n3455 , n2112 , n847 );
    nor g1542 ( n2024 , n3400 , n1102 );
    and g1543 ( n1388 , n3560 , n1656 );
    nor g1544 ( n3057 , n2497 , n1683 );
    nor g1545 ( n3844 , n2899 , n1354 );
    and g1546 ( n1018 , n3599 , n279 );
    nor g1547 ( n1479 , n289 , n3805 );
    or g1548 ( n2920 , n3161 , n370 );
    and g1549 ( n3538 , n2946 , n1755 );
    or g1550 ( n1936 , n2362 , n3271 );
    and g1551 ( n1769 , n61 , n2367 );
    nor g1552 ( n3095 , n3774 , n228 );
    not g1553 ( n483 , n3672 );
    or g1554 ( n1713 , n668 , n654 );
    or g1555 ( n1432 , n1387 , n2215 );
    or g1556 ( n909 , n805 , n1455 );
    not g1557 ( n3782 , n2097 );
    nor g1558 ( n2108 , n2143 , n2561 );
    and g1559 ( n499 , n3641 , n2996 );
    and g1560 ( n2989 , n3393 , n1597 );
    and g1561 ( n3707 , n3784 , n3529 );
    and g1562 ( n1341 , n3565 , n1953 );
    not g1563 ( n309 , n2978 );
    or g1564 ( n171 , n1684 , n2382 );
    nor g1565 ( n2716 , n2226 , n1388 );
    or g1566 ( n1301 , n3816 , n1414 );
    or g1567 ( n3617 , n634 , n1518 );
    not g1568 ( n3293 , n1467 );
    or g1569 ( n3139 , n3006 , n42 );
    and g1570 ( n7 , n3404 , n1341 );
    nor g1571 ( n2771 , n891 , n2447 );
    nor g1572 ( n3419 , n101 , n1141 );
    nor g1573 ( n3811 , n2324 , n3373 );
    nor g1574 ( n3534 , n2222 , n989 );
    not g1575 ( n726 , n700 );
    nor g1576 ( n2081 , n692 , n2874 );
    nor g1577 ( n2259 , n931 , n2298 );
    nor g1578 ( n2608 , n2853 , n1539 );
    and g1579 ( n2723 , n3649 , n3640 );
    or g1580 ( n2970 , n1800 , n3241 );
    or g1581 ( n1260 , n2856 , n1006 );
    nor g1582 ( n2348 , n1905 , n2787 );
    nor g1583 ( n3240 , n1146 , n64 );
    not g1584 ( n3228 , n2328 );
    not g1585 ( n2632 , n1596 );
    and g1586 ( n1694 , n694 , n551 );
    nor g1587 ( n3389 , n3038 , n2092 );
    nor g1588 ( n3459 , n3785 , n1072 );
    and g1589 ( n3506 , n354 , n2808 );
    or g1590 ( n1412 , n128 , n1588 );
    nor g1591 ( n703 , n413 , n3657 );
    not g1592 ( n2459 , n1427 );
    and g1593 ( n2846 , n2893 , n1917 );
    nor g1594 ( n2871 , n1671 , n1670 );
    nor g1595 ( n1088 , n3568 , n1937 );
    and g1596 ( n2927 , n2808 , n3077 );
    or g1597 ( n378 , n2669 , n1023 );
    and g1598 ( n3771 , n1065 , n1052 );
    or g1599 ( n2626 , n186 , n2105 );
    nor g1600 ( n3180 , n624 , n3453 );
    or g1601 ( n1992 , n289 , n978 );
    or g1602 ( n3126 , n1448 , n789 );
    nor g1603 ( n1706 , n215 , n2757 );
    nor g1604 ( n2446 , n822 , n2579 );
    nor g1605 ( n3132 , n1034 , n1495 );
    nor g1606 ( n3536 , n3834 , n1276 );
    not g1607 ( n1803 , n1217 );
    nor g1608 ( n709 , n239 , n2824 );
    not g1609 ( n1391 , n1476 );
    nor g1610 ( n1460 , n3144 , n3367 );
    not g1611 ( n3153 , n1314 );
    nor g1612 ( n2704 , n3821 , n49 );
    or g1613 ( n739 , n3436 , n1895 );
    not g1614 ( n3574 , n432 );
    not g1615 ( n2329 , n2635 );
    not g1616 ( n3592 , n1825 );
    or g1617 ( n2947 , n1806 , n3765 );
    or g1618 ( n3736 , n3673 , n2687 );
    nor g1619 ( n858 , n1351 , n619 );
    not g1620 ( n3832 , n1578 );
    nor g1621 ( n522 , n2222 , n136 );
    and g1622 ( n1201 , n763 , n3361 );
    nor g1623 ( n189 , n731 , n2012 );
    nor g1624 ( n1470 , n441 , n665 );
    or g1625 ( n3072 , n2900 , n1262 );
    or g1626 ( n1228 , n2492 , n17 );
    not g1627 ( n3739 , n2439 );
    or g1628 ( n2425 , n3581 , n1773 );
    and g1629 ( n1850 , n2277 , n3127 );
    not g1630 ( n704 , n1804 );
    nor g1631 ( n3757 , n3843 , n95 );
    not g1632 ( n2025 , n1582 );
    or g1633 ( n1005 , n1720 , n1126 );
    nor g1634 ( n3253 , n3491 , n2343 );
    nor g1635 ( n3105 , n3822 , n3583 );
    not g1636 ( n1085 , n3049 );
    or g1637 ( n3350 , n2506 , n1641 );
    and g1638 ( n1287 , n1233 , n1422 );
    or g1639 ( n153 , n131 , n1593 );
    nor g1640 ( n3622 , n1727 , n299 );
    or g1641 ( n1961 , n3379 , n445 );
    nor g1642 ( n1715 , n1875 , n2939 );
    and g1643 ( n2821 , n803 , n1689 );
    and g1644 ( n1326 , n1623 , n342 );
    nor g1645 ( n149 , n404 , n1977 );
    and g1646 ( n3484 , n3194 , n951 );
    or g1647 ( n2184 , n1440 , n3681 );
    and g1648 ( n2166 , n625 , n3760 );
    or g1649 ( n3211 , n1841 , n2223 );
    or g1650 ( n188 , n3758 , n3746 );
    or g1651 ( n720 , n827 , n1385 );
    or g1652 ( n234 , n2721 , n2687 );
    or g1653 ( n2713 , n2890 , n1895 );
    nor g1654 ( n3791 , n2944 , n3261 );
    not g1655 ( n157 , n1766 );
    and g1656 ( n2382 , n883 , n2869 );
    and g1657 ( n3606 , n3300 , n1313 );
    nor g1658 ( n3482 , n1950 , n3593 );
    nor g1659 ( n1997 , n2384 , n2752 );
    not g1660 ( n3362 , n981 );
    or g1661 ( n937 , n292 , n1502 );
    or g1662 ( n2533 , n3190 , n1270 );
    or g1663 ( n274 , n626 , n2815 );
    nor g1664 ( n2683 , n1359 , n2958 );
    or g1665 ( n3799 , n123 , n3840 );
    nor g1666 ( n1033 , n3125 , n640 );
    and g1667 ( n3042 , n670 , n1194 );
    nor g1668 ( n83 , n1411 , n2156 );
    and g1669 ( n3182 , n3116 , n150 );
    or g1670 ( n127 , n2841 , n1420 );
    or g1671 ( n67 , n3466 , n2760 );
    and g1672 ( n117 , n2531 , n772 );
    or g1673 ( n438 , n109 , n2168 );
    nor g1674 ( n1573 , n2882 , n2527 );
    not g1675 ( n759 , n246 );
    nor g1676 ( n1101 , n2622 , n1598 );
    nor g1677 ( n3150 , n683 , n2708 );
    nor g1678 ( n3445 , n1142 , n3518 );
    not g1679 ( n2967 , n1855 );
    not g1680 ( n1825 , n790 );
    and g1681 ( n33 , n1824 , n1114 );
    nor g1682 ( n2490 , n93 , n665 );
    not g1683 ( n1358 , n1448 );
    not g1684 ( n1960 , n2146 );
    nor g1685 ( n2615 , n3082 , n69 );
    or g1686 ( n1428 , n3410 , n3862 );
    or g1687 ( n1008 , n3275 , n3176 );
    not g1688 ( n806 , n1701 );
    not g1689 ( n3627 , n3607 );
    or g1690 ( n1303 , n40 , n2366 );
    nor g1691 ( n2177 , n174 , n2422 );
    or g1692 ( n844 , n3105 , n515 );
    or g1693 ( n289 , n601 , n1542 );
    or g1694 ( n41 , n489 , n35 );
    or g1695 ( n621 , n1888 , n380 );
    or g1696 ( n1013 , n277 , n1700 );
    and g1697 ( n971 , n3530 , n3614 );
    or g1698 ( n2582 , n2339 , n2168 );
    or g1699 ( n2586 , n3498 , n3346 );
    nor g1700 ( n2866 , n2946 , n143 );
    nor g1701 ( n2272 , n470 , n2064 );
    nor g1702 ( n1097 , n3513 , n1598 );
    nor g1703 ( n3246 , n564 , n1896 );
    and g1704 ( n687 , n467 , n3461 );
    nor g1705 ( n2270 , n3269 , n937 );
    nor g1706 ( n2914 , n1625 , n3489 );
    nor g1707 ( n2682 , n345 , n157 );
    nor g1708 ( n1438 , n3739 , n1454 );
    and g1709 ( n1964 , n2453 , n1824 );
    nor g1710 ( n702 , n1515 , n388 );
    not g1711 ( n2742 , n3125 );
    or g1712 ( n1444 , n1989 , n172 );
    nor g1713 ( n351 , n2001 , n2407 );
    nor g1714 ( n2060 , n706 , n765 );
    or g1715 ( n1987 , n259 , n2720 );
    or g1716 ( n1945 , n420 , n165 );
    or g1717 ( n910 , n1042 , n144 );
    nor g1718 ( n2462 , n3238 , n2050 );
    or g1719 ( n2316 , n1870 , n3732 );
    or g1720 ( n1749 , n1602 , n2740 );
    or g1721 ( n992 , n361 , n1263 );
    not g1722 ( n3840 , n3049 );
    nor g1723 ( n2552 , n2971 , n3598 );
    or g1724 ( n586 , n1294 , n1566 );
    nor g1725 ( n2823 , n2668 , n847 );
    or g1726 ( n2155 , n1817 , n789 );
    or g1727 ( n776 , n1486 , n3545 );
    not g1728 ( n226 , n3372 );
    nor g1729 ( n1218 , n1978 , n1817 );
    not g1730 ( n2049 , n700 );
    nor g1731 ( n2201 , n560 , n2799 );
    or g1732 ( n1848 , n2017 , n1484 );
    or g1733 ( n1413 , n1943 , n3710 );
    or g1734 ( n2314 , n835 , n242 );
    and g1735 ( n842 , n1187 , n3728 );
    and g1736 ( n3692 , n3476 , n214 );
    or g1737 ( n1923 , n261 , n3346 );
    and g1738 ( n3567 , n1617 , n771 );
    and g1739 ( n1096 , n1714 , n680 );
    or g1740 ( n2428 , n1075 , n1235 );
    and g1741 ( n1618 , n388 , n1515 );
    or g1742 ( n771 , n838 , n1385 );
    and g1743 ( n380 , n178 , n1230 );
    nor g1744 ( n1066 , n2494 , n3355 );
    or g1745 ( n8 , n2162 , n3605 );
    nor g1746 ( n953 , n2919 , n1907 );
    or g1747 ( n2499 , n110 , n1117 );
    nor g1748 ( n1192 , n2334 , n2051 );
    or g1749 ( n3268 , n1615 , n3840 );
    nor g1750 ( n2849 , n1535 , n3232 );
    and g1751 ( n338 , n3611 , n6 );
    or g1752 ( n2461 , n2510 , n2160 );
    nor g1753 ( n376 , n2210 , n769 );
    or g1754 ( n2340 , n2810 , n2507 );
    nor g1755 ( n2362 , n2031 , n691 );
    not g1756 ( n428 , n46 );
    nor g1757 ( n1261 , n3121 , n2144 );
    and g1758 ( n3406 , n1609 , n204 );
    or g1759 ( n3442 , n3825 , n1732 );
    nor g1760 ( n3020 , n2390 , n1698 );
    or g1761 ( n628 , n1644 , n2158 );
    nor g1762 ( n1153 , n348 , n3025 );
    or g1763 ( n3289 , n2932 , n1385 );
    not g1764 ( n3831 , n685 );
    not g1765 ( n2825 , n3498 );
    nor g1766 ( n3352 , n2191 , n2304 );
    nor g1767 ( n3347 , n1250 , n3069 );
    not g1768 ( n3842 , n1766 );
    not g1769 ( n3041 , n904 );
    and g1770 ( n2186 , n221 , n3332 );
    and g1771 ( n2073 , n2405 , n1175 );
    nor g1772 ( n761 , n672 , n2871 );
    or g1773 ( n1581 , n630 , n2393 );
    nor g1774 ( n3802 , n3628 , n55 );
    or g1775 ( n2630 , n1153 , n1469 );
    or g1776 ( n2634 , n729 , n549 );
    nor g1777 ( n945 , n1111 , n226 );
    nor g1778 ( n3660 , n1498 , n2592 );
    not g1779 ( n104 , n2076 );
    nor g1780 ( n1687 , n536 , n3555 );
    and g1781 ( n933 , n223 , n3141 );
    or g1782 ( n1076 , n7 , n2986 );
    or g1783 ( n3320 , n828 , n2451 );
    or g1784 ( n2686 , n1801 , n2045 );
    nor g1785 ( n2894 , n1297 , n2595 );
    nor g1786 ( n2584 , n2758 , n2799 );
    nor g1787 ( n743 , n2189 , n395 );
    or g1788 ( n1199 , n1726 , n2200 );
    not g1789 ( n1579 , n841 );
    and g1790 ( n193 , n3054 , n3717 );
    not g1791 ( n3593 , n43 );
    nor g1792 ( n2792 , n22 , n3356 );
    nor g1793 ( n967 , n528 , n639 );
    or g1794 ( n409 , n1777 , n2571 );
    or g1795 ( n1180 , n1574 , n2687 );
    nor g1796 ( n599 , n3776 , n2633 );
    nor g1797 ( n1849 , n457 , n2724 );
    nor g1798 ( n2857 , n3157 , n3683 );
    or g1799 ( n426 , n265 , n3428 );
    and g1800 ( n3006 , n2191 , n2304 );
    nor g1801 ( n573 , n3340 , n2346 );
    and g1802 ( n1016 , n2218 , n719 );
    or g1803 ( n3045 , n709 , n3767 );
    not g1804 ( n1302 , n2248 );
    nor g1805 ( n1010 , n2881 , n462 );
    or g1806 ( n2171 , n1712 , n1516 );
    nor g1807 ( n3667 , n16 , n3829 );
    not g1808 ( n468 , n317 );
    not g1809 ( n2754 , n1708 );
    or g1810 ( n1841 , n3270 , n1677 );
    nor g1811 ( n3783 , n2847 , n3253 );
    and g1812 ( n639 , n3177 , n2058 );
    and g1813 ( n1129 , n1249 , n2428 );
    nor g1814 ( n750 , n2696 , n1965 );
    and g1815 ( n3549 , n173 , n2825 );
    or g1816 ( n883 , n3786 , n3746 );
    nor g1817 ( n2434 , n531 , n3348 );
    nor g1818 ( n3653 , n3544 , n3072 );
    not g1819 ( n2824 , n1190 );
    or g1820 ( n1437 , n451 , n3080 );
    nor g1821 ( n2261 , n1132 , n1662 );
    and g1822 ( n2028 , n1689 , n1114 );
    nor g1823 ( n3501 , n3733 , n681 );
    nor g1824 ( n638 , n870 , n2555 );
    not g1825 ( n3311 , n395 );
    or g1826 ( n2402 , n1262 , n2860 );
    and g1827 ( n3733 , n457 , n2724 );
    nor g1828 ( n2867 , n521 , n2473 );
    not g1829 ( n2243 , n3578 );
    or g1830 ( n1558 , n3423 , n2227 );
    nor g1831 ( n2709 , n2328 , n1137 );
    not g1832 ( n2985 , n700 );
    or g1833 ( n2379 , n3813 , n1026 );
    not g1834 ( n2678 , n3582 );
    nor g1835 ( n1770 , n1109 , n44 );
    and g1836 ( n1939 , n3044 , n1238 );
    or g1837 ( n1418 , n181 , n182 );
    or g1838 ( n2106 , n2037 , n310 );
    or g1839 ( n3368 , n1642 , n2805 );
    and g1840 ( n929 , n2872 , n330 );
    or g1841 ( n2117 , n3716 , n2338 );
    not g1842 ( n640 , n43 );
    nor g1843 ( n1098 , n232 , n1246 );
    and g1844 ( n3321 , n3463 , n650 );
    and g1845 ( n2733 , n2400 , n1287 );
    nor g1846 ( n2111 , n1850 , n72 );
    nor g1847 ( n90 , n3076 , n1657 );
    and g1848 ( n2744 , n1395 , n1032 );
    and g1849 ( n887 , n1346 , n286 );
    or g1850 ( n1751 , n137 , n2159 );
    and g1851 ( n159 , n1699 , n854 );
    and g1852 ( n172 , n3201 , n438 );
    nor g1853 ( n1725 , n1873 , n2026 );
    nor g1854 ( n296 , n238 , n3437 );
    nor g1855 ( n2036 , n1419 , n1664 );
    nor g1856 ( n1641 , n3687 , n954 );
    or g1857 ( n991 , n2750 , n651 );
    nor g1858 ( n102 , n1311 , n210 );
    nor g1859 ( n105 , n2594 , n376 );
    or g1860 ( n985 , n775 , n641 );
    not g1861 ( n2795 , n1015 );
    nor g1862 ( n2537 , n1823 , n1 );
    or g1863 ( n1052 , n2636 , n738 );
    not g1864 ( n1555 , n683 );
    nor g1865 ( n3569 , n1548 , n418 );
    and g1866 ( n889 , n1627 , n2936 );
    or g1867 ( n1307 , n356 , n1240 );
    nor g1868 ( n3063 , n1376 , n1539 );
    not g1869 ( n919 , n700 );
    or g1870 ( n802 , n546 , n2105 );
    and g1871 ( n2067 , n2216 , n2816 );
    or g1872 ( n1782 , n872 , n18 );
    or g1873 ( n1667 , n2747 , n1074 );
    nor g1874 ( n452 , n2097 , n3593 );
    or g1875 ( n407 , n3136 , n3360 );
    and g1876 ( n2057 , n19 , n791 );
    and g1877 ( n3521 , n604 , n3587 );
    not g1878 ( n2816 , n455 );
    nor g1879 ( n2762 , n2407 , n1537 );
    not g1880 ( n3708 , n1947 );
    or g1881 ( n2869 , n732 , n1385 );
    nor g1882 ( n2269 , n2026 , n1603 );
    nor g1883 ( n1637 , n2521 , n2026 );
    or g1884 ( n1445 , n2378 , n738 );
    nor g1885 ( n1871 , n50 , n3199 );
    nor g1886 ( n2471 , n2521 , n3483 );
    and g1887 ( n1566 , n1127 , n1697 );
    or g1888 ( n2206 , n2372 , n3790 );
    or g1889 ( n2491 , n2818 , n2823 );
    and g1890 ( n568 , n2544 , n1083 );
    not g1891 ( n1404 , n176 );
    or g1892 ( n2104 , n2998 , n3844 );
    or g1893 ( n856 , n3019 , n3102 );
    not g1894 ( n1554 , n1374 );
    nor g1895 ( n2876 , n1738 , n95 );
    and g1896 ( n1055 , n2179 , n3691 );
    not g1897 ( n2129 , n2520 );
    nor g1898 ( n1672 , n2253 , n1977 );
    nor g1899 ( n207 , n510 , n2615 );
    nor g1900 ( n3117 , n1957 , n921 );
    nor g1901 ( n2641 , n1555 , n3756 );
    or g1902 ( n477 , n3670 , n3432 );
    or g1903 ( n2905 , n1517 , n2318 );
    nor g1904 ( n78 , n860 , n189 );
    not g1905 ( n2764 , n3822 );
    not g1906 ( n1477 , n1483 );
    not g1907 ( n63 , n1495 );
    and g1908 ( n1865 , n2173 , n637 );
    not g1909 ( n2256 , n2417 );
    and g1910 ( n2133 , n3721 , n2957 );
    or g1911 ( n223 , n2584 , n2429 );
    nor g1912 ( n424 , n531 , n1072 );
    nor g1913 ( n654 , n1681 , n2688 );
    and g1914 ( n30 , n1440 , n3681 );
    or g1915 ( n1226 , n1458 , n2224 );
    not g1916 ( n231 , n574 );
    or g1917 ( n2031 , n1430 , n3492 );
    nor g1918 ( n3080 , n1371 , n814 );
    and g1919 ( n369 , n1243 , n1744 );
    and g1920 ( n2088 , n3092 , n3748 );
    nor g1921 ( n913 , n1245 , n3262 );
    nor g1922 ( n1823 , n493 , n3007 );
    not g1923 ( n2190 , n3374 );
    or g1924 ( n271 , n2845 , n218 );
    and g1925 ( n2524 , n3502 , n1776 );
    nor g1926 ( n1102 , n1771 , n3651 );
    or g1927 ( n728 , n3429 , n424 );
    nor g1928 ( n3231 , n3041 , n1382 );
    nor g1929 ( n3595 , n2690 , n2258 );
    and g1930 ( n135 , n2577 , n3058 );
    or g1931 ( n1899 , n534 , n605 );
    nor g1932 ( n3047 , n3860 , n65 );
    nor g1933 ( n524 , n2837 , n2182 );
    not g1934 ( n2656 , n1389 );
    or g1935 ( n2691 , n3293 , n735 );
    nor g1936 ( n3380 , n1765 , n2700 );
    not g1937 ( n3165 , n1645 );
    not g1938 ( n2776 , n700 );
    nor g1939 ( n594 , n2549 , n3795 );
    nor g1940 ( n1750 , n851 , n2801 );
    or g1941 ( n3365 , n3098 , n2214 );
    not g1942 ( n2483 , n780 );
    or g1943 ( n2766 , n1135 , n421 );
    nor g1944 ( n2094 , n1745 , n1329 );
    nor g1945 ( n3654 , n2838 , n2370 );
    nor g1946 ( n2511 , n3627 , n3637 );
    and g1947 ( n733 , n2759 , n1300 );
    and g1948 ( n2531 , n481 , n3256 );
    or g1949 ( n2951 , n2997 , n3329 );
    or g1950 ( n921 , n1942 , n1204 );
    not g1951 ( n1662 , n1766 );
    and g1952 ( n264 , n1031 , n1155 );
    and g1953 ( n2591 , n2041 , n3829 );
    and g1954 ( n2756 , n3465 , n2757 );
    or g1955 ( n2974 , n1661 , n2923 );
    nor g1956 ( n811 , n900 , n3015 );
    and g1957 ( n1491 , n1227 , n2114 );
    not g1958 ( n3422 , n3114 );
    and g1959 ( n2813 , n401 , n2596 );
    nor g1960 ( n3661 , n3509 , n1687 );
    not g1961 ( n610 , n1938 );
    or g1962 ( n2956 , n1973 , n13 );
    and g1963 ( n1740 , n2952 , n3829 );
    nor g1964 ( n646 , n603 , n542 );
    nor g1965 ( n3650 , n3092 , n814 );
    or g1966 ( n126 , n981 , n789 );
    and g1967 ( n1198 , n3367 , n3144 );
    not g1968 ( n3215 , n2449 );
    or g1969 ( n2191 , n3447 , n2078 );
    or g1970 ( n155 , n3768 , n1663 );
    or g1971 ( n2675 , n3138 , n3693 );
    nor g1972 ( n554 , n1260 , n3805 );
    or g1973 ( n251 , n591 , n1769 );
    and g1974 ( n3423 , n502 , n269 );
    and g1975 ( n744 , n232 , n1246 );
    or g1976 ( n1889 , n3290 , n741 );
    nor g1977 ( n3235 , n1775 , n2190 );
    or g1978 ( n3566 , n1031 , n1155 );
    nor g1979 ( n2884 , n3600 , n855 );
    nor g1980 ( n25 , n1605 , n3583 );
    or g1981 ( n2195 , n2433 , n789 );
    and g1982 ( n3103 , n211 , n3559 );
    not g1983 ( n406 , n3639 );
    nor g1984 ( n3009 , n89 , n747 );
    or g1985 ( n1972 , n3432 , n2168 );
    nor g1986 ( n3494 , n3694 , n2171 );
    and g1987 ( n3166 , n121 , n1458 );
    and g1988 ( n2697 , n3340 , n2346 );
    or g1989 ( n888 , n463 , n1252 );
    nor g1990 ( n1984 , n2559 , n544 );
    nor g1991 ( n3710 , n861 , n2446 );
    or g1992 ( n2095 , n3750 , n190 );
    and g1993 ( n141 , n3183 , n1166 );
    nor g1994 ( n3075 , n1877 , n157 );
    or g1995 ( n2751 , n877 , n3823 );
    and g1996 ( n2522 , n3827 , n36 );
    or g1997 ( n280 , n79 , n3103 );
    nor g1998 ( n2961 , n3766 , n3242 );
    or g1999 ( n2198 , n1956 , n2057 );
    and g2000 ( n3462 , n3004 , n2369 );
    not g2001 ( n2169 , n1381 );
    or g2002 ( n2519 , n3638 , n393 );
    nor g2003 ( n2904 , n1851 , n2295 );
    and g2004 ( n796 , n2043 , n679 );
    or g2005 ( n2734 , n2894 , n1491 );
    not g2006 ( n2790 , n26 );
    not g2007 ( n2897 , n3539 );
    nor g2008 ( n3464 , n1293 , n691 );
    nor g2009 ( n2701 , n1545 , n1589 );
    nor g2010 ( n1113 , n1051 , n3577 );
    and g2011 ( n2978 , n707 , n1383 );
    or g2012 ( n3577 , n3499 , n1061 );
    and g2013 ( n6 , n1651 , n1398 );
    and g2014 ( n1214 , n1466 , n3737 );
    or g2015 ( n781 , n2486 , n3610 );
    or g2016 ( n2955 , n1493 , n2177 );
    nor g2017 ( n1762 , n1485 , n2111 );
    not g2018 ( n3763 , n1071 );
    nor g2019 ( n852 , n288 , n913 );
    nor g2020 ( n1619 , n764 , n3803 );
    or g2021 ( n1954 , n2635 , n1291 );
    or g2022 ( n138 , n716 , n52 );
    or g2023 ( n845 , n3005 , n2780 );
    or g2024 ( n1756 , n3733 , n2598 );
    and g2025 ( n2740 , n1840 , n1972 );
    nor g2026 ( n1354 , n372 , n1984 );
    nor g2027 ( n2960 , n2053 , n167 );
    nor g2028 ( n2628 , n897 , n1959 );
    and g2029 ( n3141 , n1188 , n2285 );
    or g2030 ( n2714 , n3536 , n498 );
    nor g2031 ( n762 , n1088 , n2811 );
    or g2032 ( n1209 , n167 , n1085 );
    and g2033 ( n1875 , n995 , n231 );
    or g2034 ( n481 , n169 , n2366 );
    or g2035 ( n1468 , n1276 , n2105 );
    nor g2036 ( n3290 , n3050 , n1137 );
    nor g2037 ( n3719 , n1529 , n2243 );
    not g2038 ( n3096 , n585 );
    not g2039 ( n1929 , n1374 );
    and g2040 ( n1970 , n3734 , n923 );
    or g2041 ( n3540 , n1172 , n1895 );
    and g2042 ( n202 , n1975 , n2254 );
    or g2043 ( n3761 , n787 , n1772 );
    not g2044 ( n3787 , n903 );
    and g2045 ( n526 , n3409 , n274 );
    or g2046 ( n2030 , n851 , n212 );
    or g2047 ( n1331 , n2170 , n1082 );
    or g2048 ( n3688 , n2546 , n2650 );
    not g2049 ( n2105 , n972 );
    nor g2050 ( n3310 , n592 , n2445 );
    or g2051 ( n2738 , n2661 , n3601 );
    and g2052 ( n2495 , n866 , n483 );
    nor g2053 ( n2078 , n3156 , n1072 );
    and g2054 ( n2549 , n1082 , n2170 );
    nor g2055 ( n49 , n1611 , n1951 );
    not g2056 ( n3621 , n1172 );
    nor g2057 ( n2275 , n1297 , n1227 );
    or g2058 ( n2725 , n3213 , n1832 );
    nor g2059 ( n2245 , n2705 , n1072 );
    nor g2060 ( n2233 , n2886 , n3181 );
    nor g2061 ( n3594 , n1578 , n3069 );
    and g2062 ( n3378 , n2457 , n535 );
    or g2063 ( n1628 , n1305 , n1798 );
    nor g2064 ( n1330 , n1868 , n3559 );
    nor g2065 ( n552 , n405 , n611 );
    or g2066 ( n755 , n3491 , n3620 );
    or g2067 ( n829 , n821 , n2042 );
    nor g2068 ( n3635 , n833 , n1114 );
    nor g2069 ( n2930 , n3002 , n3474 );
    and g2070 ( n2886 , n2951 , n3412 );
    or g2071 ( n2293 , n518 , n3727 );
    nor g2072 ( n1333 , n2946 , n1755 );
    nor g2073 ( n191 , n1275 , n226 );
    nor g2074 ( n3724 , n2733 , n3516 );
    nor g2075 ( n394 , n1695 , n1357 );
    not g2076 ( n2048 , n2855 );
    not g2077 ( n630 , n3210 );
    not g2078 ( n269 , n3673 );
    nor g2079 ( n815 , n1719 , n3339 );
    nor g2080 ( n2741 , n2124 , n2633 );
    or g2081 ( n3244 , n1293 , n513 );
    or g2082 ( n1363 , n3354 , n285 );
    not g2083 ( n1861 , n542 );
    or g2084 ( n3358 , n25 , n3455 );
    and g2085 ( n941 , n766 , n3597 );
    nor g2086 ( n661 , n2831 , n2910 );
    or g2087 ( n2260 , n1864 , n177 );
    nor g2088 ( n1017 , n3702 , n1673 );
    not g2089 ( n2352 , n790 );
    not g2090 ( n3670 , n1965 );
    nor g2091 ( n3040 , n1522 , n1372 );
    nor g2092 ( n1577 , n1213 , n1428 );
    nor g2093 ( n1196 , n2355 , n87 );
    nor g2094 ( n2558 , n2671 , n1424 );
    or g2095 ( n2994 , n3176 , n1595 );
    not g2096 ( n36 , n3475 );
    or g2097 ( n227 , n1791 , n1726 );
    and g2098 ( n1163 , n3770 , n150 );
    not g2099 ( n839 , n2422 );
    nor g2100 ( n601 , n964 , n2633 );
    nor g2101 ( n2618 , n3310 , n2558 );
    or g2102 ( n1953 , n1601 , n3765 );
    nor g2103 ( n1647 , n184 , n3093 );
    nor g2104 ( n2602 , n561 , n814 );
    and g2105 ( n87 , n1009 , n194 );
    and g2106 ( n211 , n24 , n1658 );
    nor g2107 ( n3437 , n1344 , n3775 );
    nor g2108 ( n440 , n3004 , n2369 );
    or g2109 ( n851 , n364 , n3537 );
    nor g2110 ( n374 , n1111 , n3111 );
    nor g2111 ( n1234 , n3522 , n2691 );
    and g2112 ( n2489 , n3212 , n3198 );
    nor g2113 ( n3572 , n671 , n2595 );
    not g2114 ( n1791 , n3024 );
    and g2115 ( n1901 , n1540 , n3326 );
    not g2116 ( n2170 , n1944 );
    and g2117 ( n2735 , n1120 , n2714 );
    not g2118 ( n1027 , n2990 );
    not g2119 ( n1766 , n1389 );
    or g2120 ( n3135 , n2632 , n208 );
    or g2121 ( n1609 , n248 , n789 );
    nor g2122 ( n3260 , n655 , n809 );
    nor g2123 ( n1159 , n3084 , n3849 );
    nor g2124 ( n3701 , n3203 , n2708 );
    and g2125 ( n1498 , n2268 , n1753 );
    nor g2126 ( n1827 , n1066 , n1665 );
    nor g2127 ( n822 , n456 , n479 );
    not g2128 ( n2168 , n3049 );
    and g2129 ( n1531 , n1692 , n3505 );
    nor g2130 ( n2015 , n3365 , n150 );
    nor g2131 ( n2847 , n381 , n2803 );
    and g2132 ( n2903 , n3412 , n3077 );
    nor g2133 ( n857 , n1046 , n2425 );
    nor g2134 ( n1294 , n294 , n571 );
    nor g2135 ( n520 , n942 , n628 );
    nor g2136 ( n882 , n3606 , n1436 );
    nor g2137 ( n2503 , n3478 , n2899 );
    nor g2138 ( n51 , n3278 , n847 );
    or g2139 ( n3059 , n2179 , n3691 );
    or g2140 ( n2414 , n2681 , n754 );
    and g2141 ( n110 , n187 , n1659 );
    or g2142 ( n1073 , n3641 , n3241 );
    not g2143 ( n416 , n2731 );
    nor g2144 ( n3390 , n2348 , n2406 );
    nor g2145 ( n1732 , n1099 , n665 );
    nor g2146 ( n2510 , n3404 , n1341 );
    nor g2147 ( n2109 , n3320 , n1742 );
    or g2148 ( n3837 , n276 , n373 );
    nor g2149 ( n3804 , n467 , n436 );
    or g2150 ( n1041 , n1449 , n859 );
    nor g2151 ( n752 , n2576 , n3308 );
    and g2152 ( n2385 , n3567 , n300 );
    and g2153 ( n3450 , n870 , n2555 );
    nor g2154 ( n3648 , n2773 , n3593 );
    not g2155 ( n2730 , n119 );
    or g2156 ( n3387 , n2420 , n3197 );
    nor g2157 ( n2323 , n1575 , n3090 );
    not g2158 ( n2810 , n3819 );
    nor g2159 ( n2545 , n482 , n391 );
    or g2160 ( n2040 , n3779 , n2038 );
    nor g2161 ( n3262 , n2389 , n3292 );
    and g2162 ( n1518 , n3042 , n136 );
    and g2163 ( n1569 , n1176 , n936 );
    or g2164 ( n664 , n554 , n2591 );
    or g2165 ( n1856 , n3394 , n2055 );
    or g2166 ( n1681 , n2239 , n810 );
    and g2167 ( n2512 , n1356 , n2824 );
    not g2168 ( n3302 , n3199 );
    and g2169 ( n1632 , n3415 , n1317 );
    or g2170 ( n3530 , n2732 , n3665 );
    and g2171 ( n1836 , n6 , n2421 );
    nor g2172 ( n2278 , n2589 , n2792 );
    or g2173 ( n696 , n2470 , n386 );
    nor g2174 ( n2075 , n2951 , n3412 );
    or g2175 ( n10 , n653 , n2245 );
    not g2176 ( n538 , n1259 );
    not g2177 ( n427 , n678 );
    or g2178 ( n2800 , n255 , n1157 );
    nor g2179 ( n849 , n1868 , n2952 );
    not g2180 ( n38 , n3154 );
    or g2181 ( n920 , n1976 , n57 );
    not g2182 ( n814 , n2656 );
    not g2183 ( n3265 , n3145 );
    and g2184 ( n782 , n439 , n486 );
    or g2185 ( n1679 , n2534 , n2631 );
    nor g2186 ( n2228 , n97 , n384 );
    and g2187 ( n152 , n197 , n1739 );
    nor g2188 ( n1777 , n3418 , n896 );
    or g2189 ( n446 , n54 , n3749 );
    or g2190 ( n705 , n2417 , n3749 );
    nor g2191 ( n1541 , n1964 , n171 );
    and g2192 ( n605 , n2121 , n704 );
    or g2193 ( n3375 , n2543 , n1554 );
    not g2194 ( n1229 , n2444 );
    or g2195 ( n2811 , n1590 , n2918 );
    nor g2196 ( n2214 , n1187 , n1698 );
    or g2197 ( n3685 , n1691 , n1878 );
    nor g2198 ( n1568 , n763 , n3361 );
    or g2199 ( n1029 , n2647 , n3148 );
    nor g2200 ( n1634 , n3370 , n1298 );
    nor g2201 ( n2251 , n3280 , n2017 );
    nor g2202 ( n2542 , n3570 , n3598 );
    or g2203 ( n214 , n2736 , n3241 );
    nor g2204 ( n1594 , n2857 , n1660 );
    and g2205 ( n3503 , n1597 , n3803 );
    not g2206 ( n2410 , n3214 );
    not g2207 ( n686 , n3646 );
    not g2208 ( n2149 , n301 );
    or g2209 ( n306 , n1526 , n2103 );
    or g2210 ( n1909 , n1238 , n3044 );
    nor g2211 ( n3386 , n1636 , n3546 );
    and g2212 ( n2003 , n1483 , n2483 );
    nor g2213 ( n1309 , n2934 , n2628 );
    not g2214 ( n1317 , n1640 );
    not g2215 ( n66 , n712 );
    and g2216 ( n3002 , n3628 , n55 );
    and g2217 ( n370 , n2761 , n1475 );
    nor g2218 ( n3735 , n1094 , n3590 );
    or g2219 ( n3480 , n3467 , n3407 );
    nor g2220 ( n106 , n3139 , n2891 );
    nor g2221 ( n3339 , n565 , n2718 );
    or g2222 ( n3645 , n2968 , n1360 );
    nor g2223 ( n2798 , n944 , n2421 );
    or g2224 ( n879 , n1097 , n1704 );
    and g2225 ( n1365 , n215 , n139 );
    and g2226 ( n3366 , n1988 , n1060 );
    nor g2227 ( n1854 , n1467 , n1539 );
    or g2228 ( n2946 , n2807 , n963 );
    not g2229 ( n3131 , n2806 );
    and g2230 ( n1455 , n2346 , n143 );
    nor g2231 ( n1885 , n835 , n1114 );
    and g2232 ( n303 , n2932 , n610 );
    and g2233 ( n3695 , n3323 , n3096 );
    nor g2234 ( n1949 , n3358 , n3829 );
    or g2235 ( n3568 , n2067 , n73 );
    or g2236 ( n56 , n584 , n1878 );
    and g2237 ( n205 , n55 , n2381 );
    and g2238 ( n2120 , n531 , n3215 );
    nor g2239 ( n116 , n3501 , n742 );
    nor g2240 ( n922 , n1534 , n1662 );
    and g2241 ( n1844 , n844 , n876 );
    or g2242 ( n366 , n2062 , n1008 );
    nor g2243 ( n1368 , n1731 , n640 );
    nor g2244 ( n1743 , n1692 , n2426 );
    or g2245 ( n1872 , n342 , n1056 );
    nor g2246 ( n2349 , n563 , n1606 );
    not g2247 ( n1202 , n3487 );
    not g2248 ( n3598 , n663 );
    or g2249 ( n1666 , n2659 , n1856 );
    and g2250 ( n2292 , n728 , n1760 );
    and g2251 ( n897 , n10 , n2526 );
    nor g2252 ( n1415 , n278 , n3090 );
    not g2253 ( n493 , n3248 );
    not g2254 ( n1551 , n1534 );
    and g2255 ( n3490 , n3818 , n2564 );
    or g2256 ( n1320 , n2908 , n2517 );
    and g2257 ( n2860 , n3544 , n2900 );
    nor g2258 ( n862 , n1889 , n1114 );
    and g2259 ( n3361 , n1967 , n1735 );
    and g2260 ( n3345 , n2112 , n1156 );
    and g2261 ( n331 , n1490 , n3855 );
    not g2262 ( n3559 , n726 );
    and g2263 ( n2803 , n1678 , n1912 );
    or g2264 ( n2396 , n1636 , n857 );
    not g2265 ( n2633 , n2786 );
    and g2266 ( n139 , n437 , n2209 );
    and g2267 ( n1620 , n1064 , n3022 );
    nor g2268 ( n199 , n2536 , n3042 );
    or g2269 ( n957 , n3635 , n2512 );
    nor g2270 ( n943 , n1813 , n1167 );
    not g2271 ( n2421 , n919 );
    nor g2272 ( n598 , n2519 , n1169 );
    nor g2273 ( n540 , n3442 , n1176 );
    or g2274 ( n764 , n1853 , n1900 );
    nor g2275 ( n489 , n3404 , n1603 );
    nor g2276 ( n3452 , n3067 , n3059 );
    nor g2277 ( n1416 , n2289 , n3598 );
    or g2278 ( n3364 , n1049 , n1385 );
    nor g2279 ( n2333 , n1326 , n3337 );
    not g2280 ( n2727 , n2705 );
    not g2281 ( n3396 , n361 );
    and g2282 ( n3053 , n3321 , n1652 );
    and g2283 ( n2808 , n113 , n268 );
    nor g2284 ( n969 , n2402 , n3711 );
    nor g2285 ( n2617 , n161 , n640 );
    or g2286 ( n2673 , n974 , n2492 );
    or g2287 ( n766 , n328 , n2105 );
    or g2288 ( n2152 , n1997 , n988 );
    or g2289 ( n2285 , n3656 , n859 );
    nor g2290 ( n2942 , n710 , n328 );
    and g2291 ( n312 , n3508 , n3115 );
    nor g2292 ( n684 , n3350 , n3622 );
    not g2293 ( n50 , n2636 );
    and g2294 ( n3681 , n1180 , n3799 );
    or g2295 ( n3284 , n646 , n2137 );
    or g2296 ( n3628 , n2972 , n2387 );
    and g2297 ( n1597 , n1952 , n469 );
    and g2298 ( n3516 , n2613 , n3619 );
    nor g2299 ( n2854 , n272 , n322 );
    not g2300 ( n2411 , n2721 );
    nor g2301 ( n163 , n1108 , n3472 );
    or g2302 ( n1957 , n1894 , n2765 );
    nor g2303 ( n518 , n1064 , n2447 );
    or g2304 ( n2515 , n3682 , n3665 );
    nor g2305 ( n2648 , n183 , n2026 );
    and g2306 ( n1486 , n1121 , n1162 );
    or g2307 ( n867 , n2300 , n2686 );
    nor g2308 ( n1530 , n1192 , n3671 );
    nor g2309 ( n2620 , n3717 , n3054 );
    or g2310 ( n3056 , n2754 , n3570 );
    or g2311 ( n3513 , n2876 , n3780 );
    nor g2312 ( n360 , n538 , n2767 );
    or g2313 ( n2158 , n2229 , n845 );
    or g2314 ( n2131 , n3334 , n922 );
    or g2315 ( n232 , n412 , n1181 );
    not g2316 ( n1816 , n3 );
    and g2317 ( n2159 , n2051 , n2421 );
    not g2318 ( n2645 , n278 );
    nor g2319 ( n60 , n2138 , n2531 );
    nor g2320 ( n1465 , n2279 , n2198 );
    nor g2321 ( n1006 , n1324 , n1698 );
    nor g2322 ( n2827 , n237 , n476 );
    or g2323 ( n699 , n1640 , n3601 );
    and g2324 ( n2370 , n587 , n3222 );
    or g2325 ( n459 , n478 , n3845 );
    nor g2326 ( n1729 , n3299 , n1698 );
    not g2327 ( n3031 , n333 );
    nor g2328 ( n495 , n3096 , n3323 );
    or g2329 ( n619 , n1866 , n2287 );
    or g2330 ( n3730 , n3675 , n3810 );
    not g2331 ( n2016 , n1222 );
    not g2332 ( n2026 , n390 );
    not g2333 ( n3090 , n3578 );
    or g2334 ( n2279 , n1110 , n1231 );
    or g2335 ( n3659 , n1583 , n816 );
    nor g2336 ( n2332 , n2414 , n2294 );
    or g2337 ( n1065 , n3199 , n2105 );
    or g2338 ( n1734 , n1030 , n2878 );
    nor g2339 ( n2684 , n1610 , n691 );
    and g2340 ( n1760 , n56 , n1630 );
    or g2341 ( n166 , n187 , n3241 );
    or g2342 ( n2838 , n3828 , n767 );
    or g2343 ( n2355 , n403 , n894 );
    not g2344 ( n3332 , n3325 );
    and g2345 ( n164 , n11 , n3553 );
    nor g2346 ( n1057 , n1433 , n1473 );
    nor g2347 ( n886 , n1459 , n2085 );
    and g2348 ( n363 , n1635 , n2381 );
    nor g2349 ( n1813 , n968 , n1731 );
    nor g2350 ( n2829 , n3792 , n411 );
    and g2351 ( n3434 , n2242 , n3772 );
    not g2352 ( n972 , n3294 );
    nor g2353 ( n2443 , n2627 , n2692 );
    not g2354 ( n611 , n2786 );
    nor g2355 ( n3751 , n3462 , n1148 );
    nor g2356 ( n3655 , n339 , n2585 );
    nor g2357 ( n1900 , n2559 , n1662 );
    nor g2358 ( n1685 , n2848 , n3297 );
    or g2359 ( n1840 , n1965 , n789 );
    nor g2360 ( n2638 , n3312 , n1164 );
    and g2361 ( n1774 , n1411 , n2156 );
    or g2362 ( n3642 , n3493 , n792 );
    or g2363 ( n3687 , n2846 , n1183 );
    nor g2364 ( n1290 , n370 , n2852 );
    or g2365 ( n503 , n2867 , n1969 );
    nor g2366 ( n69 , n598 , n3016 );
    nor g2367 ( n450 , n1337 , n1087 );
    and g2368 ( n527 , n139 , n3805 );
    nor g2369 ( n591 , n3131 , n841 );
    and g2370 ( n482 , n2448 , n141 );
    nor g2371 ( n1937 , n623 , n3137 );
    nor g2372 ( n2654 , n311 , n896 );
    or g2373 ( n352 , n2068 , n2687 );
    nor g2374 ( n1494 , n3231 , n2679 );
    not g2375 ( n1037 , n2248 );
    and g2376 ( n2103 , n976 , n471 );
    and g2377 ( n1369 , n3433 , n2107 );
    not g2378 ( n277 , n3308 );
    and g2379 ( n1361 , n1624 , n2025 );
    or g2380 ( n3510 , n3367 , n738 );
    nor g2381 ( n18 , n3210 , n2298 );
    and g2382 ( n2793 , n2724 , n3032 );
    not g2383 ( n2799 , n663 );
    not g2384 ( n2687 , n959 );
    nor g2385 ( n2182 , n3471 , n293 );
    or g2386 ( n1221 , n2821 , n1907 );
    nor g2387 ( n413 , n1083 , n2544 );
    and g2388 ( n2760 , n1760 , n358 );
    or g2389 ( n2194 , n63 , n3418 );
    not g2390 ( n551 , n1962 );
    or g2391 ( n239 , n1380 , n162 );
    nor g2392 ( n2299 , n2357 , n683 );
    or g2393 ( n788 , n2697 , n2966 );
    and g2394 ( n1056 , n3156 , n770 );
    or g2395 ( n1120 , n2212 , n2439 );
    and g2396 ( n2455 , n1983 , n2755 );
    and g2397 ( n1270 , n345 , n2645 );
    or g2398 ( n817 , n1490 , n2921 );
    or g2399 ( n3276 , n885 , n2434 );
    and g2400 ( n3129 , n2303 , n2335 );
    and g2401 ( n3579 , n3106 , n1767 );
    nor g2402 ( n668 , n3274 , n396 );
    nor g2403 ( n3705 , n74 , n3829 );
    nor g2404 ( n2718 , n2723 , n2024 );
    and g2405 ( n1562 , n1723 , n367 );
    nor g2406 ( n2977 , n360 , n3342 );
    or g2407 ( n3517 , n1694 , n2995 );
    and g2408 ( n1296 , n2928 , n1759 );
    and g2409 ( n2569 , n3021 , n3782 );
    nor g2410 ( n791 , n735 , n684 );
    or g2411 ( n304 , n1352 , n2219 );
    not g2412 ( n770 , n1904 );
    nor g2413 ( n3430 , n3218 , n996 );
    not g2414 ( n2980 , n3702 );
    not g2415 ( n2001 , n368 );
    nor g2416 ( n1626 , n269 , n502 );
    or g2417 ( n194 , n198 , n1895 );
    and g2418 ( n3073 , n1702 , n3070 );
    nor g2419 ( n1340 , n2989 , n3674 );
    not g2420 ( n2204 , n2812 );
    not g2421 ( n390 , n1389 );
    or g2422 ( n201 , n2291 , n819 );
    nor g2423 ( n72 , n1968 , n2827 );
    or g2424 ( n98 , n175 , n2804 );
    not g2425 ( n1776 , n3318 );
    and g2426 ( n3630 , n3178 , n1512 );
    nor g2427 ( n391 , n2356 , n3064 );
    or g2428 ( n541 , n1966 , n3646 );
    or g2429 ( n1350 , n3475 , n1929 );
    or g2430 ( n3283 , n3303 , n1538 );
    and g2431 ( n2492 , n2929 , n1803 );
    nor g2432 ( n1858 , n2796 , n2554 );
    nor g2433 ( n2859 , n3358 , n1292 );
    nor g2434 ( n1572 , n2748 , n3060 );
    or g2435 ( n3818 , n2167 , n1033 );
    nor g2436 ( n1943 , n1043 , n3252 );
    or g2437 ( n1535 , n122 , n748 );
    or g2438 ( n2265 , n1787 , n1235 );
    nor g2439 ( n2486 , n1834 , n1302 );
    or g2440 ( n924 , n944 , n1311 );
    and g2441 ( n2205 , n141 , n3077 );
    or g2442 ( n1247 , n2201 , n3650 );
    not g2443 ( n3161 , n1941 );
    and g2444 ( n3076 , n3561 , n3343 );
    and g2445 ( n2779 , n833 , n1356 );
    or g2446 ( n2401 , n2828 , n1869 );
    and g2447 ( n914 , n3514 , n1827 );
    not g2448 ( n1893 , n386 );
    or g2449 ( n1213 , n2404 , n3542 );
    and g2450 ( n2526 , n801 , n645 );
    or g2451 ( n3762 , n3705 , n3853 );
    and g2452 ( n3086 , n2008 , n115 );
    nor g2453 ( n2907 , n3001 , n796 );
    not g2454 ( n2147 , n916 );
    or g2455 ( n2085 , n59 , n2476 );
    nor g2456 ( n741 , n1051 , n1662 );
    nor g2457 ( n3777 , n1775 , n2465 );
    or g2458 ( n419 , n2077 , n2652 );
    or g2459 ( n2430 , n1210 , n359 );
    or g2460 ( n1638 , n2478 , n1554 );
    or g2461 ( n1586 , n1431 , n1173 );
    or g2462 ( n2199 , n235 , n1985 );
    or g2463 ( n1747 , n462 , n1385 );
    and g2464 ( n2346 , n3575 , n448 );
    or g2465 ( n1795 , n1645 , n2366 );
    and g2466 ( n1521 , n1913 , n3193 );
    not g2467 ( n377 , n3245 );
    nor g2468 ( n677 , n3533 , n1720 );
    nor g2469 ( n62 , n3763 , n2484 );
    nor g2470 ( n3651 , n540 , n1647 );
    nor g2471 ( n926 , n335 , n2977 );
    nor g2472 ( n29 , n685 , n896 );
    or g2473 ( n1592 , n3800 , n2485 );
    nor g2474 ( n1231 , n2046 , n682 );
    or g2475 ( n295 , n2188 , n2200 );
    or g2476 ( n2535 , n995 , n1798 );
    and g2477 ( n73 , n134 , n1229 );
    and g2478 ( n1210 , n2296 , n1358 );
    or g2479 ( n1830 , n2879 , n2320 );
    or g2480 ( n384 , n2790 , n3841 );
    or g2481 ( n1636 , n1408 , n3454 );
    nor g2482 ( n3633 , n3816 , n297 );
    nor g2483 ( n673 , n543 , n275 );
    or g2484 ( n196 , n620 , n1878 );
    nor g2485 ( n2193 , n1434 , n2392 );
    nor g2486 ( n1643 , n3362 , n2890 );
    and g2487 ( n3596 , n3287 , n2359 );
    not g2488 ( n2957 , n2002 );
    and g2489 ( n2477 , n328 , n710 );
    nor g2490 ( n449 , n1440 , n322 );
    or g2491 ( n2473 , n1497 , n1618 );
    nor g2492 ( n2419 , n3550 , n931 );
    not g2493 ( n2973 , n1220 );
    and g2494 ( n2830 , n971 , n772 );
    or g2495 ( n2872 , n511 , n3746 );
    nor g2496 ( n343 , n3548 , n3208 );
    nor g2497 ( n2908 , n1058 , n3553 );
    and g2498 ( n1189 , n3473 , n159 );
    nor g2499 ( n3713 , n3649 , n358 );
    or g2500 ( n1308 , n454 , n2648 );
    or g2501 ( n2286 , n133 , n3378 );
    and g2502 ( n1768 , n2437 , n1450 );
    not g2503 ( n1109 , n1822 );
    or g2504 ( n1653 , n1393 , n1291 );
    not g2505 ( n1295 , n2352 );
    nor g2506 ( n1387 , n381 , n2114 );
    or g2507 ( n1625 , n1756 , n1616 );
    and g2508 ( n3091 , n2172 , n399 );
    nor g2509 ( n1407 , n138 , n2941 );
    nor g2510 ( n1168 , n776 , n3414 );
    or g2511 ( n1684 , n151 , n555 );
    and g2512 ( n1821 , n3606 , n1357 );
    and g2513 ( n579 , n3725 , n2727 );
    nor g2514 ( n329 , n2327 , n3735 );
    or g2515 ( n2912 , n2917 , n33 );
    and g2516 ( n2640 , n732 , n902 );
    and g2517 ( n266 , n3839 , n3484 );
    not g2518 ( n348 , n177 );
    or g2519 ( n2880 , n2587 , n3629 );
    not g2520 ( n2900 , n2052 );
    not g2521 ( n2570 , n2590 );
    and g2522 ( n1142 , n2004 , n2221 );
    or g2523 ( n279 , n301 , n3241 );
    not g2524 ( n2875 , n3401 );
    nor g2525 ( n1373 , n178 , n2026 );
    nor g2526 ( n2343 , n3791 , n1501 );
    nor g2527 ( n3806 , n960 , n2091 );
    or g2528 ( n1070 , n1220 , n1126 );
    and g2529 ( n2513 , n1293 , n513 );
    nor g2530 ( n1525 , n2308 , n3200 );
    not g2531 ( n2335 , n3854 );
    nor g2532 ( n3760 , n3841 , n1228 );
    nor g2533 ( n1205 , n2855 , n2026 );
    or g2534 ( n3251 , n2140 , n1085 );
    nor g2535 ( n1781 , n3802 , n882 );
    not g2536 ( n701 , n2457 );
    or g2537 ( n3543 , n3535 , n1421 );
    nor g2538 ( n637 , n1361 , n3568 );
    or g2539 ( n2909 , n34 , n2739 );
    or g2540 ( n1780 , n2611 , n3346 );
    or g2541 ( n3839 , n3304 , n3648 );
    nor g2542 ( n2976 , n3522 , n847 );
    not g2543 ( n2743 , n3321 );
    not g2544 ( n2189 , n2027 );
    or g2545 ( n458 , n416 , n1361 );
    or g2546 ( n3856 , n1964 , n3745 );
    and g2547 ( n3187 , n1891 , n2447 );
    nor g2548 ( n2377 , n3284 , n1410 );
    nor g2549 ( n2070 , n3567 , n1648 );
    nor g2550 ( n1077 , n542 , n3593 );
    nor g2551 ( n79 , n3624 , n226 );
    nor g2552 ( n680 , n445 , n2306 );
    and g2553 ( n749 , n1749 , n2695 );
    or g2554 ( n1913 , n532 , n3594 );
    nor g2555 ( n899 , n267 , n358 );
    nor g2556 ( n1723 , n1054 , n508 );
    or g2557 ( n3797 , n2235 , n423 );
    and g2558 ( n2408 , n2508 , n2749 );
    or g2559 ( n2833 , n1833 , n1569 );
    and g2560 ( n3236 , n1928 , n226 );
    nor g2561 ( n1236 , n3664 , n3040 );
    or g2562 ( n940 , n191 , n164 );
    nor g2563 ( n3394 , n704 , n2121 );
    or g2564 ( n2643 , n3302 , n2636 );
    and g2565 ( n3709 , n1787 , n3422 );
    and g2566 ( n2388 , n243 , n1586 );
    and g2567 ( n2156 , n2926 , n1429 );
    or g2568 ( n1499 , n1417 , n2402 );
    or g2569 ( n2165 , n753 , n2921 );
    or g2570 ( n323 , n3123 , n329 );
    and g2571 ( n1300 , n234 , n446 );
    or g2572 ( n3742 , n2886 , n1829 );
    nor g2573 ( n1481 , n318 , n1691 );
    or g2574 ( n2509 , n1175 , n499 );
    nor g2575 ( n2022 , n3220 , n3299 );
    nor g2576 ( n2589 , n2437 , n2949 );
    nor g2577 ( n3029 , n506 , n640 );
    and g2578 ( n1122 , n2445 , n592 );
    nor g2579 ( n490 , n967 , n2884 );
    nor g2580 ( n616 , n1696 , n441 );
    nor g2581 ( n742 , n1756 , n490 );
    nor g2582 ( n1081 , n1064 , n3022 );
    nor g2583 ( n860 , n1599 , n929 );
    or g2584 ( n692 , n499 , n2073 );
    not g2585 ( n3488 , n620 );
    not g2586 ( n724 , n3001 );
    and g2587 ( n3812 , n577 , n1145 );
    or g2588 ( n2983 , n1686 , n2532 );
    and g2589 ( n1248 , n3218 , n2432 );
    nor g2590 ( n872 , n2393 , n3583 );
    nor g2591 ( n77 , n1475 , n2761 );
    or g2592 ( n3460 , n2287 , n3349 );
    and g2593 ( n1024 , n441 , n1696 );
    and g2594 ( n35 , n1341 , n1603 );
    nor g2595 ( n2870 , n803 , n1689 );
    and g2596 ( n1038 , n2834 , n3663 );
    not g2597 ( n1532 , n2712 );
    or g2598 ( n2033 , n1479 , n1299 );
    or g2599 ( n501 , n1785 , n1929 );
    and g2600 ( n1704 , n75 , n3217 );
    or g2601 ( n1353 , n231 , n303 );
    and g2602 ( n3838 , n2525 , n938 );
    nor g2603 ( n3169 , n3352 , n1921 );
    or g2604 ( n2281 , n1767 , n1503 );
    not g2605 ( n2464 , n1433 );
    and g2606 ( n1176 , n714 , n2728 );
    and g2607 ( n3773 , n1401 , n2630 );
    and g2608 ( n55 , n3174 , n2000 );
    and g2609 ( n1299 , n978 , n2595 );
    nor g2610 ( n1375 , n2588 , n2421 );
    nor g2611 ( n325 , n1944 , n1082 );
    and g2612 ( n3402 , n3127 , n3805 );
    nor g2613 ( n2013 , n3486 , n2312 );
    nor g2614 ( n3411 , n2769 , n1425 );
    not g2615 ( n1458 , n578 );
    nor g2616 ( n162 , n121 , n3842 );
    or g2617 ( n1613 , n3693 , n1085 );
    or g2618 ( n1279 , n743 , n3227 );
    nor g2619 ( n491 , n3734 , n322 );
    not g2620 ( n660 , n1865 );
    nor g2621 ( n1570 , n2118 , n1794 );
    or g2622 ( n3124 , n1776 , n1924 );
    not g2623 ( n2392 , n3743 );
    nor g2624 ( n276 , n1247 , n3217 );
    not g2625 ( n534 , n2915 );
    or g2626 ( n3611 , n2552 , n434 );
    and g2627 ( n2341 , n1442 , n1666 );
    not g2628 ( n1703 , n2068 );
    not g2629 ( n1860 , n2862 );
    or g2630 ( n382 , n4 , n2141 );
    nor g2631 ( n1754 , n432 , n95 );
    and g2632 ( n754 , n627 , n2888 );
    nor g2633 ( n975 , n2556 , n784 );
    not g2634 ( n1450 , n2014 );
    or g2635 ( n1496 , n891 , n2135 );
    or g2636 ( n1059 , n500 , n3423 );
    or g2637 ( n3136 , n3419 , n2988 );
    or g2638 ( n3836 , n1643 , n129 );
    and g2639 ( n3731 , n837 , n2540 );
    and g2640 ( n2363 , n462 , n2881 );
    nor g2641 ( n955 , n3728 , n1187 );
    or g2642 ( n1138 , n3667 , n2385 );
    nor g2643 ( n2162 , n99 , n2421 );
    nor g2644 ( n371 , n3388 , n1743 );
    or g2645 ( n1457 , n2242 , n3765 );
    nor g2646 ( n3449 , n781 , n136 );
    and g2647 ( n3349 , n1351 , n1866 );
    not g2648 ( n772 , n2985 );
    or g2649 ( n855 , n1889 , n3027 );
    nor g2650 ( n3351 , n770 , n3156 );
    nor g2651 ( n1459 , n1881 , n2820 );
    or g2652 ( n3082 , n1844 , n644 );
    or g2653 ( n1606 , n3603 , n2364 );
    and g2654 ( n11 , n715 , n3172 );
    or g2655 ( n3451 , n2129 , n1534 );
    not g2656 ( n847 , n1766 );
    and g2657 ( n1421 , n929 , n3803 );
    or g2658 ( n321 , n1934 , n3385 );
    not g2659 ( n1072 , n3374 );
    nor g2660 ( n2845 , n1925 , n1596 );
    not g2661 ( n859 , n1140 );
    nor g2662 ( n3328 , n195 , n1449 );
    nor g2663 ( n287 , n3106 , n2281 );
    or g2664 ( n2514 , n1489 , n414 );
    and g2665 ( n3116 , n94 , n3268 );
    or g2666 ( n1492 , n1881 , n3091 );
    not g2667 ( n1497 , n3776 );
    nor g2668 ( n2677 , n37 , n631 );
    or g2669 ( n2940 , n869 , n3589 );
    not g2670 ( n3485 , n2218 );
    or g2671 ( n243 , n357 , n2417 );
    or g2672 ( n2394 , n1174 , n347 );
    nor g2673 ( n410 , n2183 , n3069 );
    not g2674 ( n3112 , n2096 );
    nor g2675 ( n1245 , n2126 , n2034 );
    or g2676 ( n3565 , n2312 , n3601 );
    and g2677 ( n1155 , n1795 , n2337 );
    or g2678 ( n3003 , n1589 , n3749 );
    or g2679 ( n267 , n599 , n3439 );
    nor g2680 ( n1080 , n525 , n3842 );
    not g2681 ( n1263 , n1722 );
    and g2682 ( n2945 , n2023 , n1412 );
    nor g2683 ( n2238 , n1118 , n2956 );
    nor g2684 ( n1 , n3552 , n1253 );
    and g2685 ( n2304 , n3089 , n2565 );
    and g2686 ( n961 , n2909 , n1635 );
    or g2687 ( n3356 , n3704 , n378 );
    or g2688 ( n1237 , n582 , n1929 );
    not g2689 ( n2432 , n3682 );
    nor g2690 ( n1244 , n109 , n2920 );
    or g2691 ( n1697 , n1349 , n15 );
    not g2692 ( n1973 , n3573 );
    and g2693 ( n3537 , n835 , n242 );
    or g2694 ( n94 , n2321 , n3601 );
    not g2695 ( n2665 , n2616 );
    not g2696 ( n3772 , n2478 );
    or g2697 ( n606 , n2331 , n3380 );
    nor g2698 ( n2789 , n3709 , n1347 );
    or g2699 ( n365 , n1793 , n2702 );
    not g2700 ( n790 , n460 );
    nor g2701 ( n151 , n1962 , n1037 );
    nor g2702 ( n2831 , n2727 , n3725 );
    and g2703 ( n999 , n119 , n3317 );
    nor g2704 ( n2056 , n1841 , n2381 );
    or g2705 ( n1346 , n257 , n307 );
    or g2706 ( n1547 , n2014 , n3601 );
    or g2707 ( n2565 , n2889 , n859 );
    and g2708 ( n530 , n3630 , n2381 );
    nor g2709 ( n1890 , n2802 , n0 );
    nor g2710 ( n2670 , n3456 , n1830 );
    not g2711 ( n143 , n3372 );
    nor g2712 ( n1508 , n585 , n2190 );
    or g2713 ( n327 , n1765 , n2237 );
    nor g2714 ( n443 , n2840 , n2036 );
    nor g2715 ( n3512 , n2484 , n157 );
    or g2716 ( n1306 , n2176 , n1267 );
    or g2717 ( n562 , n3626 , n2532 );
    and g2718 ( n415 , n2468 , n3032 );
    or g2719 ( n1313 , n2651 , n1484 );
    and g2720 ( n589 , n1297 , n1227 );
    not g2721 ( n1966 , n1800 );
    or g2722 ( n340 , n2955 , n3416 );
    not g2723 ( n3728 , n474 );
    not g2724 ( n1126 , n3625 );
    and g2725 ( n1417 , n3684 , n3087 );
    and g2726 ( n3297 , n1447 , n1613 );
    and g2727 ( n745 , n1695 , n782 );
    nor g2728 ( n3591 , n2750 , n526 );
    or g2729 ( n813 , n2472 , n2666 );
    nor g2730 ( n2997 , n1822 , n68 );
    or g2731 ( n3712 , n3128 , n1808 );
    nor g2732 ( n1536 , n1918 , n20 );
    or g2733 ( n895 , n1315 , n1291 );
    nor g2734 ( n3821 , n266 , n450 );
    not g2735 ( n974 , n256 );
    or g2736 ( n2469 , n2444 , n43 );
    nor g2737 ( n609 , n3654 , n1567 );
    and g2738 ( n2089 , n399 , n2824 );
    and g2739 ( n3668 , n662 , n871 );
    and g2740 ( n3767 , n3406 , n2824 );
    nor g2741 ( n288 , n2098 , n649 );
    and g2742 ( n1820 , n2944 , n3261 );
    or g2743 ( n2777 , n38 , n1172 );
    and g2744 ( n2218 , n27 , n934 );
    nor g2745 ( n3101 , n2499 , n155 );
    or g2746 ( n1585 , n1857 , n1345 );
    or g2747 ( n2424 , n839 , n236 );
    and g2748 ( n2778 , n2424 , n695 );
    nor g2749 ( n2086 , n2737 , n361 );
    and g2750 ( n1974 , n725 , n2456 );
    or g2751 ( n1429 , n3721 , n738 );
    or g2752 ( n140 , n2993 , n3075 );
    not g2753 ( n174 , n236 );
    and g2754 ( n2782 , n3826 , n1710 );
    nor g2755 ( n1969 , n3337 , n1998 );
    not g2756 ( n3216 , n2773 );
    nor g2757 ( n1661 , n763 , n3559 );
    not g2758 ( n2317 , n878 );
    not g2759 ( n64 , n919 );
    and g2760 ( n3037 , n1547 , n1171 );
    nor g2761 ( n1461 , n354 , n143 );
    nor g2762 ( n3847 , n1580 , n611 );
    not g2763 ( n3636 , n2312 );
    nor g2764 ( n1940 , n1278 , n594 );
    nor g2765 ( n1040 , n263 , n2236 );
    nor g2766 ( n2167 , n1736 , n2243 );
    not g2767 ( n2791 , n1049 );
    or g2768 ( n3300 , n712 , n2366 );
    or g2769 ( n2479 , n987 , n2938 );
    or g2770 ( n2746 , n2896 , n3749 );
    or g2771 ( n1728 , n733 , n2123 );
    nor g2772 ( n2429 , n1420 , n3842 );
    and g2773 ( n2551 , n109 , n3161 );
    nor g2774 ( n3171 , n1085 , n3743 );
    or g2775 ( n2301 , n939 , n1541 );
    and g2776 ( n2032 , n501 , n252 );
    nor g2777 ( n1482 , n2600 , n1309 );
    nor g2778 ( n2523 , n686 , n1800 );
    nor g2779 ( n2351 , n677 , n2270 );
    or g2780 ( n3846 , n1201 , n3588 );
    and g2781 ( n1443 , n3504 , n3574 );
    or g2782 ( n3221 , n1659 , n3196 );
    or g2783 ( n1399 , n1688 , n2984 );
    nor g2784 ( n259 , n2423 , n2635 );
    not g2785 ( n3440 , n1580 );
    nor g2786 ( n1143 , n1710 , n3826 );
    nor g2787 ( n3305 , n2931 , n2207 );
    nor g2788 ( n337 , n678 , n814 );
    and g2789 ( n3416 , n762 , n39 );
    not g2790 ( n3341 , n2507 );
    or g2791 ( n3575 , n2975 , n1554 );
    nor g2792 ( n2874 , n77 , n1244 );
    nor g2793 ( n185 , n3044 , n3069 );
    and g2794 ( n3823 , n1600 , n150 );
    or g2795 ( n3616 , n2296 , n3241 );
    nor g2796 ( n2999 , n2877 , n1559 );
    or g2797 ( n2508 , n3741 , n525 );
    nor g2798 ( n2739 , n2767 , n3593 );
    nor g2799 ( n676 , n1611 , n3559 );
    nor g2800 ( n2948 , n1782 , n2447 );
    and g2801 ( n1824 , n1780 , n2819 );
    or g2802 ( n2268 , n3798 , n3104 );
    nor g2803 ( n1677 , n1623 , n3842 );
    nor g2804 ( n3160 , n1007 , n3398 );
    or g2805 ( n1130 , n177 , n1985 );
    and g2806 ( n2041 , n1104 , n3796 );
    nor g2807 ( n326 , n2605 , n487 );
    or g2808 ( n381 , n3030 , n2490 );
    and g2809 ( n1994 , n1488 , n517 );
    not g2810 ( n3744 , n688 );
    or g2811 ( n1383 , n32 , n1071 );
    not g2812 ( n1475 , n2975 );
    or g2813 ( n944 , n3719 , n1373 );
    nor g2814 ( n1167 , n966 , n2664 );
    not g2815 ( n1646 , n1575 );
    or g2816 ( n626 , n118 , n2230 );
    or g2817 ( n1359 , n440 , n1159 );
    nor g2818 ( n3137 , n2693 , n458 );
    and g2819 ( n3551 , n99 , n70 );
    not g2820 ( n1698 , n2656 );
    or g2821 ( n2769 , n2580 , n2905 );
    nor g2822 ( n3555 , n3788 , n296 );
    or g2823 ( n1289 , n932 , n2366 );
    or g2824 ( n3495 , n3313 , n1189 );
    nor g2825 ( n2933 , n1623 , n1872 );
    and g2826 ( n2802 , n2851 , n2240 );
    or g2827 ( n1256 , n3464 , n798 );
    not g2828 ( n1035 , n1268 );
    and g2829 ( n142 , n698 , n3669 );
    nor g2830 ( n2145 , n466 , n1977 );
    or g2831 ( n3206 , n1949 , n244 );
    or g2832 ( n1177 , n1101 , n1362 );
    or g2833 ( n1944 , n1477 , n2483 );
    nor g2834 ( n3556 , n1701 , n1473 );
    nor g2835 ( n934 , n1832 , n861 );
    nor g2836 ( n2153 , n387 , n317 );
    or g2837 ( n3312 , n3369 , n3152 );
    and g2838 ( n1971 , n781 , n875 );
    or g2839 ( n2944 , n2581 , n1080 );
    or g2840 ( n544 , n2204 , n1996 );
    or g2841 ( n2020 , n353 , n2096 );
    and g2842 ( n798 , n513 , n300 );
    nor g2843 ( n2452 , n3005 , n1992 );
    nor g2844 ( n748 , n1351 , n1662 );
    or g2845 ( n1611 , n2282 , n1508 );
    or g2846 ( n1658 , n2263 , n738 );
    or g2847 ( n779 , n2913 , n755 );
    nor g2848 ( n1334 , n3820 , n1072 );
    or g2849 ( n1907 , n1336 , n254 );
    or g2850 ( n662 , n223 , n3141 );
    or g2851 ( n3084 , n731 , n3479 );
    or g2852 ( n645 , n1045 , n1798 );
    or g2853 ( n3643 , n3143 , n2687 );
    nor g2854 ( n816 , n3644 , n593 );
    nor g2855 ( n871 , n2072 , n2070 );
    not g2856 ( n3601 , n959 );
    and g2857 ( n1832 , n479 , n456 );
    nor g2858 ( n1523 , n134 , n488 );
    or g2859 ( n2174 , n1011 , n2945 );
    or g2860 ( n2398 , n449 , n58 );
    and g2861 ( n3010 , n1446 , n535 );
    or g2862 ( n1020 , n2965 , n2617 );
    or g2863 ( n1602 , n2247 , n1283 );
    or g2864 ( n111 , n3855 , n1490 );
    and g2865 ( n3179 , n81 , n614 );
    nor g2866 ( n270 , n3637 , n3842 );
    or g2867 ( n1797 , n1746 , n3506 );
    not g2868 ( n2163 , n2553 );
    and g2869 ( n359 , n3157 , n2059 );
    not g2870 ( n2858 , n3250 );
    nor g2871 ( n1144 , n479 , n847 );
    and g2872 ( n4 , n1371 , n534 );
    and g2873 ( n1829 , n965 , n1778 );
    nor g2874 ( n2399 , n3301 , n3668 );
    or g2875 ( n588 , n2131 , n1721 );
    not g2876 ( n1291 , n972 );
    or g2877 ( n3441 , n2943 , n3386 );
    nor g2878 ( n2563 , n3624 , n211 );
    nor g2879 ( n247 , n91 , n1487 );
    or g2880 ( n3183 , n848 , n1929 );
    or g2881 ( n2759 , n21 , n2113 );
    or g2882 ( n1000 , n3784 , n3840 );
    or g2883 ( n61 , n1579 , n2806 );
    nor g2884 ( n220 , n3689 , n1676 );
    nor g2885 ( n28 , n836 , n2190 );
    nor g2886 ( n86 , n3787 , n1578 );
    or g2887 ( n2240 , n2671 , n2200 );
    and g2888 ( n1595 , n1909 , n943 );
    or g2889 ( n71 , n3357 , n901 );
    not g2890 ( n485 , n1726 );
    or g2891 ( n2913 , n1639 , n2217 );
    not g2892 ( n2447 , n2482 );
    or g2893 ( n3033 , n2916 , n3062 );
    nor g2894 ( n3338 , n2375 , n2431 );
    nor g2895 ( n3610 , n1975 , n665 );
    not g2896 ( n2540 , n217 );
    not g2897 ( n1894 , n2203 );
    nor g2898 ( n128 , n2678 , n1471 );
    and g2899 ( n3122 , n381 , n2803 );
    or g2900 ( n2949 , n1450 , n1198 );
    and g2901 ( n3704 , n1108 , n1048 );
    or g2902 ( n2879 , n2302 , n1763 );
    not g2903 ( n2298 , n2656 );
    nor g2904 ( n853 , n958 , n896 );
    or g2905 ( n1121 , n29 , n1100 );
    nor g2906 ( n1852 , n1143 , n2213 );
    not g2907 ( n1255 , n571 );
    and g2908 ( n2217 , n1535 , n2489 );
    or g2909 ( n1275 , n2603 , n918 );
    and g2910 ( n435 , n2157 , n1418 );
    nor g2911 ( n3360 , n3659 , n2106 );
    or g2912 ( n2231 , n3054 , n2200 );
    and g2913 ( n3189 , n2138 , n2531 );
    or g2914 ( n2273 , n2269 , n3171 );
    nor g2915 ( n1660 , n647 , n2396 );
    or g2916 ( n2536 , n3602 , n2529 );
    nor g2917 ( n2594 , n806 , n1222 );
    or g2918 ( n2071 , n3314 , n3840 );
    or g2919 ( n671 , n552 , n1057 );
    and g2920 ( n1026 , n962 , n1348 );
    nor g2921 ( n675 , n124 , n772 );
    or g2922 ( n1405 , n3154 , n3601 );
    and g2923 ( n3134 , n2407 , n2001 );
    and g2924 ( n1282 , n172 , n3032 );
    or g2925 ( n942 , n2208 , n3160 );
    nor g2926 ( n2336 , n3279 , n327 );
    and g2927 ( n3435 , n2494 , n3355 );
    nor g2928 ( n928 , n1161 , n608 );
    nor g2929 ( n1042 , n1411 , n2597 );
    nor g2930 ( n2719 , n2794 , n1504 );
    not g2931 ( n1993 , n2431 );
    and g2932 ( n373 , n2802 , n1598 );
    or g2933 ( n2958 , n3751 , n47 );
    or g2934 ( n1152 , n2120 , n1922 );
    and g2935 ( n1753 , n973 , n1209 );
    not g2936 ( n475 , n1141 );
    nor g2937 ( n496 , n1156 , n2112 );
    nor g2938 ( n1423 , n2569 , n2164 );
    and g2939 ( n3474 , n1146 , n3606 );
    nor g2940 ( n2804 , n508 , n3099 );
    nor g2941 ( n908 , n995 , n1353 );
    and g2942 ( n1091 , n2622 , n3061 );
    nor g2943 ( n3200 , n2374 , n1621 );
    or g2944 ( n840 , n1288 , n1836 );
    not g2945 ( n2921 , n1722 );
    or g2946 ( n3740 , n2553 , n3346 );
    nor g2947 ( n3677 , n2256 , n546 );
    or g2948 ( n1712 , n1218 , n750 );
    or g2949 ( n3489 , n3600 , n1649 );
    nor g2950 ( n1485 , n2622 , n3061 );
    and g2951 ( n1240 , n87 , n2447 );
    nor g2952 ( n222 , n2034 , n847 );
    nor g2953 ( n3471 , n1478 , n1285 );
    nor g2954 ( n2047 , n2832 , n2712 );
    or g2955 ( n1915 , n2898 , n3731 );
    nor g2956 ( n1288 , n3611 , n2447 );
    and g2957 ( n948 , n3009 , n112 );
    and g2958 ( n580 , n1118 , n1973 );
    or g2959 ( n22 , n2730 , n2743 );
    or g2960 ( n354 , n2145 , n2358 );
    nor g2961 ( n2100 , n1322 , n1137 );
    or g2962 ( n1676 , n2864 , n3277 );
    and g2963 ( n3344 , n608 , n1161 );
    nor g2964 ( n3229 , n2703 , n1152 );
    nor g2965 ( n3706 , n1803 , n2929 );
    nor g2966 ( n175 , n2493 , n2768 );
    or g2967 ( n2642 , n793 , n1531 );
    or g2968 ( n545 , n1826 , n1144 );
    or g2969 ( n2926 , n2002 , n1878 );
    and g2970 ( n2969 , n124 , n3630 );
    nor g2971 ( n510 , n844 , n876 );
    or g2972 ( n3409 , n76 , n3785 );
    and g2973 ( n3691 , n1831 , n3680 );
    nor g2974 ( n3011 , n2441 , n609 );
    nor g2975 ( n3815 , n785 , n622 );
    nor g2976 ( n2101 , n224 , n262 );
    or g2977 ( n2266 , n3396 , n3801 );
    or g2978 ( n2840 , n3538 , n1092 );
    nor g2979 ( n516 , n2075 , n2233 );
    and g2980 ( n2327 , n1736 , n2742 );
    nor g2981 ( n2774 , n1404 , n3188 );
    nor g2982 ( n20 , n3698 , n1961 );
    not g2983 ( n389 , n405 );
    or g2984 ( n870 , n1406 , n1286 );
    nor g2985 ( n3331 , n711 , n1137 );
    nor g2986 ( n1838 , n199 , n2301 );
    or g2987 ( n2564 , n2455 , n3048 );
    and g2988 ( n2580 , n1437 , n1446 );
    nor g2989 ( n2898 , n2317 , n667 );
    or g2990 ( n1520 , n3157 , n1484 );
    and g2991 ( n3313 , n3624 , n211 );
    nor g2992 ( n2196 , n3325 , n2298 );
    or g2993 ( n1630 , n1108 , n1895 );
    nor g2994 ( n1991 , n1091 , n1762 );
    or g2995 ( n1629 , n559 , n3503 );
    not g2996 ( n1003 , n3417 );
    nor g2997 ( n3531 , n148 , n2414 );
    nor g2998 ( n1344 , n1993 , n2971 );
    or g2999 ( n2781 , n3318 , n2532 );
    nor g3000 ( n1370 , n3835 , n575 );
    not g3001 ( n2098 , n2034 );
    and g3002 ( n2598 , n1020 , n2468 );
    or g3003 ( n3714 , n548 , n2624 );
    or g3004 ( n3689 , n1131 , n125 );
    nor g3005 ( n257 , n1504 , n2243 );
    nor g3006 ( n1716 , n223 , n3805 );
    and g3007 ( n2797 , n2361 , n1986 );
    nor g3008 ( n3238 , n3832 , n903 );
    or g3009 ( n3850 , n570 , n2602 );
    nor g3010 ( n918 , n2693 , n1473 );
    or g3011 ( n1773 , n3706 , n3117 );
    and g3012 ( n3863 , n3261 , n691 );
    not g3013 ( n2576 , n1700 );
    not g3014 ( n2006 , n557 );
    nor g3015 ( n375 , n803 , n3077 );
    or g3016 ( n252 , n1397 , n2200 );
    or g3017 ( n3315 , n74 , n1552 );
    and g3018 ( n1408 , n123 , n3376 );
    or g3019 ( n3233 , n2383 , n2904 );
    not g3020 ( n209 , n1988 );
    not g3021 ( n3190 , n2488 );
    and g3022 ( n581 , n3660 , n811 );
    and g3023 ( n2457 , n865 , n3510 );
    not g3024 ( n1759 , n3700 );
    nor g3025 ( n2837 , n3526 , n3214 );
    or g3026 ( n3222 , n2439 , n1895 );
    or g3027 ( n3814 , n1330 , n1740 );
    or g3028 ( n2750 , n120 , n1499 );
    and g3029 ( n2600 , n140 , n1191 );
    not g3030 ( n1083 , n2289 );
    or g3031 ( n2453 , n2100 , n2115 );
    nor g3032 ( n912 , n2862 , n95 );
    or g3033 ( n3405 , n1971 , n472 );
    nor g3034 ( n1430 , n994 , n611 );
    or g3035 ( n1505 , n1003 , n3718 );
    or g3036 ( n3676 , n1461 , n2927 );
    nor g3037 ( n2365 , n842 , n1105 );
    not g3038 ( n1439 , n400 );
    nor g3039 ( n1812 , n497 , n3436 );
    or g3040 ( n3722 , n509 , n1075 );
    nor g3041 ( n3789 , n275 , n2026 );
    not g3042 ( n3529 , n582 );
    nor g3043 ( n682 , n2999 , n1234 );
    nor g3044 ( n812 , n3112 , n994 );
    or g3045 ( n2707 , n245 , n3470 );
    nor g3046 ( n3588 , n1568 , n1886 );
    nor g3047 ( n253 , n2250 , n179 );
    or g3048 ( n1565 , n1053 , n1163 );
    not g3049 ( n3499 , n3050 );
    or g3050 ( n2110 , n1200 , n3665 );
    or g3051 ( n625 , n3523 , n26 );
    nor g3052 ( n666 , n3554 , n2922 );
    and g3053 ( n1381 , n846 , n435 );
    and g3054 ( n3412 , n2475 , n3289 );
    and g3055 ( n2546 , n631 , n37 );
    nor g3056 ( n1801 , n2147 , n2457 );
    and g3057 ( n3036 , n521 , n1497 );
    not g3058 ( n708 , n850 );
    or g3059 ( n3398 , n1168 , n2538 );
    nor g3060 ( n1115 , n317 , n847 );
    and g3061 ( n2135 , n3769 , n3658 );
    nor g3062 ( n2864 , n3070 , n1702 );
    nor g3063 ( n53 , n1202 , n1393 );
    nor g3064 ( n950 , n1913 , n1603 );
    or g3065 ( n880 , n1842 , n1291 );
    not g3066 ( n1230 , n1529 );
    or g3067 ( n3514 , n1748 , n3438 );
    and g3068 ( n3005 , n2588 , n1845 );
    not g3069 ( n1835 , n3026 );
    nor g3070 ( n3726 , n614 , n81 );
    nor g3071 ( n515 , n2775 , n814 );
    or g3072 ( n508 , n3344 , n316 );
    nor g3073 ( n3170 , n1472 , n2184 );
    not g3074 ( n2 , n1819 );
    nor g3075 ( n1419 , n2031 , n1129 );
    or g3076 ( n730 , n2274 , n1809 );
    nor g3077 ( n131 , n140 , n358 );
    nor g3078 ( n1367 , n1391 , n2447 );
    or g3079 ( n2116 , n1392 , n3840 );
    or g3080 ( n778 , n1206 , n2220 );
    or g3081 ( n1253 , n1646 , n1352 );
    or g3082 ( n3496 , n1818 , n1248 );
    not g3083 ( n1389 , n460 );
    and g3084 ( n1356 , n2110 , n2582 );
    nor g3085 ( n2113 , n1382 , n665 );
    and g3086 ( n2941 , n2340 , n2994 );
    or g3087 ( n182 , n3738 , n355 );
    nor g3088 ( n1789 , n833 , n1356 );
    and g3089 ( n1719 , n3365 , n1018 );
    nor g3090 ( n767 , n3672 , n640 );
    not g3091 ( n907 , n3291 );
    and g3092 ( n1311 , n1058 , n1807 );
    or g3093 ( n823 , n507 , n3034 );
    nor g3094 ( n1453 , n1707 , n519 );
    or g3095 ( n590 , n333 , n1235 );
    nor g3096 ( n125 , n3468 , n2246 );
    and g3097 ( n916 , n648 , n3793 );
    not g3098 ( n300 , n919 );
    or g3099 ( n1394 , n3699 , n1282 );
    or g3100 ( n3624 , n3063 , n1115 );
    not g3101 ( n2126 , n649 );
    or g3102 ( n3340 , n1672 , n656 );
    or g3103 ( n24 , n3732 , n1554 );
    and g3104 ( n2839 , n1339 , n315 );
    or g3105 ( n1090 , n2948 , n3187 );
    nor g3106 ( n2801 , n573 , n392 );
    not g3107 ( n1642 , n751 );
    nor g3108 ( n3444 , n389 , n1433 );
    not g3109 ( n3049 , n2616 );
    nor g3110 ( n2420 , n920 , n2595 );
    and g3111 ( n1986 , n2155 , n464 );
    and g3112 ( n2326 , n1951 , n2381 );
    or g3113 ( n1186 , n2125 , n2560 );
    nor g3114 ( n3088 , n1236 , n1883 );
    and g3115 ( n3817 , n1496 , n3389 );
    or g3116 ( n3597 , n615 , n3749 );
    nor g3117 ( n2619 , n2163 , n333 );
    or g3118 ( n124 , n2706 , n3459 );
    and g3119 ( n3363 , n3141 , n150 );
    and g3120 ( n286 , n3643 , n1070 );
    nor g3121 ( n1843 , n911 , n3245 );
    nor g3122 ( n1886 , n1620 , n3097 );
    not g3123 ( n2381 , n2985 );
    and g3124 ( n3127 , n352 , n3364 );
    or g3125 ( n2606 , n3850 , n3435 );
    nor g3126 ( n1540 , n969 , n690 );
    and g3127 ( n633 , n3111 , n3805 );
    and g3128 ( n3629 , n3355 , n150 );
    and g3129 ( n3285 , n3223 , n535 );
    nor g3130 ( n1110 , n506 , n2533 );
    nor g3131 ( n1990 , n433 , n611 );
    or g3132 ( n1272 , n1619 , n2557 );
    nor g3133 ( n2178 , n2283 , n2673 );
    or g3134 ( n1243 , n2699 , n1615 );
    or g3135 ( n2613 , n3690 , n1637 );
    nor g3136 ( n3391 , n1121 , n3803 );
    or g3137 ( n800 , n1296 , n572 );
    nor g3138 ( n1847 , n745 , n3584 );
    or g3139 ( n1067 , n2963 , n2756 );
    and g3140 ( n180 , n2236 , n263 );
    and g3141 ( n1996 , n1950 , n1860 );
    not g3142 ( n2599 , n3385 );
    or g3143 ( n2667 , n173 , n1798 );
    and g3144 ( n1616 , n3783 , n779 );
    not g3145 ( n959 , n2413 );
    nor g3146 ( n372 , n1860 , n1950 );
    or g3147 ( n865 , n1764 , n3746 );
    or g3148 ( n436 , n3461 , n180 );
    or g3149 ( n1266 , n3495 , n3033 );
    nor g3150 ( n2415 , n3189 , n3566 );
    nor g3151 ( n3443 , n3431 , n3305 );
    or g3152 ( n1733 , n1395 , n2200 );
    nor g3153 ( n1542 , n3336 , n3069 );
    not g3154 ( n738 , n2665 );
    nor g3155 ( n47 , n160 , n78 );
    nor g3156 ( n1135 , n2311 , n3583 );
    nor g3157 ( n3219 , n3756 , n1662 );
    nor g3158 ( n3469 , n2172 , n936 );
    not g3159 ( n3665 , n1374 );
    or g3160 ( n3337 , n1618 , n3036 );
    and g3161 ( n1942 , n2140 , n2472 );
    or g3162 ( n3852 , n2549 , n3655 );
    and g3163 ( n2347 , n2203 , n643 );
    or g3164 ( n1310 , n1796 , n3151 );
    and g3165 ( n3557 , n1132 , n2280 );
    or g3166 ( n3425 , n635 , n209 );
    or g3167 ( n74 , n1854 , n2976 );
    or g3168 ( n268 , n2283 , n3241 );
    nor g3169 ( n3609 , n1610 , n941 );
    and g3170 ( n641 , n3297 , n2824 );
    nor g3171 ( n1522 , n3265 , n198 );
    and g3172 ( n1390 , n3715 , n3071 );
    and g3173 ( n2313 , n1845 , n322 );
    nor g3174 ( n3759 , n561 , n2463 );
    not g3175 ( n2384 , n3693 );
    or g3176 ( n2061 , n134 , n1473 );
    not g3177 ( n136 , n2482 );
    or g3178 ( n1788 , n977 , n1584 );
    or g3179 ( n2601 , n1960 , n1980 );
    not g3180 ( n2616 , n1381 );
    not g3181 ( n3213 , n607 );
    or g3182 ( n3476 , n2726 , n1263 );
    nor g3183 ( n2505 , n496 , n2365 );
    and g3184 ( n3226 , n2775 , n2764 );
    or g3185 ( n1500 , n3502 , n1126 );
    nor g3186 ( n2128 , n657 , n2905 );
    and g3187 ( n3465 , n1544 , n1039 );
    not g3188 ( n808 , n2188 );
    nor g3189 ( n2091 , n2859 , n815 );
    or g3190 ( n3359 , n1197 , n3863 );
    not g3191 ( n893 , n298 );
    nor g3192 ( n3257 , n781 , n875 );
    and g3193 ( n156 , n239 , n3406 );
    and g3194 ( n1639 , n783 , n2032 );
    nor g3195 ( n821 , n2759 , n3077 );
    nor g3196 ( n3690 , n930 , n3090 );
    not g3197 ( n2357 , n3756 );
    nor g3198 ( n2451 , n2660 , n3057 );
    or g3199 ( n3528 , n2844 , n1223 );
    or g3200 ( n272 , n2416 , n1047 );
    and g3201 ( n2844 , n1615 , n2699 );
    not g3202 ( n1374 , n3294 );
    nor g3203 ( n1557 , n99 , n70 );
    and g3204 ( n2835 , n2069 , n3180 );
    and g3205 ( n3478 , n2559 , n2204 );
    or g3206 ( n2895 , n1062 , n807 );
    or g3207 ( n2142 , n1403 , n2593 );
    nor g3208 ( n2934 , n140 , n1191 );
    nor g3209 ( n3263 , n2427 , n143 );
    nor g3210 ( n1796 , n224 , n2114 );
    nor g3211 ( n2310 , n698 , n2190 );
    or g3212 ( n2222 , n2741 , n1205 );
    or g3213 ( n492 , n152 , n2047 );
    or g3214 ( n3348 , n3215 , n997 );
    nor g3215 ( n3043 , n2514 , n3856 );
    or g3216 ( n2021 , n3263 , n3285 );
    or g3217 ( n2132 , n1760 , n3551 );
    or g3218 ( n1831 , n26 , n2366 );
    nor g3219 ( n216 , n1071 , n2243 );
    nor g3220 ( n2922 , n3496 , n3164 );
    nor g3221 ( n179 , n1787 , n3515 );
    not g3222 ( n1866 , n2609 );
    nor g3223 ( n2246 , n1040 , n3804 );
    or g3224 ( n3491 , n3122 , n1820 );
    or g3225 ( n3463 , n636 , n2146 );
    or g3226 ( n2466 , n1596 , n1878 );
    nor g3227 ( n1968 , n2277 , n3127 );
    nor g3228 ( n137 , n2334 , n2597 );
    or g3229 ( n2851 , n688 , n3148 );
    nor g3230 ( n885 , n3440 , n1884 );
    nor g3231 ( n307 , n103 , n3842 );
    nor g3232 ( n1014 , n2885 , n1915 );
    nor g3233 ( n2717 , n1724 , n2644 );
    not g3234 ( n3748 , n560 );
    and g3235 ( n536 , n2124 , n2048 );
    nor g3236 ( n2372 , n2519 , n3217 );
    or g3237 ( n670 , n3168 , n3148 );
    nor g3238 ( n3353 , n3336 , n1906 );
    nor g3239 ( n3119 , n2838 , n136 );
    nor g3240 ( n57 , n2121 , n2298 );
    nor g3241 ( n572 , n1036 , n1994 );
    nor g3242 ( n3028 , n2733 , n3652 );
    not g3243 ( n3550 , n2711 );
    or g3244 ( n1456 , n374 , n1321 );
    or g3245 ( n1312 , n863 , n2850 );
    not g3246 ( n3834 , n1074 );
    not g3247 ( n3346 , n959 );
    not g3248 ( n868 , n2767 );
    nor g3249 ( n3679 , n3513 , n145 );
    not g3250 ( n655 , n2397 );
    or g3251 ( n3456 , n1503 , n3579 );
    and g3252 ( n2331 , n2649 , n3153 );
    and g3253 ( n1951 , n3000 , n1396 );
    or g3254 ( n1690 , n3753 , n415 );
    nor g3255 ( n3038 , n1058 , n1807 );
    nor g3256 ( n3421 , n2588 , n1845 );
    nor g3257 ( n3845 , n1908 , n382 );
    and g3258 ( n2527 , n2983 , n3003 );
    nor g3259 ( n2161 , n649 , n2243 );
    and g3260 ( n2720 , n1078 , n2379 );
    not g3261 ( n2597 , n1190 );
    nor g3262 ( n3711 , n1837 , n3777 );
    nor g3263 ( n2054 , n364 , n2314 );
    not g3264 ( n95 , n1295 );
    nor g3265 ( n9 , n232 , n322 );
    and g3266 ( n218 , n3135 , n2174 );
    or g3267 ( n0 , n1247 , n1971 );
    nor g3268 ( n1197 , n2944 , n136 );
    nor g3269 ( n539 , n1514 , n512 );
    or g3270 ( n219 , n676 , n2326 );
    nor g3271 ( n1160 , n368 , n2633 );
    or g3272 ( n181 , n53 , n291 );
    or g3273 ( n487 , n1737 , n2109 );
    or g3274 ( n1765 , n1509 , n737 );
    or g3275 ( n1219 , n3397 , n3254 );
    nor g3276 ( n265 , n2226 , n3217 );
    not g3277 ( n292 , n2732 );
    nor g3278 ( n2972 , n3248 , n896 );
    and g3279 ( n1649 , n1889 , n3027 );
    nor g3280 ( n952 , n838 , n1059 );
    nor g3281 ( n1853 , n2812 , n1137 );
    nor g3282 ( n1879 , n2939 , n2657 );
    and g3283 ( n254 , n1610 , n941 );
    or g3284 ( n3185 , n3012 , n3073 );
    nor g3285 ( n3780 , n1692 , n2026 );
    or g3286 ( n2360 , n3399 , n1147 );
    nor g3287 ( n3613 , n2090 , n1977 );
    or g3288 ( n45 , n571 , n1929 );
    and g3289 ( n2724 , n3375 , n1733 );
    or g3290 ( n2305 , n1902 , n107 );
    nor g3291 ( n65 , n3307 , n2350 );
    and g3292 ( n2842 , n2455 , n3048 );
    nor g3293 ( n3304 , n1819 , n1673 );
    or g3294 ( n2834 , n2043 , n2105 );
    or g3295 ( n3317 , n230 , n3608 );
    and g3296 ( n3727 , n3022 , n936 );
    and g3297 ( n2460 , n2474 , n383 );
    not g3298 ( n2368 , n1550 );
    not g3299 ( n456 , n3807 );
    or g3300 ( n1251 , n3539 , n3746 );
    nor g3301 ( n1833 , n3442 , n936 );
    and g3302 ( n2554 , n696 , n2568 );
    and g3303 ( n3275 , n1731 , n968 );
    and g3304 ( n237 , n1260 , n2041 );
    or g3305 ( n3301 , n3450 , n933 );
    or g3306 ( n1435 , n3558 , n2325 );
    or g3307 ( n52 , n3134 , n1604 );
    nor g3308 ( n454 , n1680 , n1673 );
    and g3309 ( n165 , n905 , n2757 );
    nor g3310 ( n305 , n2474 , n847 );
    nor g3311 ( n1022 , n2493 , n1698 );
    nor g3312 ( n1318 , n674 , n2263 );
    or g3313 ( n2005 , n3646 , n1263 );
    not g3314 ( n1934 , n1669 );
    nor g3315 ( n1564 , n3163 , n1386 );
    or g3316 ( n2046 , n1270 , n3286 );
    and g3317 ( n3858 , n2738 , n379 );
    not g3318 ( n2200 , n3625 );
    nor g3319 ( n2044 , n178 , n1802 );
    or g3320 ( n1342 , n1550 , n1554 );
    nor g3321 ( n2412 , n671 , n2813 );
    not g3322 ( n691 , n2049 );
    or g3323 ( n2058 , n2004 , n1985 );
    nor g3324 ( n884 , n980 , n746 );
    nor g3325 ( n422 , n1228 , n576 );
    nor g3326 ( n2176 , n844 , n2421 );
    nor g3327 ( n3128 , n2180 , n358 );
    and g3328 ( n1746 , n1868 , n2952 );
    and g3329 ( n1028 , n1285 , n1478 );
    not g3330 ( n2992 , n404 );
    nor g3331 ( n3828 , n866 , n1302 );
    and g3332 ( n1807 , n831 , n1005 );
    or g3333 ( n1851 , n1055 , n537 );
    nor g3334 ( n785 , n3611 , n6 );
    nor g3335 ( n2160 , n1076 , n3817 );
    or g3336 ( n1678 , n2649 , n1291 );
    nor g3337 ( n2587 , n2494 , n226 );
    or g3338 ( n2622 , n2234 , n1334 );
    or g3339 ( n1695 , n1415 , n2682 );
    nor g3340 ( n3453 , n3092 , n2252 );
    not g3341 ( n2832 , n3133 );
    and g3342 ( n2783 , n3513 , n75 );
    or g3343 ( n2235 , n2013 , n2717 );
    not g3344 ( n3058 , n773 );
    nor g3345 ( n1590 , n2816 , n2216 );
    nor g3346 ( n3518 , n606 , n2336 );
    nor g3347 ( n2234 , n1285 , n1673 );
    nor g3348 ( n805 , n3340 , n3559 );
    or g3349 ( n3247 , n945 , n633 );
    or g3350 ( n1652 , n1318 , n999 );
    or g3351 ( n1790 , n993 , n235 );
endmodule
