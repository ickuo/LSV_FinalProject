module top( n23 , n26 , n29 , n32 , n41 , n44 , n54 , n58 , n59 , 
n61 , n64 , n65 , n77 , n80 , n83 , n86 , n97 , n99 , n102 , 
n118 , n129 , n144 , n163 , n177 , n184 , n194 , n205 , n209 , n212 , 
n220 , n221 , n226 , n228 , n231 , n233 , n241 , n243 , n247 , n257 , 
n261 , n263 , n274 , n277 , n280 , n282 , n287 , n300 , n305 , n312 , 
n313 , n317 , n320 , n323 , n326 );
    input n23 , n26 , n54 , n58 , n59 , n61 , n64 , n65 , n77 , 
n86 , n97 , n102 , n118 , n129 , n144 , n184 , n205 , n209 , n220 , 
n241 , n257 , n274 , n277 , n280 , n305 , n312 , n313 , n317 , n323 ;
    output n29 , n32 , n41 , n44 , n80 , n83 , n99 , n163 , n177 , 
n194 , n212 , n221 , n226 , n228 , n231 , n233 , n243 , n247 , n261 , 
n263 , n282 , n287 , n300 , n320 , n326 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , 
n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , 
n19 , n20 , n21 , n22 , n24 , n25 , n27 , n28 , n30 , n31 , 
n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n42 , n43 , 
n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n55 , 
n56 , n57 , n60 , n62 , n63 , n66 , n67 , n68 , n69 , n70 , 
n71 , n72 , n73 , n74 , n75 , n76 , n78 , n79 , n81 , n82 , 
n84 , n85 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , 
n95 , n96 , n98 , n100 , n101 , n103 , n104 , n105 , n106 , n107 , 
n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , 
n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , 
n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
n140 , n141 , n142 , n143 , n145 , n146 , n147 , n148 , n149 , n150 , 
n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
n161 , n162 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , 
n172 , n173 , n174 , n175 , n176 , n178 , n179 , n180 , n181 , n182 , 
n183 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , 
n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , 
n206 , n207 , n208 , n210 , n211 , n213 , n214 , n215 , n216 , n217 , 
n218 , n219 , n222 , n223 , n224 , n225 , n227 , n229 , n230 , n232 , 
n234 , n235 , n236 , n237 , n238 , n239 , n240 , n242 , n244 , n245 , 
n246 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , 
n258 , n259 , n260 , n262 , n264 , n265 , n266 , n267 , n268 , n269 , 
n270 , n271 , n272 , n273 , n275 , n276 , n278 , n279 , n281 , n283 , 
n284 , n285 , n286 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , 
n295 , n296 , n297 , n298 , n299 , n301 , n302 , n303 , n304 , n306 , 
n307 , n308 , n309 , n310 , n311 , n314 , n315 , n316 , n318 , n319 , 
n321 , n322 , n324 , n325 , n327 , n328 , n329 , n330 , n331 , n332 , 
n333 ;
    not g0 ( n95 , n64 );
    and g1 ( n249 , n203 , n276 );
    not g2 ( n154 , n153 );
    and g3 ( n75 , n191 , n118 );
    not g4 ( n202 , n122 );
    or g5 ( n181 , n20 , n170 );
    and g6 ( n169 , n327 , n254 );
    nor g7 ( n248 , n186 , n92 );
    nor g8 ( n135 , n122 , n66 );
    not g9 ( n224 , n124 );
    xnor g10 ( n1 , n330 , n34 );
    nor g11 ( n68 , n114 , n324 );
    not g12 ( n128 , n183 );
    not g13 ( n69 , n111 );
    xnor g14 ( n100 , n275 , n201 );
    nor g15 ( n288 , n309 , n116 );
    and g16 ( n6 , n253 , n217 );
    xnor g17 ( n138 , n7 , n317 );
    or g18 ( n290 , n43 , n146 );
    not g19 ( n306 , n120 );
    not g20 ( n9 , n53 );
    or g21 ( n289 , n187 , n319 );
    nor g22 ( n252 , n72 , n51 );
    not g23 ( n246 , n57 );
    or g24 ( n218 , n13 , n145 );
    or g25 ( n67 , n130 , n230 );
    not g26 ( n318 , n284 );
    not g27 ( n254 , n111 );
    xnor g28 ( n127 , n211 , n294 );
    and g29 ( n255 , n179 , n217 );
    or g30 ( n24 , n95 , n333 );
    xnor g31 ( n83 , n269 , n58 );
    not g32 ( n158 , n206 );
    not g33 ( n12 , n183 );
    and g34 ( n21 , n229 , n241 );
    xnor g35 ( n101 , n236 , n199 );
    or g36 ( n258 , n75 , n128 );
    xor g37 ( n82 , n199 , n129 );
    not g38 ( n322 , n54 );
    and g39 ( n162 , n249 , n76 );
    and g40 ( n36 , n133 , n175 );
    or g41 ( n32 , n140 , n161 );
    and g42 ( n213 , n239 , n257 );
    nor g43 ( n271 , n323 , n45 );
    or g44 ( n329 , n323 , n131 );
    and g45 ( n321 , n250 , n53 );
    or g46 ( n98 , n36 , n295 );
    not g47 ( n132 , n146 );
    xnor g48 ( n103 , n174 , n241 );
    not g49 ( n108 , n72 );
    xnor g50 ( n94 , n129 , n220 );
    and g51 ( n57 , n55 , n39 );
    and g52 ( n89 , n81 , n23 );
    and g53 ( n113 , n52 , n244 );
    not g54 ( n307 , n56 );
    not g55 ( n333 , n209 );
    and g56 ( n215 , n9 , n67 );
    and g57 ( n314 , n327 , n108 );
    and g58 ( n42 , n35 , n250 );
    xnor g59 ( n90 , n272 , n102 );
    or g60 ( n96 , n256 , n264 );
    xnor g61 ( n253 , n138 , n127 );
    or g62 ( n29 , n157 , n259 );
    not g63 ( n141 , n274 );
    not g64 ( n70 , n214 );
    not g65 ( n8 , n292 );
    nor g66 ( n286 , n110 , n244 );
    and g67 ( n270 , n186 , n164 );
    not g68 ( n332 , n257 );
    not g69 ( n93 , n139 );
    or g70 ( n14 , n176 , n158 );
    or g71 ( n40 , n257 , n88 );
    and g72 ( n30 , n242 , n179 );
    and g73 ( n188 , n88 , n257 );
    xnor g74 ( n179 , n207 , n101 );
    xnor g75 ( n228 , n281 , n280 );
    not g76 ( n239 , n97 );
    not g77 ( n204 , n154 );
    xnor g78 ( n263 , n162 , n61 );
    and g79 ( n256 , n2 , n216 );
    and g80 ( n130 , n74 , n213 );
    or g81 ( n25 , n100 , n250 );
    xnor g82 ( n27 , n129 , n277 );
    nor g83 ( n200 , n150 , n70 );
    or g84 ( n208 , n227 , n301 );
    or g85 ( n56 , n205 , n182 );
    xnor g86 ( n315 , n331 , n102 );
    and g87 ( n311 , n39 , n305 );
    or g88 ( n136 , n311 , n91 );
    not g89 ( n164 , n125 );
    nor g90 ( n259 , n188 , n1 );
    nor g91 ( n268 , n257 , n313 );
    or g92 ( n92 , n51 , n62 );
    not g93 ( n49 , n266 );
    or g94 ( n237 , n42 , n98 );
    xnor g95 ( n149 , n315 , n48 );
    or g96 ( n242 , n234 , n128 );
    not g97 ( n229 , n117 );
    or g98 ( n143 , n313 , n187 );
    and g99 ( n104 , n2 , n189 );
    not g100 ( n13 , n316 );
    not g101 ( n55 , n79 );
    not g102 ( n73 , n270 );
    xnor g103 ( n151 , n280 , n129 );
    and g104 ( n244 , n141 , n257 );
    and g105 ( n173 , n227 , n189 );
    and g106 ( n227 , n119 , n172 );
    or g107 ( n166 , n257 , n322 );
    xnor g108 ( n222 , n27 , n90 );
    nor g109 ( n150 , n69 , n175 );
    and g110 ( n210 , n289 , n191 );
    nor g111 ( n109 , n305 , n253 );
    xnor g112 ( n331 , n144 , n317 );
    and g113 ( n310 , n134 , n250 );
    xnor g114 ( n172 , n289 , n271 );
    or g115 ( n111 , n164 , n103 );
    nor g116 ( n330 , n213 , n82 );
    not g117 ( n153 , n16 );
    and g118 ( n20 , n328 , n250 );
    or g119 ( n170 , n281 , n296 );
    xnor g120 ( n326 , n286 , n297 );
    or g121 ( n221 , n257 , n290 );
    and g122 ( n299 , n190 , n332 );
    xnor g123 ( n22 , n63 , n118 );
    xnor g124 ( n197 , n0 , n61 );
    not g125 ( n147 , n293 );
    not g126 ( n117 , n56 );
    or g127 ( n275 , n95 , n38 );
    nor g128 ( n78 , n275 , n202 );
    not g129 ( n39 , n307 );
    or g130 ( n301 , n192 , n46 );
    not g131 ( n230 , n13 );
    nor g132 ( n232 , n71 , n126 );
    not g133 ( n5 , n67 );
    and g134 ( n293 , n270 , n9 );
    and g135 ( n134 , n120 , n17 );
    or g136 ( n276 , n113 , n316 );
    xnor g137 ( n251 , n151 , n65 );
    and g138 ( n155 , n136 , n253 );
    and g139 ( n235 , n133 , n69 );
    not g140 ( n175 , n72 );
    and g141 ( n133 , n15 , n321 );
    and g142 ( n269 , n248 , n125 );
    nor g143 ( n161 , n45 , n156 );
    not g144 ( n183 , n292 );
    or g145 ( n62 , n206 , n283 );
    not g146 ( n266 , n172 );
    or g147 ( n279 , n162 , n137 );
    or g148 ( n84 , n303 , n194 );
    xnor g149 ( n260 , n40 , n65 );
    or g150 ( n178 , n121 , n96 );
    or g151 ( n296 , n269 , n178 );
    or g152 ( n212 , n165 , n18 );
    and g153 ( n291 , n249 , n265 );
    or g154 ( n226 , n68 , n47 );
    xnor g155 ( n80 , n310 , n144 );
    xnor g156 ( n247 , n169 , n312 );
    and g157 ( n234 , n33 , n26 );
    and g158 ( n174 , n50 , n19 );
    and g159 ( n316 , n193 , n182 );
    and g160 ( n193 , n284 , n205 );
    not g161 ( n240 , n306 );
    xnor g162 ( n297 , n238 , n299 );
    xnor g163 ( n50 , n107 , n222 );
    or g164 ( n264 , n310 , n84 );
    not g165 ( n19 , n323 );
    or g166 ( n72 , n224 , n309 );
    and g167 ( n165 , n273 , n168 );
    xnor g168 ( n163 , n256 , n317 );
    nor g169 ( n46 , n158 , n304 );
    nor g170 ( n110 , n54 , n332 );
    xnor g171 ( n148 , n139 , n166 );
    xnor g172 ( n0 , n312 , n59 );
    not g173 ( n124 , n125 );
    xnor g174 ( n233 , n314 , n59 );
    xnor g175 ( n45 , n106 , n148 );
    or g176 ( n114 , n325 , n118 );
    xnor g177 ( n125 , n6 , n305 );
    xnor g178 ( n282 , n36 , n277 );
    not g179 ( n285 , n323 );
    xnor g180 ( n261 , n295 , n129 );
    not g181 ( n225 , n215 );
    not g182 ( n219 , n313 );
    xnor g183 ( n123 , n197 , n236 );
    and g184 ( n303 , n173 , n204 );
    or g185 ( n41 , n105 , n30 );
    nor g186 ( n192 , n49 , n14 );
    xnor g187 ( n106 , n280 , n58 );
    not g188 ( n91 , n8 );
    xnor g189 ( n122 , n251 , n10 );
    nor g190 ( n17 , n5 , n147 );
    nor g191 ( n81 , n131 , n257 );
    and g192 ( n105 , n60 , n112 );
    and g193 ( n160 , n203 , n189 );
    or g194 ( n167 , n21 , n91 );
    and g195 ( n120 , n262 , n22 );
    or g196 ( n190 , n235 , n180 );
    and g197 ( n265 , n293 , n204 );
    or g198 ( n137 , n314 , n237 );
    not g199 ( n191 , n307 );
    not g200 ( n131 , n209 );
    or g201 ( n180 , n291 , n152 );
    xnor g202 ( n16 , n255 , n26 );
    or g203 ( n308 , n188 , n213 );
    not g204 ( n28 , n321 );
    not g205 ( n187 , n86 );
    nor g206 ( n156 , n210 , n292 );
    not g207 ( n298 , n276 );
    and g208 ( n327 , n249 , n214 );
    and g209 ( n267 , n198 , n77 );
    and g210 ( n272 , n268 , n77 );
    not g211 ( n2 , n306 );
    or g212 ( n284 , n219 , n333 );
    xnor g213 ( n211 , n58 , n129 );
    and g214 ( n302 , n275 , n33 );
    nor g215 ( n216 , n111 , n51 );
    xnor g216 ( n287 , n291 , n65 );
    not g217 ( n325 , n57 );
    nor g218 ( n74 , n285 , n318 );
    or g219 ( n283 , n87 , n266 );
    or g220 ( n51 , n5 , n28 );
    and g221 ( n3 , n57 , n109 );
    nor g222 ( n201 , n323 , n122 );
    and g223 ( n31 , n232 , n230 );
    xnor g224 ( n139 , n195 , n123 );
    and g225 ( n47 , n258 , n324 );
    and g226 ( n140 , n60 , n196 );
    xnor g227 ( n236 , n94 , n277 );
    not g228 ( n33 , n117 );
    not g229 ( n53 , n100 );
    xnor g230 ( n207 , n223 , n61 );
    and g231 ( n319 , n219 , n19 );
    not g232 ( n214 , n25 );
    nor g233 ( n168 , n241 , n50 );
    xnor g234 ( n294 , n94 , n312 );
    xnor g235 ( n107 , n85 , n59 );
    and g236 ( n34 , n181 , n182 );
    nor g237 ( n142 , n304 , n245 );
    not g238 ( n88 , n184 );
    xnor g239 ( n48 , n85 , n197 );
    not g240 ( n115 , n227 );
    xnor g241 ( n99 , n235 , n220 );
    or g242 ( n146 , n181 , n190 );
    and g243 ( n37 , n273 , n78 );
    or g244 ( n79 , n159 , n132 );
    xnor g245 ( n177 , n42 , n129 );
    or g246 ( n238 , n244 , n93 );
    xnor g247 ( n320 , n20 , n129 );
    nor g248 ( n223 , n257 , n143 );
    not g249 ( n60 , n325 );
    and g250 ( n4 , n218 , n71 );
    or g251 ( n243 , n37 , n135 );
    not g252 ( n217 , n323 );
    and g253 ( n295 , n288 , n224 );
    nor g254 ( n126 , n120 , n208 );
    or g255 ( n116 , n25 , n11 );
    nor g256 ( n112 , n26 , n179 );
    not g257 ( n198 , n319 );
    not g258 ( n186 , n103 );
    not g259 ( n206 , n22 );
    and g260 ( n157 , n1 , n308 );
    xnor g261 ( n324 , n260 , n149 );
    or g262 ( n231 , n3 , n155 );
    not g263 ( n273 , n246 );
    nor g264 ( n262 , n176 , n304 );
    nor g265 ( n35 , n147 , n11 );
    nor g266 ( n278 , n225 , n62 );
    nor g267 ( n196 , n289 , n171 );
    and g268 ( n189 , n108 , n215 );
    xnor g269 ( n199 , n85 , n315 );
    and g270 ( n121 , n240 , n252 );
    xnor g271 ( n300 , n121 , n102 );
    not g272 ( n309 , n103 );
    xnor g273 ( n10 , n89 , n144 );
    not g274 ( n182 , n257 );
    xnor g275 ( n195 , n129 , n65 );
    and g276 ( n176 , n329 , n23 );
    not g277 ( n15 , n11 );
    or g278 ( n11 , n298 , n115 );
    nor g279 ( n52 , n159 , n318 );
    buf g280 ( n250 , n16 );
    not g281 ( n171 , n45 );
    not g282 ( n38 , n329 );
    nor g283 ( n145 , n265 , n185 );
    and g284 ( n281 , n160 , n250 );
    nor g285 ( n66 , n302 , n12 );
    xnor g286 ( n44 , n303 , n129 );
    nor g287 ( n7 , n257 , n24 );
    not g288 ( n203 , n62 );
    and g289 ( n63 , n324 , n285 );
    or g290 ( n87 , n267 , n176 );
    and g291 ( n76 , n321 , n270 );
    or g292 ( n185 , n200 , n76 );
    or g293 ( n304 , n267 , n49 );
    or g294 ( n71 , n73 , n70 );
    and g295 ( n194 , n104 , n153 );
    and g296 ( n292 , n79 , n229 );
    or g297 ( n152 , n169 , n279 );
    or g298 ( n43 , n31 , n142 );
    xnor g299 ( n85 , n151 , n58 );
    not g300 ( n159 , n323 );
    nor g301 ( n119 , n267 , n14 );
    or g302 ( n245 , n14 , n4 );
    and g303 ( n328 , n278 , n254 );
    and g304 ( n18 , n167 , n50 );
endmodule
