module top( n3 , n10 , n12 , n21 , n24 , n25 , n26 , n27 , n28 , 
n29 , n31 , n32 , n37 , n41 , n45 , n46 , n47 , n48 , n51 , 
n52 , n54 , n55 , n60 , n62 , n64 , n70 , n76 , n77 , n83 , 
n84 , n91 , n96 , n98 , n102 , n103 , n106 , n118 , n127 , n129 , 
n139 , n140 , n143 , n153 , n155 , n160 , n163 , n164 , n168 , n169 , 
n171 , n173 , n176 , n180 , n185 , n186 , n187 , n191 , n192 , n194 , 
n197 , n198 , n202 , n210 , n216 , n220 , n221 , n222 , n235 , n242 , 
n243 , n246 , n251 , n254 );
    input n10 , n21 , n24 , n29 , n37 , n45 , n46 , n47 , n48 , 
n51 , n52 , n55 , n76 , n77 , n84 , n102 , n106 , n127 , n140 , 
n143 , n155 , n160 , n164 , n168 , n171 , n173 , n176 , n180 , n185 , 
n186 , n197 , n198 , n210 , n216 , n220 , n221 , n222 , n242 , n243 , 
n246 , n251 ;
    output n3 , n12 , n25 , n26 , n27 , n28 , n31 , n32 , n41 , 
n54 , n60 , n62 , n64 , n70 , n83 , n91 , n96 , n98 , n103 , 
n118 , n129 , n139 , n153 , n163 , n169 , n187 , n191 , n192 , n194 , 
n202 , n235 , n254 ;
    wire n0 , n1 , n2 , n4 , n5 , n6 , n7 , n8 , n9 , 
n11 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n22 , 
n23 , n30 , n33 , n34 , n35 , n36 , n38 , n39 , n40 , n42 , 
n43 , n44 , n49 , n50 , n53 , n56 , n57 , n58 , n59 , n61 , 
n63 , n65 , n66 , n67 , n68 , n69 , n71 , n72 , n73 , n74 , 
n75 , n78 , n79 , n80 , n81 , n82 , n85 , n86 , n87 , n88 , 
n89 , n90 , n92 , n93 , n94 , n95 , n97 , n99 , n100 , n101 , 
n104 , n105 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , 
n115 , n116 , n117 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , 
n126 , n128 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , 
n138 , n141 , n142 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
n151 , n152 , n154 , n156 , n157 , n158 , n159 , n161 , n162 , n165 , 
n166 , n167 , n170 , n172 , n174 , n175 , n177 , n178 , n179 , n181 , 
n182 , n183 , n184 , n188 , n189 , n190 , n193 , n195 , n196 , n199 , 
n200 , n201 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n211 , 
n212 , n213 , n214 , n215 , n217 , n218 , n219 , n223 , n224 , n225 , 
n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n236 , 
n237 , n238 , n239 , n240 , n241 , n244 , n245 , n247 , n248 , n249 , 
n250 , n252 , n253 , n255 ;
    nor g0 ( n19 , n23 , n156 );
    or g1 ( n154 , n74 , n205 );
    xnor g2 ( n163 , n59 , n197 );
    xnor g3 ( n217 , n21 , n168 );
    xnor g4 ( n80 , n29 , n164 );
    not g5 ( n209 , n220 );
    xnor g6 ( n137 , n218 , n231 );
    or g7 ( n122 , n97 , n78 );
    or g8 ( n88 , n97 , n109 );
    xnor g9 ( n56 , n140 , n52 );
    xnor g10 ( n73 , n127 , n106 );
    xor g11 ( n240 , n241 , n128 );
    or g12 ( n114 , n199 , n39 );
    xnor g13 ( n177 , n84 , n171 );
    or g14 ( n223 , n225 , n142 );
    xnor g15 ( n194 , n250 , n51 );
    or g16 ( n34 , n119 , n94 );
    or g17 ( n149 , n4 , n105 );
    nor g18 ( n42 , n133 , n232 );
    xnor g19 ( n26 , n117 , n29 );
    xnor g20 ( n207 , n106 , n102 );
    xnor g21 ( n200 , n189 , n30 );
    xnor g22 ( n75 , n196 , n217 );
    xnor g23 ( n167 , n197 , n173 );
    or g24 ( n5 , n195 , n147 );
    nor g25 ( n238 , n240 , n18 );
    or g26 ( n59 , n188 , n78 );
    xnor g27 ( n103 , n122 , n55 );
    xnor g28 ( n241 , n93 , n151 );
    nor g29 ( n232 , n199 , n239 );
    xnor g30 ( n64 , n206 , n164 );
    xnor g31 ( n255 , n246 , n222 );
    xnor g32 ( n17 , n80 , n207 );
    or g33 ( n119 , n175 , n124 );
    or g34 ( n205 , n114 , n85 );
    xnor g35 ( n22 , n249 , n131 );
    not g36 ( n33 , n45 );
    xnor g37 ( n71 , n253 , n162 );
    not g38 ( n74 , n124 );
    xnor g39 ( n187 , n53 , n46 );
    or g40 ( n43 , n159 , n252 );
    xnor g41 ( n245 , n55 , n164 );
    or g42 ( n0 , n175 , n205 );
    xnor g43 ( n138 , n171 , n10 );
    xnor g44 ( n136 , n46 , n246 );
    xnor g45 ( n254 , n63 , n127 );
    not g46 ( n40 , n77 );
    xnor g47 ( n86 , n51 , n76 );
    or g48 ( n67 , n172 , n149 );
    nor g49 ( n135 , n199 , n215 );
    xnor g50 ( n9 , n140 , n198 );
    or g51 ( n94 , n227 , n8 );
    xnor g52 ( n233 , n245 , n167 );
    xnor g53 ( n196 , n221 , n29 );
    xnor g54 ( n115 , n251 , n51 );
    nor g55 ( n183 , n19 , n135 );
    xnor g56 ( n208 , n201 , n17 );
    or g57 ( n63 , n97 , n34 );
    or g58 ( n95 , n33 , n147 );
    xnor g59 ( n235 , n14 , n10 );
    or g60 ( n134 , n188 , n109 );
    or g61 ( n190 , n61 , n240 );
    xnor g62 ( n184 , n228 , n146 );
    or g63 ( n224 , n6 , n126 );
    or g64 ( n179 , n188 , n11 );
    nor g65 ( n133 , n199 , n89 );
    xnor g66 ( n91 , n203 , n84 );
    or g67 ( n18 , n6 , n126 );
    xnor g68 ( n92 , n251 , n24 );
    xnor g69 ( n170 , n100 , n226 );
    or g70 ( n142 , n23 , n229 );
    not g71 ( n174 , n126 );
    xnor g72 ( n38 , n52 , n186 );
    or g73 ( n165 , n141 , n8 );
    xnor g74 ( n25 , n101 , n76 );
    xnor g75 ( n54 , n237 , n47 );
    xor g76 ( n126 , n71 , n58 );
    xnor g77 ( n12 , n111 , n198 );
    xnor g78 ( n249 , n168 , n173 );
    and g79 ( n8 , n42 , n183 );
    xnor g80 ( n228 , n198 , n186 );
    or g81 ( n145 , n141 , n8 );
    xnor g82 ( n153 , n154 , n24 );
    or g83 ( n182 , n193 , n147 );
    or g84 ( n253 , n40 , n147 );
    not g85 ( n248 , n240 );
    xnor g86 ( n110 , n121 , n226 );
    xnor g87 ( n58 , n138 , n255 );
    or g88 ( n227 , n172 , n126 );
    xnor g89 ( n32 , n116 , n221 );
    xnor g90 ( n128 , n9 , n115 );
    and g91 ( n72 , n61 , n211 );
    or g92 ( n225 , n1 , n39 );
    and g93 ( n81 , n61 , n158 );
    nor g94 ( n213 , n238 , n81 );
    or g95 ( n7 , n174 , n108 );
    and g96 ( n211 , n172 , n248 );
    xnor g97 ( n178 , n127 , n210 );
    or g98 ( n166 , n188 , n34 );
    xnor g99 ( n226 , n92 , n136 );
    or g100 ( n4 , n1 , n43 );
    or g101 ( n78 , n190 , n145 );
    not g102 ( n193 , n216 );
    xnor g103 ( n68 , n233 , n148 );
    or g104 ( n53 , n172 , n205 );
    xnor g105 ( n96 , n66 , n222 );
    or g106 ( n161 , n209 , n147 );
    buf g107 ( n97 , n137 );
    or g108 ( n105 , n23 , n229 );
    or g109 ( n212 , n159 , n11 );
    xnor g110 ( n146 , n155 , n10 );
    xnor g111 ( n131 , n185 , n47 );
    or g112 ( n49 , n172 , n223 );
    not g113 ( n188 , n252 );
    or g114 ( n89 , n252 , n23 );
    xnor g115 ( n27 , n0 , n251 );
    not g116 ( n159 , n112 );
    or g117 ( n237 , n159 , n109 );
    or g118 ( n14 , n174 , n149 );
    or g119 ( n156 , n252 , n112 );
    or g120 ( n104 , n82 , n147 );
    xnor g121 ( n189 , n84 , n155 );
    not g122 ( n23 , n137 );
    xnor g123 ( n214 , n24 , n76 );
    or g124 ( n157 , n1 , n34 );
    or g125 ( n250 , n175 , n223 );
    xor g126 ( n252 , n65 , n20 );
    or g127 ( n203 , n172 , n108 );
    or g128 ( n66 , n174 , n223 );
    xnor g129 ( n219 , n95 , n113 );
    or g130 ( n152 , n74 , n240 );
    or g131 ( n111 , n248 , n149 );
    xnor g132 ( n87 , n148 , n130 );
    xnor g133 ( n20 , n144 , n35 );
    not g134 ( n247 , n243 );
    or g135 ( n50 , n174 , n205 );
    xor g136 ( n112 , n219 , n22 );
    not g137 ( n147 , n160 );
    xnor g138 ( n231 , n13 , n178 );
    xnor g139 ( n65 , n104 , n110 );
    xnor g140 ( n129 , n69 , n173 );
    xnor g141 ( n123 , n176 , n47 );
    xnor g142 ( n144 , n21 , n197 );
    or g143 ( n36 , n227 , n8 );
    xnor g144 ( n148 , n57 , n123 );
    xnor g145 ( n100 , n56 , n177 );
    xnor g146 ( n236 , n242 , n185 );
    not g147 ( n61 , n124 );
    or g148 ( n206 , n1 , n78 );
    not g149 ( n175 , n240 );
    xnor g150 ( n70 , n244 , n102 );
    xnor g151 ( n41 , n50 , n246 );
    or g152 ( n234 , n247 , n147 );
    xnor g153 ( n31 , n157 , n106 );
    xnor g154 ( n202 , n88 , n210 );
    xnor g155 ( n3 , n150 , n140 );
    xnor g156 ( n15 , n184 , n121 );
    or g157 ( n150 , n175 , n108 );
    xnor g158 ( n113 , n184 , n100 );
    xnor g159 ( n169 , n166 , n242 );
    not g160 ( n195 , n37 );
    buf g161 ( n1 , n208 );
    or g162 ( n215 , n23 , n112 );
    or g163 ( n117 , n1 , n11 );
    or g164 ( n101 , n61 , n223 );
    xnor g165 ( n151 , n75 , n130 );
    xnor g166 ( n192 , n134 , n176 );
    xnor g167 ( n132 , n182 , n68 );
    or g168 ( n69 , n159 , n78 );
    or g169 ( n11 , n99 , n165 );
    not g170 ( n172 , n6 );
    or g171 ( n244 , n1 , n109 );
    or g172 ( n39 , n188 , n112 );
    xnor g173 ( n191 , n181 , n185 );
    xnor g174 ( n62 , n7 , n171 );
    or g175 ( n44 , n74 , n108 );
    or g176 ( n116 , n97 , n11 );
    xnor g177 ( n218 , n234 , n170 );
    not g178 ( n199 , n208 );
    xnor g179 ( n130 , n73 , n236 );
    xnor g180 ( n162 , n233 , n75 );
    xnor g181 ( n60 , n44 , n52 );
    xnor g182 ( n120 , n5 , n87 );
    or g183 ( n85 , n97 , n229 );
    or g184 ( n109 , n152 , n36 );
    xor g185 ( n6 , n120 , n200 );
    nor g186 ( n79 , n72 , n90 );
    xnor g187 ( n83 , n179 , n21 );
    and g188 ( n158 , n248 , n174 );
    and g189 ( n229 , n79 , n213 );
    or g190 ( n2 , n97 , n229 );
    or g191 ( n125 , n199 , n43 );
    xnor g192 ( n204 , n143 , n222 );
    xnor g193 ( n230 , n38 , n214 );
    xnor g194 ( n35 , n242 , n176 );
    xnor g195 ( n28 , n212 , n168 );
    xnor g196 ( n139 , n49 , n143 );
    xnor g197 ( n121 , n86 , n204 );
    xnor g198 ( n57 , n210 , n102 );
    not g199 ( n82 , n48 );
    or g200 ( n99 , n248 , n124 );
    not g201 ( n107 , n180 );
    xnor g202 ( n30 , n46 , n143 );
    or g203 ( n108 , n125 , n2 );
    xnor g204 ( n118 , n67 , n155 );
    or g205 ( n93 , n107 , n147 );
    xor g206 ( n124 , n132 , n230 );
    xnor g207 ( n98 , n16 , n186 );
    or g208 ( n141 , n174 , n6 );
    or g209 ( n16 , n74 , n149 );
    nor g210 ( n90 , n124 , n224 );
    xnor g211 ( n13 , n221 , n55 );
    or g212 ( n181 , n159 , n34 );
    or g213 ( n239 , n252 , n112 );
    xnor g214 ( n201 , n161 , n15 );
endmodule
