module top( n0 , n2 , n3 , n5 , n6 , n8 , n11 , n12 , n14 , 
n18 , n19 , n27 , n28 , n32 , n35 , n38 , n40 , n42 , n43 , 
n51 , n54 , n55 , n56 , n57 , n59 , n60 , n61 , n64 , n65 , 
n73 , n76 , n78 , n79 , n80 , n86 , n93 , n94 , n104 , n106 , 
n108 , n110 , n113 , n114 , n115 , n117 , n118 , n119 , n120 , n124 , 
n126 , n127 , n129 , n130 , n133 , n137 , n138 , n142 , n143 , n147 , 
n151 , n154 , n157 , n162 , n166 , n168 , n169 , n171 , n174 , n178 , 
n181 , n182 , n184 , n185 , n188 , n196 , n200 , n202 , n203 , n205 , 
n210 , n211 , n213 , n215 , n216 , n217 , n218 , n219 , n220 , n227 , 
n229 , n230 , n231 , n238 , n242 , n248 , n249 , n250 , n252 , n257 , 
n259 , n260 , n266 , n268 , n269 , n276 , n278 , n280 , n282 , n291 , 
n294 , n296 , n297 , n301 , n305 , n310 , n311 , n312 , n313 , n314 , 
n316 , n318 , n321 , n323 , n325 , n331 , n334 , n336 , n337 , n338 , 
n340 , n341 , n343 , n344 , n345 , n348 , n349 , n352 , n353 , n354 , 
n357 , n358 , n365 , n366 , n368 , n369 , n370 , n371 , n375 , n377 , 
n378 , n380 , n382 , n385 , n386 , n388 , n390 , n392 , n393 , n395 , 
n397 , n400 , n403 , n404 , n408 , n410 , n424 , n426 , n428 , n433 , 
n435 , n438 , n440 , n441 , n442 , n443 , n451 , n452 , n454 , n456 , 
n457 , n458 , n460 , n462 , n463 , n466 , n472 , n474 , n475 , n478 , 
n479 , n481 , n483 , n484 , n485 , n486 , n487 , n491 , n492 , n494 , 
n495 , n500 , n511 , n513 , n519 , n521 , n524 , n526 , n527 , n529 , 
n534 , n535 , n540 , n541 , n542 , n544 , n545 , n546 , n547 , n549 , 
n551 , n552 , n553 , n556 , n557 , n558 , n562 , n564 , n571 , n572 , 
n575 , n579 , n587 , n591 , n592 , n596 , n597 , n598 , n609 , n610 , 
n611 , n615 , n618 , n620 , n622 , n623 , n624 , n628 , n629 , n633 , 
n636 , n640 , n641 , n643 , n645 , n647 , n654 , n665 , n667 , n669 , 
n673 , n677 , n680 , n681 , n690 , n693 , n695 , n696 , n698 , n700 , 
n704 , n705 , n706 , n707 , n709 , n712 , n715 , n716 , n718 , n719 , 
n724 , n725 , n727 , n728 , n730 , n731 , n732 , n736 , n740 , n741 , 
n743 , n747 , n748 , n753 , n756 , n759 , n760 , n762 , n763 , n765 , 
n769 , n770 , n772 , n773 , n775 , n777 , n781 , n783 , n786 , n789 , 
n790 , n791 , n792 , n795 , n796 , n798 , n801 , n804 , n808 , n809 , 
n810 , n813 , n814 , n815 , n819 , n822 , n828 , n836 , n838 , n839 , 
n841 , n846 , n848 , n855 , n856 , n862 , n865 , n867 , n869 , n870 , 
n871 , n874 , n876 , n877 , n880 , n889 , n892 , n893 , n894 , n901 , 
n902 , n904 , n905 , n907 , n908 , n910 , n915 , n920 , n921 , n922 , 
n924 , n925 , n926 , n931 , n937 , n940 , n941 , n942 , n943 , n944 , 
n945 , n946 , n949 , n950 );
    input n2 , n3 , n8 , n11 , n12 , n14 , n18 , n19 , n28 , 
n32 , n38 , n40 , n42 , n43 , n51 , n54 , n57 , n64 , n76 , 
n78 , n79 , n80 , n94 , n106 , n108 , n110 , n113 , n114 , n115 , 
n117 , n119 , n120 , n124 , n127 , n130 , n133 , n137 , n142 , n143 , 
n147 , n151 , n162 , n166 , n168 , n169 , n171 , n178 , n181 , n182 , 
n185 , n203 , n205 , n211 , n213 , n216 , n218 , n219 , n220 , n227 , 
n229 , n242 , n249 , n250 , n260 , n268 , n269 , n276 , n282 , n291 , 
n294 , n296 , n297 , n310 , n311 , n312 , n314 , n316 , n321 , n336 , 
n337 , n338 , n341 , n343 , n348 , n353 , n354 , n357 , n358 , n365 , 
n366 , n369 , n370 , n371 , n382 , n385 , n388 , n390 , n397 , n400 , 
n403 , n404 , n433 , n435 , n438 , n441 , n442 , n451 , n452 , n457 , 
n458 , n462 , n463 , n472 , n478 , n479 , n483 , n484 , n485 , n486 , 
n491 , n492 , n494 , n495 , n500 , n513 , n526 , n527 , n534 , n535 , 
n540 , n541 , n542 , n544 , n545 , n546 , n549 , n552 , n553 , n556 , 
n557 , n558 , n562 , n564 , n571 , n579 , n591 , n592 , n596 , n597 , 
n598 , n609 , n610 , n611 , n615 , n620 , n623 , n624 , n633 , n636 , 
n641 , n654 , n665 , n673 , n677 , n680 , n690 , n695 , n696 , n698 , 
n700 , n704 , n705 , n715 , n718 , n719 , n724 , n727 , n736 , n747 , 
n756 , n759 , n760 , n763 , n765 , n769 , n773 , n775 , n777 , n781 , 
n783 , n790 , n791 , n795 , n796 , n798 , n801 , n808 , n809 , n810 , 
n822 , n828 , n836 , n839 , n848 , n855 , n865 , n867 , n869 , n870 , 
n874 , n876 , n877 , n880 , n889 , n892 , n893 , n901 , n902 , n904 , 
n905 , n908 , n910 , n915 , n920 , n921 , n926 , n931 , n937 , n940 , 
n941 , n943 , n945 , n950 ;
    output n0 , n5 , n6 , n27 , n35 , n55 , n56 , n59 , n60 , 
n61 , n65 , n73 , n86 , n93 , n104 , n118 , n126 , n129 , n138 , 
n154 , n157 , n174 , n184 , n188 , n196 , n200 , n202 , n210 , n215 , 
n217 , n230 , n231 , n238 , n248 , n252 , n257 , n259 , n266 , n278 , 
n280 , n301 , n305 , n313 , n318 , n323 , n325 , n331 , n334 , n340 , 
n344 , n345 , n349 , n352 , n368 , n375 , n377 , n378 , n380 , n386 , 
n392 , n393 , n395 , n408 , n410 , n424 , n426 , n428 , n440 , n443 , 
n454 , n456 , n460 , n466 , n474 , n475 , n481 , n487 , n511 , n519 , 
n521 , n524 , n529 , n547 , n551 , n572 , n575 , n587 , n618 , n622 , 
n628 , n629 , n640 , n643 , n645 , n647 , n667 , n669 , n681 , n693 , 
n706 , n707 , n709 , n712 , n716 , n725 , n728 , n730 , n731 , n732 , 
n740 , n741 , n743 , n748 , n753 , n762 , n770 , n772 , n786 , n789 , 
n792 , n804 , n813 , n814 , n815 , n819 , n838 , n841 , n846 , n856 , 
n862 , n871 , n894 , n907 , n922 , n924 , n925 , n942 , n944 , n946 , 
n949 ;
    wire n1 , n4 , n7 , n9 , n10 , n13 , n15 , n16 , n17 , 
n20 , n21 , n22 , n23 , n24 , n25 , n26 , n29 , n30 , n31 , 
n33 , n34 , n36 , n37 , n39 , n41 , n44 , n45 , n46 , n47 , 
n48 , n49 , n50 , n52 , n53 , n58 , n62 , n63 , n66 , n67 , 
n68 , n69 , n70 , n71 , n72 , n74 , n75 , n77 , n81 , n82 , 
n83 , n84 , n85 , n87 , n88 , n89 , n90 , n91 , n92 , n95 , 
n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n105 , n107 , 
n109 , n111 , n112 , n116 , n121 , n122 , n123 , n125 , n128 , n131 , 
n132 , n134 , n135 , n136 , n139 , n140 , n141 , n144 , n145 , n146 , 
n148 , n149 , n150 , n152 , n153 , n155 , n156 , n158 , n159 , n160 , 
n161 , n163 , n164 , n165 , n167 , n170 , n172 , n173 , n175 , n176 , 
n177 , n179 , n180 , n183 , n186 , n187 , n189 , n190 , n191 , n192 , 
n193 , n194 , n195 , n197 , n198 , n199 , n201 , n204 , n206 , n207 , 
n208 , n209 , n212 , n214 , n221 , n222 , n223 , n224 , n225 , n226 , 
n228 , n232 , n233 , n234 , n235 , n236 , n237 , n239 , n240 , n241 , 
n243 , n244 , n245 , n246 , n247 , n251 , n253 , n254 , n255 , n256 , 
n258 , n261 , n262 , n263 , n264 , n265 , n267 , n270 , n271 , n272 , 
n273 , n274 , n275 , n277 , n279 , n281 , n283 , n284 , n285 , n286 , 
n287 , n288 , n289 , n290 , n292 , n293 , n295 , n298 , n299 , n300 , 
n302 , n303 , n304 , n306 , n307 , n308 , n309 , n315 , n317 , n319 , 
n320 , n322 , n324 , n326 , n327 , n328 , n329 , n330 , n332 , n333 , 
n335 , n339 , n342 , n346 , n347 , n350 , n351 , n355 , n356 , n359 , 
n360 , n361 , n362 , n363 , n364 , n367 , n372 , n373 , n374 , n376 , 
n379 , n381 , n383 , n384 , n387 , n389 , n391 , n394 , n396 , n398 , 
n399 , n401 , n402 , n405 , n406 , n407 , n409 , n411 , n412 , n413 , 
n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , 
n425 , n427 , n429 , n430 , n431 , n432 , n434 , n436 , n437 , n439 , 
n444 , n445 , n446 , n447 , n448 , n449 , n450 , n453 , n455 , n459 , 
n461 , n464 , n465 , n467 , n468 , n469 , n470 , n471 , n473 , n476 , 
n477 , n480 , n482 , n488 , n489 , n490 , n493 , n496 , n497 , n498 , 
n499 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
n510 , n512 , n514 , n515 , n516 , n517 , n518 , n520 , n522 , n523 , 
n525 , n528 , n530 , n531 , n532 , n533 , n536 , n537 , n538 , n539 , 
n543 , n548 , n550 , n554 , n555 , n559 , n560 , n561 , n563 , n565 , 
n566 , n567 , n568 , n569 , n570 , n573 , n574 , n576 , n577 , n578 , 
n580 , n581 , n582 , n583 , n584 , n585 , n586 , n588 , n589 , n590 , 
n593 , n594 , n595 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , 
n606 , n607 , n608 , n612 , n613 , n614 , n616 , n617 , n619 , n621 , 
n625 , n626 , n627 , n630 , n631 , n632 , n634 , n635 , n637 , n638 , 
n639 , n642 , n644 , n646 , n648 , n649 , n650 , n651 , n652 , n653 , 
n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , 
n666 , n668 , n670 , n671 , n672 , n674 , n675 , n676 , n678 , n679 , 
n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n691 , n692 , 
n694 , n697 , n699 , n701 , n702 , n703 , n708 , n710 , n711 , n713 , 
n714 , n717 , n720 , n721 , n722 , n723 , n726 , n729 , n733 , n734 , 
n735 , n737 , n738 , n739 , n742 , n744 , n745 , n746 , n749 , n750 , 
n751 , n752 , n754 , n755 , n757 , n758 , n761 , n764 , n766 , n767 , 
n768 , n771 , n774 , n776 , n778 , n779 , n780 , n782 , n784 , n785 , 
n787 , n788 , n793 , n794 , n797 , n799 , n800 , n802 , n803 , n805 , 
n806 , n807 , n811 , n812 , n816 , n817 , n818 , n820 , n821 , n823 , 
n824 , n825 , n826 , n827 , n829 , n830 , n831 , n832 , n833 , n834 , 
n835 , n837 , n840 , n842 , n843 , n844 , n845 , n847 , n849 , n850 , 
n851 , n852 , n853 , n854 , n857 , n858 , n859 , n860 , n861 , n863 , 
n864 , n866 , n868 , n872 , n873 , n875 , n878 , n879 , n881 , n882 , 
n883 , n884 , n885 , n886 , n887 , n888 , n890 , n891 , n895 , n896 , 
n897 , n898 , n899 , n900 , n903 , n906 , n909 , n911 , n912 , n913 , 
n914 , n916 , n917 , n918 , n919 , n923 , n927 , n928 , n929 , n930 , 
n932 , n933 , n934 , n935 , n936 , n938 , n939 , n947 , n948 ;
    and g0 ( n356 , n755 , n156 );
    not g1 ( n152 , n397 );
    buf g2 ( n946 , n673 );
    xor g3 ( n195 , n475 , n629 );
    and g4 ( n538 , n2 , n928 );
    or g5 ( n62 , n849 , n360 );
    or g6 ( n764 , n726 , n360 );
    buf g7 ( n712 , n11 );
    not g8 ( n722 , n905 );
    nor g9 ( n15 , n268 , n803 );
    and g10 ( n543 , n798 , n834 );
    or g11 ( n132 , n509 , n63 );
    nor g12 ( n226 , n362 , n684 );
    and g13 ( n204 , n21 , n277 );
    nor g14 ( n482 , n585 , n69 );
    and g15 ( n4 , n845 , n800 );
    not g16 ( n272 , n260 );
    nor g17 ( n122 , n635 , n608 );
    not g18 ( n632 , n388 );
    and g19 ( n101 , n579 , n272 );
    xnor g20 ( n807 , n407 , n459 );
    buf g21 ( n257 , n795 );
    or g22 ( n295 , n244 , n476 );
    or g23 ( n179 , n649 , n204 );
    xnor g24 ( n146 , n264 , n704 );
    not g25 ( n362 , n620 );
    buf g26 ( n753 , n366 );
    buf g27 ( n647 , n321 );
    buf g28 ( n188 , n677 );
    or g29 ( n475 , n829 , n9 );
    nor g30 ( n734 , n692 , n523 );
    nor g31 ( n372 , n63 , n395 );
    xnor g32 ( n531 , n460 , n711 );
    buf g33 ( n730 , n454 );
    nor g34 ( n574 , n620 , n140 );
    or g35 ( n618 , n105 , n569 );
    xnor g36 ( n851 , n178 , n353 );
    or g37 ( n919 , n613 , n131 );
    or g38 ( n288 , n642 , n365 );
    not g39 ( n84 , n941 );
    or g40 ( n924 , n649 , n26 );
    buf g41 ( n352 , n371 );
    or g42 ( n91 , n75 , n694 );
    or g43 ( n89 , n771 , n878 );
    not g44 ( n163 , n801 );
    and g45 ( n489 , n945 , n610 );
    or g46 ( n299 , n927 , n427 );
    buf g47 ( n725 , n366 );
    not g48 ( n254 , n229 );
    or g49 ( n422 , n292 , n365 );
    and g50 ( n672 , n798 , n98 );
    buf g51 ( n154 , n218 );
    or g52 ( n454 , n328 , n903 );
    not g53 ( n439 , n40 );
    xnor g54 ( n668 , n791 , n541 );
    not g55 ( n187 , n806 );
    and g56 ( n261 , n203 , n270 );
    not g57 ( n301 , n867 );
    and g58 ( n176 , n460 , n156 );
    or g59 ( n820 , n911 , n369 );
    and g60 ( n398 , n343 , n256 );
    nor g61 ( n490 , n272 , n288 );
    not g62 ( n831 , n276 );
    or g63 ( n875 , n675 , n103 );
    buf g64 ( n375 , n915 );
    buf g65 ( n547 , n556 );
    or g66 ( n102 , n528 , n365 );
    and g67 ( n449 , n282 , n236 );
    buf g68 ( n5 , n54 );
    or g69 ( n894 , n758 , n85 );
    or g70 ( n499 , n612 , n369 );
    buf g71 ( n61 , n106 );
    or g72 ( n53 , n251 , n245 );
    not g73 ( n563 , n791 );
    buf g74 ( n862 , n760 );
    xnor g75 ( n243 , n891 , n598 );
    not g76 ( n394 , n57 );
    nor g77 ( n825 , n517 , n373 );
    or g78 ( n389 , n776 , n36 );
    not g79 ( n802 , n117 );
    buf g80 ( n118 , n119 );
    or g81 ( n933 , n929 , n369 );
    and g82 ( n584 , n372 , n465 );
    or g83 ( n277 , n705 , n928 );
    not g84 ( n528 , n546 );
    buf g85 ( n575 , n540 );
    and g86 ( n794 , n847 , n934 );
    and g87 ( n190 , n268 , n803 );
    not g88 ( n284 , n680 );
    or g89 ( n361 , n538 , n510 );
    not g90 ( n329 , n542 );
    nor g91 ( n34 , n272 , n469 );
    not g92 ( n674 , n491 );
    nor g93 ( n244 , n68 , n322 );
    nor g94 ( n568 , n362 , n607 );
    not g95 ( n686 , n18 );
    or g96 ( n646 , n152 , n365 );
    and g97 ( n69 , n98 , n156 );
    buf g98 ( n622 , n168 );
    xnor g99 ( n583 , n240 , n367 );
    not g100 ( n16 , n76 );
    nor g101 ( n746 , n362 , n499 );
    or g102 ( n566 , n906 , n744 );
    or g103 ( n731 , n284 , n392 );
    and g104 ( n447 , n545 , n588 );
    and g105 ( n833 , n649 , n204 );
    and g106 ( n315 , n763 , n256 );
    not g107 ( n550 , n432 );
    or g108 ( n628 , n766 , n721 );
    nor g109 ( n95 , n378 , n4 );
    nor g110 ( n302 , n272 , n374 );
    not g111 ( n145 , n848 );
    nor g112 ( n41 , n600 , n599 );
    or g113 ( n891 , n109 , n45 );
    or g114 ( n196 , n745 , n506 );
    not g115 ( n285 , n711 );
    or g116 ( n771 , n554 , n228 );
    buf g117 ( n313 , n877 );
    nor g118 ( n692 , n362 , n233 );
    not g119 ( n309 , n341 );
    nor g120 ( n401 , n815 , n772 );
    or g121 ( n158 , n411 , n365 );
    xnor g122 ( n701 , n173 , n682 );
    and g123 ( n666 , n452 , n365 );
    nor g124 ( n71 , n1 , n364 );
    buf g125 ( n907 , n143 );
    nor g126 ( n793 , n25 , n701 );
    not g127 ( n512 , n615 );
    or g128 ( n200 , n576 , n319 );
    and g129 ( n134 , n494 , n708 );
    nor g130 ( n532 , n620 , n23 );
    buf g131 ( n428 , n403 );
    xnor g132 ( n930 , n206 , n668 );
    and g133 ( n737 , n438 , n708 );
    not g134 ( n464 , n296 );
    nor g135 ( n275 , n272 , n646 );
    xnor g136 ( n240 , n910 , n124 );
    or g137 ( n631 , n840 , n437 );
    xnor g138 ( n473 , n467 , n216 );
    or g139 ( n207 , n275 , n797 );
    or g140 ( n85 , n477 , n750 );
    or g141 ( n23 , n376 , n360 );
    or g142 ( n283 , n588 , n833 );
    or g143 ( n177 , n702 , n369 );
    nor g144 ( n947 , n272 , n923 );
    not g145 ( n612 , n242 );
    or g146 ( n852 , n570 , n360 );
    nor g147 ( n530 , n362 , n606 );
    xnor g148 ( n206 , n297 , n8 );
    not g149 ( n419 , n920 );
    and g150 ( n648 , n507 , n525 );
    or g151 ( n279 , n512 , n290 );
    or g152 ( n585 , n705 , n471 );
    xnor g153 ( n936 , n866 , n791 );
    not g154 ( n678 , n790 );
    buf g155 ( n944 , n880 );
    or g156 ( n561 , n689 , n135 );
    or g157 ( n835 , n7 , n948 );
    xnor g158 ( n164 , n884 , n656 );
    or g159 ( n520 , n49 , n122 );
    buf g160 ( n706 , n527 );
    nor g161 ( n627 , n115 , n52 );
    and g162 ( n886 , n171 , n708 );
    or g163 ( n664 , n625 , n580 );
    not g164 ( n150 , n651 );
    or g165 ( n629 , n271 , n566 );
    nor g166 ( n67 , n601 , n263 );
    not g167 ( n170 , n549 );
    or g168 ( n460 , n844 , n881 );
    or g169 ( n46 , n663 , n536 );
    not g170 ( n408 , n834 );
    and g171 ( n537 , n777 , n708 );
    nor g172 ( n903 , n464 , n909 );
    and g173 ( n476 , n618 , n559 );
    buf g174 ( n386 , n775 );
    xnor g175 ( n367 , n769 , n908 );
    or g176 ( n914 , n153 , n713 );
    not g177 ( n693 , n521 );
    xnor g178 ( n821 , n900 , n769 );
    or g179 ( n617 , n739 , n263 );
    not g180 ( n498 , n220 );
    not g181 ( n651 , n603 );
    buf g182 ( n73 , n931 );
    or g183 ( n105 , n214 , n589 );
    or g184 ( n602 , n683 , n561 );
    nor g185 ( n412 , n864 , n31 );
    or g186 ( n48 , n947 , n888 );
    not g187 ( n210 , n552 );
    nor g188 ( n554 , n507 , n525 );
    buf g189 ( n325 , n485 );
    nor g190 ( n832 , n296 , n285 );
    buf g191 ( n0 , n166 );
    or g192 ( n761 , n757 , n365 );
    or g193 ( n853 , n144 , n360 );
    nor g194 ( n697 , n464 , n572 );
    buf g195 ( n157 , n700 );
    not g196 ( n757 , n357 );
    or g197 ( n350 , n448 , n365 );
    buf g198 ( n511 , n93 );
    or g199 ( n471 , n175 , n501 );
    and g200 ( n395 , n136 , n449 );
    nor g201 ( n663 , n272 , n717 );
    and g202 ( n818 , n337 , n256 );
    and g203 ( n548 , n798 , n289 );
    not g204 ( n378 , n305 );
    not g205 ( n770 , n492 );
    or g206 ( n899 , n739 , n263 );
    and g207 ( n97 , n798 , n785 );
    or g208 ( n720 , n826 , n735 );
    or g209 ( n838 , n751 , n835 );
    or g210 ( n324 , n112 , n365 );
    and g211 ( n247 , n110 , n256 );
    not g212 ( n308 , n719 );
    xnor g213 ( n99 , n201 , n910 );
    not g214 ( n928 , n651 );
    or g215 ( n172 , n239 , n187 );
    nor g216 ( n66 , n620 , n62 );
    buf g217 ( n871 , n458 );
    and g218 ( n461 , n545 , n649 );
    not g219 ( n175 , n354 );
    not g220 ( n274 , n32 );
    or g221 ( n149 , n720 , n898 );
    or g222 ( n829 , n101 , n708 );
    buf g223 ( n334 , n633 );
    buf g224 ( n217 , n696 );
    and g225 ( n47 , n680 , n85 );
    and g226 ( n82 , n3 , n270 );
    nor g227 ( n186 , n362 , n413 );
    or g228 ( n24 , n82 , n644 );
    or g229 ( n201 , n315 , n896 );
    or g230 ( n413 , n16 , n369 );
    and g231 ( n425 , n779 , n825 );
    or g232 ( n107 , n398 , n671 );
    or g233 ( n399 , n256 , n265 );
    or g234 ( n236 , n788 , n189 );
    or g235 ( n789 , n509 , n221 );
    not g236 ( n96 , n823 );
    or g237 ( n799 , n752 , n859 );
    or g238 ( n307 , n498 , n369 );
    not g239 ( n39 , n592 );
    not g240 ( n155 , n553 );
    or g241 ( n507 , n752 , n567 );
    buf g242 ( n741 , n623 );
    and g243 ( n328 , n464 , n588 );
    nor g244 ( n895 , n383 , n914 );
    nor g245 ( n22 , n362 , n784 );
    or g246 ( n469 , n234 , n365 );
    nor g247 ( n768 , n272 , n468 );
    not g248 ( n752 , n249 );
    xnor g249 ( n823 , n195 , n531 );
    nor g250 ( n676 , n710 , n141 );
    or g251 ( n323 , n860 , n132 );
    or g252 ( n782 , n330 , n604 );
    and g253 ( n688 , n219 , n708 );
    buf g254 ( n814 , n400 );
    not g255 ( n199 , n783 );
    buf g256 ( n349 , n182 );
    or g257 ( n271 , n581 , n537 );
    and g258 ( n153 , n378 , n4 );
    nor g259 ( n26 , n950 , n909 );
    or g260 ( n751 , n863 , n563 );
    and g261 ( n320 , n249 , n629 );
    xnor g262 ( n116 , n534 , n314 );
    buf g263 ( n60 , n169 );
    and g264 ( n303 , n937 , n270 );
    not g265 ( n138 , n698 );
    buf g266 ( n56 , n557 );
    xnor g267 ( n396 , n173 , n504 );
    or g268 ( n384 , n274 , n290 );
    xnor g269 ( n594 , n807 , n811 );
    not g270 ( n430 , n889 );
    not g271 ( n480 , n718 );
    and g272 ( n605 , n464 , n649 );
    buf g273 ( n709 , n486 );
    nor g274 ( n604 , n620 , n355 );
    buf g275 ( n443 , n558 );
    and g276 ( n896 , n798 , n91 );
    buf g277 ( n732 , n839 );
    or g278 ( n860 , n439 , n632 );
    or g279 ( n487 , n505 , n588 );
    xnor g280 ( n191 , n107 , n297 );
    nor g281 ( n934 , n950 , n148 );
    not g282 ( n812 , n133 );
    and g283 ( n859 , n791 , n938 );
    or g284 ( n180 , n416 , n365 );
    and g285 ( n729 , n545 , n618 );
    nor g286 ( n518 , n362 , n198 );
    not g287 ( n816 , n356 );
    and g288 ( n326 , n636 , n270 );
    and g289 ( n644 , n545 , n460 );
    not g290 ( n942 , n724 );
    and g291 ( n212 , n950 , n711 );
    nor g292 ( n858 , n272 , n347 );
    or g293 ( n289 , n861 , n299 );
    xnor g294 ( n658 , n695 , n855 );
    or g295 ( n576 , n121 , n919 );
    not g296 ( n339 , n641 );
    or g297 ( n515 , n450 , n461 );
    or g298 ( n824 , n27 , n210 );
    not g299 ( n573 , n42 );
    nor g300 ( n49 , n53 , n617 );
    or g301 ( n141 , n383 , n713 );
    or g302 ( n754 , n593 , n81 );
    or g303 ( n506 , n509 , n63 );
    not g304 ( n551 , n466 );
    or g305 ( n319 , n653 , n300 );
    not g306 ( n112 , n564 );
    or g307 ( n131 , n99 , n555 );
    nor g308 ( n906 , n272 , n346 );
    not g309 ( n938 , n603 );
    or g310 ( n850 , n639 , n100 );
    nor g311 ( n779 , n490 , n737 );
    xnor g312 ( n407 , n278 , n408 );
    buf g313 ( n529 , n14 );
    nor g314 ( n703 , n620 , n820 );
    or g315 ( n510 , n752 , n208 );
    not g316 ( n488 , n478 );
    buf g317 ( n440 , n269 );
    buf g318 ( n259 , n435 );
    and g319 ( n601 , n91 , n156 );
    and g320 ( n263 , n585 , n69 );
    and g321 ( n935 , n249 , n184 );
    or g322 ( n209 , n304 , n548 );
    or g323 ( n539 , n361 , n648 );
    or g324 ( n613 , n387 , n821 );
    or g325 ( n477 , n138 , n301 );
    not g326 ( n755 , n910 );
    not g327 ( n270 , n545 );
    and g328 ( n559 , n502 , n714 );
    or g329 ( n749 , n420 , n799 );
    buf g330 ( n104 , n38 );
    or g331 ( n493 , n224 , n543 );
    buf g332 ( n643 , 1'b0 );
    xnor g333 ( n432 , n909 , n173 );
    buf g334 ( n266 , n294 );
    or g335 ( n347 , n885 , n290 );
    or g336 ( n882 , n879 , n577 );
    and g337 ( n359 , n79 , n270 );
    or g338 ( n606 , n470 , n360 );
    nor g339 ( n522 , n260 , n429 );
    buf g340 ( n174 , n759 );
    buf g341 ( n846 , n370 );
    and g342 ( n735 , n317 , n434 );
    and g343 ( n420 , n211 , n928 );
    xor g344 ( n887 , n52 , n280 );
    or g345 ( n355 , n170 , n360 );
    not g346 ( n863 , n297 );
    xnor g347 ( n197 , n358 , n705 );
    and g348 ( n614 , n545 , n475 );
    nor g349 ( n864 , n58 , n830 );
    not g350 ( n778 , n535 );
    nor g351 ( n776 , n272 , n422 );
    nor g352 ( n523 , n620 , n939 );
    not g353 ( n516 , n151 );
    not g354 ( n234 , n926 );
    buf g355 ( n231 , n673 );
    or g356 ( n414 , n634 , n83 );
    not g357 ( n837 , n940 );
    and g358 ( n661 , n890 , n176 );
    and g359 ( n913 , n533 , n150 );
    or g360 ( n890 , n908 , n471 );
    or g361 ( n569 , n34 , n409 );
    or g362 ( n684 , n691 , n360 );
    nor g363 ( n655 , n620 , n391 );
    or g364 ( n603 , n175 , n172 );
    or g365 ( n567 , n704 , n938 );
    not g366 ( n448 , n227 );
    buf g367 ( n248 , n181 );
    or g368 ( n77 , n186 , n273 );
    or g369 ( n710 , n100 , n648 );
    nor g370 ( n455 , n96 , n223 );
    nor g371 ( n595 , n464 , n305 );
    not g372 ( n30 , n495 );
    or g373 ( n445 , n241 , n672 );
    not g374 ( n649 , n425 );
    xnor g375 ( n682 , n333 , n195 );
    xnor g376 ( n87 , n493 , n541 );
    or g377 ( n415 , n883 , n50 );
    buf g378 ( n716 , n336 );
    or g379 ( n653 , n159 , n37 );
    xnor g380 ( n496 , n515 , n534 );
    nor g381 ( n634 , n362 , n853 );
    or g382 ( n638 , n303 , n111 );
    and g383 ( n305 , n733 , n298 );
    or g384 ( n167 , n39 , n360 );
    or g385 ( n128 , n621 , n436 );
    or g386 ( n192 , n423 , n916 );
    or g387 ( n497 , n329 , n369 );
    or g388 ( n13 , n626 , n290 );
    and g389 ( n912 , n545 , n521 );
    or g390 ( n21 , n534 , n938 );
    xnor g391 ( n173 , n649 , n588 );
    or g392 ( n939 , n308 , n360 );
    and g393 ( n342 , n736 , n708 );
    or g394 ( n165 , n879 , n263 );
    nor g395 ( n262 , n235 , n655 );
    nor g396 ( n797 , n260 , n158 );
    xnor g397 ( n555 , n445 , n705 );
    or g398 ( n121 , n917 , n560 );
    or g399 ( n565 , n767 , n365 );
    and g400 ( n593 , n356 , n67 );
    and g401 ( n739 , n816 , n601 );
    nor g402 ( n273 , n620 , n652 );
    nor g403 ( n431 , n260 , n102 );
    and g404 ( n100 , n335 , n913 );
    or g405 ( n52 , n414 , n868 );
    not g406 ( n377 , n894 );
    or g407 ( n900 , n247 , n97 );
    buf g408 ( n238 , n596 );
    or g409 ( n306 , n823 , n396 );
    not g410 ( n292 , n796 );
    buf g411 ( n202 , n126 );
    buf g412 ( n331 , n472 );
    or g413 ( n923 , n258 , n290 );
    or g414 ( n805 , n139 , n360 );
    or g415 ( n873 , n20 , n134 );
    nor g416 ( n927 , n362 , n293 );
    nor g417 ( n322 , n910 , n928 );
    or g418 ( n861 , n226 , n444 );
    and g419 ( n109 , n213 , n270 );
    or g420 ( n327 , n573 , n360 );
    or g421 ( n619 , n199 , n290 );
    and g422 ( n766 , n115 , n52 );
    or g423 ( n136 , n738 , n780 );
    and g424 ( n466 , n584 , n401 );
    nor g425 ( n135 , n620 , n586 );
    buf g426 ( n743 , n513 );
    xnor g427 ( n387 , n24 , n908 );
    not g428 ( n509 , n19 );
    not g429 ( n290 , n365 );
    or g430 ( n742 , n488 , n369 );
    not g431 ( n255 , n348 );
    buf g432 ( n587 , n463 );
    nor g433 ( n508 , n362 , n842 );
    not g434 ( n830 , n701 );
    nor g435 ( n36 , n260 , n160 );
    or g436 ( n74 , n482 , n754 );
    or g437 ( n251 , n769 , n471 );
    or g438 ( n872 , n100 , n648 );
    and g439 ( n525 , n320 , n150 );
    or g440 ( n588 , n415 , n389 );
    nor g441 ( n364 , n283 , n295 );
    nor g442 ( n434 , n648 , n383 );
    and g443 ( n878 , n95 , n676 );
    nor g444 ( n409 , n260 , n180 );
    buf g445 ( n669 , n673 );
    or g446 ( n784 , n30 , n360 );
    and g447 ( n806 , n480 , n834 );
    or g448 ( n160 , n831 , n365 );
    or g449 ( n363 , n15 , n243 );
    or g450 ( n429 , n394 , n365 );
    xnor g451 ( n788 , n286 , n446 );
    and g452 ( n660 , n545 , n629 );
    or g453 ( n868 , n508 , n703 );
    nor g454 ( n675 , n362 , n650 );
    xnor g455 ( n17 , n2 , n211 );
    or g456 ( n714 , n358 , n150 );
    and g457 ( n713 , n935 , n749 );
    or g458 ( n586 , n232 , n369 );
    buf g459 ( n368 , n338 );
    nor g460 ( n840 , n620 , n167 );
    or g461 ( n842 , n255 , n369 );
    or g462 ( n582 , n84 , n369 );
    or g463 ( n300 , n192 , n128 );
    nor g464 ( n68 , n314 , n938 );
    or g465 ( n405 , n222 , n518 );
    not g466 ( n767 , n597 );
    nor g467 ( n657 , n260 , n565 );
    buf g468 ( n345 , n892 );
    nor g469 ( n616 , n872 , n421 );
    nand g470 ( n221 , n943 , n162 );
    not g471 ( n626 , n500 );
    or g472 ( n707 , n161 , n392 );
    nor g473 ( n418 , n272 , n685 );
    or g474 ( n918 , n568 , n574 );
    and g475 ( n304 , n94 , n256 );
    nor g476 ( n625 , n362 , n774 );
    xnor g477 ( n246 , n851 , n658 );
    or g478 ( n854 , n770 , n55 );
    nor g479 ( n20 , n272 , n13 );
    or g480 ( n721 , n836 , n627 );
    buf g481 ( n86 , n747 );
    not g482 ( n849 , n611 );
    and g483 ( n383 , n639 , n361 );
    and g484 ( n772 , n306 , n630 );
    or g485 ( n881 , n768 , n431 );
    not g486 ( n911 , n665 );
    and g487 ( n879 , n251 , n245 );
    buf g488 ( n252 , n902 );
    not g489 ( n885 , n51 );
    or g490 ( n467 , n72 , n614 );
    and g491 ( n92 , n316 , n270 );
    or g492 ( n774 , n722 , n369 );
    and g493 ( n843 , n464 , n618 );
    not g494 ( n90 , n526 );
    buf g495 ( n380 , n865 );
    or g496 ( n844 , n351 , n342 );
    not g497 ( n929 , n142 );
    nor g498 ( n517 , n272 , n619 );
    or g499 ( n685 , n837 , n365 );
    or g500 ( n578 , n858 , n886 );
    and g501 ( n421 , n514 , n71 );
    xnor g502 ( n656 , n598 , n268 );
    or g503 ( n198 , n812 , n369 );
    not g504 ( n702 , n562 );
    and g505 ( n916 , n637 , n399 );
    or g506 ( n184 , n873 , n46 );
    and g507 ( n708 , n365 , n272 );
    or g508 ( n683 , n22 , n66 );
    not g509 ( n505 , n950 );
    nor g510 ( n103 , n620 , n852 );
    or g511 ( n758 , n824 , n854 );
    nor g512 ( n536 , n260 , n350 );
    or g513 ( n267 , n661 , n882 );
    nor g514 ( n659 , n620 , n933 );
    not g515 ( n411 , n442 );
    and g516 ( n280 , n734 , n262 );
    or g517 ( n503 , n817 , n699 );
    and g518 ( n208 , n297 , n938 );
    and g519 ( n111 , n545 , n184 );
    xnor g520 ( n600 , n887 , n602 );
    buf g521 ( n925 , n715 );
    not g522 ( n281 , n108 );
    buf g523 ( n645 , n571 );
    buf g524 ( n841 , n756 );
    buf g525 ( n424 , n400 );
    buf g526 ( n922 , n822 );
    nor g527 ( n883 , n272 , n379 );
    xnor g528 ( n402 , n590 , n314 );
    xnor g529 ( n811 , n785 , n91 );
    and g530 ( n70 , n870 , n758 );
    or g531 ( n519 , n212 , n794 );
    or g532 ( n392 , n155 , n509 );
    not g533 ( n223 , n396 );
    not g534 ( n278 , n239 );
    buf g535 ( n129 , n609 );
    or g536 ( n917 , n473 , n146 );
    buf g537 ( n318 , n137 );
    or g538 ( n140 , n145 , n360 );
    nor g539 ( n630 , n43 , n455 );
    and g540 ( n450 , n147 , n270 );
    buf g541 ( n6 , n828 );
    or g542 ( n834 , n918 , n77 );
    not g543 ( n144 , n312 );
    or g544 ( n225 , n430 , n369 );
    buf g545 ( n856 , n120 );
    or g546 ( n866 , n818 , n679 );
    not g547 ( n423 , n893 );
    nor g548 ( n826 , n850 , n539 );
    not g549 ( n360 , n369 );
    xnor g550 ( n662 , n930 , n197 );
    or g551 ( n786 , n832 , n412 );
    or g552 ( n417 , n287 , n290 );
    or g553 ( n159 , n88 , n87 );
    or g554 ( n37 , n936 , n191 );
    nor g555 ( n817 , n362 , n742 );
    not g556 ( n25 , n58 );
    and g557 ( n241 , n591 , n256 );
    not g558 ( n827 , n28 );
    or g559 ( n379 , n163 , n290 );
    or g560 ( n800 , n541 , n150 );
    or g561 ( n123 , n261 , n912 );
    nor g562 ( n444 , n620 , n10 );
    or g563 ( n650 , n419 , n360 );
    or g564 ( n694 , n532 , n659 );
    buf g565 ( n410 , n400 );
    or g566 ( n514 , n476 , n179 );
    or g567 ( n785 , n782 , n664 );
    nor g568 ( n148 , n711 , n432 );
    nor g569 ( n689 , n362 , n307 );
    or g570 ( n468 , n516 , n365 );
    not g571 ( n570 , n385 );
    not g572 ( n189 , n780 );
    xnor g573 ( n237 , n115 , n836 );
    xnor g574 ( n884 , n857 , n17 );
    xnor g575 ( n446 , n78 , n80 );
    or g576 ( n521 , n578 , n453 );
    or g577 ( n264 , n92 , n660 );
    buf g578 ( n804 , n441 );
    not g579 ( n642 , n727 );
    xnor g580 ( n787 , n638 , n211 );
    not g581 ( n33 , n451 );
    and g582 ( n224 , n457 , n256 );
    nor g583 ( n723 , n272 , n332 );
    nor g584 ( n298 , n688 , n657 );
    xnor g585 ( n35 , n662 , n237 );
    buf g586 ( n681 , n544 );
    or g587 ( n803 , n359 , n729 );
    or g588 ( n711 , n48 , n207 );
    buf g589 ( n456 , n130 );
    or g590 ( n501 , n239 , n806 );
    buf g591 ( n59 , n311 );
    buf g592 ( n524 , n483 );
    nor g593 ( n744 , n260 , n324 );
    and g594 ( n50 , n390 , n708 );
    not g595 ( n232 , n64 );
    nor g596 ( n330 , n362 , n764 );
    buf g597 ( n762 , n690 );
    not g598 ( n416 , n781 );
    not g599 ( n948 , n358 );
    nor g600 ( n427 , n620 , n177 );
    not g601 ( n183 , n600 );
    or g602 ( n637 , n281 , n798 );
    not g603 ( n726 , n773 );
    not g604 ( n139 , n127 );
    or g605 ( n436 , n496 , n402 );
    not g606 ( n381 , n624 );
    buf g607 ( n640 , n291 );
    not g608 ( n265 , n52 );
    nor g609 ( n29 , n43 , n41 );
    or g610 ( n453 , n418 , n522 );
    or g611 ( n10 , n33 , n360 );
    not g612 ( n256 , n798 );
    not g613 ( n691 , n12 );
    nor g614 ( n437 , n620 , n582 );
    or g615 ( n847 , n285 , n550 );
    or g616 ( n239 , n405 , n631 );
    or g617 ( n560 , n787 , n687 );
    xnor g618 ( n857 , n704 , n216 );
    xnor g619 ( n333 , n618 , n521 );
    or g620 ( n9 , n666 , n44 );
    or g621 ( n621 , n190 , n363 );
    and g622 ( n45 , n545 , n378 );
    or g623 ( n845 , n598 , n938 );
    nor g624 ( n83 , n620 , n805 );
    nor g625 ( n671 , n256 , n280 );
    nor g626 ( n214 , n272 , n384 );
    not g627 ( n728 , n63 );
    or g628 ( n717 , n778 , n365 );
    buf g629 ( n393 , n479 );
    and g630 ( n792 , n673 , n404 );
    nor g631 ( n699 , n620 , n406 );
    nor g632 ( n580 , n620 , n225 );
    or g633 ( n98 , n875 , n503 );
    not g634 ( n738 , n788 );
    not g635 ( n470 , n874 );
    xnor g636 ( n58 , n909 , n531 );
    and g637 ( n909 , n674 , n425 );
    buf g638 ( n426 , n921 );
    or g639 ( n608 , n176 , n165 );
    not g640 ( n258 , n808 );
    or g641 ( n93 , n595 , n605 );
    xnor g642 ( n780 , n116 , n246 );
    or g643 ( n335 , n752 , n194 );
    or g644 ( n31 , n464 , n793 );
    nor g645 ( n581 , n272 , n279 );
    and g646 ( n888 , n654 , n708 );
    not g647 ( n670 , n809 );
    xnor g648 ( n504 , n184 , n193 );
    buf g649 ( n474 , n382 );
    or g650 ( n607 , n827 , n360 );
    or g651 ( n253 , n254 , n365 );
    nor g652 ( n81 , n899 , n267 );
    buf g653 ( n344 , n810 );
    or g654 ( n126 , n697 , n843 );
    not g655 ( n376 , n114 );
    or g656 ( n340 , n520 , n74 );
    and g657 ( n898 , n895 , n616 );
    and g658 ( n72 , n310 , n270 );
    nor g659 ( n228 , n125 , n648 );
    nor g660 ( n351 , n272 , n417 );
    nor g661 ( n733 , n302 , n723 );
    or g662 ( n75 , n530 , n746 );
    nor g663 ( n577 , n89 , n149 );
    or g664 ( n374 , n381 , n290 );
    buf g665 ( n667 , n869 );
    buf g666 ( n819 , n484 );
    or g667 ( n897 , n935 , n100 );
    or g668 ( n652 , n670 , n369 );
    and g669 ( n679 , n798 , n239 );
    nor g670 ( n222 , n362 , n327 );
    xnor g671 ( n230 , n164 , n583 );
    not g672 ( n161 , n870 );
    buf g673 ( n813 , n673 );
    or g674 ( n332 , n90 , n365 );
    xnor g675 ( n88 , n209 , n358 );
    or g676 ( n750 , n942 , n65 );
    nor g677 ( n1 , n618 , n559 );
    not g678 ( n55 , n250 );
    or g679 ( n406 , n802 , n369 );
    buf g680 ( n740 , n786 );
    not g681 ( n65 , n765 );
    and g682 ( n589 , n462 , n708 );
    buf g683 ( n949 , n904 );
    xnor g684 ( n286 , n205 , n185 );
    buf g685 ( n481 , n113 );
    not g686 ( n156 , n471 );
    nor g687 ( n44 , n272 , n253 );
    xnor g688 ( n193 , n378 , n333 );
    or g689 ( n233 , n339 , n360 );
    xnor g690 ( n687 , n123 , n2 );
    and g691 ( n815 , n932 , n29 );
    or g692 ( n391 , n309 , n369 );
    nor g693 ( n373 , n260 , n761 );
    and g694 ( n533 , n249 , n475 );
    and g695 ( n245 , n785 , n156 );
    not g696 ( n27 , n876 );
    or g697 ( n932 , n183 , n594 );
    or g698 ( n502 , n268 , n938 );
    or g699 ( n125 , n335 , n913 );
    or g700 ( n194 , n216 , n938 );
    and g701 ( n639 , n249 , n521 );
    xnor g702 ( n459 , n98 , n289 );
    or g703 ( n293 , n686 , n369 );
    not g704 ( n7 , n541 );
    nor g705 ( n317 , n749 , n897 );
    or g706 ( n745 , n632 , n489 );
    or g707 ( n590 , n326 , n447 );
    not g708 ( n287 , n433 );
    not g709 ( n748 , n200 );
    nor g710 ( n235 , n362 , n497 );
    or g711 ( n63 , n70 , n47 );
    not g712 ( n599 , n594 );
    nor g713 ( n465 , n35 , n230 );
    buf g714 ( n215 , n901 );
    not g715 ( n572 , n184 );
    or g716 ( n635 , n890 , n739 );
    or g717 ( n346 , n678 , n365 );
endmodule
