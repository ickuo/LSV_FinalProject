// Benchmark "top" written by ABC on Sun Dec 21 18:11:57 2025

module top ( 
    n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753, n783,
    n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333, n1353,
    n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835, n1906,
    n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433, n2464,
    n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551, n2558,
    n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172, n3342,
    n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986, n3992,
    n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312, n4370,
    n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828, n4903,
    n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212, n5240,
    n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694, n5760,
    n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126, n6254,
    n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611, n6687,
    n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159, n7160,
    n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456, n7500,
    n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862, n7891,
    n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433, n8476,
    n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195, n9241,
    n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956, n10022,
    n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451, n10510,
    n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928, n10965,
    n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407, n11423,
    n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876, n11877,
    n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044, n12069,
    n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591, n12648,
    n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826, n12925,
    n12947,
    n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807  );
  input  n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753,
    n783, n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333,
    n1353, n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835,
    n1906, n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433,
    n2464, n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551,
    n2558, n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172,
    n3342, n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986,
    n3992, n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312,
    n4370, n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828,
    n4903, n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212,
    n5240, n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694,
    n5760, n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126,
    n6254, n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611,
    n6687, n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159,
    n7160, n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456,
    n7500, n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862,
    n7891, n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433,
    n8476, n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195,
    n9241, n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956,
    n10022, n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451,
    n10510, n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928,
    n10965, n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407,
    n11423, n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876,
    n11877, n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044,
    n12069, n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591,
    n12648, n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826,
    n12925, n12947;
  output n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807;
  wire new_n377, new_n378, new_n379, new_n380, new_n381_1, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397_1,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405_1, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447_1, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503_1, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521_1, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533_1, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615_1, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658_1, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671_1, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753_1, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783_1, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806_1, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837_1, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844_1, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911_1, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992_1,
    new_n993, new_n994, new_n995, new_n996_1, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020_1, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067_1, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094_1, new_n1095,
    new_n1096, new_n1097_1, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136_1, new_n1137,
    new_n1138_1, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198_1,
    new_n1199_1, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209_1, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269_1, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1311, new_n1312,
    new_n1313, new_n1314, new_n1315, new_n1316, new_n1317, new_n1318,
    new_n1319, new_n1320, new_n1321, new_n1322, new_n1323, new_n1324,
    new_n1325, new_n1326, new_n1327, new_n1328, new_n1329, new_n1330,
    new_n1331, new_n1332, new_n1333_1, new_n1334, new_n1335, new_n1336,
    new_n1337, new_n1338, new_n1339, new_n1340, new_n1341, new_n1342,
    new_n1343, new_n1344, new_n1345, new_n1346, new_n1347, new_n1348,
    new_n1349, new_n1350, new_n1351, new_n1352, new_n1353_1, new_n1354,
    new_n1355, new_n1356, new_n1357_1, new_n1358, new_n1359, new_n1360,
    new_n1361, new_n1362, new_n1363, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369, new_n1370, new_n1371, new_n1372, new_n1373,
    new_n1374, new_n1375, new_n1376, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471_1, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478_1, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510_1, new_n1511, new_n1512_1,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523_1, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1536,
    new_n1537, new_n1538, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1547, new_n1548,
    new_n1549, new_n1550, new_n1551, new_n1552, new_n1553, new_n1554,
    new_n1555, new_n1556, new_n1557, new_n1558, new_n1559, new_n1560,
    new_n1561, new_n1562, new_n1563, new_n1564_1, new_n1565, new_n1566,
    new_n1567, new_n1568, new_n1569, new_n1570, new_n1571, new_n1572,
    new_n1573, new_n1574, new_n1575, new_n1576_1, new_n1577, new_n1578,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1583, new_n1584,
    new_n1585, new_n1586, new_n1587, new_n1588, new_n1589, new_n1590,
    new_n1591, new_n1592, new_n1593, new_n1594, new_n1595, new_n1596,
    new_n1598, new_n1599, new_n1600, new_n1601, new_n1602, new_n1603,
    new_n1604, new_n1605, new_n1606, new_n1607, new_n1608, new_n1609,
    new_n1610, new_n1611, new_n1612, new_n1613, new_n1614, new_n1615,
    new_n1616, new_n1617, new_n1618, new_n1619, new_n1620, new_n1621,
    new_n1622, new_n1623, new_n1624, new_n1625, new_n1626, new_n1627,
    new_n1628, new_n1629, new_n1630, new_n1631, new_n1632, new_n1633,
    new_n1634, new_n1635, new_n1636, new_n1637, new_n1638, new_n1639,
    new_n1640, new_n1641, new_n1642, new_n1643, new_n1644, new_n1645,
    new_n1646, new_n1647, new_n1648, new_n1649, new_n1650, new_n1651,
    new_n1652, new_n1653, new_n1654, new_n1655, new_n1656, new_n1657,
    new_n1658_1, new_n1659, new_n1660, new_n1661, new_n1662, new_n1663,
    new_n1664, new_n1665, new_n1666, new_n1667, new_n1668, new_n1669,
    new_n1670, new_n1671, new_n1672, new_n1673, new_n1674, new_n1675,
    new_n1676, new_n1677, new_n1678, new_n1679, new_n1680, new_n1681,
    new_n1682, new_n1683, new_n1684, new_n1685, new_n1686, new_n1687,
    new_n1688, new_n1689, new_n1690, new_n1691, new_n1692, new_n1693,
    new_n1694, new_n1695, new_n1696, new_n1697, new_n1698, new_n1699,
    new_n1700, new_n1701, new_n1702, new_n1703, new_n1704, new_n1705,
    new_n1706, new_n1707, new_n1708, new_n1709, new_n1710, new_n1711,
    new_n1712, new_n1713, new_n1714, new_n1715, new_n1716, new_n1717,
    new_n1718, new_n1719, new_n1720, new_n1721, new_n1722, new_n1723,
    new_n1724, new_n1725, new_n1726, new_n1727, new_n1728, new_n1729,
    new_n1730, new_n1731, new_n1732, new_n1733, new_n1734, new_n1735,
    new_n1736, new_n1737, new_n1738, new_n1739, new_n1740, new_n1741,
    new_n1742, new_n1743, new_n1744, new_n1745, new_n1746, new_n1747,
    new_n1748, new_n1749, new_n1750, new_n1751, new_n1752, new_n1753,
    new_n1754, new_n1755, new_n1756, new_n1757, new_n1758, new_n1759,
    new_n1760, new_n1761, new_n1762, new_n1763, new_n1764, new_n1765,
    new_n1766, new_n1767, new_n1768, new_n1769, new_n1770, new_n1771,
    new_n1772, new_n1773, new_n1774, new_n1775, new_n1776, new_n1777,
    new_n1778, new_n1779, new_n1780, new_n1781, new_n1782, new_n1783,
    new_n1784, new_n1785, new_n1786, new_n1787, new_n1788, new_n1789,
    new_n1790, new_n1791, new_n1792, new_n1793, new_n1794, new_n1795,
    new_n1796, new_n1797, new_n1798_1, new_n1799, new_n1800, new_n1801,
    new_n1802, new_n1803, new_n1804, new_n1805, new_n1806, new_n1807,
    new_n1808, new_n1809, new_n1810, new_n1811, new_n1812, new_n1813,
    new_n1814, new_n1815, new_n1816, new_n1817, new_n1818, new_n1819,
    new_n1820, new_n1821, new_n1822, new_n1823, new_n1824, new_n1825,
    new_n1826, new_n1827, new_n1828, new_n1829, new_n1830, new_n1831,
    new_n1832, new_n1833, new_n1834, new_n1835_1, new_n1836, new_n1837,
    new_n1838, new_n1839, new_n1840, new_n1841, new_n1842, new_n1843,
    new_n1844, new_n1845, new_n1846, new_n1847_1, new_n1848, new_n1849,
    new_n1850, new_n1851, new_n1852, new_n1853, new_n1854, new_n1855,
    new_n1856, new_n1857, new_n1858, new_n1859, new_n1860, new_n1861,
    new_n1862, new_n1863, new_n1864, new_n1865, new_n1866, new_n1867,
    new_n1868, new_n1869, new_n1870, new_n1871, new_n1872, new_n1873,
    new_n1874, new_n1875, new_n1876, new_n1877, new_n1878, new_n1879,
    new_n1880, new_n1881, new_n1882, new_n1883, new_n1884, new_n1885,
    new_n1886, new_n1887, new_n1888, new_n1889, new_n1890, new_n1891,
    new_n1892, new_n1893, new_n1894, new_n1895, new_n1896, new_n1897,
    new_n1898, new_n1899, new_n1900, new_n1901, new_n1902, new_n1903,
    new_n1904, new_n1905, new_n1906_1, new_n1907, new_n1908, new_n1909,
    new_n1910, new_n1911, new_n1912, new_n1913, new_n1914, new_n1915,
    new_n1916, new_n1917, new_n1918, new_n1919, new_n1920, new_n1921,
    new_n1922, new_n1923, new_n1924, new_n1925, new_n1926, new_n1927,
    new_n1928, new_n1929, new_n1930, new_n1931, new_n1932, new_n1933,
    new_n1934, new_n1935, new_n1936, new_n1937, new_n1938, new_n1939,
    new_n1940, new_n1941, new_n1942, new_n1943, new_n1944, new_n1945,
    new_n1946, new_n1947, new_n1948, new_n1949, new_n1950, new_n1951,
    new_n1952, new_n1953, new_n1954, new_n1955, new_n1956, new_n1957,
    new_n1958, new_n1959, new_n1960, new_n1961, new_n1962, new_n1963,
    new_n1964, new_n1965, new_n1966, new_n1967, new_n1968, new_n1969,
    new_n1970, new_n1971, new_n1972, new_n1973, new_n1974, new_n1975,
    new_n1976, new_n1977, new_n1978, new_n1979, new_n1980_1, new_n1981,
    new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024_1, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087_1, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095,
    new_n2096_1, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107,
    new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113,
    new_n2114, new_n2115, new_n2116, new_n2117, new_n2118, new_n2119,
    new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125,
    new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131_1,
    new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137,
    new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143,
    new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149,
    new_n2150, new_n2151, new_n2152, new_n2153, new_n2154, new_n2155,
    new_n2156, new_n2157, new_n2158, new_n2159, new_n2160, new_n2161,
    new_n2162, new_n2163, new_n2164, new_n2165, new_n2166, new_n2167,
    new_n2168, new_n2169, new_n2170, new_n2171, new_n2172, new_n2173,
    new_n2174, new_n2175, new_n2176, new_n2177, new_n2178, new_n2179,
    new_n2180, new_n2181, new_n2182, new_n2183, new_n2184, new_n2185,
    new_n2186, new_n2187, new_n2188, new_n2189, new_n2190, new_n2191,
    new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215,
    new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2221,
    new_n2222, new_n2223, new_n2224, new_n2225, new_n2226_1, new_n2227,
    new_n2228, new_n2229, new_n2230, new_n2231, new_n2232, new_n2233,
    new_n2234, new_n2235, new_n2236, new_n2237, new_n2238, new_n2239,
    new_n2240, new_n2241, new_n2242, new_n2243, new_n2244, new_n2245,
    new_n2246, new_n2247, new_n2248, new_n2249, new_n2250, new_n2251,
    new_n2252, new_n2253_1, new_n2254, new_n2255, new_n2256, new_n2257,
    new_n2258, new_n2259, new_n2260, new_n2261, new_n2262, new_n2263,
    new_n2264, new_n2265, new_n2266, new_n2267, new_n2268, new_n2269,
    new_n2270, new_n2271, new_n2272, new_n2273, new_n2274, new_n2275,
    new_n2276, new_n2277, new_n2278_1, new_n2279, new_n2280, new_n2281,
    new_n2282, new_n2283, new_n2284, new_n2285, new_n2286, new_n2287,
    new_n2288, new_n2289, new_n2290, new_n2291, new_n2292, new_n2293,
    new_n2294, new_n2295, new_n2296, new_n2297, new_n2298, new_n2299,
    new_n2300, new_n2301_1, new_n2302, new_n2303, new_n2304, new_n2305,
    new_n2306, new_n2307, new_n2308, new_n2309, new_n2310, new_n2311,
    new_n2312, new_n2313, new_n2314, new_n2315, new_n2316_1, new_n2317,
    new_n2318, new_n2319, new_n2320, new_n2321, new_n2322, new_n2323,
    new_n2324, new_n2325, new_n2326, new_n2327, new_n2328, new_n2329,
    new_n2330, new_n2331, new_n2332, new_n2333, new_n2334, new_n2335,
    new_n2336, new_n2337, new_n2338, new_n2339, new_n2340, new_n2341,
    new_n2342, new_n2343, new_n2344, new_n2345, new_n2346, new_n2347_1,
    new_n2348, new_n2349, new_n2350, new_n2351, new_n2352, new_n2353,
    new_n2354, new_n2355, new_n2356, new_n2357, new_n2358, new_n2359,
    new_n2360, new_n2361, new_n2362, new_n2363, new_n2364, new_n2365,
    new_n2366, new_n2367, new_n2368, new_n2369, new_n2370, new_n2371,
    new_n2372, new_n2373, new_n2374, new_n2375, new_n2376, new_n2377,
    new_n2378, new_n2379, new_n2380, new_n2381, new_n2382, new_n2383_1,
    new_n2384, new_n2385, new_n2386, new_n2387, new_n2388, new_n2389,
    new_n2390, new_n2391, new_n2392, new_n2393_1, new_n2394, new_n2395,
    new_n2396, new_n2397, new_n2398, new_n2399, new_n2400, new_n2401,
    new_n2402, new_n2403, new_n2404, new_n2405, new_n2406, new_n2407,
    new_n2408, new_n2409, new_n2410, new_n2411, new_n2412, new_n2413,
    new_n2414, new_n2415, new_n2416, new_n2417, new_n2418, new_n2419,
    new_n2420, new_n2421, new_n2422, new_n2423, new_n2424, new_n2425_1,
    new_n2426, new_n2427, new_n2428, new_n2429, new_n2430, new_n2431_1,
    new_n2432, new_n2433_1, new_n2434_1, new_n2435, new_n2436, new_n2437,
    new_n2438, new_n2439, new_n2440, new_n2441, new_n2442, new_n2443,
    new_n2444, new_n2445, new_n2446, new_n2447, new_n2448, new_n2449,
    new_n2450, new_n2451, new_n2452, new_n2453, new_n2454, new_n2455,
    new_n2456, new_n2457, new_n2458, new_n2459, new_n2460, new_n2461,
    new_n2462, new_n2463, new_n2464_1, new_n2465, new_n2466, new_n2467,
    new_n2468, new_n2469, new_n2470, new_n2471, new_n2472, new_n2473,
    new_n2474, new_n2475, new_n2476, new_n2477, new_n2478, new_n2479,
    new_n2480, new_n2481, new_n2482, new_n2483, new_n2484, new_n2485,
    new_n2486, new_n2487, new_n2488, new_n2489, new_n2490, new_n2491,
    new_n2492, new_n2493, new_n2494, new_n2495, new_n2496, new_n2497,
    new_n2498_1, new_n2499, new_n2500, new_n2501, new_n2502, new_n2503,
    new_n2504, new_n2505, new_n2506, new_n2507_1, new_n2508_1, new_n2509_1,
    new_n2510, new_n2511, new_n2512_1, new_n2513, new_n2514, new_n2515_1,
    new_n2516, new_n2517, new_n2518, new_n2519, new_n2520, new_n2521,
    new_n2522_1, new_n2523, new_n2524, new_n2525, new_n2526, new_n2527,
    new_n2528, new_n2529, new_n2530_1, new_n2531, new_n2532, new_n2533,
    new_n2534, new_n2535, new_n2536, new_n2537, new_n2538, new_n2539,
    new_n2540, new_n2541, new_n2542, new_n2543, new_n2544, new_n2545,
    new_n2546, new_n2547, new_n2548, new_n2549, new_n2550, new_n2551_1,
    new_n2552, new_n2553, new_n2554, new_n2555, new_n2556, new_n2557,
    new_n2558_1, new_n2559, new_n2560, new_n2561, new_n2562, new_n2563,
    new_n2564_1, new_n2565, new_n2566, new_n2567, new_n2568, new_n2569,
    new_n2570, new_n2571, new_n2572, new_n2573, new_n2574, new_n2575,
    new_n2576, new_n2577_1, new_n2578, new_n2579, new_n2580, new_n2581_1,
    new_n2582, new_n2583, new_n2584, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624_1,
    new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679_1, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696,
    new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702,
    new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708_1,
    new_n2709, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2720,
    new_n2721, new_n2722, new_n2723, new_n2724, new_n2725, new_n2726,
    new_n2727, new_n2728, new_n2729, new_n2730, new_n2731, new_n2732,
    new_n2733, new_n2734, new_n2735, new_n2736, new_n2737, new_n2738,
    new_n2739, new_n2740, new_n2741, new_n2742, new_n2743, new_n2744,
    new_n2745, new_n2746, new_n2747, new_n2748, new_n2749_1, new_n2750,
    new_n2751, new_n2752, new_n2753, new_n2754, new_n2755, new_n2756,
    new_n2757, new_n2758, new_n2759, new_n2760, new_n2761, new_n2762,
    new_n2763, new_n2764, new_n2765, new_n2766, new_n2767, new_n2768,
    new_n2769, new_n2770, new_n2771, new_n2772, new_n2773, new_n2774,
    new_n2775, new_n2776, new_n2777, new_n2778, new_n2779, new_n2780,
    new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792,
    new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2798,
    new_n2799, new_n2800, new_n2801, new_n2802_1, new_n2803, new_n2804,
    new_n2805, new_n2806, new_n2807, new_n2808, new_n2809, new_n2810,
    new_n2811, new_n2812, new_n2813, new_n2814, new_n2815, new_n2816,
    new_n2817, new_n2818_1, new_n2819, new_n2820, new_n2821, new_n2822,
    new_n2823, new_n2824, new_n2825, new_n2826, new_n2827, new_n2828,
    new_n2829, new_n2830, new_n2831, new_n2832, new_n2833, new_n2834,
    new_n2835, new_n2836, new_n2837, new_n2838, new_n2839, new_n2840,
    new_n2841, new_n2842, new_n2843, new_n2844, new_n2845, new_n2846,
    new_n2847, new_n2848, new_n2849, new_n2850, new_n2851, new_n2852,
    new_n2853, new_n2854, new_n2855, new_n2856, new_n2857, new_n2858,
    new_n2859, new_n2860, new_n2861, new_n2862, new_n2863, new_n2864,
    new_n2865, new_n2866, new_n2867, new_n2868, new_n2869, new_n2870,
    new_n2871, new_n2872, new_n2873, new_n2874, new_n2875, new_n2876,
    new_n2877, new_n2878, new_n2879_1, new_n2880, new_n2881, new_n2882,
    new_n2883, new_n2884, new_n2885, new_n2886, new_n2887, new_n2888,
    new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2895, new_n2896, new_n2897, new_n2898, new_n2899, new_n2900,
    new_n2901, new_n2902_1, new_n2903, new_n2904, new_n2905, new_n2906,
    new_n2907, new_n2908, new_n2909, new_n2910, new_n2911, new_n2912,
    new_n2913, new_n2914, new_n2915, new_n2916, new_n2917, new_n2918,
    new_n2919, new_n2920, new_n2921, new_n2922, new_n2923, new_n2924,
    new_n2925, new_n2926, new_n2927, new_n2928, new_n2929, new_n2930,
    new_n2931, new_n2932, new_n2933, new_n2934, new_n2935, new_n2936,
    new_n2937, new_n2938, new_n2939, new_n2940, new_n2941, new_n2942,
    new_n2943, new_n2944, new_n2945, new_n2946, new_n2947, new_n2948,
    new_n2949, new_n2950, new_n2951, new_n2952, new_n2953, new_n2954,
    new_n2955, new_n2956, new_n2957, new_n2958, new_n2959, new_n2960,
    new_n2961, new_n2962, new_n2963, new_n2964, new_n2965, new_n2966,
    new_n2967, new_n2968, new_n2969, new_n2970, new_n2971, new_n2972,
    new_n2973, new_n2974, new_n2975, new_n2976, new_n2977, new_n2978,
    new_n2979, new_n2980, new_n2981, new_n2982, new_n2983, new_n2984,
    new_n2985, new_n2986, new_n2987, new_n2988, new_n2989, new_n2990,
    new_n2991, new_n2992, new_n2993, new_n2994, new_n2995, new_n2996,
    new_n2997, new_n2998, new_n2999, new_n3000, new_n3001, new_n3002,
    new_n3003, new_n3004, new_n3005, new_n3006, new_n3007, new_n3008,
    new_n3009, new_n3010, new_n3011, new_n3012, new_n3013, new_n3014,
    new_n3015, new_n3016, new_n3017, new_n3018, new_n3019, new_n3020,
    new_n3021, new_n3022_1, new_n3023, new_n3024, new_n3025, new_n3026,
    new_n3027, new_n3028, new_n3029, new_n3030, new_n3031, new_n3032,
    new_n3033, new_n3034, new_n3035, new_n3036, new_n3037, new_n3038,
    new_n3039, new_n3040, new_n3041, new_n3042, new_n3043, new_n3044,
    new_n3045, new_n3046, new_n3047, new_n3048, new_n3049, new_n3050,
    new_n3051, new_n3052, new_n3053, new_n3054, new_n3055, new_n3056,
    new_n3057, new_n3058, new_n3059, new_n3060, new_n3061, new_n3062,
    new_n3063, new_n3064, new_n3065, new_n3066, new_n3067, new_n3068,
    new_n3069, new_n3070, new_n3071_1, new_n3072, new_n3073, new_n3074,
    new_n3075, new_n3076, new_n3077, new_n3078, new_n3079, new_n3080,
    new_n3081, new_n3082, new_n3083, new_n3084, new_n3085, new_n3086,
    new_n3087, new_n3088, new_n3089, new_n3090, new_n3091, new_n3092,
    new_n3093, new_n3094, new_n3095, new_n3096, new_n3097, new_n3098,
    new_n3099, new_n3100, new_n3101, new_n3102, new_n3103, new_n3104,
    new_n3105, new_n3106, new_n3107, new_n3108, new_n3109, new_n3110,
    new_n3111, new_n3112, new_n3113, new_n3114, new_n3115, new_n3116,
    new_n3117, new_n3118, new_n3119, new_n3120, new_n3121, new_n3122,
    new_n3123, new_n3124_1, new_n3125, new_n3126, new_n3127, new_n3128,
    new_n3129, new_n3130, new_n3131, new_n3132, new_n3133, new_n3134,
    new_n3135, new_n3136, new_n3137, new_n3138, new_n3139, new_n3140,
    new_n3141, new_n3142, new_n3143, new_n3144, new_n3145, new_n3146_1,
    new_n3147, new_n3148, new_n3149, new_n3150, new_n3151, new_n3152,
    new_n3153, new_n3154, new_n3155, new_n3156, new_n3157, new_n3158,
    new_n3159, new_n3160, new_n3161, new_n3162, new_n3163, new_n3164,
    new_n3165, new_n3166, new_n3167, new_n3168, new_n3169, new_n3170,
    new_n3171, new_n3172_1, new_n3173, new_n3174, new_n3175, new_n3176,
    new_n3177, new_n3178, new_n3179, new_n3180, new_n3181, new_n3182,
    new_n3183, new_n3184, new_n3185, new_n3186, new_n3187, new_n3188,
    new_n3189, new_n3190, new_n3191, new_n3192, new_n3193, new_n3194,
    new_n3195, new_n3196, new_n3197, new_n3198, new_n3199, new_n3200,
    new_n3201, new_n3202, new_n3203, new_n3204, new_n3205, new_n3206,
    new_n3207, new_n3208, new_n3209, new_n3210, new_n3211, new_n3212,
    new_n3213, new_n3214_1, new_n3215, new_n3216, new_n3217, new_n3218,
    new_n3219, new_n3220, new_n3221, new_n3222, new_n3223, new_n3224,
    new_n3225, new_n3226, new_n3227, new_n3228, new_n3229, new_n3230_1,
    new_n3231, new_n3232, new_n3233, new_n3234, new_n3235, new_n3236,
    new_n3237, new_n3238, new_n3239, new_n3240, new_n3241, new_n3242,
    new_n3243, new_n3244, new_n3245, new_n3246, new_n3247, new_n3248,
    new_n3249, new_n3250, new_n3251, new_n3252, new_n3253, new_n3254,
    new_n3255, new_n3256, new_n3257, new_n3258, new_n3259, new_n3260,
    new_n3261, new_n3262, new_n3263, new_n3264, new_n3265, new_n3266,
    new_n3267, new_n3268, new_n3269, new_n3270, new_n3271, new_n3272_1,
    new_n3273, new_n3274, new_n3275, new_n3276, new_n3277, new_n3278,
    new_n3279, new_n3280, new_n3281, new_n3282, new_n3283, new_n3284,
    new_n3285, new_n3286, new_n3287_1, new_n3288, new_n3289, new_n3290,
    new_n3291, new_n3292, new_n3293, new_n3294, new_n3295, new_n3296,
    new_n3297, new_n3298, new_n3299, new_n3300, new_n3301, new_n3302,
    new_n3303, new_n3304, new_n3305, new_n3306, new_n3307, new_n3308,
    new_n3309, new_n3310, new_n3311, new_n3312, new_n3313, new_n3314,
    new_n3315, new_n3316, new_n3317, new_n3318, new_n3319, new_n3320,
    new_n3321, new_n3322, new_n3323, new_n3324, new_n3325, new_n3326,
    new_n3327, new_n3328, new_n3329, new_n3330, new_n3331, new_n3332,
    new_n3333, new_n3334, new_n3335, new_n3336, new_n3337, new_n3338,
    new_n3339_1, new_n3340, new_n3341, new_n3342_1, new_n3343, new_n3344,
    new_n3345, new_n3346, new_n3347, new_n3348, new_n3349, new_n3350,
    new_n3351, new_n3352, new_n3353, new_n3354, new_n3355, new_n3356,
    new_n3357, new_n3358, new_n3359, new_n3360, new_n3361, new_n3362,
    new_n3363, new_n3364, new_n3365, new_n3366, new_n3367, new_n3368,
    new_n3369, new_n3370, new_n3371, new_n3372, new_n3373, new_n3374,
    new_n3375, new_n3376, new_n3377, new_n3378, new_n3379, new_n3380,
    new_n3381, new_n3382, new_n3383, new_n3384, new_n3385, new_n3386,
    new_n3387, new_n3388, new_n3389, new_n3390, new_n3391, new_n3392,
    new_n3393, new_n3394, new_n3395, new_n3396, new_n3397, new_n3398,
    new_n3399, new_n3400, new_n3401, new_n3402, new_n3403, new_n3404,
    new_n3405, new_n3406, new_n3407, new_n3408, new_n3409, new_n3410,
    new_n3411, new_n3412, new_n3413, new_n3414, new_n3415, new_n3416,
    new_n3417, new_n3418, new_n3419, new_n3420, new_n3421, new_n3422,
    new_n3423, new_n3424, new_n3425, new_n3426, new_n3427, new_n3428,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434,
    new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451, new_n3452,
    new_n3453, new_n3454, new_n3455, new_n3456_1, new_n3457, new_n3458,
    new_n3459, new_n3460, new_n3461, new_n3462, new_n3463, new_n3464,
    new_n3465, new_n3466, new_n3467, new_n3468, new_n3469, new_n3470,
    new_n3471, new_n3472, new_n3473, new_n3474, new_n3475, new_n3476,
    new_n3477, new_n3478, new_n3479, new_n3480, new_n3481, new_n3482,
    new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488,
    new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500,
    new_n3501, new_n3502, new_n3503, new_n3504, new_n3505, new_n3506,
    new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512,
    new_n3513, new_n3514, new_n3515, new_n3516, new_n3517, new_n3518,
    new_n3519, new_n3520, new_n3521, new_n3522, new_n3523, new_n3524,
    new_n3525, new_n3526, new_n3527, new_n3528, new_n3529, new_n3530,
    new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561, new_n3562, new_n3563, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582, new_n3584, new_n3585,
    new_n3586, new_n3587, new_n3588, new_n3589, new_n3590, new_n3591,
    new_n3592, new_n3593, new_n3594, new_n3595, new_n3596, new_n3597,
    new_n3598, new_n3599, new_n3600, new_n3601, new_n3602_1, new_n3603,
    new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609,
    new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615,
    new_n3616_1, new_n3617, new_n3618, new_n3619, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627_1,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639,
    new_n3640, new_n3641, new_n3642, new_n3643, new_n3644, new_n3645,
    new_n3646, new_n3647, new_n3648, new_n3649, new_n3650, new_n3651,
    new_n3652, new_n3653, new_n3654_1, new_n3655, new_n3656, new_n3657,
    new_n3658, new_n3659, new_n3660, new_n3661_1, new_n3662, new_n3663,
    new_n3664, new_n3665, new_n3666, new_n3667, new_n3668, new_n3669,
    new_n3670, new_n3671, new_n3672, new_n3673, new_n3674, new_n3675,
    new_n3676, new_n3677_1, new_n3678, new_n3679, new_n3680, new_n3681,
    new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687,
    new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693,
    new_n3694, new_n3695, new_n3696, new_n3697, new_n3698, new_n3699,
    new_n3700, new_n3701, new_n3702, new_n3703, new_n3704, new_n3705,
    new_n3706, new_n3707, new_n3708, new_n3709, new_n3710, new_n3711,
    new_n3712, new_n3713, new_n3714, new_n3715, new_n3716, new_n3717,
    new_n3718, new_n3719_1, new_n3720, new_n3721, new_n3722, new_n3723,
    new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754_1, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759,
    new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783,
    new_n3784, new_n3785, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794, new_n3795,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825,
    new_n3826, new_n3827, new_n3828, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842_1, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849_1,
    new_n3850, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865_1, new_n3866, new_n3867,
    new_n3868, new_n3869, new_n3870, new_n3871, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891,
    new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897,
    new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903,
    new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909,
    new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925, new_n3926, new_n3927,
    new_n3928, new_n3929, new_n3930, new_n3931, new_n3932_1, new_n3933,
    new_n3934, new_n3935, new_n3936, new_n3937, new_n3938, new_n3939,
    new_n3940, new_n3941, new_n3942, new_n3943, new_n3944, new_n3945,
    new_n3946, new_n3947, new_n3948, new_n3949, new_n3950, new_n3951,
    new_n3952, new_n3953, new_n3954, new_n3955, new_n3956, new_n3957,
    new_n3958, new_n3959, new_n3960, new_n3961, new_n3962, new_n3963,
    new_n3964, new_n3965, new_n3966, new_n3967, new_n3968, new_n3969,
    new_n3970, new_n3971, new_n3972, new_n3973, new_n3974, new_n3975,
    new_n3976, new_n3977, new_n3978, new_n3979, new_n3980, new_n3981,
    new_n3982, new_n3983, new_n3984, new_n3985, new_n3986_1, new_n3987,
    new_n3988, new_n3989, new_n3990, new_n3991, new_n3992_1, new_n3993,
    new_n3994, new_n3995, new_n3996, new_n3997, new_n3998, new_n3999,
    new_n4000, new_n4001, new_n4002, new_n4003, new_n4004, new_n4005_1,
    new_n4006, new_n4007, new_n4008, new_n4009, new_n4010, new_n4011,
    new_n4012, new_n4013, new_n4014, new_n4015, new_n4016, new_n4017,
    new_n4018, new_n4019, new_n4020, new_n4021, new_n4022, new_n4023,
    new_n4024, new_n4025, new_n4026, new_n4027, new_n4028, new_n4029,
    new_n4030, new_n4031, new_n4032, new_n4033, new_n4034, new_n4035,
    new_n4036, new_n4037, new_n4038, new_n4039, new_n4040, new_n4041,
    new_n4042, new_n4043, new_n4044, new_n4045, new_n4046, new_n4047,
    new_n4048, new_n4049, new_n4050, new_n4051, new_n4052, new_n4053,
    new_n4054, new_n4055, new_n4056, new_n4057, new_n4058, new_n4059,
    new_n4060, new_n4061, new_n4062, new_n4063, new_n4064, new_n4065,
    new_n4066, new_n4067, new_n4068, new_n4069, new_n4070, new_n4071,
    new_n4072, new_n4073, new_n4074, new_n4075, new_n4076, new_n4077,
    new_n4078, new_n4079, new_n4080, new_n4081, new_n4082, new_n4083,
    new_n4084, new_n4085, new_n4086_1, new_n4087, new_n4088_1, new_n4089,
    new_n4090, new_n4091, new_n4092, new_n4093, new_n4094_1, new_n4095,
    new_n4096, new_n4097, new_n4098, new_n4099, new_n4100, new_n4101,
    new_n4102, new_n4103, new_n4104, new_n4105, new_n4106, new_n4107,
    new_n4108, new_n4109, new_n4110, new_n4111, new_n4112, new_n4113,
    new_n4114, new_n4115, new_n4116, new_n4117, new_n4118, new_n4119,
    new_n4120, new_n4121, new_n4122, new_n4123, new_n4124, new_n4125,
    new_n4126, new_n4127, new_n4128, new_n4129, new_n4130, new_n4131,
    new_n4132, new_n4133, new_n4134, new_n4135, new_n4136, new_n4137,
    new_n4138, new_n4139, new_n4140, new_n4141_1, new_n4142, new_n4143,
    new_n4144, new_n4145, new_n4146, new_n4147, new_n4148, new_n4149,
    new_n4150, new_n4151, new_n4152, new_n4153, new_n4154, new_n4155_1,
    new_n4156, new_n4157, new_n4158, new_n4159_1, new_n4160, new_n4161,
    new_n4162, new_n4163, new_n4164, new_n4165, new_n4166, new_n4167,
    new_n4168, new_n4169, new_n4170, new_n4171, new_n4172, new_n4173,
    new_n4174, new_n4175, new_n4176, new_n4177, new_n4178, new_n4179,
    new_n4180, new_n4181, new_n4182, new_n4183, new_n4184, new_n4185,
    new_n4186, new_n4187_1, new_n4188, new_n4189_1, new_n4190_1, new_n4191,
    new_n4192, new_n4193, new_n4194, new_n4195, new_n4196, new_n4197,
    new_n4198, new_n4199, new_n4200, new_n4201, new_n4202, new_n4203_1,
    new_n4204, new_n4205, new_n4206, new_n4207, new_n4208, new_n4209,
    new_n4210, new_n4211, new_n4212, new_n4213, new_n4214, new_n4215,
    new_n4216, new_n4217, new_n4218, new_n4219, new_n4220, new_n4221,
    new_n4222, new_n4223, new_n4224, new_n4225, new_n4226_1, new_n4227,
    new_n4228, new_n4229, new_n4230_1, new_n4231, new_n4232, new_n4233,
    new_n4234, new_n4235, new_n4236, new_n4237, new_n4238, new_n4239,
    new_n4240, new_n4241, new_n4242, new_n4243, new_n4244, new_n4245,
    new_n4246, new_n4247, new_n4248, new_n4249, new_n4250, new_n4251,
    new_n4252, new_n4253, new_n4254, new_n4255, new_n4256, new_n4257,
    new_n4258, new_n4259, new_n4260, new_n4261, new_n4262, new_n4263,
    new_n4264, new_n4265, new_n4266, new_n4267, new_n4268, new_n4269,
    new_n4270, new_n4271, new_n4272, new_n4273, new_n4274, new_n4275,
    new_n4276, new_n4277, new_n4278, new_n4279, new_n4280, new_n4281,
    new_n4282, new_n4283, new_n4284, new_n4285, new_n4286, new_n4287,
    new_n4288, new_n4289, new_n4290, new_n4291, new_n4292, new_n4293,
    new_n4294, new_n4295, new_n4296, new_n4297, new_n4298, new_n4299,
    new_n4300_1, new_n4301, new_n4302, new_n4303, new_n4304, new_n4305,
    new_n4306, new_n4307, new_n4308, new_n4309, new_n4310, new_n4311,
    new_n4312_1, new_n4313, new_n4314, new_n4315, new_n4316, new_n4317,
    new_n4318, new_n4319, new_n4320, new_n4321, new_n4322, new_n4323,
    new_n4324, new_n4325, new_n4326_1, new_n4327, new_n4328, new_n4329,
    new_n4330, new_n4332, new_n4333_1, new_n4334, new_n4335, new_n4336,
    new_n4337, new_n4338, new_n4339, new_n4340, new_n4341, new_n4342,
    new_n4343, new_n4344, new_n4345, new_n4346, new_n4347, new_n4348,
    new_n4349, new_n4350, new_n4351, new_n4352, new_n4353, new_n4354,
    new_n4355, new_n4356, new_n4357, new_n4358, new_n4359, new_n4360,
    new_n4361, new_n4362, new_n4363, new_n4364, new_n4365, new_n4366,
    new_n4367, new_n4368, new_n4369, new_n4370_1, new_n4371, new_n4372,
    new_n4373, new_n4374, new_n4375, new_n4376, new_n4377, new_n4378_1,
    new_n4379, new_n4380, new_n4381, new_n4382, new_n4383, new_n4384,
    new_n4385, new_n4386, new_n4387, new_n4388, new_n4389, new_n4390,
    new_n4391, new_n4392, new_n4393, new_n4394, new_n4395, new_n4396,
    new_n4397_1, new_n4398, new_n4399, new_n4400, new_n4401, new_n4402,
    new_n4403, new_n4404, new_n4405, new_n4406, new_n4407, new_n4408,
    new_n4409, new_n4410, new_n4411, new_n4412, new_n4413, new_n4414,
    new_n4415, new_n4416, new_n4417, new_n4418, new_n4419, new_n4420,
    new_n4421, new_n4422, new_n4423, new_n4424, new_n4425, new_n4426,
    new_n4427, new_n4428, new_n4429, new_n4430, new_n4431, new_n4432,
    new_n4433, new_n4434, new_n4435, new_n4436_1, new_n4437, new_n4438,
    new_n4439, new_n4440, new_n4441, new_n4442, new_n4443, new_n4444,
    new_n4445, new_n4446, new_n4447, new_n4448, new_n4449, new_n4450,
    new_n4451, new_n4452, new_n4453, new_n4454, new_n4455, new_n4456,
    new_n4457, new_n4458, new_n4459, new_n4460, new_n4461, new_n4462,
    new_n4463, new_n4464, new_n4465, new_n4466, new_n4467, new_n4468,
    new_n4469, new_n4470, new_n4471, new_n4472, new_n4473, new_n4474,
    new_n4475, new_n4476, new_n4477, new_n4478, new_n4479, new_n4480,
    new_n4481, new_n4482, new_n4483, new_n4484, new_n4485, new_n4486,
    new_n4487, new_n4488, new_n4489, new_n4490, new_n4491, new_n4492,
    new_n4493, new_n4494, new_n4495, new_n4496, new_n4497, new_n4498,
    new_n4499_1, new_n4500, new_n4501, new_n4502, new_n4503, new_n4504,
    new_n4505, new_n4506, new_n4507, new_n4508, new_n4509, new_n4510,
    new_n4511, new_n4512, new_n4513, new_n4514, new_n4515, new_n4516_1,
    new_n4517, new_n4518, new_n4519, new_n4520, new_n4521, new_n4522,
    new_n4523, new_n4524, new_n4525, new_n4526, new_n4527, new_n4528,
    new_n4529, new_n4530, new_n4531, new_n4532, new_n4533, new_n4534,
    new_n4535, new_n4536, new_n4537, new_n4538, new_n4539, new_n4540,
    new_n4541, new_n4542, new_n4543, new_n4544, new_n4545, new_n4546,
    new_n4547, new_n4548, new_n4549, new_n4550, new_n4551, new_n4553_1,
    new_n4554, new_n4555, new_n4556, new_n4557, new_n4558, new_n4559,
    new_n4560, new_n4561, new_n4562, new_n4563, new_n4564, new_n4565,
    new_n4566, new_n4567, new_n4568, new_n4569, new_n4570, new_n4571,
    new_n4572, new_n4573, new_n4574, new_n4575, new_n4576, new_n4577,
    new_n4578, new_n4579, new_n4580, new_n4581, new_n4582, new_n4583,
    new_n4584, new_n4585, new_n4586, new_n4587, new_n4588, new_n4589,
    new_n4590, new_n4591, new_n4592, new_n4593, new_n4594, new_n4595,
    new_n4596, new_n4597, new_n4598, new_n4599, new_n4600, new_n4601,
    new_n4602, new_n4603, new_n4604, new_n4605, new_n4606, new_n4607,
    new_n4608, new_n4609, new_n4610, new_n4611, new_n4612, new_n4613,
    new_n4614, new_n4615, new_n4616, new_n4617, new_n4618, new_n4619,
    new_n4620, new_n4621, new_n4622, new_n4623, new_n4624, new_n4625,
    new_n4626, new_n4627, new_n4628, new_n4629, new_n4630, new_n4631,
    new_n4632, new_n4633, new_n4634_1, new_n4635, new_n4636, new_n4637,
    new_n4638, new_n4639, new_n4640, new_n4641, new_n4642, new_n4643,
    new_n4644, new_n4645, new_n4646, new_n4647, new_n4648, new_n4649,
    new_n4650, new_n4651, new_n4652, new_n4653, new_n4654, new_n4655,
    new_n4656, new_n4657, new_n4658, new_n4659, new_n4660, new_n4661,
    new_n4662, new_n4663, new_n4664, new_n4665, new_n4666, new_n4667,
    new_n4668, new_n4669, new_n4670, new_n4671, new_n4672, new_n4673,
    new_n4674, new_n4675, new_n4676, new_n4677, new_n4678, new_n4679,
    new_n4680, new_n4681, new_n4682, new_n4683, new_n4684, new_n4685,
    new_n4686_1, new_n4687, new_n4688, new_n4689_1, new_n4690, new_n4691,
    new_n4692, new_n4693, new_n4694, new_n4695, new_n4696, new_n4697,
    new_n4698, new_n4699, new_n4700, new_n4701, new_n4702, new_n4703,
    new_n4704, new_n4705, new_n4706, new_n4707, new_n4708, new_n4709,
    new_n4710, new_n4711, new_n4712, new_n4713, new_n4714, new_n4715,
    new_n4716, new_n4717, new_n4718, new_n4719, new_n4720, new_n4721,
    new_n4722_1, new_n4723, new_n4724, new_n4725, new_n4726, new_n4727,
    new_n4728, new_n4729, new_n4730, new_n4731, new_n4732, new_n4733_1,
    new_n4734, new_n4735, new_n4736, new_n4737, new_n4738, new_n4739,
    new_n4740, new_n4741, new_n4742, new_n4743, new_n4744, new_n4745,
    new_n4746, new_n4747, new_n4748, new_n4749, new_n4750, new_n4751,
    new_n4752, new_n4753, new_n4754, new_n4755, new_n4756, new_n4757_1,
    new_n4758, new_n4759, new_n4760, new_n4761, new_n4762, new_n4763,
    new_n4764, new_n4765, new_n4766, new_n4767, new_n4768, new_n4769,
    new_n4770, new_n4771, new_n4772, new_n4773, new_n4774, new_n4775,
    new_n4776, new_n4777, new_n4778, new_n4779, new_n4780, new_n4781,
    new_n4782, new_n4783, new_n4784, new_n4785, new_n4786, new_n4787,
    new_n4788, new_n4789, new_n4790, new_n4791, new_n4792, new_n4793,
    new_n4794, new_n4795, new_n4796, new_n4797, new_n4798, new_n4799,
    new_n4800, new_n4801, new_n4802, new_n4803, new_n4804, new_n4805_1,
    new_n4806, new_n4807, new_n4808, new_n4809, new_n4810, new_n4811,
    new_n4812, new_n4813, new_n4814, new_n4815, new_n4816, new_n4817_1,
    new_n4818, new_n4819, new_n4820, new_n4821, new_n4822, new_n4823,
    new_n4824, new_n4825, new_n4826_1, new_n4827, new_n4828_1, new_n4829,
    new_n4830, new_n4831, new_n4832, new_n4833, new_n4834, new_n4835,
    new_n4836, new_n4837, new_n4838, new_n4839, new_n4840, new_n4841,
    new_n4842, new_n4843, new_n4844, new_n4845, new_n4846, new_n4847,
    new_n4848, new_n4849, new_n4850, new_n4851, new_n4852, new_n4853,
    new_n4854, new_n4855, new_n4856, new_n4857, new_n4858, new_n4859,
    new_n4860, new_n4861, new_n4862, new_n4863, new_n4864, new_n4865,
    new_n4866, new_n4867, new_n4868, new_n4869, new_n4870, new_n4871,
    new_n4872, new_n4873, new_n4874, new_n4875, new_n4876, new_n4877,
    new_n4878, new_n4879, new_n4880, new_n4881, new_n4882, new_n4883,
    new_n4884, new_n4885, new_n4886, new_n4887, new_n4888, new_n4889,
    new_n4890, new_n4891, new_n4892, new_n4893, new_n4894, new_n4895,
    new_n4896, new_n4897, new_n4898, new_n4899, new_n4900, new_n4901,
    new_n4902, new_n4903_1, new_n4904, new_n4905, new_n4906, new_n4907,
    new_n4908, new_n4909, new_n4910, new_n4911, new_n4912, new_n4913,
    new_n4915, new_n4916, new_n4917, new_n4918, new_n4919, new_n4920,
    new_n4921_1, new_n4922, new_n4923, new_n4924, new_n4925, new_n4926,
    new_n4928_1, new_n4929, new_n4930, new_n4932, new_n4933, new_n4934,
    new_n4936, new_n4937, new_n4938_1, new_n4939, new_n4940, new_n4941,
    new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947,
    new_n4948, new_n4949, new_n4950, new_n4951, new_n4952, new_n4953,
    new_n4954, new_n4955, new_n4956, new_n4957, new_n4958, new_n4959,
    new_n4960, new_n4961, new_n4962, new_n4963, new_n4964, new_n4965,
    new_n4966, new_n4967, new_n4968, new_n4969, new_n4970_1, new_n4971_1,
    new_n4972, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983,
    new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989,
    new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020, new_n5021, new_n5022, new_n5023, new_n5024, new_n5025,
    new_n5026, new_n5027, new_n5028, new_n5029, new_n5030_1, new_n5031,
    new_n5032, new_n5033, new_n5034_1, new_n5035, new_n5036, new_n5037,
    new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043,
    new_n5044, new_n5045, new_n5046, new_n5047, new_n5048, new_n5049,
    new_n5050, new_n5051, new_n5052, new_n5053, new_n5054, new_n5055,
    new_n5056, new_n5057, new_n5058, new_n5059, new_n5060, new_n5061,
    new_n5062, new_n5063, new_n5064, new_n5065, new_n5066, new_n5067,
    new_n5068, new_n5069_1, new_n5070, new_n5071, new_n5072, new_n5073,
    new_n5074, new_n5075, new_n5076, new_n5077, new_n5078, new_n5079,
    new_n5080, new_n5081, new_n5082, new_n5083, new_n5084, new_n5085,
    new_n5086, new_n5087, new_n5088, new_n5089, new_n5090, new_n5091,
    new_n5092, new_n5093, new_n5094_1, new_n5095, new_n5096, new_n5097,
    new_n5098, new_n5099, new_n5100, new_n5101, new_n5102, new_n5103,
    new_n5104, new_n5105_1, new_n5106, new_n5107, new_n5108, new_n5109,
    new_n5110, new_n5111, new_n5112, new_n5113, new_n5114, new_n5115,
    new_n5116, new_n5117, new_n5118, new_n5119, new_n5120, new_n5121,
    new_n5122, new_n5123, new_n5124, new_n5125, new_n5126, new_n5127,
    new_n5128, new_n5129, new_n5130, new_n5131, new_n5132_1, new_n5133,
    new_n5134, new_n5135, new_n5136, new_n5137, new_n5138, new_n5139,
    new_n5140, new_n5141, new_n5142, new_n5143, new_n5144, new_n5145,
    new_n5146, new_n5147, new_n5148, new_n5149, new_n5150, new_n5151,
    new_n5152, new_n5153_1, new_n5154, new_n5155, new_n5156, new_n5157,
    new_n5158, new_n5159, new_n5160, new_n5161, new_n5162, new_n5163,
    new_n5164, new_n5165, new_n5166, new_n5167, new_n5168, new_n5169,
    new_n5170, new_n5171, new_n5172, new_n5173, new_n5174, new_n5175,
    new_n5176, new_n5177, new_n5178, new_n5179, new_n5180, new_n5181,
    new_n5182, new_n5183, new_n5184, new_n5185, new_n5186, new_n5187,
    new_n5188, new_n5189, new_n5190, new_n5191_1, new_n5192, new_n5193,
    new_n5194, new_n5195, new_n5196, new_n5197, new_n5198_1, new_n5199,
    new_n5200, new_n5201, new_n5202, new_n5203, new_n5204, new_n5205,
    new_n5206, new_n5207, new_n5208, new_n5209, new_n5210, new_n5211,
    new_n5212_1, new_n5213, new_n5214, new_n5215, new_n5216, new_n5217,
    new_n5218, new_n5219, new_n5220, new_n5221, new_n5222, new_n5223,
    new_n5224, new_n5225, new_n5226, new_n5227, new_n5228, new_n5229,
    new_n5230, new_n5231, new_n5232, new_n5233, new_n5234, new_n5235,
    new_n5236, new_n5237, new_n5238, new_n5239, new_n5240_1, new_n5241,
    new_n5242, new_n5243, new_n5244, new_n5245, new_n5246, new_n5247,
    new_n5248, new_n5249, new_n5250, new_n5251, new_n5252, new_n5253,
    new_n5254, new_n5255, new_n5256, new_n5257_1, new_n5258, new_n5259,
    new_n5260, new_n5261, new_n5262, new_n5263, new_n5264, new_n5265,
    new_n5266, new_n5267, new_n5268, new_n5269, new_n5270, new_n5271,
    new_n5272, new_n5273, new_n5274, new_n5275, new_n5276, new_n5277,
    new_n5278, new_n5279, new_n5280, new_n5281, new_n5282, new_n5283_1,
    new_n5284, new_n5285, new_n5286, new_n5287, new_n5288, new_n5289,
    new_n5290, new_n5291, new_n5292, new_n5293, new_n5294, new_n5295,
    new_n5296, new_n5297, new_n5298, new_n5299, new_n5300, new_n5301,
    new_n5302, new_n5303, new_n5304, new_n5305_1, new_n5306, new_n5307,
    new_n5308, new_n5309, new_n5310, new_n5311, new_n5312, new_n5313,
    new_n5314_1, new_n5315, new_n5316, new_n5317, new_n5318, new_n5319_1,
    new_n5320_1, new_n5321, new_n5322, new_n5323, new_n5324, new_n5325,
    new_n5326, new_n5327, new_n5328, new_n5329, new_n5330, new_n5331_1,
    new_n5332, new_n5333, new_n5334, new_n5335, new_n5336, new_n5337,
    new_n5338, new_n5339, new_n5340, new_n5341, new_n5342, new_n5343,
    new_n5344, new_n5345, new_n5346, new_n5347, new_n5348, new_n5349,
    new_n5350, new_n5351, new_n5352, new_n5353, new_n5354, new_n5355,
    new_n5356, new_n5357, new_n5358, new_n5359, new_n5360, new_n5361,
    new_n5362, new_n5363, new_n5364, new_n5365, new_n5366, new_n5367,
    new_n5368, new_n5369, new_n5370, new_n5371, new_n5372, new_n5373,
    new_n5374, new_n5375, new_n5376, new_n5377, new_n5378, new_n5379,
    new_n5380, new_n5381, new_n5382, new_n5383, new_n5384, new_n5385,
    new_n5386, new_n5387, new_n5388, new_n5389, new_n5390, new_n5391,
    new_n5392, new_n5393, new_n5394, new_n5395, new_n5396, new_n5397,
    new_n5398, new_n5399, new_n5400, new_n5401, new_n5402, new_n5403,
    new_n5404, new_n5405, new_n5406, new_n5407, new_n5408, new_n5409,
    new_n5410, new_n5411_1, new_n5412, new_n5413, new_n5414, new_n5415,
    new_n5416, new_n5417, new_n5418, new_n5419, new_n5420, new_n5421,
    new_n5422, new_n5423, new_n5424, new_n5425, new_n5426, new_n5427,
    new_n5428, new_n5429, new_n5430, new_n5431, new_n5432, new_n5433,
    new_n5434, new_n5435_1, new_n5436, new_n5437, new_n5438, new_n5439,
    new_n5440, new_n5441, new_n5442, new_n5443, new_n5444, new_n5445,
    new_n5446, new_n5447, new_n5448, new_n5449, new_n5450, new_n5451,
    new_n5452, new_n5453, new_n5454, new_n5455, new_n5456, new_n5457,
    new_n5458, new_n5459, new_n5460, new_n5461, new_n5462, new_n5463,
    new_n5464, new_n5465, new_n5466, new_n5467, new_n5468, new_n5469,
    new_n5470, new_n5471, new_n5472, new_n5473, new_n5474, new_n5475,
    new_n5476, new_n5477, new_n5478, new_n5479, new_n5480, new_n5481,
    new_n5482, new_n5483, new_n5484, new_n5485, new_n5486, new_n5487,
    new_n5488, new_n5489, new_n5490, new_n5491, new_n5492, new_n5493,
    new_n5494, new_n5495, new_n5496, new_n5497, new_n5498, new_n5499,
    new_n5500, new_n5501, new_n5502, new_n5503, new_n5504, new_n5505,
    new_n5506, new_n5507, new_n5508, new_n5509, new_n5510, new_n5511,
    new_n5512, new_n5513, new_n5514, new_n5515, new_n5516, new_n5517,
    new_n5518, new_n5519, new_n5520, new_n5521, new_n5522, new_n5523,
    new_n5524, new_n5525, new_n5526, new_n5527, new_n5528, new_n5529,
    new_n5530, new_n5531, new_n5532, new_n5533, new_n5534, new_n5535,
    new_n5536, new_n5537, new_n5538, new_n5539, new_n5540, new_n5541,
    new_n5542, new_n5543, new_n5544, new_n5545, new_n5546, new_n5547,
    new_n5548, new_n5549, new_n5550, new_n5551, new_n5552, new_n5553,
    new_n5554, new_n5555, new_n5556, new_n5557, new_n5558, new_n5559,
    new_n5560, new_n5561, new_n5562, new_n5563, new_n5564, new_n5565,
    new_n5566, new_n5567, new_n5568, new_n5569, new_n5570, new_n5571,
    new_n5572, new_n5573, new_n5574, new_n5575, new_n5576, new_n5577,
    new_n5578, new_n5579_1, new_n5580, new_n5581, new_n5582, new_n5583,
    new_n5584, new_n5585, new_n5586, new_n5587, new_n5588, new_n5589,
    new_n5590, new_n5591, new_n5592, new_n5593, new_n5594, new_n5595,
    new_n5596, new_n5597, new_n5598, new_n5599, new_n5600, new_n5601,
    new_n5602, new_n5603, new_n5604, new_n5605, new_n5606, new_n5607,
    new_n5608, new_n5609, new_n5610, new_n5611, new_n5612, new_n5613,
    new_n5614, new_n5615, new_n5616, new_n5617, new_n5618, new_n5619,
    new_n5620, new_n5621, new_n5622, new_n5623, new_n5624, new_n5625,
    new_n5626, new_n5627, new_n5628, new_n5629, new_n5630, new_n5631,
    new_n5632, new_n5633, new_n5634, new_n5635, new_n5636, new_n5637,
    new_n5638, new_n5639, new_n5640, new_n5641_1, new_n5642, new_n5643,
    new_n5644, new_n5645_1, new_n5646, new_n5647, new_n5648, new_n5649,
    new_n5650, new_n5651, new_n5652, new_n5653, new_n5654, new_n5655,
    new_n5656, new_n5657, new_n5658, new_n5659, new_n5660, new_n5661,
    new_n5662, new_n5663, new_n5664, new_n5665, new_n5666, new_n5667,
    new_n5668, new_n5669, new_n5670_1, new_n5671, new_n5672, new_n5673,
    new_n5674, new_n5675, new_n5676, new_n5677, new_n5678, new_n5679,
    new_n5680, new_n5681, new_n5682, new_n5683, new_n5684, new_n5685,
    new_n5686, new_n5687, new_n5688, new_n5689, new_n5690, new_n5691,
    new_n5692, new_n5693_1, new_n5694_1, new_n5695, new_n5696, new_n5697,
    new_n5698, new_n5699, new_n5700, new_n5701, new_n5702, new_n5703,
    new_n5704, new_n5705, new_n5706, new_n5707, new_n5708, new_n5709,
    new_n5710, new_n5711, new_n5712, new_n5713, new_n5714, new_n5715,
    new_n5716, new_n5717, new_n5718, new_n5719, new_n5720, new_n5721,
    new_n5722, new_n5723, new_n5724, new_n5725, new_n5726, new_n5727,
    new_n5728, new_n5729, new_n5730, new_n5731, new_n5732, new_n5733,
    new_n5734, new_n5735, new_n5736, new_n5737, new_n5738, new_n5739,
    new_n5740, new_n5741, new_n5742, new_n5743, new_n5744, new_n5745,
    new_n5746, new_n5747, new_n5748, new_n5749, new_n5750, new_n5751,
    new_n5752, new_n5753, new_n5754, new_n5755, new_n5756, new_n5757,
    new_n5758, new_n5759, new_n5760_1, new_n5761, new_n5762, new_n5763,
    new_n5764, new_n5765, new_n5766, new_n5767_1, new_n5768, new_n5769,
    new_n5770, new_n5771, new_n5772, new_n5773, new_n5774, new_n5775,
    new_n5776, new_n5777, new_n5778, new_n5779, new_n5780, new_n5781,
    new_n5782, new_n5783, new_n5784, new_n5785, new_n5786, new_n5787,
    new_n5788, new_n5789, new_n5790, new_n5791, new_n5792, new_n5793,
    new_n5794, new_n5795, new_n5796, new_n5797, new_n5798_1, new_n5799,
    new_n5800, new_n5801, new_n5802, new_n5803, new_n5804, new_n5805,
    new_n5806, new_n5807, new_n5808, new_n5809, new_n5810, new_n5811,
    new_n5812, new_n5813, new_n5814_1, new_n5815, new_n5816, new_n5817,
    new_n5818, new_n5819, new_n5820, new_n5821, new_n5822, new_n5823,
    new_n5824, new_n5825, new_n5826, new_n5827, new_n5828, new_n5829,
    new_n5830, new_n5831, new_n5832, new_n5833, new_n5834, new_n5835,
    new_n5836, new_n5837, new_n5838, new_n5839, new_n5840, new_n5841,
    new_n5842, new_n5843, new_n5844, new_n5845, new_n5846, new_n5847,
    new_n5848, new_n5849, new_n5850, new_n5851, new_n5852, new_n5853,
    new_n5854, new_n5855, new_n5856, new_n5857_1, new_n5858, new_n5859,
    new_n5860_1, new_n5861, new_n5862, new_n5863, new_n5864, new_n5865,
    new_n5866, new_n5867, new_n5868, new_n5869, new_n5870, new_n5871,
    new_n5872, new_n5873, new_n5874, new_n5875, new_n5876, new_n5877,
    new_n5878, new_n5879, new_n5880, new_n5881, new_n5882, new_n5883,
    new_n5884, new_n5885, new_n5886, new_n5887, new_n5888, new_n5889,
    new_n5890, new_n5891, new_n5892, new_n5893, new_n5894, new_n5895,
    new_n5896, new_n5897, new_n5898, new_n5899, new_n5900, new_n5901,
    new_n5902, new_n5903, new_n5904, new_n5905, new_n5906, new_n5907,
    new_n5908, new_n5909, new_n5910, new_n5911, new_n5912, new_n5913,
    new_n5914, new_n5915, new_n5916, new_n5917, new_n5918, new_n5919,
    new_n5920, new_n5921, new_n5922, new_n5923, new_n5924, new_n5925,
    new_n5926, new_n5927, new_n5928, new_n5929, new_n5930, new_n5931,
    new_n5932, new_n5933, new_n5934_1, new_n5936, new_n5937, new_n5938,
    new_n5939, new_n5940, new_n5941, new_n5942, new_n5943, new_n5944,
    new_n5945, new_n5946, new_n5947, new_n5948, new_n5949, new_n5950,
    new_n5951, new_n5952, new_n5953, new_n5954, new_n5955, new_n5956,
    new_n5957, new_n5958, new_n5959, new_n5960, new_n5961, new_n5962,
    new_n5963, new_n5964_1, new_n5965, new_n5966, new_n5967, new_n5968,
    new_n5969, new_n5970, new_n5971, new_n5972, new_n5973, new_n5974,
    new_n5975, new_n5976, new_n5977, new_n5978, new_n5979, new_n5980,
    new_n5981, new_n5982, new_n5983, new_n5984, new_n5985, new_n5986,
    new_n5987, new_n5988, new_n5989, new_n5990, new_n5991, new_n5992,
    new_n5993, new_n5994, new_n5995, new_n5996, new_n5997, new_n5998,
    new_n5999, new_n6000, new_n6001, new_n6002, new_n6003, new_n6004,
    new_n6005, new_n6006, new_n6007, new_n6008, new_n6009, new_n6010,
    new_n6011, new_n6012, new_n6013, new_n6014, new_n6015, new_n6016_1,
    new_n6017, new_n6018, new_n6019, new_n6020, new_n6021, new_n6022,
    new_n6023, new_n6024, new_n6025, new_n6026, new_n6027, new_n6028,
    new_n6029, new_n6030, new_n6031, new_n6032, new_n6033, new_n6034,
    new_n6035, new_n6036, new_n6037, new_n6038_1, new_n6039, new_n6040,
    new_n6041, new_n6042, new_n6043, new_n6044, new_n6045, new_n6046,
    new_n6047, new_n6048, new_n6049, new_n6050, new_n6051, new_n6052,
    new_n6053, new_n6054, new_n6055, new_n6056, new_n6057, new_n6058,
    new_n6059, new_n6060, new_n6061, new_n6062, new_n6063, new_n6064,
    new_n6065, new_n6066, new_n6067, new_n6068, new_n6069, new_n6070,
    new_n6071, new_n6072, new_n6073, new_n6074, new_n6075, new_n6076,
    new_n6077, new_n6078, new_n6079, new_n6080, new_n6081, new_n6082,
    new_n6083, new_n6084, new_n6085, new_n6086, new_n6087, new_n6088,
    new_n6089_1, new_n6090, new_n6091, new_n6092, new_n6093, new_n6094,
    new_n6095, new_n6096, new_n6097, new_n6098, new_n6099, new_n6100,
    new_n6101, new_n6102, new_n6103, new_n6104, new_n6105, new_n6106,
    new_n6107, new_n6108, new_n6109, new_n6110, new_n6111, new_n6112,
    new_n6113, new_n6114, new_n6115, new_n6116, new_n6117, new_n6118,
    new_n6119, new_n6120, new_n6121, new_n6122, new_n6123, new_n6124,
    new_n6125, new_n6126_1, new_n6127, new_n6128, new_n6129, new_n6130,
    new_n6131, new_n6132, new_n6133, new_n6134, new_n6135, new_n6136,
    new_n6137, new_n6138, new_n6139, new_n6140, new_n6141, new_n6142,
    new_n6143, new_n6144, new_n6145, new_n6146, new_n6147, new_n6148,
    new_n6149, new_n6150, new_n6151, new_n6152, new_n6153, new_n6154,
    new_n6155, new_n6156, new_n6157, new_n6158, new_n6159, new_n6160,
    new_n6161, new_n6162, new_n6163, new_n6164, new_n6165, new_n6166,
    new_n6167, new_n6168, new_n6169, new_n6170, new_n6171, new_n6172,
    new_n6173, new_n6174, new_n6175, new_n6176, new_n6177, new_n6178,
    new_n6179, new_n6180, new_n6181, new_n6182, new_n6183, new_n6184,
    new_n6185, new_n6186, new_n6187, new_n6188, new_n6189, new_n6190,
    new_n6191, new_n6192_1, new_n6193, new_n6194, new_n6195, new_n6196,
    new_n6197, new_n6198, new_n6199, new_n6200, new_n6201, new_n6202,
    new_n6203, new_n6204, new_n6205, new_n6206, new_n6207, new_n6208,
    new_n6209, new_n6210, new_n6211, new_n6212, new_n6213, new_n6214,
    new_n6215, new_n6216, new_n6217, new_n6218, new_n6219, new_n6220,
    new_n6221, new_n6222, new_n6223, new_n6224, new_n6225, new_n6226,
    new_n6227, new_n6228, new_n6229, new_n6230, new_n6231, new_n6232,
    new_n6233, new_n6234, new_n6235, new_n6236, new_n6237, new_n6238,
    new_n6239, new_n6240, new_n6241, new_n6242, new_n6243, new_n6244,
    new_n6245, new_n6246, new_n6247, new_n6248, new_n6249, new_n6250,
    new_n6251, new_n6252, new_n6253, new_n6254_1, new_n6255, new_n6256,
    new_n6257, new_n6258, new_n6259, new_n6260, new_n6261, new_n6262,
    new_n6263, new_n6264, new_n6265, new_n6266, new_n6267, new_n6268,
    new_n6269, new_n6270, new_n6271, new_n6272, new_n6273_1, new_n6274,
    new_n6275, new_n6276, new_n6277, new_n6278, new_n6279, new_n6280,
    new_n6281, new_n6282, new_n6283, new_n6284, new_n6285, new_n6286,
    new_n6287, new_n6288, new_n6289, new_n6290, new_n6291, new_n6292,
    new_n6293, new_n6294_1, new_n6295, new_n6296, new_n6297, new_n6298,
    new_n6299, new_n6300, new_n6301, new_n6302, new_n6303, new_n6304,
    new_n6305, new_n6306, new_n6307, new_n6308, new_n6309, new_n6310,
    new_n6311, new_n6312, new_n6313, new_n6314, new_n6315, new_n6316,
    new_n6317, new_n6318, new_n6319, new_n6320, new_n6321, new_n6322,
    new_n6323, new_n6324, new_n6325, new_n6326, new_n6327, new_n6328,
    new_n6329, new_n6330, new_n6331, new_n6332, new_n6333, new_n6334,
    new_n6335, new_n6336, new_n6337, new_n6338, new_n6339, new_n6340,
    new_n6341, new_n6342, new_n6343, new_n6344, new_n6345, new_n6346,
    new_n6347, new_n6348, new_n6349, new_n6350, new_n6351, new_n6352,
    new_n6353, new_n6354, new_n6355, new_n6356, new_n6357, new_n6358_1,
    new_n6359_1, new_n6360, new_n6361, new_n6362, new_n6363, new_n6364,
    new_n6365, new_n6366, new_n6367, new_n6368, new_n6369, new_n6370,
    new_n6371, new_n6372, new_n6373, new_n6374, new_n6375, new_n6376,
    new_n6377, new_n6378, new_n6379, new_n6380, new_n6381, new_n6382,
    new_n6383, new_n6384, new_n6385, new_n6386, new_n6387, new_n6388,
    new_n6389, new_n6390, new_n6391, new_n6392, new_n6393, new_n6394,
    new_n6395, new_n6396, new_n6397, new_n6398, new_n6399, new_n6400,
    new_n6401, new_n6402, new_n6403, new_n6404, new_n6405, new_n6406,
    new_n6407, new_n6408, new_n6409, new_n6410, new_n6411, new_n6412,
    new_n6413, new_n6414, new_n6415, new_n6416, new_n6417, new_n6418,
    new_n6419, new_n6420, new_n6421, new_n6422, new_n6423, new_n6424,
    new_n6425, new_n6426, new_n6427, new_n6428, new_n6429_1, new_n6430,
    new_n6431_1, new_n6432, new_n6433, new_n6434, new_n6435, new_n6436,
    new_n6437, new_n6438, new_n6439, new_n6440, new_n6441_1, new_n6442,
    new_n6443, new_n6444, new_n6445_1, new_n6446, new_n6447, new_n6448,
    new_n6449, new_n6450, new_n6451, new_n6452, new_n6453, new_n6454,
    new_n6455, new_n6456, new_n6457, new_n6458, new_n6459, new_n6460,
    new_n6461, new_n6462, new_n6463, new_n6464, new_n6465, new_n6466,
    new_n6467, new_n6469, new_n6470, new_n6471, new_n6472, new_n6473,
    new_n6474, new_n6475, new_n6476, new_n6477, new_n6478, new_n6479,
    new_n6480, new_n6481, new_n6482, new_n6483, new_n6484, new_n6485,
    new_n6486, new_n6487, new_n6488, new_n6489, new_n6490, new_n6491,
    new_n6492, new_n6493, new_n6494, new_n6495, new_n6496, new_n6497,
    new_n6498, new_n6499, new_n6500, new_n6501, new_n6502, new_n6503,
    new_n6504, new_n6505, new_n6506, new_n6507, new_n6508, new_n6509,
    new_n6510, new_n6511, new_n6512, new_n6513, new_n6514, new_n6515,
    new_n6516, new_n6517, new_n6518, new_n6519, new_n6520, new_n6521,
    new_n6522, new_n6523, new_n6524, new_n6525, new_n6526, new_n6527,
    new_n6528, new_n6529, new_n6530, new_n6531, new_n6532, new_n6533,
    new_n6534, new_n6535, new_n6536, new_n6537, new_n6538, new_n6539,
    new_n6540, new_n6541, new_n6542, new_n6543, new_n6544, new_n6545,
    new_n6546, new_n6547, new_n6548, new_n6549, new_n6550, new_n6551,
    new_n6552, new_n6553, new_n6554, new_n6555, new_n6556, new_n6557,
    new_n6558, new_n6559, new_n6560, new_n6561, new_n6562, new_n6563,
    new_n6564, new_n6565, new_n6566, new_n6567, new_n6568, new_n6569,
    new_n6570, new_n6571, new_n6572, new_n6573, new_n6574, new_n6575,
    new_n6576, new_n6577, new_n6578_1, new_n6579, new_n6580, new_n6581,
    new_n6582, new_n6583, new_n6584, new_n6585, new_n6586, new_n6587,
    new_n6588, new_n6589, new_n6590, new_n6591, new_n6592, new_n6593,
    new_n6594, new_n6595, new_n6596, new_n6597, new_n6598, new_n6599,
    new_n6600, new_n6601, new_n6602, new_n6603, new_n6604_1, new_n6605,
    new_n6606, new_n6607, new_n6608, new_n6609, new_n6610, new_n6611_1,
    new_n6612, new_n6613, new_n6614, new_n6615, new_n6616, new_n6617,
    new_n6618, new_n6619, new_n6620, new_n6621, new_n6622, new_n6623,
    new_n6624, new_n6625, new_n6626, new_n6627, new_n6628, new_n6629,
    new_n6630, new_n6631, new_n6632, new_n6633, new_n6634, new_n6635,
    new_n6636, new_n6637, new_n6638, new_n6639, new_n6640, new_n6641,
    new_n6642, new_n6643, new_n6644, new_n6645_1, new_n6646, new_n6647,
    new_n6648, new_n6649, new_n6650, new_n6651, new_n6652, new_n6653,
    new_n6654, new_n6655, new_n6656, new_n6657, new_n6658, new_n6659,
    new_n6660, new_n6661, new_n6662, new_n6663, new_n6664, new_n6665,
    new_n6666, new_n6667, new_n6668, new_n6669, new_n6670, new_n6671,
    new_n6672, new_n6673, new_n6674, new_n6675, new_n6676, new_n6677,
    new_n6678, new_n6679, new_n6680, new_n6681, new_n6682, new_n6683,
    new_n6684, new_n6685, new_n6686, new_n6687_1, new_n6688, new_n6689_1,
    new_n6690, new_n6691, new_n6692, new_n6693, new_n6694, new_n6695,
    new_n6696, new_n6697, new_n6698, new_n6699, new_n6700, new_n6701,
    new_n6702, new_n6703_1, new_n6704, new_n6705, new_n6706, new_n6707,
    new_n6708, new_n6709, new_n6710, new_n6711, new_n6712, new_n6713,
    new_n6714, new_n6715, new_n6716, new_n6717, new_n6718, new_n6719,
    new_n6720, new_n6721, new_n6722, new_n6723, new_n6724, new_n6725,
    new_n6726, new_n6727, new_n6728, new_n6729, new_n6730, new_n6731,
    new_n6732, new_n6733, new_n6734, new_n6735, new_n6736, new_n6737,
    new_n6738, new_n6739, new_n6740, new_n6741, new_n6742_1, new_n6743,
    new_n6744, new_n6745, new_n6746, new_n6747, new_n6748, new_n6749,
    new_n6750, new_n6751, new_n6752, new_n6753, new_n6754, new_n6755,
    new_n6756, new_n6757, new_n6758, new_n6759, new_n6760, new_n6761,
    new_n6762, new_n6763, new_n6764, new_n6765, new_n6766, new_n6767,
    new_n6768, new_n6769, new_n6770_1, new_n6771, new_n6772, new_n6773,
    new_n6774, new_n6775, new_n6776_1, new_n6777, new_n6778, new_n6779,
    new_n6780, new_n6781, new_n6782, new_n6783, new_n6784, new_n6785,
    new_n6786, new_n6787, new_n6788, new_n6789, new_n6790, new_n6791,
    new_n6792, new_n6793, new_n6794, new_n6795, new_n6796, new_n6797_1,
    new_n6798, new_n6799, new_n6800, new_n6801, new_n6802, new_n6803,
    new_n6804, new_n6805, new_n6806_1, new_n6807, new_n6808, new_n6809_1,
    new_n6810, new_n6811, new_n6812, new_n6813, new_n6814, new_n6815,
    new_n6816, new_n6817, new_n6818, new_n6820, new_n6821, new_n6822_1,
    new_n6823, new_n6824, new_n6825, new_n6826_1, new_n6827, new_n6828,
    new_n6829, new_n6830, new_n6831, new_n6832, new_n6833, new_n6834,
    new_n6835, new_n6836, new_n6837, new_n6838, new_n6839, new_n6840,
    new_n6841, new_n6842, new_n6843, new_n6844, new_n6845, new_n6846,
    new_n6847, new_n6848, new_n6849, new_n6850, new_n6851, new_n6852,
    new_n6853, new_n6854, new_n6855, new_n6856, new_n6857, new_n6858,
    new_n6859, new_n6860_1, new_n6861, new_n6862, new_n6863, new_n6864,
    new_n6865, new_n6866, new_n6867, new_n6868, new_n6869, new_n6870,
    new_n6871, new_n6872, new_n6873, new_n6874, new_n6875, new_n6876,
    new_n6877_1, new_n6878, new_n6879, new_n6880, new_n6881, new_n6882,
    new_n6883, new_n6884, new_n6885, new_n6886, new_n6887, new_n6888,
    new_n6889, new_n6890, new_n6891, new_n6892, new_n6893, new_n6894,
    new_n6895, new_n6896, new_n6897, new_n6898, new_n6899, new_n6900,
    new_n6901, new_n6902, new_n6903, new_n6904, new_n6905, new_n6906,
    new_n6907, new_n6908, new_n6909, new_n6910, new_n6911, new_n6912,
    new_n6913, new_n6914, new_n6915, new_n6916, new_n6917, new_n6918,
    new_n6919, new_n6920, new_n6921, new_n6922, new_n6923, new_n6924,
    new_n6925, new_n6926, new_n6927, new_n6928, new_n6929, new_n6930,
    new_n6931, new_n6932, new_n6933, new_n6934, new_n6935, new_n6936,
    new_n6937, new_n6938, new_n6939, new_n6940, new_n6941, new_n6942,
    new_n6943, new_n6944, new_n6945, new_n6946, new_n6947, new_n6948,
    new_n6949, new_n6950, new_n6951, new_n6952, new_n6953, new_n6954,
    new_n6955, new_n6956, new_n6957, new_n6958, new_n6959, new_n6960,
    new_n6961, new_n6962, new_n6963, new_n6964, new_n6965, new_n6966,
    new_n6967, new_n6968, new_n6969, new_n6970, new_n6971, new_n6972,
    new_n6973, new_n6974, new_n6975, new_n6976, new_n6977, new_n6978,
    new_n6979, new_n6980, new_n6981, new_n6982, new_n6983, new_n6984,
    new_n6985, new_n6986_1, new_n6987, new_n6988, new_n6989, new_n6990,
    new_n6991, new_n6992, new_n6993, new_n6994, new_n6995, new_n6996,
    new_n6997, new_n6998, new_n6999, new_n7000, new_n7001, new_n7002,
    new_n7003, new_n7004, new_n7005, new_n7006, new_n7007, new_n7008,
    new_n7009, new_n7010, new_n7011, new_n7012, new_n7013, new_n7014,
    new_n7015, new_n7016, new_n7017, new_n7018, new_n7019, new_n7020,
    new_n7021, new_n7022, new_n7023, new_n7024, new_n7025, new_n7026,
    new_n7027, new_n7028, new_n7029, new_n7030, new_n7031, new_n7032,
    new_n7033, new_n7034, new_n7035, new_n7036, new_n7037, new_n7038,
    new_n7039, new_n7040, new_n7041, new_n7043, new_n7044, new_n7045,
    new_n7046, new_n7047, new_n7048, new_n7049, new_n7050, new_n7051,
    new_n7052, new_n7053, new_n7054, new_n7055, new_n7056, new_n7057,
    new_n7058, new_n7059, new_n7060, new_n7061, new_n7062, new_n7063,
    new_n7064, new_n7065, new_n7066, new_n7067, new_n7068, new_n7069,
    new_n7070, new_n7071, new_n7072, new_n7073, new_n7074, new_n7075,
    new_n7076, new_n7077, new_n7078, new_n7079, new_n7080, new_n7081,
    new_n7082, new_n7083, new_n7084, new_n7085, new_n7086, new_n7087,
    new_n7088, new_n7089, new_n7090, new_n7092, new_n7093, new_n7094,
    new_n7096, new_n7097, new_n7098, new_n7099, new_n7100, new_n7101,
    new_n7102, new_n7103, new_n7104, new_n7105, new_n7106, new_n7107,
    new_n7108, new_n7109, new_n7110, new_n7111, new_n7112, new_n7113,
    new_n7114, new_n7115, new_n7116, new_n7117, new_n7118, new_n7119,
    new_n7120, new_n7121, new_n7122, new_n7123, new_n7124, new_n7125,
    new_n7126, new_n7127, new_n7128, new_n7129, new_n7130, new_n7131,
    new_n7132, new_n7133, new_n7134, new_n7135, new_n7136, new_n7137,
    new_n7138, new_n7139, new_n7140, new_n7141, new_n7142, new_n7143,
    new_n7144, new_n7145, new_n7146, new_n7147, new_n7148, new_n7149,
    new_n7150, new_n7151, new_n7152, new_n7153, new_n7154, new_n7155,
    new_n7156, new_n7157, new_n7158, new_n7159_1, new_n7160_1, new_n7161,
    new_n7162, new_n7163, new_n7164, new_n7165, new_n7166, new_n7167,
    new_n7168, new_n7169, new_n7170, new_n7171, new_n7172, new_n7173,
    new_n7174, new_n7175, new_n7176, new_n7177, new_n7178, new_n7179,
    new_n7180, new_n7181, new_n7182, new_n7183, new_n7184, new_n7185,
    new_n7186, new_n7187, new_n7188, new_n7189, new_n7190, new_n7191,
    new_n7192, new_n7193_1, new_n7194, new_n7195, new_n7196, new_n7197,
    new_n7198, new_n7199, new_n7200, new_n7201, new_n7202, new_n7203,
    new_n7204, new_n7205, new_n7206, new_n7207, new_n7208, new_n7209,
    new_n7210, new_n7211, new_n7212, new_n7213, new_n7214, new_n7215,
    new_n7216, new_n7217, new_n7218, new_n7219, new_n7220, new_n7221,
    new_n7222, new_n7223, new_n7224, new_n7225, new_n7226, new_n7227,
    new_n7228, new_n7229, new_n7230, new_n7231, new_n7232, new_n7233,
    new_n7234, new_n7235, new_n7236_1, new_n7237, new_n7238, new_n7239,
    new_n7240, new_n7241, new_n7242, new_n7243, new_n7244, new_n7245,
    new_n7246, new_n7247, new_n7248, new_n7249, new_n7250, new_n7251,
    new_n7252, new_n7253, new_n7254, new_n7255, new_n7256, new_n7257,
    new_n7258, new_n7259, new_n7260, new_n7261, new_n7262, new_n7263,
    new_n7264, new_n7265_1, new_n7266, new_n7267, new_n7268, new_n7269,
    new_n7270_1, new_n7271, new_n7272, new_n7273, new_n7274, new_n7275,
    new_n7276, new_n7277, new_n7278, new_n7279, new_n7280, new_n7281,
    new_n7282, new_n7283, new_n7284, new_n7285, new_n7286, new_n7287,
    new_n7288, new_n7289, new_n7290, new_n7291, new_n7292, new_n7293,
    new_n7294_1, new_n7295, new_n7296, new_n7297, new_n7298, new_n7299,
    new_n7300, new_n7301, new_n7302, new_n7303, new_n7304, new_n7305,
    new_n7306, new_n7307, new_n7308, new_n7309, new_n7310, new_n7311,
    new_n7312, new_n7313, new_n7314, new_n7315, new_n7316, new_n7317,
    new_n7318, new_n7319, new_n7320_1, new_n7321, new_n7322, new_n7323,
    new_n7324, new_n7325, new_n7326, new_n7327, new_n7328, new_n7329,
    new_n7330, new_n7331, new_n7332, new_n7333, new_n7334, new_n7335,
    new_n7336, new_n7337, new_n7338, new_n7339, new_n7340, new_n7341,
    new_n7342, new_n7343, new_n7344, new_n7345, new_n7346, new_n7347,
    new_n7348, new_n7349, new_n7350, new_n7351, new_n7352, new_n7353,
    new_n7354_1, new_n7355, new_n7356, new_n7357, new_n7358, new_n7359,
    new_n7360, new_n7361, new_n7362, new_n7363, new_n7364, new_n7365,
    new_n7366, new_n7367, new_n7368, new_n7369, new_n7370, new_n7371,
    new_n7372, new_n7373, new_n7374, new_n7375, new_n7376, new_n7377,
    new_n7378, new_n7379, new_n7380, new_n7381, new_n7382, new_n7383,
    new_n7384, new_n7385, new_n7386, new_n7387, new_n7388_1, new_n7389,
    new_n7390, new_n7391, new_n7392, new_n7393, new_n7394, new_n7395,
    new_n7396, new_n7397, new_n7398, new_n7399, new_n7400, new_n7401,
    new_n7402, new_n7403, new_n7404, new_n7405, new_n7406, new_n7407,
    new_n7408, new_n7409, new_n7410, new_n7411, new_n7412, new_n7413,
    new_n7414, new_n7415, new_n7416, new_n7417, new_n7418, new_n7419,
    new_n7420, new_n7421, new_n7422, new_n7423, new_n7424, new_n7425,
    new_n7426, new_n7427, new_n7428, new_n7429, new_n7430, new_n7431,
    new_n7432, new_n7433, new_n7434, new_n7435, new_n7436_1, new_n7437,
    new_n7438, new_n7439, new_n7440, new_n7441, new_n7442, new_n7443,
    new_n7444, new_n7445, new_n7446, new_n7447, new_n7448, new_n7449,
    new_n7450, new_n7451, new_n7452, new_n7453, new_n7454, new_n7455,
    new_n7456_1, new_n7457, new_n7458, new_n7459, new_n7460, new_n7461,
    new_n7462, new_n7463, new_n7464, new_n7465, new_n7466, new_n7467,
    new_n7468, new_n7469, new_n7470, new_n7471, new_n7472, new_n7473,
    new_n7474, new_n7475, new_n7476, new_n7477, new_n7478, new_n7479,
    new_n7480, new_n7481, new_n7482, new_n7483, new_n7484, new_n7485,
    new_n7486, new_n7487, new_n7488, new_n7489, new_n7490, new_n7491,
    new_n7492, new_n7493, new_n7494, new_n7495, new_n7496, new_n7497,
    new_n7498, new_n7499, new_n7500_1, new_n7501, new_n7502, new_n7503,
    new_n7504, new_n7505, new_n7506, new_n7507, new_n7508, new_n7509,
    new_n7510, new_n7511, new_n7512, new_n7513, new_n7514, new_n7515,
    new_n7516, new_n7517, new_n7518, new_n7519, new_n7520, new_n7521,
    new_n7522, new_n7523_1, new_n7524, new_n7525, new_n7526, new_n7527,
    new_n7528, new_n7529, new_n7530, new_n7531, new_n7532, new_n7533,
    new_n7534, new_n7535, new_n7536, new_n7537, new_n7538, new_n7539,
    new_n7540, new_n7541, new_n7542, new_n7543, new_n7544, new_n7545,
    new_n7546_1, new_n7547, new_n7548, new_n7549, new_n7550, new_n7551,
    new_n7552, new_n7553, new_n7554, new_n7555, new_n7556, new_n7557,
    new_n7558, new_n7559, new_n7560, new_n7561, new_n7562, new_n7563,
    new_n7564, new_n7565, new_n7566, new_n7567, new_n7568_1, new_n7569,
    new_n7570, new_n7571, new_n7572, new_n7573, new_n7574, new_n7575,
    new_n7576, new_n7577, new_n7578, new_n7579, new_n7580, new_n7581,
    new_n7582, new_n7583, new_n7584, new_n7585, new_n7586, new_n7587,
    new_n7588, new_n7589, new_n7590, new_n7591, new_n7592, new_n7593,
    new_n7594, new_n7595, new_n7596, new_n7597, new_n7598, new_n7599,
    new_n7600, new_n7601, new_n7602, new_n7603, new_n7604, new_n7605,
    new_n7606, new_n7607, new_n7608, new_n7609, new_n7610_1, new_n7611,
    new_n7612, new_n7613, new_n7614, new_n7615, new_n7616, new_n7617,
    new_n7618, new_n7619, new_n7620, new_n7621, new_n7622, new_n7623,
    new_n7624, new_n7625, new_n7626, new_n7627, new_n7628, new_n7630,
    new_n7631, new_n7632, new_n7634, new_n7635, new_n7636, new_n7637,
    new_n7638, new_n7639, new_n7640, new_n7641, new_n7642, new_n7643,
    new_n7644, new_n7645, new_n7646_1, new_n7647, new_n7648, new_n7649,
    new_n7650, new_n7651, new_n7652, new_n7653, new_n7654, new_n7655,
    new_n7656, new_n7657, new_n7658, new_n7659, new_n7660, new_n7661,
    new_n7662, new_n7663, new_n7664, new_n7665, new_n7666, new_n7667,
    new_n7668, new_n7669, new_n7670, new_n7671, new_n7672, new_n7673,
    new_n7674, new_n7675, new_n7676_1, new_n7677, new_n7678, new_n7679,
    new_n7680, new_n7681, new_n7682, new_n7683, new_n7684, new_n7685,
    new_n7686, new_n7687, new_n7688, new_n7689, new_n7690_1, new_n7691,
    new_n7692, new_n7693, new_n7694, new_n7695, new_n7696, new_n7697,
    new_n7698, new_n7699, new_n7700, new_n7701, new_n7702, new_n7703,
    new_n7704, new_n7705, new_n7706, new_n7707, new_n7708, new_n7709,
    new_n7710, new_n7711, new_n7712, new_n7713, new_n7714, new_n7715,
    new_n7716, new_n7717, new_n7718, new_n7719, new_n7720, new_n7721,
    new_n7722, new_n7723, new_n7724, new_n7725, new_n7726, new_n7727,
    new_n7728, new_n7729, new_n7730_1, new_n7731, new_n7732, new_n7733_1,
    new_n7734, new_n7735, new_n7736, new_n7737, new_n7738, new_n7739,
    new_n7740, new_n7741, new_n7742, new_n7743, new_n7744, new_n7745,
    new_n7746, new_n7747, new_n7748, new_n7749, new_n7750, new_n7751,
    new_n7752, new_n7753, new_n7754, new_n7755, new_n7756, new_n7757,
    new_n7758, new_n7759, new_n7760, new_n7761, new_n7762, new_n7763,
    new_n7764, new_n7765, new_n7766, new_n7767, new_n7768, new_n7769,
    new_n7770, new_n7771, new_n7772, new_n7773, new_n7774, new_n7775,
    new_n7776, new_n7777, new_n7778, new_n7779, new_n7780, new_n7781,
    new_n7782, new_n7783, new_n7784, new_n7785, new_n7786, new_n7787,
    new_n7788, new_n7789, new_n7790, new_n7791, new_n7792, new_n7793,
    new_n7794, new_n7795, new_n7796, new_n7797, new_n7798, new_n7799,
    new_n7800, new_n7801, new_n7802, new_n7803, new_n7804, new_n7805,
    new_n7806, new_n7807, new_n7808, new_n7809, new_n7810, new_n7811,
    new_n7812, new_n7813, new_n7814, new_n7815, new_n7816, new_n7817,
    new_n7818, new_n7819, new_n7820, new_n7821, new_n7822, new_n7823_1,
    new_n7824, new_n7825, new_n7826, new_n7827, new_n7828, new_n7829,
    new_n7830, new_n7831, new_n7832, new_n7833, new_n7834, new_n7835,
    new_n7836, new_n7837, new_n7838, new_n7839, new_n7840, new_n7841,
    new_n7842, new_n7843, new_n7844, new_n7845, new_n7846, new_n7847,
    new_n7848, new_n7849, new_n7850, new_n7851, new_n7852, new_n7853,
    new_n7854, new_n7855, new_n7856, new_n7857, new_n7858, new_n7859,
    new_n7860, new_n7861, new_n7862_1, new_n7863, new_n7864, new_n7865,
    new_n7866, new_n7867, new_n7868, new_n7869, new_n7870, new_n7871,
    new_n7872, new_n7873, new_n7874, new_n7875, new_n7876, new_n7877,
    new_n7878, new_n7879, new_n7880, new_n7881, new_n7882, new_n7883,
    new_n7884, new_n7885, new_n7886, new_n7887, new_n7888, new_n7889,
    new_n7890, new_n7891_1, new_n7892, new_n7893, new_n7894, new_n7895,
    new_n7896, new_n7897, new_n7898, new_n7899, new_n7900, new_n7901,
    new_n7902, new_n7903, new_n7904, new_n7905, new_n7906, new_n7907,
    new_n7908, new_n7909, new_n7910, new_n7911, new_n7912, new_n7913,
    new_n7914, new_n7915, new_n7916, new_n7917, new_n7918, new_n7919,
    new_n7920, new_n7921, new_n7922, new_n7923, new_n7924, new_n7925,
    new_n7926, new_n7927, new_n7928, new_n7929, new_n7930, new_n7931,
    new_n7932, new_n7933, new_n7934, new_n7935, new_n7936, new_n7937,
    new_n7938, new_n7939, new_n7940, new_n7941, new_n7942, new_n7943,
    new_n7944, new_n7945, new_n7946_1, new_n7947, new_n7948, new_n7949,
    new_n7950, new_n7951, new_n7952, new_n7953, new_n7954, new_n7955,
    new_n7956, new_n7957, new_n7958, new_n7959, new_n7960, new_n7961,
    new_n7962, new_n7963, new_n7964, new_n7965_1, new_n7966_1, new_n7967,
    new_n7968, new_n7969, new_n7970, new_n7971, new_n7972, new_n7973,
    new_n7974, new_n7975, new_n7976, new_n7977, new_n7978, new_n7979,
    new_n7980, new_n7981_1, new_n7982, new_n7983, new_n7984, new_n7985,
    new_n7986, new_n7987, new_n7988, new_n7989, new_n7990, new_n7991,
    new_n7992, new_n7993, new_n7994, new_n7995, new_n7996, new_n7997,
    new_n7998, new_n7999, new_n8000, new_n8001, new_n8002, new_n8003,
    new_n8004, new_n8005, new_n8006, new_n8007, new_n8008, new_n8009,
    new_n8010, new_n8011, new_n8012, new_n8013, new_n8014, new_n8015,
    new_n8016, new_n8017, new_n8018, new_n8019, new_n8020, new_n8021,
    new_n8022, new_n8023, new_n8024, new_n8025, new_n8026, new_n8027,
    new_n8028_1, new_n8029, new_n8030, new_n8031, new_n8032, new_n8033,
    new_n8034, new_n8035, new_n8036, new_n8037, new_n8038, new_n8039,
    new_n8040, new_n8041, new_n8042, new_n8043, new_n8044, new_n8045,
    new_n8046, new_n8047, new_n8048, new_n8049, new_n8050, new_n8051,
    new_n8052, new_n8053, new_n8054, new_n8055, new_n8056, new_n8057,
    new_n8058, new_n8059, new_n8060, new_n8061, new_n8062, new_n8063,
    new_n8064, new_n8065_1, new_n8066, new_n8067, new_n8068, new_n8069,
    new_n8070, new_n8071, new_n8072, new_n8073, new_n8074, new_n8075,
    new_n8076, new_n8077, new_n8078, new_n8079, new_n8080, new_n8081,
    new_n8082, new_n8083, new_n8084, new_n8085, new_n8086, new_n8087,
    new_n8088, new_n8089, new_n8090, new_n8091, new_n8092, new_n8093,
    new_n8094, new_n8095, new_n8096, new_n8097, new_n8098, new_n8099,
    new_n8100_1, new_n8101, new_n8102, new_n8103, new_n8104, new_n8105,
    new_n8106, new_n8107, new_n8108, new_n8109, new_n8110, new_n8111,
    new_n8112, new_n8113, new_n8114, new_n8115, new_n8116, new_n8117,
    new_n8118, new_n8119, new_n8120, new_n8121, new_n8122, new_n8123,
    new_n8124, new_n8125, new_n8126, new_n8127, new_n8128, new_n8129,
    new_n8130, new_n8131, new_n8132, new_n8133, new_n8134, new_n8135,
    new_n8136, new_n8137, new_n8138_1, new_n8139, new_n8140, new_n8141,
    new_n8142, new_n8143, new_n8144, new_n8145, new_n8146, new_n8147,
    new_n8148, new_n8149, new_n8150, new_n8151, new_n8152, new_n8153,
    new_n8154, new_n8155, new_n8156, new_n8157, new_n8158, new_n8159,
    new_n8160, new_n8161, new_n8162, new_n8163, new_n8164, new_n8165,
    new_n8166, new_n8167, new_n8168, new_n8169, new_n8170, new_n8171,
    new_n8172, new_n8173, new_n8174, new_n8175, new_n8176, new_n8177,
    new_n8178, new_n8179, new_n8180, new_n8181, new_n8182, new_n8183,
    new_n8184, new_n8185, new_n8186, new_n8187, new_n8188, new_n8189,
    new_n8190, new_n8191, new_n8192, new_n8193, new_n8194, new_n8195,
    new_n8196, new_n8197, new_n8198, new_n8199, new_n8200, new_n8201,
    new_n8202_1, new_n8203, new_n8204, new_n8205, new_n8206, new_n8207,
    new_n8208, new_n8209, new_n8210, new_n8211, new_n8212, new_n8213,
    new_n8214, new_n8215, new_n8216, new_n8217, new_n8218, new_n8219,
    new_n8220, new_n8221, new_n8222, new_n8223, new_n8224, new_n8225,
    new_n8226, new_n8227, new_n8228, new_n8229, new_n8230, new_n8231,
    new_n8232, new_n8233, new_n8234, new_n8235, new_n8236_1, new_n8237,
    new_n8238, new_n8239, new_n8240, new_n8241, new_n8242, new_n8243,
    new_n8244, new_n8245, new_n8246, new_n8247, new_n8248, new_n8249,
    new_n8250, new_n8251, new_n8252, new_n8253, new_n8254, new_n8255,
    new_n8256, new_n8257, new_n8258, new_n8259, new_n8260, new_n8261,
    new_n8262, new_n8263, new_n8264, new_n8265, new_n8266, new_n8267,
    new_n8268, new_n8269, new_n8270, new_n8271, new_n8272, new_n8273,
    new_n8274, new_n8275, new_n8276_1, new_n8277, new_n8278, new_n8279,
    new_n8280, new_n8281, new_n8282, new_n8283, new_n8284, new_n8285,
    new_n8286, new_n8287, new_n8288, new_n8289, new_n8290, new_n8291,
    new_n8292, new_n8293, new_n8294, new_n8295, new_n8296, new_n8297,
    new_n8298, new_n8299, new_n8300, new_n8301, new_n8302, new_n8303_1,
    new_n8304, new_n8305, new_n8306, new_n8307, new_n8308, new_n8309,
    new_n8310, new_n8311, new_n8312, new_n8313, new_n8314, new_n8315,
    new_n8316, new_n8317, new_n8318, new_n8319, new_n8320, new_n8321,
    new_n8322, new_n8323, new_n8324, new_n8325, new_n8326, new_n8327,
    new_n8328, new_n8329, new_n8330, new_n8331, new_n8332, new_n8333,
    new_n8334, new_n8335, new_n8336_1, new_n8337, new_n8338, new_n8339,
    new_n8340, new_n8341, new_n8342, new_n8343, new_n8344, new_n8345,
    new_n8346, new_n8347, new_n8348, new_n8349, new_n8350, new_n8351,
    new_n8352, new_n8353, new_n8354, new_n8355, new_n8356, new_n8357,
    new_n8358, new_n8359, new_n8360, new_n8361, new_n8362, new_n8363,
    new_n8364, new_n8365, new_n8366, new_n8367, new_n8368, new_n8369,
    new_n8370, new_n8371, new_n8372, new_n8373, new_n8374, new_n8375,
    new_n8376, new_n8377, new_n8378, new_n8379, new_n8380, new_n8381,
    new_n8382, new_n8383, new_n8384_1, new_n8385, new_n8386, new_n8387,
    new_n8388, new_n8389, new_n8390, new_n8391, new_n8392, new_n8393,
    new_n8394, new_n8395, new_n8396, new_n8397, new_n8398_1, new_n8399,
    new_n8400, new_n8401, new_n8402, new_n8403, new_n8404, new_n8405,
    new_n8406, new_n8407, new_n8408, new_n8409, new_n8410, new_n8411,
    new_n8412, new_n8414, new_n8415, new_n8416, new_n8418, new_n8419,
    new_n8420, new_n8422, new_n8423, new_n8424, new_n8426, new_n8427,
    new_n8428, new_n8430, new_n8431, new_n8432, new_n8434, new_n8435,
    new_n8436, new_n8437, new_n8438, new_n8439, new_n8440, new_n8441,
    new_n8442, new_n8443, new_n8444, new_n8445, new_n8446, new_n8447,
    new_n8448, new_n8449, new_n8450, new_n8451, new_n8452, new_n8453,
    new_n8454, new_n8455, new_n8456, new_n8457, new_n8458, new_n8459,
    new_n8460, new_n8461, new_n8462, new_n8463, new_n8464, new_n8465,
    new_n8466, new_n8467, new_n8468, new_n8469, new_n8470, new_n8471,
    new_n8472, new_n8473, new_n8474, new_n8475, new_n8476_1, new_n8477,
    new_n8478, new_n8479, new_n8480, new_n8481, new_n8482, new_n8483,
    new_n8484, new_n8485, new_n8486, new_n8487, new_n8488, new_n8489,
    new_n8490, new_n8491, new_n8492, new_n8493, new_n8494, new_n8495,
    new_n8496, new_n8497, new_n8498, new_n8499, new_n8500, new_n8501,
    new_n8502, new_n8503, new_n8504, new_n8505, new_n8506, new_n8507,
    new_n8508, new_n8509, new_n8510, new_n8511, new_n8512, new_n8513,
    new_n8514, new_n8515, new_n8516, new_n8517, new_n8518, new_n8519,
    new_n8520, new_n8521, new_n8522, new_n8523, new_n8524, new_n8525,
    new_n8526, new_n8527, new_n8528, new_n8529, new_n8530, new_n8531,
    new_n8532, new_n8533, new_n8534, new_n8535, new_n8536, new_n8537,
    new_n8538, new_n8539, new_n8540, new_n8541, new_n8542, new_n8543,
    new_n8544, new_n8545, new_n8546, new_n8547, new_n8548, new_n8549,
    new_n8550, new_n8551, new_n8552, new_n8553, new_n8554, new_n8555,
    new_n8556, new_n8557, new_n8558, new_n8559, new_n8560, new_n8561,
    new_n8562, new_n8563, new_n8564, new_n8565, new_n8566, new_n8567,
    new_n8568, new_n8569, new_n8570, new_n8571, new_n8572, new_n8573,
    new_n8574, new_n8575, new_n8576, new_n8577, new_n8578, new_n8579,
    new_n8580, new_n8581, new_n8582, new_n8583, new_n8584, new_n8585,
    new_n8586, new_n8587, new_n8588, new_n8589, new_n8590, new_n8591,
    new_n8592, new_n8593, new_n8594, new_n8595_1, new_n8596, new_n8597,
    new_n8598, new_n8599, new_n8600, new_n8601, new_n8602, new_n8603,
    new_n8604, new_n8605, new_n8606, new_n8607, new_n8608, new_n8609,
    new_n8610, new_n8611, new_n8612, new_n8613, new_n8614, new_n8615,
    new_n8616, new_n8617, new_n8618, new_n8619, new_n8620, new_n8621,
    new_n8622, new_n8623, new_n8624, new_n8625, new_n8626, new_n8627,
    new_n8628, new_n8629, new_n8630, new_n8631, new_n8632, new_n8633,
    new_n8634, new_n8635, new_n8636, new_n8637, new_n8638, new_n8639,
    new_n8640, new_n8641, new_n8642, new_n8643, new_n8644, new_n8645,
    new_n8646, new_n8647, new_n8648, new_n8649, new_n8650, new_n8651,
    new_n8652, new_n8653, new_n8654, new_n8655, new_n8656, new_n8657,
    new_n8658, new_n8659, new_n8660, new_n8661, new_n8662, new_n8663,
    new_n8664, new_n8665_1, new_n8666, new_n8667, new_n8668, new_n8669,
    new_n8670, new_n8671, new_n8672, new_n8673, new_n8674, new_n8675,
    new_n8676, new_n8677, new_n8678, new_n8679, new_n8680, new_n8681,
    new_n8682, new_n8683, new_n8684, new_n8685, new_n8686, new_n8687,
    new_n8688, new_n8689, new_n8690, new_n8691, new_n8692, new_n8693,
    new_n8694, new_n8695, new_n8696, new_n8697, new_n8698, new_n8699,
    new_n8700, new_n8701, new_n8702, new_n8703, new_n8704, new_n8705,
    new_n8706, new_n8707, new_n8708, new_n8709, new_n8710, new_n8711,
    new_n8712, new_n8713, new_n8714, new_n8715, new_n8716, new_n8717_1,
    new_n8718, new_n8719, new_n8720, new_n8721, new_n8722, new_n8723,
    new_n8724, new_n8725, new_n8726, new_n8727, new_n8728, new_n8729,
    new_n8730, new_n8731, new_n8732, new_n8733, new_n8734, new_n8735,
    new_n8736, new_n8737, new_n8738, new_n8739, new_n8740, new_n8741,
    new_n8742, new_n8743, new_n8744, new_n8745, new_n8746, new_n8747,
    new_n8748, new_n8749, new_n8750, new_n8751, new_n8752, new_n8753,
    new_n8754, new_n8755, new_n8756, new_n8757, new_n8758, new_n8759_1,
    new_n8760, new_n8761, new_n8762, new_n8763, new_n8764, new_n8765,
    new_n8766, new_n8767, new_n8768, new_n8769, new_n8770, new_n8771,
    new_n8772, new_n8773, new_n8774, new_n8775, new_n8776, new_n8777,
    new_n8778, new_n8779, new_n8780, new_n8781, new_n8782, new_n8783,
    new_n8784, new_n8785, new_n8786, new_n8787, new_n8788, new_n8789,
    new_n8790, new_n8791, new_n8792, new_n8793, new_n8794, new_n8795,
    new_n8796, new_n8797, new_n8798, new_n8799, new_n8800, new_n8801,
    new_n8802, new_n8803, new_n8804, new_n8805, new_n8806, new_n8807,
    new_n8808, new_n8809, new_n8810, new_n8811, new_n8812, new_n8813,
    new_n8814, new_n8815, new_n8816, new_n8817, new_n8818, new_n8819_1,
    new_n8820, new_n8821, new_n8822, new_n8823, new_n8824, new_n8825,
    new_n8826, new_n8827, new_n8828, new_n8829, new_n8830, new_n8831,
    new_n8832, new_n8833, new_n8834, new_n8835, new_n8836, new_n8837,
    new_n8838, new_n8839, new_n8840, new_n8841, new_n8842, new_n8843,
    new_n8844, new_n8845, new_n8846, new_n8847, new_n8848, new_n8849,
    new_n8850, new_n8851, new_n8852, new_n8853, new_n8854, new_n8855,
    new_n8856, new_n8857, new_n8858, new_n8859, new_n8860, new_n8861,
    new_n8862, new_n8863, new_n8864, new_n8865, new_n8866, new_n8867,
    new_n8868, new_n8869, new_n8870, new_n8871, new_n8872, new_n8873,
    new_n8874, new_n8875, new_n8876, new_n8877, new_n8878, new_n8879,
    new_n8880, new_n8881, new_n8882, new_n8883, new_n8884, new_n8885,
    new_n8886, new_n8887, new_n8888, new_n8889, new_n8890, new_n8891,
    new_n8892, new_n8893, new_n8894, new_n8895, new_n8896, new_n8897,
    new_n8898, new_n8899, new_n8900, new_n8901, new_n8902, new_n8903,
    new_n8904, new_n8905, new_n8906, new_n8907, new_n8908, new_n8909,
    new_n8910, new_n8911, new_n8912, new_n8913, new_n8914, new_n8915,
    new_n8916, new_n8917, new_n8918, new_n8919, new_n8920, new_n8921,
    new_n8922, new_n8923, new_n8924, new_n8925, new_n8926, new_n8927,
    new_n8928, new_n8929, new_n8930, new_n8931, new_n8932, new_n8933,
    new_n8934, new_n8935, new_n8936, new_n8937, new_n8938, new_n8939,
    new_n8940, new_n8941, new_n8942, new_n8943, new_n8944, new_n8945,
    new_n8946, new_n8947, new_n8948, new_n8949, new_n8950, new_n8951,
    new_n8952, new_n8953, new_n8954, new_n8955, new_n8956, new_n8957,
    new_n8958, new_n8959, new_n8960, new_n8961, new_n8962, new_n8963,
    new_n8964, new_n8965, new_n8966, new_n8967, new_n8968, new_n8969,
    new_n8970, new_n8971, new_n8972, new_n8973, new_n8974, new_n8975,
    new_n8976, new_n8977, new_n8978, new_n8979, new_n8980, new_n8981,
    new_n8982, new_n8983, new_n8984, new_n8985, new_n8986, new_n8987,
    new_n8988, new_n8989, new_n8990, new_n8991, new_n8992, new_n8993,
    new_n8994, new_n8995, new_n8996, new_n8997, new_n8998, new_n8999,
    new_n9000, new_n9001, new_n9002, new_n9003, new_n9004, new_n9005,
    new_n9006, new_n9007, new_n9008, new_n9009, new_n9010, new_n9011,
    new_n9012, new_n9013, new_n9014, new_n9015, new_n9016, new_n9017,
    new_n9018, new_n9019, new_n9020, new_n9021, new_n9022, new_n9023,
    new_n9024, new_n9025, new_n9026, new_n9027, new_n9028, new_n9029,
    new_n9030, new_n9031, new_n9032, new_n9033, new_n9034, new_n9035,
    new_n9036, new_n9037, new_n9038, new_n9039, new_n9040, new_n9041,
    new_n9042, new_n9043, new_n9044, new_n9045, new_n9046, new_n9047,
    new_n9048, new_n9049, new_n9050, new_n9051, new_n9052, new_n9053,
    new_n9054, new_n9055, new_n9056, new_n9057, new_n9058, new_n9059,
    new_n9060, new_n9061, new_n9062, new_n9063, new_n9064, new_n9065,
    new_n9066, new_n9067, new_n9068, new_n9069, new_n9070, new_n9071,
    new_n9072, new_n9073, new_n9074, new_n9076, new_n9077, new_n9078,
    new_n9079, new_n9080_1, new_n9081, new_n9082, new_n9083, new_n9084,
    new_n9085, new_n9086, new_n9087, new_n9088, new_n9089, new_n9090,
    new_n9091, new_n9092, new_n9093, new_n9094, new_n9095, new_n9096,
    new_n9097, new_n9098, new_n9099, new_n9100, new_n9101, new_n9102,
    new_n9103, new_n9104, new_n9105, new_n9106, new_n9107, new_n9108,
    new_n9109, new_n9110, new_n9111_1, new_n9112, new_n9113, new_n9114,
    new_n9115, new_n9116, new_n9117, new_n9118, new_n9119, new_n9120,
    new_n9121, new_n9122, new_n9123, new_n9124, new_n9125, new_n9126,
    new_n9127, new_n9128, new_n9129, new_n9130, new_n9131, new_n9132,
    new_n9133, new_n9134, new_n9135, new_n9136, new_n9137_1, new_n9138,
    new_n9139, new_n9140, new_n9141, new_n9142, new_n9143, new_n9144,
    new_n9145, new_n9146, new_n9147, new_n9148, new_n9149, new_n9150,
    new_n9151, new_n9152, new_n9153, new_n9154, new_n9155, new_n9156,
    new_n9157, new_n9158, new_n9159, new_n9160, new_n9161, new_n9162,
    new_n9163, new_n9164, new_n9165, new_n9166, new_n9167, new_n9168,
    new_n9169, new_n9170, new_n9171, new_n9172, new_n9173, new_n9174,
    new_n9175, new_n9176, new_n9177, new_n9178, new_n9179, new_n9180,
    new_n9181, new_n9182, new_n9183, new_n9184, new_n9185, new_n9186,
    new_n9187, new_n9188, new_n9189_1, new_n9190, new_n9191, new_n9192,
    new_n9193, new_n9194, new_n9195_1, new_n9196, new_n9197, new_n9198,
    new_n9199, new_n9200, new_n9201, new_n9202, new_n9203, new_n9204,
    new_n9205, new_n9206, new_n9207, new_n9208, new_n9209, new_n9210,
    new_n9211, new_n9212, new_n9213, new_n9214, new_n9215, new_n9216,
    new_n9217, new_n9218, new_n9219, new_n9220, new_n9221, new_n9222,
    new_n9223, new_n9224, new_n9225, new_n9226, new_n9227, new_n9228,
    new_n9229, new_n9230, new_n9231, new_n9232, new_n9233, new_n9234,
    new_n9235, new_n9236, new_n9237, new_n9238, new_n9239, new_n9240,
    new_n9241_1, new_n9242, new_n9243, new_n9244, new_n9245, new_n9246,
    new_n9247, new_n9248, new_n9249, new_n9250, new_n9251, new_n9252,
    new_n9253, new_n9254, new_n9256, new_n9257, new_n9258, new_n9260,
    new_n9261, new_n9262, new_n9264, new_n9265, new_n9266, new_n9267,
    new_n9268, new_n9269, new_n9270, new_n9271, new_n9272, new_n9273,
    new_n9274, new_n9275, new_n9277, new_n9278, new_n9279, new_n9281,
    new_n9282, new_n9283, new_n9284, new_n9285, new_n9286, new_n9287,
    new_n9288, new_n9289, new_n9290, new_n9291, new_n9292, new_n9293,
    new_n9294, new_n9295, new_n9296, new_n9297, new_n9298, new_n9299,
    new_n9300, new_n9301, new_n9302, new_n9303, new_n9304, new_n9305,
    new_n9306, new_n9307, new_n9308, new_n9309, new_n9310, new_n9311,
    new_n9312, new_n9313, new_n9314, new_n9315, new_n9316, new_n9317,
    new_n9318, new_n9319, new_n9320, new_n9321, new_n9322, new_n9323,
    new_n9324, new_n9325, new_n9326, new_n9327, new_n9328, new_n9329,
    new_n9330, new_n9331, new_n9332, new_n9333, new_n9334, new_n9335,
    new_n9336, new_n9337, new_n9338, new_n9339, new_n9340, new_n9341,
    new_n9342, new_n9343, new_n9344, new_n9345, new_n9346, new_n9347,
    new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353,
    new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359,
    new_n9360, new_n9361, new_n9362, new_n9363, new_n9364, new_n9365,
    new_n9366, new_n9367, new_n9368, new_n9369, new_n9370, new_n9371,
    new_n9372, new_n9373, new_n9374, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380, new_n9381, new_n9382, new_n9383,
    new_n9384, new_n9386, new_n9387_1, new_n9388, new_n9390, new_n9391,
    new_n9392, new_n9394, new_n9395, new_n9396, new_n9397, new_n9398,
    new_n9399, new_n9400_1, new_n9401, new_n9402, new_n9403, new_n9404,
    new_n9405, new_n9406, new_n9407, new_n9408, new_n9409, new_n9410,
    new_n9411, new_n9412, new_n9413, new_n9414, new_n9415, new_n9416,
    new_n9417, new_n9418, new_n9419, new_n9420, new_n9421, new_n9422,
    new_n9423, new_n9424, new_n9425, new_n9426, new_n9427, new_n9428,
    new_n9429, new_n9430, new_n9431, new_n9432, new_n9433, new_n9434,
    new_n9435, new_n9436, new_n9437, new_n9438, new_n9439, new_n9440,
    new_n9441, new_n9442, new_n9443, new_n9444, new_n9445, new_n9446,
    new_n9447, new_n9448, new_n9449, new_n9450, new_n9451, new_n9452,
    new_n9453, new_n9454, new_n9455, new_n9456, new_n9457_1, new_n9458,
    new_n9459, new_n9460, new_n9461, new_n9462, new_n9463, new_n9464,
    new_n9465, new_n9466, new_n9467, new_n9468, new_n9469, new_n9470,
    new_n9471, new_n9472, new_n9473, new_n9474, new_n9475, new_n9476,
    new_n9477, new_n9478, new_n9479, new_n9480, new_n9481, new_n9482,
    new_n9483, new_n9484, new_n9485, new_n9486, new_n9487, new_n9488,
    new_n9489, new_n9490, new_n9491, new_n9492, new_n9493, new_n9494,
    new_n9495, new_n9496, new_n9497, new_n9498, new_n9499, new_n9500,
    new_n9501, new_n9502, new_n9503, new_n9504, new_n9505, new_n9506,
    new_n9507, new_n9508, new_n9509, new_n9510, new_n9511, new_n9512,
    new_n9513, new_n9514, new_n9515, new_n9516, new_n9517, new_n9518,
    new_n9519, new_n9520, new_n9521, new_n9522, new_n9523, new_n9524,
    new_n9525, new_n9526, new_n9527, new_n9528, new_n9529, new_n9530,
    new_n9531, new_n9532, new_n9533, new_n9534, new_n9535, new_n9536,
    new_n9537, new_n9538, new_n9539, new_n9540, new_n9541, new_n9542,
    new_n9543, new_n9544, new_n9545, new_n9546, new_n9547, new_n9548,
    new_n9549, new_n9550, new_n9551, new_n9552, new_n9553, new_n9554,
    new_n9555, new_n9556, new_n9557, new_n9558, new_n9559, new_n9560,
    new_n9561, new_n9562, new_n9563, new_n9564, new_n9565, new_n9566,
    new_n9567, new_n9568, new_n9569, new_n9570, new_n9571_1, new_n9572,
    new_n9573, new_n9574, new_n9575, new_n9576, new_n9577, new_n9578_1,
    new_n9579, new_n9580, new_n9581, new_n9582, new_n9583_1, new_n9584,
    new_n9585, new_n9586, new_n9587, new_n9588, new_n9589, new_n9590,
    new_n9591, new_n9592, new_n9593, new_n9594, new_n9595, new_n9596,
    new_n9597, new_n9598, new_n9599, new_n9600, new_n9601, new_n9602,
    new_n9603, new_n9604, new_n9605, new_n9606, new_n9607, new_n9608,
    new_n9609, new_n9610, new_n9611, new_n9612, new_n9613, new_n9614,
    new_n9615, new_n9616, new_n9617, new_n9618, new_n9619, new_n9620,
    new_n9621, new_n9622, new_n9623, new_n9624, new_n9625, new_n9626,
    new_n9627, new_n9628, new_n9629, new_n9630, new_n9631, new_n9632,
    new_n9633, new_n9634, new_n9635, new_n9636, new_n9637_1, new_n9638,
    new_n9639, new_n9640_1, new_n9641, new_n9642, new_n9643, new_n9644,
    new_n9645, new_n9646, new_n9647, new_n9648, new_n9649, new_n9650,
    new_n9651, new_n9652, new_n9653, new_n9654, new_n9655, new_n9656,
    new_n9657, new_n9658, new_n9659, new_n9660, new_n9661, new_n9662,
    new_n9663, new_n9664, new_n9665, new_n9666, new_n9667, new_n9668,
    new_n9669, new_n9670, new_n9671, new_n9672, new_n9673, new_n9674,
    new_n9675, new_n9676, new_n9677, new_n9678, new_n9679, new_n9680,
    new_n9681, new_n9682, new_n9683, new_n9684, new_n9685, new_n9686,
    new_n9687, new_n9688, new_n9689, new_n9690, new_n9691, new_n9692,
    new_n9693, new_n9694, new_n9695, new_n9696, new_n9697, new_n9698,
    new_n9699, new_n9700, new_n9701, new_n9702, new_n9703, new_n9704,
    new_n9705, new_n9706_1, new_n9707, new_n9708, new_n9709, new_n9710,
    new_n9711, new_n9712, new_n9713, new_n9714, new_n9715, new_n9716,
    new_n9717, new_n9718, new_n9719, new_n9720, new_n9721, new_n9722,
    new_n9723, new_n9724, new_n9725_1, new_n9726, new_n9727, new_n9728,
    new_n9729, new_n9730, new_n9731, new_n9732, new_n9733, new_n9734,
    new_n9735, new_n9736, new_n9737, new_n9738, new_n9739, new_n9740,
    new_n9741, new_n9742, new_n9743, new_n9744, new_n9745, new_n9746,
    new_n9747, new_n9748, new_n9749, new_n9750, new_n9751, new_n9752,
    new_n9753, new_n9754, new_n9755, new_n9756_1, new_n9757, new_n9758,
    new_n9759, new_n9760, new_n9761, new_n9762, new_n9763_1, new_n9764,
    new_n9765, new_n9766, new_n9767_1, new_n9768, new_n9769, new_n9770,
    new_n9771, new_n9772, new_n9773, new_n9774, new_n9775, new_n9776,
    new_n9777, new_n9778, new_n9779, new_n9780, new_n9781, new_n9782,
    new_n9783, new_n9784, new_n9785, new_n9786, new_n9787, new_n9788,
    new_n9789, new_n9790, new_n9791, new_n9792, new_n9793, new_n9794,
    new_n9795, new_n9796, new_n9797, new_n9798, new_n9799, new_n9800,
    new_n9801, new_n9802, new_n9803, new_n9804, new_n9805, new_n9806,
    new_n9807, new_n9808, new_n9809, new_n9810, new_n9811, new_n9812,
    new_n9813, new_n9814, new_n9815, new_n9816, new_n9817, new_n9818,
    new_n9819, new_n9820_1, new_n9821, new_n9822, new_n9823, new_n9824,
    new_n9825, new_n9826, new_n9827, new_n9828, new_n9829, new_n9830,
    new_n9831, new_n9832, new_n9833, new_n9834, new_n9835, new_n9836,
    new_n9837, new_n9838, new_n9839, new_n9840, new_n9841, new_n9842,
    new_n9843, new_n9844, new_n9845, new_n9846, new_n9847, new_n9848,
    new_n9849, new_n9850, new_n9851, new_n9852, new_n9853, new_n9854,
    new_n9855, new_n9856, new_n9857, new_n9858, new_n9859, new_n9860,
    new_n9861, new_n9862, new_n9863, new_n9864, new_n9865, new_n9866,
    new_n9867, new_n9868, new_n9869, new_n9870, new_n9871, new_n9872,
    new_n9873, new_n9874, new_n9875, new_n9876, new_n9877, new_n9878,
    new_n9879, new_n9880, new_n9881, new_n9882, new_n9883, new_n9884,
    new_n9885, new_n9886, new_n9887, new_n9888, new_n9889, new_n9890,
    new_n9891, new_n9892, new_n9893, new_n9894, new_n9895, new_n9896,
    new_n9897, new_n9898, new_n9899, new_n9900, new_n9901, new_n9902,
    new_n9903, new_n9904, new_n9905, new_n9906, new_n9907, new_n9908,
    new_n9909, new_n9910, new_n9911, new_n9912, new_n9913, new_n9914,
    new_n9915, new_n9916, new_n9917, new_n9918, new_n9919, new_n9920_1,
    new_n9921, new_n9922, new_n9923, new_n9924, new_n9925, new_n9926,
    new_n9927, new_n9928, new_n9929, new_n9930, new_n9931, new_n9932,
    new_n9933, new_n9934, new_n9935, new_n9936, new_n9937, new_n9938_1,
    new_n9939, new_n9940, new_n9941, new_n9942, new_n9943, new_n9944,
    new_n9945, new_n9946, new_n9947, new_n9948, new_n9949, new_n9950,
    new_n9951, new_n9952, new_n9953, new_n9954, new_n9955, new_n9956_1,
    new_n9957, new_n9958, new_n9959, new_n9960, new_n9961, new_n9962,
    new_n9963, new_n9964, new_n9965, new_n9966, new_n9967, new_n9968,
    new_n9969, new_n9970, new_n9971, new_n9972, new_n9973, new_n9974,
    new_n9975, new_n9976, new_n9977, new_n9978, new_n9979, new_n9980,
    new_n9981, new_n9982, new_n9983, new_n9984, new_n9985, new_n9986,
    new_n9987, new_n9988, new_n9989, new_n9990, new_n9991, new_n9992,
    new_n9993, new_n9994, new_n9995, new_n9996, new_n9997, new_n9998,
    new_n9999, new_n10000, new_n10001, new_n10002, new_n10003, new_n10004,
    new_n10005, new_n10006, new_n10007, new_n10008, new_n10009, new_n10010,
    new_n10011, new_n10012, new_n10013, new_n10014, new_n10015, new_n10016,
    new_n10017, new_n10018, new_n10019, new_n10020, new_n10021,
    new_n10022_1, new_n10023, new_n10024, new_n10025, new_n10026,
    new_n10027, new_n10028, new_n10029, new_n10030, new_n10031, new_n10032,
    new_n10033, new_n10034, new_n10035, new_n10036, new_n10037, new_n10038,
    new_n10039, new_n10040, new_n10041, new_n10042, new_n10043, new_n10044,
    new_n10045, new_n10046, new_n10047, new_n10048, new_n10049, new_n10050,
    new_n10051, new_n10052, new_n10053, new_n10054, new_n10055, new_n10056,
    new_n10057, new_n10058, new_n10059, new_n10060, new_n10061, new_n10062,
    new_n10063, new_n10064, new_n10065, new_n10066, new_n10067, new_n10068,
    new_n10069, new_n10070, new_n10071, new_n10072, new_n10073, new_n10074,
    new_n10075, new_n10076, new_n10077, new_n10078, new_n10079, new_n10080,
    new_n10081, new_n10082, new_n10083, new_n10084, new_n10085, new_n10086,
    new_n10087, new_n10088, new_n10089, new_n10090, new_n10091, new_n10092,
    new_n10093, new_n10094, new_n10095, new_n10096, new_n10097, new_n10098,
    new_n10099, new_n10100, new_n10101, new_n10102, new_n10103, new_n10104,
    new_n10105, new_n10106, new_n10107, new_n10108, new_n10109, new_n10110,
    new_n10111, new_n10112, new_n10113, new_n10114, new_n10115, new_n10116,
    new_n10117, new_n10118, new_n10119, new_n10120, new_n10121, new_n10122,
    new_n10123, new_n10124, new_n10125, new_n10126, new_n10127, new_n10128,
    new_n10129, new_n10130, new_n10131, new_n10132, new_n10133, new_n10134,
    new_n10135, new_n10136, new_n10137, new_n10138, new_n10139, new_n10140,
    new_n10141, new_n10142, new_n10143, new_n10144, new_n10145, new_n10146,
    new_n10147, new_n10148, new_n10149, new_n10150, new_n10151, new_n10152,
    new_n10153, new_n10154, new_n10155, new_n10156, new_n10157, new_n10158,
    new_n10159, new_n10160, new_n10161, new_n10162, new_n10163, new_n10164,
    new_n10165, new_n10166, new_n10167, new_n10168, new_n10169, new_n10170,
    new_n10171, new_n10172, new_n10173, new_n10174_1, new_n10175,
    new_n10176, new_n10177, new_n10178, new_n10179, new_n10180, new_n10181,
    new_n10182, new_n10183, new_n10184, new_n10185, new_n10186, new_n10187,
    new_n10188, new_n10189, new_n10190, new_n10191, new_n10192, new_n10193,
    new_n10194, new_n10195, new_n10196, new_n10197, new_n10198, new_n10199,
    new_n10200, new_n10201, new_n10202, new_n10203, new_n10204, new_n10205,
    new_n10206, new_n10207, new_n10208, new_n10209, new_n10210, new_n10211,
    new_n10212, new_n10213, new_n10214, new_n10215, new_n10216,
    new_n10217_1, new_n10218, new_n10219, new_n10220, new_n10221,
    new_n10222, new_n10223_1, new_n10224, new_n10225, new_n10226,
    new_n10227, new_n10228, new_n10229, new_n10230, new_n10231, new_n10232,
    new_n10233, new_n10234, new_n10235, new_n10236, new_n10237, new_n10238,
    new_n10239, new_n10240, new_n10241, new_n10242, new_n10243, new_n10244,
    new_n10245, new_n10246, new_n10247, new_n10248, new_n10249, new_n10250,
    new_n10251, new_n10252, new_n10253, new_n10254, new_n10255, new_n10256,
    new_n10257, new_n10258, new_n10259, new_n10260, new_n10261, new_n10262,
    new_n10263, new_n10264, new_n10265, new_n10266, new_n10267, new_n10268,
    new_n10269, new_n10270, new_n10271, new_n10272, new_n10273, new_n10274,
    new_n10275, new_n10276, new_n10277, new_n10278_1, new_n10280,
    new_n10281, new_n10282, new_n10284, new_n10285, new_n10286, new_n10288,
    new_n10289, new_n10290, new_n10291, new_n10292, new_n10293, new_n10294,
    new_n10295, new_n10296, new_n10297, new_n10298, new_n10299, new_n10300,
    new_n10301, new_n10302, new_n10303, new_n10304, new_n10305, new_n10306,
    new_n10307, new_n10308, new_n10309, new_n10310, new_n10311, new_n10312,
    new_n10313, new_n10314, new_n10315, new_n10316, new_n10317, new_n10318,
    new_n10319, new_n10320, new_n10321, new_n10322, new_n10323, new_n10324,
    new_n10325, new_n10326, new_n10327_1, new_n10328, new_n10329,
    new_n10330, new_n10331, new_n10332, new_n10333, new_n10334, new_n10335,
    new_n10336, new_n10337, new_n10338, new_n10339, new_n10340, new_n10341,
    new_n10342, new_n10343, new_n10344, new_n10345, new_n10346, new_n10347,
    new_n10348, new_n10349, new_n10350, new_n10351, new_n10352, new_n10353,
    new_n10354, new_n10355, new_n10356, new_n10357, new_n10358, new_n10359,
    new_n10360, new_n10361, new_n10362, new_n10363, new_n10364, new_n10365,
    new_n10366, new_n10367, new_n10368, new_n10369, new_n10370, new_n10371,
    new_n10372, new_n10373, new_n10374, new_n10375, new_n10376, new_n10377,
    new_n10378, new_n10379, new_n10380, new_n10381, new_n10382, new_n10383,
    new_n10384, new_n10385, new_n10386, new_n10387, new_n10388, new_n10389,
    new_n10390, new_n10391_1, new_n10392, new_n10393, new_n10394,
    new_n10395, new_n10396, new_n10397, new_n10398, new_n10399, new_n10400,
    new_n10401, new_n10402, new_n10403, new_n10404, new_n10405, new_n10406,
    new_n10407, new_n10408, new_n10409, new_n10410, new_n10411, new_n10412,
    new_n10413, new_n10414, new_n10415, new_n10416, new_n10417, new_n10418,
    new_n10419, new_n10420, new_n10421, new_n10422, new_n10423, new_n10424,
    new_n10425, new_n10426, new_n10427, new_n10428, new_n10429, new_n10430,
    new_n10431, new_n10432, new_n10433, new_n10434, new_n10435, new_n10436,
    new_n10437, new_n10438, new_n10439_1, new_n10440, new_n10441,
    new_n10442, new_n10443, new_n10444, new_n10445, new_n10446, new_n10447,
    new_n10448, new_n10449, new_n10450, new_n10451_1, new_n10452,
    new_n10453, new_n10454, new_n10455, new_n10456, new_n10457, new_n10458,
    new_n10459, new_n10460, new_n10461, new_n10462, new_n10463, new_n10464,
    new_n10465, new_n10466, new_n10467, new_n10468, new_n10469, new_n10470,
    new_n10471, new_n10472, new_n10473, new_n10474, new_n10475,
    new_n10476_1, new_n10477, new_n10478, new_n10479, new_n10480,
    new_n10481, new_n10482, new_n10483, new_n10484, new_n10485, new_n10486,
    new_n10487, new_n10488, new_n10489, new_n10490, new_n10491, new_n10492,
    new_n10493, new_n10494, new_n10495, new_n10496, new_n10497, new_n10498,
    new_n10499, new_n10500, new_n10501, new_n10502, new_n10503, new_n10504,
    new_n10505, new_n10506, new_n10507, new_n10508, new_n10509,
    new_n10510_1, new_n10511, new_n10512, new_n10513, new_n10514,
    new_n10515, new_n10516, new_n10517, new_n10518, new_n10519, new_n10520,
    new_n10521, new_n10522, new_n10523, new_n10524, new_n10525, new_n10526,
    new_n10527, new_n10528, new_n10529, new_n10530, new_n10531, new_n10532,
    new_n10533, new_n10534, new_n10535, new_n10536, new_n10537, new_n10538,
    new_n10539, new_n10540, new_n10541, new_n10542, new_n10543, new_n10544,
    new_n10545_1, new_n10546, new_n10547_1, new_n10548, new_n10549,
    new_n10550, new_n10551, new_n10552, new_n10553, new_n10554, new_n10555,
    new_n10556, new_n10557, new_n10558, new_n10559, new_n10560, new_n10561,
    new_n10562, new_n10563, new_n10564, new_n10565, new_n10566, new_n10567,
    new_n10568, new_n10569, new_n10570, new_n10571, new_n10572, new_n10573,
    new_n10574, new_n10575, new_n10576, new_n10577, new_n10578, new_n10579,
    new_n10580, new_n10581, new_n10582, new_n10583, new_n10584, new_n10585,
    new_n10586, new_n10587, new_n10588, new_n10589_1, new_n10590,
    new_n10591, new_n10592, new_n10593, new_n10594, new_n10595, new_n10596,
    new_n10597, new_n10598, new_n10599, new_n10600, new_n10601, new_n10602,
    new_n10603, new_n10604, new_n10605, new_n10606, new_n10607, new_n10608,
    new_n10609, new_n10610, new_n10611, new_n10612, new_n10613, new_n10614,
    new_n10615, new_n10616, new_n10617, new_n10618, new_n10619, new_n10620,
    new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626,
    new_n10627, new_n10628, new_n10629, new_n10630, new_n10631, new_n10632,
    new_n10633, new_n10634, new_n10635, new_n10636, new_n10637, new_n10638,
    new_n10639, new_n10640, new_n10641, new_n10642, new_n10643,
    new_n10644_1, new_n10645, new_n10646, new_n10647, new_n10648,
    new_n10649, new_n10650, new_n10651, new_n10652, new_n10653, new_n10654,
    new_n10655, new_n10656, new_n10657, new_n10658, new_n10659, new_n10660,
    new_n10661, new_n10662, new_n10663, new_n10664, new_n10665, new_n10666,
    new_n10667, new_n10668, new_n10669, new_n10670, new_n10671, new_n10672,
    new_n10673, new_n10674, new_n10675, new_n10676, new_n10677,
    new_n10678_1, new_n10679, new_n10680, new_n10681, new_n10682,
    new_n10683, new_n10684, new_n10685_1, new_n10686, new_n10687,
    new_n10688, new_n10689, new_n10690, new_n10691, new_n10692, new_n10693,
    new_n10694, new_n10695_1, new_n10696, new_n10697, new_n10698,
    new_n10699, new_n10700, new_n10701, new_n10702, new_n10703, new_n10704,
    new_n10705, new_n10706, new_n10707, new_n10708, new_n10709, new_n10710,
    new_n10711, new_n10712, new_n10713, new_n10714, new_n10715, new_n10716,
    new_n10717, new_n10718, new_n10719, new_n10720, new_n10721, new_n10722,
    new_n10723, new_n10724, new_n10725, new_n10726, new_n10727, new_n10728,
    new_n10729, new_n10730, new_n10731, new_n10732, new_n10733, new_n10734,
    new_n10735, new_n10736, new_n10737, new_n10738, new_n10739, new_n10740,
    new_n10741, new_n10742, new_n10743, new_n10744, new_n10745, new_n10746,
    new_n10747, new_n10748, new_n10749, new_n10750, new_n10751, new_n10752,
    new_n10753, new_n10754, new_n10755, new_n10756, new_n10757, new_n10758,
    new_n10759, new_n10760, new_n10761, new_n10762, new_n10763, new_n10764,
    new_n10765, new_n10766, new_n10767, new_n10768, new_n10769, new_n10770,
    new_n10771, new_n10772, new_n10773, new_n10774, new_n10775, new_n10776,
    new_n10777, new_n10778, new_n10779, new_n10780, new_n10781, new_n10782,
    new_n10783, new_n10784, new_n10785, new_n10786, new_n10787, new_n10788,
    new_n10789_1, new_n10790, new_n10791, new_n10792, new_n10793,
    new_n10794, new_n10795, new_n10796, new_n10797, new_n10798, new_n10799,
    new_n10800, new_n10801, new_n10802, new_n10803, new_n10804, new_n10805,
    new_n10806, new_n10807, new_n10808, new_n10809, new_n10810, new_n10811,
    new_n10812, new_n10813, new_n10814, new_n10815, new_n10816, new_n10817,
    new_n10818, new_n10819, new_n10820, new_n10821, new_n10822, new_n10823,
    new_n10824, new_n10825, new_n10826, new_n10827, new_n10828, new_n10829,
    new_n10830, new_n10831, new_n10832, new_n10833, new_n10834, new_n10835,
    new_n10836, new_n10837, new_n10838, new_n10839, new_n10840, new_n10841,
    new_n10842, new_n10843, new_n10844, new_n10845, new_n10846, new_n10847,
    new_n10848_1, new_n10849, new_n10850, new_n10851_1, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864,
    new_n10865, new_n10866, new_n10867, new_n10868, new_n10869, new_n10870,
    new_n10871, new_n10872, new_n10873, new_n10874, new_n10875, new_n10876,
    new_n10877, new_n10878, new_n10879, new_n10880, new_n10881, new_n10882,
    new_n10883, new_n10884, new_n10885, new_n10886, new_n10887, new_n10888,
    new_n10889, new_n10890, new_n10891, new_n10892, new_n10893, new_n10894,
    new_n10895, new_n10896, new_n10897, new_n10898_1, new_n10899,
    new_n10900, new_n10901, new_n10902, new_n10903, new_n10904, new_n10905,
    new_n10906, new_n10907, new_n10908, new_n10909, new_n10910, new_n10911,
    new_n10912, new_n10913_1, new_n10914, new_n10915, new_n10916,
    new_n10917, new_n10918, new_n10919, new_n10920, new_n10921, new_n10922,
    new_n10923, new_n10924, new_n10925, new_n10926, new_n10927,
    new_n10928_1, new_n10929, new_n10930, new_n10931, new_n10932,
    new_n10933, new_n10934, new_n10935, new_n10936, new_n10937, new_n10938,
    new_n10939, new_n10940, new_n10941, new_n10942, new_n10943, new_n10944,
    new_n10945, new_n10946, new_n10947, new_n10948, new_n10949_1,
    new_n10950, new_n10951, new_n10952, new_n10953, new_n10954, new_n10955,
    new_n10956, new_n10957, new_n10958, new_n10959, new_n10960, new_n10961,
    new_n10962, new_n10963, new_n10964, new_n10965_1, new_n10966,
    new_n10967, new_n10968, new_n10969, new_n10970, new_n10971, new_n10972,
    new_n10973, new_n10974, new_n10975, new_n10976, new_n10977, new_n10978,
    new_n10979, new_n10980, new_n10981, new_n10982, new_n10983, new_n10984,
    new_n10985, new_n10986, new_n10987, new_n10988, new_n10989,
    new_n10990_1, new_n10991, new_n10992, new_n10993, new_n10994,
    new_n10995, new_n10996, new_n10997, new_n10998, new_n10999, new_n11000,
    new_n11001, new_n11002, new_n11003, new_n11004, new_n11005, new_n11006,
    new_n11007, new_n11008, new_n11009, new_n11010, new_n11011, new_n11012,
    new_n11013, new_n11014, new_n11015, new_n11016, new_n11017, new_n11018,
    new_n11019, new_n11020, new_n11021, new_n11022, new_n11023_1,
    new_n11024, new_n11025, new_n11026, new_n11027, new_n11028, new_n11029,
    new_n11030, new_n11031, new_n11032, new_n11033, new_n11034, new_n11035,
    new_n11036, new_n11037, new_n11038, new_n11039, new_n11040, new_n11041,
    new_n11042, new_n11043, new_n11044, new_n11045, new_n11046, new_n11047,
    new_n11048, new_n11049, new_n11050, new_n11051, new_n11052, new_n11053,
    new_n11054, new_n11055, new_n11056, new_n11057, new_n11058, new_n11059,
    new_n11060, new_n11061, new_n11062, new_n11063, new_n11064, new_n11065,
    new_n11066, new_n11067, new_n11068, new_n11069, new_n11070, new_n11071,
    new_n11072, new_n11073, new_n11074, new_n11075, new_n11076, new_n11077,
    new_n11078, new_n11079, new_n11080, new_n11081, new_n11082, new_n11083,
    new_n11084, new_n11085, new_n11086, new_n11087, new_n11088, new_n11089,
    new_n11090, new_n11091, new_n11092, new_n11093, new_n11094, new_n11095,
    new_n11096, new_n11097, new_n11098, new_n11099, new_n11100, new_n11101,
    new_n11102, new_n11103, new_n11104, new_n11105, new_n11106, new_n11107,
    new_n11108, new_n11109, new_n11110, new_n11111, new_n11112, new_n11113,
    new_n11114, new_n11115, new_n11116, new_n11117, new_n11118, new_n11119,
    new_n11120, new_n11121, new_n11122, new_n11123, new_n11124, new_n11125,
    new_n11126, new_n11127, new_n11128, new_n11129, new_n11130, new_n11131,
    new_n11132, new_n11133, new_n11134, new_n11135, new_n11136, new_n11137,
    new_n11138, new_n11139, new_n11140, new_n11141, new_n11142, new_n11143,
    new_n11144, new_n11145, new_n11146, new_n11147, new_n11148, new_n11149,
    new_n11150, new_n11151, new_n11152, new_n11153_1, new_n11154,
    new_n11155, new_n11156, new_n11157, new_n11158, new_n11159, new_n11160,
    new_n11161, new_n11162, new_n11163, new_n11164, new_n11165, new_n11166,
    new_n11167, new_n11168, new_n11169, new_n11170, new_n11171, new_n11172,
    new_n11173, new_n11174, new_n11175, new_n11176, new_n11177, new_n11178,
    new_n11179, new_n11180, new_n11181, new_n11182, new_n11183, new_n11184,
    new_n11185, new_n11186, new_n11187, new_n11188, new_n11189, new_n11190,
    new_n11191, new_n11192, new_n11193, new_n11194, new_n11195, new_n11196,
    new_n11197, new_n11198, new_n11199, new_n11200, new_n11201, new_n11202,
    new_n11203, new_n11204, new_n11205, new_n11206, new_n11207, new_n11208,
    new_n11209, new_n11210, new_n11211, new_n11212, new_n11213, new_n11214,
    new_n11215, new_n11216_1, new_n11217, new_n11218, new_n11219,
    new_n11220, new_n11221, new_n11222_1, new_n11223, new_n11224,
    new_n11225, new_n11226, new_n11227, new_n11228, new_n11229, new_n11230,
    new_n11231, new_n11232, new_n11233, new_n11234, new_n11235, new_n11236,
    new_n11237, new_n11238, new_n11239, new_n11240, new_n11241, new_n11242,
    new_n11243, new_n11244, new_n11245, new_n11246, new_n11247, new_n11248,
    new_n11249, new_n11250, new_n11251, new_n11252, new_n11253, new_n11254,
    new_n11255, new_n11256, new_n11257_1, new_n11258, new_n11259,
    new_n11260, new_n11261, new_n11262, new_n11263, new_n11264, new_n11265,
    new_n11266, new_n11267, new_n11268, new_n11269, new_n11270, new_n11271,
    new_n11272, new_n11273, new_n11274, new_n11276, new_n11277, new_n11278,
    new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285,
    new_n11286, new_n11287, new_n11288, new_n11289, new_n11290, new_n11291,
    new_n11292, new_n11293, new_n11294, new_n11295, new_n11296_1,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301, new_n11302,
    new_n11303, new_n11304, new_n11305, new_n11306, new_n11307, new_n11308,
    new_n11309, new_n11310, new_n11311_1, new_n11312, new_n11313,
    new_n11314, new_n11315, new_n11316, new_n11317, new_n11318, new_n11319,
    new_n11320, new_n11321, new_n11322, new_n11323, new_n11324, new_n11325,
    new_n11326_1, new_n11327, new_n11328, new_n11329, new_n11330,
    new_n11331, new_n11332, new_n11333, new_n11334, new_n11335, new_n11336,
    new_n11337, new_n11338, new_n11339, new_n11340, new_n11341, new_n11342,
    new_n11343, new_n11344, new_n11345, new_n11346, new_n11347, new_n11348,
    new_n11349, new_n11350, new_n11351, new_n11352, new_n11353, new_n11354,
    new_n11355, new_n11356, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375, new_n11376, new_n11377, new_n11378,
    new_n11379, new_n11380, new_n11381, new_n11382, new_n11383, new_n11384,
    new_n11385, new_n11386, new_n11387, new_n11388, new_n11389, new_n11390,
    new_n11391, new_n11392, new_n11393, new_n11394, new_n11395, new_n11396,
    new_n11397, new_n11398, new_n11399, new_n11400, new_n11401, new_n11402,
    new_n11403, new_n11404, new_n11405, new_n11406, new_n11407_1,
    new_n11408, new_n11409, new_n11410, new_n11411, new_n11412, new_n11413,
    new_n11414, new_n11415, new_n11416, new_n11417, new_n11418, new_n11419,
    new_n11420, new_n11421, new_n11422, new_n11423_1, new_n11424,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439, new_n11440, new_n11441, new_n11442,
    new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448,
    new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455, new_n11456, new_n11457, new_n11458, new_n11459, new_n11460,
    new_n11461, new_n11462, new_n11463, new_n11464, new_n11465, new_n11466,
    new_n11467, new_n11468, new_n11469, new_n11470, new_n11471, new_n11472,
    new_n11473, new_n11474, new_n11475, new_n11476, new_n11477,
    new_n11478_1, new_n11479, new_n11480, new_n11481, new_n11482,
    new_n11483, new_n11484, new_n11485, new_n11486, new_n11487, new_n11488,
    new_n11489, new_n11490, new_n11491, new_n11492, new_n11493, new_n11494,
    new_n11495, new_n11496, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503, new_n11504, new_n11505, new_n11506,
    new_n11507, new_n11508, new_n11509, new_n11510, new_n11511, new_n11512,
    new_n11513, new_n11514, new_n11515, new_n11516, new_n11517, new_n11518,
    new_n11519, new_n11520, new_n11521, new_n11522, new_n11523, new_n11524,
    new_n11525, new_n11526, new_n11527, new_n11528, new_n11529, new_n11530,
    new_n11531, new_n11532, new_n11533, new_n11534, new_n11535,
    new_n11536_1, new_n11537, new_n11538, new_n11539, new_n11540,
    new_n11541, new_n11542, new_n11543, new_n11544, new_n11545, new_n11546,
    new_n11547, new_n11548, new_n11549, new_n11550, new_n11551, new_n11552,
    new_n11553, new_n11554, new_n11555, new_n11556, new_n11557, new_n11558,
    new_n11559, new_n11560, new_n11561, new_n11562, new_n11563, new_n11564,
    new_n11565, new_n11566, new_n11567, new_n11568, new_n11569, new_n11570,
    new_n11571, new_n11572, new_n11573, new_n11574, new_n11575, new_n11576,
    new_n11577, new_n11578, new_n11579, new_n11580, new_n11581, new_n11582,
    new_n11583, new_n11584, new_n11585, new_n11586, new_n11587, new_n11588,
    new_n11589, new_n11590, new_n11591, new_n11592, new_n11593, new_n11594,
    new_n11595, new_n11596, new_n11598, new_n11599, new_n11600, new_n11602,
    new_n11603, new_n11604, new_n11606, new_n11608, new_n11609, new_n11610,
    new_n11612, new_n11614, new_n11615, new_n11616, new_n11617, new_n11618,
    new_n11619, new_n11620, new_n11621, new_n11622, new_n11623, new_n11624,
    new_n11625, new_n11626, new_n11627, new_n11628, new_n11629, new_n11630,
    new_n11631, new_n11632, new_n11633, new_n11634, new_n11635, new_n11636,
    new_n11637, new_n11638, new_n11639, new_n11640, new_n11641, new_n11642,
    new_n11643, new_n11644, new_n11645, new_n11646, new_n11647, new_n11648,
    new_n11649, new_n11650, new_n11651, new_n11652, new_n11653, new_n11654,
    new_n11655, new_n11656, new_n11657, new_n11658, new_n11659, new_n11660,
    new_n11661, new_n11662_1, new_n11663, new_n11664, new_n11665,
    new_n11666, new_n11667, new_n11668, new_n11669, new_n11670, new_n11671,
    new_n11672, new_n11673, new_n11674, new_n11675, new_n11676, new_n11677,
    new_n11678, new_n11679, new_n11680, new_n11681, new_n11682, new_n11683,
    new_n11684, new_n11685, new_n11686, new_n11687, new_n11688, new_n11689,
    new_n11690, new_n11691, new_n11692, new_n11693, new_n11694, new_n11695,
    new_n11696, new_n11697, new_n11698, new_n11699, new_n11700, new_n11701,
    new_n11702, new_n11703, new_n11704, new_n11705, new_n11706,
    new_n11707_1, new_n11708, new_n11709, new_n11710, new_n11711,
    new_n11712, new_n11713, new_n11714, new_n11715, new_n11716, new_n11717,
    new_n11718, new_n11719, new_n11720, new_n11721, new_n11722, new_n11723,
    new_n11724, new_n11725, new_n11726, new_n11727, new_n11728_1,
    new_n11729, new_n11730, new_n11731, new_n11732, new_n11733, new_n11734,
    new_n11735, new_n11736, new_n11737, new_n11738, new_n11739, new_n11740,
    new_n11741, new_n11742, new_n11743, new_n11744, new_n11745, new_n11746,
    new_n11747, new_n11748, new_n11749, new_n11750, new_n11751, new_n11752,
    new_n11753, new_n11754, new_n11755_1, new_n11756, new_n11757_1,
    new_n11758, new_n11759, new_n11760, new_n11761, new_n11762, new_n11763,
    new_n11764, new_n11765, new_n11766, new_n11767, new_n11768, new_n11769,
    new_n11770, new_n11771, new_n11772, new_n11773, new_n11774, new_n11775,
    new_n11776, new_n11777, new_n11778, new_n11779, new_n11780_1,
    new_n11781, new_n11782, new_n11783, new_n11784, new_n11785, new_n11786,
    new_n11787, new_n11788, new_n11789, new_n11790, new_n11791_1,
    new_n11792, new_n11793, new_n11794, new_n11795, new_n11796, new_n11797,
    new_n11798, new_n11799, new_n11800, new_n11801, new_n11802, new_n11803,
    new_n11804, new_n11805, new_n11806, new_n11807, new_n11808, new_n11809,
    new_n11810, new_n11811, new_n11812, new_n11813, new_n11814, new_n11815,
    new_n11816, new_n11817, new_n11818, new_n11819, new_n11820,
    new_n11821_1, new_n11822, new_n11823, new_n11824, new_n11825,
    new_n11826, new_n11827, new_n11828, new_n11829, new_n11830, new_n11831,
    new_n11832, new_n11833, new_n11834, new_n11835, new_n11836, new_n11837,
    new_n11838, new_n11839, new_n11840, new_n11841, new_n11842, new_n11843,
    new_n11844, new_n11845, new_n11846, new_n11847, new_n11848, new_n11849,
    new_n11850, new_n11851, new_n11852, new_n11853, new_n11854, new_n11855,
    new_n11856, new_n11857, new_n11858, new_n11859, new_n11860, new_n11861,
    new_n11862, new_n11863, new_n11864, new_n11865, new_n11866, new_n11867,
    new_n11868, new_n11869, new_n11870, new_n11871, new_n11872, new_n11873,
    new_n11874, new_n11875, new_n11876_1, new_n11877_1, new_n11878,
    new_n11879, new_n11880, new_n11881, new_n11882, new_n11883, new_n11884,
    new_n11885, new_n11886, new_n11887, new_n11888, new_n11889, new_n11890,
    new_n11891, new_n11892_1, new_n11893, new_n11894, new_n11895,
    new_n11896, new_n11897, new_n11898, new_n11899, new_n11900, new_n11901,
    new_n11902, new_n11903, new_n11904, new_n11905, new_n11906, new_n11907,
    new_n11908, new_n11909, new_n11910, new_n11911, new_n11912, new_n11913,
    new_n11914, new_n11915, new_n11916, new_n11917_1, new_n11918,
    new_n11919_1, new_n11920, new_n11921, new_n11922_1, new_n11923,
    new_n11924, new_n11925, new_n11926, new_n11927, new_n11928, new_n11929,
    new_n11930, new_n11931, new_n11932, new_n11933, new_n11934, new_n11935,
    new_n11936, new_n11937, new_n11938, new_n11939, new_n11940, new_n11941,
    new_n11942, new_n11943, new_n11944, new_n11945, new_n11946, new_n11947,
    new_n11948, new_n11949, new_n11950, new_n11951, new_n11952, new_n11953,
    new_n11954, new_n11955, new_n11956, new_n11957, new_n11958, new_n11959,
    new_n11960, new_n11961, new_n11962, new_n11963, new_n11964, new_n11965,
    new_n11966, new_n11967_1, new_n11968, new_n11969, new_n11970,
    new_n11971, new_n11972, new_n11973, new_n11974, new_n11975, new_n11976,
    new_n11977, new_n11978, new_n11979, new_n11980, new_n11981, new_n11982,
    new_n11983, new_n11984, new_n11985, new_n11986, new_n11987, new_n11988,
    new_n11989, new_n11990, new_n11991, new_n11992, new_n11993, new_n11994,
    new_n11995, new_n11996, new_n11997, new_n11998, new_n11999_1,
    new_n12000_1, new_n12001, new_n12002, new_n12003, new_n12004,
    new_n12005_1, new_n12006, new_n12007, new_n12008, new_n12009,
    new_n12010, new_n12011, new_n12012, new_n12013, new_n12014_1,
    new_n12015, new_n12016, new_n12017, new_n12018, new_n12019,
    new_n12020_1, new_n12021, new_n12022, new_n12023, new_n12024,
    new_n12025_1, new_n12026, new_n12027, new_n12028, new_n12029,
    new_n12030, new_n12031, new_n12032, new_n12033, new_n12034, new_n12035,
    new_n12036, new_n12037, new_n12038, new_n12039, new_n12040, new_n12041,
    new_n12042, new_n12043, new_n12044_1, new_n12045, new_n12046,
    new_n12047, new_n12048, new_n12049, new_n12050, new_n12051, new_n12052,
    new_n12053, new_n12054, new_n12055, new_n12056, new_n12057, new_n12058,
    new_n12059, new_n12060, new_n12061, new_n12062, new_n12063, new_n12064,
    new_n12065, new_n12066, new_n12067, new_n12068, new_n12069_1,
    new_n12070, new_n12071, new_n12072, new_n12073, new_n12074, new_n12075,
    new_n12076_1, new_n12077, new_n12078, new_n12079, new_n12080,
    new_n12081, new_n12082, new_n12083, new_n12084, new_n12085, new_n12086,
    new_n12087, new_n12088, new_n12089, new_n12090, new_n12091, new_n12092,
    new_n12093, new_n12094, new_n12095, new_n12096, new_n12097, new_n12098,
    new_n12099, new_n12100, new_n12101, new_n12102, new_n12103, new_n12104,
    new_n12105, new_n12106, new_n12107, new_n12108, new_n12109, new_n12110,
    new_n12111_1, new_n12112, new_n12113, new_n12114, new_n12115,
    new_n12116, new_n12117, new_n12118, new_n12119, new_n12120, new_n12121,
    new_n12122, new_n12123, new_n12124, new_n12125, new_n12126, new_n12127,
    new_n12128, new_n12129, new_n12130, new_n12131, new_n12132, new_n12133,
    new_n12134, new_n12135, new_n12136, new_n12137, new_n12138, new_n12139,
    new_n12140, new_n12141, new_n12142, new_n12143, new_n12144,
    new_n12145_1, new_n12146, new_n12147, new_n12148, new_n12149,
    new_n12150, new_n12151, new_n12152, new_n12153, new_n12154, new_n12155,
    new_n12156, new_n12157, new_n12158, new_n12159, new_n12160, new_n12161,
    new_n12162, new_n12163, new_n12164, new_n12165, new_n12166, new_n12167,
    new_n12168, new_n12169, new_n12170, new_n12171, new_n12172, new_n12173,
    new_n12174, new_n12175, new_n12176, new_n12177, new_n12178, new_n12179,
    new_n12180, new_n12181, new_n12182, new_n12183, new_n12184, new_n12185,
    new_n12186, new_n12187, new_n12188, new_n12189, new_n12190, new_n12191,
    new_n12192, new_n12193, new_n12194, new_n12195, new_n12196, new_n12197,
    new_n12198, new_n12199, new_n12200, new_n12201, new_n12202, new_n12203,
    new_n12204, new_n12205, new_n12206, new_n12207, new_n12208, new_n12209,
    new_n12210, new_n12211, new_n12212, new_n12213, new_n12214, new_n12215,
    new_n12216, new_n12217, new_n12218, new_n12219, new_n12220,
    new_n12221_1, new_n12222, new_n12223, new_n12224, new_n12225,
    new_n12226, new_n12227, new_n12228, new_n12229, new_n12230, new_n12231,
    new_n12232, new_n12233, new_n12234, new_n12235, new_n12236, new_n12237,
    new_n12238, new_n12239, new_n12240, new_n12241, new_n12242, new_n12243,
    new_n12244, new_n12245, new_n12246, new_n12247_1, new_n12248,
    new_n12249, new_n12250, new_n12251, new_n12252, new_n12253, new_n12255,
    new_n12256, new_n12257, new_n12259, new_n12260, new_n12261, new_n12263,
    new_n12264, new_n12265, new_n12266, new_n12267, new_n12268, new_n12269,
    new_n12270, new_n12271, new_n12272, new_n12273, new_n12274, new_n12275,
    new_n12276, new_n12277, new_n12278, new_n12279, new_n12280, new_n12281,
    new_n12282, new_n12283, new_n12284, new_n12285, new_n12286, new_n12287,
    new_n12288, new_n12289, new_n12290, new_n12291, new_n12292, new_n12293,
    new_n12294, new_n12295, new_n12296, new_n12297, new_n12298,
    new_n12299_1, new_n12300, new_n12301, new_n12302, new_n12303,
    new_n12304, new_n12305, new_n12306, new_n12307, new_n12308, new_n12309,
    new_n12310, new_n12311, new_n12312, new_n12313, new_n12314, new_n12315,
    new_n12316, new_n12317, new_n12318, new_n12319, new_n12320, new_n12321,
    new_n12322, new_n12323, new_n12324, new_n12325, new_n12326, new_n12327,
    new_n12328, new_n12329, new_n12330, new_n12331, new_n12332, new_n12333,
    new_n12334, new_n12335, new_n12336, new_n12337, new_n12338, new_n12339,
    new_n12340, new_n12341, new_n12342, new_n12343, new_n12344, new_n12345,
    new_n12346, new_n12347, new_n12348, new_n12349, new_n12350, new_n12351,
    new_n12352, new_n12353, new_n12354, new_n12355, new_n12356, new_n12357,
    new_n12358, new_n12359, new_n12360, new_n12361, new_n12362, new_n12363,
    new_n12364, new_n12365, new_n12366, new_n12367, new_n12368, new_n12369,
    new_n12370, new_n12371, new_n12372, new_n12373, new_n12374, new_n12375,
    new_n12376, new_n12377, new_n12378, new_n12379, new_n12380, new_n12381,
    new_n12382, new_n12383, new_n12384, new_n12385, new_n12386, new_n12387,
    new_n12388, new_n12389, new_n12390, new_n12391_1, new_n12392,
    new_n12393, new_n12394, new_n12395, new_n12396, new_n12397, new_n12398,
    new_n12399, new_n12400, new_n12401, new_n12402, new_n12403, new_n12405,
    new_n12406, new_n12407, new_n12408, new_n12409, new_n12410, new_n12411,
    new_n12412, new_n12413, new_n12414, new_n12415, new_n12416, new_n12417,
    new_n12418, new_n12419, new_n12420, new_n12421, new_n12422, new_n12423,
    new_n12424, new_n12425, new_n12426, new_n12427, new_n12428, new_n12429,
    new_n12430, new_n12431, new_n12432, new_n12433, new_n12434, new_n12435,
    new_n12436, new_n12437, new_n12438, new_n12439, new_n12440, new_n12441,
    new_n12442, new_n12443, new_n12444_1, new_n12445, new_n12446,
    new_n12447, new_n12448, new_n12449, new_n12450, new_n12451, new_n12452,
    new_n12453, new_n12454, new_n12455, new_n12456, new_n12457, new_n12458,
    new_n12459, new_n12460, new_n12461, new_n12462, new_n12463, new_n12464,
    new_n12465, new_n12466, new_n12467, new_n12468, new_n12469, new_n12470,
    new_n12471, new_n12472, new_n12473, new_n12474, new_n12475, new_n12476,
    new_n12477, new_n12478, new_n12479, new_n12480, new_n12481, new_n12482,
    new_n12483, new_n12484, new_n12485, new_n12486, new_n12487, new_n12488,
    new_n12489_1, new_n12490, new_n12491, new_n12492, new_n12493,
    new_n12494, new_n12495, new_n12496, new_n12497, new_n12498, new_n12499,
    new_n12500, new_n12501, new_n12502, new_n12503, new_n12504, new_n12505,
    new_n12506, new_n12507, new_n12508, new_n12509, new_n12510,
    new_n12511_1, new_n12512, new_n12513, new_n12514, new_n12515,
    new_n12516, new_n12517, new_n12518, new_n12519, new_n12520, new_n12521,
    new_n12522, new_n12523, new_n12524, new_n12525, new_n12526, new_n12527,
    new_n12528, new_n12529, new_n12530, new_n12531, new_n12532, new_n12533,
    new_n12534, new_n12535, new_n12536, new_n12537, new_n12538, new_n12539,
    new_n12540, new_n12541, new_n12542, new_n12543, new_n12544, new_n12545,
    new_n12546, new_n12547, new_n12548, new_n12549, new_n12550, new_n12551,
    new_n12552, new_n12553, new_n12554, new_n12555, new_n12556, new_n12557,
    new_n12558, new_n12559, new_n12560, new_n12561, new_n12562, new_n12563,
    new_n12564, new_n12565, new_n12566, new_n12567, new_n12568, new_n12569,
    new_n12570, new_n12571, new_n12572, new_n12573, new_n12574, new_n12575,
    new_n12576, new_n12577, new_n12578, new_n12579, new_n12580, new_n12581,
    new_n12582, new_n12583, new_n12584, new_n12585, new_n12586, new_n12587,
    new_n12588, new_n12589, new_n12590, new_n12591_1, new_n12592,
    new_n12593, new_n12594, new_n12595, new_n12596, new_n12597, new_n12598,
    new_n12599, new_n12600, new_n12601, new_n12602, new_n12603, new_n12604,
    new_n12605, new_n12606, new_n12607, new_n12608, new_n12609, new_n12610,
    new_n12611, new_n12612, new_n12613, new_n12614, new_n12615, new_n12616,
    new_n12617, new_n12618, new_n12619, new_n12620, new_n12621, new_n12622,
    new_n12623, new_n12624, new_n12625, new_n12626, new_n12627, new_n12628,
    new_n12629, new_n12630, new_n12631, new_n12632, new_n12633, new_n12634,
    new_n12635, new_n12636, new_n12637, new_n12638, new_n12639, new_n12640,
    new_n12641, new_n12642, new_n12643, new_n12644, new_n12645, new_n12646,
    new_n12647, new_n12648_1, new_n12649, new_n12650, new_n12651,
    new_n12652, new_n12653, new_n12654, new_n12655, new_n12656, new_n12657,
    new_n12658, new_n12659, new_n12660, new_n12661, new_n12662, new_n12663,
    new_n12664, new_n12665, new_n12666, new_n12667, new_n12668, new_n12669,
    new_n12670, new_n12671, new_n12672, new_n12673, new_n12674, new_n12675,
    new_n12676, new_n12677, new_n12678, new_n12679, new_n12680, new_n12681,
    new_n12682, new_n12683, new_n12684, new_n12685, new_n12686, new_n12687,
    new_n12688, new_n12689, new_n12690, new_n12691, new_n12692, new_n12693,
    new_n12694, new_n12695, new_n12696, new_n12697, new_n12698, new_n12699,
    new_n12700, new_n12701, new_n12702, new_n12703, new_n12704_1,
    new_n12705_1, new_n12706_1, new_n12707, new_n12708, new_n12709_1,
    new_n12710, new_n12711, new_n12712, new_n12713, new_n12714, new_n12715,
    new_n12716, new_n12717, new_n12718, new_n12719, new_n12720_1,
    new_n12721, new_n12722, new_n12723, new_n12724, new_n12725, new_n12726,
    new_n12727, new_n12728, new_n12729, new_n12730, new_n12731, new_n12732,
    new_n12733, new_n12734, new_n12735, new_n12736, new_n12737, new_n12738,
    new_n12739, new_n12740, new_n12741, new_n12742, new_n12743, new_n12744,
    new_n12745, new_n12746, new_n12747, new_n12748, new_n12749, new_n12750,
    new_n12751, new_n12752, new_n12753_1, new_n12754, new_n12755,
    new_n12756, new_n12757, new_n12758, new_n12759, new_n12760, new_n12761,
    new_n12762, new_n12763, new_n12764, new_n12765, new_n12766, new_n12767,
    new_n12768, new_n12769, new_n12770, new_n12771, new_n12772, new_n12773,
    new_n12774, new_n12775, new_n12776, new_n12777_1, new_n12778,
    new_n12779, new_n12780, new_n12781, new_n12782, new_n12783, new_n12784,
    new_n12785, new_n12786, new_n12787, new_n12788, new_n12789, new_n12790,
    new_n12791, new_n12792, new_n12793, new_n12794, new_n12795, new_n12796,
    new_n12797, new_n12798, new_n12799, new_n12800, new_n12801, new_n12802,
    new_n12803, new_n12804, new_n12805, new_n12806, new_n12807_1,
    new_n12808, new_n12809, new_n12810, new_n12811, new_n12812, new_n12813,
    new_n12814, new_n12815, new_n12816, new_n12817, new_n12818, new_n12819,
    new_n12820, new_n12821, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826_1, new_n12827, new_n12828, new_n12829, new_n12830,
    new_n12831, new_n12832, new_n12833, new_n12834, new_n12835, new_n12836,
    new_n12837, new_n12838, new_n12839, new_n12840, new_n12841, new_n12842,
    new_n12843, new_n12844, new_n12845, new_n12846, new_n12847, new_n12848,
    new_n12849, new_n12850, new_n12851, new_n12852, new_n12853, new_n12854,
    new_n12855, new_n12856, new_n12857, new_n12858, new_n12859, new_n12860,
    new_n12861, new_n12862, new_n12863, new_n12864, new_n12865, new_n12866,
    new_n12867, new_n12868, new_n12869, new_n12870, new_n12871, new_n12872,
    new_n12873, new_n12874, new_n12875, new_n12876, new_n12877, new_n12878,
    new_n12879, new_n12880, new_n12881, new_n12882, new_n12883, new_n12884,
    new_n12885, new_n12886, new_n12887, new_n12888, new_n12889, new_n12890,
    new_n12891, new_n12892, new_n12893, new_n12894, new_n12895, new_n12896,
    new_n12897, new_n12898, new_n12899, new_n12900, new_n12901, new_n12902,
    new_n12903, new_n12904, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914,
    new_n12915, new_n12916, new_n12917, new_n12918, new_n12919, new_n12920,
    new_n12921, new_n12922, new_n12923, new_n12924, new_n12925_1,
    new_n12926, new_n12927, new_n12928, new_n12929, new_n12930, new_n12931,
    new_n12932, new_n12933, new_n12934, new_n12935, new_n12936, new_n12937,
    new_n12938, new_n12939, new_n12940, new_n12941, new_n12942, new_n12943,
    new_n12944, new_n12945, new_n12946, new_n12947_1, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956, new_n12957, new_n12958, new_n12959, new_n12960,
    new_n12961, new_n12962, new_n12963, new_n12964, new_n12965, new_n12966,
    new_n12967, new_n12968, new_n12969, new_n12970, new_n12971, new_n12972,
    new_n12973, new_n12974, new_n12975, new_n12976, new_n12977, new_n12978,
    new_n12979, new_n12980, new_n12981, new_n12982, new_n12983, new_n12984,
    new_n12985, new_n12986, new_n12987, new_n12988, new_n12989, new_n12990,
    new_n12991, new_n12992, new_n12993, new_n12994, new_n12995, new_n12996,
    new_n12997, new_n12998, new_n12999, new_n13000, new_n13001, new_n13002,
    new_n13003, new_n13004, new_n13005, new_n13006, new_n13007, new_n13008,
    new_n13009, new_n13010, new_n13011, new_n13012, new_n13013, new_n13014,
    new_n13015, new_n13016, new_n13017, new_n13018, new_n13019, new_n13020,
    new_n13021, new_n13022, new_n13023, new_n13024, new_n13025, new_n13026,
    new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032,
    new_n13033, new_n13034, new_n13035, new_n13036, new_n13037, new_n13038,
    new_n13039, new_n13040, new_n13041, new_n13042, new_n13043, new_n13044,
    new_n13045, new_n13046, new_n13047, new_n13048, new_n13049, new_n13050,
    new_n13051, new_n13052, new_n13053, new_n13054, new_n13055, new_n13056,
    new_n13057, new_n13058, new_n13059, new_n13060, new_n13061, new_n13062,
    new_n13063, new_n13064, new_n13065, new_n13066, new_n13067, new_n13068,
    new_n13069, new_n13070, new_n13071, new_n13072, new_n13073, new_n13074,
    new_n13075, new_n13076, new_n13077, new_n13078, new_n13079, new_n13080,
    new_n13081, new_n13082, new_n13083, new_n13084, new_n13085, new_n13086,
    new_n13087, new_n13088, new_n13089, new_n13090, new_n13091, new_n13092,
    new_n13093, new_n13094, new_n13095, new_n13096, new_n13097, new_n13098,
    new_n13099, new_n13100, new_n13101, new_n13102, new_n13103, new_n13104,
    new_n13105, new_n13106, new_n13107, new_n13108, new_n13109, new_n13110,
    new_n13111, new_n13112, new_n13113, new_n13114, new_n13115, new_n13116,
    new_n13117, new_n13118, new_n13119, new_n13120, new_n13121, new_n13122,
    new_n13123, new_n13124, new_n13125, new_n13126, new_n13127, new_n13128,
    new_n13129, new_n13130, new_n13131, new_n13132, new_n13133, new_n13134,
    new_n13135, new_n13136, new_n13137, new_n13138, new_n13139, new_n13140,
    new_n13141, new_n13142, new_n13143, new_n13144, new_n13145, new_n13146,
    new_n13147, new_n13148, new_n13149, new_n13150, new_n13151, new_n13152,
    new_n13153, new_n13154, new_n13155, new_n13156, new_n13157, new_n13158,
    new_n13159, new_n13160, new_n13161, new_n13162, new_n13163, new_n13164,
    new_n13165, new_n13166, new_n13167, new_n13168, new_n13169, new_n13170,
    new_n13171, new_n13172, new_n13173, new_n13174, new_n13175, new_n13176,
    new_n13177, new_n13178, new_n13179, new_n13180, new_n13181, new_n13182,
    new_n13183, new_n13184, new_n13185, new_n13186, new_n13187, new_n13188,
    new_n13189, new_n13190, new_n13191, new_n13192, new_n13193, new_n13194,
    new_n13195, new_n13196, new_n13197, new_n13198, new_n13199, new_n13200,
    new_n13201, new_n13202, new_n13203, new_n13204, new_n13205, new_n13206,
    new_n13207, new_n13208, new_n13209, new_n13210, new_n13211, new_n13212,
    new_n13213, new_n13214, new_n13215, new_n13216, new_n13217, new_n13218,
    new_n13219, new_n13220, new_n13221, new_n13222, new_n13223, new_n13224,
    new_n13225, new_n13226, new_n13227, new_n13228, new_n13229, new_n13230,
    new_n13231, new_n13232, new_n13233, new_n13234, new_n13235, new_n13236,
    new_n13237, new_n13238, new_n13239, new_n13240, new_n13241, new_n13242,
    new_n13243, new_n13244, new_n13245, new_n13246, new_n13247, new_n13248,
    new_n13249, new_n13250, new_n13251, new_n13252, new_n13253, new_n13254,
    new_n13255, new_n13256, new_n13257, new_n13258, new_n13259, new_n13260,
    new_n13261, new_n13262, new_n13263, new_n13264, new_n13265, new_n13266,
    new_n13267, new_n13268, new_n13269, new_n13270, new_n13271, new_n13272,
    new_n13273, new_n13274, new_n13275, new_n13276, new_n13277, new_n13278,
    new_n13279, new_n13280, new_n13281, new_n13282, new_n13283, new_n13284,
    new_n13285, new_n13286, new_n13287, new_n13288, new_n13289, new_n13290,
    new_n13291, new_n13292, new_n13293, new_n13294, new_n13295, new_n13296,
    new_n13297, new_n13298, new_n13299, new_n13300, new_n13301, new_n13302,
    new_n13303, new_n13304, new_n13305, new_n13306, new_n13307, new_n13308,
    new_n13309, new_n13310, new_n13311, new_n13312, new_n13313, new_n13314,
    new_n13315, new_n13316, new_n13317, new_n13318, new_n13319, new_n13320,
    new_n13321, new_n13322, new_n13323, new_n13324, new_n13325, new_n13326,
    new_n13327, new_n13328, new_n13329, new_n13330, new_n13331, new_n13332,
    new_n13333, new_n13334, new_n13335, new_n13336, new_n13337, new_n13338,
    new_n13339, new_n13340, new_n13341, new_n13342, new_n13343, new_n13344,
    new_n13345, new_n13346, new_n13347, new_n13348, new_n13349, new_n13350,
    new_n13351, new_n13352, new_n13353, new_n13354, new_n13355, new_n13356,
    new_n13357, new_n13358, new_n13359, new_n13360, new_n13361, new_n13362,
    new_n13363, new_n13364, new_n13365, new_n13366, new_n13367, new_n13368,
    new_n13369, new_n13370, new_n13371, new_n13372, new_n13373, new_n13374,
    new_n13375, new_n13376, new_n13377, new_n13378, new_n13379, new_n13380,
    new_n13381, new_n13382, new_n13383, new_n13384, new_n13385, new_n13386,
    new_n13387, new_n13388, new_n13389, new_n13390, new_n13391, new_n13392,
    new_n13393, new_n13394, new_n13395, new_n13396, new_n13397, new_n13398,
    new_n13399, new_n13400, new_n13401, new_n13403, new_n13405, new_n13407,
    new_n13409, new_n13410, new_n13411, new_n13413, new_n13414, new_n13415,
    new_n13417, new_n13418, new_n13419, new_n13421, new_n13422, new_n13423,
    new_n13425, new_n13426, new_n13427, new_n13429, new_n13430, new_n13431,
    new_n13433, new_n13434, new_n13435, new_n13437, new_n13438, new_n13439,
    new_n13440, new_n13441, new_n13442, new_n13443, new_n13444, new_n13445,
    new_n13446, new_n13447, new_n13448, new_n13449, new_n13450, new_n13451,
    new_n13452, new_n13453, new_n13454, new_n13455, new_n13456, new_n13457,
    new_n13458, new_n13459, new_n13460, new_n13461, new_n13462, new_n13463,
    new_n13464, new_n13465, new_n13466, new_n13467, new_n13468, new_n13469,
    new_n13470, new_n13471, new_n13472, new_n13473, new_n13474, new_n13475,
    new_n13476, new_n13477, new_n13478, new_n13479, new_n13480, new_n13481,
    new_n13482, new_n13483, new_n13484, new_n13485, new_n13486, new_n13487,
    new_n13488, new_n13489, new_n13490, new_n13491, new_n13492, new_n13493,
    new_n13494, new_n13495, new_n13496, new_n13497, new_n13498, new_n13499,
    new_n13500, new_n13501, new_n13502, new_n13503, new_n13504, new_n13505,
    new_n13506, new_n13507, new_n13508, new_n13509, new_n13510, new_n13511,
    new_n13512, new_n13513, new_n13514, new_n13515, new_n13516, new_n13517,
    new_n13518, new_n13519, new_n13520, new_n13521, new_n13522, new_n13523,
    new_n13524, new_n13525, new_n13526, new_n13527, new_n13528, new_n13529,
    new_n13530, new_n13531, new_n13532, new_n13533, new_n13534, new_n13535,
    new_n13536, new_n13537, new_n13538, new_n13539, new_n13540, new_n13541,
    new_n13542, new_n13543, new_n13544, new_n13545, new_n13546, new_n13547,
    new_n13548, new_n13549, new_n13550, new_n13551, new_n13552, new_n13553,
    new_n13554, new_n13555, new_n13556, new_n13557, new_n13558, new_n13559,
    new_n13560, new_n13561, new_n13562, new_n13563, new_n13564, new_n13565,
    new_n13566, new_n13567, new_n13568, new_n13569, new_n13570, new_n13571,
    new_n13572, new_n13573, new_n13574, new_n13575, new_n13576, new_n13577,
    new_n13578, new_n13579, new_n13580, new_n13581, new_n13582, new_n13583,
    new_n13584, new_n13585, new_n13586, new_n13587, new_n13588, new_n13589,
    new_n13590, new_n13591, new_n13592, new_n13593, new_n13594, new_n13595,
    new_n13596, new_n13597, new_n13598, new_n13599, new_n13600, new_n13601,
    new_n13602, new_n13603, new_n13604, new_n13605, new_n13606, new_n13607,
    new_n13608, new_n13609, new_n13610, new_n13611, new_n13612, new_n13613,
    new_n13614, new_n13615, new_n13616, new_n13617, new_n13618, new_n13619,
    new_n13620, new_n13621, new_n13622, new_n13623, new_n13624, new_n13625,
    new_n13626, new_n13627, new_n13628, new_n13629, new_n13630, new_n13631,
    new_n13632, new_n13633, new_n13634, new_n13635, new_n13636, new_n13637,
    new_n13638, new_n13639, new_n13640, new_n13641, new_n13642, new_n13643,
    new_n13644, new_n13645, new_n13646, new_n13647, new_n13648, new_n13649,
    new_n13650, new_n13651, new_n13652, new_n13653, new_n13654, new_n13655,
    new_n13656, new_n13657, new_n13658, new_n13659, new_n13660, new_n13661,
    new_n13662, new_n13663, new_n13664, new_n13665, new_n13666, new_n13667,
    new_n13668, new_n13669, new_n13670, new_n13671, new_n13672, new_n13673,
    new_n13674, new_n13675, new_n13676, new_n13677, new_n13678, new_n13679,
    new_n13680, new_n13681, new_n13682, new_n13683, new_n13684, new_n13685,
    new_n13686, new_n13687, new_n13688, new_n13689, new_n13690, new_n13691,
    new_n13692, new_n13693, new_n13694, new_n13695, new_n13696, new_n13697,
    new_n13698, new_n13699, new_n13700, new_n13701, new_n13702, new_n13703,
    new_n13704, new_n13705, new_n13706, new_n13707, new_n13708, new_n13709,
    new_n13710, new_n13711, new_n13712, new_n13713, new_n13714, new_n13715,
    new_n13716, new_n13717, new_n13718, new_n13719, new_n13720, new_n13721,
    new_n13722, new_n13723, new_n13724, new_n13725, new_n13726, new_n13727,
    new_n13728, new_n13729, new_n13730, new_n13731, new_n13732, new_n13733,
    new_n13734, new_n13735, new_n13736, new_n13737, new_n13738, new_n13739,
    new_n13740, new_n13741, new_n13742, new_n13743, new_n13744, new_n13745,
    new_n13746, new_n13747, new_n13748, new_n13749, new_n13750, new_n13751,
    new_n13752, new_n13753, new_n13754, new_n13755, new_n13756, new_n13757,
    new_n13758, new_n13759, new_n13760, new_n13761, new_n13762, new_n13763,
    new_n13764, new_n13765, new_n13766, new_n13767, new_n13768, new_n13769,
    new_n13770, new_n13771, new_n13772, new_n13773, new_n13774, new_n13775,
    new_n13776, new_n13777, new_n13778, new_n13779, new_n13780, new_n13781,
    new_n13782, new_n13783, new_n13784, new_n13785, new_n13786, new_n13787,
    new_n13788, new_n13789, new_n13790, new_n13791, new_n13792, new_n13793,
    new_n13794, new_n13795, new_n13796, new_n13797, new_n13798, new_n13799,
    new_n13800, new_n13801, new_n13802, new_n13803, new_n13804, new_n13805,
    new_n13806, new_n13807, new_n13808, new_n13809, new_n13810, new_n13811,
    new_n13812, new_n13813, new_n13814, new_n13815, new_n13816, new_n13817,
    new_n13818, new_n13819, new_n13820, new_n13821, new_n13822, new_n13823,
    new_n13824, new_n13825, new_n13826, new_n13827, new_n13828, new_n13829,
    new_n13830, new_n13832, new_n13834, new_n13835, new_n13836, new_n13837,
    new_n13838, new_n13839, new_n13840, new_n13841, new_n13842, new_n13843,
    new_n13844, new_n13845, new_n13846, new_n13847, new_n13848, new_n13849,
    new_n13850, new_n13851, new_n13852, new_n13853, new_n13854, new_n13855,
    new_n13856, new_n13857, new_n13858, new_n13859, new_n13860, new_n13861,
    new_n13862, new_n13863, new_n13864, new_n13865, new_n13866, new_n13867,
    new_n13868, new_n13869, new_n13870, new_n13871, new_n13872, new_n13873,
    new_n13874, new_n13875, new_n13876, new_n13877, new_n13878, new_n13879,
    new_n13880, new_n13881, new_n13882, new_n13883, new_n13884, new_n13885,
    new_n13886, new_n13887, new_n13888, new_n13889, new_n13890, new_n13891,
    new_n13892, new_n13893, new_n13894, new_n13895, new_n13896, new_n13897,
    new_n13898, new_n13899, new_n13900, new_n13901, new_n13902, new_n13903,
    new_n13904, new_n13905, new_n13906, new_n13907, new_n13908, new_n13909,
    new_n13910, new_n13911, new_n13912, new_n13913, new_n13914, new_n13915,
    new_n13916, new_n13917, new_n13918, new_n13919, new_n13920, new_n13921,
    new_n13922, new_n13923, new_n13924, new_n13925, new_n13926, new_n13927,
    new_n13928, new_n13929, new_n13930, new_n13931, new_n13932, new_n13933,
    new_n13934, new_n13935, new_n13936, new_n13937, new_n13938, new_n13939,
    new_n13940, new_n13941, new_n13942, new_n13943, new_n13944, new_n13945,
    new_n13946, new_n13947, new_n13948, new_n13949, new_n13950, new_n13951,
    new_n13952, new_n13953, new_n13954, new_n13955, new_n13956, new_n13957,
    new_n13958, new_n13959, new_n13960, new_n13961, new_n13962, new_n13963,
    new_n13964, new_n13965, new_n13966, new_n13967, new_n13968, new_n13969,
    new_n13970, new_n13971, new_n13972, new_n13973, new_n13974, new_n13975,
    new_n13976, new_n13977, new_n13978, new_n13979, new_n13980, new_n13981,
    new_n13982, new_n13983, new_n13984, new_n13985, new_n13986, new_n13987,
    new_n13988, new_n13989, new_n13990, new_n13991, new_n13992, new_n13993,
    new_n13994, new_n13995, new_n13996, new_n13997, new_n13998, new_n13999,
    new_n14000, new_n14001, new_n14002, new_n14003, new_n14004, new_n14005,
    new_n14006, new_n14007, new_n14008, new_n14009, new_n14010, new_n14011,
    new_n14012, new_n14013, new_n14014, new_n14015, new_n14016, new_n14017,
    new_n14018, new_n14019, new_n14020, new_n14021, new_n14022, new_n14023,
    new_n14024, new_n14025, new_n14026, new_n14027, new_n14028, new_n14029,
    new_n14030, new_n14031, new_n14032, new_n14033, new_n14034, new_n14035,
    new_n14036, new_n14037, new_n14038, new_n14039, new_n14040, new_n14041,
    new_n14042, new_n14043, new_n14044, new_n14045, new_n14046, new_n14047,
    new_n14048, new_n14049, new_n14050, new_n14051, new_n14052, new_n14053,
    new_n14054, new_n14055, new_n14056, new_n14057, new_n14058, new_n14059,
    new_n14060, new_n14061, new_n14062, new_n14063, new_n14064, new_n14065,
    new_n14066, new_n14067, new_n14068, new_n14069, new_n14070, new_n14071,
    new_n14072, new_n14073, new_n14074, new_n14075, new_n14076, new_n14077,
    new_n14078, new_n14079, new_n14080, new_n14081, new_n14082, new_n14083,
    new_n14084, new_n14085, new_n14086, new_n14088, new_n14089, new_n14090,
    new_n14092, new_n14093, new_n14094, new_n14096, new_n14098, new_n14099,
    new_n14100, new_n14102, new_n14103, new_n14104, new_n14106, new_n14107,
    new_n14108, new_n14110, new_n14111, new_n14112, new_n14114, new_n14115,
    new_n14116, new_n14117, new_n14118, new_n14119, new_n14120, new_n14121,
    new_n14122, new_n14123, new_n14124, new_n14125, new_n14126, new_n14127,
    new_n14128, new_n14129, new_n14130, new_n14131, new_n14132, new_n14133,
    new_n14134, new_n14135, new_n14136, new_n14137, new_n14138, new_n14139,
    new_n14140, new_n14141, new_n14142, new_n14143, new_n14144, new_n14145,
    new_n14146, new_n14147, new_n14148, new_n14149, new_n14150, new_n14151,
    new_n14152, new_n14153, new_n14154, new_n14155, new_n14156, new_n14157,
    new_n14158, new_n14159, new_n14160, new_n14161, new_n14162, new_n14163,
    new_n14164, new_n14165, new_n14166, new_n14167, new_n14168, new_n14169,
    new_n14170, new_n14171, new_n14172, new_n14173, new_n14174, new_n14175,
    new_n14176, new_n14177, new_n14178, new_n14179, new_n14180, new_n14181,
    new_n14182, new_n14183, new_n14184, new_n14185, new_n14186, new_n14187,
    new_n14188, new_n14189, new_n14190, new_n14191, new_n14192, new_n14193,
    new_n14194, new_n14195, new_n14196, new_n14197, new_n14198, new_n14199,
    new_n14200, new_n14201, new_n14202, new_n14203, new_n14204, new_n14205,
    new_n14206, new_n14207, new_n14208, new_n14209, new_n14210, new_n14211,
    new_n14212, new_n14213, new_n14214, new_n14215, new_n14216, new_n14217,
    new_n14218, new_n14219, new_n14220, new_n14221, new_n14222, new_n14223,
    new_n14224, new_n14225, new_n14226, new_n14227, new_n14228, new_n14229,
    new_n14230, new_n14231, new_n14232, new_n14233, new_n14234, new_n14235,
    new_n14236, new_n14237, new_n14238, new_n14239, new_n14240, new_n14241,
    new_n14242, new_n14243, new_n14244, new_n14245, new_n14246, new_n14247,
    new_n14248, new_n14249, new_n14250, new_n14251, new_n14252, new_n14253,
    new_n14254, new_n14255, new_n14256, new_n14257, new_n14258, new_n14259,
    new_n14260, new_n14261, new_n14262, new_n14263, new_n14264, new_n14265,
    new_n14266, new_n14267, new_n14268, new_n14269, new_n14270, new_n14271,
    new_n14272, new_n14273, new_n14274, new_n14275, new_n14276, new_n14277,
    new_n14278, new_n14279, new_n14280, new_n14281, new_n14282, new_n14283,
    new_n14284, new_n14285, new_n14286, new_n14287, new_n14288, new_n14289,
    new_n14290, new_n14291, new_n14292, new_n14293, new_n14294, new_n14295,
    new_n14296, new_n14297, new_n14298, new_n14299, new_n14300, new_n14301,
    new_n14302, new_n14303, new_n14304, new_n14305, new_n14306, new_n14307,
    new_n14308, new_n14309, new_n14310, new_n14311, new_n14312, new_n14313,
    new_n14314, new_n14315, new_n14316, new_n14317, new_n14318, new_n14319,
    new_n14320, new_n14321, new_n14322, new_n14323, new_n14324, new_n14325,
    new_n14326, new_n14327, new_n14328, new_n14329, new_n14330, new_n14331,
    new_n14332, new_n14333, new_n14334, new_n14335, new_n14336, new_n14337,
    new_n14338, new_n14339, new_n14340, new_n14341, new_n14342, new_n14343,
    new_n14344, new_n14345, new_n14346, new_n14347, new_n14348, new_n14349,
    new_n14350, new_n14351, new_n14352, new_n14353, new_n14354, new_n14355,
    new_n14356, new_n14357, new_n14358, new_n14359, new_n14360, new_n14361,
    new_n14362, new_n14363, new_n14364, new_n14365, new_n14366, new_n14367,
    new_n14368, new_n14369, new_n14370, new_n14371, new_n14372, new_n14373,
    new_n14374, new_n14375, new_n14376, new_n14377, new_n14378, new_n14379,
    new_n14380, new_n14381, new_n14382, new_n14383, new_n14384, new_n14385,
    new_n14386, new_n14387, new_n14388, new_n14389, new_n14390, new_n14391,
    new_n14392, new_n14393, new_n14394, new_n14395, new_n14396, new_n14397,
    new_n14398, new_n14399, new_n14400, new_n14401, new_n14402, new_n14403,
    new_n14404, new_n14405, new_n14406, new_n14407, new_n14408, new_n14409,
    new_n14410, new_n14411, new_n14412, new_n14413, new_n14414, new_n14415,
    new_n14416, new_n14417, new_n14418, new_n14419, new_n14420, new_n14421,
    new_n14422, new_n14423, new_n14424, new_n14425, new_n14426, new_n14427,
    new_n14428, new_n14429, new_n14430, new_n14431, new_n14432, new_n14433,
    new_n14434, new_n14435, new_n14436, new_n14437, new_n14438, new_n14439,
    new_n14440, new_n14441, new_n14442, new_n14443, new_n14444, new_n14445,
    new_n14446, new_n14447, new_n14448, new_n14449, new_n14450, new_n14451,
    new_n14452, new_n14453, new_n14454, new_n14455, new_n14456, new_n14457,
    new_n14458, new_n14459, new_n14460, new_n14461, new_n14462, new_n14463,
    new_n14464, new_n14465, new_n14466, new_n14467, new_n14468, new_n14469,
    new_n14470, new_n14471, new_n14472, new_n14473, new_n14474, new_n14475,
    new_n14476, new_n14477, new_n14478, new_n14479, new_n14480, new_n14481,
    new_n14482, new_n14483, new_n14484, new_n14485, new_n14486, new_n14487,
    new_n14488, new_n14489, new_n14490, new_n14491, new_n14492, new_n14493,
    new_n14494, new_n14495, new_n14496, new_n14497, new_n14498, new_n14499,
    new_n14500, new_n14501, new_n14502, new_n14503, new_n14504, new_n14505,
    new_n14506, new_n14507, new_n14508, new_n14509, new_n14510, new_n14511,
    new_n14512, new_n14513, new_n14514, new_n14515, new_n14516, new_n14517,
    new_n14518, new_n14519, new_n14520, new_n14521, new_n14522, new_n14523,
    new_n14524, new_n14525, new_n14526, new_n14527, new_n14528, new_n14529,
    new_n14530, new_n14531, new_n14532, new_n14533, new_n14534, new_n14535,
    new_n14536, new_n14537, new_n14538, new_n14539, new_n14540, new_n14541,
    new_n14542, new_n14543, new_n14544, new_n14545, new_n14546, new_n14547,
    new_n14548, new_n14549, new_n14550, new_n14551, new_n14552, new_n14553,
    new_n14554, new_n14555, new_n14556, new_n14557, new_n14558, new_n14559,
    new_n14560, new_n14561, new_n14562, new_n14563, new_n14564, new_n14565,
    new_n14566, new_n14567, new_n14568, new_n14569, new_n14570, new_n14571,
    new_n14572, new_n14573, new_n14574, new_n14575, new_n14576, new_n14577,
    new_n14578, new_n14579, new_n14581, new_n14582, new_n14583, new_n14585,
    new_n14586, new_n14587, new_n14589, new_n14590, new_n14591, new_n14593,
    new_n14594, new_n14595, new_n14597, new_n14599, new_n14600, new_n14601,
    new_n14603, new_n14604, new_n14605, new_n14607, new_n14608, new_n14609,
    new_n14611, new_n14612, new_n14613, new_n14615, new_n14616, new_n14617,
    new_n14619, new_n14620, new_n14621, new_n14623, new_n14624, new_n14625,
    new_n14626, new_n14627, new_n14628, new_n14629, new_n14630, new_n14631,
    new_n14632, new_n14633, new_n14634, new_n14635, new_n14636, new_n14637,
    new_n14638, new_n14639, new_n14640, new_n14641, new_n14642, new_n14643,
    new_n14644, new_n14645, new_n14646, new_n14647, new_n14648, new_n14649,
    new_n14650, new_n14651, new_n14652, new_n14653, new_n14654, new_n14655,
    new_n14656, new_n14657, new_n14658, new_n14659, new_n14660, new_n14661,
    new_n14662, new_n14663, new_n14664, new_n14665, new_n14666, new_n14667,
    new_n14668, new_n14669, new_n14670, new_n14671, new_n14672, new_n14673,
    new_n14674, new_n14675, new_n14676, new_n14677, new_n14678, new_n14679,
    new_n14680, new_n14681, new_n14682, new_n14683, new_n14684, new_n14685,
    new_n14686, new_n14687, new_n14688, new_n14689, new_n14690, new_n14691,
    new_n14692, new_n14693, new_n14694, new_n14695, new_n14696, new_n14697,
    new_n14698, new_n14699, new_n14700, new_n14701, new_n14702, new_n14703,
    new_n14704, new_n14705, new_n14706, new_n14707, new_n14708, new_n14709,
    new_n14710, new_n14711, new_n14712, new_n14713, new_n14714, new_n14715,
    new_n14716, new_n14717, new_n14718, new_n14719, new_n14720, new_n14721,
    new_n14722, new_n14723, new_n14724, new_n14725, new_n14726, new_n14727,
    new_n14728, new_n14729, new_n14730, new_n14731, new_n14732, new_n14733,
    new_n14734, new_n14735, new_n14736, new_n14737, new_n14738, new_n14739,
    new_n14740, new_n14741, new_n14742, new_n14743, new_n14744, new_n14745,
    new_n14746, new_n14747, new_n14748, new_n14749, new_n14750, new_n14751,
    new_n14752, new_n14753, new_n14754, new_n14755, new_n14756, new_n14757,
    new_n14758, new_n14759, new_n14760, new_n14761, new_n14762, new_n14763,
    new_n14764, new_n14765, new_n14766, new_n14767, new_n14768, new_n14769,
    new_n14770, new_n14771, new_n14772, new_n14773, new_n14774, new_n14775,
    new_n14776, new_n14777, new_n14778, new_n14779, new_n14780, new_n14781,
    new_n14782, new_n14783, new_n14784, new_n14785, new_n14786, new_n14787,
    new_n14788, new_n14789, new_n14790, new_n14791, new_n14792, new_n14793,
    new_n14794, new_n14795, new_n14796, new_n14797, new_n14798, new_n14799,
    new_n14800, new_n14801, new_n14802, new_n14803, new_n14804, new_n14805,
    new_n14806, new_n14807, new_n14808, new_n14809, new_n14810, new_n14811,
    new_n14812, new_n14813, new_n14814, new_n14815, new_n14816, new_n14817,
    new_n14818, new_n14819, new_n14820, new_n14821, new_n14822, new_n14823,
    new_n14824, new_n14825, new_n14826, new_n14827, new_n14828, new_n14829,
    new_n14830, new_n14831, new_n14832, new_n14833, new_n14834, new_n14835,
    new_n14836, new_n14837, new_n14838, new_n14839, new_n14840, new_n14841,
    new_n14842, new_n14843, new_n14844, new_n14845, new_n14846, new_n14847,
    new_n14848, new_n14849, new_n14850, new_n14851, new_n14852, new_n14853,
    new_n14854, new_n14855, new_n14856, new_n14857, new_n14858, new_n14859,
    new_n14860, new_n14861, new_n14862, new_n14863, new_n14864, new_n14865,
    new_n14866, new_n14867, new_n14868, new_n14869, new_n14870, new_n14871,
    new_n14872, new_n14874, new_n14875, new_n14876, new_n14878, new_n14879,
    new_n14880, new_n14881, new_n14882, new_n14883, new_n14884, new_n14885,
    new_n14886, new_n14887, new_n14888, new_n14889, new_n14890, new_n14891,
    new_n14892, new_n14893, new_n14894, new_n14895, new_n14896, new_n14897,
    new_n14898, new_n14899, new_n14900, new_n14901, new_n14902, new_n14903,
    new_n14904, new_n14905, new_n14906, new_n14907, new_n14908, new_n14909,
    new_n14910, new_n14911, new_n14912, new_n14913, new_n14914, new_n14915,
    new_n14916, new_n14917, new_n14918, new_n14919, new_n14920, new_n14921,
    new_n14922, new_n14923, new_n14924, new_n14925, new_n14926, new_n14927,
    new_n14928, new_n14929, new_n14930, new_n14931, new_n14932, new_n14933,
    new_n14934, new_n14935, new_n14936, new_n14937, new_n14938, new_n14939,
    new_n14940, new_n14941, new_n14942, new_n14943, new_n14944, new_n14945,
    new_n14946, new_n14947, new_n14948, new_n14949, new_n14950, new_n14951,
    new_n14952, new_n14953, new_n14954, new_n14955, new_n14956, new_n14957,
    new_n14958, new_n14959, new_n14960, new_n14961, new_n14962, new_n14963,
    new_n14964, new_n14965, new_n14966, new_n14967, new_n14968, new_n14969,
    new_n14970, new_n14971, new_n14972, new_n14973, new_n14974, new_n14975,
    new_n14976, new_n14977, new_n14978, new_n14979, new_n14980, new_n14981,
    new_n14982, new_n14983, new_n14984, new_n14985, new_n14986, new_n14987,
    new_n14988, new_n14989, new_n14990, new_n14991, new_n14992, new_n14993,
    new_n14994, new_n14995, new_n14996, new_n14997, new_n14998, new_n14999,
    new_n15000, new_n15001, new_n15002, new_n15003, new_n15004, new_n15005,
    new_n15006, new_n15007, new_n15008, new_n15009, new_n15010, new_n15011,
    new_n15012, new_n15013, new_n15014, new_n15015, new_n15016, new_n15017,
    new_n15018, new_n15019, new_n15020, new_n15021, new_n15022, new_n15023,
    new_n15024, new_n15025, new_n15026, new_n15027, new_n15028, new_n15029,
    new_n15030, new_n15031, new_n15032, new_n15033, new_n15034, new_n15035,
    new_n15036, new_n15037, new_n15038, new_n15039, new_n15040, new_n15041,
    new_n15042, new_n15043, new_n15044, new_n15045, new_n15046, new_n15047,
    new_n15048, new_n15049, new_n15050, new_n15051, new_n15052, new_n15053,
    new_n15054, new_n15055, new_n15056, new_n15057, new_n15058, new_n15059,
    new_n15060, new_n15061, new_n15062, new_n15063, new_n15064, new_n15065,
    new_n15066, new_n15067, new_n15068, new_n15069, new_n15070, new_n15071,
    new_n15072, new_n15073, new_n15074, new_n15075, new_n15076, new_n15077,
    new_n15078, new_n15079, new_n15080, new_n15081, new_n15082, new_n15083,
    new_n15084, new_n15085, new_n15086, new_n15087, new_n15088, new_n15089,
    new_n15090, new_n15091, new_n15092, new_n15093, new_n15094, new_n15095,
    new_n15096, new_n15097, new_n15098, new_n15099, new_n15100, new_n15101,
    new_n15102, new_n15103, new_n15104, new_n15105, new_n15106, new_n15107,
    new_n15108, new_n15109, new_n15110, new_n15111, new_n15112, new_n15113,
    new_n15114, new_n15115, new_n15116, new_n15117, new_n15118, new_n15119,
    new_n15120, new_n15121, new_n15122, new_n15123, new_n15124, new_n15125,
    new_n15126, new_n15127, new_n15128, new_n15129, new_n15131, new_n15132,
    new_n15133, new_n15135, new_n15136, new_n15137, new_n15139, new_n15141,
    new_n15142, new_n15143, new_n15145, new_n15146, new_n15147, new_n15149,
    new_n15150, new_n15151, new_n15153, new_n15154, new_n15155, new_n15157,
    new_n15158, new_n15159, new_n15161, new_n15162, new_n15163, new_n15165,
    new_n15166, new_n15167, new_n15169, new_n15170, new_n15171, new_n15172,
    new_n15173, new_n15174, new_n15175, new_n15176, new_n15177, new_n15178,
    new_n15179, new_n15180, new_n15181, new_n15182, new_n15183, new_n15184,
    new_n15185, new_n15186, new_n15187, new_n15188, new_n15189, new_n15190,
    new_n15191, new_n15192, new_n15193, new_n15194, new_n15195, new_n15196,
    new_n15197, new_n15198, new_n15199, new_n15200, new_n15201, new_n15202,
    new_n15203, new_n15204, new_n15205, new_n15206, new_n15207, new_n15208,
    new_n15209, new_n15210, new_n15211, new_n15212, new_n15213, new_n15214,
    new_n15215, new_n15216, new_n15217, new_n15218, new_n15219, new_n15220,
    new_n15221, new_n15222, new_n15223, new_n15224, new_n15225, new_n15226,
    new_n15227, new_n15228, new_n15229, new_n15230, new_n15231, new_n15232,
    new_n15233, new_n15234, new_n15235, new_n15236, new_n15237, new_n15238,
    new_n15239, new_n15240, new_n15241, new_n15242, new_n15243, new_n15244,
    new_n15245, new_n15246, new_n15247, new_n15248, new_n15249, new_n15250,
    new_n15251, new_n15252, new_n15253, new_n15254, new_n15255, new_n15256,
    new_n15257, new_n15258, new_n15259, new_n15260, new_n15261, new_n15262,
    new_n15263, new_n15264, new_n15265, new_n15266, new_n15267, new_n15268,
    new_n15269, new_n15270, new_n15271, new_n15272, new_n15273, new_n15274,
    new_n15275, new_n15276, new_n15277, new_n15278, new_n15279, new_n15280,
    new_n15281, new_n15282, new_n15283, new_n15284, new_n15285, new_n15286,
    new_n15287, new_n15288, new_n15289, new_n15290, new_n15291, new_n15292,
    new_n15293, new_n15294, new_n15295, new_n15296, new_n15297, new_n15298,
    new_n15299, new_n15300, new_n15301, new_n15302, new_n15303, new_n15304,
    new_n15305, new_n15306, new_n15307, new_n15308, new_n15309, new_n15310,
    new_n15311, new_n15312, new_n15313, new_n15314, new_n15315, new_n15316,
    new_n15317, new_n15318, new_n15319, new_n15320, new_n15321, new_n15322,
    new_n15323, new_n15324, new_n15325, new_n15326, new_n15327, new_n15328,
    new_n15329, new_n15330, new_n15331, new_n15332, new_n15333, new_n15334,
    new_n15335, new_n15336, new_n15337, new_n15338, new_n15339, new_n15340,
    new_n15341, new_n15342, new_n15343, new_n15344, new_n15345, new_n15346,
    new_n15347, new_n15348, new_n15349, new_n15350, new_n15351, new_n15352,
    new_n15353, new_n15354, new_n15355, new_n15356, new_n15357, new_n15358,
    new_n15359, new_n15360, new_n15361, new_n15362, new_n15363, new_n15364,
    new_n15365, new_n15366, new_n15367, new_n15368, new_n15369, new_n15370,
    new_n15371, new_n15372, new_n15373, new_n15374, new_n15375, new_n15376,
    new_n15377, new_n15378, new_n15379, new_n15380, new_n15381, new_n15382,
    new_n15383, new_n15384, new_n15385, new_n15386, new_n15387, new_n15388,
    new_n15389, new_n15390, new_n15391, new_n15392, new_n15393, new_n15394,
    new_n15395, new_n15396, new_n15397, new_n15398, new_n15399, new_n15400,
    new_n15401, new_n15402, new_n15403, new_n15404, new_n15405, new_n15406,
    new_n15407, new_n15408, new_n15409, new_n15410, new_n15411, new_n15412,
    new_n15413, new_n15414, new_n15415, new_n15416, new_n15417, new_n15418,
    new_n15419, new_n15420, new_n15421, new_n15423, new_n15424, new_n15425,
    new_n15427, new_n15428, new_n15429, new_n15431, new_n15432, new_n15433,
    new_n15435, new_n15436, new_n15437, new_n15439, new_n15440, new_n15441,
    new_n15443, new_n15444, new_n15445, new_n15447, new_n15449, new_n15450,
    new_n15451, new_n15453, new_n15454, new_n15455, new_n15457, new_n15458,
    new_n15459, new_n15461, new_n15463, new_n15464, new_n15465, new_n15466,
    new_n15467, new_n15468, new_n15469, new_n15470, new_n15471, new_n15472,
    new_n15473, new_n15474, new_n15475, new_n15476, new_n15477, new_n15478,
    new_n15479, new_n15480, new_n15481, new_n15482, new_n15483, new_n15484,
    new_n15485, new_n15486, new_n15487, new_n15488, new_n15489, new_n15490,
    new_n15491, new_n15492, new_n15493, new_n15494, new_n15495, new_n15496,
    new_n15497, new_n15498, new_n15499, new_n15500, new_n15501, new_n15502,
    new_n15503, new_n15504, new_n15505, new_n15506, new_n15507, new_n15508,
    new_n15509, new_n15510, new_n15511, new_n15512, new_n15513, new_n15514,
    new_n15515, new_n15516, new_n15517, new_n15518, new_n15519, new_n15520,
    new_n15521, new_n15522, new_n15523, new_n15524, new_n15525, new_n15526,
    new_n15527, new_n15528, new_n15529, new_n15530, new_n15531, new_n15532,
    new_n15533, new_n15534, new_n15535, new_n15536, new_n15537, new_n15538,
    new_n15539, new_n15540, new_n15541, new_n15542, new_n15543, new_n15544,
    new_n15545, new_n15546, new_n15547, new_n15548, new_n15549, new_n15550,
    new_n15551, new_n15552, new_n15553, new_n15554, new_n15555, new_n15556,
    new_n15557, new_n15558, new_n15559, new_n15560, new_n15561, new_n15562,
    new_n15563, new_n15564, new_n15565, new_n15566, new_n15567, new_n15568,
    new_n15569, new_n15570, new_n15571, new_n15572, new_n15573, new_n15574,
    new_n15575, new_n15576, new_n15577, new_n15578, new_n15579, new_n15580,
    new_n15581, new_n15582, new_n15583, new_n15584, new_n15585, new_n15586,
    new_n15587, new_n15588, new_n15589, new_n15590, new_n15591, new_n15592,
    new_n15593, new_n15594, new_n15595, new_n15596, new_n15597, new_n15598,
    new_n15599, new_n15600, new_n15601, new_n15602, new_n15603, new_n15604,
    new_n15605, new_n15606, new_n15607, new_n15608, new_n15609, new_n15610,
    new_n15611, new_n15612, new_n15613, new_n15614, new_n15615, new_n15616,
    new_n15617, new_n15618, new_n15619, new_n15620, new_n15621, new_n15622,
    new_n15623, new_n15624, new_n15625, new_n15626, new_n15627, new_n15628,
    new_n15629, new_n15630, new_n15631, new_n15632, new_n15633, new_n15634,
    new_n15635, new_n15636, new_n15637, new_n15638, new_n15639, new_n15640,
    new_n15641, new_n15642, new_n15643, new_n15644, new_n15645, new_n15646,
    new_n15647, new_n15648, new_n15649, new_n15650, new_n15651, new_n15652,
    new_n15653, new_n15654, new_n15655, new_n15656, new_n15657, new_n15658,
    new_n15659, new_n15660, new_n15661, new_n15662, new_n15663, new_n15664,
    new_n15665, new_n15666, new_n15667, new_n15668, new_n15669, new_n15670,
    new_n15671, new_n15672, new_n15673, new_n15674, new_n15675, new_n15676,
    new_n15677, new_n15678, new_n15679, new_n15680, new_n15681, new_n15682,
    new_n15683, new_n15684, new_n15685, new_n15686, new_n15687, new_n15688,
    new_n15689, new_n15690, new_n15691, new_n15692, new_n15693, new_n15694,
    new_n15695, new_n15696, new_n15697, new_n15698, new_n15699, new_n15700,
    new_n15701, new_n15702, new_n15703, new_n15704, new_n15705, new_n15706,
    new_n15707, new_n15708, new_n15709, new_n15710, new_n15711, new_n15712,
    new_n15713, new_n15715, new_n15716, new_n15717, new_n15719, new_n15720,
    new_n15721, new_n15723, new_n15724, new_n15725, new_n15727, new_n15728,
    new_n15729, new_n15731, new_n15732, new_n15733, new_n15735, new_n15736,
    new_n15737, new_n15739, new_n15740, new_n15741, new_n15743, new_n15744,
    new_n15745, new_n15747, new_n15748, new_n15749, new_n15751, new_n15752,
    new_n15753;
  assign new_n377 = n6038 & n6687;
  assign new_n378 = n7354 & n8336;
  assign new_n379 = n8028 & n11222;
  assign new_n380 = n1564 & n12069;
  assign new_n381_1 = new_n379 & new_n380;
  assign new_n382 = ~new_n379 & ~new_n380;
  assign new_n383 = ~new_n381_1 & ~new_n382;
  assign new_n384 = new_n378 & new_n383;
  assign new_n385 = ~new_n378 & ~new_n383;
  assign new_n386 = ~new_n384 & ~new_n385;
  assign new_n387 = new_n377 & new_n386;
  assign new_n388 = ~new_n377 & ~new_n386;
  assign n112 = ~new_n387 & ~new_n388;
  assign new_n390 = n4005 & n5305;
  assign new_n391 = n2585 & n5305;
  assign new_n392 = n2508 & n5964;
  assign new_n393 = n2509 & n4312;
  assign new_n394 = n1097 & n12720;
  assign new_n395 = n6038 & n12705;
  assign new_n396 = ~new_n394 & ~new_n395;
  assign new_n397_1 = new_n394 & new_n395;
  assign new_n398 = ~new_n396 & ~new_n397_1;
  assign new_n399 = new_n393 & ~new_n398;
  assign new_n400 = ~new_n393 & new_n398;
  assign new_n401 = ~new_n399 & ~new_n400;
  assign new_n402 = ~new_n392 & new_n401;
  assign new_n403 = new_n392 & ~new_n401;
  assign new_n404 = ~new_n402 & ~new_n403;
  assign new_n405_1 = n5964 & n12720;
  assign new_n406 = n1097 & n2509;
  assign new_n407 = new_n405_1 & new_n406;
  assign new_n408 = ~new_n405_1 & ~new_n406;
  assign new_n409 = n4312 & n6038;
  assign new_n410 = ~new_n408 & new_n409;
  assign new_n411 = ~new_n407 & ~new_n410;
  assign new_n412 = new_n404 & ~new_n411;
  assign new_n413 = ~new_n404 & new_n411;
  assign new_n414 = ~new_n412 & ~new_n413;
  assign new_n415 = new_n391 & new_n414;
  assign new_n416 = ~new_n391 & ~new_n414;
  assign new_n417 = n2508 & n5305;
  assign new_n418 = n2509 & n5964;
  assign new_n419 = n5305 & n12720;
  assign new_n420 = new_n418 & new_n419;
  assign new_n421 = n1097 & n6038;
  assign new_n422 = ~new_n418 & ~new_n419;
  assign new_n423 = new_n421 & ~new_n422;
  assign new_n424 = ~new_n420 & ~new_n423;
  assign new_n425 = ~new_n417 & new_n424;
  assign new_n426 = new_n417 & ~new_n424;
  assign new_n427 = ~new_n407 & ~new_n408;
  assign new_n428 = ~new_n409 & ~new_n427;
  assign new_n429 = new_n409 & new_n427;
  assign new_n430 = ~new_n428 & ~new_n429;
  assign new_n431 = ~new_n426 & ~new_n430;
  assign new_n432 = ~new_n425 & ~new_n431;
  assign new_n433 = ~new_n416 & new_n432;
  assign new_n434 = ~new_n415 & ~new_n433;
  assign new_n435 = n1097 & n2508;
  assign new_n436 = n2585 & n5964;
  assign new_n437 = ~new_n435 & ~new_n436;
  assign new_n438 = new_n435 & new_n436;
  assign new_n439 = ~new_n437 & ~new_n438;
  assign new_n440 = n4312 & n12720;
  assign new_n441 = n6038 & n12025;
  assign new_n442 = n2509 & n12705;
  assign new_n443 = ~new_n441 & ~new_n442;
  assign new_n444 = new_n441 & new_n442;
  assign new_n445 = ~new_n443 & ~new_n444;
  assign new_n446 = ~new_n440 & ~new_n445;
  assign new_n447_1 = new_n393 & ~new_n396;
  assign new_n448 = ~new_n397_1 & ~new_n447_1;
  assign new_n449 = new_n446 & new_n448;
  assign new_n450 = new_n440 & new_n445;
  assign new_n451 = new_n448 & ~new_n450;
  assign new_n452 = ~new_n446 & ~new_n451;
  assign new_n453 = ~new_n449 & ~new_n452;
  assign new_n454 = ~new_n448 & new_n450;
  assign new_n455 = ~new_n453 & ~new_n454;
  assign new_n456 = new_n439 & ~new_n455;
  assign new_n457 = ~new_n439 & new_n455;
  assign new_n458 = ~new_n456 & ~new_n457;
  assign new_n459 = ~new_n402 & ~new_n411;
  assign new_n460 = ~new_n403 & ~new_n459;
  assign new_n461 = ~new_n458 & ~new_n460;
  assign new_n462 = new_n458 & new_n460;
  assign new_n463 = ~new_n461 & ~new_n462;
  assign new_n464 = ~new_n434 & ~new_n463;
  assign new_n465 = new_n434 & new_n463;
  assign new_n466 = ~new_n464 & ~new_n465;
  assign new_n467 = new_n390 & new_n466;
  assign new_n468 = n2509 & n5305;
  assign new_n469 = n5964 & n6038;
  assign new_n470 = new_n468 & new_n469;
  assign new_n471 = ~new_n420 & ~new_n422;
  assign new_n472 = ~new_n421 & ~new_n471;
  assign new_n473 = new_n421 & new_n471;
  assign new_n474 = ~new_n472 & ~new_n473;
  assign new_n475 = new_n470 & new_n474;
  assign new_n476 = ~new_n425 & ~new_n426;
  assign new_n477 = new_n430 & ~new_n476;
  assign new_n478 = ~new_n430 & new_n476;
  assign new_n479 = ~new_n477 & ~new_n478;
  assign new_n480 = new_n475 & ~new_n479;
  assign new_n481 = ~new_n415 & new_n433;
  assign new_n482 = ~new_n415 & ~new_n416;
  assign new_n483 = ~new_n432 & ~new_n482;
  assign new_n484 = ~new_n481 & ~new_n483;
  assign new_n485 = new_n480 & new_n484;
  assign new_n486 = ~new_n390 & ~new_n466;
  assign new_n487 = ~new_n467 & ~new_n486;
  assign new_n488 = new_n485 & new_n487;
  assign new_n489 = ~new_n467 & ~new_n488;
  assign new_n490 = ~new_n457 & ~new_n460;
  assign new_n491 = ~new_n438 & ~new_n490;
  assign new_n492 = ~new_n456 & new_n491;
  assign new_n493 = new_n438 & new_n490;
  assign new_n494 = ~new_n492 & ~new_n493;
  assign new_n495 = n1097 & n2585;
  assign new_n496 = n5305 & n12706;
  assign new_n497 = n4005 & n5964;
  assign new_n498 = ~new_n496 & ~new_n497;
  assign new_n499 = new_n496 & new_n497;
  assign new_n500 = ~new_n498 & ~new_n499;
  assign new_n501 = new_n495 & ~new_n500;
  assign new_n502 = ~new_n495 & new_n500;
  assign new_n503_1 = ~new_n501 & ~new_n502;
  assign new_n504 = new_n452 & ~new_n503_1;
  assign new_n505 = ~new_n452 & new_n503_1;
  assign new_n506 = ~new_n504 & ~new_n505;
  assign new_n507 = n2508 & n4312;
  assign new_n508 = new_n444 & new_n507;
  assign new_n509 = ~new_n444 & ~new_n507;
  assign new_n510 = ~new_n508 & ~new_n509;
  assign new_n511 = n2509 & n12025;
  assign new_n512 = n12705 & n12720;
  assign new_n513 = n6038 & n11257;
  assign new_n514 = ~new_n512 & ~new_n513;
  assign new_n515 = new_n512 & new_n513;
  assign new_n516 = ~new_n514 & ~new_n515;
  assign new_n517 = ~new_n511 & ~new_n516;
  assign new_n518 = new_n511 & new_n516;
  assign new_n519 = ~new_n517 & ~new_n518;
  assign new_n520 = new_n510 & ~new_n519;
  assign new_n521_1 = ~new_n510 & new_n519;
  assign new_n522 = ~new_n520 & ~new_n521_1;
  assign new_n523 = ~new_n506 & ~new_n522;
  assign new_n524 = new_n506 & new_n522;
  assign new_n525 = ~new_n523 & ~new_n524;
  assign new_n526 = ~new_n494 & new_n525;
  assign new_n527 = new_n494 & ~new_n525;
  assign new_n528 = ~new_n526 & ~new_n527;
  assign new_n529 = ~new_n464 & ~new_n528;
  assign new_n530 = new_n464 & new_n528;
  assign new_n531 = ~new_n529 & ~new_n530;
  assign new_n532 = ~new_n489 & new_n531;
  assign new_n533_1 = new_n489 & ~new_n531;
  assign new_n534 = ~new_n532 & ~new_n533_1;
  assign new_n535 = ~new_n485 & ~new_n487;
  assign new_n536 = ~new_n488 & ~new_n535;
  assign new_n537 = n1564 & n8476;
  assign new_n538 = n1512 & n5331;
  assign new_n539 = new_n537 & new_n538;
  assign new_n540 = n1564 & n2530;
  assign new_n541 = n533 & n5331;
  assign new_n542 = ~new_n540 & ~new_n541;
  assign new_n543 = n1564 & n5331;
  assign new_n544 = n533 & n2530;
  assign new_n545 = new_n543 & new_n544;
  assign new_n546 = ~new_n542 & ~new_n545;
  assign new_n547 = new_n539 & ~new_n546;
  assign new_n548 = n2802 & n5331;
  assign new_n549 = n1512 & n8476;
  assign new_n550 = ~new_n545 & ~new_n549;
  assign new_n551 = ~new_n542 & ~new_n550;
  assign new_n552 = new_n548 & new_n551;
  assign new_n553 = ~new_n548 & ~new_n551;
  assign new_n554 = ~new_n552 & ~new_n553;
  assign new_n555 = n1512 & n2530;
  assign new_n556 = n1564 & n12648;
  assign new_n557 = n533 & n8476;
  assign new_n558 = ~new_n556 & ~new_n557;
  assign new_n559 = new_n556 & new_n557;
  assign new_n560 = ~new_n558 & ~new_n559;
  assign new_n561 = new_n555 & ~new_n560;
  assign new_n562 = ~new_n555 & new_n560;
  assign new_n563 = ~new_n561 & ~new_n562;
  assign new_n564 = ~new_n554 & ~new_n563;
  assign new_n565 = new_n554 & new_n563;
  assign new_n566 = ~new_n564 & ~new_n565;
  assign new_n567 = new_n547 & ~new_n566;
  assign new_n568 = n5331 & n6806;
  assign new_n569 = n2802 & n8476;
  assign new_n570 = new_n555 & ~new_n558;
  assign new_n571 = ~new_n559 & ~new_n570;
  assign new_n572 = new_n569 & ~new_n571;
  assign new_n573 = ~new_n569 & new_n571;
  assign new_n574 = ~new_n572 & ~new_n573;
  assign new_n575 = n1512 & n12648;
  assign new_n576 = n1564 & n10545;
  assign new_n577 = ~new_n544 & ~new_n576;
  assign new_n578 = n533 & n10545;
  assign new_n579 = new_n540 & new_n578;
  assign new_n580 = ~new_n577 & ~new_n579;
  assign new_n581 = ~new_n575 & new_n580;
  assign new_n582 = new_n575 & ~new_n580;
  assign new_n583 = ~new_n581 & ~new_n582;
  assign new_n584 = ~new_n574 & ~new_n583;
  assign new_n585 = new_n574 & new_n583;
  assign new_n586 = ~new_n584 & ~new_n585;
  assign new_n587 = new_n568 & ~new_n586;
  assign new_n588 = ~new_n568 & new_n586;
  assign new_n589 = ~new_n587 & ~new_n588;
  assign new_n590 = ~new_n553 & ~new_n563;
  assign new_n591 = ~new_n552 & ~new_n590;
  assign new_n592 = ~new_n589 & ~new_n591;
  assign new_n593 = new_n589 & new_n591;
  assign new_n594 = ~new_n592 & ~new_n593;
  assign new_n595 = new_n567 & ~new_n594;
  assign new_n596 = n5069 & n5331;
  assign new_n597 = ~new_n588 & ~new_n591;
  assign new_n598 = ~new_n587 & ~new_n597;
  assign new_n599 = n6806 & n8476;
  assign new_n600 = n2530 & n2802;
  assign new_n601 = ~new_n599 & ~new_n600;
  assign new_n602 = new_n599 & new_n600;
  assign new_n603 = ~new_n601 & ~new_n602;
  assign new_n604 = n533 & n12648;
  assign new_n605 = n1512 & n10545;
  assign new_n606 = n1564 & n7690;
  assign new_n607 = ~new_n605 & ~new_n606;
  assign new_n608 = new_n605 & new_n606;
  assign new_n609 = ~new_n607 & ~new_n608;
  assign new_n610 = new_n604 & new_n609;
  assign new_n611 = ~new_n604 & ~new_n609;
  assign new_n612 = ~new_n610 & ~new_n611;
  assign new_n613 = ~new_n575 & ~new_n579;
  assign new_n614 = ~new_n577 & ~new_n613;
  assign new_n615_1 = ~new_n612 & ~new_n614;
  assign new_n616 = new_n612 & new_n614;
  assign new_n617 = ~new_n615_1 & ~new_n616;
  assign new_n618 = new_n603 & new_n617;
  assign new_n619 = ~new_n603 & ~new_n617;
  assign new_n620 = ~new_n618 & ~new_n619;
  assign new_n621 = ~new_n573 & ~new_n583;
  assign new_n622 = ~new_n572 & ~new_n621;
  assign new_n623 = ~new_n620 & ~new_n622;
  assign new_n624 = new_n620 & new_n622;
  assign new_n625 = ~new_n623 & ~new_n624;
  assign new_n626 = ~new_n598 & ~new_n625;
  assign new_n627 = new_n598 & new_n625;
  assign new_n628 = ~new_n626 & ~new_n627;
  assign new_n629 = new_n596 & new_n628;
  assign new_n630 = ~new_n596 & ~new_n628;
  assign new_n631 = ~new_n629 & ~new_n630;
  assign new_n632 = new_n595 & new_n631;
  assign new_n633 = ~new_n595 & ~new_n631;
  assign new_n634 = ~new_n632 & ~new_n633;
  assign new_n635 = ~new_n567 & new_n594;
  assign new_n636 = ~new_n595 & ~new_n635;
  assign new_n637 = ~new_n547 & new_n566;
  assign new_n638 = ~new_n567 & ~new_n637;
  assign new_n639 = n7965 & n10848;
  assign new_n640 = n7388 & n8028;
  assign new_n641 = new_n639 & new_n640;
  assign new_n642 = n8028 & n11892;
  assign new_n643 = n7388 & n10848;
  assign new_n644 = n1980 & n7965;
  assign new_n645 = ~new_n643 & ~new_n644;
  assign new_n646 = new_n643 & new_n644;
  assign new_n647 = ~new_n645 & ~new_n646;
  assign new_n648 = new_n642 & ~new_n647;
  assign new_n649 = ~new_n642 & new_n647;
  assign new_n650 = ~new_n648 & ~new_n649;
  assign new_n651 = new_n641 & ~new_n650;
  assign new_n652 = n7294 & n7965;
  assign new_n653 = new_n642 & ~new_n645;
  assign new_n654 = ~new_n646 & ~new_n653;
  assign new_n655 = ~new_n652 & new_n654;
  assign new_n656 = new_n652 & ~new_n654;
  assign new_n657 = ~new_n655 & ~new_n656;
  assign new_n658_1 = n2393 & n8028;
  assign new_n659 = n1980 & n7388;
  assign new_n660 = n10848 & n11892;
  assign new_n661 = ~new_n659 & ~new_n660;
  assign new_n662 = new_n659 & new_n660;
  assign new_n663 = ~new_n661 & ~new_n662;
  assign new_n664 = new_n658_1 & ~new_n663;
  assign new_n665 = ~new_n658_1 & new_n663;
  assign new_n666 = ~new_n664 & ~new_n665;
  assign new_n667 = ~new_n657 & new_n666;
  assign new_n668 = new_n657 & ~new_n666;
  assign new_n669 = ~new_n667 & ~new_n668;
  assign new_n670 = new_n651 & new_n669;
  assign new_n671_1 = ~new_n651 & ~new_n669;
  assign new_n672 = ~new_n670 & ~new_n671_1;
  assign new_n673 = ~new_n638 & ~new_n672;
  assign new_n674 = new_n638 & new_n672;
  assign new_n675 = ~new_n641 & new_n650;
  assign new_n676 = ~new_n651 & ~new_n675;
  assign new_n677 = ~new_n543 & new_n549;
  assign new_n678 = ~new_n546 & ~new_n677;
  assign new_n679 = ~new_n542 & new_n677;
  assign new_n680 = ~new_n678 & ~new_n679;
  assign new_n681 = ~new_n676 & ~new_n680;
  assign new_n682 = new_n676 & new_n680;
  assign new_n683 = n7965 & n8028;
  assign new_n684 = new_n543 & new_n683;
  assign new_n685 = ~new_n537 & ~new_n538;
  assign new_n686 = ~new_n539 & ~new_n685;
  assign new_n687 = new_n684 & new_n686;
  assign new_n688 = ~new_n684 & ~new_n686;
  assign new_n689 = ~new_n639 & ~new_n640;
  assign new_n690 = ~new_n641 & ~new_n689;
  assign new_n691 = ~new_n688 & new_n690;
  assign new_n692 = ~new_n687 & ~new_n691;
  assign new_n693 = ~new_n682 & new_n692;
  assign new_n694 = ~new_n681 & ~new_n693;
  assign new_n695 = ~new_n674 & ~new_n694;
  assign new_n696 = ~new_n673 & ~new_n695;
  assign new_n697 = new_n636 & new_n696;
  assign new_n698 = ~new_n636 & ~new_n696;
  assign new_n699 = n7965 & n12704;
  assign new_n700 = n7294 & n7388;
  assign new_n701 = new_n658_1 & ~new_n661;
  assign new_n702 = ~new_n662 & ~new_n701;
  assign new_n703 = new_n700 & ~new_n702;
  assign new_n704 = ~new_n700 & new_n702;
  assign new_n705 = ~new_n703 & ~new_n704;
  assign new_n706 = n5860 & n8028;
  assign new_n707 = n1980 & n11892;
  assign new_n708 = n2393 & n10848;
  assign new_n709 = ~new_n707 & ~new_n708;
  assign new_n710 = new_n707 & new_n708;
  assign new_n711 = ~new_n709 & ~new_n710;
  assign new_n712 = new_n706 & ~new_n711;
  assign new_n713 = ~new_n706 & new_n711;
  assign new_n714 = ~new_n712 & ~new_n713;
  assign new_n715 = ~new_n705 & ~new_n714;
  assign new_n716 = new_n705 & new_n714;
  assign new_n717 = ~new_n715 & ~new_n716;
  assign new_n718 = new_n699 & ~new_n717;
  assign new_n719 = ~new_n699 & new_n717;
  assign new_n720 = ~new_n718 & ~new_n719;
  assign new_n721 = ~new_n655 & ~new_n666;
  assign new_n722 = ~new_n656 & ~new_n721;
  assign new_n723 = ~new_n720 & ~new_n722;
  assign new_n724 = new_n720 & new_n722;
  assign new_n725 = ~new_n723 & ~new_n724;
  assign new_n726 = ~new_n670 & new_n725;
  assign new_n727 = new_n670 & ~new_n725;
  assign new_n728 = ~new_n726 & ~new_n727;
  assign new_n729 = ~new_n698 & new_n728;
  assign new_n730 = ~new_n697 & ~new_n729;
  assign new_n731 = new_n634 & ~new_n730;
  assign new_n732 = ~new_n634 & new_n730;
  assign new_n733 = ~new_n731 & ~new_n732;
  assign new_n734 = n5814 & n7965;
  assign new_n735 = ~new_n718 & new_n722;
  assign new_n736 = ~new_n719 & ~new_n735;
  assign new_n737 = n7388 & n12704;
  assign new_n738 = n7294 & n11892;
  assign new_n739 = ~new_n737 & ~new_n738;
  assign new_n740 = new_n737 & new_n738;
  assign new_n741 = ~new_n739 & ~new_n740;
  assign new_n742 = n1980 & n2393;
  assign new_n743 = n3986 & n8028;
  assign new_n744 = n5860 & n10848;
  assign new_n745 = ~new_n743 & ~new_n744;
  assign new_n746 = new_n743 & new_n744;
  assign new_n747 = ~new_n745 & ~new_n746;
  assign new_n748 = new_n742 & new_n747;
  assign new_n749 = ~new_n742 & ~new_n747;
  assign new_n750 = ~new_n748 & ~new_n749;
  assign new_n751 = ~new_n706 & ~new_n710;
  assign new_n752 = ~new_n709 & ~new_n751;
  assign new_n753_1 = ~new_n750 & new_n752;
  assign new_n754 = new_n750 & ~new_n752;
  assign new_n755 = ~new_n753_1 & ~new_n754;
  assign new_n756 = new_n741 & ~new_n755;
  assign new_n757 = ~new_n741 & new_n755;
  assign new_n758 = ~new_n756 & ~new_n757;
  assign new_n759 = ~new_n703 & new_n714;
  assign new_n760 = ~new_n704 & ~new_n759;
  assign new_n761 = ~new_n758 & new_n760;
  assign new_n762 = new_n758 & ~new_n760;
  assign new_n763 = ~new_n761 & ~new_n762;
  assign new_n764 = new_n736 & ~new_n763;
  assign new_n765 = ~new_n736 & new_n763;
  assign new_n766 = ~new_n764 & ~new_n765;
  assign new_n767 = new_n734 & new_n766;
  assign new_n768 = ~new_n734 & ~new_n766;
  assign new_n769 = ~new_n767 & ~new_n768;
  assign new_n770 = new_n727 & new_n769;
  assign new_n771 = ~new_n727 & ~new_n769;
  assign new_n772 = ~new_n770 & ~new_n771;
  assign new_n773 = ~new_n733 & new_n772;
  assign new_n774 = new_n733 & ~new_n772;
  assign new_n775 = ~new_n773 & ~new_n774;
  assign new_n776 = n7354 & n12299;
  assign new_n777 = n1209 & n8759;
  assign new_n778 = ~new_n776 & ~new_n777;
  assign new_n779 = n7354 & n8759;
  assign new_n780 = n1209 & n12299;
  assign new_n781 = new_n779 & new_n780;
  assign new_n782 = ~new_n778 & ~new_n781;
  assign new_n783_1 = n6776 & n7354;
  assign new_n784 = n7500 & n8759;
  assign new_n785 = new_n783_1 & new_n784;
  assign new_n786 = ~new_n782 & new_n785;
  assign new_n787 = n5105 & n8759;
  assign new_n788 = n6776 & n7500;
  assign new_n789 = ~new_n778 & new_n788;
  assign new_n790 = ~new_n781 & ~new_n789;
  assign new_n791 = new_n787 & ~new_n790;
  assign new_n792 = ~new_n787 & new_n790;
  assign new_n793 = ~new_n791 & ~new_n792;
  assign new_n794 = n7500 & n12299;
  assign new_n795 = n7354 & n7436;
  assign new_n796 = n1209 & n6776;
  assign new_n797 = ~new_n795 & ~new_n796;
  assign new_n798 = new_n795 & new_n796;
  assign new_n799 = ~new_n797 & ~new_n798;
  assign new_n800 = new_n794 & ~new_n799;
  assign new_n801 = ~new_n794 & new_n799;
  assign new_n802 = ~new_n800 & ~new_n801;
  assign new_n803 = new_n793 & new_n802;
  assign new_n804 = ~new_n793 & ~new_n802;
  assign new_n805 = ~new_n803 & ~new_n804;
  assign new_n806_1 = new_n786 & ~new_n805;
  assign new_n807 = n4141 & n8759;
  assign new_n808 = n5105 & n6776;
  assign new_n809 = new_n794 & ~new_n797;
  assign new_n810 = ~new_n798 & ~new_n809;
  assign new_n811 = new_n808 & ~new_n810;
  assign new_n812 = ~new_n808 & new_n810;
  assign new_n813 = ~new_n811 & ~new_n812;
  assign new_n814 = n7436 & n7500;
  assign new_n815 = n7354 & n8276;
  assign new_n816 = ~new_n780 & ~new_n815;
  assign new_n817 = new_n780 & new_n815;
  assign new_n818 = ~new_n816 & ~new_n817;
  assign new_n819 = new_n814 & ~new_n818;
  assign new_n820 = ~new_n814 & new_n818;
  assign new_n821 = ~new_n819 & ~new_n820;
  assign new_n822 = ~new_n813 & ~new_n821;
  assign new_n823 = new_n813 & new_n821;
  assign new_n824 = ~new_n822 & ~new_n823;
  assign new_n825 = new_n807 & ~new_n824;
  assign new_n826 = ~new_n807 & new_n824;
  assign new_n827 = ~new_n825 & ~new_n826;
  assign new_n828 = ~new_n792 & ~new_n802;
  assign new_n829 = ~new_n791 & ~new_n828;
  assign new_n830 = ~new_n827 & ~new_n829;
  assign new_n831 = new_n827 & new_n829;
  assign new_n832 = ~new_n830 & ~new_n831;
  assign new_n833 = new_n806_1 & ~new_n832;
  assign new_n834 = n4928 & n8759;
  assign new_n835 = ~new_n826 & ~new_n829;
  assign new_n836 = ~new_n825 & ~new_n835;
  assign new_n837_1 = n4141 & n6776;
  assign new_n838 = n5105 & n12299;
  assign new_n839 = ~new_n837_1 & ~new_n838;
  assign new_n840 = new_n837_1 & new_n838;
  assign new_n841 = ~new_n839 & ~new_n840;
  assign new_n842 = n1209 & n7436;
  assign new_n843 = n7500 & n8276;
  assign new_n844_1 = n7354 & n9241;
  assign new_n845 = ~new_n843 & ~new_n844_1;
  assign new_n846 = new_n843 & new_n844_1;
  assign new_n847 = ~new_n845 & ~new_n846;
  assign new_n848 = new_n842 & new_n847;
  assign new_n849 = ~new_n842 & ~new_n847;
  assign new_n850 = ~new_n848 & ~new_n849;
  assign new_n851 = new_n814 & ~new_n816;
  assign new_n852 = ~new_n817 & ~new_n851;
  assign new_n853 = ~new_n850 & ~new_n852;
  assign new_n854 = new_n850 & new_n852;
  assign new_n855 = ~new_n853 & ~new_n854;
  assign new_n856 = new_n841 & ~new_n855;
  assign new_n857 = ~new_n841 & new_n855;
  assign new_n858 = ~new_n856 & ~new_n857;
  assign new_n859 = ~new_n812 & ~new_n821;
  assign new_n860 = ~new_n811 & ~new_n859;
  assign new_n861 = new_n858 & new_n860;
  assign new_n862 = ~new_n858 & ~new_n860;
  assign new_n863 = ~new_n861 & ~new_n862;
  assign new_n864 = ~new_n836 & ~new_n863;
  assign new_n865 = new_n836 & new_n863;
  assign new_n866 = ~new_n864 & ~new_n865;
  assign new_n867 = new_n834 & new_n866;
  assign new_n868 = ~new_n834 & ~new_n866;
  assign new_n869 = ~new_n867 & ~new_n868;
  assign new_n870 = new_n833 & new_n869;
  assign new_n871 = ~new_n833 & ~new_n869;
  assign new_n872 = ~new_n870 & ~new_n871;
  assign new_n873 = ~new_n806_1 & new_n832;
  assign new_n874 = ~new_n833 & ~new_n873;
  assign new_n875 = ~new_n786 & new_n805;
  assign new_n876 = ~new_n806_1 & ~new_n875;
  assign new_n877 = ~new_n543 & ~new_n683;
  assign new_n878 = ~new_n684 & ~new_n877;
  assign new_n879 = new_n779 & new_n878;
  assign new_n880 = ~new_n783_1 & ~new_n784;
  assign new_n881 = ~new_n785 & ~new_n880;
  assign new_n882 = new_n879 & new_n881;
  assign new_n883 = ~new_n879 & ~new_n881;
  assign new_n884 = ~new_n687 & ~new_n688;
  assign new_n885 = new_n690 & ~new_n884;
  assign new_n886 = ~new_n690 & new_n884;
  assign new_n887 = ~new_n885 & ~new_n886;
  assign new_n888 = ~new_n883 & ~new_n887;
  assign new_n889 = ~new_n882 & ~new_n888;
  assign new_n890 = ~new_n779 & new_n788;
  assign new_n891 = ~new_n778 & new_n890;
  assign new_n892 = ~new_n782 & ~new_n890;
  assign new_n893 = ~new_n891 & ~new_n892;
  assign new_n894 = new_n889 & ~new_n893;
  assign new_n895 = ~new_n889 & new_n893;
  assign new_n896 = ~new_n681 & ~new_n682;
  assign new_n897 = new_n692 & ~new_n896;
  assign new_n898 = ~new_n692 & new_n896;
  assign new_n899 = ~new_n897 & ~new_n898;
  assign new_n900 = ~new_n895 & ~new_n899;
  assign new_n901 = ~new_n894 & ~new_n900;
  assign new_n902 = ~new_n876 & ~new_n901;
  assign new_n903 = new_n876 & new_n901;
  assign new_n904 = ~new_n673 & ~new_n674;
  assign new_n905 = new_n694 & ~new_n904;
  assign new_n906 = ~new_n673 & new_n695;
  assign new_n907 = ~new_n905 & ~new_n906;
  assign new_n908 = ~new_n903 & new_n907;
  assign new_n909 = ~new_n902 & ~new_n908;
  assign new_n910 = new_n874 & new_n909;
  assign new_n911_1 = ~new_n874 & ~new_n909;
  assign new_n912 = ~new_n697 & ~new_n698;
  assign new_n913 = new_n728 & new_n912;
  assign new_n914 = ~new_n728 & ~new_n912;
  assign new_n915 = ~new_n913 & ~new_n914;
  assign new_n916 = ~new_n911_1 & new_n915;
  assign new_n917 = ~new_n910 & ~new_n916;
  assign new_n918 = ~new_n872 & new_n917;
  assign new_n919 = new_n872 & ~new_n917;
  assign new_n920 = ~new_n918 & ~new_n919;
  assign new_n921 = ~new_n775 & ~new_n920;
  assign new_n922 = new_n775 & new_n920;
  assign new_n923 = ~new_n921 & ~new_n922;
  assign new_n924 = new_n536 & ~new_n923;
  assign new_n925 = ~new_n536 & new_n923;
  assign new_n926 = ~new_n480 & ~new_n484;
  assign new_n927 = ~new_n485 & ~new_n926;
  assign new_n928 = ~new_n910 & ~new_n911_1;
  assign new_n929 = ~new_n915 & new_n928;
  assign new_n930 = new_n915 & ~new_n928;
  assign new_n931 = ~new_n929 & ~new_n930;
  assign new_n932 = ~new_n927 & new_n931;
  assign new_n933 = new_n927 & ~new_n931;
  assign new_n934 = ~new_n475 & new_n479;
  assign new_n935 = ~new_n480 & ~new_n934;
  assign new_n936 = ~new_n902 & ~new_n903;
  assign new_n937 = new_n907 & ~new_n936;
  assign new_n938 = ~new_n907 & new_n936;
  assign new_n939 = ~new_n937 & ~new_n938;
  assign new_n940 = ~new_n935 & ~new_n939;
  assign new_n941 = new_n935 & new_n939;
  assign new_n942 = ~new_n470 & ~new_n474;
  assign new_n943 = ~new_n475 & ~new_n942;
  assign new_n944 = ~new_n894 & ~new_n895;
  assign new_n945 = ~new_n899 & ~new_n944;
  assign new_n946 = new_n899 & new_n944;
  assign new_n947 = ~new_n945 & ~new_n946;
  assign new_n948 = new_n943 & new_n947;
  assign new_n949 = ~new_n943 & ~new_n947;
  assign new_n950 = n5305 & n6038;
  assign new_n951 = ~new_n779 & ~new_n878;
  assign new_n952 = ~new_n879 & ~new_n951;
  assign new_n953 = new_n950 & new_n952;
  assign new_n954 = ~new_n468 & ~new_n469;
  assign new_n955 = ~new_n470 & ~new_n954;
  assign new_n956 = new_n953 & new_n955;
  assign new_n957 = ~new_n953 & ~new_n955;
  assign new_n958 = ~new_n882 & ~new_n883;
  assign new_n959 = ~new_n887 & new_n958;
  assign new_n960 = new_n887 & ~new_n958;
  assign new_n961 = ~new_n959 & ~new_n960;
  assign new_n962 = ~new_n957 & new_n961;
  assign new_n963 = ~new_n956 & ~new_n962;
  assign new_n964 = ~new_n949 & ~new_n963;
  assign new_n965 = ~new_n948 & ~new_n964;
  assign new_n966 = ~new_n941 & new_n965;
  assign new_n967 = ~new_n940 & ~new_n966;
  assign new_n968 = ~new_n933 & ~new_n967;
  assign new_n969 = ~new_n932 & ~new_n968;
  assign new_n970 = ~new_n925 & new_n969;
  assign new_n971 = ~new_n924 & ~new_n970;
  assign new_n972 = ~new_n534 & new_n971;
  assign new_n973 = new_n534 & ~new_n971;
  assign new_n974 = ~new_n972 & ~new_n973;
  assign new_n975 = ~new_n857 & ~new_n860;
  assign new_n976 = ~new_n840 & ~new_n975;
  assign new_n977 = ~new_n856 & new_n976;
  assign new_n978 = new_n840 & new_n975;
  assign new_n979 = ~new_n977 & ~new_n978;
  assign new_n980 = n4928 & n6776;
  assign new_n981 = n4141 & n12299;
  assign new_n982 = n8236 & n8759;
  assign new_n983 = ~new_n981 & ~new_n982;
  assign new_n984 = new_n981 & new_n982;
  assign new_n985 = ~new_n983 & ~new_n984;
  assign new_n986 = ~new_n980 & ~new_n985;
  assign new_n987 = new_n980 & new_n985;
  assign new_n988 = ~new_n986 & ~new_n987;
  assign new_n989 = ~new_n848 & new_n852;
  assign new_n990 = ~new_n849 & ~new_n989;
  assign new_n991 = ~new_n988 & ~new_n990;
  assign new_n992_1 = n5105 & n7436;
  assign new_n993 = new_n846 & new_n992_1;
  assign new_n994 = ~new_n846 & ~new_n992_1;
  assign new_n995 = ~new_n993 & ~new_n994;
  assign new_n996_1 = n7354 & n10510;
  assign new_n997 = n1209 & n8276;
  assign new_n998 = n7500 & n9241;
  assign new_n999 = ~new_n997 & ~new_n998;
  assign new_n1000 = new_n997 & new_n998;
  assign new_n1001 = ~new_n999 & ~new_n1000;
  assign new_n1002 = new_n996_1 & ~new_n1001;
  assign new_n1003 = ~new_n996_1 & new_n1001;
  assign new_n1004 = ~new_n1002 & ~new_n1003;
  assign new_n1005 = new_n995 & new_n1004;
  assign new_n1006 = ~new_n995 & ~new_n1004;
  assign new_n1007 = ~new_n1005 & ~new_n1006;
  assign new_n1008 = new_n991 & new_n1007;
  assign new_n1009 = new_n988 & new_n990;
  assign new_n1010 = new_n1007 & ~new_n1009;
  assign new_n1011 = ~new_n991 & ~new_n1010;
  assign new_n1012 = ~new_n1008 & ~new_n1011;
  assign new_n1013 = ~new_n1007 & new_n1009;
  assign new_n1014 = ~new_n1012 & ~new_n1013;
  assign new_n1015 = ~new_n979 & new_n1014;
  assign new_n1016 = new_n979 & ~new_n1014;
  assign new_n1017 = ~new_n1015 & ~new_n1016;
  assign new_n1018 = ~new_n864 & ~new_n1017;
  assign new_n1019 = new_n864 & new_n1017;
  assign new_n1020_1 = ~new_n1018 & ~new_n1019;
  assign new_n1021 = ~new_n867 & ~new_n870;
  assign new_n1022 = ~new_n1020_1 & new_n1021;
  assign new_n1023 = new_n1020_1 & ~new_n1021;
  assign new_n1024 = ~new_n1022 & ~new_n1023;
  assign new_n1025 = ~new_n619 & ~new_n622;
  assign new_n1026 = ~new_n602 & ~new_n1025;
  assign new_n1027 = ~new_n618 & new_n1026;
  assign new_n1028 = new_n602 & new_n1025;
  assign new_n1029 = ~new_n1027 & ~new_n1028;
  assign new_n1030 = n5069 & n8476;
  assign new_n1031 = n2530 & n6806;
  assign new_n1032 = n5331 & n12044;
  assign new_n1033 = ~new_n1031 & ~new_n1032;
  assign new_n1034 = new_n1031 & new_n1032;
  assign new_n1035 = ~new_n1033 & ~new_n1034;
  assign new_n1036 = ~new_n1030 & ~new_n1035;
  assign new_n1037 = new_n1030 & new_n1035;
  assign new_n1038 = ~new_n1036 & ~new_n1037;
  assign new_n1039 = ~new_n611 & new_n614;
  assign new_n1040 = ~new_n610 & ~new_n1039;
  assign new_n1041 = new_n1038 & ~new_n1040;
  assign new_n1042 = ~new_n1038 & new_n1040;
  assign new_n1043 = ~new_n1041 & ~new_n1042;
  assign new_n1044 = n2802 & n12648;
  assign new_n1045 = ~new_n608 & ~new_n1044;
  assign new_n1046 = new_n608 & new_n1044;
  assign new_n1047 = ~new_n1045 & ~new_n1046;
  assign new_n1048 = n1512 & n7690;
  assign new_n1049 = n1564 & n3616;
  assign new_n1050 = ~new_n578 & ~new_n1049;
  assign new_n1051 = new_n578 & new_n1049;
  assign new_n1052 = ~new_n1050 & ~new_n1051;
  assign new_n1053 = ~new_n1048 & ~new_n1052;
  assign new_n1054 = new_n1048 & new_n1052;
  assign new_n1055 = ~new_n1053 & ~new_n1054;
  assign new_n1056 = new_n1047 & ~new_n1055;
  assign new_n1057 = ~new_n1047 & new_n1055;
  assign new_n1058 = ~new_n1056 & ~new_n1057;
  assign new_n1059 = ~new_n1043 & ~new_n1058;
  assign new_n1060 = new_n1043 & new_n1058;
  assign new_n1061 = ~new_n1059 & ~new_n1060;
  assign new_n1062 = ~new_n1029 & new_n1061;
  assign new_n1063 = new_n1029 & ~new_n1061;
  assign new_n1064 = ~new_n1062 & ~new_n1063;
  assign new_n1065 = ~new_n626 & ~new_n1064;
  assign new_n1066 = new_n626 & new_n1064;
  assign new_n1067_1 = ~new_n1065 & ~new_n1066;
  assign new_n1068 = ~new_n629 & ~new_n632;
  assign new_n1069 = ~new_n1067_1 & new_n1068;
  assign new_n1070 = new_n1067_1 & ~new_n1068;
  assign new_n1071 = ~new_n1069 & ~new_n1070;
  assign new_n1072 = ~new_n757 & new_n760;
  assign new_n1073 = ~new_n740 & ~new_n1072;
  assign new_n1074 = ~new_n756 & new_n1073;
  assign new_n1075 = new_n740 & new_n1072;
  assign new_n1076 = ~new_n1074 & ~new_n1075;
  assign new_n1077 = n5814 & n7388;
  assign new_n1078 = n11892 & n12704;
  assign new_n1079 = n4903 & n7965;
  assign new_n1080 = ~new_n1078 & ~new_n1079;
  assign new_n1081 = new_n1078 & new_n1079;
  assign new_n1082 = ~new_n1080 & ~new_n1081;
  assign new_n1083 = ~new_n1077 & ~new_n1082;
  assign new_n1084 = new_n1077 & new_n1082;
  assign new_n1085 = ~new_n1083 & ~new_n1084;
  assign new_n1086 = ~new_n748 & ~new_n752;
  assign new_n1087 = ~new_n749 & ~new_n1086;
  assign new_n1088 = ~new_n1085 & ~new_n1087;
  assign new_n1089 = n2393 & n7294;
  assign new_n1090 = ~new_n746 & ~new_n1089;
  assign new_n1091 = new_n746 & new_n1089;
  assign new_n1092 = ~new_n1090 & ~new_n1091;
  assign new_n1093 = n3986 & n10848;
  assign new_n1094_1 = n5857 & n8028;
  assign new_n1095 = n1980 & n5860;
  assign new_n1096 = ~new_n1094_1 & ~new_n1095;
  assign new_n1097_1 = new_n1094_1 & new_n1095;
  assign new_n1098 = ~new_n1096 & ~new_n1097_1;
  assign new_n1099 = ~new_n1093 & ~new_n1098;
  assign new_n1100 = new_n1093 & new_n1098;
  assign new_n1101 = ~new_n1099 & ~new_n1100;
  assign new_n1102 = ~new_n1092 & new_n1101;
  assign new_n1103 = ~new_n1091 & ~new_n1101;
  assign new_n1104 = ~new_n1090 & new_n1103;
  assign new_n1105 = ~new_n1102 & ~new_n1104;
  assign new_n1106 = new_n1088 & new_n1105;
  assign new_n1107 = new_n1085 & new_n1087;
  assign new_n1108 = ~new_n1105 & new_n1107;
  assign new_n1109 = ~new_n1088 & ~new_n1105;
  assign new_n1110 = ~new_n1107 & ~new_n1109;
  assign new_n1111 = ~new_n1108 & ~new_n1110;
  assign new_n1112 = ~new_n1106 & ~new_n1111;
  assign new_n1113 = new_n1076 & ~new_n1112;
  assign new_n1114 = ~new_n1076 & new_n1112;
  assign new_n1115 = ~new_n1113 & ~new_n1114;
  assign new_n1116 = ~new_n764 & new_n1115;
  assign new_n1117 = new_n764 & ~new_n1115;
  assign new_n1118 = ~new_n1116 & ~new_n1117;
  assign new_n1119 = ~new_n767 & ~new_n770;
  assign new_n1120 = ~new_n1118 & new_n1119;
  assign new_n1121 = new_n1118 & ~new_n1119;
  assign new_n1122 = ~new_n1120 & ~new_n1121;
  assign new_n1123 = new_n1071 & new_n1122;
  assign new_n1124 = ~new_n1071 & ~new_n1122;
  assign new_n1125 = ~new_n1123 & ~new_n1124;
  assign new_n1126 = ~new_n732 & new_n772;
  assign new_n1127 = ~new_n731 & ~new_n1126;
  assign new_n1128 = new_n1125 & new_n1127;
  assign new_n1129 = ~new_n1125 & ~new_n1127;
  assign new_n1130 = ~new_n1128 & ~new_n1129;
  assign new_n1131 = ~new_n1024 & new_n1130;
  assign new_n1132 = new_n1024 & ~new_n1130;
  assign new_n1133 = ~new_n1131 & ~new_n1132;
  assign new_n1134 = ~new_n775 & ~new_n918;
  assign new_n1135 = ~new_n919 & ~new_n1134;
  assign new_n1136_1 = new_n1133 & new_n1135;
  assign new_n1137 = ~new_n1133 & ~new_n1135;
  assign new_n1138_1 = ~new_n1136_1 & ~new_n1137;
  assign new_n1139 = new_n974 & ~new_n1138_1;
  assign new_n1140 = ~new_n974 & new_n1138_1;
  assign n226 = ~new_n1139 & ~new_n1140;
  assign new_n1142 = n2879 & n5305;
  assign new_n1143 = n5964 & n7265;
  assign new_n1144 = new_n1142 & new_n1143;
  assign new_n1145 = n1097 & n7265;
  assign new_n1146 = n2879 & n5964;
  assign new_n1147 = n5305 & n10223;
  assign new_n1148 = ~new_n1146 & ~new_n1147;
  assign new_n1149 = new_n1146 & new_n1147;
  assign new_n1150 = ~new_n1148 & ~new_n1149;
  assign new_n1151 = new_n1145 & ~new_n1150;
  assign new_n1152 = ~new_n1145 & new_n1150;
  assign new_n1153 = ~new_n1151 & ~new_n1152;
  assign new_n1154 = new_n1144 & ~new_n1153;
  assign new_n1155 = n4634 & n5305;
  assign new_n1156 = new_n1145 & ~new_n1148;
  assign new_n1157 = ~new_n1149 & ~new_n1156;
  assign new_n1158 = ~new_n1155 & new_n1157;
  assign new_n1159 = new_n1155 & ~new_n1157;
  assign new_n1160 = ~new_n1158 & ~new_n1159;
  assign new_n1161 = n4312 & n7265;
  assign new_n1162 = n5964 & n10223;
  assign new_n1163 = n1097 & n2879;
  assign new_n1164 = ~new_n1162 & ~new_n1163;
  assign new_n1165 = new_n1162 & new_n1163;
  assign new_n1166 = ~new_n1164 & ~new_n1165;
  assign new_n1167 = new_n1161 & ~new_n1166;
  assign new_n1168 = ~new_n1161 & new_n1166;
  assign new_n1169 = ~new_n1167 & ~new_n1168;
  assign new_n1170 = ~new_n1160 & new_n1169;
  assign new_n1171 = new_n1160 & ~new_n1169;
  assign new_n1172 = ~new_n1170 & ~new_n1171;
  assign new_n1173 = new_n1154 & new_n1172;
  assign new_n1174 = ~new_n1154 & ~new_n1172;
  assign new_n1175 = ~new_n1173 & ~new_n1174;
  assign new_n1176 = ~new_n1144 & new_n1153;
  assign new_n1177 = ~new_n1154 & ~new_n1176;
  assign new_n1178 = n7946 & n12299;
  assign new_n1179 = n8759 & n9189;
  assign new_n1180 = ~new_n1178 & ~new_n1179;
  assign new_n1181 = n7946 & n8759;
  assign new_n1182 = n9189 & n12299;
  assign new_n1183 = new_n1181 & new_n1182;
  assign new_n1184 = ~new_n1180 & ~new_n1183;
  assign new_n1185 = n2024 & n6776;
  assign new_n1186 = ~new_n1181 & new_n1185;
  assign new_n1187 = ~new_n1184 & ~new_n1186;
  assign new_n1188 = ~new_n1180 & new_n1185;
  assign new_n1189 = ~new_n1181 & new_n1188;
  assign new_n1190 = ~new_n1187 & ~new_n1189;
  assign new_n1191 = n2558 & n5331;
  assign new_n1192 = n7965 & n9763;
  assign new_n1193 = new_n1191 & new_n1192;
  assign new_n1194 = ~new_n1191 & ~new_n1192;
  assign new_n1195 = ~new_n1193 & ~new_n1194;
  assign new_n1196 = new_n1181 & new_n1195;
  assign new_n1197 = n6776 & n7946;
  assign new_n1198_1 = n2024 & n8759;
  assign new_n1199_1 = ~new_n1197 & ~new_n1198_1;
  assign new_n1200 = new_n1197 & new_n1198_1;
  assign new_n1201 = ~new_n1199_1 & ~new_n1200;
  assign new_n1202 = new_n1196 & new_n1201;
  assign new_n1203 = ~new_n1196 & ~new_n1201;
  assign new_n1204 = n2498 & n5331;
  assign new_n1205 = n2558 & n8476;
  assign new_n1206 = ~new_n1204 & ~new_n1205;
  assign new_n1207 = new_n1204 & new_n1205;
  assign new_n1208 = ~new_n1206 & ~new_n1207;
  assign new_n1209_1 = n7965 & n9111;
  assign new_n1210 = n7388 & n9763;
  assign new_n1211 = ~new_n1209_1 & ~new_n1210;
  assign new_n1212 = new_n1209_1 & new_n1210;
  assign new_n1213 = ~new_n1211 & ~new_n1212;
  assign new_n1214 = new_n1193 & new_n1213;
  assign new_n1215 = ~new_n1193 & ~new_n1213;
  assign new_n1216 = ~new_n1214 & ~new_n1215;
  assign new_n1217 = new_n1208 & ~new_n1216;
  assign new_n1218 = ~new_n1208 & new_n1216;
  assign new_n1219 = ~new_n1217 & ~new_n1218;
  assign new_n1220 = ~new_n1203 & ~new_n1219;
  assign new_n1221 = ~new_n1202 & ~new_n1220;
  assign new_n1222 = new_n1190 & ~new_n1221;
  assign new_n1223 = ~new_n1190 & new_n1221;
  assign new_n1224 = ~new_n1222 & ~new_n1223;
  assign new_n1225 = n2530 & n2558;
  assign new_n1226 = n2498 & n8476;
  assign new_n1227 = n5331 & n5579;
  assign new_n1228 = ~new_n1226 & ~new_n1227;
  assign new_n1229 = new_n1226 & new_n1227;
  assign new_n1230 = ~new_n1228 & ~new_n1229;
  assign new_n1231 = new_n1225 & ~new_n1230;
  assign new_n1232 = ~new_n1225 & new_n1230;
  assign new_n1233 = ~new_n1231 & ~new_n1232;
  assign new_n1234 = ~new_n1207 & new_n1233;
  assign new_n1235 = new_n1207 & ~new_n1233;
  assign new_n1236 = ~new_n1234 & ~new_n1235;
  assign new_n1237 = n9763 & n11892;
  assign new_n1238 = n7388 & n9111;
  assign new_n1239 = n3342 & n7965;
  assign new_n1240 = ~new_n1238 & ~new_n1239;
  assign new_n1241 = new_n1238 & new_n1239;
  assign new_n1242 = ~new_n1240 & ~new_n1241;
  assign new_n1243 = new_n1237 & ~new_n1242;
  assign new_n1244 = ~new_n1237 & new_n1242;
  assign new_n1245 = ~new_n1243 & ~new_n1244;
  assign new_n1246 = new_n1212 & ~new_n1245;
  assign new_n1247 = ~new_n1212 & new_n1245;
  assign new_n1248 = ~new_n1246 & ~new_n1247;
  assign new_n1249 = ~new_n1208 & ~new_n1214;
  assign new_n1250 = ~new_n1215 & ~new_n1249;
  assign new_n1251 = new_n1248 & new_n1250;
  assign new_n1252 = ~new_n1248 & ~new_n1250;
  assign new_n1253 = ~new_n1251 & ~new_n1252;
  assign new_n1254 = ~new_n1236 & new_n1253;
  assign new_n1255 = new_n1236 & ~new_n1253;
  assign new_n1256 = ~new_n1254 & ~new_n1255;
  assign new_n1257 = ~new_n1224 & ~new_n1256;
  assign new_n1258 = new_n1224 & new_n1256;
  assign new_n1259 = ~new_n1257 & ~new_n1258;
  assign new_n1260 = new_n1177 & ~new_n1259;
  assign new_n1261 = ~new_n1177 & new_n1259;
  assign new_n1262 = n5305 & n7265;
  assign new_n1263 = ~new_n1181 & ~new_n1195;
  assign new_n1264 = ~new_n1196 & ~new_n1263;
  assign new_n1265 = new_n1262 & new_n1264;
  assign new_n1266 = ~new_n1142 & ~new_n1143;
  assign new_n1267 = ~new_n1144 & ~new_n1266;
  assign new_n1268 = new_n1265 & new_n1267;
  assign new_n1269_1 = ~new_n1265 & ~new_n1267;
  assign new_n1270 = ~new_n1202 & ~new_n1203;
  assign new_n1271 = new_n1219 & ~new_n1270;
  assign new_n1272 = ~new_n1219 & new_n1270;
  assign new_n1273 = ~new_n1271 & ~new_n1272;
  assign new_n1274 = ~new_n1269_1 & new_n1273;
  assign new_n1275 = ~new_n1268 & ~new_n1274;
  assign new_n1276 = ~new_n1261 & ~new_n1275;
  assign new_n1277 = ~new_n1260 & ~new_n1276;
  assign new_n1278 = new_n1175 & ~new_n1277;
  assign new_n1279 = ~new_n1175 & new_n1277;
  assign new_n1280 = ~new_n1278 & ~new_n1279;
  assign new_n1281 = ~new_n1184 & new_n1200;
  assign new_n1282 = n2522 & n8759;
  assign new_n1283 = ~new_n1183 & ~new_n1188;
  assign new_n1284 = new_n1282 & ~new_n1283;
  assign new_n1285 = ~new_n1282 & new_n1283;
  assign new_n1286 = ~new_n1284 & ~new_n1285;
  assign new_n1287 = n7436 & n7946;
  assign new_n1288 = n6776 & n9189;
  assign new_n1289 = n2024 & n12299;
  assign new_n1290 = ~new_n1288 & ~new_n1289;
  assign new_n1291 = new_n1288 & new_n1289;
  assign new_n1292 = ~new_n1290 & ~new_n1291;
  assign new_n1293 = new_n1287 & ~new_n1292;
  assign new_n1294 = ~new_n1287 & new_n1292;
  assign new_n1295 = ~new_n1293 & ~new_n1294;
  assign new_n1296 = ~new_n1286 & ~new_n1295;
  assign new_n1297 = new_n1286 & new_n1295;
  assign new_n1298 = ~new_n1296 & ~new_n1297;
  assign new_n1299 = ~new_n1281 & new_n1298;
  assign new_n1300 = new_n1281 & ~new_n1298;
  assign new_n1301 = ~new_n1299 & ~new_n1300;
  assign new_n1302 = ~new_n1222 & new_n1256;
  assign new_n1303 = ~new_n1223 & ~new_n1302;
  assign new_n1304 = new_n1301 & new_n1303;
  assign new_n1305 = ~new_n1301 & ~new_n1303;
  assign new_n1306 = ~new_n1304 & ~new_n1305;
  assign new_n1307 = n521 & n5331;
  assign new_n1308 = new_n1225 & ~new_n1228;
  assign new_n1309 = ~new_n1229 & ~new_n1308;
  assign new_n1310 = new_n1307 & ~new_n1309;
  assign new_n1311 = ~new_n1307 & new_n1309;
  assign new_n1312 = ~new_n1310 & ~new_n1311;
  assign new_n1313 = n2558 & n12648;
  assign new_n1314 = n5579 & n8476;
  assign new_n1315 = n2498 & n2530;
  assign new_n1316 = ~new_n1314 & ~new_n1315;
  assign new_n1317 = new_n1314 & new_n1315;
  assign new_n1318 = ~new_n1316 & ~new_n1317;
  assign new_n1319 = new_n1313 & ~new_n1318;
  assign new_n1320 = ~new_n1313 & new_n1318;
  assign new_n1321 = ~new_n1319 & ~new_n1320;
  assign new_n1322 = ~new_n1312 & ~new_n1321;
  assign new_n1323 = new_n1312 & new_n1321;
  assign new_n1324 = ~new_n1322 & ~new_n1323;
  assign new_n1325 = ~new_n1235 & new_n1324;
  assign new_n1326 = new_n1235 & ~new_n1324;
  assign new_n1327 = ~new_n1325 & ~new_n1326;
  assign new_n1328 = n806 & n7965;
  assign new_n1329 = new_n1237 & ~new_n1240;
  assign new_n1330 = ~new_n1241 & ~new_n1329;
  assign new_n1331 = new_n1328 & ~new_n1330;
  assign new_n1332 = ~new_n1328 & new_n1330;
  assign new_n1333_1 = ~new_n1331 & ~new_n1332;
  assign new_n1334 = n2393 & n9763;
  assign new_n1335 = n3342 & n7388;
  assign new_n1336 = n9111 & n11892;
  assign new_n1337 = ~new_n1335 & ~new_n1336;
  assign new_n1338 = new_n1335 & new_n1336;
  assign new_n1339 = ~new_n1337 & ~new_n1338;
  assign new_n1340 = new_n1334 & ~new_n1339;
  assign new_n1341 = ~new_n1334 & new_n1339;
  assign new_n1342 = ~new_n1340 & ~new_n1341;
  assign new_n1343 = ~new_n1333_1 & ~new_n1342;
  assign new_n1344 = new_n1333_1 & new_n1342;
  assign new_n1345 = ~new_n1343 & ~new_n1344;
  assign new_n1346 = new_n1246 & ~new_n1345;
  assign new_n1347 = ~new_n1246 & new_n1345;
  assign new_n1348 = ~new_n1346 & ~new_n1347;
  assign new_n1349 = ~new_n1327 & ~new_n1348;
  assign new_n1350 = new_n1236 & ~new_n1252;
  assign new_n1351 = ~new_n1251 & ~new_n1350;
  assign new_n1352 = new_n1349 & new_n1351;
  assign new_n1353_1 = new_n1327 & new_n1348;
  assign new_n1354 = ~new_n1351 & new_n1353_1;
  assign new_n1355 = ~new_n1349 & ~new_n1351;
  assign new_n1356 = ~new_n1353_1 & ~new_n1355;
  assign new_n1357_1 = ~new_n1354 & ~new_n1356;
  assign new_n1358 = ~new_n1352 & ~new_n1357_1;
  assign new_n1359 = ~new_n1306 & new_n1358;
  assign new_n1360 = new_n1306 & ~new_n1358;
  assign new_n1361 = ~new_n1359 & ~new_n1360;
  assign new_n1362 = new_n1280 & new_n1361;
  assign new_n1363 = ~new_n1280 & ~new_n1361;
  assign n381 = new_n1362 | new_n1363;
  assign new_n1365 = n6038 & n7862;
  assign new_n1366 = n6877 & n7354;
  assign new_n1367 = n1564 & n4805;
  assign new_n1368 = n7236 & n8028;
  assign new_n1369 = new_n1367 & new_n1368;
  assign new_n1370 = ~new_n1367 & ~new_n1368;
  assign new_n1371 = ~new_n1369 & ~new_n1370;
  assign new_n1372 = new_n1366 & new_n1371;
  assign new_n1373 = ~new_n1366 & ~new_n1371;
  assign new_n1374 = ~new_n1372 & ~new_n1373;
  assign new_n1375 = new_n1365 & new_n1374;
  assign new_n1376 = ~new_n1365 & ~new_n1374;
  assign n397 = ~new_n1375 & ~new_n1376;
  assign new_n1378 = n4189 & n11407;
  assign new_n1379 = n6687 & n11877;
  assign new_n1380 = ~new_n1378 & ~new_n1379;
  assign new_n1381 = n6687 & n11407;
  assign new_n1382 = n4189 & n11877;
  assign new_n1383 = new_n1381 & new_n1382;
  assign new_n1384 = ~new_n1380 & ~new_n1383;
  assign new_n1385 = n2564 & n11407;
  assign new_n1386 = n5212 & n6687;
  assign new_n1387 = new_n1385 & new_n1386;
  assign new_n1388 = ~new_n1384 & new_n1387;
  assign new_n1389 = n4370 & n6687;
  assign new_n1390 = n2564 & n5212;
  assign new_n1391 = ~new_n1383 & ~new_n1390;
  assign new_n1392 = ~new_n1380 & ~new_n1391;
  assign new_n1393 = new_n1389 & new_n1392;
  assign new_n1394 = ~new_n1389 & ~new_n1392;
  assign new_n1395 = ~new_n1393 & ~new_n1394;
  assign new_n1396 = n4189 & n5212;
  assign new_n1397 = n6770 & n11407;
  assign new_n1398 = n2564 & n11877;
  assign new_n1399 = ~new_n1397 & ~new_n1398;
  assign new_n1400 = new_n1397 & new_n1398;
  assign new_n1401 = ~new_n1399 & ~new_n1400;
  assign new_n1402 = new_n1396 & ~new_n1401;
  assign new_n1403 = ~new_n1396 & new_n1401;
  assign new_n1404 = ~new_n1402 & ~new_n1403;
  assign new_n1405 = ~new_n1395 & ~new_n1404;
  assign new_n1406 = new_n1395 & new_n1404;
  assign new_n1407 = ~new_n1405 & ~new_n1406;
  assign new_n1408 = new_n1388 & ~new_n1407;
  assign new_n1409 = ~new_n1388 & new_n1407;
  assign new_n1410 = ~new_n1408 & ~new_n1409;
  assign new_n1411 = n5314 & n10990;
  assign new_n1412 = n1478 & n11222;
  assign new_n1413 = ~new_n1411 & ~new_n1412;
  assign new_n1414 = new_n1411 & new_n1412;
  assign new_n1415 = ~new_n1413 & ~new_n1414;
  assign new_n1416 = n10990 & n11222;
  assign new_n1417 = n5760 & n11153;
  assign new_n1418 = ~new_n1416 & new_n1417;
  assign new_n1419 = ~new_n1415 & ~new_n1418;
  assign new_n1420 = ~new_n1413 & new_n1417;
  assign new_n1421 = ~new_n1416 & new_n1420;
  assign new_n1422 = ~new_n1419 & ~new_n1421;
  assign new_n1423 = n12069 & n12489;
  assign new_n1424 = n7159 & n12391;
  assign new_n1425 = ~new_n1423 & new_n1424;
  assign new_n1426 = n7891 & n12489;
  assign new_n1427 = n12069 & n12777;
  assign new_n1428 = ~new_n1426 & ~new_n1427;
  assign new_n1429 = n7891 & n12777;
  assign new_n1430 = new_n1423 & new_n1429;
  assign new_n1431 = ~new_n1428 & ~new_n1430;
  assign new_n1432 = ~new_n1425 & ~new_n1431;
  assign new_n1433 = new_n1425 & ~new_n1428;
  assign new_n1434 = ~new_n1432 & ~new_n1433;
  assign new_n1435 = new_n1422 & new_n1434;
  assign new_n1436 = ~new_n1422 & ~new_n1434;
  assign new_n1437 = ~new_n1435 & ~new_n1436;
  assign new_n1438 = new_n1416 & new_n1423;
  assign new_n1439 = n5760 & n11222;
  assign new_n1440 = n10990 & n11153;
  assign new_n1441 = ~new_n1439 & ~new_n1440;
  assign new_n1442 = new_n1439 & new_n1440;
  assign new_n1443 = ~new_n1441 & ~new_n1442;
  assign new_n1444 = new_n1438 & new_n1443;
  assign new_n1445 = ~new_n1438 & ~new_n1443;
  assign new_n1446 = n7159 & n12069;
  assign new_n1447 = n12391 & n12489;
  assign new_n1448 = ~new_n1446 & ~new_n1447;
  assign new_n1449 = new_n1446 & new_n1447;
  assign new_n1450 = ~new_n1448 & ~new_n1449;
  assign new_n1451 = ~new_n1445 & new_n1450;
  assign new_n1452 = ~new_n1444 & ~new_n1451;
  assign new_n1453 = new_n1437 & new_n1452;
  assign new_n1454 = ~new_n1437 & ~new_n1452;
  assign new_n1455 = ~new_n1453 & ~new_n1454;
  assign new_n1456 = n8336 & n11728;
  assign new_n1457 = n10928 & n12709;
  assign new_n1458 = new_n1456 & new_n1457;
  assign new_n1459 = n6986 & n12709;
  assign new_n1460 = n10928 & n11728;
  assign new_n1461 = n6429 & n8336;
  assign new_n1462 = ~new_n1460 & ~new_n1461;
  assign new_n1463 = new_n1460 & new_n1461;
  assign new_n1464 = ~new_n1462 & ~new_n1463;
  assign new_n1465 = new_n1459 & ~new_n1464;
  assign new_n1466 = ~new_n1459 & new_n1464;
  assign new_n1467 = ~new_n1465 & ~new_n1466;
  assign new_n1468 = new_n1458 & ~new_n1467;
  assign new_n1469 = ~new_n1458 & new_n1467;
  assign new_n1470 = ~new_n1468 & ~new_n1469;
  assign new_n1471_1 = n8336 & n12709;
  assign new_n1472 = ~new_n1416 & ~new_n1423;
  assign new_n1473 = ~new_n1438 & ~new_n1472;
  assign new_n1474 = new_n1471_1 & new_n1473;
  assign new_n1475 = ~new_n1456 & ~new_n1457;
  assign new_n1476 = ~new_n1458 & ~new_n1475;
  assign new_n1477 = new_n1474 & new_n1476;
  assign new_n1478_1 = ~new_n1474 & ~new_n1476;
  assign new_n1479 = ~new_n1444 & ~new_n1445;
  assign new_n1480 = new_n1450 & ~new_n1479;
  assign new_n1481 = ~new_n1450 & new_n1479;
  assign new_n1482 = ~new_n1480 & ~new_n1481;
  assign new_n1483 = ~new_n1478_1 & ~new_n1482;
  assign new_n1484 = ~new_n1477 & ~new_n1483;
  assign new_n1485 = ~new_n1470 & new_n1484;
  assign new_n1486 = new_n1470 & ~new_n1484;
  assign new_n1487 = ~new_n1485 & ~new_n1486;
  assign new_n1488 = new_n1455 & ~new_n1487;
  assign new_n1489 = ~new_n1455 & new_n1487;
  assign new_n1490 = ~new_n1488 & ~new_n1489;
  assign new_n1491 = ~new_n1381 & new_n1390;
  assign new_n1492 = new_n1384 & ~new_n1491;
  assign new_n1493 = ~new_n1384 & new_n1491;
  assign new_n1494 = ~new_n1492 & ~new_n1493;
  assign new_n1495 = new_n1490 & ~new_n1494;
  assign new_n1496 = ~new_n1490 & new_n1494;
  assign new_n1497 = ~new_n1471_1 & ~new_n1473;
  assign new_n1498 = ~new_n1474 & ~new_n1497;
  assign new_n1499 = new_n1381 & new_n1498;
  assign new_n1500 = ~new_n1385 & ~new_n1386;
  assign new_n1501 = ~new_n1387 & ~new_n1500;
  assign new_n1502 = new_n1499 & new_n1501;
  assign new_n1503 = ~new_n1499 & ~new_n1501;
  assign new_n1504 = ~new_n1477 & ~new_n1478_1;
  assign new_n1505 = ~new_n1482 & new_n1504;
  assign new_n1506 = new_n1482 & ~new_n1504;
  assign new_n1507 = ~new_n1505 & ~new_n1506;
  assign new_n1508 = ~new_n1503 & new_n1507;
  assign new_n1509 = ~new_n1502 & ~new_n1508;
  assign new_n1510_1 = ~new_n1496 & ~new_n1509;
  assign new_n1511 = ~new_n1495 & ~new_n1510_1;
  assign new_n1512_1 = new_n1410 & ~new_n1511;
  assign new_n1513 = ~new_n1410 & new_n1511;
  assign new_n1514 = ~new_n1512_1 & ~new_n1513;
  assign new_n1515 = n8336 & n8819;
  assign new_n1516 = n2226 & n12709;
  assign new_n1517 = n6429 & n10928;
  assign new_n1518 = n6986 & n11728;
  assign new_n1519 = ~new_n1517 & ~new_n1518;
  assign new_n1520 = new_n1517 & new_n1518;
  assign new_n1521 = ~new_n1519 & ~new_n1520;
  assign new_n1522 = new_n1516 & ~new_n1521;
  assign new_n1523_1 = ~new_n1516 & new_n1521;
  assign new_n1524 = ~new_n1522 & ~new_n1523_1;
  assign new_n1525 = new_n1515 & ~new_n1524;
  assign new_n1526 = ~new_n1515 & new_n1524;
  assign new_n1527 = ~new_n1525 & ~new_n1526;
  assign new_n1528 = new_n1459 & ~new_n1462;
  assign new_n1529 = ~new_n1463 & ~new_n1528;
  assign new_n1530 = ~new_n1527 & ~new_n1529;
  assign new_n1531 = new_n1527 & new_n1529;
  assign new_n1532 = ~new_n1530 & ~new_n1531;
  assign new_n1533 = ~new_n1468 & new_n1532;
  assign new_n1534 = new_n1468 & ~new_n1532;
  assign new_n1535 = ~new_n1533 & ~new_n1534;
  assign new_n1536 = ~new_n1431 & new_n1449;
  assign new_n1537 = n6254 & n12069;
  assign new_n1538 = ~new_n1424 & ~new_n1430;
  assign new_n1539 = ~new_n1428 & ~new_n1538;
  assign new_n1540 = new_n1537 & new_n1539;
  assign new_n1541 = ~new_n1537 & ~new_n1539;
  assign new_n1542 = ~new_n1540 & ~new_n1541;
  assign new_n1543 = n7160 & n12489;
  assign new_n1544 = n12391 & n12777;
  assign new_n1545 = n7159 & n7891;
  assign new_n1546 = ~new_n1544 & ~new_n1545;
  assign new_n1547 = new_n1544 & new_n1545;
  assign new_n1548 = ~new_n1546 & ~new_n1547;
  assign new_n1549 = new_n1543 & ~new_n1548;
  assign new_n1550 = ~new_n1543 & new_n1548;
  assign new_n1551 = ~new_n1549 & ~new_n1550;
  assign new_n1552 = ~new_n1542 & ~new_n1551;
  assign new_n1553 = new_n1542 & new_n1551;
  assign new_n1554 = ~new_n1552 & ~new_n1553;
  assign new_n1555 = ~new_n1536 & new_n1554;
  assign new_n1556 = new_n1536 & ~new_n1554;
  assign new_n1557 = ~new_n1555 & ~new_n1556;
  assign new_n1558 = ~new_n1415 & new_n1442;
  assign new_n1559 = n11222 & n11791;
  assign new_n1560 = ~new_n1414 & ~new_n1420;
  assign new_n1561 = new_n1559 & ~new_n1560;
  assign new_n1562 = ~new_n1559 & new_n1560;
  assign new_n1563 = ~new_n1561 & ~new_n1562;
  assign new_n1564_1 = n5314 & n5760;
  assign new_n1565 = n996 & n10990;
  assign new_n1566 = n1478 & n11153;
  assign new_n1567 = ~new_n1565 & ~new_n1566;
  assign new_n1568 = new_n1565 & new_n1566;
  assign new_n1569 = ~new_n1567 & ~new_n1568;
  assign new_n1570 = new_n1564_1 & ~new_n1569;
  assign new_n1571 = ~new_n1564_1 & new_n1569;
  assign new_n1572 = ~new_n1570 & ~new_n1571;
  assign new_n1573 = ~new_n1563 & ~new_n1572;
  assign new_n1574 = new_n1563 & new_n1572;
  assign new_n1575 = ~new_n1573 & ~new_n1574;
  assign new_n1576_1 = new_n1558 & ~new_n1575;
  assign new_n1577 = ~new_n1558 & new_n1575;
  assign new_n1578 = ~new_n1576_1 & ~new_n1577;
  assign new_n1579 = new_n1557 & new_n1578;
  assign new_n1580 = ~new_n1557 & ~new_n1578;
  assign new_n1581 = ~new_n1579 & ~new_n1580;
  assign new_n1582 = ~new_n1436 & ~new_n1452;
  assign new_n1583 = ~new_n1435 & ~new_n1582;
  assign new_n1584 = new_n1581 & new_n1583;
  assign new_n1585 = ~new_n1581 & ~new_n1583;
  assign new_n1586 = ~new_n1584 & ~new_n1585;
  assign new_n1587 = new_n1535 & ~new_n1586;
  assign new_n1588 = ~new_n1535 & new_n1586;
  assign new_n1589 = ~new_n1587 & ~new_n1588;
  assign new_n1590 = ~new_n1455 & ~new_n1485;
  assign new_n1591 = ~new_n1486 & ~new_n1590;
  assign new_n1592 = ~new_n1589 & ~new_n1591;
  assign new_n1593 = new_n1589 & new_n1591;
  assign new_n1594 = ~new_n1592 & ~new_n1593;
  assign new_n1595 = new_n1514 & ~new_n1594;
  assign new_n1596 = ~new_n1514 & new_n1594;
  assign n658 = ~new_n1595 & ~new_n1596;
  assign new_n1598 = n1333 & n2585;
  assign new_n1599 = n2508 & n3172;
  assign new_n1600 = ~new_n1598 & ~new_n1599;
  assign new_n1601 = new_n1598 & new_n1599;
  assign new_n1602 = ~new_n1600 & ~new_n1601;
  assign new_n1603 = n1333 & n2508;
  assign new_n1604 = n1333 & n12720;
  assign new_n1605 = n2509 & n3172;
  assign new_n1606 = new_n1604 & new_n1605;
  assign new_n1607 = ~new_n1604 & ~new_n1605;
  assign new_n1608 = n6038 & n11757;
  assign new_n1609 = ~new_n1607 & new_n1608;
  assign new_n1610 = ~new_n1606 & ~new_n1609;
  assign new_n1611 = ~new_n1603 & new_n1610;
  assign new_n1612 = new_n1603 & ~new_n1610;
  assign new_n1613 = n2509 & n11757;
  assign new_n1614 = n3172 & n12720;
  assign new_n1615 = n5240 & n6038;
  assign new_n1616 = ~new_n1614 & ~new_n1615;
  assign new_n1617 = n3172 & n6038;
  assign new_n1618 = n5240 & n12720;
  assign new_n1619 = new_n1617 & new_n1618;
  assign new_n1620 = ~new_n1616 & ~new_n1619;
  assign new_n1621 = ~new_n1613 & ~new_n1620;
  assign new_n1622 = new_n1613 & new_n1620;
  assign new_n1623 = ~new_n1621 & ~new_n1622;
  assign new_n1624 = ~new_n1612 & ~new_n1623;
  assign new_n1625 = ~new_n1611 & ~new_n1624;
  assign new_n1626 = ~new_n1602 & ~new_n1625;
  assign new_n1627 = new_n1602 & new_n1625;
  assign new_n1628 = ~new_n1626 & ~new_n1627;
  assign new_n1629 = n11757 & n12720;
  assign new_n1630 = n2509 & n5240;
  assign new_n1631 = n6038 & n11821;
  assign new_n1632 = ~new_n1630 & ~new_n1631;
  assign new_n1633 = new_n1630 & new_n1631;
  assign new_n1634 = ~new_n1632 & ~new_n1633;
  assign new_n1635 = ~new_n1629 & ~new_n1634;
  assign new_n1636 = new_n1629 & new_n1634;
  assign new_n1637 = ~new_n1635 & ~new_n1636;
  assign new_n1638 = new_n1613 & ~new_n1616;
  assign new_n1639 = ~new_n1619 & ~new_n1638;
  assign new_n1640 = ~new_n1637 & new_n1639;
  assign new_n1641 = new_n1637 & ~new_n1639;
  assign new_n1642 = ~new_n1640 & ~new_n1641;
  assign new_n1643 = ~new_n1628 & ~new_n1642;
  assign new_n1644 = new_n1628 & new_n1642;
  assign new_n1645 = ~new_n1643 & ~new_n1644;
  assign new_n1646 = n2585 & n7862;
  assign new_n1647 = ~new_n1611 & ~new_n1612;
  assign new_n1648 = new_n1623 & ~new_n1647;
  assign new_n1649 = ~new_n1623 & new_n1647;
  assign new_n1650 = ~new_n1648 & ~new_n1649;
  assign new_n1651 = new_n1646 & ~new_n1650;
  assign new_n1652 = ~new_n1646 & new_n1650;
  assign new_n1653 = n2508 & n7862;
  assign new_n1654 = new_n1365 & new_n1614;
  assign new_n1655 = n1333 & n2509;
  assign new_n1656 = n7862 & n12720;
  assign new_n1657 = ~new_n1617 & ~new_n1656;
  assign new_n1658_1 = new_n1655 & ~new_n1657;
  assign new_n1659 = ~new_n1654 & ~new_n1658_1;
  assign new_n1660 = ~new_n1653 & new_n1659;
  assign new_n1661 = new_n1653 & ~new_n1659;
  assign new_n1662 = ~new_n1606 & ~new_n1607;
  assign new_n1663 = ~new_n1608 & ~new_n1662;
  assign new_n1664 = new_n1608 & new_n1662;
  assign new_n1665 = ~new_n1663 & ~new_n1664;
  assign new_n1666 = ~new_n1661 & ~new_n1665;
  assign new_n1667 = ~new_n1660 & ~new_n1666;
  assign new_n1668 = ~new_n1652 & new_n1667;
  assign new_n1669 = ~new_n1651 & ~new_n1668;
  assign new_n1670 = new_n1645 & ~new_n1669;
  assign new_n1671 = ~new_n1626 & new_n1642;
  assign new_n1672 = ~new_n1601 & ~new_n1671;
  assign new_n1673 = ~new_n1627 & new_n1672;
  assign new_n1674 = new_n1601 & new_n1671;
  assign new_n1675 = ~new_n1673 & ~new_n1674;
  assign new_n1676 = n2509 & n11821;
  assign new_n1677 = n6038 & n9080;
  assign new_n1678 = new_n1618 & new_n1677;
  assign new_n1679 = ~new_n1618 & ~new_n1677;
  assign new_n1680 = ~new_n1678 & ~new_n1679;
  assign new_n1681 = ~new_n1676 & ~new_n1680;
  assign new_n1682 = new_n1676 & new_n1680;
  assign new_n1683 = ~new_n1681 & ~new_n1682;
  assign new_n1684 = n2508 & n11757;
  assign new_n1685 = ~new_n1633 & ~new_n1684;
  assign new_n1686 = new_n1633 & new_n1684;
  assign new_n1687 = ~new_n1685 & ~new_n1686;
  assign new_n1688 = ~new_n1683 & new_n1687;
  assign new_n1689 = new_n1683 & ~new_n1687;
  assign new_n1690 = ~new_n1688 & ~new_n1689;
  assign new_n1691 = ~new_n1636 & new_n1639;
  assign new_n1692 = ~new_n1635 & ~new_n1691;
  assign new_n1693 = n2585 & n3172;
  assign new_n1694 = n7862 & n12706;
  assign new_n1695 = n1333 & n4005;
  assign new_n1696 = ~new_n1694 & ~new_n1695;
  assign new_n1697 = new_n1694 & new_n1695;
  assign new_n1698 = ~new_n1696 & ~new_n1697;
  assign new_n1699 = new_n1693 & ~new_n1698;
  assign new_n1700 = ~new_n1693 & new_n1698;
  assign new_n1701 = ~new_n1699 & ~new_n1700;
  assign new_n1702 = new_n1692 & ~new_n1701;
  assign new_n1703 = ~new_n1692 & new_n1701;
  assign new_n1704 = ~new_n1702 & ~new_n1703;
  assign new_n1705 = ~new_n1690 & ~new_n1704;
  assign new_n1706 = new_n1690 & new_n1704;
  assign new_n1707 = ~new_n1705 & ~new_n1706;
  assign new_n1708 = ~new_n1675 & new_n1707;
  assign new_n1709 = new_n1675 & ~new_n1707;
  assign new_n1710 = ~new_n1708 & ~new_n1709;
  assign new_n1711 = new_n1670 & new_n1710;
  assign new_n1712 = ~new_n1670 & ~new_n1710;
  assign new_n1713 = ~new_n1711 & ~new_n1712;
  assign new_n1714 = n4005 & n7862;
  assign new_n1715 = ~new_n1645 & new_n1669;
  assign new_n1716 = ~new_n1670 & ~new_n1715;
  assign new_n1717 = new_n1714 & new_n1716;
  assign new_n1718 = ~new_n1654 & ~new_n1657;
  assign new_n1719 = n2509 & n7862;
  assign new_n1720 = n1333 & n6038;
  assign new_n1721 = new_n1719 & new_n1720;
  assign new_n1722 = ~new_n1718 & new_n1721;
  assign new_n1723 = ~new_n1660 & ~new_n1661;
  assign new_n1724 = ~new_n1665 & ~new_n1723;
  assign new_n1725 = new_n1665 & new_n1723;
  assign new_n1726 = ~new_n1724 & ~new_n1725;
  assign new_n1727 = new_n1722 & new_n1726;
  assign new_n1728 = ~new_n1651 & ~new_n1652;
  assign new_n1729 = ~new_n1667 & ~new_n1728;
  assign new_n1730 = new_n1667 & new_n1728;
  assign new_n1731 = ~new_n1729 & ~new_n1730;
  assign new_n1732 = new_n1727 & new_n1731;
  assign new_n1733 = ~new_n1714 & ~new_n1716;
  assign new_n1734 = ~new_n1717 & ~new_n1733;
  assign new_n1735 = new_n1732 & new_n1734;
  assign new_n1736 = ~new_n1717 & ~new_n1735;
  assign new_n1737 = new_n1713 & ~new_n1736;
  assign new_n1738 = ~new_n1713 & new_n1736;
  assign new_n1739 = ~new_n1737 & ~new_n1738;
  assign new_n1740 = n4141 & n9400;
  assign new_n1741 = n2464 & n5105;
  assign new_n1742 = new_n1740 & new_n1741;
  assign new_n1743 = ~new_n1740 & ~new_n1741;
  assign new_n1744 = ~new_n1742 & ~new_n1743;
  assign new_n1745 = n5105 & n9400;
  assign new_n1746 = n1209 & n9400;
  assign new_n1747 = n2464 & n7500;
  assign new_n1748 = new_n1746 & new_n1747;
  assign new_n1749 = ~new_n1746 & ~new_n1747;
  assign new_n1750 = n7354 & n11311;
  assign new_n1751 = ~new_n1749 & new_n1750;
  assign new_n1752 = ~new_n1748 & ~new_n1751;
  assign new_n1753 = new_n1745 & ~new_n1752;
  assign new_n1754 = ~new_n1745 & new_n1752;
  assign new_n1755 = n7500 & n11311;
  assign new_n1756 = n1209 & n2464;
  assign new_n1757 = n4187 & n7354;
  assign new_n1758 = ~new_n1756 & ~new_n1757;
  assign new_n1759 = new_n1756 & new_n1757;
  assign new_n1760 = ~new_n1758 & ~new_n1759;
  assign new_n1761 = new_n1755 & ~new_n1760;
  assign new_n1762 = ~new_n1755 & new_n1760;
  assign new_n1763 = ~new_n1761 & ~new_n1762;
  assign new_n1764 = ~new_n1754 & ~new_n1763;
  assign new_n1765 = ~new_n1753 & ~new_n1764;
  assign new_n1766 = ~new_n1744 & new_n1765;
  assign new_n1767 = new_n1744 & ~new_n1765;
  assign new_n1768 = ~new_n1766 & ~new_n1767;
  assign new_n1769 = n1209 & n11311;
  assign new_n1770 = n4187 & n7500;
  assign new_n1771 = n4203 & n7354;
  assign new_n1772 = ~new_n1770 & ~new_n1771;
  assign new_n1773 = new_n1770 & new_n1771;
  assign new_n1774 = ~new_n1772 & ~new_n1773;
  assign new_n1775 = new_n1769 & new_n1774;
  assign new_n1776 = ~new_n1769 & ~new_n1774;
  assign new_n1777 = ~new_n1775 & ~new_n1776;
  assign new_n1778 = new_n1755 & ~new_n1758;
  assign new_n1779 = ~new_n1759 & ~new_n1778;
  assign new_n1780 = ~new_n1777 & ~new_n1779;
  assign new_n1781 = new_n1777 & new_n1779;
  assign new_n1782 = ~new_n1780 & ~new_n1781;
  assign new_n1783 = new_n1768 & ~new_n1782;
  assign new_n1784 = ~new_n1768 & new_n1782;
  assign new_n1785 = ~new_n1783 & ~new_n1784;
  assign new_n1786 = n4141 & n6877;
  assign new_n1787 = n5105 & n6877;
  assign new_n1788 = n7500 & n9400;
  assign new_n1789 = n1209 & n6877;
  assign new_n1790 = new_n1788 & new_n1789;
  assign new_n1791 = n2464 & n7354;
  assign new_n1792 = ~new_n1788 & ~new_n1789;
  assign new_n1793 = new_n1791 & ~new_n1792;
  assign new_n1794 = ~new_n1790 & ~new_n1793;
  assign new_n1795 = ~new_n1787 & new_n1794;
  assign new_n1796 = new_n1787 & ~new_n1794;
  assign new_n1797 = ~new_n1748 & ~new_n1749;
  assign new_n1798_1 = ~new_n1750 & ~new_n1797;
  assign new_n1799 = new_n1750 & new_n1797;
  assign new_n1800 = ~new_n1798_1 & ~new_n1799;
  assign new_n1801 = ~new_n1796 & ~new_n1800;
  assign new_n1802 = ~new_n1795 & ~new_n1801;
  assign new_n1803 = new_n1786 & new_n1802;
  assign new_n1804 = ~new_n1786 & ~new_n1802;
  assign new_n1805 = ~new_n1753 & ~new_n1754;
  assign new_n1806 = new_n1763 & new_n1805;
  assign new_n1807 = ~new_n1763 & ~new_n1805;
  assign new_n1808 = ~new_n1806 & ~new_n1807;
  assign new_n1809 = ~new_n1804 & ~new_n1808;
  assign new_n1810 = ~new_n1803 & ~new_n1809;
  assign new_n1811 = new_n1785 & ~new_n1810;
  assign new_n1812 = ~new_n1766 & ~new_n1782;
  assign new_n1813 = new_n1742 & new_n1812;
  assign new_n1814 = ~new_n1742 & ~new_n1812;
  assign new_n1815 = ~new_n1767 & new_n1814;
  assign new_n1816 = n2464 & n4141;
  assign new_n1817 = n6877 & n8236;
  assign new_n1818 = n4928 & n9400;
  assign new_n1819 = ~new_n1817 & ~new_n1818;
  assign new_n1820 = new_n1817 & new_n1818;
  assign new_n1821 = ~new_n1819 & ~new_n1820;
  assign new_n1822 = new_n1816 & ~new_n1821;
  assign new_n1823 = ~new_n1816 & new_n1821;
  assign new_n1824 = ~new_n1822 & ~new_n1823;
  assign new_n1825 = ~new_n1775 & new_n1779;
  assign new_n1826 = ~new_n1776 & ~new_n1825;
  assign new_n1827 = ~new_n1824 & new_n1826;
  assign new_n1828 = new_n1824 & ~new_n1826;
  assign new_n1829 = ~new_n1827 & ~new_n1828;
  assign new_n1830 = n5105 & n11311;
  assign new_n1831 = new_n1773 & new_n1830;
  assign new_n1832 = ~new_n1773 & ~new_n1830;
  assign new_n1833 = ~new_n1831 & ~new_n1832;
  assign new_n1834 = n4203 & n7500;
  assign new_n1835_1 = n1209 & n4187;
  assign new_n1836 = n7354 & n12753;
  assign new_n1837 = ~new_n1835_1 & ~new_n1836;
  assign new_n1838 = new_n1835_1 & new_n1836;
  assign new_n1839 = ~new_n1837 & ~new_n1838;
  assign new_n1840 = ~new_n1834 & ~new_n1839;
  assign new_n1841 = new_n1834 & new_n1839;
  assign new_n1842 = ~new_n1840 & ~new_n1841;
  assign new_n1843 = new_n1833 & ~new_n1842;
  assign new_n1844 = ~new_n1833 & new_n1842;
  assign new_n1845 = ~new_n1843 & ~new_n1844;
  assign new_n1846 = new_n1829 & new_n1845;
  assign new_n1847_1 = ~new_n1829 & ~new_n1845;
  assign new_n1848 = ~new_n1846 & ~new_n1847_1;
  assign new_n1849 = ~new_n1815 & ~new_n1848;
  assign new_n1850 = ~new_n1813 & ~new_n1849;
  assign new_n1851 = new_n1815 & new_n1848;
  assign new_n1852 = new_n1850 & ~new_n1851;
  assign new_n1853 = new_n1813 & ~new_n1848;
  assign new_n1854 = ~new_n1852 & ~new_n1853;
  assign new_n1855 = new_n1811 & ~new_n1854;
  assign new_n1856 = ~new_n1811 & new_n1854;
  assign new_n1857 = ~new_n1855 & ~new_n1856;
  assign new_n1858 = n4928 & n6877;
  assign new_n1859 = ~new_n1785 & new_n1810;
  assign new_n1860 = ~new_n1811 & ~new_n1859;
  assign new_n1861 = new_n1858 & new_n1860;
  assign new_n1862 = n6877 & n7500;
  assign new_n1863 = n7354 & n9400;
  assign new_n1864 = new_n1862 & new_n1863;
  assign new_n1865 = ~new_n1790 & ~new_n1792;
  assign new_n1866 = ~new_n1791 & ~new_n1865;
  assign new_n1867 = new_n1791 & new_n1865;
  assign new_n1868 = ~new_n1866 & ~new_n1867;
  assign new_n1869 = new_n1864 & new_n1868;
  assign new_n1870 = ~new_n1795 & ~new_n1796;
  assign new_n1871 = ~new_n1800 & new_n1870;
  assign new_n1872 = new_n1800 & ~new_n1870;
  assign new_n1873 = ~new_n1871 & ~new_n1872;
  assign new_n1874 = new_n1869 & ~new_n1873;
  assign new_n1875 = ~new_n1803 & ~new_n1804;
  assign new_n1876 = ~new_n1808 & new_n1875;
  assign new_n1877 = new_n1808 & ~new_n1875;
  assign new_n1878 = ~new_n1876 & ~new_n1877;
  assign new_n1879 = new_n1874 & new_n1878;
  assign new_n1880 = ~new_n1858 & ~new_n1860;
  assign new_n1881 = ~new_n1861 & ~new_n1880;
  assign new_n1882 = new_n1879 & new_n1881;
  assign new_n1883 = ~new_n1861 & ~new_n1882;
  assign new_n1884 = new_n1857 & ~new_n1883;
  assign new_n1885 = ~new_n1857 & new_n1883;
  assign new_n1886 = ~new_n1884 & ~new_n1885;
  assign new_n1887 = n7236 & n12704;
  assign new_n1888 = n7236 & n7294;
  assign new_n1889 = n1980 & n8384;
  assign new_n1890 = new_n1368 & new_n1889;
  assign new_n1891 = n3992 & n10848;
  assign new_n1892 = n8028 & n8384;
  assign new_n1893 = n1980 & n7236;
  assign new_n1894 = ~new_n1892 & ~new_n1893;
  assign new_n1895 = new_n1891 & ~new_n1894;
  assign new_n1896 = ~new_n1890 & ~new_n1895;
  assign new_n1897 = new_n1888 & ~new_n1896;
  assign new_n1898 = ~new_n1888 & new_n1896;
  assign new_n1899 = n6358 & n8028;
  assign new_n1900 = n1980 & n3992;
  assign new_n1901 = n8384 & n10848;
  assign new_n1902 = ~new_n1900 & ~new_n1901;
  assign new_n1903 = new_n1900 & new_n1901;
  assign new_n1904 = ~new_n1902 & ~new_n1903;
  assign new_n1905 = new_n1899 & ~new_n1904;
  assign new_n1906_1 = ~new_n1899 & new_n1904;
  assign new_n1907 = ~new_n1905 & ~new_n1906_1;
  assign new_n1908 = ~new_n1898 & ~new_n1907;
  assign new_n1909 = ~new_n1897 & ~new_n1908;
  assign new_n1910 = new_n1887 & ~new_n1909;
  assign new_n1911 = ~new_n1887 & new_n1909;
  assign new_n1912 = n3992 & n7294;
  assign new_n1913 = new_n1899 & ~new_n1902;
  assign new_n1914 = ~new_n1903 & ~new_n1913;
  assign new_n1915 = ~new_n1912 & new_n1914;
  assign new_n1916 = new_n1912 & ~new_n1914;
  assign new_n1917 = ~new_n1915 & ~new_n1916;
  assign new_n1918 = n6358 & n10848;
  assign new_n1919 = n5198 & n8028;
  assign new_n1920 = ~new_n1889 & ~new_n1919;
  assign new_n1921 = new_n1889 & new_n1919;
  assign new_n1922 = ~new_n1920 & ~new_n1921;
  assign new_n1923 = new_n1918 & ~new_n1922;
  assign new_n1924 = ~new_n1918 & new_n1922;
  assign new_n1925 = ~new_n1923 & ~new_n1924;
  assign new_n1926 = ~new_n1917 & ~new_n1925;
  assign new_n1927 = new_n1917 & new_n1925;
  assign new_n1928 = ~new_n1926 & ~new_n1927;
  assign new_n1929 = ~new_n1911 & ~new_n1928;
  assign new_n1930 = ~new_n1910 & ~new_n1929;
  assign new_n1931 = n7294 & n8384;
  assign new_n1932 = n3992 & n12704;
  assign new_n1933 = ~new_n1931 & ~new_n1932;
  assign new_n1934 = new_n1931 & new_n1932;
  assign new_n1935 = ~new_n1933 & ~new_n1934;
  assign new_n1936 = ~new_n1915 & ~new_n1925;
  assign new_n1937 = ~new_n1916 & ~new_n1936;
  assign new_n1938 = new_n1935 & ~new_n1937;
  assign new_n1939 = ~new_n1935 & new_n1937;
  assign new_n1940 = ~new_n1938 & ~new_n1939;
  assign new_n1941 = n5198 & n10848;
  assign new_n1942 = n1471 & n8028;
  assign new_n1943 = ~new_n1941 & ~new_n1942;
  assign new_n1944 = new_n1941 & new_n1942;
  assign new_n1945 = ~new_n1943 & ~new_n1944;
  assign new_n1946 = n1980 & n6358;
  assign new_n1947 = new_n1918 & ~new_n1920;
  assign new_n1948 = ~new_n1921 & ~new_n1947;
  assign new_n1949 = new_n1946 & ~new_n1948;
  assign new_n1950 = ~new_n1946 & new_n1948;
  assign new_n1951 = ~new_n1949 & ~new_n1950;
  assign new_n1952 = ~new_n1945 & new_n1951;
  assign new_n1953 = new_n1945 & ~new_n1951;
  assign new_n1954 = ~new_n1952 & ~new_n1953;
  assign new_n1955 = new_n1940 & new_n1954;
  assign new_n1956 = ~new_n1940 & ~new_n1954;
  assign new_n1957 = ~new_n1955 & ~new_n1956;
  assign new_n1958 = ~new_n1930 & ~new_n1957;
  assign new_n1959 = ~new_n1939 & ~new_n1954;
  assign new_n1960 = ~new_n1934 & ~new_n1959;
  assign new_n1961 = ~new_n1938 & new_n1960;
  assign new_n1962 = new_n1934 & new_n1959;
  assign new_n1963 = ~new_n1961 & ~new_n1962;
  assign new_n1964 = n3992 & n5814;
  assign new_n1965 = n8384 & n12704;
  assign new_n1966 = n4903 & n7236;
  assign new_n1967 = ~new_n1965 & ~new_n1966;
  assign new_n1968 = new_n1965 & new_n1966;
  assign new_n1969 = ~new_n1967 & ~new_n1968;
  assign new_n1970 = ~new_n1964 & ~new_n1969;
  assign new_n1971 = new_n1964 & new_n1969;
  assign new_n1972 = ~new_n1970 & ~new_n1971;
  assign new_n1973 = new_n1945 & ~new_n1950;
  assign new_n1974 = ~new_n1949 & ~new_n1973;
  assign new_n1975 = new_n1972 & ~new_n1974;
  assign new_n1976 = ~new_n1972 & new_n1974;
  assign new_n1977 = ~new_n1975 & ~new_n1976;
  assign new_n1978 = n6358 & n7294;
  assign new_n1979 = ~new_n1944 & ~new_n1978;
  assign new_n1980_1 = new_n1944 & new_n1978;
  assign new_n1981 = ~new_n1979 & ~new_n1980_1;
  assign new_n1982 = n1471 & n10848;
  assign new_n1983 = n1980 & n5198;
  assign new_n1984 = n7646 & n8028;
  assign new_n1985 = ~new_n1983 & ~new_n1984;
  assign new_n1986 = new_n1983 & new_n1984;
  assign new_n1987 = ~new_n1985 & ~new_n1986;
  assign new_n1988 = ~new_n1982 & ~new_n1987;
  assign new_n1989 = new_n1982 & new_n1987;
  assign new_n1990 = ~new_n1988 & ~new_n1989;
  assign new_n1991 = new_n1981 & ~new_n1990;
  assign new_n1992 = ~new_n1981 & new_n1990;
  assign new_n1993 = ~new_n1991 & ~new_n1992;
  assign new_n1994 = ~new_n1977 & ~new_n1993;
  assign new_n1995 = new_n1977 & new_n1993;
  assign new_n1996 = ~new_n1994 & ~new_n1995;
  assign new_n1997 = ~new_n1963 & new_n1996;
  assign new_n1998 = new_n1963 & ~new_n1996;
  assign new_n1999 = ~new_n1997 & ~new_n1998;
  assign new_n2000 = ~new_n1958 & ~new_n1999;
  assign new_n2001 = new_n1958 & new_n1999;
  assign new_n2002 = ~new_n2000 & ~new_n2001;
  assign new_n2003 = n5814 & n7236;
  assign new_n2004 = new_n1930 & new_n1957;
  assign new_n2005 = ~new_n1958 & ~new_n2004;
  assign new_n2006 = new_n2003 & new_n2005;
  assign new_n2007 = ~new_n1890 & ~new_n1894;
  assign new_n2008 = n7236 & n10848;
  assign new_n2009 = n3992 & n8028;
  assign new_n2010 = new_n2008 & new_n2009;
  assign new_n2011 = ~new_n2007 & new_n2010;
  assign new_n2012 = ~new_n1897 & ~new_n1898;
  assign new_n2013 = new_n1907 & ~new_n2012;
  assign new_n2014 = ~new_n1907 & new_n2012;
  assign new_n2015 = ~new_n2013 & ~new_n2014;
  assign new_n2016 = new_n2011 & new_n2015;
  assign new_n2017 = ~new_n1910 & ~new_n1911;
  assign new_n2018 = new_n1928 & ~new_n2017;
  assign new_n2019 = ~new_n1928 & new_n2017;
  assign new_n2020 = ~new_n2018 & ~new_n2019;
  assign new_n2021 = new_n2016 & new_n2020;
  assign new_n2022 = ~new_n2003 & ~new_n2005;
  assign new_n2023 = ~new_n2006 & ~new_n2022;
  assign new_n2024_1 = new_n2021 & new_n2023;
  assign new_n2025 = ~new_n2006 & ~new_n2024_1;
  assign new_n2026 = ~new_n2002 & new_n2025;
  assign new_n2027 = new_n2002 & ~new_n2025;
  assign new_n2028 = ~new_n2026 & ~new_n2027;
  assign new_n2029 = n4805 & n5069;
  assign new_n2030 = n4805 & n6806;
  assign new_n2031 = n2802 & n11478;
  assign new_n2032 = n533 & n11478;
  assign new_n2033 = n1512 & n5283;
  assign new_n2034 = new_n2032 & new_n2033;
  assign new_n2035 = ~new_n2032 & ~new_n2033;
  assign new_n2036 = n137 & n1564;
  assign new_n2037 = ~new_n2035 & new_n2036;
  assign new_n2038 = ~new_n2034 & ~new_n2037;
  assign new_n2039 = new_n2031 & ~new_n2038;
  assign new_n2040 = ~new_n2031 & new_n2038;
  assign new_n2041 = ~new_n2039 & ~new_n2040;
  assign new_n2042 = n137 & n1512;
  assign new_n2043 = n533 & n5283;
  assign new_n2044 = n1564 & n6294;
  assign new_n2045 = ~new_n2043 & ~new_n2044;
  assign new_n2046 = new_n2043 & new_n2044;
  assign new_n2047 = ~new_n2045 & ~new_n2046;
  assign new_n2048 = new_n2042 & ~new_n2047;
  assign new_n2049 = ~new_n2042 & new_n2047;
  assign new_n2050 = ~new_n2048 & ~new_n2049;
  assign new_n2051 = ~new_n2041 & ~new_n2050;
  assign new_n2052 = new_n2041 & new_n2050;
  assign new_n2053 = ~new_n2051 & ~new_n2052;
  assign new_n2054 = new_n2030 & ~new_n2053;
  assign new_n2055 = ~new_n2030 & new_n2053;
  assign new_n2056 = n2802 & n4805;
  assign new_n2057 = n1512 & n11478;
  assign new_n2058 = n533 & n4805;
  assign new_n2059 = new_n2057 & new_n2058;
  assign new_n2060 = n1564 & n5283;
  assign new_n2061 = ~new_n2057 & ~new_n2058;
  assign new_n2062 = new_n2060 & ~new_n2061;
  assign new_n2063 = ~new_n2059 & ~new_n2062;
  assign new_n2064 = ~new_n2056 & new_n2063;
  assign new_n2065 = new_n2056 & ~new_n2063;
  assign new_n2066 = ~new_n2034 & ~new_n2035;
  assign new_n2067 = ~new_n2036 & ~new_n2066;
  assign new_n2068 = new_n2036 & new_n2066;
  assign new_n2069 = ~new_n2067 & ~new_n2068;
  assign new_n2070 = ~new_n2065 & ~new_n2069;
  assign new_n2071 = ~new_n2064 & ~new_n2070;
  assign new_n2072 = ~new_n2055 & new_n2071;
  assign new_n2073 = ~new_n2054 & ~new_n2072;
  assign new_n2074 = n6806 & n11478;
  assign new_n2075 = n2802 & n5283;
  assign new_n2076 = ~new_n2074 & ~new_n2075;
  assign new_n2077 = new_n2074 & new_n2075;
  assign new_n2078 = ~new_n2076 & ~new_n2077;
  assign new_n2079 = n137 & n533;
  assign new_n2080 = n1512 & n6294;
  assign new_n2081 = n1564 & n6797;
  assign new_n2082 = ~new_n2080 & ~new_n2081;
  assign new_n2083 = new_n2080 & new_n2081;
  assign new_n2084 = ~new_n2082 & ~new_n2083;
  assign new_n2085 = new_n2079 & new_n2084;
  assign new_n2086 = ~new_n2079 & ~new_n2084;
  assign new_n2087_1 = ~new_n2085 & ~new_n2086;
  assign new_n2088 = new_n2042 & ~new_n2045;
  assign new_n2089 = ~new_n2046 & ~new_n2088;
  assign new_n2090 = ~new_n2087_1 & ~new_n2089;
  assign new_n2091 = new_n2087_1 & new_n2089;
  assign new_n2092 = ~new_n2090 & ~new_n2091;
  assign new_n2093 = new_n2078 & ~new_n2092;
  assign new_n2094 = ~new_n2078 & new_n2092;
  assign new_n2095 = ~new_n2093 & ~new_n2094;
  assign new_n2096_1 = ~new_n2040 & ~new_n2050;
  assign new_n2097 = ~new_n2039 & ~new_n2096_1;
  assign new_n2098 = new_n2095 & new_n2097;
  assign new_n2099 = ~new_n2095 & ~new_n2097;
  assign new_n2100 = ~new_n2098 & ~new_n2099;
  assign new_n2101 = ~new_n2073 & ~new_n2100;
  assign new_n2102 = new_n2073 & new_n2100;
  assign new_n2103 = ~new_n2101 & ~new_n2102;
  assign new_n2104 = new_n2029 & new_n2103;
  assign new_n2105 = n1512 & n4805;
  assign new_n2106 = n1564 & n11478;
  assign new_n2107 = new_n2105 & new_n2106;
  assign new_n2108 = ~new_n2059 & ~new_n2061;
  assign new_n2109 = ~new_n2060 & ~new_n2108;
  assign new_n2110 = new_n2060 & new_n2108;
  assign new_n2111 = ~new_n2109 & ~new_n2110;
  assign new_n2112 = new_n2107 & new_n2111;
  assign new_n2113 = ~new_n2064 & ~new_n2065;
  assign new_n2114 = new_n2069 & ~new_n2113;
  assign new_n2115 = ~new_n2069 & new_n2113;
  assign new_n2116 = ~new_n2114 & ~new_n2115;
  assign new_n2117 = new_n2112 & ~new_n2116;
  assign new_n2118 = ~new_n2054 & ~new_n2055;
  assign new_n2119 = new_n2071 & new_n2118;
  assign new_n2120 = ~new_n2071 & ~new_n2118;
  assign new_n2121 = ~new_n2119 & ~new_n2120;
  assign new_n2122 = new_n2117 & new_n2121;
  assign new_n2123 = ~new_n2029 & ~new_n2103;
  assign new_n2124 = ~new_n2104 & ~new_n2123;
  assign new_n2125 = new_n2122 & new_n2124;
  assign new_n2126 = ~new_n2104 & ~new_n2125;
  assign new_n2127 = ~new_n2094 & ~new_n2097;
  assign new_n2128 = ~new_n2077 & ~new_n2127;
  assign new_n2129 = ~new_n2093 & new_n2128;
  assign new_n2130 = new_n2077 & new_n2127;
  assign new_n2131_1 = ~new_n2129 & ~new_n2130;
  assign new_n2132 = n5283 & n6806;
  assign new_n2133 = n4805 & n12044;
  assign new_n2134 = n5069 & n11478;
  assign new_n2135 = ~new_n2133 & ~new_n2134;
  assign new_n2136 = new_n2133 & new_n2134;
  assign new_n2137 = ~new_n2135 & ~new_n2136;
  assign new_n2138 = new_n2132 & ~new_n2137;
  assign new_n2139 = ~new_n2132 & new_n2137;
  assign new_n2140 = ~new_n2138 & ~new_n2139;
  assign new_n2141 = ~new_n2085 & new_n2089;
  assign new_n2142 = ~new_n2086 & ~new_n2141;
  assign new_n2143 = ~new_n2140 & new_n2142;
  assign new_n2144 = new_n2140 & ~new_n2142;
  assign new_n2145 = ~new_n2143 & ~new_n2144;
  assign new_n2146 = n137 & n2802;
  assign new_n2147 = ~new_n2083 & ~new_n2146;
  assign new_n2148 = new_n2083 & new_n2146;
  assign new_n2149 = ~new_n2147 & ~new_n2148;
  assign new_n2150 = n1512 & n6797;
  assign new_n2151 = n533 & n6294;
  assign new_n2152 = n1564 & n3146;
  assign new_n2153 = ~new_n2151 & ~new_n2152;
  assign new_n2154 = new_n2151 & new_n2152;
  assign new_n2155 = ~new_n2153 & ~new_n2154;
  assign new_n2156 = ~new_n2150 & ~new_n2155;
  assign new_n2157 = new_n2150 & new_n2155;
  assign new_n2158 = ~new_n2156 & ~new_n2157;
  assign new_n2159 = new_n2149 & ~new_n2158;
  assign new_n2160 = ~new_n2149 & new_n2158;
  assign new_n2161 = ~new_n2159 & ~new_n2160;
  assign new_n2162 = ~new_n2145 & ~new_n2161;
  assign new_n2163 = new_n2145 & new_n2161;
  assign new_n2164 = ~new_n2162 & ~new_n2163;
  assign new_n2165 = ~new_n2131_1 & new_n2164;
  assign new_n2166 = new_n2131_1 & ~new_n2164;
  assign new_n2167 = ~new_n2165 & ~new_n2166;
  assign new_n2168 = new_n2101 & new_n2167;
  assign new_n2169 = ~new_n2101 & ~new_n2167;
  assign new_n2170 = ~new_n2168 & ~new_n2169;
  assign new_n2171 = ~new_n2126 & new_n2170;
  assign new_n2172 = new_n2126 & ~new_n2170;
  assign new_n2173 = ~new_n2171 & ~new_n2172;
  assign new_n2174 = new_n2028 & new_n2173;
  assign new_n2175 = ~new_n2028 & ~new_n2173;
  assign new_n2176 = ~new_n2174 & ~new_n2175;
  assign new_n2177 = ~new_n2021 & ~new_n2023;
  assign new_n2178 = ~new_n2024_1 & ~new_n2177;
  assign new_n2179 = ~new_n2122 & ~new_n2124;
  assign new_n2180 = ~new_n2125 & ~new_n2179;
  assign new_n2181 = new_n2178 & new_n2180;
  assign new_n2182 = ~new_n2178 & ~new_n2180;
  assign new_n2183 = ~new_n2016 & ~new_n2020;
  assign new_n2184 = ~new_n2021 & ~new_n2183;
  assign new_n2185 = ~new_n2112 & new_n2116;
  assign new_n2186 = ~new_n2117 & ~new_n2185;
  assign new_n2187 = ~new_n2011 & ~new_n2015;
  assign new_n2188 = ~new_n2016 & ~new_n2187;
  assign new_n2189 = new_n2186 & new_n2188;
  assign new_n2190 = ~new_n2186 & ~new_n2188;
  assign new_n2191 = ~new_n2107 & ~new_n2111;
  assign new_n2192 = ~new_n2112 & ~new_n2191;
  assign new_n2193 = ~new_n2105 & ~new_n2106;
  assign new_n2194 = ~new_n2107 & ~new_n2193;
  assign new_n2195 = new_n1369 & new_n2194;
  assign new_n2196 = ~new_n1369 & ~new_n2194;
  assign new_n2197 = ~new_n2008 & ~new_n2009;
  assign new_n2198 = ~new_n2010 & ~new_n2197;
  assign new_n2199 = ~new_n2196 & new_n2198;
  assign new_n2200 = ~new_n2195 & ~new_n2199;
  assign new_n2201 = new_n2192 & ~new_n2200;
  assign new_n2202 = ~new_n2192 & new_n2200;
  assign new_n2203 = ~new_n1368 & new_n1891;
  assign new_n2204 = ~new_n2007 & ~new_n2203;
  assign new_n2205 = ~new_n1368 & new_n1895;
  assign new_n2206 = ~new_n2204 & ~new_n2205;
  assign new_n2207 = ~new_n2202 & new_n2206;
  assign new_n2208 = ~new_n2201 & ~new_n2207;
  assign new_n2209 = ~new_n2190 & ~new_n2208;
  assign new_n2210 = ~new_n2189 & ~new_n2209;
  assign new_n2211 = new_n2184 & ~new_n2210;
  assign new_n2212 = ~new_n2184 & new_n2210;
  assign new_n2213 = ~new_n2117 & ~new_n2121;
  assign new_n2214 = ~new_n2122 & ~new_n2213;
  assign new_n2215 = ~new_n2212 & new_n2214;
  assign new_n2216 = ~new_n2211 & ~new_n2215;
  assign new_n2217 = ~new_n2182 & ~new_n2216;
  assign new_n2218 = ~new_n2181 & ~new_n2217;
  assign new_n2219 = new_n2176 & new_n2218;
  assign new_n2220 = ~new_n2176 & ~new_n2218;
  assign new_n2221 = ~new_n2219 & ~new_n2220;
  assign new_n2222 = new_n1886 & ~new_n2221;
  assign new_n2223 = ~new_n1879 & ~new_n1881;
  assign new_n2224 = ~new_n1882 & ~new_n2223;
  assign new_n2225 = ~new_n2181 & ~new_n2182;
  assign new_n2226_1 = new_n2216 & ~new_n2225;
  assign new_n2227 = ~new_n2216 & new_n2225;
  assign new_n2228 = ~new_n2226_1 & ~new_n2227;
  assign new_n2229 = ~new_n2224 & ~new_n2228;
  assign new_n2230 = new_n2224 & new_n2228;
  assign new_n2231 = ~new_n1874 & ~new_n1878;
  assign new_n2232 = ~new_n1879 & ~new_n2231;
  assign new_n2233 = ~new_n2211 & ~new_n2212;
  assign new_n2234 = ~new_n2214 & ~new_n2233;
  assign new_n2235 = new_n2214 & new_n2233;
  assign new_n2236 = ~new_n2234 & ~new_n2235;
  assign new_n2237 = ~new_n2232 & ~new_n2236;
  assign new_n2238 = new_n2232 & new_n2236;
  assign new_n2239 = ~new_n1869 & new_n1873;
  assign new_n2240 = ~new_n1874 & ~new_n2239;
  assign new_n2241 = ~new_n2189 & ~new_n2190;
  assign new_n2242 = new_n2208 & ~new_n2241;
  assign new_n2243 = ~new_n2208 & new_n2241;
  assign new_n2244 = ~new_n2242 & ~new_n2243;
  assign new_n2245 = ~new_n2240 & ~new_n2244;
  assign new_n2246 = new_n2240 & new_n2244;
  assign new_n2247 = ~new_n1864 & ~new_n1868;
  assign new_n2248 = ~new_n1869 & ~new_n2247;
  assign new_n2249 = ~new_n2201 & ~new_n2202;
  assign new_n2250 = ~new_n2206 & ~new_n2249;
  assign new_n2251 = new_n2206 & new_n2249;
  assign new_n2252 = ~new_n2250 & ~new_n2251;
  assign new_n2253_1 = ~new_n2248 & ~new_n2252;
  assign new_n2254 = new_n2248 & new_n2252;
  assign new_n2255 = ~new_n1862 & ~new_n1863;
  assign new_n2256 = ~new_n1864 & ~new_n2255;
  assign new_n2257 = ~new_n2195 & ~new_n2196;
  assign new_n2258 = new_n2198 & ~new_n2257;
  assign new_n2259 = ~new_n2198 & new_n2257;
  assign new_n2260 = ~new_n2258 & ~new_n2259;
  assign new_n2261 = new_n2256 & ~new_n2260;
  assign new_n2262 = ~new_n2256 & new_n2260;
  assign new_n2263 = new_n1372 & ~new_n2262;
  assign new_n2264 = ~new_n2261 & ~new_n2263;
  assign new_n2265 = ~new_n2254 & new_n2264;
  assign new_n2266 = ~new_n2253_1 & ~new_n2265;
  assign new_n2267 = ~new_n2246 & ~new_n2266;
  assign new_n2268 = ~new_n2245 & ~new_n2267;
  assign new_n2269 = ~new_n2238 & ~new_n2268;
  assign new_n2270 = ~new_n2237 & ~new_n2269;
  assign new_n2271 = ~new_n2230 & ~new_n2270;
  assign new_n2272 = ~new_n2229 & ~new_n2271;
  assign new_n2273 = new_n2222 & new_n2272;
  assign new_n2274 = ~new_n1886 & new_n2221;
  assign new_n2275 = ~new_n2272 & new_n2274;
  assign new_n2276 = ~new_n2222 & ~new_n2272;
  assign new_n2277 = ~new_n2274 & ~new_n2276;
  assign new_n2278_1 = ~new_n2275 & ~new_n2277;
  assign new_n2279 = ~new_n2273 & ~new_n2278_1;
  assign new_n2280 = new_n1739 & ~new_n2279;
  assign new_n2281 = ~new_n1739 & new_n2279;
  assign new_n2282 = ~new_n1732 & ~new_n1734;
  assign new_n2283 = ~new_n1735 & ~new_n2282;
  assign new_n2284 = ~new_n2229 & ~new_n2230;
  assign new_n2285 = new_n2270 & ~new_n2284;
  assign new_n2286 = ~new_n2270 & new_n2284;
  assign new_n2287 = ~new_n2285 & ~new_n2286;
  assign new_n2288 = new_n2283 & ~new_n2287;
  assign new_n2289 = ~new_n2283 & new_n2287;
  assign new_n2290 = ~new_n1727 & ~new_n1731;
  assign new_n2291 = ~new_n1732 & ~new_n2290;
  assign new_n2292 = ~new_n2237 & ~new_n2238;
  assign new_n2293 = new_n2268 & ~new_n2292;
  assign new_n2294 = ~new_n2268 & new_n2292;
  assign new_n2295 = ~new_n2293 & ~new_n2294;
  assign new_n2296 = new_n2291 & ~new_n2295;
  assign new_n2297 = ~new_n2291 & new_n2295;
  assign new_n2298 = ~new_n1722 & ~new_n1726;
  assign new_n2299 = ~new_n1727 & ~new_n2298;
  assign new_n2300 = ~new_n2245 & ~new_n2246;
  assign new_n2301_1 = new_n2266 & ~new_n2300;
  assign new_n2302 = ~new_n2266 & new_n2300;
  assign new_n2303 = ~new_n2301_1 & ~new_n2302;
  assign new_n2304 = new_n2299 & ~new_n2303;
  assign new_n2305 = ~new_n2299 & new_n2303;
  assign new_n2306 = ~new_n1365 & new_n1655;
  assign new_n2307 = new_n1657 & new_n2306;
  assign new_n2308 = new_n1718 & ~new_n2306;
  assign new_n2309 = ~new_n2307 & ~new_n2308;
  assign new_n2310 = ~new_n2253_1 & ~new_n2254;
  assign new_n2311 = new_n2264 & new_n2310;
  assign new_n2312 = ~new_n2264 & ~new_n2310;
  assign new_n2313 = ~new_n2311 & ~new_n2312;
  assign new_n2314 = ~new_n2309 & ~new_n2313;
  assign new_n2315 = new_n2309 & new_n2313;
  assign new_n2316_1 = ~new_n1719 & ~new_n1720;
  assign new_n2317 = ~new_n1721 & ~new_n2316_1;
  assign new_n2318 = new_n1375 & new_n2317;
  assign new_n2319 = ~new_n1375 & ~new_n2317;
  assign new_n2320 = ~new_n2261 & ~new_n2262;
  assign new_n2321 = ~new_n1372 & ~new_n2320;
  assign new_n2322 = new_n1372 & new_n2320;
  assign new_n2323 = ~new_n2321 & ~new_n2322;
  assign new_n2324 = ~new_n2319 & new_n2323;
  assign new_n2325 = ~new_n2318 & ~new_n2324;
  assign new_n2326 = ~new_n2315 & ~new_n2325;
  assign new_n2327 = ~new_n2314 & ~new_n2326;
  assign new_n2328 = ~new_n2305 & ~new_n2327;
  assign new_n2329 = ~new_n2304 & ~new_n2328;
  assign new_n2330 = ~new_n2297 & ~new_n2329;
  assign new_n2331 = ~new_n2296 & ~new_n2330;
  assign new_n2332 = ~new_n2289 & ~new_n2331;
  assign new_n2333 = ~new_n2288 & ~new_n2332;
  assign new_n2334 = ~new_n2281 & ~new_n2333;
  assign new_n2335 = ~new_n2280 & ~new_n2334;
  assign new_n2336 = ~new_n2175 & ~new_n2218;
  assign new_n2337 = ~new_n2174 & ~new_n2336;
  assign new_n2338 = ~new_n1828 & ~new_n1845;
  assign new_n2339 = ~new_n1827 & ~new_n2338;
  assign new_n2340 = n4141 & n11311;
  assign new_n2341 = ~new_n1834 & ~new_n1838;
  assign new_n2342 = ~new_n1837 & ~new_n2341;
  assign new_n2343 = ~new_n2340 & new_n2342;
  assign new_n2344 = new_n2340 & ~new_n2342;
  assign new_n2345 = ~new_n2343 & ~new_n2344;
  assign new_n2346 = new_n2339 & ~new_n2345;
  assign new_n2347_1 = ~new_n2339 & new_n2345;
  assign new_n2348 = ~new_n2346 & ~new_n2347_1;
  assign new_n2349 = ~new_n1831 & ~new_n1842;
  assign new_n2350 = ~new_n1832 & ~new_n2349;
  assign new_n2351 = n4187 & n5105;
  assign new_n2352 = n1209 & n4203;
  assign new_n2353 = ~new_n2351 & new_n2352;
  assign new_n2354 = new_n2351 & ~new_n2352;
  assign new_n2355 = ~new_n2353 & ~new_n2354;
  assign new_n2356 = n8236 & n9400;
  assign new_n2357 = n2464 & n4928;
  assign new_n2358 = ~new_n2356 & new_n2357;
  assign new_n2359 = new_n2356 & ~new_n2357;
  assign new_n2360 = ~new_n2358 & ~new_n2359;
  assign new_n2361 = ~new_n2355 & ~new_n2360;
  assign new_n2362 = new_n2355 & new_n2360;
  assign new_n2363 = ~new_n2361 & ~new_n2362;
  assign new_n2364 = ~new_n2350 & new_n2363;
  assign new_n2365 = new_n2350 & ~new_n2363;
  assign new_n2366 = ~new_n2364 & ~new_n2365;
  assign new_n2367 = new_n2348 & ~new_n2366;
  assign new_n2368 = ~new_n2348 & new_n2366;
  assign new_n2369 = ~new_n2367 & ~new_n2368;
  assign new_n2370 = new_n2337 & new_n2369;
  assign new_n2371 = ~new_n2337 & ~new_n2369;
  assign new_n2372 = ~new_n2370 & ~new_n2371;
  assign new_n2373 = ~new_n2168 & ~new_n2171;
  assign new_n2374 = ~new_n1711 & ~new_n1737;
  assign new_n2375 = new_n2373 & new_n2374;
  assign new_n2376 = ~new_n2373 & ~new_n2374;
  assign new_n2377 = ~new_n2375 & ~new_n2376;
  assign new_n2378 = ~new_n2129 & ~new_n2164;
  assign new_n2379 = ~new_n2130 & ~new_n2378;
  assign new_n2380 = n137 & n6806;
  assign new_n2381 = n2802 & n6294;
  assign new_n2382 = ~new_n2380 & ~new_n2381;
  assign new_n2383_1 = new_n2380 & new_n2381;
  assign new_n2384 = ~new_n2382 & ~new_n2383_1;
  assign new_n2385 = n533 & n6797;
  assign new_n2386 = n1512 & n3146;
  assign new_n2387 = new_n2385 & ~new_n2386;
  assign new_n2388 = ~new_n2385 & new_n2386;
  assign new_n2389 = ~new_n2387 & ~new_n2388;
  assign new_n2390 = ~new_n2384 & ~new_n2389;
  assign new_n2391 = new_n2384 & new_n2389;
  assign new_n2392 = ~new_n2390 & ~new_n2391;
  assign new_n2393_1 = ~new_n2379 & ~new_n2392;
  assign new_n2394 = new_n2379 & new_n2392;
  assign new_n2395 = ~new_n2393_1 & ~new_n2394;
  assign new_n2396 = n1564 & n4938;
  assign new_n2397 = n5814 & n8384;
  assign new_n2398 = ~new_n1980_1 & ~new_n1990;
  assign new_n2399 = ~new_n1979 & ~new_n2398;
  assign new_n2400 = new_n2397 & new_n2399;
  assign new_n2401 = ~new_n2397 & ~new_n2399;
  assign new_n2402 = ~new_n2400 & ~new_n2401;
  assign new_n2403 = ~new_n1975 & new_n1993;
  assign new_n2404 = ~new_n1976 & ~new_n2403;
  assign new_n2405 = ~new_n2402 & new_n2404;
  assign new_n2406 = new_n2402 & ~new_n2404;
  assign new_n2407 = ~new_n2405 & ~new_n2406;
  assign new_n2408 = n4805 & n5694;
  assign new_n2409 = n3992 & n4903;
  assign new_n2410 = n6358 & n12704;
  assign new_n2411 = n5198 & n7294;
  assign new_n2412 = ~new_n2410 & new_n2411;
  assign new_n2413 = new_n2410 & ~new_n2411;
  assign new_n2414 = ~new_n2412 & ~new_n2413;
  assign new_n2415 = new_n2409 & new_n2414;
  assign new_n2416 = ~new_n2409 & ~new_n2414;
  assign new_n2417 = ~new_n2415 & ~new_n2416;
  assign new_n2418 = ~new_n1964 & ~new_n1968;
  assign new_n2419 = ~new_n1967 & ~new_n2418;
  assign new_n2420 = ~new_n2417 & new_n2419;
  assign new_n2421 = new_n2417 & ~new_n2419;
  assign new_n2422 = ~new_n2420 & ~new_n2421;
  assign new_n2423 = ~new_n1982 & ~new_n1986;
  assign new_n2424 = ~new_n1985 & ~new_n2423;
  assign new_n2425_1 = ~new_n2422 & new_n2424;
  assign new_n2426 = new_n2422 & ~new_n2424;
  assign new_n2427 = ~new_n2425_1 & ~new_n2426;
  assign new_n2428 = new_n2408 & new_n2427;
  assign new_n2429 = ~new_n2408 & ~new_n2427;
  assign new_n2430 = ~new_n2428 & ~new_n2429;
  assign new_n2431_1 = ~new_n2407 & new_n2430;
  assign new_n2432 = new_n2407 & ~new_n2430;
  assign new_n2433_1 = ~new_n2431_1 & ~new_n2432;
  assign new_n2434_1 = ~new_n2396 & new_n2433_1;
  assign new_n2435 = new_n2396 & ~new_n2433_1;
  assign new_n2436 = ~new_n2434_1 & ~new_n2435;
  assign new_n2437 = new_n2395 & ~new_n2436;
  assign new_n2438 = ~new_n2395 & new_n2436;
  assign new_n2439 = ~new_n2437 & ~new_n2438;
  assign new_n2440 = ~new_n1673 & ~new_n1707;
  assign new_n2441 = ~new_n1674 & ~new_n2440;
  assign new_n2442 = new_n2132 & ~new_n2135;
  assign new_n2443 = ~new_n2136 & ~new_n2442;
  assign new_n2444 = n615 & n7862;
  assign new_n2445 = n6038 & n6826;
  assign new_n2446 = new_n2444 & ~new_n2445;
  assign new_n2447 = ~new_n2444 & new_n2445;
  assign new_n2448 = ~new_n2446 & ~new_n2447;
  assign new_n2449 = ~new_n2443 & new_n2448;
  assign new_n2450 = new_n2443 & ~new_n2448;
  assign new_n2451 = ~new_n2449 & ~new_n2450;
  assign new_n2452 = ~new_n2144 & ~new_n2161;
  assign new_n2453 = ~new_n2143 & ~new_n2452;
  assign new_n2454 = ~new_n2451 & new_n2453;
  assign new_n2455 = new_n2451 & ~new_n2453;
  assign new_n2456 = ~new_n2454 & ~new_n2455;
  assign new_n2457 = new_n2441 & ~new_n2456;
  assign new_n2458 = ~new_n2441 & new_n2456;
  assign new_n2459 = ~new_n2457 & ~new_n2458;
  assign new_n2460 = ~new_n2150 & ~new_n2154;
  assign new_n2461 = ~new_n2153 & ~new_n2460;
  assign new_n2462 = n11478 & n12044;
  assign new_n2463 = n5069 & n5283;
  assign new_n2464_1 = new_n2462 & ~new_n2463;
  assign new_n2465 = ~new_n2462 & new_n2463;
  assign new_n2466 = ~new_n2464_1 & ~new_n2465;
  assign new_n2467 = ~new_n2461 & ~new_n2466;
  assign new_n2468 = new_n2461 & new_n2466;
  assign new_n2469 = ~new_n2467 & ~new_n2468;
  assign new_n2470 = ~new_n2147 & new_n2158;
  assign new_n2471 = ~new_n2148 & ~new_n2470;
  assign new_n2472 = ~new_n2469 & ~new_n2471;
  assign new_n2473 = new_n2469 & new_n2471;
  assign new_n2474 = ~new_n2472 & ~new_n2473;
  assign new_n2475 = ~new_n2459 & new_n2474;
  assign new_n2476 = new_n2459 & ~new_n2474;
  assign new_n2477 = ~new_n2475 & ~new_n2476;
  assign new_n2478 = ~new_n2439 & new_n2477;
  assign new_n2479 = new_n2439 & ~new_n2477;
  assign new_n2480 = ~new_n2478 & ~new_n2479;
  assign new_n2481 = ~new_n2001 & ~new_n2027;
  assign new_n2482 = ~new_n1816 & ~new_n1820;
  assign new_n2483 = ~new_n1819 & ~new_n2482;
  assign new_n2484 = new_n2481 & new_n2483;
  assign new_n2485 = ~new_n2481 & ~new_n2483;
  assign new_n2486 = ~new_n2484 & ~new_n2485;
  assign new_n2487 = new_n2480 & ~new_n2486;
  assign new_n2488 = ~new_n2480 & new_n2486;
  assign new_n2489 = ~new_n2487 & ~new_n2488;
  assign new_n2490 = ~new_n2377 & new_n2489;
  assign new_n2491 = new_n2377 & ~new_n2489;
  assign new_n2492 = ~new_n2490 & ~new_n2491;
  assign new_n2493 = ~new_n2372 & ~new_n2492;
  assign new_n2494 = new_n2372 & new_n2492;
  assign new_n2495 = ~new_n2493 & ~new_n2494;
  assign new_n2496 = n1471 & n1980;
  assign new_n2497 = n7646 & n10848;
  assign new_n2498_1 = ~new_n2496 & ~new_n2497;
  assign new_n2499 = new_n2496 & new_n2497;
  assign new_n2500 = ~new_n2498_1 & ~new_n2499;
  assign new_n2501 = n1906 & n7236;
  assign new_n2502 = n4722 & n8028;
  assign new_n2503 = new_n2501 & ~new_n2502;
  assign new_n2504 = ~new_n2501 & new_n2502;
  assign new_n2505 = ~new_n2503 & ~new_n2504;
  assign new_n2506 = ~new_n2500 & ~new_n2505;
  assign new_n2507_1 = new_n2500 & new_n2505;
  assign new_n2508_1 = ~new_n2506 & ~new_n2507_1;
  assign new_n2509_1 = ~new_n1855 & ~new_n1884;
  assign new_n2510 = ~new_n1693 & ~new_n1697;
  assign new_n2511 = ~new_n1696 & ~new_n2510;
  assign new_n2512_1 = ~new_n1690 & ~new_n1703;
  assign new_n2513 = ~new_n1702 & ~new_n2512_1;
  assign new_n2514 = ~new_n2511 & new_n2513;
  assign new_n2515_1 = new_n2511 & ~new_n2513;
  assign new_n2516 = ~new_n2514 & ~new_n2515_1;
  assign new_n2517 = new_n2509_1 & ~new_n2516;
  assign new_n2518 = ~new_n2509_1 & new_n2516;
  assign new_n2519 = ~new_n2517 & ~new_n2518;
  assign new_n2520 = ~new_n1961 & ~new_n1996;
  assign new_n2521 = ~new_n1962 & ~new_n2520;
  assign new_n2522_1 = n2508 & n5240;
  assign new_n2523 = n1333 & n12706;
  assign new_n2524 = n3172 & n4005;
  assign new_n2525 = new_n2523 & new_n2524;
  assign new_n2526 = ~new_n2523 & ~new_n2524;
  assign new_n2527 = ~new_n2525 & ~new_n2526;
  assign new_n2528 = new_n2522_1 & ~new_n2527;
  assign new_n2529 = ~new_n2522_1 & new_n2527;
  assign new_n2530_1 = ~new_n2528 & ~new_n2529;
  assign new_n2531 = n2585 & n11757;
  assign new_n2532 = ~new_n1676 & ~new_n1678;
  assign new_n2533 = ~new_n1679 & ~new_n2532;
  assign new_n2534 = new_n2531 & new_n2533;
  assign new_n2535 = ~new_n2531 & ~new_n2533;
  assign new_n2536 = ~new_n2534 & ~new_n2535;
  assign new_n2537 = new_n2530_1 & ~new_n2536;
  assign new_n2538 = ~new_n2530_1 & new_n2536;
  assign new_n2539 = ~new_n2537 & ~new_n2538;
  assign new_n2540 = ~new_n1683 & ~new_n1686;
  assign new_n2541 = ~new_n1685 & ~new_n2540;
  assign new_n2542 = n11821 & n12720;
  assign new_n2543 = n2509 & n9080;
  assign new_n2544 = new_n2542 & new_n2543;
  assign new_n2545 = ~new_n2542 & ~new_n2543;
  assign new_n2546 = ~new_n2544 & ~new_n2545;
  assign new_n2547 = new_n2541 & ~new_n2546;
  assign new_n2548 = ~new_n2541 & new_n2546;
  assign new_n2549 = ~new_n2547 & ~new_n2548;
  assign new_n2550 = ~new_n2539 & ~new_n2549;
  assign new_n2551_1 = new_n2539 & new_n2549;
  assign new_n2552 = ~new_n2550 & ~new_n2551_1;
  assign new_n2553 = n7500 & n12753;
  assign new_n2554 = n7354 & n10174;
  assign new_n2555 = n783 & n6877;
  assign new_n2556 = new_n2554 & ~new_n2555;
  assign new_n2557 = ~new_n2554 & new_n2555;
  assign new_n2558_1 = ~new_n2556 & ~new_n2557;
  assign new_n2559 = new_n2553 & ~new_n2558_1;
  assign new_n2560 = ~new_n2553 & new_n2558_1;
  assign new_n2561 = ~new_n2559 & ~new_n2560;
  assign new_n2562 = new_n1850 & new_n2561;
  assign new_n2563 = ~new_n1850 & ~new_n2561;
  assign new_n2564_1 = ~new_n2562 & ~new_n2563;
  assign new_n2565 = new_n2552 & ~new_n2564_1;
  assign new_n2566 = ~new_n2552 & new_n2564_1;
  assign new_n2567 = ~new_n2565 & ~new_n2566;
  assign new_n2568 = ~new_n2521 & new_n2567;
  assign new_n2569 = new_n2521 & ~new_n2567;
  assign new_n2570 = ~new_n2568 & ~new_n2569;
  assign new_n2571 = new_n2519 & new_n2570;
  assign new_n2572 = ~new_n2519 & ~new_n2570;
  assign new_n2573 = ~new_n2571 & ~new_n2572;
  assign new_n2574 = new_n2508_1 & ~new_n2573;
  assign new_n2575 = ~new_n2508_1 & new_n2573;
  assign new_n2576 = ~new_n2574 & ~new_n2575;
  assign new_n2577_1 = ~new_n2277 & ~new_n2576;
  assign new_n2578 = new_n2277 & new_n2576;
  assign new_n2579 = ~new_n2577_1 & ~new_n2578;
  assign new_n2580 = ~new_n2495 & new_n2579;
  assign new_n2581_1 = new_n2495 & ~new_n2579;
  assign new_n2582 = ~new_n2580 & ~new_n2581_1;
  assign new_n2583 = new_n2335 & ~new_n2582;
  assign new_n2584 = ~new_n2335 & new_n2582;
  assign n671 = new_n2583 | new_n2584;
  assign new_n2586 = n2577 & n5305;
  assign new_n2587 = n3842 & n5964;
  assign new_n2588 = n1097 & n4921;
  assign new_n2589 = n5964 & n11917;
  assign new_n2590 = new_n2588 & new_n2589;
  assign new_n2591 = ~new_n2588 & ~new_n2589;
  assign new_n2592 = n4312 & n9956;
  assign new_n2593 = ~new_n2591 & new_n2592;
  assign new_n2594 = ~new_n2590 & ~new_n2593;
  assign new_n2595 = new_n2587 & ~new_n2594;
  assign new_n2596 = ~new_n2587 & new_n2594;
  assign new_n2597 = ~new_n2595 & ~new_n2596;
  assign new_n2598 = n9956 & n12705;
  assign new_n2599 = n1097 & n11917;
  assign new_n2600 = n4312 & n4921;
  assign new_n2601 = ~new_n2599 & ~new_n2600;
  assign new_n2602 = new_n2599 & new_n2600;
  assign new_n2603 = ~new_n2601 & ~new_n2602;
  assign new_n2604 = new_n2598 & ~new_n2603;
  assign new_n2605 = ~new_n2598 & new_n2603;
  assign new_n2606 = ~new_n2604 & ~new_n2605;
  assign new_n2607 = ~new_n2597 & ~new_n2606;
  assign new_n2608 = new_n2597 & new_n2606;
  assign new_n2609 = ~new_n2607 & ~new_n2608;
  assign new_n2610 = new_n2586 & ~new_n2609;
  assign new_n2611 = ~new_n2586 & new_n2609;
  assign new_n2612 = n3842 & n5305;
  assign new_n2613 = n4921 & n5964;
  assign new_n2614 = n5305 & n11917;
  assign new_n2615 = new_n2613 & new_n2614;
  assign new_n2616 = ~new_n2613 & ~new_n2614;
  assign new_n2617 = n1097 & n9956;
  assign new_n2618 = ~new_n2616 & new_n2617;
  assign new_n2619 = ~new_n2615 & ~new_n2618;
  assign new_n2620 = ~new_n2612 & new_n2619;
  assign new_n2621 = new_n2612 & ~new_n2619;
  assign new_n2622 = ~new_n2590 & ~new_n2591;
  assign new_n2623 = ~new_n2592 & ~new_n2622;
  assign new_n2624_1 = new_n2592 & new_n2622;
  assign new_n2625 = ~new_n2623 & ~new_n2624_1;
  assign new_n2626 = ~new_n2621 & ~new_n2625;
  assign new_n2627 = ~new_n2620 & ~new_n2626;
  assign new_n2628 = ~new_n2611 & new_n2627;
  assign new_n2629 = ~new_n2610 & ~new_n2628;
  assign new_n2630 = n2577 & n5964;
  assign new_n2631 = n1097 & n3842;
  assign new_n2632 = ~new_n2630 & ~new_n2631;
  assign new_n2633 = new_n2630 & new_n2631;
  assign new_n2634 = ~new_n2632 & ~new_n2633;
  assign new_n2635 = n4312 & n11917;
  assign new_n2636 = n4921 & n12705;
  assign new_n2637 = n9956 & n12025;
  assign new_n2638 = ~new_n2636 & ~new_n2637;
  assign new_n2639 = new_n2636 & new_n2637;
  assign new_n2640 = ~new_n2638 & ~new_n2639;
  assign new_n2641 = new_n2635 & new_n2640;
  assign new_n2642 = ~new_n2635 & ~new_n2640;
  assign new_n2643 = ~new_n2641 & ~new_n2642;
  assign new_n2644 = ~new_n2598 & ~new_n2602;
  assign new_n2645 = ~new_n2601 & ~new_n2644;
  assign new_n2646 = ~new_n2643 & ~new_n2645;
  assign new_n2647 = new_n2643 & new_n2645;
  assign new_n2648 = ~new_n2646 & ~new_n2647;
  assign new_n2649 = new_n2634 & new_n2648;
  assign new_n2650 = ~new_n2634 & ~new_n2648;
  assign new_n2651 = ~new_n2649 & ~new_n2650;
  assign new_n2652 = ~new_n2595 & new_n2606;
  assign new_n2653 = ~new_n2596 & ~new_n2652;
  assign new_n2654 = ~new_n2651 & new_n2653;
  assign new_n2655 = new_n2651 & ~new_n2653;
  assign new_n2656 = ~new_n2654 & ~new_n2655;
  assign new_n2657 = ~new_n2629 & ~new_n2656;
  assign new_n2658 = ~new_n2650 & new_n2653;
  assign new_n2659 = ~new_n2633 & ~new_n2658;
  assign new_n2660 = ~new_n2649 & new_n2659;
  assign new_n2661 = new_n2633 & new_n2658;
  assign new_n2662 = ~new_n2660 & ~new_n2661;
  assign new_n2663 = n5964 & n9637;
  assign new_n2664 = n1097 & n2577;
  assign new_n2665 = n1835 & n5305;
  assign new_n2666 = ~new_n2664 & ~new_n2665;
  assign new_n2667 = new_n2664 & new_n2665;
  assign new_n2668 = ~new_n2666 & ~new_n2667;
  assign new_n2669 = ~new_n2663 & ~new_n2668;
  assign new_n2670 = new_n2663 & new_n2668;
  assign new_n2671 = ~new_n2669 & ~new_n2670;
  assign new_n2672 = ~new_n2642 & new_n2645;
  assign new_n2673 = ~new_n2641 & ~new_n2672;
  assign new_n2674 = new_n2671 & ~new_n2673;
  assign new_n2675 = ~new_n2671 & new_n2673;
  assign new_n2676 = ~new_n2674 & ~new_n2675;
  assign new_n2677 = n3842 & n4312;
  assign new_n2678 = new_n2639 & new_n2677;
  assign new_n2679_1 = ~new_n2639 & ~new_n2677;
  assign new_n2680 = ~new_n2678 & ~new_n2679_1;
  assign new_n2681 = n4921 & n12025;
  assign new_n2682 = n11917 & n12705;
  assign new_n2683 = n9956 & n11257;
  assign new_n2684 = ~new_n2682 & ~new_n2683;
  assign new_n2685 = new_n2682 & new_n2683;
  assign new_n2686 = ~new_n2684 & ~new_n2685;
  assign new_n2687 = ~new_n2681 & ~new_n2686;
  assign new_n2688 = new_n2681 & new_n2686;
  assign new_n2689 = ~new_n2687 & ~new_n2688;
  assign new_n2690 = new_n2680 & ~new_n2689;
  assign new_n2691 = ~new_n2680 & new_n2689;
  assign new_n2692 = ~new_n2690 & ~new_n2691;
  assign new_n2693 = new_n2676 & new_n2692;
  assign new_n2694 = ~new_n2676 & ~new_n2692;
  assign new_n2695 = ~new_n2693 & ~new_n2694;
  assign new_n2696 = new_n2662 & new_n2695;
  assign new_n2697 = ~new_n2662 & ~new_n2695;
  assign new_n2698 = ~new_n2696 & ~new_n2697;
  assign new_n2699 = ~new_n2657 & new_n2698;
  assign new_n2700 = new_n2657 & ~new_n2698;
  assign new_n2701 = ~new_n2699 & ~new_n2700;
  assign new_n2702 = n5305 & n9637;
  assign new_n2703 = new_n2629 & new_n2656;
  assign new_n2704 = ~new_n2657 & ~new_n2703;
  assign new_n2705 = new_n2702 & new_n2704;
  assign new_n2706 = n4921 & n5305;
  assign new_n2707 = n5964 & n9956;
  assign new_n2708_1 = new_n2706 & new_n2707;
  assign new_n2709 = ~new_n2615 & ~new_n2616;
  assign new_n2710 = ~new_n2617 & ~new_n2709;
  assign new_n2711 = new_n2617 & new_n2709;
  assign new_n2712 = ~new_n2710 & ~new_n2711;
  assign new_n2713 = new_n2708_1 & new_n2712;
  assign new_n2714 = ~new_n2620 & ~new_n2621;
  assign new_n2715 = ~new_n2625 & ~new_n2714;
  assign new_n2716 = new_n2625 & new_n2714;
  assign new_n2717 = ~new_n2715 & ~new_n2716;
  assign new_n2718 = new_n2713 & new_n2717;
  assign new_n2719 = ~new_n2610 & ~new_n2611;
  assign new_n2720 = ~new_n2627 & ~new_n2719;
  assign new_n2721 = new_n2627 & new_n2719;
  assign new_n2722 = ~new_n2720 & ~new_n2721;
  assign new_n2723 = new_n2718 & new_n2722;
  assign new_n2724 = ~new_n2702 & ~new_n2704;
  assign new_n2725 = ~new_n2705 & ~new_n2724;
  assign new_n2726 = new_n2723 & new_n2725;
  assign new_n2727 = ~new_n2705 & ~new_n2726;
  assign new_n2728 = ~new_n2701 & new_n2727;
  assign new_n2729 = new_n2701 & ~new_n2727;
  assign new_n2730 = ~new_n2728 & ~new_n2729;
  assign new_n2731 = n8065 & n8759;
  assign new_n2732 = n8759 & n10439;
  assign new_n2733 = n6776 & n8595;
  assign new_n2734 = n3602 & n12299;
  assign new_n2735 = n6126 & n6776;
  assign new_n2736 = new_n2734 & new_n2735;
  assign new_n2737 = ~new_n2734 & ~new_n2735;
  assign new_n2738 = n3719 & n7436;
  assign new_n2739 = ~new_n2737 & new_n2738;
  assign new_n2740 = ~new_n2736 & ~new_n2739;
  assign new_n2741 = new_n2733 & ~new_n2740;
  assign new_n2742 = ~new_n2733 & new_n2740;
  assign new_n2743 = ~new_n2741 & ~new_n2742;
  assign new_n2744 = n3719 & n8276;
  assign new_n2745 = n6126 & n12299;
  assign new_n2746 = n3602 & n7436;
  assign new_n2747 = ~new_n2745 & ~new_n2746;
  assign new_n2748 = new_n2745 & new_n2746;
  assign new_n2749_1 = ~new_n2747 & ~new_n2748;
  assign new_n2750 = new_n2744 & ~new_n2749_1;
  assign new_n2751 = ~new_n2744 & new_n2749_1;
  assign new_n2752 = ~new_n2750 & ~new_n2751;
  assign new_n2753 = ~new_n2743 & ~new_n2752;
  assign new_n2754 = new_n2743 & new_n2752;
  assign new_n2755 = ~new_n2753 & ~new_n2754;
  assign new_n2756 = new_n2732 & ~new_n2755;
  assign new_n2757 = ~new_n2732 & new_n2755;
  assign new_n2758 = n8595 & n8759;
  assign new_n2759 = n3719 & n8759;
  assign new_n2760 = new_n2745 & new_n2759;
  assign new_n2761 = n3602 & n6776;
  assign new_n2762 = n6126 & n8759;
  assign new_n2763 = n3719 & n12299;
  assign new_n2764 = ~new_n2762 & ~new_n2763;
  assign new_n2765 = new_n2761 & ~new_n2764;
  assign new_n2766 = ~new_n2760 & ~new_n2765;
  assign new_n2767 = ~new_n2758 & new_n2766;
  assign new_n2768 = new_n2758 & ~new_n2766;
  assign new_n2769 = ~new_n2736 & ~new_n2737;
  assign new_n2770 = ~new_n2738 & ~new_n2769;
  assign new_n2771 = new_n2738 & new_n2769;
  assign new_n2772 = ~new_n2770 & ~new_n2771;
  assign new_n2773 = ~new_n2768 & ~new_n2772;
  assign new_n2774 = ~new_n2767 & ~new_n2773;
  assign new_n2775 = ~new_n2757 & new_n2774;
  assign new_n2776 = ~new_n2756 & ~new_n2775;
  assign new_n2777 = n6776 & n10439;
  assign new_n2778 = n8595 & n12299;
  assign new_n2779 = ~new_n2777 & ~new_n2778;
  assign new_n2780 = new_n2777 & new_n2778;
  assign new_n2781 = ~new_n2779 & ~new_n2780;
  assign new_n2782 = n6126 & n7436;
  assign new_n2783 = n3719 & n9241;
  assign new_n2784 = n3602 & n8276;
  assign new_n2785 = ~new_n2783 & ~new_n2784;
  assign new_n2786 = new_n2783 & new_n2784;
  assign new_n2787 = ~new_n2785 & ~new_n2786;
  assign new_n2788 = new_n2782 & new_n2787;
  assign new_n2789 = ~new_n2782 & ~new_n2787;
  assign new_n2790 = ~new_n2788 & ~new_n2789;
  assign new_n2791 = new_n2744 & ~new_n2747;
  assign new_n2792 = ~new_n2748 & ~new_n2791;
  assign new_n2793 = ~new_n2790 & new_n2792;
  assign new_n2794 = new_n2790 & ~new_n2792;
  assign new_n2795 = ~new_n2793 & ~new_n2794;
  assign new_n2796 = new_n2781 & new_n2795;
  assign new_n2797 = ~new_n2781 & ~new_n2795;
  assign new_n2798 = ~new_n2796 & ~new_n2797;
  assign new_n2799 = ~new_n2741 & new_n2752;
  assign new_n2800 = ~new_n2742 & ~new_n2799;
  assign new_n2801 = ~new_n2798 & new_n2800;
  assign new_n2802_1 = new_n2798 & ~new_n2800;
  assign new_n2803 = ~new_n2801 & ~new_n2802_1;
  assign new_n2804 = ~new_n2776 & ~new_n2803;
  assign new_n2805 = new_n2776 & new_n2803;
  assign new_n2806 = ~new_n2804 & ~new_n2805;
  assign new_n2807 = new_n2731 & new_n2806;
  assign new_n2808 = ~new_n2760 & ~new_n2764;
  assign new_n2809 = n3602 & n8759;
  assign new_n2810 = n3719 & n6776;
  assign new_n2811 = new_n2809 & new_n2810;
  assign new_n2812 = ~new_n2808 & new_n2811;
  assign new_n2813 = ~new_n2767 & ~new_n2768;
  assign new_n2814 = ~new_n2772 & ~new_n2813;
  assign new_n2815 = new_n2772 & new_n2813;
  assign new_n2816 = ~new_n2814 & ~new_n2815;
  assign new_n2817 = new_n2812 & new_n2816;
  assign new_n2818_1 = ~new_n2756 & ~new_n2757;
  assign new_n2819 = ~new_n2774 & ~new_n2818_1;
  assign new_n2820 = new_n2774 & new_n2818_1;
  assign new_n2821 = ~new_n2819 & ~new_n2820;
  assign new_n2822 = new_n2817 & new_n2821;
  assign new_n2823 = ~new_n2731 & ~new_n2806;
  assign new_n2824 = ~new_n2807 & ~new_n2823;
  assign new_n2825 = new_n2822 & new_n2824;
  assign new_n2826 = ~new_n2807 & ~new_n2825;
  assign new_n2827 = ~new_n2797 & new_n2800;
  assign new_n2828 = new_n2780 & new_n2827;
  assign new_n2829 = ~new_n2780 & ~new_n2827;
  assign new_n2830 = ~new_n2796 & new_n2829;
  assign new_n2831 = ~new_n2828 & ~new_n2830;
  assign new_n2832 = n7436 & n8595;
  assign new_n2833 = new_n2786 & new_n2832;
  assign new_n2834 = ~new_n2786 & ~new_n2832;
  assign new_n2835 = ~new_n2833 & ~new_n2834;
  assign new_n2836 = n3719 & n10510;
  assign new_n2837 = n3602 & n9241;
  assign new_n2838 = n6126 & n8276;
  assign new_n2839 = ~new_n2837 & ~new_n2838;
  assign new_n2840 = new_n2837 & new_n2838;
  assign new_n2841 = ~new_n2839 & ~new_n2840;
  assign new_n2842 = new_n2836 & ~new_n2841;
  assign new_n2843 = ~new_n2836 & new_n2841;
  assign new_n2844 = ~new_n2842 & ~new_n2843;
  assign new_n2845 = new_n2835 & new_n2844;
  assign new_n2846 = ~new_n2835 & ~new_n2844;
  assign new_n2847 = ~new_n2845 & ~new_n2846;
  assign new_n2848 = n6776 & n8065;
  assign new_n2849 = n10439 & n12299;
  assign new_n2850 = n8759 & n10391;
  assign new_n2851 = ~new_n2849 & ~new_n2850;
  assign new_n2852 = new_n2849 & new_n2850;
  assign new_n2853 = ~new_n2851 & ~new_n2852;
  assign new_n2854 = ~new_n2848 & ~new_n2853;
  assign new_n2855 = new_n2848 & new_n2853;
  assign new_n2856 = ~new_n2854 & ~new_n2855;
  assign new_n2857 = ~new_n2789 & ~new_n2792;
  assign new_n2858 = ~new_n2788 & ~new_n2857;
  assign new_n2859 = ~new_n2856 & new_n2858;
  assign new_n2860 = new_n2856 & ~new_n2858;
  assign new_n2861 = ~new_n2859 & ~new_n2860;
  assign new_n2862 = ~new_n2847 & ~new_n2861;
  assign new_n2863 = new_n2847 & new_n2861;
  assign new_n2864 = ~new_n2862 & ~new_n2863;
  assign new_n2865 = new_n2831 & new_n2864;
  assign new_n2866 = ~new_n2831 & ~new_n2864;
  assign new_n2867 = ~new_n2865 & ~new_n2866;
  assign new_n2868 = new_n2804 & ~new_n2867;
  assign new_n2869 = ~new_n2804 & new_n2867;
  assign new_n2870 = ~new_n2868 & ~new_n2869;
  assign new_n2871 = ~new_n2826 & new_n2870;
  assign new_n2872 = new_n2826 & ~new_n2870;
  assign new_n2873 = ~new_n2871 & ~new_n2872;
  assign new_n2874 = n4970 & n8476;
  assign new_n2875 = n2530 & n7610;
  assign new_n2876 = ~new_n2874 & ~new_n2875;
  assign new_n2877 = new_n2874 & new_n2875;
  assign new_n2878 = ~new_n2876 & ~new_n2877;
  assign new_n2879_1 = n4826 & n12648;
  assign new_n2880 = n7733 & n10545;
  assign new_n2881 = n7690 & n12925;
  assign new_n2882 = new_n2880 & new_n2881;
  assign new_n2883 = ~new_n2880 & ~new_n2881;
  assign new_n2884 = ~new_n2882 & ~new_n2883;
  assign new_n2885 = new_n2879_1 & new_n2884;
  assign new_n2886 = ~new_n2879_1 & ~new_n2884;
  assign new_n2887 = ~new_n2885 & ~new_n2886;
  assign new_n2888 = n2530 & n12925;
  assign new_n2889 = n4826 & n10545;
  assign new_n2890 = new_n2888 & new_n2889;
  assign new_n2891 = n7733 & n12648;
  assign new_n2892 = n10545 & n12925;
  assign new_n2893 = n2530 & n4826;
  assign new_n2894 = ~new_n2892 & ~new_n2893;
  assign new_n2895 = new_n2891 & ~new_n2894;
  assign new_n2896 = ~new_n2890 & ~new_n2895;
  assign new_n2897 = new_n2887 & new_n2896;
  assign new_n2898 = ~new_n2887 & ~new_n2896;
  assign new_n2899 = ~new_n2897 & ~new_n2898;
  assign new_n2900 = ~new_n2878 & new_n2899;
  assign new_n2901 = new_n2878 & ~new_n2899;
  assign new_n2902_1 = ~new_n2900 & ~new_n2901;
  assign new_n2903 = n7610 & n8476;
  assign new_n2904 = n8476 & n12925;
  assign new_n2905 = new_n2879_1 & new_n2904;
  assign new_n2906 = n2530 & n7733;
  assign new_n2907 = n12648 & n12925;
  assign new_n2908 = n4826 & n8476;
  assign new_n2909 = ~new_n2907 & ~new_n2908;
  assign new_n2910 = new_n2906 & ~new_n2909;
  assign new_n2911 = ~new_n2905 & ~new_n2910;
  assign new_n2912 = ~new_n2903 & new_n2911;
  assign new_n2913 = new_n2903 & ~new_n2911;
  assign new_n2914 = ~new_n2890 & ~new_n2894;
  assign new_n2915 = ~new_n2891 & ~new_n2914;
  assign new_n2916 = new_n2891 & new_n2914;
  assign new_n2917 = ~new_n2915 & ~new_n2916;
  assign new_n2918 = ~new_n2913 & ~new_n2917;
  assign new_n2919 = ~new_n2912 & ~new_n2918;
  assign new_n2920 = ~new_n2902_1 & ~new_n2919;
  assign new_n2921 = new_n2902_1 & new_n2919;
  assign new_n2922 = ~new_n2920 & ~new_n2921;
  assign new_n2923 = n4970 & n5331;
  assign new_n2924 = n5331 & n7610;
  assign new_n2925 = n5331 & n12925;
  assign new_n2926 = new_n2893 & new_n2925;
  assign new_n2927 = n4826 & n5331;
  assign new_n2928 = ~new_n2888 & ~new_n2927;
  assign new_n2929 = n7733 & n8476;
  assign new_n2930 = ~new_n2928 & new_n2929;
  assign new_n2931 = ~new_n2926 & ~new_n2930;
  assign new_n2932 = ~new_n2924 & new_n2931;
  assign new_n2933 = new_n2924 & ~new_n2931;
  assign new_n2934 = ~new_n2905 & ~new_n2909;
  assign new_n2935 = ~new_n2906 & ~new_n2934;
  assign new_n2936 = new_n2906 & new_n2934;
  assign new_n2937 = ~new_n2935 & ~new_n2936;
  assign new_n2938 = ~new_n2933 & ~new_n2937;
  assign new_n2939 = ~new_n2932 & ~new_n2938;
  assign new_n2940 = new_n2923 & new_n2939;
  assign new_n2941 = ~new_n2923 & ~new_n2939;
  assign new_n2942 = ~new_n2912 & ~new_n2913;
  assign new_n2943 = ~new_n2917 & ~new_n2942;
  assign new_n2944 = new_n2917 & new_n2942;
  assign new_n2945 = ~new_n2943 & ~new_n2944;
  assign new_n2946 = ~new_n2941 & new_n2945;
  assign new_n2947 = ~new_n2940 & ~new_n2946;
  assign new_n2948 = new_n2922 & ~new_n2947;
  assign new_n2949 = ~new_n2900 & new_n2919;
  assign new_n2950 = ~new_n2877 & ~new_n2949;
  assign new_n2951 = ~new_n2901 & new_n2950;
  assign new_n2952 = new_n2877 & new_n2949;
  assign new_n2953 = ~new_n2951 & ~new_n2952;
  assign new_n2954 = n503 & n8476;
  assign new_n2955 = n2530 & n4970;
  assign new_n2956 = n5331 & n10965;
  assign new_n2957 = ~new_n2955 & ~new_n2956;
  assign new_n2958 = new_n2955 & new_n2956;
  assign new_n2959 = ~new_n2957 & ~new_n2958;
  assign new_n2960 = ~new_n2954 & ~new_n2959;
  assign new_n2961 = new_n2954 & new_n2959;
  assign new_n2962 = ~new_n2960 & ~new_n2961;
  assign new_n2963 = ~new_n2885 & new_n2896;
  assign new_n2964 = ~new_n2886 & ~new_n2963;
  assign new_n2965 = new_n2962 & new_n2964;
  assign new_n2966 = ~new_n2962 & ~new_n2964;
  assign new_n2967 = ~new_n2965 & ~new_n2966;
  assign new_n2968 = n7690 & n7733;
  assign new_n2969 = n3616 & n12925;
  assign new_n2970 = ~new_n2889 & ~new_n2969;
  assign new_n2971 = new_n2889 & new_n2969;
  assign new_n2972 = ~new_n2970 & ~new_n2971;
  assign new_n2973 = ~new_n2968 & ~new_n2972;
  assign new_n2974 = new_n2968 & new_n2972;
  assign new_n2975 = ~new_n2973 & ~new_n2974;
  assign new_n2976 = n7610 & n12648;
  assign new_n2977 = new_n2882 & new_n2976;
  assign new_n2978 = ~new_n2882 & ~new_n2976;
  assign new_n2979 = ~new_n2977 & ~new_n2978;
  assign new_n2980 = new_n2975 & ~new_n2979;
  assign new_n2981 = ~new_n2975 & new_n2979;
  assign new_n2982 = ~new_n2980 & ~new_n2981;
  assign new_n2983 = new_n2967 & new_n2982;
  assign new_n2984 = ~new_n2967 & ~new_n2982;
  assign new_n2985 = ~new_n2983 & ~new_n2984;
  assign new_n2986 = new_n2953 & ~new_n2985;
  assign new_n2987 = ~new_n2953 & new_n2985;
  assign new_n2988 = ~new_n2986 & ~new_n2987;
  assign new_n2989 = new_n2948 & new_n2988;
  assign new_n2990 = ~new_n2948 & ~new_n2988;
  assign new_n2991 = ~new_n2989 & ~new_n2990;
  assign new_n2992 = n503 & n5331;
  assign new_n2993 = ~new_n2922 & new_n2947;
  assign new_n2994 = ~new_n2948 & ~new_n2993;
  assign new_n2995 = new_n2992 & new_n2994;
  assign new_n2996 = ~new_n2926 & ~new_n2928;
  assign new_n2997 = n5331 & n7733;
  assign new_n2998 = new_n2904 & new_n2997;
  assign new_n2999 = ~new_n2996 & new_n2998;
  assign new_n3000 = ~new_n2932 & ~new_n2933;
  assign new_n3001 = ~new_n2937 & ~new_n3000;
  assign new_n3002 = new_n2937 & new_n3000;
  assign new_n3003 = ~new_n3001 & ~new_n3002;
  assign new_n3004 = new_n2999 & new_n3003;
  assign new_n3005 = new_n2940 & new_n2945;
  assign new_n3006 = new_n2941 & ~new_n2945;
  assign new_n3007 = new_n2947 & ~new_n3006;
  assign new_n3008 = ~new_n3005 & ~new_n3007;
  assign new_n3009 = new_n3004 & ~new_n3008;
  assign new_n3010 = ~new_n2992 & ~new_n2994;
  assign new_n3011 = ~new_n2995 & ~new_n3010;
  assign new_n3012 = new_n3009 & new_n3011;
  assign new_n3013 = ~new_n2995 & ~new_n3012;
  assign new_n3014 = new_n2991 & ~new_n3013;
  assign new_n3015 = ~new_n2991 & new_n3013;
  assign new_n3016 = ~new_n3014 & ~new_n3015;
  assign new_n3017 = n6611 & n7965;
  assign new_n3018 = n217 & n7388;
  assign new_n3019 = n2393 & n4086;
  assign new_n3020 = n7388 & n8433;
  assign new_n3021 = new_n3019 & new_n3020;
  assign new_n3022_1 = n2393 & n8433;
  assign new_n3023 = n4086 & n7388;
  assign new_n3024 = ~new_n3022_1 & ~new_n3023;
  assign new_n3025 = n405 & n11892;
  assign new_n3026 = ~new_n3024 & new_n3025;
  assign new_n3027 = ~new_n3021 & ~new_n3026;
  assign new_n3028 = new_n3018 & ~new_n3027;
  assign new_n3029 = ~new_n3018 & new_n3027;
  assign new_n3030 = ~new_n3028 & ~new_n3029;
  assign new_n3031 = n405 & n2393;
  assign new_n3032 = n5860 & n8433;
  assign new_n3033 = n4086 & n11892;
  assign new_n3034 = ~new_n3032 & ~new_n3033;
  assign new_n3035 = n8433 & n11892;
  assign new_n3036 = n4086 & n5860;
  assign new_n3037 = new_n3035 & new_n3036;
  assign new_n3038 = ~new_n3034 & ~new_n3037;
  assign new_n3039 = ~new_n3031 & ~new_n3038;
  assign new_n3040 = new_n3031 & new_n3038;
  assign new_n3041 = ~new_n3039 & ~new_n3040;
  assign new_n3042 = ~new_n3030 & new_n3041;
  assign new_n3043 = new_n3030 & ~new_n3041;
  assign new_n3044 = ~new_n3042 & ~new_n3043;
  assign new_n3045 = new_n3017 & ~new_n3044;
  assign new_n3046 = ~new_n3017 & new_n3044;
  assign new_n3047 = n217 & n7965;
  assign new_n3048 = n7965 & n8433;
  assign new_n3049 = new_n3033 & new_n3048;
  assign new_n3050 = n4086 & n7965;
  assign new_n3051 = ~new_n3035 & ~new_n3050;
  assign new_n3052 = n405 & n7388;
  assign new_n3053 = ~new_n3051 & new_n3052;
  assign new_n3054 = ~new_n3049 & ~new_n3053;
  assign new_n3055 = ~new_n3047 & new_n3054;
  assign new_n3056 = new_n3047 & ~new_n3054;
  assign new_n3057 = ~new_n3021 & ~new_n3024;
  assign new_n3058 = ~new_n3025 & ~new_n3057;
  assign new_n3059 = new_n3025 & new_n3057;
  assign new_n3060 = ~new_n3058 & ~new_n3059;
  assign new_n3061 = ~new_n3056 & ~new_n3060;
  assign new_n3062 = ~new_n3055 & ~new_n3061;
  assign new_n3063 = ~new_n3046 & new_n3062;
  assign new_n3064 = ~new_n3045 & ~new_n3063;
  assign new_n3065 = n6611 & n7388;
  assign new_n3066 = n217 & n11892;
  assign new_n3067 = ~new_n3065 & ~new_n3066;
  assign new_n3068 = new_n3065 & new_n3066;
  assign new_n3069 = ~new_n3067 & ~new_n3068;
  assign new_n3070 = n405 & n5860;
  assign new_n3071_1 = n3986 & n8433;
  assign new_n3072 = new_n3070 & new_n3071_1;
  assign new_n3073 = ~new_n3070 & ~new_n3071_1;
  assign new_n3074 = ~new_n3072 & ~new_n3073;
  assign new_n3075 = ~new_n3019 & ~new_n3074;
  assign new_n3076 = new_n3019 & new_n3074;
  assign new_n3077 = ~new_n3075 & ~new_n3076;
  assign new_n3078 = new_n3031 & ~new_n3034;
  assign new_n3079 = ~new_n3037 & ~new_n3078;
  assign new_n3080 = ~new_n3077 & new_n3079;
  assign new_n3081 = new_n3077 & ~new_n3079;
  assign new_n3082 = ~new_n3080 & ~new_n3081;
  assign new_n3083 = new_n3069 & new_n3082;
  assign new_n3084 = ~new_n3069 & ~new_n3082;
  assign new_n3085 = ~new_n3083 & ~new_n3084;
  assign new_n3086 = ~new_n3028 & ~new_n3041;
  assign new_n3087 = ~new_n3029 & ~new_n3086;
  assign new_n3088 = new_n3085 & ~new_n3087;
  assign new_n3089 = ~new_n3085 & new_n3087;
  assign new_n3090 = ~new_n3088 & ~new_n3089;
  assign new_n3091 = ~new_n3064 & ~new_n3090;
  assign new_n3092 = ~new_n3084 & new_n3087;
  assign new_n3093 = ~new_n3068 & ~new_n3092;
  assign new_n3094 = ~new_n3083 & new_n3093;
  assign new_n3095 = new_n3068 & new_n3092;
  assign new_n3096 = ~new_n3094 & ~new_n3095;
  assign new_n3097 = n217 & n2393;
  assign new_n3098 = ~new_n3072 & ~new_n3097;
  assign new_n3099 = new_n3072 & new_n3097;
  assign new_n3100 = ~new_n3098 & ~new_n3099;
  assign new_n3101 = n405 & n3986;
  assign new_n3102 = n5857 & n8433;
  assign new_n3103 = new_n3036 & new_n3102;
  assign new_n3104 = ~new_n3036 & ~new_n3102;
  assign new_n3105 = ~new_n3103 & ~new_n3104;
  assign new_n3106 = ~new_n3101 & ~new_n3105;
  assign new_n3107 = new_n3101 & new_n3105;
  assign new_n3108 = ~new_n3106 & ~new_n3107;
  assign new_n3109 = new_n3100 & ~new_n3108;
  assign new_n3110 = ~new_n3100 & new_n3108;
  assign new_n3111 = ~new_n3109 & ~new_n3110;
  assign new_n3112 = n7965 & n11296;
  assign new_n3113 = n6611 & n11892;
  assign new_n3114 = n6359 & n7388;
  assign new_n3115 = ~new_n3113 & ~new_n3114;
  assign new_n3116 = n6359 & n11892;
  assign new_n3117 = new_n3065 & new_n3116;
  assign new_n3118 = ~new_n3115 & ~new_n3117;
  assign new_n3119 = ~new_n3112 & ~new_n3118;
  assign new_n3120 = new_n3112 & new_n3118;
  assign new_n3121 = ~new_n3119 & ~new_n3120;
  assign new_n3122 = ~new_n3076 & new_n3079;
  assign new_n3123 = ~new_n3075 & ~new_n3122;
  assign new_n3124_1 = new_n3121 & new_n3123;
  assign new_n3125 = ~new_n3121 & ~new_n3123;
  assign new_n3126 = ~new_n3124_1 & ~new_n3125;
  assign new_n3127 = ~new_n3111 & ~new_n3126;
  assign new_n3128 = new_n3111 & new_n3126;
  assign new_n3129 = ~new_n3127 & ~new_n3128;
  assign new_n3130 = ~new_n3096 & new_n3129;
  assign new_n3131 = new_n3096 & ~new_n3129;
  assign new_n3132 = ~new_n3130 & ~new_n3131;
  assign new_n3133 = ~new_n3091 & ~new_n3132;
  assign new_n3134 = new_n3091 & new_n3132;
  assign new_n3135 = ~new_n3133 & ~new_n3134;
  assign new_n3136 = n6359 & n7965;
  assign new_n3137 = new_n3064 & new_n3090;
  assign new_n3138 = ~new_n3091 & ~new_n3137;
  assign new_n3139 = new_n3136 & new_n3138;
  assign new_n3140 = ~new_n3049 & ~new_n3051;
  assign new_n3141 = n405 & n7965;
  assign new_n3142 = new_n3020 & new_n3141;
  assign new_n3143 = ~new_n3140 & new_n3142;
  assign new_n3144 = ~new_n3055 & ~new_n3056;
  assign new_n3145 = ~new_n3060 & ~new_n3144;
  assign new_n3146_1 = new_n3060 & new_n3144;
  assign new_n3147 = ~new_n3145 & ~new_n3146_1;
  assign new_n3148 = new_n3143 & new_n3147;
  assign new_n3149 = ~new_n3045 & ~new_n3046;
  assign new_n3150 = ~new_n3062 & ~new_n3149;
  assign new_n3151 = new_n3062 & new_n3149;
  assign new_n3152 = ~new_n3150 & ~new_n3151;
  assign new_n3153 = new_n3148 & new_n3152;
  assign new_n3154 = ~new_n3136 & ~new_n3138;
  assign new_n3155 = ~new_n3139 & ~new_n3154;
  assign new_n3156 = new_n3153 & new_n3155;
  assign new_n3157 = ~new_n3139 & ~new_n3156;
  assign new_n3158 = ~new_n3135 & new_n3157;
  assign new_n3159 = new_n3135 & ~new_n3157;
  assign new_n3160 = ~new_n3158 & ~new_n3159;
  assign new_n3161 = new_n3016 & new_n3160;
  assign new_n3162 = ~new_n3016 & ~new_n3160;
  assign new_n3163 = ~new_n3161 & ~new_n3162;
  assign new_n3164 = ~new_n3009 & ~new_n3011;
  assign new_n3165 = ~new_n3012 & ~new_n3164;
  assign new_n3166 = ~new_n3153 & ~new_n3155;
  assign new_n3167 = ~new_n3156 & ~new_n3166;
  assign new_n3168 = new_n3165 & new_n3167;
  assign new_n3169 = ~new_n3165 & ~new_n3167;
  assign new_n3170 = ~new_n3148 & ~new_n3152;
  assign new_n3171 = ~new_n3153 & ~new_n3170;
  assign new_n3172_1 = ~new_n2999 & ~new_n3003;
  assign new_n3173 = ~new_n3004 & ~new_n3172_1;
  assign new_n3174 = ~new_n3143 & ~new_n3147;
  assign new_n3175 = ~new_n3148 & ~new_n3174;
  assign new_n3176 = new_n3173 & new_n3175;
  assign new_n3177 = ~new_n3173 & ~new_n3175;
  assign new_n3178 = new_n2925 & new_n3048;
  assign new_n3179 = ~new_n3020 & ~new_n3141;
  assign new_n3180 = ~new_n3142 & ~new_n3179;
  assign new_n3181 = new_n3178 & new_n3180;
  assign new_n3182 = ~new_n3178 & ~new_n3180;
  assign new_n3183 = ~new_n2904 & ~new_n2997;
  assign new_n3184 = ~new_n2998 & ~new_n3183;
  assign new_n3185 = ~new_n3182 & new_n3184;
  assign new_n3186 = ~new_n3181 & ~new_n3185;
  assign new_n3187 = ~new_n2925 & new_n2929;
  assign new_n3188 = ~new_n2996 & new_n3187;
  assign new_n3189 = new_n2996 & ~new_n3187;
  assign new_n3190 = ~new_n3188 & ~new_n3189;
  assign new_n3191 = ~new_n3186 & ~new_n3190;
  assign new_n3192 = new_n3186 & new_n3190;
  assign new_n3193 = ~new_n3048 & new_n3052;
  assign new_n3194 = new_n3051 & new_n3193;
  assign new_n3195 = new_n3140 & ~new_n3193;
  assign new_n3196 = ~new_n3194 & ~new_n3195;
  assign new_n3197 = ~new_n3192 & ~new_n3196;
  assign new_n3198 = ~new_n3191 & ~new_n3197;
  assign new_n3199 = ~new_n3177 & ~new_n3198;
  assign new_n3200 = ~new_n3176 & ~new_n3199;
  assign new_n3201 = new_n3171 & ~new_n3200;
  assign new_n3202 = ~new_n3171 & new_n3200;
  assign new_n3203 = ~new_n3004 & new_n3008;
  assign new_n3204 = ~new_n3009 & ~new_n3203;
  assign new_n3205 = ~new_n3202 & new_n3204;
  assign new_n3206 = ~new_n3201 & ~new_n3205;
  assign new_n3207 = ~new_n3169 & ~new_n3206;
  assign new_n3208 = ~new_n3168 & ~new_n3207;
  assign new_n3209 = ~new_n3163 & ~new_n3208;
  assign new_n3210 = new_n3163 & new_n3208;
  assign new_n3211 = ~new_n3209 & ~new_n3210;
  assign new_n3212 = ~new_n2873 & new_n3211;
  assign new_n3213 = new_n2873 & ~new_n3211;
  assign new_n3214_1 = ~new_n3212 & ~new_n3213;
  assign new_n3215 = ~new_n2822 & ~new_n2824;
  assign new_n3216 = ~new_n2825 & ~new_n3215;
  assign new_n3217 = ~new_n2817 & ~new_n2821;
  assign new_n3218 = ~new_n2822 & ~new_n3217;
  assign new_n3219 = ~new_n3201 & ~new_n3202;
  assign new_n3220 = new_n3204 & new_n3219;
  assign new_n3221 = ~new_n3204 & ~new_n3219;
  assign new_n3222 = ~new_n3220 & ~new_n3221;
  assign new_n3223 = ~new_n3218 & ~new_n3222;
  assign new_n3224 = new_n3218 & new_n3222;
  assign new_n3225 = ~new_n2812 & ~new_n2816;
  assign new_n3226 = ~new_n2817 & ~new_n3225;
  assign new_n3227 = ~new_n3176 & ~new_n3177;
  assign new_n3228 = new_n3198 & ~new_n3227;
  assign new_n3229 = ~new_n3198 & new_n3227;
  assign new_n3230_1 = ~new_n3228 & ~new_n3229;
  assign new_n3231 = ~new_n3226 & ~new_n3230_1;
  assign new_n3232 = new_n3226 & new_n3230_1;
  assign new_n3233 = ~new_n2759 & new_n2761;
  assign new_n3234 = new_n2764 & new_n3233;
  assign new_n3235 = new_n2808 & ~new_n3233;
  assign new_n3236 = ~new_n3234 & ~new_n3235;
  assign new_n3237 = ~new_n3191 & ~new_n3192;
  assign new_n3238 = new_n3196 & ~new_n3237;
  assign new_n3239 = ~new_n3196 & new_n3237;
  assign new_n3240 = ~new_n3238 & ~new_n3239;
  assign new_n3241 = new_n3236 & ~new_n3240;
  assign new_n3242 = ~new_n3236 & new_n3240;
  assign new_n3243 = ~new_n2809 & ~new_n2810;
  assign new_n3244 = ~new_n2811 & ~new_n3243;
  assign new_n3245 = ~new_n3181 & ~new_n3182;
  assign new_n3246 = new_n3184 & ~new_n3245;
  assign new_n3247 = ~new_n3184 & new_n3245;
  assign new_n3248 = ~new_n3246 & ~new_n3247;
  assign new_n3249 = new_n3244 & ~new_n3248;
  assign new_n3250 = ~new_n3244 & new_n3248;
  assign new_n3251 = ~new_n2925 & ~new_n3048;
  assign new_n3252 = ~new_n3178 & ~new_n3251;
  assign new_n3253 = new_n2759 & new_n3252;
  assign new_n3254 = ~new_n3250 & new_n3253;
  assign new_n3255 = ~new_n3249 & ~new_n3254;
  assign new_n3256 = ~new_n3242 & new_n3255;
  assign new_n3257 = ~new_n3241 & ~new_n3256;
  assign new_n3258 = ~new_n3232 & ~new_n3257;
  assign new_n3259 = ~new_n3231 & ~new_n3258;
  assign new_n3260 = ~new_n3224 & ~new_n3259;
  assign new_n3261 = ~new_n3223 & ~new_n3260;
  assign new_n3262 = ~new_n3216 & ~new_n3261;
  assign new_n3263 = new_n3216 & new_n3261;
  assign new_n3264 = ~new_n3168 & ~new_n3169;
  assign new_n3265 = new_n3206 & ~new_n3264;
  assign new_n3266 = ~new_n3206 & new_n3264;
  assign new_n3267 = ~new_n3265 & ~new_n3266;
  assign new_n3268 = ~new_n3263 & ~new_n3267;
  assign new_n3269 = ~new_n3262 & ~new_n3268;
  assign new_n3270 = ~new_n3214_1 & ~new_n3269;
  assign new_n3271 = new_n3214_1 & new_n3269;
  assign new_n3272_1 = ~new_n3270 & ~new_n3271;
  assign new_n3273 = new_n2730 & new_n3272_1;
  assign new_n3274 = ~new_n2730 & ~new_n3272_1;
  assign new_n3275 = ~new_n2723 & ~new_n2725;
  assign new_n3276 = ~new_n2726 & ~new_n3275;
  assign new_n3277 = ~new_n3262 & ~new_n3263;
  assign new_n3278 = ~new_n3267 & new_n3277;
  assign new_n3279 = new_n3267 & ~new_n3277;
  assign new_n3280 = ~new_n3278 & ~new_n3279;
  assign new_n3281 = new_n3276 & ~new_n3280;
  assign new_n3282 = ~new_n3276 & new_n3280;
  assign new_n3283 = ~new_n2718 & ~new_n2722;
  assign new_n3284 = ~new_n2723 & ~new_n3283;
  assign new_n3285 = ~new_n3223 & ~new_n3224;
  assign new_n3286 = new_n3259 & ~new_n3285;
  assign new_n3287_1 = ~new_n3259 & new_n3285;
  assign new_n3288 = ~new_n3286 & ~new_n3287_1;
  assign new_n3289 = new_n3284 & ~new_n3288;
  assign new_n3290 = ~new_n3284 & new_n3288;
  assign new_n3291 = ~new_n2713 & ~new_n2717;
  assign new_n3292 = ~new_n2718 & ~new_n3291;
  assign new_n3293 = ~new_n3231 & ~new_n3232;
  assign new_n3294 = new_n3257 & ~new_n3293;
  assign new_n3295 = ~new_n3257 & new_n3293;
  assign new_n3296 = ~new_n3294 & ~new_n3295;
  assign new_n3297 = new_n3292 & ~new_n3296;
  assign new_n3298 = ~new_n3292 & new_n3296;
  assign new_n3299 = ~new_n2708_1 & ~new_n2712;
  assign new_n3300 = ~new_n2713 & ~new_n3299;
  assign new_n3301 = ~new_n3241 & ~new_n3242;
  assign new_n3302 = new_n3255 & new_n3301;
  assign new_n3303 = ~new_n3255 & ~new_n3301;
  assign new_n3304 = ~new_n3302 & ~new_n3303;
  assign new_n3305 = new_n3300 & ~new_n3304;
  assign new_n3306 = ~new_n3300 & new_n3304;
  assign new_n3307 = n5305 & n9956;
  assign new_n3308 = ~new_n2759 & ~new_n3252;
  assign new_n3309 = ~new_n3253 & ~new_n3308;
  assign new_n3310 = new_n3307 & new_n3309;
  assign new_n3311 = ~new_n2706 & ~new_n2707;
  assign new_n3312 = ~new_n2708_1 & ~new_n3311;
  assign new_n3313 = new_n3310 & new_n3312;
  assign new_n3314 = ~new_n3310 & ~new_n3312;
  assign new_n3315 = ~new_n3249 & ~new_n3250;
  assign new_n3316 = new_n3253 & new_n3315;
  assign new_n3317 = ~new_n3253 & ~new_n3315;
  assign new_n3318 = ~new_n3316 & ~new_n3317;
  assign new_n3319 = ~new_n3314 & new_n3318;
  assign new_n3320 = ~new_n3313 & ~new_n3319;
  assign new_n3321 = ~new_n3306 & ~new_n3320;
  assign new_n3322 = ~new_n3305 & ~new_n3321;
  assign new_n3323 = ~new_n3298 & ~new_n3322;
  assign new_n3324 = ~new_n3297 & ~new_n3323;
  assign new_n3325 = ~new_n3290 & ~new_n3324;
  assign new_n3326 = ~new_n3289 & ~new_n3325;
  assign new_n3327 = ~new_n3282 & ~new_n3326;
  assign new_n3328 = ~new_n3281 & ~new_n3327;
  assign new_n3329 = ~new_n3274 & ~new_n3328;
  assign new_n3330 = ~new_n3273 & ~new_n3329;
  assign new_n3331 = ~new_n2989 & ~new_n3014;
  assign new_n3332 = n7388 & n11296;
  assign new_n3333 = ~new_n3116 & ~new_n3332;
  assign new_n3334 = new_n3116 & new_n3332;
  assign new_n3335 = ~new_n3333 & ~new_n3334;
  assign new_n3336 = n2393 & n6611;
  assign new_n3337 = n217 & n5860;
  assign new_n3338 = new_n3336 & ~new_n3337;
  assign new_n3339_1 = ~new_n3336 & new_n3337;
  assign new_n3340 = ~new_n3338 & ~new_n3339_1;
  assign new_n3341 = ~new_n3335 & ~new_n3340;
  assign new_n3342_1 = new_n3335 & new_n3340;
  assign new_n3343 = ~new_n3341 & ~new_n3342_1;
  assign new_n3344 = ~new_n3098 & new_n3108;
  assign new_n3345 = ~new_n3099 & ~new_n3344;
  assign new_n3346 = ~new_n3343 & new_n3345;
  assign new_n3347 = new_n3343 & ~new_n3345;
  assign new_n3348 = ~new_n3346 & ~new_n3347;
  assign new_n3349 = n4970 & n12648;
  assign new_n3350 = n7610 & n10545;
  assign new_n3351 = ~new_n3349 & ~new_n3350;
  assign new_n3352 = new_n3349 & new_n3350;
  assign new_n3353 = ~new_n3351 & ~new_n3352;
  assign new_n3354 = n4826 & n7690;
  assign new_n3355 = n3616 & n7733;
  assign new_n3356 = new_n3354 & ~new_n3355;
  assign new_n3357 = ~new_n3354 & new_n3355;
  assign new_n3358 = ~new_n3356 & ~new_n3357;
  assign new_n3359 = ~new_n3353 & ~new_n3358;
  assign new_n3360 = new_n3353 & new_n3358;
  assign new_n3361 = ~new_n3359 & ~new_n3360;
  assign new_n3362 = ~new_n3348 & new_n3361;
  assign new_n3363 = new_n3348 & ~new_n3361;
  assign new_n3364 = ~new_n3362 & ~new_n3363;
  assign new_n3365 = ~new_n2951 & ~new_n2985;
  assign new_n3366 = ~new_n2952 & ~new_n3365;
  assign new_n3367 = ~new_n3111 & ~new_n3125;
  assign new_n3368 = ~new_n3124_1 & ~new_n3367;
  assign new_n3369 = n5331 & n7546;
  assign new_n3370 = n4499 & n12925;
  assign new_n3371 = ~new_n3369 & new_n3370;
  assign new_n3372 = new_n3369 & ~new_n3370;
  assign new_n3373 = ~new_n3371 & ~new_n3372;
  assign new_n3374 = new_n3112 & ~new_n3115;
  assign new_n3375 = ~new_n3117 & ~new_n3374;
  assign new_n3376 = ~new_n3101 & ~new_n3103;
  assign new_n3377 = ~new_n3104 & ~new_n3376;
  assign new_n3378 = ~new_n3375 & new_n3377;
  assign new_n3379 = new_n3375 & ~new_n3377;
  assign new_n3380 = ~new_n3378 & ~new_n3379;
  assign new_n3381 = ~new_n3373 & new_n3380;
  assign new_n3382 = new_n3373 & ~new_n3380;
  assign new_n3383 = ~new_n3381 & ~new_n3382;
  assign new_n3384 = ~new_n3368 & ~new_n3383;
  assign new_n3385 = new_n3368 & new_n3383;
  assign new_n3386 = ~new_n3384 & ~new_n3385;
  assign new_n3387 = new_n3366 & new_n3386;
  assign new_n3388 = ~new_n3366 & ~new_n3386;
  assign new_n3389 = ~new_n3387 & ~new_n3388;
  assign new_n3390 = new_n3364 & new_n3389;
  assign new_n3391 = ~new_n3364 & ~new_n3389;
  assign new_n3392 = ~new_n3390 & ~new_n3391;
  assign new_n3393 = ~new_n2954 & ~new_n2958;
  assign new_n3394 = ~new_n2957 & ~new_n3393;
  assign new_n3395 = ~new_n2966 & ~new_n2982;
  assign new_n3396 = ~new_n2965 & ~new_n3395;
  assign new_n3397 = ~new_n3394 & ~new_n3396;
  assign new_n3398 = new_n3394 & new_n3396;
  assign new_n3399 = ~new_n3397 & ~new_n3398;
  assign new_n3400 = ~new_n3392 & new_n3399;
  assign new_n3401 = new_n3392 & ~new_n3399;
  assign new_n3402 = ~new_n3400 & ~new_n3401;
  assign new_n3403 = ~new_n3331 & new_n3402;
  assign new_n3404 = new_n3331 & ~new_n3402;
  assign new_n3405 = ~new_n3403 & ~new_n3404;
  assign new_n3406 = ~new_n3330 & new_n3405;
  assign new_n3407 = new_n3330 & ~new_n3405;
  assign new_n3408 = ~new_n3406 & ~new_n3407;
  assign new_n3409 = ~new_n2975 & ~new_n2977;
  assign new_n3410 = ~new_n2978 & ~new_n3409;
  assign new_n3411 = ~new_n2968 & ~new_n2971;
  assign new_n3412 = ~new_n2970 & ~new_n3411;
  assign new_n3413 = n8476 & n10965;
  assign new_n3414 = n503 & n2530;
  assign new_n3415 = new_n3413 & ~new_n3414;
  assign new_n3416 = ~new_n3413 & new_n3414;
  assign new_n3417 = ~new_n3415 & ~new_n3416;
  assign new_n3418 = ~new_n3412 & new_n3417;
  assign new_n3419 = new_n3412 & ~new_n3417;
  assign new_n3420 = ~new_n3418 & ~new_n3419;
  assign new_n3421 = new_n3410 & ~new_n3420;
  assign new_n3422 = ~new_n3410 & new_n3420;
  assign new_n3423 = ~new_n3421 & ~new_n3422;
  assign new_n3424 = ~new_n3213 & ~new_n3269;
  assign new_n3425 = ~new_n3212 & ~new_n3424;
  assign new_n3426 = n1357 & n7965;
  assign new_n3427 = n45 & n8433;
  assign new_n3428 = new_n3426 & ~new_n3427;
  assign new_n3429 = ~new_n3426 & new_n3427;
  assign new_n3430 = ~new_n3428 & ~new_n3429;
  assign new_n3431 = ~new_n3162 & ~new_n3208;
  assign new_n3432 = ~new_n3161 & ~new_n3431;
  assign new_n3433 = n3986 & n4086;
  assign new_n3434 = n405 & n5857;
  assign new_n3435 = ~new_n3433 & ~new_n3434;
  assign new_n3436 = new_n3433 & new_n3434;
  assign new_n3437 = ~new_n3435 & ~new_n3436;
  assign new_n3438 = new_n3432 & new_n3437;
  assign new_n3439 = ~new_n3432 & ~new_n3437;
  assign new_n3440 = ~new_n3438 & ~new_n3439;
  assign new_n3441 = new_n3430 & ~new_n3440;
  assign new_n3442 = ~new_n3430 & new_n3440;
  assign new_n3443 = ~new_n3441 & ~new_n3442;
  assign new_n3444 = ~new_n3425 & ~new_n3443;
  assign new_n3445 = new_n3425 & new_n3443;
  assign new_n3446 = ~new_n3444 & ~new_n3445;
  assign new_n3447 = ~new_n3134 & ~new_n3159;
  assign new_n3448 = ~new_n3094 & ~new_n3129;
  assign new_n3449 = ~new_n3095 & ~new_n3448;
  assign new_n3450 = n6126 & n9241;
  assign new_n3451 = n8276 & n8595;
  assign new_n3452 = ~new_n3450 & new_n3451;
  assign new_n3453 = new_n3450 & ~new_n3451;
  assign new_n3454 = ~new_n3452 & ~new_n3453;
  assign new_n3455 = n8065 & n12299;
  assign new_n3456_1 = n6776 & n10391;
  assign new_n3457 = ~new_n3455 & new_n3456_1;
  assign new_n3458 = new_n3455 & ~new_n3456_1;
  assign new_n3459 = ~new_n3457 & ~new_n3458;
  assign new_n3460 = new_n3454 & ~new_n3459;
  assign new_n3461 = ~new_n3454 & new_n3459;
  assign new_n3462 = ~new_n3460 & ~new_n3461;
  assign new_n3463 = ~new_n2833 & new_n2844;
  assign new_n3464 = ~new_n2834 & ~new_n3463;
  assign new_n3465 = ~new_n3462 & new_n3464;
  assign new_n3466 = new_n3462 & ~new_n3464;
  assign new_n3467 = ~new_n3465 & ~new_n3466;
  assign new_n3468 = new_n2836 & ~new_n2839;
  assign new_n3469 = ~new_n2840 & ~new_n3468;
  assign new_n3470 = ~new_n3467 & new_n3469;
  assign new_n3471 = new_n3467 & ~new_n3469;
  assign new_n3472 = ~new_n3470 & ~new_n3471;
  assign new_n3473 = n7436 & n10439;
  assign new_n3474 = ~new_n2847 & ~new_n2859;
  assign new_n3475 = ~new_n2860 & ~new_n3474;
  assign new_n3476 = new_n3473 & new_n3475;
  assign new_n3477 = ~new_n3473 & ~new_n3475;
  assign new_n3478 = ~new_n3476 & ~new_n3477;
  assign new_n3479 = new_n3472 & new_n3478;
  assign new_n3480 = ~new_n3472 & ~new_n3478;
  assign new_n3481 = ~new_n3479 & ~new_n3480;
  assign new_n3482 = ~new_n2848 & ~new_n2852;
  assign new_n3483 = ~new_n2851 & ~new_n3482;
  assign new_n3484 = ~new_n3481 & new_n3483;
  assign new_n3485 = new_n3481 & ~new_n3483;
  assign new_n3486 = ~new_n3484 & ~new_n3485;
  assign new_n3487 = new_n3449 & ~new_n3486;
  assign new_n3488 = ~new_n3449 & new_n3486;
  assign new_n3489 = ~new_n3487 & ~new_n3488;
  assign new_n3490 = new_n3447 & ~new_n3489;
  assign new_n3491 = ~new_n3447 & new_n3489;
  assign new_n3492 = ~new_n3490 & ~new_n3491;
  assign new_n3493 = ~new_n2868 & ~new_n2871;
  assign new_n3494 = ~new_n2830 & ~new_n2864;
  assign new_n3495 = ~new_n2828 & ~new_n3494;
  assign new_n3496 = n3719 & n10644;
  assign new_n3497 = new_n3495 & ~new_n3496;
  assign new_n3498 = ~new_n3495 & new_n3496;
  assign new_n3499 = ~new_n3497 & ~new_n3498;
  assign new_n3500 = n11917 & n12025;
  assign new_n3501 = n4921 & n11257;
  assign new_n3502 = ~new_n3500 & new_n3501;
  assign new_n3503 = new_n3500 & ~new_n3501;
  assign new_n3504 = ~new_n3502 & ~new_n3503;
  assign new_n3505 = n1835 & n5964;
  assign new_n3506 = n2577 & n4312;
  assign new_n3507 = n3842 & n12705;
  assign new_n3508 = new_n3506 & new_n3507;
  assign new_n3509 = ~new_n3506 & ~new_n3507;
  assign new_n3510 = ~new_n3508 & ~new_n3509;
  assign new_n3511 = new_n3505 & ~new_n3510;
  assign new_n3512 = ~new_n3505 & new_n3510;
  assign new_n3513 = ~new_n3511 & ~new_n3512;
  assign new_n3514 = ~new_n3504 & ~new_n3513;
  assign new_n3515 = new_n3504 & new_n3513;
  assign new_n3516 = ~new_n3514 & ~new_n3515;
  assign new_n3517 = ~new_n2681 & ~new_n2685;
  assign new_n3518 = ~new_n2684 & ~new_n3517;
  assign new_n3519 = ~new_n2663 & ~new_n2667;
  assign new_n3520 = ~new_n2666 & ~new_n3519;
  assign new_n3521 = ~new_n3518 & new_n3520;
  assign new_n3522 = new_n3518 & ~new_n3520;
  assign new_n3523 = ~new_n3521 & ~new_n3522;
  assign new_n3524 = ~new_n3516 & new_n3523;
  assign new_n3525 = new_n3516 & ~new_n3523;
  assign new_n3526 = ~new_n3524 & ~new_n3525;
  assign new_n3527 = n1097 & n9637;
  assign new_n3528 = ~new_n2678 & ~new_n2689;
  assign new_n3529 = ~new_n2679_1 & ~new_n3528;
  assign new_n3530 = new_n3527 & new_n3529;
  assign new_n3531 = ~new_n3527 & ~new_n3529;
  assign new_n3532 = ~new_n3530 & ~new_n3531;
  assign new_n3533 = new_n3526 & new_n3532;
  assign new_n3534 = ~new_n3526 & ~new_n3532;
  assign new_n3535 = ~new_n3533 & ~new_n3534;
  assign new_n3536 = ~new_n2675 & ~new_n2692;
  assign new_n3537 = ~new_n2674 & ~new_n3536;
  assign new_n3538 = ~new_n3535 & new_n3537;
  assign new_n3539 = new_n3535 & ~new_n3537;
  assign new_n3540 = ~new_n3538 & ~new_n3539;
  assign new_n3541 = n4190 & n8759;
  assign new_n3542 = n3602 & n10510;
  assign new_n3543 = ~new_n3541 & ~new_n3542;
  assign new_n3544 = new_n3541 & new_n3542;
  assign new_n3545 = ~new_n3543 & ~new_n3544;
  assign new_n3546 = ~new_n3540 & new_n3545;
  assign new_n3547 = new_n3540 & ~new_n3545;
  assign new_n3548 = ~new_n3546 & ~new_n3547;
  assign new_n3549 = ~new_n3499 & new_n3548;
  assign new_n3550 = new_n3499 & ~new_n3548;
  assign new_n3551 = ~new_n3549 & ~new_n3550;
  assign new_n3552 = new_n3493 & new_n3551;
  assign new_n3553 = ~new_n3493 & ~new_n3551;
  assign new_n3554 = ~new_n3552 & ~new_n3553;
  assign new_n3555 = ~new_n2700 & ~new_n2729;
  assign new_n3556 = ~new_n2660 & ~new_n2695;
  assign new_n3557 = ~new_n2661 & ~new_n3556;
  assign new_n3558 = n9956 & n10547;
  assign new_n3559 = n5305 & n11536;
  assign new_n3560 = ~new_n3558 & new_n3559;
  assign new_n3561 = new_n3558 & ~new_n3559;
  assign new_n3562 = ~new_n3560 & ~new_n3561;
  assign new_n3563 = ~new_n3557 & ~new_n3562;
  assign new_n3564 = new_n3557 & new_n3562;
  assign new_n3565 = ~new_n3563 & ~new_n3564;
  assign new_n3566 = ~new_n3555 & new_n3565;
  assign new_n3567 = new_n3555 & ~new_n3565;
  assign new_n3568 = ~new_n3566 & ~new_n3567;
  assign new_n3569 = ~new_n3554 & new_n3568;
  assign new_n3570 = new_n3554 & ~new_n3568;
  assign new_n3571 = ~new_n3569 & ~new_n3570;
  assign new_n3572 = ~new_n3492 & new_n3571;
  assign new_n3573 = new_n3492 & ~new_n3571;
  assign new_n3574 = ~new_n3572 & ~new_n3573;
  assign new_n3575 = new_n3446 & new_n3574;
  assign new_n3576 = ~new_n3446 & ~new_n3574;
  assign new_n3577 = ~new_n3575 & ~new_n3576;
  assign new_n3578 = new_n3423 & new_n3577;
  assign new_n3579 = ~new_n3423 & ~new_n3577;
  assign new_n3580 = ~new_n3578 & ~new_n3579;
  assign new_n3581 = new_n3408 & new_n3580;
  assign new_n3582 = ~new_n3408 & ~new_n3580;
  assign n837 = ~new_n3581 & ~new_n3582;
  assign new_n3584 = n2577 & n7862;
  assign new_n3585 = n5240 & n9956;
  assign new_n3586 = n3172 & n11917;
  assign new_n3587 = n4921 & n11757;
  assign new_n3588 = ~new_n3586 & ~new_n3587;
  assign new_n3589 = new_n3586 & new_n3587;
  assign new_n3590 = ~new_n3588 & ~new_n3589;
  assign new_n3591 = ~new_n3585 & ~new_n3590;
  assign new_n3592 = new_n3585 & new_n3590;
  assign new_n3593 = ~new_n3591 & ~new_n3592;
  assign new_n3594 = n1333 & n3842;
  assign new_n3595 = n3172 & n4921;
  assign new_n3596 = n1333 & n11917;
  assign new_n3597 = new_n3595 & new_n3596;
  assign new_n3598 = ~new_n3595 & ~new_n3596;
  assign new_n3599 = n9956 & n11757;
  assign new_n3600 = ~new_n3598 & new_n3599;
  assign new_n3601 = ~new_n3597 & ~new_n3600;
  assign new_n3602_1 = ~new_n3594 & new_n3601;
  assign new_n3603 = new_n3594 & ~new_n3601;
  assign new_n3604 = ~new_n3602_1 & ~new_n3603;
  assign new_n3605 = ~new_n3593 & ~new_n3604;
  assign new_n3606 = new_n3593 & new_n3604;
  assign new_n3607 = ~new_n3605 & ~new_n3606;
  assign new_n3608 = ~new_n3584 & ~new_n3607;
  assign new_n3609 = new_n3584 & new_n3607;
  assign new_n3610 = n3842 & n7862;
  assign new_n3611 = n7862 & n9956;
  assign new_n3612 = new_n3586 & new_n3611;
  assign new_n3613 = n1333 & n4921;
  assign new_n3614 = n3172 & n9956;
  assign new_n3615 = n7862 & n11917;
  assign new_n3616_1 = ~new_n3614 & ~new_n3615;
  assign new_n3617 = new_n3613 & ~new_n3616_1;
  assign new_n3618 = ~new_n3612 & ~new_n3617;
  assign new_n3619 = new_n3610 & ~new_n3618;
  assign new_n3620 = ~new_n3610 & new_n3618;
  assign new_n3621 = ~new_n3597 & ~new_n3598;
  assign new_n3622 = new_n3599 & ~new_n3621;
  assign new_n3623 = ~new_n3599 & new_n3621;
  assign new_n3624 = ~new_n3622 & ~new_n3623;
  assign new_n3625 = ~new_n3620 & ~new_n3624;
  assign new_n3626 = ~new_n3619 & ~new_n3625;
  assign new_n3627_1 = ~new_n3609 & new_n3626;
  assign new_n3628 = ~new_n3608 & ~new_n3627_1;
  assign new_n3629 = n1333 & n2577;
  assign new_n3630 = n3172 & n3842;
  assign new_n3631 = ~new_n3629 & ~new_n3630;
  assign new_n3632 = new_n3629 & new_n3630;
  assign new_n3633 = ~new_n3631 & ~new_n3632;
  assign new_n3634 = n11757 & n11917;
  assign new_n3635 = new_n3585 & ~new_n3588;
  assign new_n3636 = ~new_n3595 & ~new_n3635;
  assign new_n3637 = new_n3634 & ~new_n3636;
  assign new_n3638 = ~new_n3634 & ~new_n3635;
  assign new_n3639 = ~new_n3637 & ~new_n3638;
  assign new_n3640 = n4921 & n5240;
  assign new_n3641 = n9956 & n11821;
  assign new_n3642 = ~new_n3640 & ~new_n3641;
  assign new_n3643 = new_n3640 & new_n3641;
  assign new_n3644 = ~new_n3642 & ~new_n3643;
  assign new_n3645 = ~new_n3639 & new_n3644;
  assign new_n3646 = new_n3639 & ~new_n3644;
  assign new_n3647 = ~new_n3645 & ~new_n3646;
  assign new_n3648 = new_n3633 & ~new_n3647;
  assign new_n3649 = ~new_n3633 & new_n3647;
  assign new_n3650 = ~new_n3648 & ~new_n3649;
  assign new_n3651 = ~new_n3593 & ~new_n3603;
  assign new_n3652 = ~new_n3602_1 & ~new_n3651;
  assign new_n3653 = new_n3650 & ~new_n3652;
  assign new_n3654_1 = ~new_n3650 & new_n3652;
  assign new_n3655 = ~new_n3653 & ~new_n3654_1;
  assign new_n3656 = new_n3628 & ~new_n3655;
  assign new_n3657 = ~new_n3648 & ~new_n3652;
  assign new_n3658 = ~new_n3649 & ~new_n3657;
  assign new_n3659 = ~new_n3632 & ~new_n3658;
  assign new_n3660 = new_n3632 & new_n3658;
  assign new_n3661_1 = ~new_n3659 & ~new_n3660;
  assign new_n3662 = ~new_n3638 & new_n3644;
  assign new_n3663 = ~new_n3637 & ~new_n3662;
  assign new_n3664 = n2577 & n3172;
  assign new_n3665 = n1835 & n7862;
  assign new_n3666 = n1333 & n9637;
  assign new_n3667 = ~new_n3665 & ~new_n3666;
  assign new_n3668 = new_n3665 & new_n3666;
  assign new_n3669 = ~new_n3667 & ~new_n3668;
  assign new_n3670 = new_n3664 & ~new_n3669;
  assign new_n3671 = ~new_n3664 & new_n3669;
  assign new_n3672 = ~new_n3670 & ~new_n3671;
  assign new_n3673 = ~new_n3663 & ~new_n3672;
  assign new_n3674 = new_n3663 & new_n3672;
  assign new_n3675 = ~new_n3673 & ~new_n3674;
  assign new_n3676 = n3842 & n11757;
  assign new_n3677_1 = new_n3643 & new_n3676;
  assign new_n3678 = ~new_n3643 & ~new_n3676;
  assign new_n3679 = ~new_n3677_1 & ~new_n3678;
  assign new_n3680 = n4921 & n11821;
  assign new_n3681 = n9080 & n9956;
  assign new_n3682 = n5240 & n11917;
  assign new_n3683 = ~new_n3681 & ~new_n3682;
  assign new_n3684 = new_n3681 & new_n3682;
  assign new_n3685 = ~new_n3683 & ~new_n3684;
  assign new_n3686 = ~new_n3680 & ~new_n3685;
  assign new_n3687 = new_n3680 & new_n3685;
  assign new_n3688 = ~new_n3686 & ~new_n3687;
  assign new_n3689 = new_n3679 & ~new_n3688;
  assign new_n3690 = ~new_n3679 & new_n3688;
  assign new_n3691 = ~new_n3689 & ~new_n3690;
  assign new_n3692 = new_n3675 & new_n3691;
  assign new_n3693 = ~new_n3675 & ~new_n3691;
  assign new_n3694 = ~new_n3692 & ~new_n3693;
  assign new_n3695 = ~new_n3661_1 & new_n3694;
  assign new_n3696 = new_n3661_1 & ~new_n3694;
  assign new_n3697 = ~new_n3695 & ~new_n3696;
  assign new_n3698 = ~new_n3656 & ~new_n3697;
  assign new_n3699 = new_n3656 & new_n3697;
  assign new_n3700 = ~new_n3698 & ~new_n3699;
  assign new_n3701 = n7862 & n9637;
  assign new_n3702 = ~new_n3628 & new_n3655;
  assign new_n3703 = ~new_n3656 & ~new_n3702;
  assign new_n3704 = new_n3701 & new_n3703;
  assign new_n3705 = ~new_n3612 & ~new_n3616_1;
  assign new_n3706 = n4921 & n7862;
  assign new_n3707 = n1333 & n9956;
  assign new_n3708 = new_n3706 & new_n3707;
  assign new_n3709 = ~new_n3705 & new_n3708;
  assign new_n3710 = ~new_n3619 & ~new_n3620;
  assign new_n3711 = new_n3624 & ~new_n3710;
  assign new_n3712 = ~new_n3624 & new_n3710;
  assign new_n3713 = ~new_n3711 & ~new_n3712;
  assign new_n3714 = new_n3709 & new_n3713;
  assign new_n3715 = ~new_n3608 & ~new_n3609;
  assign new_n3716 = ~new_n3626 & ~new_n3715;
  assign new_n3717 = ~new_n3608 & new_n3627_1;
  assign new_n3718 = ~new_n3716 & ~new_n3717;
  assign new_n3719_1 = new_n3714 & ~new_n3718;
  assign new_n3720 = ~new_n3701 & ~new_n3703;
  assign new_n3721 = ~new_n3704 & ~new_n3720;
  assign new_n3722 = new_n3719_1 & new_n3721;
  assign new_n3723 = ~new_n3704 & ~new_n3722;
  assign new_n3724 = ~new_n3700 & new_n3723;
  assign new_n3725 = new_n3700 & ~new_n3723;
  assign new_n3726 = ~new_n3724 & ~new_n3725;
  assign new_n3727 = ~new_n3719_1 & ~new_n3721;
  assign new_n3728 = ~new_n3722 & ~new_n3727;
  assign new_n3729 = ~new_n3714 & new_n3718;
  assign new_n3730 = ~new_n3719_1 & ~new_n3729;
  assign new_n3731 = n3602 & n6877;
  assign new_n3732 = n3719 & n9400;
  assign new_n3733 = new_n3731 & new_n3732;
  assign new_n3734 = n2464 & n3719;
  assign new_n3735 = n3602 & n9400;
  assign new_n3736 = n6126 & n6877;
  assign new_n3737 = ~new_n3735 & ~new_n3736;
  assign new_n3738 = new_n3735 & new_n3736;
  assign new_n3739 = ~new_n3737 & ~new_n3738;
  assign new_n3740 = new_n3734 & ~new_n3739;
  assign new_n3741 = ~new_n3734 & new_n3739;
  assign new_n3742 = ~new_n3740 & ~new_n3741;
  assign new_n3743 = new_n3733 & ~new_n3742;
  assign new_n3744 = n6877 & n8595;
  assign new_n3745 = new_n3734 & ~new_n3737;
  assign new_n3746 = ~new_n3738 & ~new_n3745;
  assign new_n3747 = ~new_n3744 & new_n3746;
  assign new_n3748 = new_n3744 & ~new_n3746;
  assign new_n3749 = ~new_n3747 & ~new_n3748;
  assign new_n3750 = n3719 & n11311;
  assign new_n3751 = n6126 & n9400;
  assign new_n3752 = n2464 & n3602;
  assign new_n3753 = ~new_n3751 & ~new_n3752;
  assign new_n3754_1 = new_n3751 & new_n3752;
  assign new_n3755 = ~new_n3753 & ~new_n3754_1;
  assign new_n3756 = new_n3750 & ~new_n3755;
  assign new_n3757 = ~new_n3750 & new_n3755;
  assign new_n3758 = ~new_n3756 & ~new_n3757;
  assign new_n3759 = ~new_n3749 & new_n3758;
  assign new_n3760 = new_n3749 & ~new_n3758;
  assign new_n3761 = ~new_n3759 & ~new_n3760;
  assign new_n3762 = new_n3743 & new_n3761;
  assign new_n3763 = n6877 & n10439;
  assign new_n3764 = n8595 & n9400;
  assign new_n3765 = new_n3750 & ~new_n3753;
  assign new_n3766 = ~new_n3754_1 & ~new_n3765;
  assign new_n3767 = new_n3764 & ~new_n3766;
  assign new_n3768 = ~new_n3764 & new_n3766;
  assign new_n3769 = ~new_n3767 & ~new_n3768;
  assign new_n3770 = n3602 & n11311;
  assign new_n3771 = n2464 & n6126;
  assign new_n3772 = n3719 & n4187;
  assign new_n3773 = ~new_n3771 & ~new_n3772;
  assign new_n3774 = new_n3771 & new_n3772;
  assign new_n3775 = ~new_n3773 & ~new_n3774;
  assign new_n3776 = new_n3770 & ~new_n3775;
  assign new_n3777 = ~new_n3770 & new_n3775;
  assign new_n3778 = ~new_n3776 & ~new_n3777;
  assign new_n3779 = ~new_n3769 & ~new_n3778;
  assign new_n3780 = new_n3769 & new_n3778;
  assign new_n3781 = ~new_n3779 & ~new_n3780;
  assign new_n3782 = new_n3763 & ~new_n3781;
  assign new_n3783 = ~new_n3763 & new_n3781;
  assign new_n3784 = ~new_n3782 & ~new_n3783;
  assign new_n3785 = ~new_n3747 & ~new_n3758;
  assign new_n3786 = ~new_n3748 & ~new_n3785;
  assign new_n3787 = ~new_n3784 & ~new_n3786;
  assign new_n3788 = new_n3784 & new_n3786;
  assign new_n3789 = ~new_n3787 & ~new_n3788;
  assign new_n3790 = new_n3762 & ~new_n3789;
  assign new_n3791 = ~new_n3762 & new_n3789;
  assign new_n3792 = ~new_n3790 & ~new_n3791;
  assign new_n3793 = ~new_n3743 & ~new_n3761;
  assign new_n3794 = ~new_n3762 & ~new_n3793;
  assign new_n3795 = ~new_n3733 & new_n3742;
  assign new_n3796 = ~new_n3743 & ~new_n3795;
  assign new_n3797 = n5283 & n12925;
  assign new_n3798 = n4805 & n4826;
  assign new_n3799 = ~new_n3797 & ~new_n3798;
  assign new_n3800 = n4805 & n12925;
  assign new_n3801 = n7733 & n11478;
  assign new_n3802 = ~new_n3800 & new_n3801;
  assign new_n3803 = ~new_n3799 & new_n3802;
  assign new_n3804 = n4826 & n5283;
  assign new_n3805 = new_n3800 & new_n3804;
  assign new_n3806 = ~new_n3799 & ~new_n3805;
  assign new_n3807 = ~new_n3802 & ~new_n3806;
  assign new_n3808 = ~new_n3803 & ~new_n3807;
  assign new_n3809 = n8384 & n8433;
  assign new_n3810 = n4086 & n7236;
  assign new_n3811 = ~new_n3809 & ~new_n3810;
  assign new_n3812 = n7236 & n8433;
  assign new_n3813 = n4086 & n8384;
  assign new_n3814 = new_n3812 & new_n3813;
  assign new_n3815 = ~new_n3811 & ~new_n3814;
  assign new_n3816 = n405 & n3992;
  assign new_n3817 = ~new_n3812 & new_n3816;
  assign new_n3818 = new_n3815 & ~new_n3817;
  assign new_n3819 = ~new_n3815 & new_n3817;
  assign new_n3820 = ~new_n3818 & ~new_n3819;
  assign new_n3821 = new_n3800 & new_n3812;
  assign new_n3822 = n4805 & n7733;
  assign new_n3823 = n11478 & n12925;
  assign new_n3824 = ~new_n3822 & ~new_n3823;
  assign new_n3825 = new_n3822 & new_n3823;
  assign new_n3826 = ~new_n3824 & ~new_n3825;
  assign new_n3827 = new_n3821 & new_n3826;
  assign new_n3828 = ~new_n3821 & ~new_n3826;
  assign new_n3829 = n405 & n7236;
  assign new_n3830 = n3992 & n8433;
  assign new_n3831 = ~new_n3829 & ~new_n3830;
  assign new_n3832 = new_n3829 & new_n3830;
  assign new_n3833 = ~new_n3831 & ~new_n3832;
  assign new_n3834 = ~new_n3828 & new_n3833;
  assign new_n3835 = ~new_n3827 & ~new_n3834;
  assign new_n3836 = ~new_n3820 & ~new_n3835;
  assign new_n3837 = new_n3820 & new_n3835;
  assign new_n3838 = ~new_n3836 & ~new_n3837;
  assign new_n3839 = ~new_n3808 & ~new_n3838;
  assign new_n3840 = new_n3808 & new_n3838;
  assign new_n3841 = ~new_n3839 & ~new_n3840;
  assign new_n3842_1 = new_n3796 & new_n3841;
  assign new_n3843 = ~new_n3796 & ~new_n3841;
  assign new_n3844 = ~new_n3731 & ~new_n3732;
  assign new_n3845 = ~new_n3733 & ~new_n3844;
  assign new_n3846 = ~new_n3827 & ~new_n3828;
  assign new_n3847 = new_n3833 & ~new_n3846;
  assign new_n3848 = ~new_n3833 & new_n3846;
  assign new_n3849_1 = ~new_n3847 & ~new_n3848;
  assign new_n3850 = new_n3845 & ~new_n3849_1;
  assign new_n3851 = ~new_n3845 & new_n3849_1;
  assign new_n3852 = n3719 & n6877;
  assign new_n3853 = ~new_n3800 & ~new_n3812;
  assign new_n3854 = ~new_n3821 & ~new_n3853;
  assign new_n3855 = new_n3852 & new_n3854;
  assign new_n3856 = ~new_n3851 & new_n3855;
  assign new_n3857 = ~new_n3850 & ~new_n3856;
  assign new_n3858 = ~new_n3843 & ~new_n3857;
  assign new_n3859 = ~new_n3842_1 & ~new_n3858;
  assign new_n3860 = ~new_n3794 & new_n3859;
  assign new_n3861 = new_n3794 & ~new_n3859;
  assign new_n3862 = ~new_n3806 & new_n3825;
  assign new_n3863 = n4805 & n7610;
  assign new_n3864 = ~new_n3801 & ~new_n3805;
  assign new_n3865_1 = ~new_n3799 & ~new_n3864;
  assign new_n3866 = new_n3863 & new_n3865_1;
  assign new_n3867 = ~new_n3863 & ~new_n3865_1;
  assign new_n3868 = ~new_n3866 & ~new_n3867;
  assign new_n3869 = n5283 & n7733;
  assign new_n3870 = n137 & n12925;
  assign new_n3871 = n4826 & n11478;
  assign new_n3872 = ~new_n3870 & ~new_n3871;
  assign new_n3873 = new_n3870 & new_n3871;
  assign new_n3874 = ~new_n3872 & ~new_n3873;
  assign new_n3875 = new_n3869 & ~new_n3874;
  assign new_n3876 = ~new_n3869 & new_n3874;
  assign new_n3877 = ~new_n3875 & ~new_n3876;
  assign new_n3878 = ~new_n3868 & ~new_n3877;
  assign new_n3879 = new_n3868 & new_n3877;
  assign new_n3880 = ~new_n3878 & ~new_n3879;
  assign new_n3881 = new_n3862 & ~new_n3880;
  assign new_n3882 = ~new_n3862 & new_n3880;
  assign new_n3883 = ~new_n3881 & ~new_n3882;
  assign new_n3884 = ~new_n3815 & new_n3832;
  assign new_n3885 = n217 & n7236;
  assign new_n3886 = ~new_n3814 & ~new_n3816;
  assign new_n3887 = ~new_n3811 & ~new_n3886;
  assign new_n3888 = new_n3885 & new_n3887;
  assign new_n3889 = ~new_n3885 & ~new_n3887;
  assign new_n3890 = ~new_n3888 & ~new_n3889;
  assign new_n3891 = n405 & n8384;
  assign new_n3892 = n6358 & n8433;
  assign new_n3893 = n3992 & n4086;
  assign new_n3894 = ~new_n3892 & ~new_n3893;
  assign new_n3895 = new_n3892 & new_n3893;
  assign new_n3896 = ~new_n3894 & ~new_n3895;
  assign new_n3897 = new_n3891 & ~new_n3896;
  assign new_n3898 = ~new_n3891 & new_n3896;
  assign new_n3899 = ~new_n3897 & ~new_n3898;
  assign new_n3900 = ~new_n3890 & ~new_n3899;
  assign new_n3901 = new_n3890 & new_n3899;
  assign new_n3902 = ~new_n3900 & ~new_n3901;
  assign new_n3903 = new_n3884 & ~new_n3902;
  assign new_n3904 = ~new_n3884 & new_n3902;
  assign new_n3905 = ~new_n3903 & ~new_n3904;
  assign new_n3906 = new_n3883 & new_n3905;
  assign new_n3907 = ~new_n3883 & ~new_n3905;
  assign new_n3908 = ~new_n3906 & ~new_n3907;
  assign new_n3909 = ~new_n3808 & ~new_n3836;
  assign new_n3910 = ~new_n3837 & ~new_n3909;
  assign new_n3911 = ~new_n3908 & ~new_n3910;
  assign new_n3912 = new_n3908 & new_n3910;
  assign new_n3913 = ~new_n3911 & ~new_n3912;
  assign new_n3914 = ~new_n3861 & ~new_n3913;
  assign new_n3915 = ~new_n3860 & ~new_n3914;
  assign new_n3916 = new_n3792 & new_n3915;
  assign new_n3917 = ~new_n3792 & ~new_n3915;
  assign new_n3918 = ~new_n3916 & ~new_n3917;
  assign new_n3919 = n6611 & n7236;
  assign new_n3920 = n217 & n3992;
  assign new_n3921 = new_n3891 & ~new_n3894;
  assign new_n3922 = ~new_n3895 & ~new_n3921;
  assign new_n3923 = new_n3920 & ~new_n3922;
  assign new_n3924 = ~new_n3920 & new_n3922;
  assign new_n3925 = ~new_n3923 & ~new_n3924;
  assign new_n3926 = n405 & n6358;
  assign new_n3927 = n5198 & n8433;
  assign new_n3928 = ~new_n3813 & ~new_n3927;
  assign new_n3929 = new_n3813 & new_n3927;
  assign new_n3930 = ~new_n3928 & ~new_n3929;
  assign new_n3931 = new_n3926 & ~new_n3930;
  assign new_n3932_1 = ~new_n3926 & new_n3930;
  assign new_n3933 = ~new_n3931 & ~new_n3932_1;
  assign new_n3934 = ~new_n3925 & ~new_n3933;
  assign new_n3935 = new_n3925 & new_n3933;
  assign new_n3936 = ~new_n3934 & ~new_n3935;
  assign new_n3937 = new_n3919 & ~new_n3936;
  assign new_n3938 = ~new_n3919 & new_n3936;
  assign new_n3939 = ~new_n3937 & ~new_n3938;
  assign new_n3940 = ~new_n3889 & ~new_n3899;
  assign new_n3941 = ~new_n3888 & ~new_n3940;
  assign new_n3942 = ~new_n3939 & ~new_n3941;
  assign new_n3943 = new_n3939 & new_n3941;
  assign new_n3944 = ~new_n3942 & ~new_n3943;
  assign new_n3945 = new_n3903 & ~new_n3944;
  assign new_n3946 = ~new_n3903 & new_n3944;
  assign new_n3947 = ~new_n3945 & ~new_n3946;
  assign new_n3948 = n4805 & n4970;
  assign new_n3949 = n7610 & n11478;
  assign new_n3950 = new_n3869 & ~new_n3872;
  assign new_n3951 = ~new_n3873 & ~new_n3950;
  assign new_n3952 = new_n3949 & ~new_n3951;
  assign new_n3953 = ~new_n3949 & new_n3951;
  assign new_n3954 = ~new_n3952 & ~new_n3953;
  assign new_n3955 = n137 & n7733;
  assign new_n3956 = n6294 & n12925;
  assign new_n3957 = ~new_n3804 & ~new_n3956;
  assign new_n3958 = new_n3804 & new_n3956;
  assign new_n3959 = ~new_n3957 & ~new_n3958;
  assign new_n3960 = new_n3955 & ~new_n3959;
  assign new_n3961 = ~new_n3955 & new_n3959;
  assign new_n3962 = ~new_n3960 & ~new_n3961;
  assign new_n3963 = ~new_n3954 & ~new_n3962;
  assign new_n3964 = new_n3954 & new_n3962;
  assign new_n3965 = ~new_n3963 & ~new_n3964;
  assign new_n3966 = new_n3948 & ~new_n3965;
  assign new_n3967 = ~new_n3948 & new_n3965;
  assign new_n3968 = ~new_n3966 & ~new_n3967;
  assign new_n3969 = ~new_n3867 & ~new_n3877;
  assign new_n3970 = ~new_n3866 & ~new_n3969;
  assign new_n3971 = ~new_n3968 & ~new_n3970;
  assign new_n3972 = new_n3968 & new_n3970;
  assign new_n3973 = ~new_n3971 & ~new_n3972;
  assign new_n3974 = new_n3881 & ~new_n3973;
  assign new_n3975 = ~new_n3881 & new_n3973;
  assign new_n3976 = ~new_n3974 & ~new_n3975;
  assign new_n3977 = ~new_n3906 & ~new_n3910;
  assign new_n3978 = ~new_n3907 & ~new_n3977;
  assign new_n3979 = new_n3976 & new_n3978;
  assign new_n3980 = ~new_n3976 & ~new_n3978;
  assign new_n3981 = ~new_n3979 & ~new_n3980;
  assign new_n3982 = ~new_n3947 & new_n3981;
  assign new_n3983 = new_n3947 & ~new_n3981;
  assign new_n3984 = ~new_n3982 & ~new_n3983;
  assign new_n3985 = new_n3918 & new_n3984;
  assign new_n3986_1 = ~new_n3918 & ~new_n3984;
  assign new_n3987 = ~new_n3985 & ~new_n3986_1;
  assign new_n3988 = new_n3730 & ~new_n3987;
  assign new_n3989 = ~new_n3730 & new_n3987;
  assign new_n3990 = ~new_n3709 & ~new_n3713;
  assign new_n3991 = ~new_n3714 & ~new_n3990;
  assign new_n3992_1 = ~new_n3860 & ~new_n3861;
  assign new_n3993 = ~new_n3913 & new_n3992_1;
  assign new_n3994 = new_n3913 & ~new_n3992_1;
  assign new_n3995 = ~new_n3993 & ~new_n3994;
  assign new_n3996 = new_n3991 & ~new_n3995;
  assign new_n3997 = ~new_n3991 & new_n3995;
  assign new_n3998 = ~new_n3611 & new_n3613;
  assign new_n3999 = ~new_n3705 & ~new_n3998;
  assign new_n4000 = ~new_n3616_1 & new_n3998;
  assign new_n4001 = ~new_n3999 & ~new_n4000;
  assign new_n4002 = ~new_n3842_1 & ~new_n3843;
  assign new_n4003 = new_n3857 & ~new_n4002;
  assign new_n4004 = ~new_n3857 & new_n4002;
  assign new_n4005_1 = ~new_n4003 & ~new_n4004;
  assign new_n4006 = new_n4001 & new_n4005_1;
  assign new_n4007 = ~new_n4001 & ~new_n4005_1;
  assign new_n4008 = ~new_n3852 & ~new_n3854;
  assign new_n4009 = ~new_n3855 & ~new_n4008;
  assign new_n4010 = new_n3611 & new_n4009;
  assign new_n4011 = ~new_n3706 & ~new_n3707;
  assign new_n4012 = ~new_n3708 & ~new_n4011;
  assign new_n4013 = ~new_n4010 & ~new_n4012;
  assign new_n4014 = new_n4010 & new_n4012;
  assign new_n4015 = ~new_n3850 & ~new_n3851;
  assign new_n4016 = ~new_n3855 & ~new_n4015;
  assign new_n4017 = new_n3855 & new_n4015;
  assign new_n4018 = ~new_n4016 & ~new_n4017;
  assign new_n4019 = ~new_n4014 & ~new_n4018;
  assign new_n4020 = ~new_n4013 & ~new_n4019;
  assign new_n4021 = ~new_n4007 & new_n4020;
  assign new_n4022 = ~new_n4006 & ~new_n4021;
  assign new_n4023 = ~new_n3997 & ~new_n4022;
  assign new_n4024 = ~new_n3996 & ~new_n4023;
  assign new_n4025 = ~new_n3989 & ~new_n4024;
  assign new_n4026 = ~new_n3988 & ~new_n4025;
  assign new_n4027 = ~new_n3728 & new_n4026;
  assign new_n4028 = new_n3728 & ~new_n4026;
  assign new_n4029 = n6877 & n8065;
  assign new_n4030 = ~new_n3783 & ~new_n3786;
  assign new_n4031 = ~new_n3782 & ~new_n4030;
  assign new_n4032 = n9400 & n10439;
  assign new_n4033 = n2464 & n8595;
  assign new_n4034 = ~new_n4032 & ~new_n4033;
  assign new_n4035 = new_n4032 & new_n4033;
  assign new_n4036 = ~new_n4034 & ~new_n4035;
  assign new_n4037 = n6126 & n11311;
  assign new_n4038 = n3719 & n4203;
  assign new_n4039 = n3602 & n4187;
  assign new_n4040 = ~new_n4038 & ~new_n4039;
  assign new_n4041 = new_n4038 & new_n4039;
  assign new_n4042 = ~new_n4040 & ~new_n4041;
  assign new_n4043 = new_n4037 & new_n4042;
  assign new_n4044 = ~new_n4037 & ~new_n4042;
  assign new_n4045 = ~new_n4043 & ~new_n4044;
  assign new_n4046 = new_n3770 & ~new_n3773;
  assign new_n4047 = ~new_n3774 & ~new_n4046;
  assign new_n4048 = ~new_n4045 & ~new_n4047;
  assign new_n4049 = new_n4045 & new_n4047;
  assign new_n4050 = ~new_n4048 & ~new_n4049;
  assign new_n4051 = new_n4036 & ~new_n4050;
  assign new_n4052 = ~new_n4036 & new_n4050;
  assign new_n4053 = ~new_n4051 & ~new_n4052;
  assign new_n4054 = ~new_n3768 & ~new_n3778;
  assign new_n4055 = ~new_n3767 & ~new_n4054;
  assign new_n4056 = new_n4053 & new_n4055;
  assign new_n4057 = ~new_n4053 & ~new_n4055;
  assign new_n4058 = ~new_n4056 & ~new_n4057;
  assign new_n4059 = ~new_n4031 & ~new_n4058;
  assign new_n4060 = new_n4031 & new_n4058;
  assign new_n4061 = ~new_n4059 & ~new_n4060;
  assign new_n4062 = new_n4029 & new_n4061;
  assign new_n4063 = ~new_n4029 & ~new_n4061;
  assign new_n4064 = ~new_n4062 & ~new_n4063;
  assign new_n4065 = new_n3790 & new_n4064;
  assign new_n4066 = ~new_n3790 & ~new_n4064;
  assign new_n4067 = ~new_n4065 & ~new_n4066;
  assign new_n4068 = ~new_n3917 & ~new_n3984;
  assign new_n4069 = ~new_n3916 & ~new_n4068;
  assign new_n4070 = ~new_n4067 & new_n4069;
  assign new_n4071 = new_n4067 & ~new_n4069;
  assign new_n4072 = ~new_n4070 & ~new_n4071;
  assign new_n4073 = n6359 & n7236;
  assign new_n4074 = ~new_n3937 & new_n3941;
  assign new_n4075 = ~new_n3938 & ~new_n4074;
  assign new_n4076 = n217 & n8384;
  assign new_n4077 = n3992 & n6611;
  assign new_n4078 = ~new_n4076 & ~new_n4077;
  assign new_n4079 = new_n4076 & new_n4077;
  assign new_n4080 = ~new_n4078 & ~new_n4079;
  assign new_n4081 = n4086 & n6358;
  assign new_n4082 = new_n3926 & ~new_n3928;
  assign new_n4083 = ~new_n3929 & ~new_n4082;
  assign new_n4084 = ~new_n4081 & new_n4083;
  assign new_n4085 = new_n4081 & ~new_n4083;
  assign new_n4086_1 = n405 & n5198;
  assign new_n4087 = n1471 & n8433;
  assign new_n4088_1 = ~new_n4086_1 & ~new_n4087;
  assign new_n4089 = new_n4086_1 & new_n4087;
  assign new_n4090 = ~new_n4088_1 & ~new_n4089;
  assign new_n4091 = ~new_n4085 & ~new_n4090;
  assign new_n4092 = ~new_n4084 & new_n4091;
  assign new_n4093 = ~new_n4084 & ~new_n4085;
  assign new_n4094_1 = new_n4090 & ~new_n4093;
  assign new_n4095 = ~new_n4092 & ~new_n4094_1;
  assign new_n4096 = new_n4080 & ~new_n4095;
  assign new_n4097 = ~new_n4080 & new_n4095;
  assign new_n4098 = ~new_n4096 & ~new_n4097;
  assign new_n4099 = ~new_n3924 & ~new_n3933;
  assign new_n4100 = ~new_n3923 & ~new_n4099;
  assign new_n4101 = new_n4098 & new_n4100;
  assign new_n4102 = ~new_n4098 & ~new_n4100;
  assign new_n4103 = ~new_n4101 & ~new_n4102;
  assign new_n4104 = new_n4075 & ~new_n4103;
  assign new_n4105 = ~new_n4075 & new_n4103;
  assign new_n4106 = ~new_n4104 & ~new_n4105;
  assign new_n4107 = new_n4073 & new_n4106;
  assign new_n4108 = ~new_n4073 & ~new_n4106;
  assign new_n4109 = ~new_n4107 & ~new_n4108;
  assign new_n4110 = new_n3945 & new_n4109;
  assign new_n4111 = ~new_n3945 & ~new_n4109;
  assign new_n4112 = ~new_n4110 & ~new_n4111;
  assign new_n4113 = n503 & n4805;
  assign new_n4114 = ~new_n3967 & ~new_n3970;
  assign new_n4115 = ~new_n3966 & ~new_n4114;
  assign new_n4116 = n4970 & n11478;
  assign new_n4117 = n5283 & n7610;
  assign new_n4118 = ~new_n4116 & ~new_n4117;
  assign new_n4119 = new_n4116 & new_n4117;
  assign new_n4120 = ~new_n4118 & ~new_n4119;
  assign new_n4121 = n137 & n4826;
  assign new_n4122 = n6294 & n7733;
  assign new_n4123 = n6797 & n12925;
  assign new_n4124 = ~new_n4122 & ~new_n4123;
  assign new_n4125 = new_n4122 & new_n4123;
  assign new_n4126 = ~new_n4124 & ~new_n4125;
  assign new_n4127 = new_n4121 & new_n4126;
  assign new_n4128 = ~new_n4121 & ~new_n4126;
  assign new_n4129 = ~new_n4127 & ~new_n4128;
  assign new_n4130 = new_n3955 & ~new_n3957;
  assign new_n4131 = ~new_n3958 & ~new_n4130;
  assign new_n4132 = ~new_n4129 & ~new_n4131;
  assign new_n4133 = new_n4129 & new_n4131;
  assign new_n4134 = ~new_n4132 & ~new_n4133;
  assign new_n4135 = new_n4120 & ~new_n4134;
  assign new_n4136 = ~new_n4120 & new_n4134;
  assign new_n4137 = ~new_n4135 & ~new_n4136;
  assign new_n4138 = ~new_n3953 & ~new_n3962;
  assign new_n4139 = ~new_n3952 & ~new_n4138;
  assign new_n4140 = new_n4137 & new_n4139;
  assign new_n4141_1 = ~new_n4137 & ~new_n4139;
  assign new_n4142 = ~new_n4140 & ~new_n4141_1;
  assign new_n4143 = ~new_n4115 & ~new_n4142;
  assign new_n4144 = new_n4115 & new_n4142;
  assign new_n4145 = ~new_n4143 & ~new_n4144;
  assign new_n4146 = new_n4113 & new_n4145;
  assign new_n4147 = ~new_n4113 & ~new_n4145;
  assign new_n4148 = ~new_n4146 & ~new_n4147;
  assign new_n4149 = new_n3974 & new_n4148;
  assign new_n4150 = ~new_n3974 & ~new_n4148;
  assign new_n4151 = ~new_n4149 & ~new_n4150;
  assign new_n4152 = new_n4112 & new_n4151;
  assign new_n4153 = ~new_n4112 & ~new_n4151;
  assign new_n4154 = ~new_n4152 & ~new_n4153;
  assign new_n4155_1 = new_n3947 & ~new_n3980;
  assign new_n4156 = ~new_n3979 & ~new_n4155_1;
  assign new_n4157 = ~new_n4154 & ~new_n4156;
  assign new_n4158 = new_n4154 & new_n4156;
  assign new_n4159_1 = ~new_n4157 & ~new_n4158;
  assign new_n4160 = new_n4072 & ~new_n4159_1;
  assign new_n4161 = ~new_n4072 & new_n4159_1;
  assign new_n4162 = ~new_n4160 & ~new_n4161;
  assign new_n4163 = ~new_n4028 & ~new_n4162;
  assign new_n4164 = ~new_n4027 & ~new_n4163;
  assign new_n4165 = ~new_n3726 & ~new_n4164;
  assign new_n4166 = new_n3726 & new_n4164;
  assign new_n4167 = ~new_n4165 & ~new_n4166;
  assign new_n4168 = ~new_n4062 & ~new_n4065;
  assign new_n4169 = ~new_n4052 & ~new_n4055;
  assign new_n4170 = ~new_n4035 & ~new_n4169;
  assign new_n4171 = ~new_n4051 & new_n4170;
  assign new_n4172 = new_n4035 & new_n4169;
  assign new_n4173 = ~new_n4171 & ~new_n4172;
  assign new_n4174 = ~new_n4044 & ~new_n4047;
  assign new_n4175 = ~new_n4043 & ~new_n4174;
  assign new_n4176 = n2464 & n10439;
  assign new_n4177 = n6877 & n10391;
  assign new_n4178 = n8065 & n9400;
  assign new_n4179 = ~new_n4177 & ~new_n4178;
  assign new_n4180 = new_n4177 & new_n4178;
  assign new_n4181 = ~new_n4179 & ~new_n4180;
  assign new_n4182 = new_n4176 & ~new_n4181;
  assign new_n4183 = ~new_n4176 & new_n4181;
  assign new_n4184 = ~new_n4182 & ~new_n4183;
  assign new_n4185 = ~new_n4175 & ~new_n4184;
  assign new_n4186 = new_n4175 & new_n4184;
  assign new_n4187_1 = ~new_n4185 & ~new_n4186;
  assign new_n4188 = n8595 & n11311;
  assign new_n4189_1 = new_n4041 & new_n4188;
  assign new_n4190_1 = ~new_n4041 & ~new_n4188;
  assign new_n4191 = ~new_n4189_1 & ~new_n4190_1;
  assign new_n4192 = n3602 & n4203;
  assign new_n4193 = n4187 & n6126;
  assign new_n4194 = n3719 & n12753;
  assign new_n4195 = ~new_n4193 & ~new_n4194;
  assign new_n4196 = new_n4193 & new_n4194;
  assign new_n4197 = ~new_n4195 & ~new_n4196;
  assign new_n4198 = ~new_n4192 & ~new_n4197;
  assign new_n4199 = new_n4192 & new_n4197;
  assign new_n4200 = ~new_n4198 & ~new_n4199;
  assign new_n4201 = new_n4191 & ~new_n4200;
  assign new_n4202 = ~new_n4191 & new_n4200;
  assign new_n4203_1 = ~new_n4201 & ~new_n4202;
  assign new_n4204 = new_n4187_1 & new_n4203_1;
  assign new_n4205 = ~new_n4187_1 & ~new_n4203_1;
  assign new_n4206 = ~new_n4204 & ~new_n4205;
  assign new_n4207 = ~new_n4173 & new_n4206;
  assign new_n4208 = new_n4173 & ~new_n4206;
  assign new_n4209 = ~new_n4207 & ~new_n4208;
  assign new_n4210 = ~new_n4059 & ~new_n4209;
  assign new_n4211 = new_n4059 & new_n4209;
  assign new_n4212 = ~new_n4210 & ~new_n4211;
  assign new_n4213 = ~new_n4168 & new_n4212;
  assign new_n4214 = new_n4168 & ~new_n4212;
  assign new_n4215 = ~new_n4213 & ~new_n4214;
  assign new_n4216 = ~new_n4136 & ~new_n4139;
  assign new_n4217 = ~new_n4119 & ~new_n4216;
  assign new_n4218 = ~new_n4135 & new_n4217;
  assign new_n4219 = new_n4119 & new_n4216;
  assign new_n4220 = ~new_n4218 & ~new_n4219;
  assign new_n4221 = ~new_n4128 & ~new_n4131;
  assign new_n4222 = ~new_n4127 & ~new_n4221;
  assign new_n4223 = n4805 & n10965;
  assign new_n4224 = n4970 & n5283;
  assign new_n4225 = n503 & n11478;
  assign new_n4226_1 = ~new_n4224 & ~new_n4225;
  assign new_n4227 = new_n4224 & new_n4225;
  assign new_n4228 = ~new_n4226_1 & ~new_n4227;
  assign new_n4229 = new_n4223 & ~new_n4228;
  assign new_n4230_1 = ~new_n4223 & new_n4228;
  assign new_n4231 = ~new_n4229 & ~new_n4230_1;
  assign new_n4232 = new_n4222 & new_n4231;
  assign new_n4233 = n137 & n7610;
  assign new_n4234 = ~new_n4125 & ~new_n4233;
  assign new_n4235 = new_n4125 & new_n4233;
  assign new_n4236 = ~new_n4234 & ~new_n4235;
  assign new_n4237 = n3146 & n12925;
  assign new_n4238 = n4826 & n6294;
  assign new_n4239 = n6797 & n7733;
  assign new_n4240 = ~new_n4238 & ~new_n4239;
  assign new_n4241 = new_n4238 & new_n4239;
  assign new_n4242 = ~new_n4240 & ~new_n4241;
  assign new_n4243 = new_n4237 & ~new_n4242;
  assign new_n4244 = ~new_n4237 & new_n4242;
  assign new_n4245 = ~new_n4243 & ~new_n4244;
  assign new_n4246 = new_n4236 & new_n4245;
  assign new_n4247 = ~new_n4236 & ~new_n4245;
  assign new_n4248 = ~new_n4246 & ~new_n4247;
  assign new_n4249 = new_n4232 & new_n4248;
  assign new_n4250 = ~new_n4222 & ~new_n4231;
  assign new_n4251 = new_n4248 & ~new_n4250;
  assign new_n4252 = ~new_n4232 & ~new_n4251;
  assign new_n4253 = ~new_n4249 & ~new_n4252;
  assign new_n4254 = ~new_n4248 & new_n4250;
  assign new_n4255 = ~new_n4253 & ~new_n4254;
  assign new_n4256 = ~new_n4220 & ~new_n4255;
  assign new_n4257 = new_n4220 & new_n4255;
  assign new_n4258 = ~new_n4256 & ~new_n4257;
  assign new_n4259 = ~new_n4143 & new_n4258;
  assign new_n4260 = new_n4143 & ~new_n4258;
  assign new_n4261 = ~new_n4259 & ~new_n4260;
  assign new_n4262 = ~new_n4146 & ~new_n4149;
  assign new_n4263 = ~new_n4261 & new_n4262;
  assign new_n4264 = new_n4261 & ~new_n4262;
  assign new_n4265 = ~new_n4263 & ~new_n4264;
  assign new_n4266 = ~new_n4097 & ~new_n4100;
  assign new_n4267 = ~new_n4079 & ~new_n4266;
  assign new_n4268 = ~new_n4096 & new_n4267;
  assign new_n4269 = new_n4079 & new_n4266;
  assign new_n4270 = ~new_n4268 & ~new_n4269;
  assign new_n4271 = ~new_n4084 & ~new_n4091;
  assign new_n4272 = n7236 & n11296;
  assign new_n4273 = n6611 & n8384;
  assign new_n4274 = n3992 & n6359;
  assign new_n4275 = ~new_n4273 & ~new_n4274;
  assign new_n4276 = new_n4273 & new_n4274;
  assign new_n4277 = ~new_n4275 & ~new_n4276;
  assign new_n4278 = new_n4272 & ~new_n4277;
  assign new_n4279 = ~new_n4272 & new_n4277;
  assign new_n4280 = ~new_n4278 & ~new_n4279;
  assign new_n4281 = new_n4271 & ~new_n4280;
  assign new_n4282 = ~new_n4271 & new_n4280;
  assign new_n4283 = ~new_n4281 & ~new_n4282;
  assign new_n4284 = n217 & n6358;
  assign new_n4285 = ~new_n4089 & ~new_n4284;
  assign new_n4286 = new_n4089 & new_n4284;
  assign new_n4287 = ~new_n4285 & ~new_n4286;
  assign new_n4288 = n7646 & n8433;
  assign new_n4289 = n4086 & n5198;
  assign new_n4290 = n405 & n1471;
  assign new_n4291 = ~new_n4289 & ~new_n4290;
  assign new_n4292 = new_n4289 & new_n4290;
  assign new_n4293 = ~new_n4291 & ~new_n4292;
  assign new_n4294 = new_n4288 & ~new_n4293;
  assign new_n4295 = ~new_n4288 & new_n4293;
  assign new_n4296 = ~new_n4294 & ~new_n4295;
  assign new_n4297 = new_n4287 & ~new_n4296;
  assign new_n4298 = ~new_n4287 & new_n4296;
  assign new_n4299 = ~new_n4297 & ~new_n4298;
  assign new_n4300_1 = ~new_n4283 & ~new_n4299;
  assign new_n4301 = new_n4283 & new_n4299;
  assign new_n4302 = ~new_n4300_1 & ~new_n4301;
  assign new_n4303 = new_n4270 & ~new_n4302;
  assign new_n4304 = ~new_n4270 & new_n4302;
  assign new_n4305 = ~new_n4303 & ~new_n4304;
  assign new_n4306 = ~new_n4104 & new_n4305;
  assign new_n4307 = new_n4104 & ~new_n4305;
  assign new_n4308 = ~new_n4306 & ~new_n4307;
  assign new_n4309 = ~new_n4107 & ~new_n4110;
  assign new_n4310 = ~new_n4308 & new_n4309;
  assign new_n4311 = new_n4308 & ~new_n4309;
  assign new_n4312_1 = ~new_n4310 & ~new_n4311;
  assign new_n4313 = new_n4265 & new_n4312_1;
  assign new_n4314 = ~new_n4265 & ~new_n4312_1;
  assign new_n4315 = ~new_n4313 & ~new_n4314;
  assign new_n4316 = ~new_n4153 & ~new_n4156;
  assign new_n4317 = ~new_n4152 & ~new_n4316;
  assign new_n4318 = new_n4315 & new_n4317;
  assign new_n4319 = ~new_n4315 & ~new_n4317;
  assign new_n4320 = ~new_n4318 & ~new_n4319;
  assign new_n4321 = new_n4215 & ~new_n4320;
  assign new_n4322 = ~new_n4215 & new_n4320;
  assign new_n4323 = ~new_n4321 & ~new_n4322;
  assign new_n4324 = ~new_n4071 & new_n4159_1;
  assign new_n4325 = ~new_n4070 & ~new_n4324;
  assign new_n4326_1 = ~new_n4323 & new_n4325;
  assign new_n4327 = new_n4323 & ~new_n4325;
  assign new_n4328 = ~new_n4326_1 & ~new_n4327;
  assign new_n4329 = new_n4167 & ~new_n4328;
  assign new_n4330 = ~new_n4167 & new_n4328;
  assign n844 = ~new_n4329 & ~new_n4330;
  assign new_n4332 = n3932 & n6687;
  assign new_n4333_1 = n1798 & n2564;
  assign new_n4334 = new_n4332 & new_n4333_1;
  assign new_n4335 = n1798 & n4189;
  assign new_n4336 = n2564 & n3932;
  assign new_n4337 = n6687 & n12591;
  assign new_n4338 = ~new_n4336 & ~new_n4337;
  assign new_n4339 = new_n4336 & new_n4337;
  assign new_n4340 = ~new_n4338 & ~new_n4339;
  assign new_n4341 = new_n4335 & ~new_n4340;
  assign new_n4342 = ~new_n4335 & new_n4340;
  assign new_n4343 = ~new_n4341 & ~new_n4342;
  assign new_n4344 = new_n4334 & ~new_n4343;
  assign new_n4345 = n6687 & n7456;
  assign new_n4346 = new_n4335 & ~new_n4338;
  assign new_n4347 = ~new_n4339 & ~new_n4346;
  assign new_n4348 = ~new_n4345 & new_n4347;
  assign new_n4349 = new_n4345 & ~new_n4347;
  assign new_n4350 = ~new_n4348 & ~new_n4349;
  assign new_n4351 = n1798 & n6770;
  assign new_n4352 = n2564 & n12591;
  assign new_n4353 = n3932 & n4189;
  assign new_n4354 = ~new_n4352 & ~new_n4353;
  assign new_n4355 = new_n4352 & new_n4353;
  assign new_n4356 = ~new_n4354 & ~new_n4355;
  assign new_n4357 = new_n4351 & ~new_n4356;
  assign new_n4358 = ~new_n4351 & new_n4356;
  assign new_n4359 = ~new_n4357 & ~new_n4358;
  assign new_n4360 = ~new_n4350 & new_n4359;
  assign new_n4361 = new_n4350 & ~new_n4359;
  assign new_n4362 = ~new_n4360 & ~new_n4361;
  assign new_n4363 = new_n4344 & new_n4362;
  assign new_n4364 = ~new_n4344 & ~new_n4362;
  assign new_n4365 = ~new_n4363 & ~new_n4364;
  assign new_n4366 = ~new_n4334 & new_n4343;
  assign new_n4367 = ~new_n4344 & ~new_n4366;
  assign new_n4368 = n5645 & n12391;
  assign new_n4369 = n1067 & n12069;
  assign new_n4370_1 = new_n4368 & new_n4369;
  assign new_n4371 = n8665 & n12069;
  assign new_n4372 = n1067 & n12391;
  assign new_n4373 = n5645 & n7891;
  assign new_n4374 = ~new_n4372 & ~new_n4373;
  assign new_n4375 = new_n4372 & new_n4373;
  assign new_n4376 = ~new_n4374 & ~new_n4375;
  assign new_n4377 = new_n4371 & ~new_n4376;
  assign new_n4378_1 = ~new_n4371 & new_n4376;
  assign new_n4379 = ~new_n4377 & ~new_n4378_1;
  assign new_n4380 = ~new_n4370_1 & new_n4379;
  assign new_n4381 = new_n4370_1 & ~new_n4379;
  assign new_n4382 = ~new_n4380 & ~new_n4381;
  assign new_n4383 = n10898 & n11222;
  assign new_n4384 = n11153 & n11876;
  assign new_n4385 = new_n4383 & new_n4384;
  assign new_n4386 = n5314 & n11876;
  assign new_n4387 = n10898 & n11153;
  assign new_n4388 = n3754 & n11222;
  assign new_n4389 = ~new_n4387 & ~new_n4388;
  assign new_n4390 = new_n4387 & new_n4388;
  assign new_n4391 = ~new_n4389 & ~new_n4390;
  assign new_n4392 = new_n4386 & ~new_n4391;
  assign new_n4393 = ~new_n4386 & new_n4391;
  assign new_n4394 = ~new_n4392 & ~new_n4393;
  assign new_n4395 = new_n4385 & ~new_n4394;
  assign new_n4396 = ~new_n4385 & new_n4394;
  assign new_n4397_1 = ~new_n4395 & ~new_n4396;
  assign new_n4398 = n5645 & n12069;
  assign new_n4399 = n11222 & n11876;
  assign new_n4400 = new_n4398 & new_n4399;
  assign new_n4401 = ~new_n4368 & ~new_n4369;
  assign new_n4402 = ~new_n4370_1 & ~new_n4401;
  assign new_n4403 = ~new_n4400 & ~new_n4402;
  assign new_n4404 = new_n4400 & new_n4402;
  assign new_n4405 = ~new_n4383 & ~new_n4384;
  assign new_n4406 = ~new_n4385 & ~new_n4405;
  assign new_n4407 = ~new_n4404 & ~new_n4406;
  assign new_n4408 = ~new_n4403 & ~new_n4407;
  assign new_n4409 = new_n4397_1 & new_n4408;
  assign new_n4410 = ~new_n4397_1 & ~new_n4408;
  assign new_n4411 = ~new_n4409 & ~new_n4410;
  assign new_n4412 = ~new_n4382 & new_n4411;
  assign new_n4413 = new_n4382 & ~new_n4411;
  assign new_n4414 = ~new_n4412 & ~new_n4413;
  assign new_n4415 = n8336 & n9640;
  assign new_n4416 = n6703 & n10928;
  assign new_n4417 = new_n4415 & new_n4416;
  assign new_n4418 = n6703 & n6986;
  assign new_n4419 = n9640 & n10928;
  assign new_n4420 = n3022 & n8336;
  assign new_n4421 = ~new_n4419 & ~new_n4420;
  assign new_n4422 = new_n4419 & new_n4420;
  assign new_n4423 = ~new_n4421 & ~new_n4422;
  assign new_n4424 = new_n4418 & ~new_n4423;
  assign new_n4425 = ~new_n4418 & new_n4423;
  assign new_n4426 = ~new_n4424 & ~new_n4425;
  assign new_n4427 = new_n4417 & ~new_n4426;
  assign new_n4428 = ~new_n4417 & new_n4426;
  assign new_n4429 = ~new_n4427 & ~new_n4428;
  assign new_n4430 = n6703 & n8336;
  assign new_n4431 = ~new_n4398 & ~new_n4399;
  assign new_n4432 = ~new_n4400 & ~new_n4431;
  assign new_n4433 = new_n4430 & new_n4432;
  assign new_n4434 = ~new_n4415 & ~new_n4416;
  assign new_n4435 = ~new_n4417 & ~new_n4434;
  assign new_n4436_1 = new_n4433 & new_n4435;
  assign new_n4437 = ~new_n4433 & ~new_n4435;
  assign new_n4438 = ~new_n4403 & ~new_n4404;
  assign new_n4439 = ~new_n4406 & new_n4438;
  assign new_n4440 = new_n4406 & ~new_n4438;
  assign new_n4441 = ~new_n4439 & ~new_n4440;
  assign new_n4442 = ~new_n4437 & ~new_n4441;
  assign new_n4443 = ~new_n4436_1 & ~new_n4442;
  assign new_n4444 = ~new_n4429 & new_n4443;
  assign new_n4445 = new_n4429 & ~new_n4443;
  assign new_n4446 = ~new_n4444 & ~new_n4445;
  assign new_n4447 = new_n4414 & new_n4446;
  assign new_n4448 = ~new_n4414 & ~new_n4446;
  assign new_n4449 = ~new_n4447 & ~new_n4448;
  assign new_n4450 = new_n4367 & ~new_n4449;
  assign new_n4451 = ~new_n4367 & new_n4449;
  assign new_n4452 = n1798 & n6687;
  assign new_n4453 = ~new_n4430 & ~new_n4432;
  assign new_n4454 = ~new_n4433 & ~new_n4453;
  assign new_n4455 = new_n4452 & new_n4454;
  assign new_n4456 = ~new_n4332 & ~new_n4333_1;
  assign new_n4457 = ~new_n4334 & ~new_n4456;
  assign new_n4458 = new_n4455 & new_n4457;
  assign new_n4459 = ~new_n4455 & ~new_n4457;
  assign new_n4460 = ~new_n4436_1 & ~new_n4437;
  assign new_n4461 = ~new_n4441 & new_n4460;
  assign new_n4462 = new_n4441 & ~new_n4460;
  assign new_n4463 = ~new_n4461 & ~new_n4462;
  assign new_n4464 = ~new_n4459 & new_n4463;
  assign new_n4465 = ~new_n4458 & ~new_n4464;
  assign new_n4466 = ~new_n4451 & ~new_n4465;
  assign new_n4467 = ~new_n4450 & ~new_n4466;
  assign new_n4468 = new_n4365 & ~new_n4467;
  assign new_n4469 = ~new_n4365 & new_n4467;
  assign new_n4470 = ~new_n4468 & ~new_n4469;
  assign new_n4471 = n8336 & n11023;
  assign new_n4472 = new_n4418 & ~new_n4421;
  assign new_n4473 = ~new_n4422 & ~new_n4472;
  assign new_n4474 = ~new_n4471 & new_n4473;
  assign new_n4475 = new_n4471 & ~new_n4473;
  assign new_n4476 = ~new_n4474 & ~new_n4475;
  assign new_n4477 = n2226 & n6703;
  assign new_n4478 = n3022 & n10928;
  assign new_n4479 = n6986 & n9640;
  assign new_n4480 = ~new_n4478 & ~new_n4479;
  assign new_n4481 = new_n4478 & new_n4479;
  assign new_n4482 = ~new_n4480 & ~new_n4481;
  assign new_n4483 = new_n4477 & ~new_n4482;
  assign new_n4484 = ~new_n4477 & new_n4482;
  assign new_n4485 = ~new_n4483 & ~new_n4484;
  assign new_n4486 = ~new_n4476 & new_n4485;
  assign new_n4487 = new_n4476 & ~new_n4485;
  assign new_n4488 = ~new_n4486 & ~new_n4487;
  assign new_n4489 = ~new_n4427 & ~new_n4488;
  assign new_n4490 = new_n4427 & new_n4488;
  assign new_n4491 = ~new_n4489 & ~new_n4490;
  assign new_n4492 = ~new_n4414 & ~new_n4444;
  assign new_n4493 = ~new_n4445 & ~new_n4492;
  assign new_n4494 = new_n4491 & ~new_n4493;
  assign new_n4495 = ~new_n4491 & new_n4493;
  assign new_n4496 = ~new_n4494 & ~new_n4495;
  assign new_n4497 = n11922 & n12069;
  assign new_n4498 = new_n4371 & ~new_n4374;
  assign new_n4499_1 = ~new_n4375 & ~new_n4498;
  assign new_n4500 = new_n4497 & ~new_n4499_1;
  assign new_n4501 = ~new_n4497 & new_n4499_1;
  assign new_n4502 = ~new_n4500 & ~new_n4501;
  assign new_n4503 = n5645 & n7160;
  assign new_n4504 = n1067 & n7891;
  assign new_n4505 = n8665 & n12391;
  assign new_n4506 = ~new_n4504 & ~new_n4505;
  assign new_n4507 = new_n4504 & new_n4505;
  assign new_n4508 = ~new_n4506 & ~new_n4507;
  assign new_n4509 = new_n4503 & ~new_n4508;
  assign new_n4510 = ~new_n4503 & new_n4508;
  assign new_n4511 = ~new_n4509 & ~new_n4510;
  assign new_n4512 = ~new_n4502 & ~new_n4511;
  assign new_n4513 = new_n4502 & new_n4511;
  assign new_n4514 = ~new_n4512 & ~new_n4513;
  assign new_n4515 = ~new_n4381 & new_n4514;
  assign new_n4516_1 = new_n4381 & ~new_n4514;
  assign new_n4517 = ~new_n4515 & ~new_n4516_1;
  assign new_n4518 = n2749 & n11222;
  assign new_n4519 = new_n4386 & ~new_n4389;
  assign new_n4520 = ~new_n4390 & ~new_n4519;
  assign new_n4521 = new_n4518 & ~new_n4520;
  assign new_n4522 = ~new_n4518 & new_n4520;
  assign new_n4523 = ~new_n4521 & ~new_n4522;
  assign new_n4524 = n5314 & n10898;
  assign new_n4525 = n3754 & n11153;
  assign new_n4526 = n996 & n11876;
  assign new_n4527 = ~new_n4525 & ~new_n4526;
  assign new_n4528 = new_n4525 & new_n4526;
  assign new_n4529 = ~new_n4527 & ~new_n4528;
  assign new_n4530 = new_n4524 & ~new_n4529;
  assign new_n4531 = ~new_n4524 & new_n4529;
  assign new_n4532 = ~new_n4530 & ~new_n4531;
  assign new_n4533 = ~new_n4523 & ~new_n4532;
  assign new_n4534 = new_n4523 & new_n4532;
  assign new_n4535 = ~new_n4533 & ~new_n4534;
  assign new_n4536 = new_n4395 & ~new_n4535;
  assign new_n4537 = ~new_n4395 & new_n4535;
  assign new_n4538 = ~new_n4536 & ~new_n4537;
  assign new_n4539 = new_n4517 & new_n4538;
  assign new_n4540 = ~new_n4517 & ~new_n4538;
  assign new_n4541 = ~new_n4539 & ~new_n4540;
  assign new_n4542 = new_n4382 & ~new_n4410;
  assign new_n4543 = ~new_n4409 & ~new_n4542;
  assign new_n4544 = new_n4541 & new_n4543;
  assign new_n4545 = ~new_n4541 & ~new_n4543;
  assign new_n4546 = ~new_n4544 & ~new_n4545;
  assign new_n4547 = new_n4496 & ~new_n4546;
  assign new_n4548 = ~new_n4496 & new_n4546;
  assign new_n4549 = ~new_n4547 & ~new_n4548;
  assign new_n4550 = new_n4470 & ~new_n4549;
  assign new_n4551 = ~new_n4470 & new_n4549;
  assign n911 = new_n4550 | new_n4551;
  assign new_n4553_1 = n4921 & n6687;
  assign new_n4554 = n2564 & n9956;
  assign new_n4555 = new_n4553_1 & new_n4554;
  assign new_n4556 = n4189 & n9956;
  assign new_n4557 = n2564 & n4921;
  assign new_n4558 = n6687 & n11917;
  assign new_n4559 = ~new_n4557 & ~new_n4558;
  assign new_n4560 = new_n4557 & new_n4558;
  assign new_n4561 = ~new_n4559 & ~new_n4560;
  assign new_n4562 = new_n4556 & ~new_n4561;
  assign new_n4563 = ~new_n4556 & new_n4561;
  assign new_n4564 = ~new_n4562 & ~new_n4563;
  assign new_n4565 = new_n4555 & ~new_n4564;
  assign new_n4566 = n3842 & n6687;
  assign new_n4567 = new_n4556 & ~new_n4559;
  assign new_n4568 = ~new_n4560 & ~new_n4567;
  assign new_n4569 = ~new_n4566 & new_n4568;
  assign new_n4570 = new_n4566 & ~new_n4568;
  assign new_n4571 = ~new_n4569 & ~new_n4570;
  assign new_n4572 = n6770 & n9956;
  assign new_n4573 = n2564 & n11917;
  assign new_n4574 = n4189 & n4921;
  assign new_n4575 = ~new_n4573 & ~new_n4574;
  assign new_n4576 = new_n4573 & new_n4574;
  assign new_n4577 = ~new_n4575 & ~new_n4576;
  assign new_n4578 = new_n4572 & ~new_n4577;
  assign new_n4579 = ~new_n4572 & new_n4577;
  assign new_n4580 = ~new_n4578 & ~new_n4579;
  assign new_n4581 = ~new_n4571 & new_n4580;
  assign new_n4582 = new_n4571 & ~new_n4580;
  assign new_n4583 = ~new_n4581 & ~new_n4582;
  assign new_n4584 = new_n4565 & new_n4583;
  assign new_n4585 = n2577 & n6687;
  assign new_n4586 = ~new_n4569 & ~new_n4580;
  assign new_n4587 = ~new_n4570 & ~new_n4586;
  assign new_n4588 = new_n4585 & ~new_n4587;
  assign new_n4589 = ~new_n4585 & new_n4587;
  assign new_n4590 = ~new_n4588 & ~new_n4589;
  assign new_n4591 = n2564 & n3842;
  assign new_n4592 = new_n4572 & ~new_n4575;
  assign new_n4593 = ~new_n4576 & ~new_n4592;
  assign new_n4594 = new_n4591 & ~new_n4593;
  assign new_n4595 = ~new_n4591 & new_n4593;
  assign new_n4596 = ~new_n4594 & ~new_n4595;
  assign new_n4597 = n4921 & n6770;
  assign new_n4598 = n4189 & n11917;
  assign new_n4599 = n9920 & n9956;
  assign new_n4600 = ~new_n4598 & ~new_n4599;
  assign new_n4601 = new_n4598 & new_n4599;
  assign new_n4602 = ~new_n4600 & ~new_n4601;
  assign new_n4603 = new_n4597 & ~new_n4602;
  assign new_n4604 = ~new_n4597 & new_n4602;
  assign new_n4605 = ~new_n4603 & ~new_n4604;
  assign new_n4606 = ~new_n4596 & ~new_n4605;
  assign new_n4607 = new_n4596 & new_n4605;
  assign new_n4608 = ~new_n4606 & ~new_n4607;
  assign new_n4609 = ~new_n4590 & ~new_n4608;
  assign new_n4610 = new_n4590 & new_n4608;
  assign new_n4611 = ~new_n4609 & ~new_n4610;
  assign new_n4612 = new_n4584 & ~new_n4611;
  assign new_n4613 = ~new_n4584 & new_n4611;
  assign new_n4614 = ~new_n4612 & ~new_n4613;
  assign new_n4615 = ~new_n4565 & ~new_n4583;
  assign new_n4616 = ~new_n4584 & ~new_n4615;
  assign new_n4617 = n3602 & n8336;
  assign new_n4618 = n3719 & n10928;
  assign new_n4619 = new_n4617 & new_n4618;
  assign new_n4620 = n3719 & n6986;
  assign new_n4621 = n3602 & n10928;
  assign new_n4622 = n6126 & n8336;
  assign new_n4623 = ~new_n4621 & ~new_n4622;
  assign new_n4624 = new_n4621 & new_n4622;
  assign new_n4625 = ~new_n4623 & ~new_n4624;
  assign new_n4626 = new_n4620 & ~new_n4625;
  assign new_n4627 = ~new_n4620 & new_n4625;
  assign new_n4628 = ~new_n4626 & ~new_n4627;
  assign new_n4629 = new_n4619 & ~new_n4628;
  assign new_n4630 = n8336 & n8595;
  assign new_n4631 = new_n4620 & ~new_n4623;
  assign new_n4632 = ~new_n4624 & ~new_n4631;
  assign new_n4633 = ~new_n4630 & new_n4632;
  assign new_n4634_1 = new_n4630 & ~new_n4632;
  assign new_n4635 = ~new_n4633 & ~new_n4634_1;
  assign new_n4636 = n2226 & n3719;
  assign new_n4637 = n6126 & n10928;
  assign new_n4638 = n3602 & n6986;
  assign new_n4639 = ~new_n4637 & ~new_n4638;
  assign new_n4640 = new_n4637 & new_n4638;
  assign new_n4641 = ~new_n4639 & ~new_n4640;
  assign new_n4642 = new_n4636 & ~new_n4641;
  assign new_n4643 = ~new_n4636 & new_n4641;
  assign new_n4644 = ~new_n4642 & ~new_n4643;
  assign new_n4645 = ~new_n4635 & new_n4644;
  assign new_n4646 = new_n4635 & ~new_n4644;
  assign new_n4647 = ~new_n4645 & ~new_n4646;
  assign new_n4648 = ~new_n4629 & ~new_n4647;
  assign new_n4649 = new_n4629 & new_n4647;
  assign new_n4650 = ~new_n4648 & ~new_n4649;
  assign new_n4651 = n7733 & n12069;
  assign new_n4652 = n12391 & n12925;
  assign new_n4653 = new_n4651 & new_n4652;
  assign new_n4654 = n7891 & n12925;
  assign new_n4655 = n7733 & n12391;
  assign new_n4656 = n4826 & n12069;
  assign new_n4657 = ~new_n4655 & ~new_n4656;
  assign new_n4658 = new_n4655 & new_n4656;
  assign new_n4659 = ~new_n4657 & ~new_n4658;
  assign new_n4660 = new_n4654 & ~new_n4659;
  assign new_n4661 = ~new_n4654 & new_n4659;
  assign new_n4662 = ~new_n4660 & ~new_n4661;
  assign new_n4663 = new_n4653 & ~new_n4662;
  assign new_n4664 = n7610 & n12069;
  assign new_n4665 = new_n4654 & ~new_n4657;
  assign new_n4666 = ~new_n4658 & ~new_n4665;
  assign new_n4667 = ~new_n4664 & new_n4666;
  assign new_n4668 = new_n4664 & ~new_n4666;
  assign new_n4669 = ~new_n4667 & ~new_n4668;
  assign new_n4670 = n7160 & n12925;
  assign new_n4671 = n4826 & n12391;
  assign new_n4672 = n7733 & n7891;
  assign new_n4673 = ~new_n4671 & ~new_n4672;
  assign new_n4674 = new_n4671 & new_n4672;
  assign new_n4675 = ~new_n4673 & ~new_n4674;
  assign new_n4676 = new_n4670 & ~new_n4675;
  assign new_n4677 = ~new_n4670 & new_n4675;
  assign new_n4678 = ~new_n4676 & ~new_n4677;
  assign new_n4679 = ~new_n4669 & new_n4678;
  assign new_n4680 = new_n4669 & ~new_n4678;
  assign new_n4681 = ~new_n4679 & ~new_n4680;
  assign new_n4682 = ~new_n4663 & ~new_n4681;
  assign new_n4683 = new_n4663 & new_n4681;
  assign new_n4684 = ~new_n4682 & ~new_n4683;
  assign new_n4685 = n5314 & n8433;
  assign new_n4686_1 = n4086 & n11222;
  assign new_n4687 = ~new_n4685 & ~new_n4686_1;
  assign new_n4688 = n8433 & n11222;
  assign new_n4689_1 = n4086 & n5314;
  assign new_n4690 = new_n4688 & new_n4689_1;
  assign new_n4691 = ~new_n4687 & ~new_n4690;
  assign new_n4692 = n405 & n11222;
  assign new_n4693 = n8433 & n11153;
  assign new_n4694 = new_n4692 & new_n4693;
  assign new_n4695 = ~new_n4691 & new_n4694;
  assign new_n4696 = n217 & n11222;
  assign new_n4697 = n405 & n11153;
  assign new_n4698 = ~new_n4687 & new_n4697;
  assign new_n4699 = ~new_n4690 & ~new_n4698;
  assign new_n4700 = new_n4696 & ~new_n4699;
  assign new_n4701 = ~new_n4696 & new_n4699;
  assign new_n4702 = ~new_n4700 & ~new_n4701;
  assign new_n4703 = n996 & n8433;
  assign new_n4704 = n4086 & n11153;
  assign new_n4705 = n405 & n5314;
  assign new_n4706 = ~new_n4704 & ~new_n4705;
  assign new_n4707 = new_n4704 & new_n4705;
  assign new_n4708 = ~new_n4706 & ~new_n4707;
  assign new_n4709 = new_n4703 & ~new_n4708;
  assign new_n4710 = ~new_n4703 & new_n4708;
  assign new_n4711 = ~new_n4709 & ~new_n4710;
  assign new_n4712 = ~new_n4702 & ~new_n4711;
  assign new_n4713 = new_n4702 & new_n4711;
  assign new_n4714 = ~new_n4712 & ~new_n4713;
  assign new_n4715 = new_n4695 & ~new_n4714;
  assign new_n4716 = ~new_n4695 & new_n4714;
  assign new_n4717 = ~new_n4715 & ~new_n4716;
  assign new_n4718 = new_n4684 & new_n4717;
  assign new_n4719 = ~new_n4684 & ~new_n4717;
  assign new_n4720 = ~new_n4718 & ~new_n4719;
  assign new_n4721 = n12069 & n12925;
  assign new_n4722_1 = new_n4688 & new_n4721;
  assign new_n4723 = ~new_n4692 & ~new_n4693;
  assign new_n4724 = ~new_n4694 & ~new_n4723;
  assign new_n4725 = new_n4722_1 & new_n4724;
  assign new_n4726 = ~new_n4722_1 & ~new_n4724;
  assign new_n4727 = ~new_n4651 & ~new_n4652;
  assign new_n4728 = ~new_n4653 & ~new_n4727;
  assign new_n4729 = ~new_n4726 & new_n4728;
  assign new_n4730 = ~new_n4725 & ~new_n4729;
  assign new_n4731 = ~new_n4688 & new_n4697;
  assign new_n4732 = ~new_n4687 & new_n4731;
  assign new_n4733_1 = ~new_n4691 & ~new_n4731;
  assign new_n4734 = ~new_n4732 & ~new_n4733_1;
  assign new_n4735 = ~new_n4730 & new_n4734;
  assign new_n4736 = new_n4730 & ~new_n4734;
  assign new_n4737 = ~new_n4653 & new_n4662;
  assign new_n4738 = ~new_n4663 & ~new_n4737;
  assign new_n4739 = ~new_n4736 & new_n4738;
  assign new_n4740 = ~new_n4735 & ~new_n4739;
  assign new_n4741 = new_n4720 & new_n4740;
  assign new_n4742 = ~new_n4720 & ~new_n4740;
  assign new_n4743 = ~new_n4741 & ~new_n4742;
  assign new_n4744 = new_n4650 & ~new_n4743;
  assign new_n4745 = ~new_n4650 & new_n4743;
  assign new_n4746 = ~new_n4744 & ~new_n4745;
  assign new_n4747 = ~new_n4619 & new_n4628;
  assign new_n4748 = ~new_n4629 & ~new_n4747;
  assign new_n4749 = ~new_n4735 & ~new_n4736;
  assign new_n4750 = new_n4738 & new_n4749;
  assign new_n4751 = ~new_n4738 & ~new_n4749;
  assign new_n4752 = ~new_n4750 & ~new_n4751;
  assign new_n4753 = ~new_n4748 & ~new_n4752;
  assign new_n4754 = new_n4748 & new_n4752;
  assign new_n4755 = ~new_n4617 & ~new_n4618;
  assign new_n4756 = ~new_n4619 & ~new_n4755;
  assign new_n4757_1 = ~new_n4725 & ~new_n4726;
  assign new_n4758 = new_n4728 & ~new_n4757_1;
  assign new_n4759 = ~new_n4728 & new_n4757_1;
  assign new_n4760 = ~new_n4758 & ~new_n4759;
  assign new_n4761 = new_n4756 & ~new_n4760;
  assign new_n4762 = ~new_n4756 & new_n4760;
  assign new_n4763 = n3719 & n8336;
  assign new_n4764 = ~new_n4688 & ~new_n4721;
  assign new_n4765 = ~new_n4722_1 & ~new_n4764;
  assign new_n4766 = new_n4763 & new_n4765;
  assign new_n4767 = ~new_n4762 & new_n4766;
  assign new_n4768 = ~new_n4761 & ~new_n4767;
  assign new_n4769 = ~new_n4754 & new_n4768;
  assign new_n4770 = ~new_n4753 & ~new_n4769;
  assign new_n4771 = ~new_n4746 & new_n4770;
  assign new_n4772 = new_n4746 & ~new_n4770;
  assign new_n4773 = ~new_n4771 & ~new_n4772;
  assign new_n4774 = new_n4616 & ~new_n4773;
  assign new_n4775 = ~new_n4616 & new_n4773;
  assign new_n4776 = ~new_n4555 & new_n4564;
  assign new_n4777 = ~new_n4565 & ~new_n4776;
  assign new_n4778 = ~new_n4753 & ~new_n4754;
  assign new_n4779 = new_n4768 & new_n4778;
  assign new_n4780 = ~new_n4768 & ~new_n4778;
  assign new_n4781 = ~new_n4779 & ~new_n4780;
  assign new_n4782 = new_n4777 & ~new_n4781;
  assign new_n4783 = ~new_n4777 & new_n4781;
  assign new_n4784 = n6687 & n9956;
  assign new_n4785 = ~new_n4763 & ~new_n4765;
  assign new_n4786 = ~new_n4766 & ~new_n4785;
  assign new_n4787 = new_n4784 & new_n4786;
  assign new_n4788 = ~new_n4553_1 & ~new_n4554;
  assign new_n4789 = ~new_n4555 & ~new_n4788;
  assign new_n4790 = new_n4787 & new_n4789;
  assign new_n4791 = ~new_n4787 & ~new_n4789;
  assign new_n4792 = ~new_n4761 & ~new_n4762;
  assign new_n4793 = ~new_n4766 & ~new_n4792;
  assign new_n4794 = new_n4766 & new_n4792;
  assign new_n4795 = ~new_n4793 & ~new_n4794;
  assign new_n4796 = ~new_n4791 & new_n4795;
  assign new_n4797 = ~new_n4790 & ~new_n4796;
  assign new_n4798 = ~new_n4783 & ~new_n4797;
  assign new_n4799 = ~new_n4782 & ~new_n4798;
  assign new_n4800 = ~new_n4775 & ~new_n4799;
  assign new_n4801 = ~new_n4774 & ~new_n4800;
  assign new_n4802 = ~new_n4614 & new_n4801;
  assign new_n4803 = new_n4614 & ~new_n4801;
  assign new_n4804 = ~new_n4802 & ~new_n4803;
  assign new_n4805_1 = n8336 & n10439;
  assign new_n4806 = ~new_n4633 & ~new_n4644;
  assign new_n4807 = ~new_n4634_1 & ~new_n4806;
  assign new_n4808 = ~new_n4805_1 & new_n4807;
  assign new_n4809 = n8595 & n10928;
  assign new_n4810 = new_n4636 & ~new_n4639;
  assign new_n4811 = ~new_n4640 & ~new_n4810;
  assign new_n4812 = new_n4809 & ~new_n4811;
  assign new_n4813 = ~new_n4809 & new_n4811;
  assign new_n4814 = ~new_n4812 & ~new_n4813;
  assign new_n4815 = n2226 & n3602;
  assign new_n4816 = n6126 & n6986;
  assign new_n4817_1 = n1094 & n3719;
  assign new_n4818 = ~new_n4816 & ~new_n4817_1;
  assign new_n4819 = new_n4816 & new_n4817_1;
  assign new_n4820 = ~new_n4818 & ~new_n4819;
  assign new_n4821 = new_n4815 & ~new_n4820;
  assign new_n4822 = ~new_n4815 & new_n4820;
  assign new_n4823 = ~new_n4821 & ~new_n4822;
  assign new_n4824 = ~new_n4814 & ~new_n4823;
  assign new_n4825 = new_n4814 & new_n4823;
  assign new_n4826_1 = ~new_n4824 & ~new_n4825;
  assign new_n4827 = new_n4808 & new_n4826_1;
  assign new_n4828_1 = new_n4805_1 & ~new_n4807;
  assign new_n4829 = new_n4826_1 & ~new_n4828_1;
  assign new_n4830 = ~new_n4808 & ~new_n4829;
  assign new_n4831 = ~new_n4827 & ~new_n4830;
  assign new_n4832 = ~new_n4826_1 & new_n4828_1;
  assign new_n4833 = ~new_n4831 & ~new_n4832;
  assign new_n4834 = new_n4649 & ~new_n4833;
  assign new_n4835 = ~new_n4649 & new_n4833;
  assign new_n4836 = ~new_n4834 & ~new_n4835;
  assign new_n4837 = n6611 & n11222;
  assign new_n4838 = n217 & n11153;
  assign new_n4839 = n5767 & n8433;
  assign new_n4840 = n405 & n996;
  assign new_n4841 = ~new_n4689_1 & ~new_n4840;
  assign new_n4842 = new_n4689_1 & new_n4840;
  assign new_n4843 = ~new_n4841 & ~new_n4842;
  assign new_n4844 = new_n4839 & ~new_n4843;
  assign new_n4845 = ~new_n4839 & new_n4843;
  assign new_n4846 = ~new_n4844 & ~new_n4845;
  assign new_n4847 = new_n4838 & ~new_n4846;
  assign new_n4848 = ~new_n4838 & new_n4846;
  assign new_n4849 = ~new_n4847 & ~new_n4848;
  assign new_n4850 = new_n4703 & ~new_n4706;
  assign new_n4851 = ~new_n4707 & ~new_n4850;
  assign new_n4852 = ~new_n4849 & ~new_n4851;
  assign new_n4853 = new_n4849 & new_n4851;
  assign new_n4854 = ~new_n4852 & ~new_n4853;
  assign new_n4855 = new_n4837 & ~new_n4854;
  assign new_n4856 = ~new_n4837 & new_n4854;
  assign new_n4857 = ~new_n4855 & ~new_n4856;
  assign new_n4858 = ~new_n4701 & ~new_n4711;
  assign new_n4859 = ~new_n4700 & ~new_n4858;
  assign new_n4860 = ~new_n4857 & ~new_n4859;
  assign new_n4861 = new_n4857 & new_n4859;
  assign new_n4862 = ~new_n4860 & ~new_n4861;
  assign new_n4863 = ~new_n4715 & new_n4862;
  assign new_n4864 = new_n4715 & ~new_n4862;
  assign new_n4865 = ~new_n4863 & ~new_n4864;
  assign new_n4866 = n4970 & n12069;
  assign new_n4867 = n7610 & n12391;
  assign new_n4868 = new_n4670 & ~new_n4673;
  assign new_n4869 = ~new_n4674 & ~new_n4868;
  assign new_n4870 = new_n4867 & ~new_n4869;
  assign new_n4871 = ~new_n4867 & new_n4869;
  assign new_n4872 = ~new_n4870 & ~new_n4871;
  assign new_n4873 = n7160 & n7733;
  assign new_n4874 = n4826 & n7891;
  assign new_n4875 = n4828 & n12925;
  assign new_n4876 = ~new_n4874 & ~new_n4875;
  assign new_n4877 = new_n4874 & new_n4875;
  assign new_n4878 = ~new_n4876 & ~new_n4877;
  assign new_n4879 = new_n4873 & ~new_n4878;
  assign new_n4880 = ~new_n4873 & new_n4878;
  assign new_n4881 = ~new_n4879 & ~new_n4880;
  assign new_n4882 = ~new_n4872 & ~new_n4881;
  assign new_n4883 = new_n4872 & new_n4881;
  assign new_n4884 = ~new_n4882 & ~new_n4883;
  assign new_n4885 = new_n4866 & ~new_n4884;
  assign new_n4886 = ~new_n4866 & new_n4884;
  assign new_n4887 = ~new_n4885 & ~new_n4886;
  assign new_n4888 = ~new_n4667 & ~new_n4678;
  assign new_n4889 = ~new_n4668 & ~new_n4888;
  assign new_n4890 = ~new_n4887 & ~new_n4889;
  assign new_n4891 = new_n4887 & new_n4889;
  assign new_n4892 = ~new_n4890 & ~new_n4891;
  assign new_n4893 = new_n4683 & ~new_n4892;
  assign new_n4894 = ~new_n4683 & new_n4892;
  assign new_n4895 = ~new_n4893 & ~new_n4894;
  assign new_n4896 = ~new_n4719 & ~new_n4740;
  assign new_n4897 = ~new_n4718 & ~new_n4896;
  assign new_n4898 = new_n4895 & ~new_n4897;
  assign new_n4899 = ~new_n4895 & new_n4897;
  assign new_n4900 = ~new_n4898 & ~new_n4899;
  assign new_n4901 = new_n4865 & new_n4900;
  assign new_n4902 = ~new_n4865 & ~new_n4900;
  assign new_n4903_1 = ~new_n4901 & ~new_n4902;
  assign new_n4904 = new_n4836 & new_n4903_1;
  assign new_n4905 = ~new_n4836 & ~new_n4903_1;
  assign new_n4906 = ~new_n4904 & ~new_n4905;
  assign new_n4907 = ~new_n4744 & ~new_n4770;
  assign new_n4908 = ~new_n4745 & ~new_n4907;
  assign new_n4909 = new_n4906 & ~new_n4908;
  assign new_n4910 = ~new_n4906 & new_n4908;
  assign new_n4911 = ~new_n4909 & ~new_n4910;
  assign new_n4912 = new_n4804 & ~new_n4911;
  assign new_n4913 = ~new_n4804 & new_n4911;
  assign n992 = ~new_n4912 & ~new_n4913;
  assign new_n4915 = n6687 & n7265;
  assign new_n4916 = n7946 & n8336;
  assign new_n4917 = n9763 & n11222;
  assign new_n4918 = n2558 & n12069;
  assign new_n4919 = new_n4917 & new_n4918;
  assign new_n4920 = ~new_n4917 & ~new_n4918;
  assign new_n4921_1 = ~new_n4919 & ~new_n4920;
  assign new_n4922 = new_n4916 & new_n4921_1;
  assign new_n4923 = ~new_n4916 & ~new_n4921_1;
  assign new_n4924 = ~new_n4922 & ~new_n4923;
  assign new_n4925 = new_n4915 & new_n4924;
  assign new_n4926 = ~new_n4915 & ~new_n4924;
  assign n1020 = ~new_n4925 & ~new_n4926;
  assign new_n4928_1 = ~new_n2288 & ~new_n2289;
  assign new_n4929 = new_n2331 & ~new_n4928_1;
  assign new_n4930 = ~new_n2331 & new_n4928_1;
  assign n1136 = ~new_n4929 & ~new_n4930;
  assign new_n4932 = ~new_n4774 & ~new_n4775;
  assign new_n4933 = new_n4799 & ~new_n4932;
  assign new_n4934 = ~new_n4799 & new_n4932;
  assign n1138 = ~new_n4933 & ~new_n4934;
  assign new_n4936 = n159 & n7236;
  assign new_n4937 = n2749 & n7236;
  assign new_n4938_1 = n3754 & n7236;
  assign new_n4939 = n3992 & n10898;
  assign new_n4940 = new_n4938_1 & new_n4939;
  assign new_n4941 = ~new_n4938_1 & ~new_n4939;
  assign new_n4942 = n8384 & n11876;
  assign new_n4943 = ~new_n4941 & new_n4942;
  assign new_n4944 = ~new_n4940 & ~new_n4943;
  assign new_n4945 = ~new_n4937 & new_n4944;
  assign new_n4946 = new_n4937 & ~new_n4944;
  assign new_n4947 = n8384 & n10898;
  assign new_n4948 = n3754 & n6358;
  assign new_n4949 = n3992 & n11876;
  assign new_n4950 = new_n4948 & new_n4949;
  assign new_n4951 = n6358 & n11876;
  assign new_n4952 = n3754 & n3992;
  assign new_n4953 = ~new_n4951 & ~new_n4952;
  assign new_n4954 = ~new_n4950 & ~new_n4953;
  assign new_n4955 = ~new_n4947 & ~new_n4954;
  assign new_n4956 = new_n4947 & new_n4954;
  assign new_n4957 = ~new_n4955 & ~new_n4956;
  assign new_n4958 = ~new_n4946 & ~new_n4957;
  assign new_n4959 = ~new_n4945 & ~new_n4958;
  assign new_n4960 = ~new_n4936 & ~new_n4959;
  assign new_n4961 = new_n4936 & new_n4959;
  assign new_n4962 = n6358 & n10898;
  assign new_n4963 = n5198 & n11876;
  assign new_n4964 = n3754 & n8384;
  assign new_n4965 = ~new_n4963 & ~new_n4964;
  assign new_n4966 = n3754 & n5198;
  assign new_n4967 = new_n4942 & new_n4966;
  assign new_n4968 = ~new_n4965 & ~new_n4967;
  assign new_n4969 = ~new_n4962 & ~new_n4968;
  assign new_n4970_1 = new_n4962 & new_n4968;
  assign new_n4971_1 = ~new_n4969 & ~new_n4970_1;
  assign new_n4972 = n2749 & n3992;
  assign new_n4973 = new_n4947 & ~new_n4953;
  assign new_n4974 = ~new_n4950 & ~new_n4973;
  assign new_n4975 = ~new_n4972 & new_n4974;
  assign new_n4976 = new_n4972 & ~new_n4974;
  assign new_n4977 = ~new_n4975 & ~new_n4976;
  assign new_n4978 = new_n4971_1 & ~new_n4977;
  assign new_n4979 = ~new_n4971_1 & new_n4977;
  assign new_n4980 = ~new_n4978 & ~new_n4979;
  assign new_n4981 = ~new_n4961 & new_n4980;
  assign new_n4982 = ~new_n4960 & ~new_n4981;
  assign new_n4983 = n2749 & n8384;
  assign new_n4984 = n159 & n3992;
  assign new_n4985 = ~new_n4983 & ~new_n4984;
  assign new_n4986 = new_n4983 & new_n4984;
  assign new_n4987 = ~new_n4985 & ~new_n4986;
  assign new_n4988 = ~new_n4971_1 & ~new_n4976;
  assign new_n4989 = ~new_n4975 & ~new_n4988;
  assign new_n4990 = new_n4987 & new_n4989;
  assign new_n4991 = ~new_n4987 & ~new_n4989;
  assign new_n4992 = ~new_n4990 & ~new_n4991;
  assign new_n4993 = n5198 & n10898;
  assign new_n4994 = n1471 & n11876;
  assign new_n4995 = ~new_n4993 & ~new_n4994;
  assign new_n4996 = new_n4993 & new_n4994;
  assign new_n4997 = ~new_n4995 & ~new_n4996;
  assign new_n4998 = ~new_n4948 & ~new_n4997;
  assign new_n4999 = new_n4948 & new_n4997;
  assign new_n5000 = ~new_n4998 & ~new_n4999;
  assign new_n5001 = new_n4962 & ~new_n4965;
  assign new_n5002 = ~new_n4967 & ~new_n5001;
  assign new_n5003 = ~new_n5000 & new_n5002;
  assign new_n5004 = new_n5000 & ~new_n5002;
  assign new_n5005 = ~new_n5003 & ~new_n5004;
  assign new_n5006 = ~new_n4992 & new_n5005;
  assign new_n5007 = new_n4992 & ~new_n5005;
  assign new_n5008 = ~new_n5006 & ~new_n5007;
  assign new_n5009 = new_n4982 & ~new_n5008;
  assign new_n5010 = ~new_n4991 & new_n5005;
  assign new_n5011 = ~new_n4986 & ~new_n5010;
  assign new_n5012 = ~new_n4990 & new_n5011;
  assign new_n5013 = new_n4986 & new_n5010;
  assign new_n5014 = ~new_n5012 & ~new_n5013;
  assign new_n5015 = n1510 & n3992;
  assign new_n5016 = n159 & n8384;
  assign new_n5017 = n7236 & n12247;
  assign new_n5018 = ~new_n5016 & ~new_n5017;
  assign new_n5019 = new_n5016 & new_n5017;
  assign new_n5020 = ~new_n5018 & ~new_n5019;
  assign new_n5021 = ~new_n5015 & ~new_n5020;
  assign new_n5022 = new_n5015 & new_n5020;
  assign new_n5023 = ~new_n5021 & ~new_n5022;
  assign new_n5024 = ~new_n4999 & new_n5002;
  assign new_n5025 = ~new_n4998 & ~new_n5024;
  assign new_n5026 = ~new_n5023 & ~new_n5025;
  assign new_n5027 = new_n5023 & new_n5025;
  assign new_n5028 = ~new_n5026 & ~new_n5027;
  assign new_n5029 = n2749 & n6358;
  assign new_n5030_1 = ~new_n4996 & ~new_n5029;
  assign new_n5031 = new_n4996 & new_n5029;
  assign new_n5032 = ~new_n5030_1 & ~new_n5031;
  assign new_n5033 = n1471 & n10898;
  assign new_n5034_1 = n7646 & n11876;
  assign new_n5035 = ~new_n4966 & ~new_n5034_1;
  assign new_n5036 = new_n4966 & new_n5034_1;
  assign new_n5037 = ~new_n5035 & ~new_n5036;
  assign new_n5038 = ~new_n5033 & ~new_n5037;
  assign new_n5039 = new_n5033 & new_n5037;
  assign new_n5040 = ~new_n5038 & ~new_n5039;
  assign new_n5041 = new_n5032 & ~new_n5040;
  assign new_n5042 = ~new_n5032 & new_n5040;
  assign new_n5043 = ~new_n5041 & ~new_n5042;
  assign new_n5044 = new_n5028 & ~new_n5043;
  assign new_n5045 = ~new_n5028 & new_n5043;
  assign new_n5046 = ~new_n5044 & ~new_n5045;
  assign new_n5047 = new_n5014 & ~new_n5046;
  assign new_n5048 = ~new_n5014 & new_n5046;
  assign new_n5049 = ~new_n5047 & ~new_n5048;
  assign new_n5050 = new_n5009 & ~new_n5049;
  assign new_n5051 = ~new_n5009 & new_n5049;
  assign new_n5052 = ~new_n5050 & ~new_n5051;
  assign new_n5053 = n1510 & n7236;
  assign new_n5054 = ~new_n4982 & new_n5008;
  assign new_n5055 = ~new_n5009 & ~new_n5054;
  assign new_n5056 = new_n5053 & new_n5055;
  assign new_n5057 = n7236 & n10898;
  assign new_n5058 = new_n4949 & new_n5057;
  assign new_n5059 = ~new_n4940 & ~new_n4941;
  assign new_n5060 = ~new_n4942 & ~new_n5059;
  assign new_n5061 = new_n4942 & new_n5059;
  assign new_n5062 = ~new_n5060 & ~new_n5061;
  assign new_n5063 = new_n5058 & new_n5062;
  assign new_n5064 = ~new_n4945 & ~new_n4946;
  assign new_n5065 = new_n4957 & ~new_n5064;
  assign new_n5066 = ~new_n4957 & new_n5064;
  assign new_n5067 = ~new_n5065 & ~new_n5066;
  assign new_n5068 = new_n5063 & ~new_n5067;
  assign new_n5069_1 = ~new_n4960 & ~new_n4961;
  assign new_n5070 = ~new_n4980 & ~new_n5069_1;
  assign new_n5071 = new_n4980 & new_n5069_1;
  assign new_n5072 = ~new_n5070 & ~new_n5071;
  assign new_n5073 = new_n5068 & ~new_n5072;
  assign new_n5074 = ~new_n5053 & ~new_n5055;
  assign new_n5075 = ~new_n5056 & ~new_n5074;
  assign new_n5076 = new_n5073 & new_n5075;
  assign new_n5077 = ~new_n5056 & ~new_n5076;
  assign new_n5078 = new_n5052 & ~new_n5077;
  assign new_n5079 = ~new_n5050 & ~new_n5078;
  assign new_n5080 = n7862 & n11662;
  assign new_n5081 = n1333 & n7456;
  assign new_n5082 = n1333 & n12591;
  assign new_n5083 = n3172 & n3932;
  assign new_n5084 = new_n5082 & new_n5083;
  assign new_n5085 = ~new_n5082 & ~new_n5083;
  assign new_n5086 = n1798 & n11757;
  assign new_n5087 = ~new_n5085 & new_n5086;
  assign new_n5088 = ~new_n5084 & ~new_n5087;
  assign new_n5089 = ~new_n5081 & new_n5088;
  assign new_n5090 = new_n5081 & ~new_n5088;
  assign new_n5091 = ~new_n5089 & ~new_n5090;
  assign new_n5092 = n1798 & n5240;
  assign new_n5093 = n3172 & n12591;
  assign new_n5094_1 = n3932 & n11757;
  assign new_n5095 = ~new_n5093 & ~new_n5094_1;
  assign new_n5096 = new_n5093 & new_n5094_1;
  assign new_n5097 = ~new_n5095 & ~new_n5096;
  assign new_n5098 = new_n5092 & ~new_n5097;
  assign new_n5099 = ~new_n5092 & new_n5097;
  assign new_n5100 = ~new_n5098 & ~new_n5099;
  assign new_n5101 = ~new_n5091 & new_n5100;
  assign new_n5102 = new_n5091 & ~new_n5100;
  assign new_n5103 = ~new_n5101 & ~new_n5102;
  assign new_n5104 = new_n5080 & new_n5103;
  assign new_n5105_1 = ~new_n5080 & ~new_n5103;
  assign new_n5106 = n7456 & n7862;
  assign new_n5107 = n1333 & n3932;
  assign new_n5108 = n7862 & n12591;
  assign new_n5109 = new_n5107 & new_n5108;
  assign new_n5110 = ~new_n5107 & ~new_n5108;
  assign new_n5111 = n1798 & n3172;
  assign new_n5112 = ~new_n5110 & new_n5111;
  assign new_n5113 = ~new_n5109 & ~new_n5112;
  assign new_n5114 = ~new_n5106 & new_n5113;
  assign new_n5115 = new_n5106 & ~new_n5113;
  assign new_n5116 = ~new_n5084 & ~new_n5085;
  assign new_n5117 = ~new_n5086 & ~new_n5116;
  assign new_n5118 = new_n5086 & new_n5116;
  assign new_n5119 = ~new_n5117 & ~new_n5118;
  assign new_n5120 = ~new_n5115 & ~new_n5119;
  assign new_n5121 = ~new_n5114 & ~new_n5120;
  assign new_n5122 = ~new_n5105_1 & new_n5121;
  assign new_n5123 = ~new_n5104 & ~new_n5122;
  assign new_n5124 = n1333 & n11662;
  assign new_n5125 = n3172 & n7456;
  assign new_n5126 = ~new_n5124 & ~new_n5125;
  assign new_n5127 = new_n5124 & new_n5125;
  assign new_n5128 = ~new_n5126 & ~new_n5127;
  assign new_n5129 = ~new_n5089 & ~new_n5100;
  assign new_n5130 = ~new_n5090 & ~new_n5129;
  assign new_n5131 = ~new_n5128 & new_n5130;
  assign new_n5132_1 = new_n5128 & ~new_n5130;
  assign new_n5133 = ~new_n5131 & ~new_n5132_1;
  assign new_n5134 = ~new_n5092 & ~new_n5096;
  assign new_n5135 = ~new_n5095 & ~new_n5134;
  assign new_n5136 = n11757 & n12591;
  assign new_n5137 = n3932 & n5240;
  assign new_n5138 = n1798 & n11821;
  assign new_n5139 = ~new_n5137 & ~new_n5138;
  assign new_n5140 = new_n5137 & new_n5138;
  assign new_n5141 = ~new_n5139 & ~new_n5140;
  assign new_n5142 = ~new_n5136 & ~new_n5141;
  assign new_n5143 = new_n5136 & new_n5141;
  assign new_n5144 = ~new_n5142 & ~new_n5143;
  assign new_n5145 = ~new_n5135 & ~new_n5144;
  assign new_n5146 = new_n5135 & new_n5144;
  assign new_n5147 = ~new_n5145 & ~new_n5146;
  assign new_n5148 = ~new_n5133 & ~new_n5147;
  assign new_n5149 = new_n5133 & new_n5147;
  assign new_n5150 = ~new_n5148 & ~new_n5149;
  assign new_n5151 = ~new_n5123 & new_n5150;
  assign new_n5152 = n7456 & n11757;
  assign new_n5153_1 = new_n5140 & new_n5152;
  assign new_n5154 = ~new_n5140 & ~new_n5152;
  assign new_n5155 = ~new_n5153_1 & ~new_n5154;
  assign new_n5156 = n1798 & n9080;
  assign new_n5157 = n3932 & n11821;
  assign new_n5158 = n5240 & n12591;
  assign new_n5159 = ~new_n5157 & ~new_n5158;
  assign new_n5160 = new_n5157 & new_n5158;
  assign new_n5161 = ~new_n5159 & ~new_n5160;
  assign new_n5162 = new_n5156 & ~new_n5161;
  assign new_n5163 = ~new_n5156 & new_n5161;
  assign new_n5164 = ~new_n5162 & ~new_n5163;
  assign new_n5165 = new_n5155 & new_n5164;
  assign new_n5166 = ~new_n5155 & ~new_n5164;
  assign new_n5167 = ~new_n5165 & ~new_n5166;
  assign new_n5168 = n1333 & n10327;
  assign new_n5169 = n3172 & n11662;
  assign new_n5170 = n7862 & n9583;
  assign new_n5171 = ~new_n5169 & ~new_n5170;
  assign new_n5172 = new_n5169 & new_n5170;
  assign new_n5173 = ~new_n5171 & ~new_n5172;
  assign new_n5174 = ~new_n5168 & ~new_n5173;
  assign new_n5175 = new_n5168 & new_n5173;
  assign new_n5176 = ~new_n5174 & ~new_n5175;
  assign new_n5177 = new_n5135 & ~new_n5142;
  assign new_n5178 = ~new_n5143 & ~new_n5177;
  assign new_n5179 = ~new_n5176 & new_n5178;
  assign new_n5180 = new_n5176 & ~new_n5178;
  assign new_n5181 = ~new_n5179 & ~new_n5180;
  assign new_n5182 = ~new_n5167 & new_n5181;
  assign new_n5183 = new_n5167 & ~new_n5181;
  assign new_n5184 = ~new_n5182 & ~new_n5183;
  assign new_n5185 = ~new_n5131 & new_n5147;
  assign new_n5186 = new_n5127 & new_n5185;
  assign new_n5187 = ~new_n5127 & ~new_n5185;
  assign new_n5188 = ~new_n5132_1 & new_n5187;
  assign new_n5189 = ~new_n5186 & ~new_n5188;
  assign new_n5190 = new_n5184 & new_n5189;
  assign new_n5191_1 = ~new_n5184 & ~new_n5189;
  assign new_n5192 = ~new_n5190 & ~new_n5191_1;
  assign new_n5193 = new_n5151 & new_n5192;
  assign new_n5194 = ~new_n5151 & ~new_n5192;
  assign new_n5195 = ~new_n5193 & ~new_n5194;
  assign new_n5196 = n7862 & n10327;
  assign new_n5197 = new_n5123 & ~new_n5150;
  assign new_n5198_1 = ~new_n5151 & ~new_n5197;
  assign new_n5199 = new_n5196 & new_n5198_1;
  assign new_n5200 = n3932 & n7862;
  assign new_n5201 = n1333 & n1798;
  assign new_n5202 = new_n5200 & new_n5201;
  assign new_n5203 = ~new_n5109 & ~new_n5110;
  assign new_n5204 = ~new_n5111 & ~new_n5203;
  assign new_n5205 = new_n5111 & new_n5203;
  assign new_n5206 = ~new_n5204 & ~new_n5205;
  assign new_n5207 = new_n5202 & new_n5206;
  assign new_n5208 = ~new_n5114 & ~new_n5115;
  assign new_n5209 = new_n5119 & ~new_n5208;
  assign new_n5210 = ~new_n5119 & new_n5208;
  assign new_n5211 = ~new_n5209 & ~new_n5210;
  assign new_n5212_1 = new_n5207 & ~new_n5211;
  assign new_n5213 = ~new_n5104 & ~new_n5105_1;
  assign new_n5214 = new_n5121 & new_n5213;
  assign new_n5215 = ~new_n5121 & ~new_n5213;
  assign new_n5216 = ~new_n5214 & ~new_n5215;
  assign new_n5217 = new_n5212_1 & new_n5216;
  assign new_n5218 = ~new_n5196 & ~new_n5198_1;
  assign new_n5219 = ~new_n5199 & ~new_n5218;
  assign new_n5220 = new_n5217 & new_n5219;
  assign new_n5221 = ~new_n5199 & ~new_n5220;
  assign new_n5222 = new_n5195 & ~new_n5221;
  assign new_n5223 = ~new_n5195 & new_n5221;
  assign new_n5224 = ~new_n5222 & ~new_n5223;
  assign new_n5225 = n6877 & n10451;
  assign new_n5226 = n9400 & n11023;
  assign new_n5227 = n2464 & n9640;
  assign new_n5228 = n3022 & n9400;
  assign new_n5229 = new_n5227 & new_n5228;
  assign new_n5230 = ~new_n5227 & ~new_n5228;
  assign new_n5231 = n6703 & n11311;
  assign new_n5232 = ~new_n5230 & new_n5231;
  assign new_n5233 = ~new_n5229 & ~new_n5232;
  assign new_n5234 = ~new_n5226 & new_n5233;
  assign new_n5235 = new_n5226 & ~new_n5233;
  assign new_n5236 = ~new_n5234 & ~new_n5235;
  assign new_n5237 = n4187 & n6703;
  assign new_n5238 = n2464 & n3022;
  assign new_n5239 = n9640 & n11311;
  assign new_n5240_1 = ~new_n5238 & ~new_n5239;
  assign new_n5241 = new_n5238 & new_n5239;
  assign new_n5242 = ~new_n5240_1 & ~new_n5241;
  assign new_n5243 = new_n5237 & ~new_n5242;
  assign new_n5244 = ~new_n5237 & new_n5242;
  assign new_n5245 = ~new_n5243 & ~new_n5244;
  assign new_n5246 = ~new_n5236 & new_n5245;
  assign new_n5247 = new_n5236 & ~new_n5245;
  assign new_n5248 = ~new_n5246 & ~new_n5247;
  assign new_n5249 = new_n5225 & new_n5248;
  assign new_n5250 = ~new_n5225 & ~new_n5248;
  assign new_n5251 = n6877 & n11023;
  assign new_n5252 = n9400 & n9640;
  assign new_n5253 = n3022 & n6877;
  assign new_n5254 = new_n5252 & new_n5253;
  assign new_n5255 = ~new_n5252 & ~new_n5253;
  assign new_n5256 = n2464 & n6703;
  assign new_n5257_1 = ~new_n5255 & new_n5256;
  assign new_n5258 = ~new_n5254 & ~new_n5257_1;
  assign new_n5259 = ~new_n5251 & new_n5258;
  assign new_n5260 = new_n5251 & ~new_n5258;
  assign new_n5261 = ~new_n5229 & ~new_n5230;
  assign new_n5262 = ~new_n5231 & ~new_n5261;
  assign new_n5263 = new_n5231 & new_n5261;
  assign new_n5264 = ~new_n5262 & ~new_n5263;
  assign new_n5265 = ~new_n5260 & ~new_n5264;
  assign new_n5266 = ~new_n5259 & ~new_n5265;
  assign new_n5267 = ~new_n5250 & new_n5266;
  assign new_n5268 = ~new_n5249 & ~new_n5267;
  assign new_n5269 = n9400 & n10451;
  assign new_n5270 = n2464 & n11023;
  assign new_n5271 = ~new_n5269 & ~new_n5270;
  assign new_n5272 = new_n5269 & new_n5270;
  assign new_n5273 = ~new_n5271 & ~new_n5272;
  assign new_n5274 = n3022 & n11311;
  assign new_n5275 = n4187 & n9640;
  assign new_n5276 = n4203 & n6703;
  assign new_n5277 = ~new_n5275 & ~new_n5276;
  assign new_n5278 = new_n5275 & new_n5276;
  assign new_n5279 = ~new_n5277 & ~new_n5278;
  assign new_n5280 = new_n5274 & new_n5279;
  assign new_n5281 = ~new_n5274 & ~new_n5279;
  assign new_n5282 = ~new_n5280 & ~new_n5281;
  assign new_n5283_1 = ~new_n5237 & ~new_n5241;
  assign new_n5284 = ~new_n5240_1 & ~new_n5283_1;
  assign new_n5285 = ~new_n5282 & new_n5284;
  assign new_n5286 = new_n5282 & ~new_n5284;
  assign new_n5287 = ~new_n5285 & ~new_n5286;
  assign new_n5288 = new_n5273 & ~new_n5287;
  assign new_n5289 = ~new_n5273 & new_n5287;
  assign new_n5290 = ~new_n5288 & ~new_n5289;
  assign new_n5291 = ~new_n5234 & ~new_n5245;
  assign new_n5292 = ~new_n5235 & ~new_n5291;
  assign new_n5293 = new_n5290 & new_n5292;
  assign new_n5294 = ~new_n5290 & ~new_n5292;
  assign new_n5295 = ~new_n5293 & ~new_n5294;
  assign new_n5296 = ~new_n5268 & ~new_n5295;
  assign new_n5297 = ~new_n5289 & ~new_n5292;
  assign new_n5298 = ~new_n5272 & ~new_n5297;
  assign new_n5299 = ~new_n5288 & new_n5298;
  assign new_n5300 = new_n5272 & new_n5297;
  assign new_n5301 = ~new_n5299 & ~new_n5300;
  assign new_n5302 = n2464 & n10451;
  assign new_n5303 = n6877 & n11423;
  assign new_n5304 = n9400 & n10278;
  assign new_n5305_1 = ~new_n5303 & ~new_n5304;
  assign new_n5306 = new_n5303 & new_n5304;
  assign new_n5307 = ~new_n5305_1 & ~new_n5306;
  assign new_n5308 = new_n5302 & ~new_n5307;
  assign new_n5309 = ~new_n5302 & new_n5307;
  assign new_n5310 = ~new_n5308 & ~new_n5309;
  assign new_n5311 = ~new_n5280 & ~new_n5284;
  assign new_n5312 = ~new_n5281 & ~new_n5311;
  assign new_n5313 = new_n5310 & ~new_n5312;
  assign new_n5314_1 = n11023 & n11311;
  assign new_n5315 = new_n5278 & new_n5314_1;
  assign new_n5316 = ~new_n5278 & ~new_n5314_1;
  assign new_n5317 = ~new_n5315 & ~new_n5316;
  assign new_n5318 = n6703 & n12753;
  assign new_n5319_1 = n4203 & n9640;
  assign new_n5320_1 = n3022 & n4187;
  assign new_n5321 = ~new_n5319_1 & ~new_n5320_1;
  assign new_n5322 = new_n5319_1 & new_n5320_1;
  assign new_n5323 = ~new_n5321 & ~new_n5322;
  assign new_n5324 = new_n5318 & ~new_n5323;
  assign new_n5325 = ~new_n5318 & new_n5323;
  assign new_n5326 = ~new_n5324 & ~new_n5325;
  assign new_n5327 = new_n5317 & new_n5326;
  assign new_n5328 = ~new_n5317 & ~new_n5326;
  assign new_n5329 = ~new_n5327 & ~new_n5328;
  assign new_n5330 = new_n5313 & new_n5329;
  assign new_n5331_1 = ~new_n5310 & new_n5312;
  assign new_n5332 = ~new_n5329 & new_n5331_1;
  assign new_n5333 = ~new_n5313 & ~new_n5329;
  assign new_n5334 = ~new_n5331_1 & ~new_n5333;
  assign new_n5335 = ~new_n5332 & ~new_n5334;
  assign new_n5336 = ~new_n5330 & ~new_n5335;
  assign new_n5337 = new_n5301 & ~new_n5336;
  assign new_n5338 = ~new_n5301 & new_n5336;
  assign new_n5339 = ~new_n5337 & ~new_n5338;
  assign new_n5340 = ~new_n5296 & new_n5339;
  assign new_n5341 = new_n5296 & ~new_n5339;
  assign new_n5342 = ~new_n5340 & ~new_n5341;
  assign new_n5343 = n6877 & n10278;
  assign new_n5344 = new_n5268 & new_n5295;
  assign new_n5345 = ~new_n5296 & ~new_n5344;
  assign new_n5346 = new_n5343 & new_n5345;
  assign new_n5347 = n6877 & n9640;
  assign new_n5348 = n6703 & n9400;
  assign new_n5349 = new_n5347 & new_n5348;
  assign new_n5350 = ~new_n5254 & ~new_n5255;
  assign new_n5351 = ~new_n5256 & ~new_n5350;
  assign new_n5352 = new_n5256 & new_n5350;
  assign new_n5353 = ~new_n5351 & ~new_n5352;
  assign new_n5354 = new_n5349 & new_n5353;
  assign new_n5355 = ~new_n5259 & ~new_n5260;
  assign new_n5356 = ~new_n5264 & ~new_n5355;
  assign new_n5357 = new_n5264 & new_n5355;
  assign new_n5358 = ~new_n5356 & ~new_n5357;
  assign new_n5359 = new_n5354 & new_n5358;
  assign new_n5360 = ~new_n5249 & ~new_n5250;
  assign new_n5361 = ~new_n5266 & ~new_n5360;
  assign new_n5362 = new_n5266 & new_n5360;
  assign new_n5363 = ~new_n5361 & ~new_n5362;
  assign new_n5364 = new_n5359 & new_n5363;
  assign new_n5365 = ~new_n5343 & ~new_n5345;
  assign new_n5366 = ~new_n5346 & ~new_n5365;
  assign new_n5367 = new_n5364 & new_n5366;
  assign new_n5368 = ~new_n5346 & ~new_n5367;
  assign new_n5369 = ~new_n5342 & new_n5368;
  assign new_n5370 = new_n5342 & ~new_n5368;
  assign new_n5371 = ~new_n5369 & ~new_n5370;
  assign new_n5372 = n4805 & n12826;
  assign new_n5373 = n2551 & n11478;
  assign new_n5374 = n5283 & n11922;
  assign new_n5375 = ~new_n5373 & ~new_n5374;
  assign new_n5376 = new_n5373 & new_n5374;
  assign new_n5377 = ~new_n5375 & ~new_n5376;
  assign new_n5378 = n11478 & n11922;
  assign new_n5379 = n8665 & n11478;
  assign new_n5380 = n1067 & n5283;
  assign new_n5381 = ~new_n5379 & ~new_n5380;
  assign new_n5382 = n137 & n5645;
  assign new_n5383 = new_n5379 & new_n5380;
  assign new_n5384 = ~new_n5382 & ~new_n5383;
  assign new_n5385 = ~new_n5381 & ~new_n5384;
  assign new_n5386 = new_n5378 & new_n5385;
  assign new_n5387 = ~new_n5378 & ~new_n5385;
  assign new_n5388 = n137 & n1067;
  assign new_n5389 = n5283 & n8665;
  assign new_n5390 = n5645 & n6294;
  assign new_n5391 = ~new_n5389 & ~new_n5390;
  assign new_n5392 = new_n5389 & new_n5390;
  assign new_n5393 = ~new_n5391 & ~new_n5392;
  assign new_n5394 = new_n5388 & ~new_n5393;
  assign new_n5395 = ~new_n5388 & new_n5393;
  assign new_n5396 = ~new_n5394 & ~new_n5395;
  assign new_n5397 = ~new_n5387 & ~new_n5396;
  assign new_n5398 = ~new_n5386 & ~new_n5397;
  assign new_n5399 = ~new_n5377 & new_n5398;
  assign new_n5400 = new_n5377 & ~new_n5398;
  assign new_n5401 = ~new_n5399 & ~new_n5400;
  assign new_n5402 = n137 & n8665;
  assign new_n5403 = n1067 & n6294;
  assign new_n5404 = n5645 & n6797;
  assign new_n5405 = ~new_n5403 & ~new_n5404;
  assign new_n5406 = new_n5403 & new_n5404;
  assign new_n5407 = ~new_n5405 & ~new_n5406;
  assign new_n5408 = new_n5402 & new_n5407;
  assign new_n5409 = ~new_n5402 & ~new_n5407;
  assign new_n5410 = ~new_n5408 & ~new_n5409;
  assign new_n5411_1 = new_n5388 & ~new_n5391;
  assign new_n5412 = ~new_n5392 & ~new_n5411_1;
  assign new_n5413 = ~new_n5410 & ~new_n5412;
  assign new_n5414 = new_n5410 & new_n5412;
  assign new_n5415 = ~new_n5413 & ~new_n5414;
  assign new_n5416 = ~new_n5401 & ~new_n5415;
  assign new_n5417 = new_n5401 & new_n5415;
  assign new_n5418 = ~new_n5416 & ~new_n5417;
  assign new_n5419 = n2551 & n4805;
  assign new_n5420 = n4805 & n11922;
  assign new_n5421 = n4805 & n5645;
  assign new_n5422 = new_n5389 & new_n5421;
  assign new_n5423 = n1067 & n11478;
  assign new_n5424 = n5283 & n5645;
  assign new_n5425 = n4805 & n8665;
  assign new_n5426 = ~new_n5424 & ~new_n5425;
  assign new_n5427 = new_n5423 & ~new_n5426;
  assign new_n5428 = ~new_n5422 & ~new_n5427;
  assign new_n5429 = new_n5420 & ~new_n5428;
  assign new_n5430 = ~new_n5420 & new_n5428;
  assign new_n5431 = ~new_n5381 & ~new_n5383;
  assign new_n5432 = new_n5382 & ~new_n5431;
  assign new_n5433 = ~new_n5382 & new_n5431;
  assign new_n5434 = ~new_n5432 & ~new_n5433;
  assign new_n5435_1 = ~new_n5430 & ~new_n5434;
  assign new_n5436 = ~new_n5429 & ~new_n5435_1;
  assign new_n5437 = new_n5419 & ~new_n5436;
  assign new_n5438 = ~new_n5419 & new_n5436;
  assign new_n5439 = ~new_n5386 & ~new_n5387;
  assign new_n5440 = ~new_n5396 & ~new_n5439;
  assign new_n5441 = new_n5396 & new_n5439;
  assign new_n5442 = ~new_n5440 & ~new_n5441;
  assign new_n5443 = ~new_n5438 & ~new_n5442;
  assign new_n5444 = ~new_n5437 & ~new_n5443;
  assign new_n5445 = ~new_n5418 & ~new_n5444;
  assign new_n5446 = new_n5418 & new_n5444;
  assign new_n5447 = ~new_n5445 & ~new_n5446;
  assign new_n5448 = new_n5372 & new_n5447;
  assign new_n5449 = ~new_n5422 & ~new_n5426;
  assign new_n5450 = n1067 & n4805;
  assign new_n5451 = n5645 & n11478;
  assign new_n5452 = new_n5450 & new_n5451;
  assign new_n5453 = ~new_n5449 & new_n5452;
  assign new_n5454 = ~new_n5429 & ~new_n5430;
  assign new_n5455 = new_n5434 & ~new_n5454;
  assign new_n5456 = ~new_n5434 & new_n5454;
  assign new_n5457 = ~new_n5455 & ~new_n5456;
  assign new_n5458 = new_n5453 & new_n5457;
  assign new_n5459 = ~new_n5437 & ~new_n5438;
  assign new_n5460 = new_n5442 & ~new_n5459;
  assign new_n5461 = ~new_n5442 & new_n5459;
  assign new_n5462 = ~new_n5460 & ~new_n5461;
  assign new_n5463 = new_n5458 & new_n5462;
  assign new_n5464 = ~new_n5372 & ~new_n5447;
  assign new_n5465 = ~new_n5448 & ~new_n5464;
  assign new_n5466 = new_n5463 & new_n5465;
  assign new_n5467 = ~new_n5448 & ~new_n5466;
  assign new_n5468 = ~new_n5399 & ~new_n5415;
  assign new_n5469 = ~new_n5376 & ~new_n5468;
  assign new_n5470 = ~new_n5400 & new_n5469;
  assign new_n5471 = new_n5376 & new_n5468;
  assign new_n5472 = ~new_n5470 & ~new_n5471;
  assign new_n5473 = n2551 & n5283;
  assign new_n5474 = n4094 & n4805;
  assign new_n5475 = n11478 & n12826;
  assign new_n5476 = ~new_n5474 & ~new_n5475;
  assign new_n5477 = new_n5474 & new_n5475;
  assign new_n5478 = ~new_n5476 & ~new_n5477;
  assign new_n5479 = new_n5473 & ~new_n5478;
  assign new_n5480 = ~new_n5473 & new_n5478;
  assign new_n5481 = ~new_n5479 & ~new_n5480;
  assign new_n5482 = ~new_n5408 & new_n5412;
  assign new_n5483 = ~new_n5409 & ~new_n5482;
  assign new_n5484 = ~new_n5481 & new_n5483;
  assign new_n5485 = new_n5481 & ~new_n5483;
  assign new_n5486 = ~new_n5484 & ~new_n5485;
  assign new_n5487 = n137 & n11922;
  assign new_n5488 = ~new_n5406 & ~new_n5487;
  assign new_n5489 = new_n5406 & new_n5487;
  assign new_n5490 = ~new_n5488 & ~new_n5489;
  assign new_n5491 = n1067 & n6797;
  assign new_n5492 = n6294 & n8665;
  assign new_n5493 = n3146 & n5645;
  assign new_n5494 = ~new_n5492 & ~new_n5493;
  assign new_n5495 = new_n5492 & new_n5493;
  assign new_n5496 = ~new_n5494 & ~new_n5495;
  assign new_n5497 = ~new_n5491 & ~new_n5496;
  assign new_n5498 = new_n5491 & new_n5496;
  assign new_n5499 = ~new_n5497 & ~new_n5498;
  assign new_n5500 = new_n5490 & ~new_n5499;
  assign new_n5501 = ~new_n5490 & new_n5499;
  assign new_n5502 = ~new_n5500 & ~new_n5501;
  assign new_n5503 = ~new_n5486 & ~new_n5502;
  assign new_n5504 = new_n5486 & new_n5502;
  assign new_n5505 = ~new_n5503 & ~new_n5504;
  assign new_n5506 = ~new_n5472 & new_n5505;
  assign new_n5507 = new_n5472 & ~new_n5505;
  assign new_n5508 = ~new_n5506 & ~new_n5507;
  assign new_n5509 = new_n5445 & new_n5508;
  assign new_n5510 = ~new_n5445 & ~new_n5508;
  assign new_n5511 = ~new_n5509 & ~new_n5510;
  assign new_n5512 = ~new_n5467 & new_n5511;
  assign new_n5513 = new_n5467 & ~new_n5511;
  assign new_n5514 = ~new_n5512 & ~new_n5513;
  assign new_n5515 = ~new_n5052 & new_n5077;
  assign new_n5516 = ~new_n5078 & ~new_n5515;
  assign new_n5517 = new_n5514 & new_n5516;
  assign new_n5518 = ~new_n5514 & ~new_n5516;
  assign new_n5519 = ~new_n5517 & ~new_n5518;
  assign new_n5520 = ~new_n5463 & ~new_n5465;
  assign new_n5521 = ~new_n5466 & ~new_n5520;
  assign new_n5522 = ~new_n5073 & ~new_n5075;
  assign new_n5523 = ~new_n5076 & ~new_n5522;
  assign new_n5524 = new_n5521 & new_n5523;
  assign new_n5525 = ~new_n5521 & ~new_n5523;
  assign new_n5526 = ~new_n5068 & new_n5072;
  assign new_n5527 = ~new_n5073 & ~new_n5526;
  assign new_n5528 = ~new_n5453 & ~new_n5457;
  assign new_n5529 = ~new_n5458 & ~new_n5528;
  assign new_n5530 = ~new_n5063 & new_n5067;
  assign new_n5531 = ~new_n5068 & ~new_n5530;
  assign new_n5532 = new_n5529 & new_n5531;
  assign new_n5533 = ~new_n5529 & ~new_n5531;
  assign new_n5534 = ~new_n5421 & new_n5423;
  assign new_n5535 = ~new_n5449 & ~new_n5534;
  assign new_n5536 = ~new_n5426 & new_n5534;
  assign new_n5537 = ~new_n5535 & ~new_n5536;
  assign new_n5538 = ~new_n4949 & ~new_n5057;
  assign new_n5539 = ~new_n5058 & ~new_n5538;
  assign new_n5540 = ~new_n5450 & ~new_n5451;
  assign new_n5541 = ~new_n5452 & ~new_n5540;
  assign new_n5542 = ~new_n5539 & ~new_n5541;
  assign new_n5543 = new_n5539 & new_n5541;
  assign new_n5544 = n7236 & n11876;
  assign new_n5545 = new_n5421 & new_n5544;
  assign new_n5546 = ~new_n5543 & ~new_n5545;
  assign new_n5547 = ~new_n5542 & ~new_n5546;
  assign new_n5548 = new_n5537 & new_n5547;
  assign new_n5549 = ~new_n5537 & ~new_n5547;
  assign new_n5550 = ~new_n5058 & ~new_n5062;
  assign new_n5551 = ~new_n5063 & ~new_n5550;
  assign new_n5552 = ~new_n5549 & new_n5551;
  assign new_n5553 = ~new_n5548 & ~new_n5552;
  assign new_n5554 = ~new_n5533 & ~new_n5553;
  assign new_n5555 = ~new_n5532 & ~new_n5554;
  assign new_n5556 = new_n5527 & ~new_n5555;
  assign new_n5557 = ~new_n5527 & new_n5555;
  assign new_n5558 = ~new_n5458 & ~new_n5462;
  assign new_n5559 = ~new_n5463 & ~new_n5558;
  assign new_n5560 = ~new_n5557 & new_n5559;
  assign new_n5561 = ~new_n5556 & ~new_n5560;
  assign new_n5562 = ~new_n5525 & ~new_n5561;
  assign new_n5563 = ~new_n5524 & ~new_n5562;
  assign new_n5564 = ~new_n5519 & ~new_n5563;
  assign new_n5565 = new_n5519 & new_n5563;
  assign new_n5566 = ~new_n5564 & ~new_n5565;
  assign new_n5567 = ~new_n5371 & new_n5566;
  assign new_n5568 = ~new_n5364 & ~new_n5366;
  assign new_n5569 = ~new_n5367 & ~new_n5568;
  assign new_n5570 = ~new_n5524 & ~new_n5525;
  assign new_n5571 = new_n5561 & ~new_n5570;
  assign new_n5572 = ~new_n5561 & new_n5570;
  assign new_n5573 = ~new_n5571 & ~new_n5572;
  assign new_n5574 = new_n5569 & new_n5573;
  assign new_n5575 = ~new_n5569 & ~new_n5573;
  assign new_n5576 = ~new_n5359 & ~new_n5363;
  assign new_n5577 = ~new_n5364 & ~new_n5576;
  assign new_n5578 = ~new_n5354 & ~new_n5358;
  assign new_n5579_1 = ~new_n5359 & ~new_n5578;
  assign new_n5580 = ~new_n5532 & ~new_n5533;
  assign new_n5581 = new_n5553 & ~new_n5580;
  assign new_n5582 = ~new_n5553 & new_n5580;
  assign new_n5583 = ~new_n5581 & ~new_n5582;
  assign new_n5584 = ~new_n5579_1 & ~new_n5583;
  assign new_n5585 = new_n5579_1 & new_n5583;
  assign new_n5586 = ~new_n5349 & ~new_n5353;
  assign new_n5587 = ~new_n5354 & ~new_n5586;
  assign new_n5588 = ~new_n5548 & ~new_n5549;
  assign new_n5589 = ~new_n5551 & ~new_n5588;
  assign new_n5590 = new_n5551 & new_n5588;
  assign new_n5591 = ~new_n5589 & ~new_n5590;
  assign new_n5592 = ~new_n5587 & ~new_n5591;
  assign new_n5593 = new_n5587 & new_n5591;
  assign new_n5594 = ~new_n5347 & ~new_n5348;
  assign new_n5595 = ~new_n5349 & ~new_n5594;
  assign new_n5596 = ~new_n5542 & ~new_n5543;
  assign new_n5597 = ~new_n5545 & new_n5596;
  assign new_n5598 = new_n5545 & ~new_n5596;
  assign new_n5599 = ~new_n5597 & ~new_n5598;
  assign new_n5600 = ~new_n5595 & new_n5599;
  assign new_n5601 = new_n5595 & ~new_n5599;
  assign new_n5602 = n6703 & n6877;
  assign new_n5603 = ~new_n5421 & ~new_n5544;
  assign new_n5604 = ~new_n5545 & ~new_n5603;
  assign new_n5605 = new_n5602 & new_n5604;
  assign new_n5606 = ~new_n5601 & ~new_n5605;
  assign new_n5607 = ~new_n5600 & ~new_n5606;
  assign new_n5608 = ~new_n5593 & ~new_n5607;
  assign new_n5609 = ~new_n5592 & ~new_n5608;
  assign new_n5610 = ~new_n5585 & ~new_n5609;
  assign new_n5611 = ~new_n5584 & ~new_n5610;
  assign new_n5612 = new_n5577 & new_n5611;
  assign new_n5613 = ~new_n5577 & ~new_n5611;
  assign new_n5614 = ~new_n5556 & ~new_n5557;
  assign new_n5615 = ~new_n5559 & ~new_n5614;
  assign new_n5616 = new_n5559 & new_n5614;
  assign new_n5617 = ~new_n5615 & ~new_n5616;
  assign new_n5618 = ~new_n5613 & new_n5617;
  assign new_n5619 = ~new_n5612 & ~new_n5618;
  assign new_n5620 = ~new_n5575 & ~new_n5619;
  assign new_n5621 = ~new_n5574 & ~new_n5620;
  assign new_n5622 = new_n5567 & new_n5621;
  assign new_n5623 = new_n5371 & ~new_n5566;
  assign new_n5624 = ~new_n5621 & new_n5623;
  assign new_n5625 = ~new_n5567 & ~new_n5621;
  assign new_n5626 = ~new_n5623 & ~new_n5625;
  assign new_n5627 = ~new_n5624 & ~new_n5626;
  assign new_n5628 = ~new_n5622 & ~new_n5627;
  assign new_n5629 = ~new_n5224 & ~new_n5628;
  assign new_n5630 = new_n5224 & new_n5628;
  assign new_n5631 = ~new_n5217 & ~new_n5219;
  assign new_n5632 = ~new_n5220 & ~new_n5631;
  assign new_n5633 = ~new_n5212_1 & ~new_n5216;
  assign new_n5634 = ~new_n5217 & ~new_n5633;
  assign new_n5635 = ~new_n5612 & ~new_n5613;
  assign new_n5636 = ~new_n5617 & new_n5635;
  assign new_n5637 = new_n5617 & ~new_n5635;
  assign new_n5638 = ~new_n5636 & ~new_n5637;
  assign new_n5639 = ~new_n5634 & new_n5638;
  assign new_n5640 = new_n5634 & ~new_n5638;
  assign new_n5641_1 = ~new_n5207 & new_n5211;
  assign new_n5642 = ~new_n5212_1 & ~new_n5641_1;
  assign new_n5643 = ~new_n5584 & ~new_n5585;
  assign new_n5644 = new_n5609 & ~new_n5643;
  assign new_n5645_1 = ~new_n5609 & new_n5643;
  assign new_n5646 = ~new_n5644 & ~new_n5645_1;
  assign new_n5647 = new_n5642 & ~new_n5646;
  assign new_n5648 = ~new_n5642 & new_n5646;
  assign new_n5649 = ~new_n5202 & ~new_n5206;
  assign new_n5650 = ~new_n5207 & ~new_n5649;
  assign new_n5651 = ~new_n5592 & ~new_n5593;
  assign new_n5652 = new_n5607 & ~new_n5651;
  assign new_n5653 = ~new_n5607 & new_n5651;
  assign new_n5654 = ~new_n5652 & ~new_n5653;
  assign new_n5655 = new_n5650 & ~new_n5654;
  assign new_n5656 = ~new_n5650 & new_n5654;
  assign new_n5657 = n1798 & n7862;
  assign new_n5658 = ~new_n5602 & ~new_n5604;
  assign new_n5659 = ~new_n5605 & ~new_n5658;
  assign new_n5660 = new_n5657 & new_n5659;
  assign new_n5661 = ~new_n5200 & ~new_n5201;
  assign new_n5662 = ~new_n5202 & ~new_n5661;
  assign new_n5663 = new_n5660 & new_n5662;
  assign new_n5664 = ~new_n5660 & ~new_n5662;
  assign new_n5665 = ~new_n5600 & ~new_n5601;
  assign new_n5666 = ~new_n5605 & new_n5665;
  assign new_n5667 = new_n5605 & ~new_n5665;
  assign new_n5668 = ~new_n5666 & ~new_n5667;
  assign new_n5669 = ~new_n5664 & ~new_n5668;
  assign new_n5670_1 = ~new_n5663 & ~new_n5669;
  assign new_n5671 = ~new_n5656 & ~new_n5670_1;
  assign new_n5672 = ~new_n5655 & ~new_n5671;
  assign new_n5673 = ~new_n5648 & ~new_n5672;
  assign new_n5674 = ~new_n5647 & ~new_n5673;
  assign new_n5675 = ~new_n5640 & new_n5674;
  assign new_n5676 = ~new_n5639 & ~new_n5675;
  assign new_n5677 = ~new_n5632 & ~new_n5676;
  assign new_n5678 = new_n5632 & new_n5676;
  assign new_n5679 = ~new_n5574 & ~new_n5575;
  assign new_n5680 = new_n5619 & ~new_n5679;
  assign new_n5681 = ~new_n5619 & new_n5679;
  assign new_n5682 = ~new_n5680 & ~new_n5681;
  assign new_n5683 = ~new_n5678 & ~new_n5682;
  assign new_n5684 = ~new_n5677 & ~new_n5683;
  assign new_n5685 = ~new_n5630 & ~new_n5684;
  assign new_n5686 = ~new_n5629 & ~new_n5685;
  assign new_n5687 = ~new_n5518 & ~new_n5563;
  assign new_n5688 = ~new_n5517 & ~new_n5687;
  assign new_n5689 = n10451 & n11311;
  assign new_n5690 = ~new_n5318 & ~new_n5322;
  assign new_n5691 = ~new_n5321 & ~new_n5690;
  assign new_n5692 = ~new_n5689 & new_n5691;
  assign new_n5693_1 = new_n5689 & ~new_n5691;
  assign new_n5694_1 = ~new_n5692 & ~new_n5693_1;
  assign new_n5695 = ~new_n5316 & ~new_n5326;
  assign new_n5696 = ~new_n5315 & ~new_n5695;
  assign new_n5697 = n3022 & n4203;
  assign new_n5698 = n4187 & n11023;
  assign new_n5699 = ~new_n5697 & new_n5698;
  assign new_n5700 = new_n5697 & ~new_n5698;
  assign new_n5701 = ~new_n5699 & ~new_n5700;
  assign new_n5702 = n9400 & n11423;
  assign new_n5703 = n2464 & n10278;
  assign new_n5704 = ~new_n5702 & new_n5703;
  assign new_n5705 = new_n5702 & ~new_n5703;
  assign new_n5706 = ~new_n5704 & ~new_n5705;
  assign new_n5707 = ~new_n5701 & ~new_n5706;
  assign new_n5708 = new_n5701 & new_n5706;
  assign new_n5709 = ~new_n5707 & ~new_n5708;
  assign new_n5710 = new_n5696 & new_n5709;
  assign new_n5711 = ~new_n5696 & ~new_n5709;
  assign new_n5712 = ~new_n5710 & ~new_n5711;
  assign new_n5713 = new_n5694_1 & ~new_n5712;
  assign new_n5714 = ~new_n5694_1 & new_n5712;
  assign new_n5715 = ~new_n5713 & ~new_n5714;
  assign new_n5716 = ~new_n5334 & ~new_n5715;
  assign new_n5717 = new_n5334 & new_n5715;
  assign new_n5718 = ~new_n5716 & ~new_n5717;
  assign new_n5719 = new_n5688 & ~new_n5718;
  assign new_n5720 = ~new_n5688 & new_n5718;
  assign new_n5721 = ~new_n5719 & ~new_n5720;
  assign new_n5722 = ~new_n5341 & ~new_n5370;
  assign new_n5723 = n6703 & n10174;
  assign new_n5724 = n2278 & n6877;
  assign new_n5725 = n9640 & n12753;
  assign new_n5726 = ~new_n5724 & new_n5725;
  assign new_n5727 = new_n5724 & ~new_n5725;
  assign new_n5728 = ~new_n5726 & ~new_n5727;
  assign new_n5729 = new_n5723 & new_n5728;
  assign new_n5730 = ~new_n5723 & ~new_n5728;
  assign new_n5731 = ~new_n5729 & ~new_n5730;
  assign new_n5732 = new_n5167 & ~new_n5180;
  assign new_n5733 = ~new_n5179 & ~new_n5732;
  assign new_n5734 = ~new_n5168 & ~new_n5172;
  assign new_n5735 = ~new_n5171 & ~new_n5734;
  assign new_n5736 = ~new_n5733 & new_n5735;
  assign new_n5737 = new_n5733 & ~new_n5735;
  assign new_n5738 = ~new_n5736 & ~new_n5737;
  assign new_n5739 = n11821 & n12591;
  assign new_n5740 = n3932 & n9080;
  assign new_n5741 = new_n5739 & new_n5740;
  assign new_n5742 = ~new_n5739 & ~new_n5740;
  assign new_n5743 = ~new_n5741 & ~new_n5742;
  assign new_n5744 = new_n5738 & ~new_n5743;
  assign new_n5745 = ~new_n5738 & new_n5743;
  assign new_n5746 = ~new_n5744 & ~new_n5745;
  assign new_n5747 = ~new_n5731 & new_n5746;
  assign new_n5748 = new_n5731 & ~new_n5746;
  assign new_n5749 = ~new_n5747 & ~new_n5748;
  assign new_n5750 = ~new_n5299 & new_n5336;
  assign new_n5751 = ~new_n5300 & ~new_n5750;
  assign new_n5752 = ~new_n5154 & ~new_n5164;
  assign new_n5753 = ~new_n5153_1 & ~new_n5752;
  assign new_n5754 = n11662 & n11757;
  assign new_n5755 = n3172 & n10327;
  assign new_n5756 = n1333 & n9583;
  assign new_n5757 = ~new_n5755 & new_n5756;
  assign new_n5758 = new_n5755 & ~new_n5756;
  assign new_n5759 = ~new_n5757 & ~new_n5758;
  assign new_n5760_1 = new_n5754 & new_n5759;
  assign new_n5761 = ~new_n5754 & ~new_n5759;
  assign new_n5762 = ~new_n5760_1 & ~new_n5761;
  assign new_n5763 = ~new_n5156 & ~new_n5160;
  assign new_n5764 = ~new_n5159 & ~new_n5763;
  assign new_n5765 = n5240 & n7456;
  assign new_n5766 = new_n5764 & ~new_n5765;
  assign new_n5767_1 = ~new_n5764 & new_n5765;
  assign new_n5768 = ~new_n5766 & ~new_n5767_1;
  assign new_n5769 = new_n5762 & ~new_n5768;
  assign new_n5770 = ~new_n5762 & new_n5768;
  assign new_n5771 = ~new_n5769 & ~new_n5770;
  assign new_n5772 = ~new_n5753 & new_n5771;
  assign new_n5773 = new_n5753 & ~new_n5771;
  assign new_n5774 = ~new_n5772 & ~new_n5773;
  assign new_n5775 = ~new_n5751 & ~new_n5774;
  assign new_n5776 = new_n5751 & new_n5774;
  assign new_n5777 = ~new_n5775 & ~new_n5776;
  assign new_n5778 = ~new_n5749 & new_n5777;
  assign new_n5779 = new_n5749 & ~new_n5777;
  assign new_n5780 = ~new_n5778 & ~new_n5779;
  assign new_n5781 = new_n5722 & new_n5780;
  assign new_n5782 = ~new_n5722 & ~new_n5780;
  assign new_n5783 = ~new_n5781 & ~new_n5782;
  assign new_n5784 = new_n5721 & ~new_n5783;
  assign new_n5785 = ~new_n5721 & new_n5783;
  assign new_n5786 = ~new_n5784 & ~new_n5785;
  assign new_n5787 = ~new_n5509 & ~new_n5512;
  assign new_n5788 = ~new_n5470 & ~new_n5505;
  assign new_n5789 = ~new_n5471 & ~new_n5788;
  assign new_n5790 = n137 & n2551;
  assign new_n5791 = n6294 & n11922;
  assign new_n5792 = ~new_n5790 & ~new_n5791;
  assign new_n5793 = new_n5790 & new_n5791;
  assign new_n5794 = ~new_n5792 & ~new_n5793;
  assign new_n5795 = n6797 & n8665;
  assign new_n5796 = n1067 & n3146;
  assign new_n5797 = new_n5795 & ~new_n5796;
  assign new_n5798_1 = ~new_n5795 & new_n5796;
  assign new_n5799 = ~new_n5797 & ~new_n5798_1;
  assign new_n5800 = ~new_n5794 & ~new_n5799;
  assign new_n5801 = new_n5794 & new_n5799;
  assign new_n5802 = ~new_n5800 & ~new_n5801;
  assign new_n5803 = new_n5789 & ~new_n5802;
  assign new_n5804 = ~new_n5789 & new_n5802;
  assign new_n5805 = ~new_n5803 & ~new_n5804;
  assign new_n5806 = n3992 & n12247;
  assign new_n5807 = n159 & n6358;
  assign new_n5808 = n2749 & n5198;
  assign new_n5809 = ~new_n5807 & new_n5808;
  assign new_n5810 = new_n5807 & ~new_n5808;
  assign new_n5811 = ~new_n5809 & ~new_n5810;
  assign new_n5812 = new_n5806 & new_n5811;
  assign new_n5813 = ~new_n5806 & ~new_n5811;
  assign new_n5814_1 = ~new_n5812 & ~new_n5813;
  assign new_n5815 = ~new_n5015 & ~new_n5019;
  assign new_n5816 = ~new_n5018 & ~new_n5815;
  assign new_n5817 = ~new_n5814_1 & new_n5816;
  assign new_n5818 = new_n5814_1 & ~new_n5816;
  assign new_n5819 = ~new_n5817 & ~new_n5818;
  assign new_n5820 = ~new_n5033 & ~new_n5036;
  assign new_n5821 = ~new_n5035 & ~new_n5820;
  assign new_n5822 = n1510 & n8384;
  assign new_n5823 = n4805 & n10685;
  assign new_n5824 = n4938 & n5645;
  assign new_n5825 = new_n5823 & ~new_n5824;
  assign new_n5826 = ~new_n5823 & new_n5824;
  assign new_n5827 = ~new_n5825 & ~new_n5826;
  assign new_n5828 = new_n5822 & ~new_n5827;
  assign new_n5829 = ~new_n5822 & new_n5827;
  assign new_n5830 = ~new_n5828 & ~new_n5829;
  assign new_n5831 = ~new_n5821 & ~new_n5830;
  assign new_n5832 = new_n5821 & new_n5830;
  assign new_n5833 = ~new_n5831 & ~new_n5832;
  assign new_n5834 = ~new_n5819 & new_n5833;
  assign new_n5835 = new_n5819 & ~new_n5833;
  assign new_n5836 = ~new_n5834 & ~new_n5835;
  assign new_n5837 = ~new_n5026 & ~new_n5043;
  assign new_n5838 = ~new_n5027 & ~new_n5837;
  assign new_n5839 = ~new_n5031 & ~new_n5040;
  assign new_n5840 = ~new_n5030_1 & ~new_n5839;
  assign new_n5841 = new_n5838 & new_n5840;
  assign new_n5842 = ~new_n5838 & ~new_n5840;
  assign new_n5843 = ~new_n5841 & ~new_n5842;
  assign new_n5844 = new_n5836 & ~new_n5843;
  assign new_n5845 = ~new_n5836 & new_n5843;
  assign new_n5846 = ~new_n5844 & ~new_n5845;
  assign new_n5847 = ~new_n5805 & ~new_n5846;
  assign new_n5848 = new_n5805 & new_n5846;
  assign new_n5849 = ~new_n5847 & ~new_n5848;
  assign new_n5850 = new_n5473 & ~new_n5476;
  assign new_n5851 = ~new_n5477 & ~new_n5850;
  assign new_n5852 = ~new_n5485 & ~new_n5502;
  assign new_n5853 = ~new_n5484 & ~new_n5852;
  assign new_n5854 = new_n5851 & new_n5853;
  assign new_n5855 = ~new_n5851 & ~new_n5853;
  assign new_n5856 = ~new_n5854 & ~new_n5855;
  assign new_n5857_1 = ~new_n5849 & new_n5856;
  assign new_n5858 = new_n5849 & ~new_n5856;
  assign new_n5859 = ~new_n5857_1 & ~new_n5858;
  assign new_n5860_1 = new_n5787 & ~new_n5859;
  assign new_n5861 = ~new_n5787 & new_n5859;
  assign new_n5862 = ~new_n5860_1 & ~new_n5861;
  assign new_n5863 = ~new_n5302 & ~new_n5306;
  assign new_n5864 = ~new_n5305_1 & ~new_n5863;
  assign new_n5865 = n1471 & n3754;
  assign new_n5866 = n7646 & n10898;
  assign new_n5867 = ~new_n5865 & ~new_n5866;
  assign new_n5868 = new_n5865 & new_n5866;
  assign new_n5869 = ~new_n5867 & ~new_n5868;
  assign new_n5870 = n7236 & n12511;
  assign new_n5871 = n4722 & n11876;
  assign new_n5872 = new_n5870 & ~new_n5871;
  assign new_n5873 = ~new_n5870 & new_n5871;
  assign new_n5874 = ~new_n5872 & ~new_n5873;
  assign new_n5875 = ~new_n5869 & ~new_n5874;
  assign new_n5876 = new_n5869 & new_n5874;
  assign new_n5877 = ~new_n5875 & ~new_n5876;
  assign new_n5878 = ~new_n5864 & new_n5877;
  assign new_n5879 = new_n5864 & ~new_n5877;
  assign new_n5880 = ~new_n5878 & ~new_n5879;
  assign new_n5881 = ~new_n5862 & new_n5880;
  assign new_n5882 = new_n5862 & ~new_n5880;
  assign new_n5883 = ~new_n5881 & ~new_n5882;
  assign new_n5884 = ~new_n5012 & new_n5046;
  assign new_n5885 = ~new_n5013 & ~new_n5884;
  assign new_n5886 = ~new_n5193 & ~new_n5222;
  assign new_n5887 = new_n5184 & ~new_n5188;
  assign new_n5888 = ~new_n5186 & ~new_n5887;
  assign new_n5889 = ~new_n5491 & ~new_n5495;
  assign new_n5890 = ~new_n5494 & ~new_n5889;
  assign new_n5891 = n4094 & n11478;
  assign new_n5892 = n5283 & n12826;
  assign new_n5893 = ~new_n5891 & new_n5892;
  assign new_n5894 = new_n5891 & ~new_n5892;
  assign new_n5895 = ~new_n5893 & ~new_n5894;
  assign new_n5896 = ~new_n5890 & ~new_n5895;
  assign new_n5897 = new_n5890 & new_n5895;
  assign new_n5898 = ~new_n5896 & ~new_n5897;
  assign new_n5899 = ~new_n5488 & new_n5499;
  assign new_n5900 = ~new_n5489 & ~new_n5899;
  assign new_n5901 = ~new_n5898 & ~new_n5900;
  assign new_n5902 = new_n5898 & new_n5900;
  assign new_n5903 = ~new_n5901 & ~new_n5902;
  assign new_n5904 = n753 & n7862;
  assign new_n5905 = n1798 & n6826;
  assign new_n5906 = ~new_n5904 & new_n5905;
  assign new_n5907 = new_n5904 & ~new_n5905;
  assign new_n5908 = ~new_n5906 & ~new_n5907;
  assign new_n5909 = ~new_n5903 & new_n5908;
  assign new_n5910 = new_n5903 & ~new_n5908;
  assign new_n5911 = ~new_n5909 & ~new_n5910;
  assign new_n5912 = new_n5888 & ~new_n5911;
  assign new_n5913 = ~new_n5888 & new_n5911;
  assign new_n5914 = ~new_n5912 & ~new_n5913;
  assign new_n5915 = new_n5886 & ~new_n5914;
  assign new_n5916 = ~new_n5886 & new_n5914;
  assign new_n5917 = ~new_n5915 & ~new_n5916;
  assign new_n5918 = new_n5885 & new_n5917;
  assign new_n5919 = ~new_n5885 & ~new_n5917;
  assign new_n5920 = ~new_n5918 & ~new_n5919;
  assign new_n5921 = new_n5883 & new_n5920;
  assign new_n5922 = ~new_n5883 & ~new_n5920;
  assign new_n5923 = ~new_n5921 & ~new_n5922;
  assign new_n5924 = new_n5626 & ~new_n5923;
  assign new_n5925 = ~new_n5626 & new_n5923;
  assign new_n5926 = ~new_n5924 & ~new_n5925;
  assign new_n5927 = ~new_n5786 & ~new_n5926;
  assign new_n5928 = new_n5786 & new_n5926;
  assign new_n5929 = ~new_n5927 & ~new_n5928;
  assign new_n5930 = ~new_n5686 & new_n5929;
  assign new_n5931 = new_n5686 & ~new_n5929;
  assign new_n5932 = ~new_n5930 & ~new_n5931;
  assign new_n5933 = new_n5079 & new_n5932;
  assign new_n5934_1 = ~new_n5079 & ~new_n5932;
  assign n1269 = ~new_n5933 & ~new_n5934_1;
  assign new_n5936 = n5305 & n9195;
  assign new_n5937 = ~new_n1158 & ~new_n1169;
  assign new_n5938 = ~new_n1159 & ~new_n5937;
  assign new_n5939 = ~new_n5936 & new_n5938;
  assign new_n5940 = new_n5936 & ~new_n5938;
  assign new_n5941 = n7265 & n12705;
  assign new_n5942 = n1097 & n10223;
  assign new_n5943 = n2879 & n4312;
  assign new_n5944 = ~new_n5942 & ~new_n5943;
  assign new_n5945 = new_n5942 & new_n5943;
  assign new_n5946 = ~new_n5944 & ~new_n5945;
  assign new_n5947 = ~new_n5941 & ~new_n5946;
  assign new_n5948 = new_n5941 & new_n5946;
  assign new_n5949 = ~new_n5947 & ~new_n5948;
  assign new_n5950 = n4634 & n5964;
  assign new_n5951 = new_n1161 & ~new_n1164;
  assign new_n5952 = ~new_n1165 & ~new_n5951;
  assign new_n5953 = ~new_n5950 & new_n5952;
  assign new_n5954 = new_n5950 & ~new_n5952;
  assign new_n5955 = ~new_n5953 & ~new_n5954;
  assign new_n5956 = ~new_n5949 & ~new_n5955;
  assign new_n5957 = new_n5949 & new_n5955;
  assign new_n5958 = ~new_n5956 & ~new_n5957;
  assign new_n5959 = ~new_n5940 & ~new_n5958;
  assign new_n5960 = ~new_n5939 & ~new_n5959;
  assign new_n5961 = n5964 & n9195;
  assign new_n5962 = n1097 & n4634;
  assign new_n5963 = ~new_n5961 & ~new_n5962;
  assign new_n5964_1 = new_n5961 & new_n5962;
  assign new_n5965 = ~new_n5963 & ~new_n5964_1;
  assign new_n5966 = n4312 & n10223;
  assign new_n5967 = new_n5941 & ~new_n5944;
  assign new_n5968 = ~new_n1163 & ~new_n5967;
  assign new_n5969 = new_n5966 & ~new_n5968;
  assign new_n5970 = ~new_n5966 & ~new_n5967;
  assign new_n5971 = ~new_n5969 & ~new_n5970;
  assign new_n5972 = n7265 & n12025;
  assign new_n5973 = n2879 & n12705;
  assign new_n5974 = ~new_n5972 & ~new_n5973;
  assign new_n5975 = new_n5972 & new_n5973;
  assign new_n5976 = ~new_n5974 & ~new_n5975;
  assign new_n5977 = ~new_n5971 & new_n5976;
  assign new_n5978 = new_n5971 & ~new_n5976;
  assign new_n5979 = ~new_n5977 & ~new_n5978;
  assign new_n5980 = new_n5965 & ~new_n5979;
  assign new_n5981 = ~new_n5965 & new_n5979;
  assign new_n5982 = ~new_n5980 & ~new_n5981;
  assign new_n5983 = ~new_n5949 & ~new_n5954;
  assign new_n5984 = ~new_n5953 & ~new_n5983;
  assign new_n5985 = new_n5982 & ~new_n5984;
  assign new_n5986 = ~new_n5982 & new_n5984;
  assign new_n5987 = ~new_n5985 & ~new_n5986;
  assign new_n5988 = new_n5960 & ~new_n5987;
  assign new_n5989 = ~new_n5980 & ~new_n5984;
  assign new_n5990 = ~new_n5981 & ~new_n5989;
  assign new_n5991 = ~new_n5964_1 & ~new_n5990;
  assign new_n5992 = new_n5964_1 & new_n5990;
  assign new_n5993 = ~new_n5991 & ~new_n5992;
  assign new_n5994 = n2253 & n5964;
  assign new_n5995 = n1097 & n9195;
  assign new_n5996 = n3865 & n5305;
  assign new_n5997 = ~new_n5995 & ~new_n5996;
  assign new_n5998 = new_n5995 & new_n5996;
  assign new_n5999 = ~new_n5997 & ~new_n5998;
  assign new_n6000 = ~new_n5994 & ~new_n5999;
  assign new_n6001 = new_n5994 & new_n5999;
  assign new_n6002 = ~new_n6000 & ~new_n6001;
  assign new_n6003 = ~new_n5970 & new_n5976;
  assign new_n6004 = ~new_n5969 & ~new_n6003;
  assign new_n6005 = new_n6002 & ~new_n6004;
  assign new_n6006 = ~new_n6002 & new_n6004;
  assign new_n6007 = ~new_n6005 & ~new_n6006;
  assign new_n6008 = n4312 & n4634;
  assign new_n6009 = ~new_n5975 & ~new_n6008;
  assign new_n6010 = new_n5975 & new_n6008;
  assign new_n6011 = ~new_n6009 & ~new_n6010;
  assign new_n6012 = n2879 & n12025;
  assign new_n6013 = n7265 & n11257;
  assign new_n6014 = n10223 & n12705;
  assign new_n6015 = ~new_n6013 & ~new_n6014;
  assign new_n6016_1 = new_n6013 & new_n6014;
  assign new_n6017 = ~new_n6015 & ~new_n6016_1;
  assign new_n6018 = ~new_n6012 & ~new_n6017;
  assign new_n6019 = new_n6012 & new_n6017;
  assign new_n6020 = ~new_n6018 & ~new_n6019;
  assign new_n6021 = new_n6011 & ~new_n6020;
  assign new_n6022 = ~new_n6011 & new_n6020;
  assign new_n6023 = ~new_n6021 & ~new_n6022;
  assign new_n6024 = ~new_n6007 & ~new_n6023;
  assign new_n6025 = new_n6007 & new_n6023;
  assign new_n6026 = ~new_n6024 & ~new_n6025;
  assign new_n6027 = ~new_n5993 & ~new_n6026;
  assign new_n6028 = ~new_n5992 & new_n6026;
  assign new_n6029 = ~new_n5991 & new_n6028;
  assign new_n6030 = ~new_n6027 & ~new_n6029;
  assign new_n6031 = ~new_n5988 & new_n6030;
  assign new_n6032 = new_n5988 & ~new_n6030;
  assign new_n6033 = ~new_n6031 & ~new_n6032;
  assign new_n6034 = n2253 & n5305;
  assign new_n6035 = ~new_n5960 & new_n5987;
  assign new_n6036 = ~new_n5988 & ~new_n6035;
  assign new_n6037 = new_n6034 & new_n6036;
  assign new_n6038_1 = ~new_n5939 & ~new_n5940;
  assign new_n6039 = new_n5958 & ~new_n6038_1;
  assign new_n6040 = ~new_n5958 & new_n6038_1;
  assign new_n6041 = ~new_n6039 & ~new_n6040;
  assign new_n6042 = new_n1173 & ~new_n6041;
  assign new_n6043 = ~new_n6034 & ~new_n6036;
  assign new_n6044 = ~new_n6037 & ~new_n6043;
  assign new_n6045 = new_n6042 & new_n6044;
  assign new_n6046 = ~new_n6037 & ~new_n6045;
  assign new_n6047 = ~new_n6033 & new_n6046;
  assign new_n6048 = new_n6033 & ~new_n6046;
  assign new_n6049 = ~new_n6047 & ~new_n6048;
  assign new_n6050 = ~new_n6042 & ~new_n6044;
  assign new_n6051 = ~new_n6045 & ~new_n6050;
  assign new_n6052 = n8759 & n12145;
  assign new_n6053 = ~new_n1285 & ~new_n1295;
  assign new_n6054 = ~new_n1284 & ~new_n6053;
  assign new_n6055 = new_n6052 & ~new_n6054;
  assign new_n6056 = ~new_n6052 & new_n6054;
  assign new_n6057 = ~new_n6055 & ~new_n6056;
  assign new_n6058 = n7946 & n8276;
  assign new_n6059 = n2024 & n7436;
  assign new_n6060 = ~new_n1182 & ~new_n6059;
  assign new_n6061 = new_n1182 & new_n6059;
  assign new_n6062 = ~new_n6060 & ~new_n6061;
  assign new_n6063 = ~new_n6058 & ~new_n6062;
  assign new_n6064 = new_n6058 & new_n6062;
  assign new_n6065 = ~new_n6063 & ~new_n6064;
  assign new_n6066 = n2522 & n6776;
  assign new_n6067 = new_n1287 & ~new_n1290;
  assign new_n6068 = ~new_n1291 & ~new_n6067;
  assign new_n6069 = ~new_n6066 & new_n6068;
  assign new_n6070 = new_n6066 & ~new_n6068;
  assign new_n6071 = ~new_n6069 & ~new_n6070;
  assign new_n6072 = ~new_n6065 & ~new_n6071;
  assign new_n6073 = new_n6065 & new_n6071;
  assign new_n6074 = ~new_n6072 & ~new_n6073;
  assign new_n6075 = ~new_n6057 & new_n6074;
  assign new_n6076 = new_n6057 & ~new_n6074;
  assign new_n6077 = ~new_n6075 & ~new_n6076;
  assign new_n6078 = new_n1300 & ~new_n6077;
  assign new_n6079 = n8759 & n12221;
  assign new_n6080 = ~new_n6055 & ~new_n6074;
  assign new_n6081 = ~new_n6056 & ~new_n6080;
  assign new_n6082 = n6776 & n12145;
  assign new_n6083 = n2522 & n12299;
  assign new_n6084 = ~new_n6082 & ~new_n6083;
  assign new_n6085 = new_n6082 & new_n6083;
  assign new_n6086 = ~new_n6084 & ~new_n6085;
  assign new_n6087 = ~new_n6065 & ~new_n6070;
  assign new_n6088 = ~new_n6069 & ~new_n6087;
  assign new_n6089_1 = ~new_n6086 & ~new_n6088;
  assign new_n6090 = new_n6086 & new_n6088;
  assign new_n6091 = ~new_n6089_1 & ~new_n6090;
  assign new_n6092 = n7436 & n9189;
  assign new_n6093 = new_n6058 & ~new_n6060;
  assign new_n6094 = ~new_n1289 & ~new_n6093;
  assign new_n6095 = new_n6092 & ~new_n6094;
  assign new_n6096 = ~new_n6092 & ~new_n6093;
  assign new_n6097 = ~new_n6095 & ~new_n6096;
  assign new_n6098 = n2024 & n8276;
  assign new_n6099 = n7946 & n9241;
  assign new_n6100 = ~new_n6098 & ~new_n6099;
  assign new_n6101 = new_n6098 & new_n6099;
  assign new_n6102 = ~new_n6100 & ~new_n6101;
  assign new_n6103 = new_n6097 & ~new_n6102;
  assign new_n6104 = ~new_n6097 & new_n6102;
  assign new_n6105 = ~new_n6103 & ~new_n6104;
  assign new_n6106 = new_n6091 & ~new_n6105;
  assign new_n6107 = ~new_n6091 & new_n6105;
  assign new_n6108 = ~new_n6106 & ~new_n6107;
  assign new_n6109 = new_n6081 & new_n6108;
  assign new_n6110 = ~new_n6081 & ~new_n6108;
  assign new_n6111 = ~new_n6109 & ~new_n6110;
  assign new_n6112 = new_n6079 & new_n6111;
  assign new_n6113 = ~new_n6079 & ~new_n6111;
  assign new_n6114 = ~new_n6112 & ~new_n6113;
  assign new_n6115 = new_n6078 & new_n6114;
  assign new_n6116 = ~new_n6078 & ~new_n6114;
  assign new_n6117 = ~new_n6115 & ~new_n6116;
  assign new_n6118 = ~new_n1300 & new_n6077;
  assign new_n6119 = ~new_n6078 & ~new_n6118;
  assign new_n6120 = n5331 & n6016;
  assign new_n6121 = n521 & n8476;
  assign new_n6122 = new_n1313 & ~new_n1316;
  assign new_n6123 = ~new_n1317 & ~new_n6122;
  assign new_n6124 = new_n6121 & ~new_n6123;
  assign new_n6125 = ~new_n6121 & new_n6123;
  assign new_n6126_1 = ~new_n6124 & ~new_n6125;
  assign new_n6127 = n2558 & n10545;
  assign new_n6128 = n2530 & n5579;
  assign new_n6129 = n2498 & n12648;
  assign new_n6130 = ~new_n6128 & ~new_n6129;
  assign new_n6131 = new_n6128 & new_n6129;
  assign new_n6132 = ~new_n6130 & ~new_n6131;
  assign new_n6133 = new_n6127 & ~new_n6132;
  assign new_n6134 = ~new_n6127 & new_n6132;
  assign new_n6135 = ~new_n6133 & ~new_n6134;
  assign new_n6136 = ~new_n6126_1 & ~new_n6135;
  assign new_n6137 = new_n6126_1 & new_n6135;
  assign new_n6138 = ~new_n6136 & ~new_n6137;
  assign new_n6139 = new_n6120 & ~new_n6138;
  assign new_n6140 = ~new_n6120 & new_n6138;
  assign new_n6141 = ~new_n6139 & ~new_n6140;
  assign new_n6142 = ~new_n1310 & new_n1321;
  assign new_n6143 = ~new_n1311 & ~new_n6142;
  assign new_n6144 = ~new_n6141 & new_n6143;
  assign new_n6145 = new_n6141 & ~new_n6143;
  assign new_n6146 = ~new_n6144 & ~new_n6145;
  assign new_n6147 = new_n1326 & ~new_n6146;
  assign new_n6148 = ~new_n1326 & new_n6146;
  assign new_n6149 = ~new_n6147 & ~new_n6148;
  assign new_n6150 = n7270 & n7965;
  assign new_n6151 = n806 & n7388;
  assign new_n6152 = new_n1334 & ~new_n1337;
  assign new_n6153 = ~new_n1338 & ~new_n6152;
  assign new_n6154 = ~new_n6151 & new_n6153;
  assign new_n6155 = new_n6151 & ~new_n6153;
  assign new_n6156 = ~new_n6154 & ~new_n6155;
  assign new_n6157 = n5860 & n9763;
  assign new_n6158 = n3342 & n11892;
  assign new_n6159 = n2393 & n9111;
  assign new_n6160 = ~new_n6158 & ~new_n6159;
  assign new_n6161 = new_n6158 & new_n6159;
  assign new_n6162 = ~new_n6160 & ~new_n6161;
  assign new_n6163 = new_n6157 & ~new_n6162;
  assign new_n6164 = ~new_n6157 & new_n6162;
  assign new_n6165 = ~new_n6163 & ~new_n6164;
  assign new_n6166 = ~new_n6156 & new_n6165;
  assign new_n6167 = new_n6156 & ~new_n6165;
  assign new_n6168 = ~new_n6166 & ~new_n6167;
  assign new_n6169 = new_n6150 & new_n6168;
  assign new_n6170 = ~new_n6150 & ~new_n6168;
  assign new_n6171 = ~new_n6169 & ~new_n6170;
  assign new_n6172 = ~new_n1331 & new_n1342;
  assign new_n6173 = ~new_n1332 & ~new_n6172;
  assign new_n6174 = ~new_n6171 & new_n6173;
  assign new_n6175 = new_n6171 & ~new_n6173;
  assign new_n6176 = ~new_n6174 & ~new_n6175;
  assign new_n6177 = new_n1346 & ~new_n6176;
  assign new_n6178 = ~new_n1346 & new_n6176;
  assign new_n6179 = ~new_n6177 & ~new_n6178;
  assign new_n6180 = new_n6149 & new_n6179;
  assign new_n6181 = ~new_n6149 & ~new_n6179;
  assign new_n6182 = ~new_n6180 & ~new_n6181;
  assign new_n6183 = new_n1356 & new_n6182;
  assign new_n6184 = ~new_n1356 & ~new_n6182;
  assign new_n6185 = ~new_n6183 & ~new_n6184;
  assign new_n6186 = new_n6119 & ~new_n6185;
  assign new_n6187 = ~new_n6119 & new_n6185;
  assign new_n6188 = ~new_n1305 & new_n1358;
  assign new_n6189 = ~new_n1304 & ~new_n6188;
  assign new_n6190 = ~new_n6187 & ~new_n6189;
  assign new_n6191 = ~new_n6186 & ~new_n6190;
  assign new_n6192_1 = ~new_n6117 & new_n6191;
  assign new_n6193 = new_n6117 & ~new_n6191;
  assign new_n6194 = ~new_n6192_1 & ~new_n6193;
  assign new_n6195 = n5331 & n5798;
  assign new_n6196 = ~new_n6140 & new_n6143;
  assign new_n6197 = ~new_n6139 & ~new_n6196;
  assign new_n6198 = n6016 & n8476;
  assign new_n6199 = n521 & n2530;
  assign new_n6200 = ~new_n6198 & ~new_n6199;
  assign new_n6201 = new_n6198 & new_n6199;
  assign new_n6202 = ~new_n6200 & ~new_n6201;
  assign new_n6203 = n5579 & n12648;
  assign new_n6204 = n2498 & n10545;
  assign new_n6205 = n2558 & n7690;
  assign new_n6206 = ~new_n6204 & ~new_n6205;
  assign new_n6207 = new_n6204 & new_n6205;
  assign new_n6208 = ~new_n6206 & ~new_n6207;
  assign new_n6209 = new_n6203 & new_n6208;
  assign new_n6210 = ~new_n6203 & ~new_n6208;
  assign new_n6211 = ~new_n6209 & ~new_n6210;
  assign new_n6212 = new_n6127 & ~new_n6130;
  assign new_n6213 = ~new_n6131 & ~new_n6212;
  assign new_n6214 = ~new_n6211 & ~new_n6213;
  assign new_n6215 = new_n6211 & new_n6213;
  assign new_n6216 = ~new_n6214 & ~new_n6215;
  assign new_n6217 = new_n6202 & ~new_n6216;
  assign new_n6218 = ~new_n6202 & new_n6216;
  assign new_n6219 = ~new_n6217 & ~new_n6218;
  assign new_n6220 = ~new_n6124 & new_n6135;
  assign new_n6221 = ~new_n6125 & ~new_n6220;
  assign new_n6222 = ~new_n6219 & new_n6221;
  assign new_n6223 = new_n6219 & ~new_n6221;
  assign new_n6224 = ~new_n6222 & ~new_n6223;
  assign new_n6225 = ~new_n6197 & ~new_n6224;
  assign new_n6226 = new_n6197 & new_n6224;
  assign new_n6227 = ~new_n6225 & ~new_n6226;
  assign new_n6228 = new_n6195 & new_n6227;
  assign new_n6229 = ~new_n6195 & ~new_n6227;
  assign new_n6230 = ~new_n6228 & ~new_n6229;
  assign new_n6231 = new_n6147 & new_n6230;
  assign new_n6232 = ~new_n6147 & ~new_n6230;
  assign new_n6233 = ~new_n6231 & ~new_n6232;
  assign new_n6234 = n5153 & n7965;
  assign new_n6235 = ~new_n6170 & new_n6173;
  assign new_n6236 = ~new_n6169 & ~new_n6235;
  assign new_n6237 = n7270 & n7388;
  assign new_n6238 = n806 & n11892;
  assign new_n6239 = ~new_n6237 & ~new_n6238;
  assign new_n6240 = new_n6237 & new_n6238;
  assign new_n6241 = ~new_n6239 & ~new_n6240;
  assign new_n6242 = n2393 & n3342;
  assign new_n6243 = n3986 & n9763;
  assign new_n6244 = n5860 & n9111;
  assign new_n6245 = ~new_n6243 & ~new_n6244;
  assign new_n6246 = new_n6243 & new_n6244;
  assign new_n6247 = ~new_n6245 & ~new_n6246;
  assign new_n6248 = new_n6242 & new_n6247;
  assign new_n6249 = ~new_n6242 & ~new_n6247;
  assign new_n6250 = ~new_n6248 & ~new_n6249;
  assign new_n6251 = ~new_n6157 & ~new_n6161;
  assign new_n6252 = ~new_n6160 & ~new_n6251;
  assign new_n6253 = ~new_n6250 & new_n6252;
  assign new_n6254_1 = new_n6250 & ~new_n6252;
  assign new_n6255 = ~new_n6253 & ~new_n6254_1;
  assign new_n6256 = new_n6241 & ~new_n6255;
  assign new_n6257 = ~new_n6241 & new_n6255;
  assign new_n6258 = ~new_n6256 & ~new_n6257;
  assign new_n6259 = ~new_n6154 & ~new_n6165;
  assign new_n6260 = ~new_n6155 & ~new_n6259;
  assign new_n6261 = new_n6258 & new_n6260;
  assign new_n6262 = ~new_n6258 & ~new_n6260;
  assign new_n6263 = ~new_n6261 & ~new_n6262;
  assign new_n6264 = ~new_n6236 & ~new_n6263;
  assign new_n6265 = new_n6236 & new_n6263;
  assign new_n6266 = ~new_n6264 & ~new_n6265;
  assign new_n6267 = new_n6234 & new_n6266;
  assign new_n6268 = ~new_n6234 & ~new_n6266;
  assign new_n6269 = ~new_n6267 & ~new_n6268;
  assign new_n6270 = new_n6177 & new_n6269;
  assign new_n6271 = ~new_n6177 & ~new_n6269;
  assign new_n6272 = ~new_n6270 & ~new_n6271;
  assign new_n6273_1 = ~new_n6233 & ~new_n6272;
  assign new_n6274 = ~new_n1356 & ~new_n6181;
  assign new_n6275 = ~new_n6180 & ~new_n6274;
  assign new_n6276 = new_n6273_1 & new_n6275;
  assign new_n6277 = new_n6233 & new_n6272;
  assign new_n6278 = ~new_n6275 & new_n6277;
  assign new_n6279 = ~new_n6273_1 & ~new_n6275;
  assign new_n6280 = ~new_n6277 & ~new_n6279;
  assign new_n6281 = ~new_n6278 & ~new_n6280;
  assign new_n6282 = ~new_n6276 & ~new_n6281;
  assign new_n6283 = ~new_n6194 & ~new_n6282;
  assign new_n6284 = new_n6194 & new_n6282;
  assign new_n6285 = ~new_n6283 & ~new_n6284;
  assign new_n6286 = new_n6051 & new_n6285;
  assign new_n6287 = ~new_n6051 & ~new_n6285;
  assign new_n6288 = ~new_n1173 & new_n6041;
  assign new_n6289 = ~new_n6042 & ~new_n6288;
  assign new_n6290 = new_n6186 & ~new_n6189;
  assign new_n6291 = new_n6187 & new_n6189;
  assign new_n6292 = new_n6191 & ~new_n6291;
  assign new_n6293 = ~new_n6290 & ~new_n6292;
  assign new_n6294_1 = ~new_n6289 & new_n6293;
  assign new_n6295 = new_n6289 & ~new_n6293;
  assign new_n6296 = ~new_n1279 & ~new_n1361;
  assign new_n6297 = ~new_n1278 & ~new_n6296;
  assign new_n6298 = ~new_n6295 & new_n6297;
  assign new_n6299 = ~new_n6294_1 & ~new_n6298;
  assign new_n6300 = ~new_n6287 & new_n6299;
  assign new_n6301 = ~new_n6286 & ~new_n6300;
  assign new_n6302 = new_n6049 & ~new_n6301;
  assign new_n6303 = ~new_n6049 & new_n6301;
  assign new_n6304 = ~new_n6302 & ~new_n6303;
  assign new_n6305 = ~new_n6112 & ~new_n6115;
  assign new_n6306 = ~new_n6090 & new_n6105;
  assign new_n6307 = ~new_n6089_1 & ~new_n6306;
  assign new_n6308 = ~new_n6085 & ~new_n6307;
  assign new_n6309 = new_n6085 & new_n6307;
  assign new_n6310 = ~new_n6308 & ~new_n6309;
  assign new_n6311 = n6776 & n12221;
  assign new_n6312 = n12145 & n12299;
  assign new_n6313 = n8759 & n10217;
  assign new_n6314 = ~new_n6312 & ~new_n6313;
  assign new_n6315 = new_n6312 & new_n6313;
  assign new_n6316 = ~new_n6314 & ~new_n6315;
  assign new_n6317 = ~new_n6311 & ~new_n6316;
  assign new_n6318 = new_n6311 & new_n6316;
  assign new_n6319 = ~new_n6317 & ~new_n6318;
  assign new_n6320 = ~new_n6096 & new_n6102;
  assign new_n6321 = ~new_n6095 & ~new_n6320;
  assign new_n6322 = new_n6319 & ~new_n6321;
  assign new_n6323 = ~new_n6319 & new_n6321;
  assign new_n6324 = ~new_n6322 & ~new_n6323;
  assign new_n6325 = n2522 & n7436;
  assign new_n6326 = new_n6101 & new_n6325;
  assign new_n6327 = ~new_n6101 & ~new_n6325;
  assign new_n6328 = ~new_n6326 & ~new_n6327;
  assign new_n6329 = n7946 & n10510;
  assign new_n6330 = n2024 & n9241;
  assign new_n6331 = n8276 & n9189;
  assign new_n6332 = ~new_n6330 & ~new_n6331;
  assign new_n6333 = new_n6330 & new_n6331;
  assign new_n6334 = ~new_n6332 & ~new_n6333;
  assign new_n6335 = new_n6329 & ~new_n6334;
  assign new_n6336 = ~new_n6329 & new_n6334;
  assign new_n6337 = ~new_n6335 & ~new_n6336;
  assign new_n6338 = new_n6328 & new_n6337;
  assign new_n6339 = ~new_n6328 & ~new_n6337;
  assign new_n6340 = ~new_n6338 & ~new_n6339;
  assign new_n6341 = ~new_n6324 & new_n6340;
  assign new_n6342 = new_n6324 & ~new_n6340;
  assign new_n6343 = ~new_n6341 & ~new_n6342;
  assign new_n6344 = new_n6310 & new_n6343;
  assign new_n6345 = ~new_n6310 & ~new_n6343;
  assign new_n6346 = ~new_n6344 & ~new_n6345;
  assign new_n6347 = ~new_n6109 & ~new_n6346;
  assign new_n6348 = new_n6109 & new_n6346;
  assign new_n6349 = ~new_n6347 & ~new_n6348;
  assign new_n6350 = ~new_n6305 & new_n6349;
  assign new_n6351 = new_n6305 & ~new_n6349;
  assign new_n6352 = ~new_n6350 & ~new_n6351;
  assign new_n6353 = ~new_n6192_1 & new_n6282;
  assign new_n6354 = ~new_n6193 & ~new_n6353;
  assign new_n6355 = ~new_n6352 & new_n6354;
  assign new_n6356 = new_n6352 & ~new_n6354;
  assign new_n6357 = ~new_n6355 & ~new_n6356;
  assign new_n6358_1 = ~new_n6218 & new_n6221;
  assign new_n6359_1 = ~new_n6201 & ~new_n6358_1;
  assign new_n6360 = ~new_n6217 & new_n6359_1;
  assign new_n6361 = new_n6201 & new_n6358_1;
  assign new_n6362 = ~new_n6360 & ~new_n6361;
  assign new_n6363 = n2530 & n6016;
  assign new_n6364 = n2347 & n5331;
  assign new_n6365 = n5798 & n8476;
  assign new_n6366 = ~new_n6364 & ~new_n6365;
  assign new_n6367 = new_n6364 & new_n6365;
  assign new_n6368 = ~new_n6366 & ~new_n6367;
  assign new_n6369 = new_n6363 & ~new_n6368;
  assign new_n6370 = ~new_n6363 & new_n6368;
  assign new_n6371 = ~new_n6369 & ~new_n6370;
  assign new_n6372 = ~new_n6209 & new_n6213;
  assign new_n6373 = ~new_n6210 & ~new_n6372;
  assign new_n6374 = ~new_n6371 & new_n6373;
  assign new_n6375 = new_n6371 & ~new_n6373;
  assign new_n6376 = ~new_n6374 & ~new_n6375;
  assign new_n6377 = n521 & n12648;
  assign new_n6378 = ~new_n6207 & ~new_n6377;
  assign new_n6379 = new_n6207 & new_n6377;
  assign new_n6380 = ~new_n6378 & ~new_n6379;
  assign new_n6381 = n2498 & n7690;
  assign new_n6382 = n2558 & n3616;
  assign new_n6383 = n5579 & n10545;
  assign new_n6384 = ~new_n6382 & ~new_n6383;
  assign new_n6385 = new_n6382 & new_n6383;
  assign new_n6386 = ~new_n6384 & ~new_n6385;
  assign new_n6387 = ~new_n6381 & ~new_n6386;
  assign new_n6388 = new_n6381 & new_n6386;
  assign new_n6389 = ~new_n6387 & ~new_n6388;
  assign new_n6390 = ~new_n6380 & ~new_n6389;
  assign new_n6391 = ~new_n6378 & new_n6389;
  assign new_n6392 = ~new_n6379 & new_n6391;
  assign new_n6393 = ~new_n6390 & ~new_n6392;
  assign new_n6394 = ~new_n6376 & new_n6393;
  assign new_n6395 = new_n6376 & ~new_n6393;
  assign new_n6396 = ~new_n6394 & ~new_n6395;
  assign new_n6397 = ~new_n6362 & new_n6396;
  assign new_n6398 = new_n6362 & ~new_n6396;
  assign new_n6399 = ~new_n6397 & ~new_n6398;
  assign new_n6400 = ~new_n6225 & ~new_n6399;
  assign new_n6401 = new_n6225 & new_n6399;
  assign new_n6402 = ~new_n6400 & ~new_n6401;
  assign new_n6403 = ~new_n6228 & ~new_n6231;
  assign new_n6404 = ~new_n6402 & new_n6403;
  assign new_n6405 = new_n6402 & ~new_n6403;
  assign new_n6406 = ~new_n6404 & ~new_n6405;
  assign new_n6407 = ~new_n6257 & ~new_n6260;
  assign new_n6408 = ~new_n6240 & ~new_n6407;
  assign new_n6409 = ~new_n6256 & new_n6408;
  assign new_n6410 = new_n6240 & new_n6407;
  assign new_n6411 = ~new_n6409 & ~new_n6410;
  assign new_n6412 = n5153 & n7388;
  assign new_n6413 = n7270 & n11892;
  assign new_n6414 = n2507 & n7965;
  assign new_n6415 = ~new_n6413 & ~new_n6414;
  assign new_n6416 = new_n6413 & new_n6414;
  assign new_n6417 = ~new_n6415 & ~new_n6416;
  assign new_n6418 = ~new_n6412 & ~new_n6417;
  assign new_n6419 = new_n6412 & new_n6417;
  assign new_n6420 = ~new_n6418 & ~new_n6419;
  assign new_n6421 = ~new_n6248 & ~new_n6252;
  assign new_n6422 = ~new_n6249 & ~new_n6421;
  assign new_n6423 = new_n6420 & new_n6422;
  assign new_n6424 = ~new_n6420 & ~new_n6422;
  assign new_n6425 = ~new_n6423 & ~new_n6424;
  assign new_n6426 = n806 & n2393;
  assign new_n6427 = new_n6246 & new_n6426;
  assign new_n6428 = ~new_n6246 & ~new_n6426;
  assign new_n6429_1 = ~new_n6427 & ~new_n6428;
  assign new_n6430 = n3986 & n9111;
  assign new_n6431_1 = n5857 & n9763;
  assign new_n6432 = n3342 & n5860;
  assign new_n6433 = ~new_n6431_1 & ~new_n6432;
  assign new_n6434 = new_n6431_1 & new_n6432;
  assign new_n6435 = ~new_n6433 & ~new_n6434;
  assign new_n6436 = ~new_n6430 & ~new_n6435;
  assign new_n6437 = new_n6430 & new_n6435;
  assign new_n6438 = ~new_n6436 & ~new_n6437;
  assign new_n6439 = new_n6429_1 & ~new_n6438;
  assign new_n6440 = ~new_n6429_1 & new_n6438;
  assign new_n6441_1 = ~new_n6439 & ~new_n6440;
  assign new_n6442 = new_n6425 & new_n6441_1;
  assign new_n6443 = ~new_n6425 & ~new_n6441_1;
  assign new_n6444 = ~new_n6442 & ~new_n6443;
  assign new_n6445_1 = new_n6411 & new_n6444;
  assign new_n6446 = ~new_n6411 & ~new_n6444;
  assign new_n6447 = ~new_n6445_1 & ~new_n6446;
  assign new_n6448 = ~new_n6264 & new_n6447;
  assign new_n6449 = new_n6264 & ~new_n6447;
  assign new_n6450 = ~new_n6448 & ~new_n6449;
  assign new_n6451 = ~new_n6267 & ~new_n6270;
  assign new_n6452 = ~new_n6450 & new_n6451;
  assign new_n6453 = new_n6450 & ~new_n6451;
  assign new_n6454 = ~new_n6452 & ~new_n6453;
  assign new_n6455 = ~new_n6406 & ~new_n6454;
  assign new_n6456 = new_n6280 & new_n6455;
  assign new_n6457 = new_n6406 & new_n6454;
  assign new_n6458 = ~new_n6280 & new_n6457;
  assign new_n6459 = ~new_n6280 & ~new_n6455;
  assign new_n6460 = ~new_n6457 & ~new_n6459;
  assign new_n6461 = ~new_n6458 & ~new_n6460;
  assign new_n6462 = ~new_n6456 & ~new_n6461;
  assign new_n6463 = new_n6357 & new_n6462;
  assign new_n6464 = ~new_n6357 & ~new_n6462;
  assign new_n6465 = ~new_n6463 & ~new_n6464;
  assign new_n6466 = ~new_n6304 & new_n6465;
  assign new_n6467 = new_n6304 & ~new_n6465;
  assign n1523 = new_n6466 | new_n6467;
  assign new_n6469 = n2879 & n6687;
  assign new_n6470 = n2564 & n7265;
  assign new_n6471 = new_n6469 & new_n6470;
  assign new_n6472 = n4189 & n7265;
  assign new_n6473 = n2564 & n2879;
  assign new_n6474 = n6687 & n10223;
  assign new_n6475 = ~new_n6473 & ~new_n6474;
  assign new_n6476 = new_n6473 & new_n6474;
  assign new_n6477 = ~new_n6475 & ~new_n6476;
  assign new_n6478 = new_n6472 & ~new_n6477;
  assign new_n6479 = ~new_n6472 & new_n6477;
  assign new_n6480 = ~new_n6478 & ~new_n6479;
  assign new_n6481 = new_n6471 & ~new_n6480;
  assign new_n6482 = n4634 & n6687;
  assign new_n6483 = new_n6472 & ~new_n6475;
  assign new_n6484 = ~new_n6476 & ~new_n6483;
  assign new_n6485 = new_n6482 & ~new_n6484;
  assign new_n6486 = ~new_n6482 & new_n6484;
  assign new_n6487 = ~new_n6485 & ~new_n6486;
  assign new_n6488 = n2879 & n4189;
  assign new_n6489 = n2564 & n10223;
  assign new_n6490 = n6770 & n7265;
  assign new_n6491 = ~new_n6489 & ~new_n6490;
  assign new_n6492 = new_n6489 & new_n6490;
  assign new_n6493 = ~new_n6491 & ~new_n6492;
  assign new_n6494 = new_n6488 & ~new_n6493;
  assign new_n6495 = ~new_n6488 & new_n6493;
  assign new_n6496 = ~new_n6494 & ~new_n6495;
  assign new_n6497 = ~new_n6487 & ~new_n6496;
  assign new_n6498 = new_n6487 & new_n6496;
  assign new_n6499 = ~new_n6497 & ~new_n6498;
  assign new_n6500 = new_n6481 & ~new_n6499;
  assign new_n6501 = ~new_n6481 & new_n6499;
  assign new_n6502 = ~new_n6500 & ~new_n6501;
  assign new_n6503 = n2024 & n8336;
  assign new_n6504 = n7946 & n10928;
  assign new_n6505 = new_n6503 & new_n6504;
  assign new_n6506 = n6986 & n7946;
  assign new_n6507 = n2024 & n10928;
  assign new_n6508 = n8336 & n9189;
  assign new_n6509 = ~new_n6507 & ~new_n6508;
  assign new_n6510 = new_n6507 & new_n6508;
  assign new_n6511 = ~new_n6509 & ~new_n6510;
  assign new_n6512 = new_n6506 & ~new_n6511;
  assign new_n6513 = ~new_n6506 & new_n6511;
  assign new_n6514 = ~new_n6512 & ~new_n6513;
  assign new_n6515 = new_n6505 & ~new_n6514;
  assign new_n6516 = n2522 & n8336;
  assign new_n6517 = new_n6506 & ~new_n6509;
  assign new_n6518 = ~new_n6510 & ~new_n6517;
  assign new_n6519 = new_n6516 & ~new_n6518;
  assign new_n6520 = ~new_n6516 & new_n6518;
  assign new_n6521 = ~new_n6519 & ~new_n6520;
  assign new_n6522 = n2226 & n7946;
  assign new_n6523 = n9189 & n10928;
  assign new_n6524 = n2024 & n6986;
  assign new_n6525 = ~new_n6523 & ~new_n6524;
  assign new_n6526 = new_n6523 & new_n6524;
  assign new_n6527 = ~new_n6525 & ~new_n6526;
  assign new_n6528 = new_n6522 & ~new_n6527;
  assign new_n6529 = ~new_n6522 & new_n6527;
  assign new_n6530 = ~new_n6528 & ~new_n6529;
  assign new_n6531 = ~new_n6521 & ~new_n6530;
  assign new_n6532 = new_n6521 & new_n6530;
  assign new_n6533 = ~new_n6531 & ~new_n6532;
  assign new_n6534 = new_n6515 & ~new_n6533;
  assign new_n6535 = ~new_n6515 & new_n6533;
  assign new_n6536 = ~new_n6534 & ~new_n6535;
  assign new_n6537 = n2498 & n12069;
  assign new_n6538 = n2558 & n12391;
  assign new_n6539 = new_n6537 & new_n6538;
  assign new_n6540 = n2558 & n7891;
  assign new_n6541 = n2498 & n12391;
  assign new_n6542 = n5579 & n12069;
  assign new_n6543 = ~new_n6541 & ~new_n6542;
  assign new_n6544 = new_n6541 & new_n6542;
  assign new_n6545 = ~new_n6543 & ~new_n6544;
  assign new_n6546 = new_n6540 & ~new_n6545;
  assign new_n6547 = ~new_n6540 & new_n6545;
  assign new_n6548 = ~new_n6546 & ~new_n6547;
  assign new_n6549 = new_n6539 & ~new_n6548;
  assign new_n6550 = n521 & n12069;
  assign new_n6551 = new_n6540 & ~new_n6543;
  assign new_n6552 = ~new_n6544 & ~new_n6551;
  assign new_n6553 = ~new_n6550 & new_n6552;
  assign new_n6554 = new_n6550 & ~new_n6552;
  assign new_n6555 = ~new_n6553 & ~new_n6554;
  assign new_n6556 = n2558 & n7160;
  assign new_n6557 = n5579 & n12391;
  assign new_n6558 = n2498 & n7891;
  assign new_n6559 = ~new_n6557 & ~new_n6558;
  assign new_n6560 = new_n6557 & new_n6558;
  assign new_n6561 = ~new_n6559 & ~new_n6560;
  assign new_n6562 = new_n6556 & ~new_n6561;
  assign new_n6563 = ~new_n6556 & new_n6561;
  assign new_n6564 = ~new_n6562 & ~new_n6563;
  assign new_n6565 = ~new_n6555 & new_n6564;
  assign new_n6566 = new_n6555 & ~new_n6564;
  assign new_n6567 = ~new_n6565 & ~new_n6566;
  assign new_n6568 = ~new_n6549 & ~new_n6567;
  assign new_n6569 = new_n6549 & new_n6567;
  assign new_n6570 = ~new_n6568 & ~new_n6569;
  assign new_n6571 = n9111 & n11222;
  assign new_n6572 = n9763 & n11153;
  assign new_n6573 = new_n6571 & new_n6572;
  assign new_n6574 = n5314 & n9763;
  assign new_n6575 = n9111 & n11153;
  assign new_n6576 = n3342 & n11222;
  assign new_n6577 = ~new_n6575 & ~new_n6576;
  assign new_n6578_1 = new_n6575 & new_n6576;
  assign new_n6579 = ~new_n6577 & ~new_n6578_1;
  assign new_n6580 = new_n6574 & ~new_n6579;
  assign new_n6581 = ~new_n6574 & new_n6579;
  assign new_n6582 = ~new_n6580 & ~new_n6581;
  assign new_n6583 = new_n6573 & ~new_n6582;
  assign new_n6584 = n806 & n11222;
  assign new_n6585 = new_n6574 & ~new_n6577;
  assign new_n6586 = ~new_n6578_1 & ~new_n6585;
  assign new_n6587 = new_n6584 & ~new_n6586;
  assign new_n6588 = ~new_n6584 & new_n6586;
  assign new_n6589 = ~new_n6587 & ~new_n6588;
  assign new_n6590 = n996 & n9763;
  assign new_n6591 = n3342 & n11153;
  assign new_n6592 = n5314 & n9111;
  assign new_n6593 = ~new_n6591 & ~new_n6592;
  assign new_n6594 = new_n6591 & new_n6592;
  assign new_n6595 = ~new_n6593 & ~new_n6594;
  assign new_n6596 = new_n6590 & ~new_n6595;
  assign new_n6597 = ~new_n6590 & new_n6595;
  assign new_n6598 = ~new_n6596 & ~new_n6597;
  assign new_n6599 = ~new_n6589 & ~new_n6598;
  assign new_n6600 = new_n6589 & new_n6598;
  assign new_n6601 = ~new_n6599 & ~new_n6600;
  assign new_n6602 = new_n6583 & ~new_n6601;
  assign new_n6603 = ~new_n6583 & new_n6601;
  assign new_n6604_1 = ~new_n6602 & ~new_n6603;
  assign new_n6605 = new_n6570 & new_n6604_1;
  assign new_n6606 = ~new_n6570 & ~new_n6604_1;
  assign new_n6607 = ~new_n6605 & ~new_n6606;
  assign new_n6608 = ~new_n6573 & new_n6582;
  assign new_n6609 = ~new_n6583 & ~new_n6608;
  assign new_n6610 = ~new_n6537 & ~new_n6538;
  assign new_n6611_1 = ~new_n6539 & ~new_n6610;
  assign new_n6612 = new_n4919 & new_n6611_1;
  assign new_n6613 = ~new_n4919 & ~new_n6611_1;
  assign new_n6614 = ~new_n6571 & ~new_n6572;
  assign new_n6615 = ~new_n6573 & ~new_n6614;
  assign new_n6616 = ~new_n6613 & new_n6615;
  assign new_n6617 = ~new_n6612 & ~new_n6616;
  assign new_n6618 = new_n6609 & ~new_n6617;
  assign new_n6619 = ~new_n6539 & new_n6548;
  assign new_n6620 = ~new_n6549 & ~new_n6619;
  assign new_n6621 = ~new_n6609 & new_n6617;
  assign new_n6622 = new_n6620 & ~new_n6621;
  assign new_n6623 = ~new_n6618 & ~new_n6622;
  assign new_n6624 = new_n6607 & new_n6623;
  assign new_n6625 = ~new_n6607 & ~new_n6623;
  assign new_n6626 = ~new_n6624 & ~new_n6625;
  assign new_n6627 = new_n6536 & ~new_n6626;
  assign new_n6628 = ~new_n6536 & new_n6626;
  assign new_n6629 = ~new_n6627 & ~new_n6628;
  assign new_n6630 = ~new_n6505 & new_n6514;
  assign new_n6631 = ~new_n6515 & ~new_n6630;
  assign new_n6632 = ~new_n6618 & ~new_n6621;
  assign new_n6633 = ~new_n6620 & ~new_n6632;
  assign new_n6634 = new_n6620 & new_n6632;
  assign new_n6635 = ~new_n6633 & ~new_n6634;
  assign new_n6636 = ~new_n6631 & ~new_n6635;
  assign new_n6637 = new_n6631 & new_n6635;
  assign new_n6638 = ~new_n6503 & ~new_n6504;
  assign new_n6639 = ~new_n6505 & ~new_n6638;
  assign new_n6640 = ~new_n6612 & ~new_n6613;
  assign new_n6641 = new_n6615 & ~new_n6640;
  assign new_n6642 = ~new_n6615 & new_n6640;
  assign new_n6643 = ~new_n6641 & ~new_n6642;
  assign new_n6644 = new_n6639 & ~new_n6643;
  assign new_n6645_1 = ~new_n6639 & new_n6643;
  assign new_n6646 = new_n4922 & ~new_n6645_1;
  assign new_n6647 = ~new_n6644 & ~new_n6646;
  assign new_n6648 = ~new_n6637 & new_n6647;
  assign new_n6649 = ~new_n6636 & ~new_n6648;
  assign new_n6650 = ~new_n6629 & ~new_n6649;
  assign new_n6651 = new_n6629 & new_n6649;
  assign new_n6652 = ~new_n6650 & ~new_n6651;
  assign new_n6653 = new_n6502 & new_n6652;
  assign new_n6654 = ~new_n6502 & ~new_n6652;
  assign new_n6655 = ~new_n6471 & new_n6480;
  assign new_n6656 = ~new_n6481 & ~new_n6655;
  assign new_n6657 = ~new_n6636 & ~new_n6637;
  assign new_n6658 = ~new_n6647 & ~new_n6657;
  assign new_n6659 = new_n6647 & new_n6657;
  assign new_n6660 = ~new_n6658 & ~new_n6659;
  assign new_n6661 = new_n6656 & ~new_n6660;
  assign new_n6662 = ~new_n6656 & new_n6660;
  assign new_n6663 = ~new_n6469 & ~new_n6470;
  assign new_n6664 = ~new_n6471 & ~new_n6663;
  assign new_n6665 = new_n4925 & new_n6664;
  assign new_n6666 = ~new_n4925 & ~new_n6664;
  assign new_n6667 = ~new_n6644 & ~new_n6645_1;
  assign new_n6668 = ~new_n4922 & ~new_n6667;
  assign new_n6669 = new_n4922 & new_n6667;
  assign new_n6670 = ~new_n6668 & ~new_n6669;
  assign new_n6671 = ~new_n6666 & new_n6670;
  assign new_n6672 = ~new_n6665 & ~new_n6671;
  assign new_n6673 = ~new_n6662 & ~new_n6672;
  assign new_n6674 = ~new_n6661 & ~new_n6673;
  assign new_n6675 = ~new_n6654 & ~new_n6674;
  assign new_n6676 = ~new_n6653 & ~new_n6675;
  assign new_n6677 = n6687 & n9195;
  assign new_n6678 = n2564 & n4634;
  assign new_n6679 = n2879 & n6770;
  assign new_n6680 = n7265 & n9920;
  assign new_n6681 = n4189 & n10223;
  assign new_n6682 = ~new_n6680 & ~new_n6681;
  assign new_n6683 = n9920 & n10223;
  assign new_n6684 = new_n6472 & new_n6683;
  assign new_n6685 = ~new_n6682 & ~new_n6684;
  assign new_n6686 = ~new_n6679 & new_n6685;
  assign new_n6687_1 = new_n6679 & ~new_n6685;
  assign new_n6688 = ~new_n6686 & ~new_n6687_1;
  assign new_n6689_1 = new_n6678 & ~new_n6688;
  assign new_n6690 = ~new_n6678 & new_n6688;
  assign new_n6691 = ~new_n6689_1 & ~new_n6690;
  assign new_n6692 = new_n6488 & ~new_n6491;
  assign new_n6693 = ~new_n6492 & ~new_n6692;
  assign new_n6694 = ~new_n6691 & ~new_n6693;
  assign new_n6695 = new_n6691 & new_n6693;
  assign new_n6696 = ~new_n6694 & ~new_n6695;
  assign new_n6697 = new_n6677 & ~new_n6696;
  assign new_n6698 = ~new_n6677 & new_n6696;
  assign new_n6699 = ~new_n6697 & ~new_n6698;
  assign new_n6700 = ~new_n6486 & ~new_n6496;
  assign new_n6701 = ~new_n6485 & ~new_n6700;
  assign new_n6702 = ~new_n6699 & ~new_n6701;
  assign new_n6703_1 = new_n6699 & new_n6701;
  assign new_n6704 = ~new_n6702 & ~new_n6703_1;
  assign new_n6705 = new_n6500 & ~new_n6704;
  assign new_n6706 = ~new_n6500 & new_n6704;
  assign new_n6707 = ~new_n6705 & ~new_n6706;
  assign new_n6708 = n6016 & n12069;
  assign new_n6709 = n2558 & n4828;
  assign new_n6710 = n5579 & n7891;
  assign new_n6711 = n2498 & n7160;
  assign new_n6712 = ~new_n6710 & ~new_n6711;
  assign new_n6713 = new_n6710 & new_n6711;
  assign new_n6714 = ~new_n6712 & ~new_n6713;
  assign new_n6715 = ~new_n6709 & ~new_n6714;
  assign new_n6716 = new_n6709 & new_n6714;
  assign new_n6717 = ~new_n6715 & ~new_n6716;
  assign new_n6718 = n521 & n12391;
  assign new_n6719 = new_n6556 & ~new_n6559;
  assign new_n6720 = ~new_n6560 & ~new_n6719;
  assign new_n6721 = ~new_n6718 & new_n6720;
  assign new_n6722 = new_n6718 & ~new_n6720;
  assign new_n6723 = ~new_n6721 & ~new_n6722;
  assign new_n6724 = ~new_n6717 & ~new_n6723;
  assign new_n6725 = new_n6717 & new_n6723;
  assign new_n6726 = ~new_n6724 & ~new_n6725;
  assign new_n6727 = new_n6708 & new_n6726;
  assign new_n6728 = ~new_n6708 & ~new_n6726;
  assign new_n6729 = ~new_n6727 & ~new_n6728;
  assign new_n6730 = ~new_n6553 & ~new_n6564;
  assign new_n6731 = ~new_n6554 & ~new_n6730;
  assign new_n6732 = ~new_n6729 & ~new_n6731;
  assign new_n6733 = new_n6729 & new_n6731;
  assign new_n6734 = ~new_n6732 & ~new_n6733;
  assign new_n6735 = new_n6569 & ~new_n6734;
  assign new_n6736 = ~new_n6569 & new_n6734;
  assign new_n6737 = ~new_n6735 & ~new_n6736;
  assign new_n6738 = n7270 & n11222;
  assign new_n6739 = n806 & n11153;
  assign new_n6740 = new_n6590 & ~new_n6593;
  assign new_n6741 = ~new_n6594 & ~new_n6740;
  assign new_n6742_1 = ~new_n6739 & new_n6741;
  assign new_n6743 = new_n6739 & ~new_n6741;
  assign new_n6744 = ~new_n6742_1 & ~new_n6743;
  assign new_n6745 = n5767 & n9763;
  assign new_n6746 = n3342 & n5314;
  assign new_n6747 = n996 & n9111;
  assign new_n6748 = ~new_n6746 & ~new_n6747;
  assign new_n6749 = new_n6746 & new_n6747;
  assign new_n6750 = ~new_n6748 & ~new_n6749;
  assign new_n6751 = new_n6745 & ~new_n6750;
  assign new_n6752 = ~new_n6745 & new_n6750;
  assign new_n6753 = ~new_n6751 & ~new_n6752;
  assign new_n6754 = ~new_n6744 & new_n6753;
  assign new_n6755 = new_n6744 & ~new_n6753;
  assign new_n6756 = ~new_n6754 & ~new_n6755;
  assign new_n6757 = new_n6738 & new_n6756;
  assign new_n6758 = ~new_n6738 & ~new_n6756;
  assign new_n6759 = ~new_n6757 & ~new_n6758;
  assign new_n6760 = ~new_n6587 & new_n6598;
  assign new_n6761 = ~new_n6588 & ~new_n6760;
  assign new_n6762 = ~new_n6759 & new_n6761;
  assign new_n6763 = new_n6759 & ~new_n6761;
  assign new_n6764 = ~new_n6762 & ~new_n6763;
  assign new_n6765 = new_n6602 & ~new_n6764;
  assign new_n6766 = ~new_n6602 & new_n6764;
  assign new_n6767 = ~new_n6765 & ~new_n6766;
  assign new_n6768 = new_n6737 & new_n6767;
  assign new_n6769 = ~new_n6737 & ~new_n6767;
  assign new_n6770_1 = ~new_n6768 & ~new_n6769;
  assign new_n6771 = ~new_n6606 & ~new_n6623;
  assign new_n6772 = ~new_n6605 & ~new_n6771;
  assign new_n6773 = new_n6770_1 & new_n6772;
  assign new_n6774 = ~new_n6770_1 & ~new_n6772;
  assign new_n6775 = ~new_n6773 & ~new_n6774;
  assign new_n6776_1 = n8336 & n12145;
  assign new_n6777 = n2522 & n10928;
  assign new_n6778 = new_n6522 & ~new_n6525;
  assign new_n6779 = ~new_n6526 & ~new_n6778;
  assign new_n6780 = new_n6777 & ~new_n6779;
  assign new_n6781 = ~new_n6777 & new_n6779;
  assign new_n6782 = ~new_n6780 & ~new_n6781;
  assign new_n6783 = n2024 & n2226;
  assign new_n6784 = n6986 & n9189;
  assign new_n6785 = n1094 & n7946;
  assign new_n6786 = ~new_n6784 & ~new_n6785;
  assign new_n6787 = new_n6784 & new_n6785;
  assign new_n6788 = ~new_n6786 & ~new_n6787;
  assign new_n6789 = new_n6783 & ~new_n6788;
  assign new_n6790 = ~new_n6783 & new_n6788;
  assign new_n6791 = ~new_n6789 & ~new_n6790;
  assign new_n6792 = ~new_n6782 & ~new_n6791;
  assign new_n6793 = new_n6782 & new_n6791;
  assign new_n6794 = ~new_n6792 & ~new_n6793;
  assign new_n6795 = new_n6776_1 & ~new_n6794;
  assign new_n6796 = ~new_n6776_1 & new_n6794;
  assign new_n6797_1 = ~new_n6795 & ~new_n6796;
  assign new_n6798 = ~new_n6519 & new_n6530;
  assign new_n6799 = ~new_n6520 & ~new_n6798;
  assign new_n6800 = ~new_n6797_1 & new_n6799;
  assign new_n6801 = new_n6797_1 & ~new_n6799;
  assign new_n6802 = ~new_n6800 & ~new_n6801;
  assign new_n6803 = new_n6534 & ~new_n6802;
  assign new_n6804 = ~new_n6534 & new_n6802;
  assign new_n6805 = ~new_n6803 & ~new_n6804;
  assign new_n6806_1 = ~new_n6627 & ~new_n6649;
  assign new_n6807 = ~new_n6628 & ~new_n6806_1;
  assign new_n6808 = ~new_n6805 & ~new_n6807;
  assign new_n6809_1 = new_n6805 & new_n6807;
  assign new_n6810 = ~new_n6808 & ~new_n6809_1;
  assign new_n6811 = new_n6775 & ~new_n6810;
  assign new_n6812 = ~new_n6775 & new_n6810;
  assign new_n6813 = ~new_n6811 & ~new_n6812;
  assign new_n6814 = ~new_n6707 & ~new_n6813;
  assign new_n6815 = new_n6707 & new_n6813;
  assign new_n6816 = ~new_n6814 & ~new_n6815;
  assign new_n6817 = new_n6676 & new_n6816;
  assign new_n6818 = ~new_n6676 & ~new_n6816;
  assign n1658 = new_n6817 | new_n6818;
  assign new_n6820 = n2879 & n7862;
  assign new_n6821 = n1333 & n7265;
  assign new_n6822_1 = new_n6820 & new_n6821;
  assign new_n6823 = n3172 & n7265;
  assign new_n6824 = n1333 & n2879;
  assign new_n6825 = n7862 & n10223;
  assign new_n6826_1 = ~new_n6824 & ~new_n6825;
  assign new_n6827 = new_n6824 & new_n6825;
  assign new_n6828 = ~new_n6826_1 & ~new_n6827;
  assign new_n6829 = new_n6823 & ~new_n6828;
  assign new_n6830 = ~new_n6823 & new_n6828;
  assign new_n6831 = ~new_n6829 & ~new_n6830;
  assign new_n6832 = new_n6822_1 & ~new_n6831;
  assign new_n6833 = n4634 & n7862;
  assign new_n6834 = new_n6823 & ~new_n6826_1;
  assign new_n6835 = ~new_n6827 & ~new_n6834;
  assign new_n6836 = ~new_n6833 & new_n6835;
  assign new_n6837 = new_n6833 & ~new_n6835;
  assign new_n6838 = ~new_n6836 & ~new_n6837;
  assign new_n6839 = n7265 & n11757;
  assign new_n6840 = n1333 & n10223;
  assign new_n6841 = n2879 & n3172;
  assign new_n6842 = ~new_n6840 & ~new_n6841;
  assign new_n6843 = new_n6840 & new_n6841;
  assign new_n6844 = ~new_n6842 & ~new_n6843;
  assign new_n6845 = new_n6839 & ~new_n6844;
  assign new_n6846 = ~new_n6839 & new_n6844;
  assign new_n6847 = ~new_n6845 & ~new_n6846;
  assign new_n6848 = ~new_n6838 & new_n6847;
  assign new_n6849 = new_n6838 & ~new_n6847;
  assign new_n6850 = ~new_n6848 & ~new_n6849;
  assign new_n6851 = new_n6832 & new_n6850;
  assign new_n6852 = ~new_n6832 & ~new_n6850;
  assign new_n6853 = ~new_n6851 & ~new_n6852;
  assign new_n6854 = n2024 & n6877;
  assign new_n6855 = n7946 & n9400;
  assign new_n6856 = new_n6854 & new_n6855;
  assign new_n6857 = n2464 & n7946;
  assign new_n6858 = n2024 & n9400;
  assign new_n6859 = n6877 & n9189;
  assign new_n6860_1 = ~new_n6858 & ~new_n6859;
  assign new_n6861 = new_n6858 & new_n6859;
  assign new_n6862 = ~new_n6860_1 & ~new_n6861;
  assign new_n6863 = new_n6857 & ~new_n6862;
  assign new_n6864 = ~new_n6857 & new_n6862;
  assign new_n6865 = ~new_n6863 & ~new_n6864;
  assign new_n6866 = new_n6856 & ~new_n6865;
  assign new_n6867 = n2522 & n6877;
  assign new_n6868 = n2024 & n2464;
  assign new_n6869 = n9189 & n9400;
  assign new_n6870 = n7946 & n11311;
  assign new_n6871 = ~new_n6869 & ~new_n6870;
  assign new_n6872 = new_n6869 & new_n6870;
  assign new_n6873 = ~new_n6871 & ~new_n6872;
  assign new_n6874 = new_n6868 & ~new_n6873;
  assign new_n6875 = ~new_n6868 & new_n6873;
  assign new_n6876 = ~new_n6874 & ~new_n6875;
  assign new_n6877_1 = new_n6867 & ~new_n6876;
  assign new_n6878 = ~new_n6867 & new_n6876;
  assign new_n6879 = ~new_n6877_1 & ~new_n6878;
  assign new_n6880 = new_n6857 & ~new_n6860_1;
  assign new_n6881 = ~new_n6861 & ~new_n6880;
  assign new_n6882 = ~new_n6879 & ~new_n6881;
  assign new_n6883 = new_n6879 & new_n6881;
  assign new_n6884 = ~new_n6882 & ~new_n6883;
  assign new_n6885 = ~new_n6866 & new_n6884;
  assign new_n6886 = new_n6866 & ~new_n6884;
  assign new_n6887 = ~new_n6885 & ~new_n6886;
  assign new_n6888 = ~new_n6856 & new_n6865;
  assign new_n6889 = ~new_n6866 & ~new_n6888;
  assign new_n6890 = n6877 & n7946;
  assign new_n6891 = n2558 & n4805;
  assign new_n6892 = n7236 & n9763;
  assign new_n6893 = new_n6891 & new_n6892;
  assign new_n6894 = ~new_n6891 & ~new_n6892;
  assign new_n6895 = ~new_n6893 & ~new_n6894;
  assign new_n6896 = new_n6890 & new_n6895;
  assign new_n6897 = ~new_n6854 & ~new_n6855;
  assign new_n6898 = ~new_n6856 & ~new_n6897;
  assign new_n6899 = new_n6896 & new_n6898;
  assign new_n6900 = ~new_n6896 & ~new_n6898;
  assign new_n6901 = n2498 & n4805;
  assign new_n6902 = n2558 & n11478;
  assign new_n6903 = ~new_n6901 & ~new_n6902;
  assign new_n6904 = new_n6901 & new_n6902;
  assign new_n6905 = ~new_n6903 & ~new_n6904;
  assign new_n6906 = n7236 & n9111;
  assign new_n6907 = n3992 & n9763;
  assign new_n6908 = ~new_n6906 & ~new_n6907;
  assign new_n6909 = new_n6906 & new_n6907;
  assign new_n6910 = ~new_n6908 & ~new_n6909;
  assign new_n6911 = new_n6893 & new_n6910;
  assign new_n6912 = ~new_n6893 & ~new_n6910;
  assign new_n6913 = ~new_n6911 & ~new_n6912;
  assign new_n6914 = new_n6905 & ~new_n6913;
  assign new_n6915 = ~new_n6905 & new_n6913;
  assign new_n6916 = ~new_n6914 & ~new_n6915;
  assign new_n6917 = ~new_n6900 & ~new_n6916;
  assign new_n6918 = ~new_n6899 & ~new_n6917;
  assign new_n6919 = new_n6889 & ~new_n6918;
  assign new_n6920 = ~new_n6889 & new_n6918;
  assign new_n6921 = ~new_n6905 & ~new_n6911;
  assign new_n6922 = ~new_n6912 & ~new_n6921;
  assign new_n6923 = n2498 & n11478;
  assign new_n6924 = ~new_n6891 & new_n6923;
  assign new_n6925 = n2558 & n5283;
  assign new_n6926 = n4805 & n5579;
  assign new_n6927 = ~new_n6925 & ~new_n6926;
  assign new_n6928 = n5283 & n5579;
  assign new_n6929 = new_n6891 & new_n6928;
  assign new_n6930 = ~new_n6927 & ~new_n6929;
  assign new_n6931 = ~new_n6924 & ~new_n6930;
  assign new_n6932 = new_n6924 & ~new_n6927;
  assign new_n6933 = ~new_n6931 & ~new_n6932;
  assign new_n6934 = ~new_n6922 & ~new_n6933;
  assign new_n6935 = n8384 & n9763;
  assign new_n6936 = n3342 & n7236;
  assign new_n6937 = ~new_n6935 & ~new_n6936;
  assign new_n6938 = n3342 & n8384;
  assign new_n6939 = new_n6892 & new_n6938;
  assign new_n6940 = ~new_n6937 & ~new_n6939;
  assign new_n6941 = n3992 & n9111;
  assign new_n6942 = ~new_n6892 & new_n6941;
  assign new_n6943 = ~new_n6940 & ~new_n6942;
  assign new_n6944 = ~new_n6937 & new_n6941;
  assign new_n6945 = ~new_n6892 & new_n6944;
  assign new_n6946 = ~new_n6943 & ~new_n6945;
  assign new_n6947 = new_n6934 & ~new_n6946;
  assign new_n6948 = new_n6922 & new_n6933;
  assign new_n6949 = ~new_n6946 & ~new_n6948;
  assign new_n6950 = ~new_n6934 & ~new_n6949;
  assign new_n6951 = ~new_n6947 & ~new_n6950;
  assign new_n6952 = new_n6946 & new_n6948;
  assign new_n6953 = ~new_n6951 & ~new_n6952;
  assign new_n6954 = ~new_n6920 & ~new_n6953;
  assign new_n6955 = ~new_n6919 & ~new_n6954;
  assign new_n6956 = new_n6887 & ~new_n6955;
  assign new_n6957 = ~new_n6887 & new_n6955;
  assign new_n6958 = ~new_n6956 & ~new_n6957;
  assign new_n6959 = new_n6904 & ~new_n6930;
  assign new_n6960 = n521 & n4805;
  assign new_n6961 = ~new_n6923 & ~new_n6929;
  assign new_n6962 = ~new_n6927 & ~new_n6961;
  assign new_n6963 = new_n6960 & new_n6962;
  assign new_n6964 = ~new_n6960 & ~new_n6962;
  assign new_n6965 = ~new_n6963 & ~new_n6964;
  assign new_n6966 = n137 & n2558;
  assign new_n6967 = n5579 & n11478;
  assign new_n6968 = n2498 & n5283;
  assign new_n6969 = ~new_n6967 & ~new_n6968;
  assign new_n6970 = new_n6967 & new_n6968;
  assign new_n6971 = ~new_n6969 & ~new_n6970;
  assign new_n6972 = new_n6966 & ~new_n6971;
  assign new_n6973 = ~new_n6966 & new_n6971;
  assign new_n6974 = ~new_n6972 & ~new_n6973;
  assign new_n6975 = ~new_n6965 & ~new_n6974;
  assign new_n6976 = new_n6965 & new_n6974;
  assign new_n6977 = ~new_n6975 & ~new_n6976;
  assign new_n6978 = new_n6959 & ~new_n6977;
  assign new_n6979 = ~new_n6959 & new_n6977;
  assign new_n6980 = ~new_n6978 & ~new_n6979;
  assign new_n6981 = new_n6909 & ~new_n6940;
  assign new_n6982 = n806 & n7236;
  assign new_n6983 = ~new_n6939 & ~new_n6944;
  assign new_n6984 = new_n6982 & ~new_n6983;
  assign new_n6985 = ~new_n6982 & new_n6983;
  assign new_n6986_1 = ~new_n6984 & ~new_n6985;
  assign new_n6987 = n6358 & n9763;
  assign new_n6988 = n3342 & n3992;
  assign new_n6989 = n8384 & n9111;
  assign new_n6990 = ~new_n6988 & ~new_n6989;
  assign new_n6991 = new_n6988 & new_n6989;
  assign new_n6992 = ~new_n6990 & ~new_n6991;
  assign new_n6993 = new_n6987 & ~new_n6992;
  assign new_n6994 = ~new_n6987 & new_n6992;
  assign new_n6995 = ~new_n6993 & ~new_n6994;
  assign new_n6996 = ~new_n6986_1 & ~new_n6995;
  assign new_n6997 = new_n6986_1 & new_n6995;
  assign new_n6998 = ~new_n6996 & ~new_n6997;
  assign new_n6999 = new_n6981 & ~new_n6998;
  assign new_n7000 = ~new_n6981 & new_n6998;
  assign new_n7001 = ~new_n6999 & ~new_n7000;
  assign new_n7002 = ~new_n6980 & ~new_n7001;
  assign new_n7003 = ~new_n6950 & new_n7002;
  assign new_n7004 = new_n6980 & new_n7001;
  assign new_n7005 = ~new_n6950 & ~new_n7004;
  assign new_n7006 = ~new_n7002 & ~new_n7005;
  assign new_n7007 = ~new_n7003 & ~new_n7006;
  assign new_n7008 = new_n6950 & new_n7004;
  assign new_n7009 = ~new_n7007 & ~new_n7008;
  assign new_n7010 = new_n6958 & new_n7009;
  assign new_n7011 = ~new_n6958 & ~new_n7009;
  assign new_n7012 = ~new_n7010 & ~new_n7011;
  assign new_n7013 = new_n6853 & ~new_n7012;
  assign new_n7014 = ~new_n6853 & new_n7012;
  assign new_n7015 = ~new_n7013 & ~new_n7014;
  assign new_n7016 = ~new_n6822_1 & new_n6831;
  assign new_n7017 = ~new_n6832 & ~new_n7016;
  assign new_n7018 = ~new_n6919 & ~new_n6920;
  assign new_n7019 = new_n6953 & ~new_n7018;
  assign new_n7020 = ~new_n6953 & new_n7018;
  assign new_n7021 = ~new_n7019 & ~new_n7020;
  assign new_n7022 = ~new_n7017 & ~new_n7021;
  assign new_n7023 = new_n7017 & new_n7021;
  assign new_n7024 = n7265 & n7862;
  assign new_n7025 = ~new_n6890 & ~new_n6895;
  assign new_n7026 = ~new_n6896 & ~new_n7025;
  assign new_n7027 = new_n7024 & new_n7026;
  assign new_n7028 = ~new_n6820 & ~new_n6821;
  assign new_n7029 = ~new_n6822_1 & ~new_n7028;
  assign new_n7030 = new_n7027 & new_n7029;
  assign new_n7031 = ~new_n7027 & ~new_n7029;
  assign new_n7032 = ~new_n6899 & ~new_n6900;
  assign new_n7033 = new_n6916 & ~new_n7032;
  assign new_n7034 = ~new_n6916 & new_n7032;
  assign new_n7035 = ~new_n7033 & ~new_n7034;
  assign new_n7036 = ~new_n7031 & new_n7035;
  assign new_n7037 = ~new_n7030 & ~new_n7036;
  assign new_n7038 = ~new_n7023 & new_n7037;
  assign new_n7039 = ~new_n7022 & ~new_n7038;
  assign new_n7040 = ~new_n7015 & new_n7039;
  assign new_n7041 = new_n7015 & ~new_n7039;
  assign n1847 = new_n7040 | new_n7041;
  assign new_n7043 = n1798 & n5305;
  assign new_n7044 = n6703 & n8759;
  assign new_n7045 = n5331 & n5645;
  assign new_n7046 = n7965 & n11876;
  assign new_n7047 = new_n7045 & new_n7046;
  assign new_n7048 = ~new_n7045 & ~new_n7046;
  assign new_n7049 = ~new_n7047 & ~new_n7048;
  assign new_n7050 = new_n7044 & new_n7049;
  assign new_n7051 = ~new_n7044 & ~new_n7049;
  assign new_n7052 = ~new_n7050 & ~new_n7051;
  assign new_n7053 = new_n7043 & new_n7052;
  assign new_n7054 = n3932 & n5305;
  assign new_n7055 = n1798 & n5964;
  assign new_n7056 = ~new_n7054 & ~new_n7055;
  assign new_n7057 = new_n7054 & new_n7055;
  assign new_n7058 = ~new_n7056 & ~new_n7057;
  assign new_n7059 = new_n7053 & new_n7058;
  assign new_n7060 = ~new_n7053 & ~new_n7058;
  assign new_n7061 = ~new_n7059 & ~new_n7060;
  assign new_n7062 = n8759 & n9640;
  assign new_n7063 = n6703 & n6776;
  assign new_n7064 = ~new_n7062 & ~new_n7063;
  assign new_n7065 = new_n7062 & new_n7063;
  assign new_n7066 = ~new_n7064 & ~new_n7065;
  assign new_n7067 = new_n7050 & new_n7066;
  assign new_n7068 = ~new_n7050 & ~new_n7066;
  assign new_n7069 = ~new_n7067 & ~new_n7068;
  assign new_n7070 = n7965 & n10898;
  assign new_n7071 = n7388 & n11876;
  assign new_n7072 = ~new_n7070 & ~new_n7071;
  assign new_n7073 = new_n7070 & new_n7071;
  assign new_n7074 = ~new_n7072 & ~new_n7073;
  assign new_n7075 = new_n7047 & new_n7074;
  assign new_n7076 = ~new_n7047 & ~new_n7074;
  assign new_n7077 = ~new_n7075 & ~new_n7076;
  assign new_n7078 = n1067 & n5331;
  assign new_n7079 = n5645 & n8476;
  assign new_n7080 = ~new_n7078 & ~new_n7079;
  assign new_n7081 = new_n7078 & new_n7079;
  assign new_n7082 = ~new_n7080 & ~new_n7081;
  assign new_n7083 = ~new_n7077 & new_n7082;
  assign new_n7084 = new_n7077 & ~new_n7082;
  assign new_n7085 = ~new_n7083 & ~new_n7084;
  assign new_n7086 = new_n7069 & new_n7085;
  assign new_n7087 = ~new_n7069 & ~new_n7085;
  assign new_n7088 = ~new_n7086 & ~new_n7087;
  assign new_n7089 = new_n7061 & ~new_n7088;
  assign new_n7090 = ~new_n7061 & new_n7088;
  assign n2096 = ~new_n7089 & ~new_n7090;
  assign new_n7092 = ~new_n3988 & ~new_n3989;
  assign new_n7093 = new_n4024 & ~new_n7092;
  assign new_n7094 = ~new_n4024 & new_n7092;
  assign n2131 = ~new_n7093 & ~new_n7094;
  assign new_n7096 = n2564 & n11662;
  assign new_n7097 = n4189 & n7456;
  assign new_n7098 = ~new_n7096 & ~new_n7097;
  assign new_n7099 = new_n7096 & new_n7097;
  assign new_n7100 = ~new_n7098 & ~new_n7099;
  assign new_n7101 = n2564 & n7456;
  assign new_n7102 = new_n4351 & ~new_n4354;
  assign new_n7103 = ~new_n4355 & ~new_n7102;
  assign new_n7104 = ~new_n7101 & new_n7103;
  assign new_n7105 = new_n7101 & ~new_n7103;
  assign new_n7106 = n1798 & n9920;
  assign new_n7107 = n4189 & n12591;
  assign new_n7108 = n3932 & n6770;
  assign new_n7109 = ~new_n7107 & ~new_n7108;
  assign new_n7110 = new_n7107 & new_n7108;
  assign new_n7111 = ~new_n7109 & ~new_n7110;
  assign new_n7112 = new_n7106 & ~new_n7111;
  assign new_n7113 = ~new_n7106 & new_n7111;
  assign new_n7114 = ~new_n7112 & ~new_n7113;
  assign new_n7115 = ~new_n7105 & new_n7114;
  assign new_n7116 = ~new_n7104 & ~new_n7115;
  assign new_n7117 = new_n7100 & new_n7116;
  assign new_n7118 = ~new_n7100 & ~new_n7116;
  assign new_n7119 = ~new_n7117 & ~new_n7118;
  assign new_n7120 = n6770 & n12591;
  assign new_n7121 = n1798 & n3627;
  assign new_n7122 = n3932 & n9920;
  assign new_n7123 = ~new_n7121 & ~new_n7122;
  assign new_n7124 = new_n7121 & new_n7122;
  assign new_n7125 = ~new_n7123 & ~new_n7124;
  assign new_n7126 = new_n7120 & new_n7125;
  assign new_n7127 = ~new_n7120 & ~new_n7125;
  assign new_n7128 = ~new_n7126 & ~new_n7127;
  assign new_n7129 = ~new_n7106 & ~new_n7110;
  assign new_n7130 = ~new_n7109 & ~new_n7129;
  assign new_n7131 = ~new_n7128 & new_n7130;
  assign new_n7132 = new_n7128 & ~new_n7130;
  assign new_n7133 = ~new_n7131 & ~new_n7132;
  assign new_n7134 = new_n7119 & new_n7133;
  assign new_n7135 = ~new_n7119 & ~new_n7133;
  assign new_n7136 = ~new_n7134 & ~new_n7135;
  assign new_n7137 = n6687 & n11662;
  assign new_n7138 = ~new_n4348 & ~new_n4359;
  assign new_n7139 = ~new_n4349 & ~new_n7138;
  assign new_n7140 = new_n7137 & ~new_n7139;
  assign new_n7141 = ~new_n7137 & new_n7139;
  assign new_n7142 = ~new_n7104 & ~new_n7105;
  assign new_n7143 = new_n7114 & ~new_n7142;
  assign new_n7144 = ~new_n7114 & new_n7142;
  assign new_n7145 = ~new_n7143 & ~new_n7144;
  assign new_n7146 = ~new_n7141 & new_n7145;
  assign new_n7147 = ~new_n7140 & ~new_n7146;
  assign new_n7148 = ~new_n7136 & ~new_n7147;
  assign new_n7149 = ~new_n7118 & ~new_n7133;
  assign new_n7150 = ~new_n7099 & ~new_n7149;
  assign new_n7151 = ~new_n7117 & new_n7150;
  assign new_n7152 = new_n7099 & new_n7149;
  assign new_n7153 = ~new_n7151 & ~new_n7152;
  assign new_n7154 = n2564 & n10327;
  assign new_n7155 = n4189 & n11662;
  assign new_n7156 = n6687 & n9583;
  assign new_n7157 = ~new_n7155 & ~new_n7156;
  assign new_n7158 = new_n7155 & new_n7156;
  assign new_n7159_1 = ~new_n7157 & ~new_n7158;
  assign new_n7160_1 = ~new_n7154 & ~new_n7159_1;
  assign new_n7161 = new_n7154 & new_n7159_1;
  assign new_n7162 = ~new_n7160_1 & ~new_n7161;
  assign new_n7163 = ~new_n7126 & ~new_n7130;
  assign new_n7164 = ~new_n7127 & ~new_n7163;
  assign new_n7165 = ~new_n7162 & ~new_n7164;
  assign new_n7166 = n6770 & n7456;
  assign new_n7167 = new_n7124 & new_n7166;
  assign new_n7168 = ~new_n7124 & ~new_n7166;
  assign new_n7169 = ~new_n7167 & ~new_n7168;
  assign new_n7170 = n1798 & n4516;
  assign new_n7171 = n3627 & n3932;
  assign new_n7172 = n9920 & n12591;
  assign new_n7173 = ~new_n7171 & ~new_n7172;
  assign new_n7174 = new_n7171 & new_n7172;
  assign new_n7175 = ~new_n7173 & ~new_n7174;
  assign new_n7176 = new_n7170 & ~new_n7175;
  assign new_n7177 = ~new_n7170 & new_n7175;
  assign new_n7178 = ~new_n7176 & ~new_n7177;
  assign new_n7179 = new_n7169 & new_n7178;
  assign new_n7180 = ~new_n7169 & ~new_n7178;
  assign new_n7181 = ~new_n7179 & ~new_n7180;
  assign new_n7182 = new_n7165 & new_n7181;
  assign new_n7183 = new_n7162 & new_n7164;
  assign new_n7184 = new_n7181 & ~new_n7183;
  assign new_n7185 = ~new_n7165 & ~new_n7184;
  assign new_n7186 = ~new_n7182 & ~new_n7185;
  assign new_n7187 = ~new_n7181 & new_n7183;
  assign new_n7188 = ~new_n7186 & ~new_n7187;
  assign new_n7189 = ~new_n7153 & ~new_n7188;
  assign new_n7190 = new_n7153 & new_n7188;
  assign new_n7191 = ~new_n7189 & ~new_n7190;
  assign new_n7192 = ~new_n7148 & new_n7191;
  assign new_n7193_1 = new_n7148 & ~new_n7191;
  assign new_n7194 = ~new_n7192 & ~new_n7193_1;
  assign new_n7195 = n6687 & n10327;
  assign new_n7196 = new_n7136 & new_n7147;
  assign new_n7197 = ~new_n7148 & ~new_n7196;
  assign new_n7198 = new_n7195 & new_n7197;
  assign new_n7199 = ~new_n7140 & ~new_n7141;
  assign new_n7200 = ~new_n7145 & ~new_n7199;
  assign new_n7201 = new_n7145 & new_n7199;
  assign new_n7202 = ~new_n7200 & ~new_n7201;
  assign new_n7203 = new_n4363 & new_n7202;
  assign new_n7204 = ~new_n7195 & ~new_n7197;
  assign new_n7205 = ~new_n7198 & ~new_n7204;
  assign new_n7206 = new_n7203 & new_n7205;
  assign new_n7207 = ~new_n7198 & ~new_n7206;
  assign new_n7208 = ~new_n7194 & new_n7207;
  assign new_n7209 = new_n7194 & ~new_n7207;
  assign new_n7210 = ~new_n7208 & ~new_n7209;
  assign new_n7211 = n8336 & n10278;
  assign new_n7212 = n8336 & n10451;
  assign new_n7213 = n10928 & n11023;
  assign new_n7214 = new_n4477 & ~new_n4480;
  assign new_n7215 = ~new_n4481 & ~new_n7214;
  assign new_n7216 = ~new_n7213 & new_n7215;
  assign new_n7217 = new_n7213 & ~new_n7215;
  assign new_n7218 = ~new_n7216 & ~new_n7217;
  assign new_n7219 = n1094 & n6703;
  assign new_n7220 = n3022 & n6986;
  assign new_n7221 = n2226 & n9640;
  assign new_n7222 = ~new_n7220 & ~new_n7221;
  assign new_n7223 = new_n7220 & new_n7221;
  assign new_n7224 = ~new_n7222 & ~new_n7223;
  assign new_n7225 = new_n7219 & ~new_n7224;
  assign new_n7226 = ~new_n7219 & new_n7224;
  assign new_n7227 = ~new_n7225 & ~new_n7226;
  assign new_n7228 = ~new_n7218 & new_n7227;
  assign new_n7229 = new_n7218 & ~new_n7227;
  assign new_n7230 = ~new_n7228 & ~new_n7229;
  assign new_n7231 = ~new_n7212 & ~new_n7230;
  assign new_n7232 = new_n7212 & new_n7230;
  assign new_n7233 = ~new_n4474 & ~new_n4485;
  assign new_n7234 = ~new_n4475 & ~new_n7233;
  assign new_n7235 = ~new_n7232 & new_n7234;
  assign new_n7236_1 = ~new_n7231 & ~new_n7235;
  assign new_n7237 = n10451 & n10928;
  assign new_n7238 = n6986 & n11023;
  assign new_n7239 = ~new_n7237 & ~new_n7238;
  assign new_n7240 = new_n7237 & new_n7238;
  assign new_n7241 = ~new_n7239 & ~new_n7240;
  assign new_n7242 = n2226 & n3022;
  assign new_n7243 = n1094 & n9640;
  assign new_n7244 = n6703 & n10678;
  assign new_n7245 = ~new_n7243 & ~new_n7244;
  assign new_n7246 = new_n7243 & new_n7244;
  assign new_n7247 = ~new_n7245 & ~new_n7246;
  assign new_n7248 = new_n7242 & new_n7247;
  assign new_n7249 = ~new_n7242 & ~new_n7247;
  assign new_n7250 = ~new_n7248 & ~new_n7249;
  assign new_n7251 = ~new_n7219 & ~new_n7223;
  assign new_n7252 = ~new_n7222 & ~new_n7251;
  assign new_n7253 = ~new_n7250 & new_n7252;
  assign new_n7254 = new_n7250 & ~new_n7252;
  assign new_n7255 = ~new_n7253 & ~new_n7254;
  assign new_n7256 = new_n7241 & ~new_n7255;
  assign new_n7257 = ~new_n7241 & new_n7255;
  assign new_n7258 = ~new_n7256 & ~new_n7257;
  assign new_n7259 = ~new_n7216 & ~new_n7227;
  assign new_n7260 = ~new_n7217 & ~new_n7259;
  assign new_n7261 = new_n7258 & new_n7260;
  assign new_n7262 = ~new_n7258 & ~new_n7260;
  assign new_n7263 = ~new_n7261 & ~new_n7262;
  assign new_n7264 = new_n7236_1 & ~new_n7263;
  assign new_n7265_1 = ~new_n7236_1 & new_n7263;
  assign new_n7266 = ~new_n7264 & ~new_n7265_1;
  assign new_n7267 = new_n7211 & new_n7266;
  assign new_n7268 = ~new_n7231 & ~new_n7232;
  assign new_n7269 = ~new_n7234 & ~new_n7268;
  assign new_n7270_1 = ~new_n7231 & new_n7235;
  assign new_n7271 = ~new_n7269 & ~new_n7270_1;
  assign new_n7272 = new_n4490 & ~new_n7271;
  assign new_n7273 = ~new_n7211 & ~new_n7266;
  assign new_n7274 = ~new_n7267 & ~new_n7273;
  assign new_n7275 = new_n7272 & new_n7274;
  assign new_n7276 = ~new_n7267 & ~new_n7275;
  assign new_n7277 = ~new_n7257 & ~new_n7260;
  assign new_n7278 = ~new_n7240 & ~new_n7277;
  assign new_n7279 = ~new_n7256 & new_n7278;
  assign new_n7280 = new_n7240 & new_n7277;
  assign new_n7281 = ~new_n7279 & ~new_n7280;
  assign new_n7282 = n10278 & n10928;
  assign new_n7283 = n6986 & n10451;
  assign new_n7284 = n8336 & n11423;
  assign new_n7285 = ~new_n7283 & ~new_n7284;
  assign new_n7286 = new_n7283 & new_n7284;
  assign new_n7287 = ~new_n7285 & ~new_n7286;
  assign new_n7288 = ~new_n7282 & ~new_n7287;
  assign new_n7289 = new_n7282 & new_n7287;
  assign new_n7290 = ~new_n7288 & ~new_n7289;
  assign new_n7291 = ~new_n7248 & ~new_n7252;
  assign new_n7292 = ~new_n7249 & ~new_n7291;
  assign new_n7293 = new_n7290 & new_n7292;
  assign new_n7294_1 = ~new_n7290 & ~new_n7292;
  assign new_n7295 = ~new_n7293 & ~new_n7294_1;
  assign new_n7296 = n2226 & n11023;
  assign new_n7297 = new_n7246 & new_n7296;
  assign new_n7298 = ~new_n7246 & ~new_n7296;
  assign new_n7299 = ~new_n7297 & ~new_n7298;
  assign new_n7300 = n9640 & n10678;
  assign new_n7301 = n6703 & n7320;
  assign new_n7302 = n1094 & n3022;
  assign new_n7303 = ~new_n7301 & ~new_n7302;
  assign new_n7304 = new_n7301 & new_n7302;
  assign new_n7305 = ~new_n7303 & ~new_n7304;
  assign new_n7306 = ~new_n7300 & ~new_n7305;
  assign new_n7307 = new_n7300 & new_n7305;
  assign new_n7308 = ~new_n7306 & ~new_n7307;
  assign new_n7309 = new_n7299 & ~new_n7308;
  assign new_n7310 = ~new_n7299 & new_n7308;
  assign new_n7311 = ~new_n7309 & ~new_n7310;
  assign new_n7312 = new_n7295 & new_n7311;
  assign new_n7313 = ~new_n7295 & ~new_n7311;
  assign new_n7314 = ~new_n7312 & ~new_n7313;
  assign new_n7315 = ~new_n7281 & new_n7314;
  assign new_n7316 = new_n7281 & ~new_n7314;
  assign new_n7317 = ~new_n7315 & ~new_n7316;
  assign new_n7318 = ~new_n7264 & ~new_n7317;
  assign new_n7319 = new_n7264 & new_n7317;
  assign new_n7320_1 = ~new_n7318 & ~new_n7319;
  assign new_n7321 = ~new_n7276 & new_n7320_1;
  assign new_n7322 = new_n7276 & ~new_n7320_1;
  assign new_n7323 = ~new_n7321 & ~new_n7322;
  assign new_n7324 = n12069 & n12826;
  assign new_n7325 = n2551 & n12069;
  assign new_n7326 = n11922 & n12391;
  assign new_n7327 = new_n4503 & ~new_n4506;
  assign new_n7328 = ~new_n4507 & ~new_n7327;
  assign new_n7329 = new_n7326 & ~new_n7328;
  assign new_n7330 = ~new_n7326 & new_n7328;
  assign new_n7331 = ~new_n7329 & ~new_n7330;
  assign new_n7332 = n1067 & n7160;
  assign new_n7333 = n7891 & n8665;
  assign new_n7334 = n4828 & n5645;
  assign new_n7335 = ~new_n7333 & ~new_n7334;
  assign new_n7336 = new_n7333 & new_n7334;
  assign new_n7337 = ~new_n7335 & ~new_n7336;
  assign new_n7338 = new_n7332 & ~new_n7337;
  assign new_n7339 = ~new_n7332 & new_n7337;
  assign new_n7340 = ~new_n7338 & ~new_n7339;
  assign new_n7341 = ~new_n7331 & ~new_n7340;
  assign new_n7342 = new_n7331 & new_n7340;
  assign new_n7343 = ~new_n7341 & ~new_n7342;
  assign new_n7344 = new_n7325 & ~new_n7343;
  assign new_n7345 = ~new_n7325 & new_n7343;
  assign new_n7346 = ~new_n4500 & new_n4511;
  assign new_n7347 = ~new_n4501 & ~new_n7346;
  assign new_n7348 = ~new_n7345 & new_n7347;
  assign new_n7349 = ~new_n7344 & ~new_n7348;
  assign new_n7350 = n2551 & n12391;
  assign new_n7351 = n7891 & n11922;
  assign new_n7352 = ~new_n7350 & ~new_n7351;
  assign new_n7353 = new_n7350 & new_n7351;
  assign new_n7354_1 = ~new_n7352 & ~new_n7353;
  assign new_n7355 = n7160 & n8665;
  assign new_n7356 = n1067 & n4828;
  assign new_n7357 = n2515 & n5645;
  assign new_n7358 = ~new_n7356 & ~new_n7357;
  assign new_n7359 = new_n7356 & new_n7357;
  assign new_n7360 = ~new_n7358 & ~new_n7359;
  assign new_n7361 = new_n7355 & new_n7360;
  assign new_n7362 = ~new_n7355 & ~new_n7360;
  assign new_n7363 = ~new_n7361 & ~new_n7362;
  assign new_n7364 = new_n7332 & ~new_n7335;
  assign new_n7365 = ~new_n7336 & ~new_n7364;
  assign new_n7366 = ~new_n7363 & ~new_n7365;
  assign new_n7367 = new_n7363 & new_n7365;
  assign new_n7368 = ~new_n7366 & ~new_n7367;
  assign new_n7369 = new_n7354_1 & ~new_n7368;
  assign new_n7370 = ~new_n7354_1 & new_n7368;
  assign new_n7371 = ~new_n7369 & ~new_n7370;
  assign new_n7372 = ~new_n7330 & ~new_n7340;
  assign new_n7373 = ~new_n7329 & ~new_n7372;
  assign new_n7374 = new_n7371 & new_n7373;
  assign new_n7375 = ~new_n7371 & ~new_n7373;
  assign new_n7376 = ~new_n7374 & ~new_n7375;
  assign new_n7377 = ~new_n7349 & ~new_n7376;
  assign new_n7378 = new_n7349 & new_n7376;
  assign new_n7379 = ~new_n7377 & ~new_n7378;
  assign new_n7380 = new_n7324 & new_n7379;
  assign new_n7381 = ~new_n7344 & ~new_n7345;
  assign new_n7382 = ~new_n7347 & ~new_n7381;
  assign new_n7383 = new_n7347 & new_n7381;
  assign new_n7384 = ~new_n7382 & ~new_n7383;
  assign new_n7385 = new_n4516_1 & new_n7384;
  assign new_n7386 = ~new_n7324 & ~new_n7379;
  assign new_n7387 = ~new_n7380 & ~new_n7386;
  assign new_n7388_1 = new_n7385 & new_n7387;
  assign new_n7389 = ~new_n7380 & ~new_n7388_1;
  assign new_n7390 = ~new_n7370 & ~new_n7373;
  assign new_n7391 = ~new_n7353 & ~new_n7390;
  assign new_n7392 = ~new_n7369 & new_n7391;
  assign new_n7393 = new_n7353 & new_n7390;
  assign new_n7394 = ~new_n7392 & ~new_n7393;
  assign new_n7395 = n12391 & n12826;
  assign new_n7396 = n2551 & n7891;
  assign new_n7397 = n4094 & n12069;
  assign new_n7398 = ~new_n7396 & ~new_n7397;
  assign new_n7399 = new_n7396 & new_n7397;
  assign new_n7400 = ~new_n7398 & ~new_n7399;
  assign new_n7401 = ~new_n7395 & ~new_n7400;
  assign new_n7402 = new_n7395 & new_n7400;
  assign new_n7403 = ~new_n7401 & ~new_n7402;
  assign new_n7404 = ~new_n7362 & ~new_n7365;
  assign new_n7405 = ~new_n7361 & ~new_n7404;
  assign new_n7406 = new_n7403 & ~new_n7405;
  assign new_n7407 = ~new_n7403 & new_n7405;
  assign new_n7408 = ~new_n7406 & ~new_n7407;
  assign new_n7409 = n7160 & n11922;
  assign new_n7410 = ~new_n7359 & ~new_n7409;
  assign new_n7411 = new_n7359 & new_n7409;
  assign new_n7412 = ~new_n7410 & ~new_n7411;
  assign new_n7413 = n1199 & n5645;
  assign new_n7414 = n4828 & n8665;
  assign new_n7415 = n1067 & n2515;
  assign new_n7416 = ~new_n7414 & ~new_n7415;
  assign new_n7417 = new_n7414 & new_n7415;
  assign new_n7418 = ~new_n7416 & ~new_n7417;
  assign new_n7419 = new_n7413 & ~new_n7418;
  assign new_n7420 = ~new_n7413 & new_n7418;
  assign new_n7421 = ~new_n7419 & ~new_n7420;
  assign new_n7422 = new_n7412 & new_n7421;
  assign new_n7423 = ~new_n7412 & ~new_n7421;
  assign new_n7424 = ~new_n7422 & ~new_n7423;
  assign new_n7425 = ~new_n7408 & ~new_n7424;
  assign new_n7426 = new_n7408 & new_n7424;
  assign new_n7427 = ~new_n7425 & ~new_n7426;
  assign new_n7428 = ~new_n7394 & new_n7427;
  assign new_n7429 = new_n7394 & ~new_n7427;
  assign new_n7430 = ~new_n7428 & ~new_n7429;
  assign new_n7431 = ~new_n7377 & ~new_n7430;
  assign new_n7432 = new_n7377 & new_n7430;
  assign new_n7433 = ~new_n7431 & ~new_n7432;
  assign new_n7434 = ~new_n7389 & new_n7433;
  assign new_n7435 = new_n7389 & ~new_n7433;
  assign new_n7436_1 = ~new_n7434 & ~new_n7435;
  assign new_n7437 = n1510 & n11222;
  assign new_n7438 = n159 & n11222;
  assign new_n7439 = n2749 & n11153;
  assign new_n7440 = new_n4524 & ~new_n4527;
  assign new_n7441 = ~new_n4528 & ~new_n7440;
  assign new_n7442 = ~new_n7439 & new_n7441;
  assign new_n7443 = new_n7439 & ~new_n7441;
  assign new_n7444 = ~new_n7442 & ~new_n7443;
  assign new_n7445 = n5767 & n11876;
  assign new_n7446 = n3754 & n5314;
  assign new_n7447 = n996 & n10898;
  assign new_n7448 = ~new_n7446 & ~new_n7447;
  assign new_n7449 = new_n7446 & new_n7447;
  assign new_n7450 = ~new_n7448 & ~new_n7449;
  assign new_n7451 = new_n7445 & ~new_n7450;
  assign new_n7452 = ~new_n7445 & new_n7450;
  assign new_n7453 = ~new_n7451 & ~new_n7452;
  assign new_n7454 = ~new_n7444 & new_n7453;
  assign new_n7455 = new_n7444 & ~new_n7453;
  assign new_n7456_1 = ~new_n7454 & ~new_n7455;
  assign new_n7457 = ~new_n7438 & ~new_n7456_1;
  assign new_n7458 = new_n7438 & new_n7456_1;
  assign new_n7459 = ~new_n4522 & ~new_n4532;
  assign new_n7460 = ~new_n4521 & ~new_n7459;
  assign new_n7461 = ~new_n7458 & new_n7460;
  assign new_n7462 = ~new_n7457 & ~new_n7461;
  assign new_n7463 = n159 & n11153;
  assign new_n7464 = n2749 & n5314;
  assign new_n7465 = ~new_n7463 & ~new_n7464;
  assign new_n7466 = new_n7463 & new_n7464;
  assign new_n7467 = ~new_n7465 & ~new_n7466;
  assign new_n7468 = n996 & n3754;
  assign new_n7469 = n5767 & n10898;
  assign new_n7470 = n5319 & n11876;
  assign new_n7471 = ~new_n7469 & ~new_n7470;
  assign new_n7472 = new_n7469 & new_n7470;
  assign new_n7473 = ~new_n7471 & ~new_n7472;
  assign new_n7474 = new_n7468 & new_n7473;
  assign new_n7475 = ~new_n7468 & ~new_n7473;
  assign new_n7476 = ~new_n7474 & ~new_n7475;
  assign new_n7477 = new_n7445 & ~new_n7448;
  assign new_n7478 = ~new_n7449 & ~new_n7477;
  assign new_n7479 = ~new_n7476 & ~new_n7478;
  assign new_n7480 = new_n7476 & new_n7478;
  assign new_n7481 = ~new_n7479 & ~new_n7480;
  assign new_n7482 = new_n7467 & ~new_n7481;
  assign new_n7483 = ~new_n7467 & new_n7481;
  assign new_n7484 = ~new_n7482 & ~new_n7483;
  assign new_n7485 = ~new_n7442 & ~new_n7453;
  assign new_n7486 = ~new_n7443 & ~new_n7485;
  assign new_n7487 = new_n7484 & new_n7486;
  assign new_n7488 = ~new_n7484 & ~new_n7486;
  assign new_n7489 = ~new_n7487 & ~new_n7488;
  assign new_n7490 = new_n7462 & ~new_n7489;
  assign new_n7491 = ~new_n7462 & new_n7489;
  assign new_n7492 = ~new_n7490 & ~new_n7491;
  assign new_n7493 = new_n7437 & new_n7492;
  assign new_n7494 = ~new_n7457 & ~new_n7458;
  assign new_n7495 = ~new_n7460 & ~new_n7494;
  assign new_n7496 = new_n7460 & new_n7494;
  assign new_n7497 = ~new_n7495 & ~new_n7496;
  assign new_n7498 = new_n4536 & ~new_n7497;
  assign new_n7499 = ~new_n7437 & ~new_n7492;
  assign new_n7500_1 = ~new_n7493 & ~new_n7499;
  assign new_n7501 = new_n7498 & new_n7500_1;
  assign new_n7502 = ~new_n7493 & ~new_n7501;
  assign new_n7503 = ~new_n7483 & ~new_n7486;
  assign new_n7504 = ~new_n7466 & ~new_n7503;
  assign new_n7505 = ~new_n7482 & new_n7504;
  assign new_n7506 = new_n7466 & new_n7503;
  assign new_n7507 = ~new_n7505 & ~new_n7506;
  assign new_n7508 = n1510 & n11153;
  assign new_n7509 = n159 & n5314;
  assign new_n7510 = n11222 & n12247;
  assign new_n7511 = ~new_n7509 & ~new_n7510;
  assign new_n7512 = new_n7509 & new_n7510;
  assign new_n7513 = ~new_n7511 & ~new_n7512;
  assign new_n7514 = ~new_n7508 & ~new_n7513;
  assign new_n7515 = new_n7508 & new_n7513;
  assign new_n7516 = ~new_n7514 & ~new_n7515;
  assign new_n7517 = ~new_n7474 & new_n7478;
  assign new_n7518 = ~new_n7475 & ~new_n7517;
  assign new_n7519 = new_n7516 & new_n7518;
  assign new_n7520 = ~new_n7516 & ~new_n7518;
  assign new_n7521 = ~new_n7519 & ~new_n7520;
  assign new_n7522 = n996 & n2749;
  assign new_n7523_1 = new_n7472 & new_n7522;
  assign new_n7524 = ~new_n7472 & ~new_n7522;
  assign new_n7525 = ~new_n7523_1 & ~new_n7524;
  assign new_n7526 = n5319 & n10898;
  assign new_n7527 = n9457 & n11876;
  assign new_n7528 = n3754 & n5767;
  assign new_n7529 = ~new_n7527 & ~new_n7528;
  assign new_n7530 = new_n7527 & new_n7528;
  assign new_n7531 = ~new_n7529 & ~new_n7530;
  assign new_n7532 = ~new_n7526 & ~new_n7531;
  assign new_n7533 = new_n7526 & new_n7531;
  assign new_n7534 = ~new_n7532 & ~new_n7533;
  assign new_n7535 = new_n7525 & ~new_n7534;
  assign new_n7536 = ~new_n7525 & new_n7534;
  assign new_n7537 = ~new_n7535 & ~new_n7536;
  assign new_n7538 = new_n7521 & new_n7537;
  assign new_n7539 = ~new_n7521 & ~new_n7537;
  assign new_n7540 = ~new_n7538 & ~new_n7539;
  assign new_n7541 = ~new_n7507 & new_n7540;
  assign new_n7542 = new_n7507 & ~new_n7540;
  assign new_n7543 = ~new_n7541 & ~new_n7542;
  assign new_n7544 = ~new_n7490 & ~new_n7543;
  assign new_n7545 = new_n7490 & new_n7543;
  assign new_n7546_1 = ~new_n7544 & ~new_n7545;
  assign new_n7547 = ~new_n7502 & new_n7546_1;
  assign new_n7548 = new_n7502 & ~new_n7546_1;
  assign new_n7549 = ~new_n7547 & ~new_n7548;
  assign new_n7550 = ~new_n7498 & ~new_n7500_1;
  assign new_n7551 = ~new_n7501 & ~new_n7550;
  assign new_n7552 = ~new_n7385 & ~new_n7387;
  assign new_n7553 = ~new_n7388_1 & ~new_n7552;
  assign new_n7554 = new_n7551 & new_n7553;
  assign new_n7555 = ~new_n7551 & ~new_n7553;
  assign new_n7556 = ~new_n4516_1 & ~new_n7384;
  assign new_n7557 = ~new_n7385 & ~new_n7556;
  assign new_n7558 = ~new_n4540 & ~new_n4543;
  assign new_n7559 = ~new_n4539 & ~new_n7558;
  assign new_n7560 = new_n7557 & ~new_n7559;
  assign new_n7561 = ~new_n7557 & new_n7559;
  assign new_n7562 = ~new_n4536 & new_n7497;
  assign new_n7563 = ~new_n7498 & ~new_n7562;
  assign new_n7564 = ~new_n7561 & new_n7563;
  assign new_n7565 = ~new_n7560 & ~new_n7564;
  assign new_n7566 = ~new_n7555 & ~new_n7565;
  assign new_n7567 = ~new_n7554 & ~new_n7566;
  assign new_n7568_1 = new_n7549 & ~new_n7567;
  assign new_n7569 = ~new_n7549 & new_n7567;
  assign new_n7570 = ~new_n7568_1 & ~new_n7569;
  assign new_n7571 = ~new_n7436_1 & new_n7570;
  assign new_n7572 = new_n7436_1 & ~new_n7570;
  assign new_n7573 = ~new_n7571 & ~new_n7572;
  assign new_n7574 = new_n7323 & ~new_n7573;
  assign new_n7575 = ~new_n7323 & new_n7573;
  assign new_n7576 = ~new_n7574 & ~new_n7575;
  assign new_n7577 = ~new_n7272 & ~new_n7274;
  assign new_n7578 = ~new_n7275 & ~new_n7577;
  assign new_n7579 = ~new_n4490 & new_n7271;
  assign new_n7580 = ~new_n7272 & ~new_n7579;
  assign new_n7581 = ~new_n7560 & ~new_n7561;
  assign new_n7582 = new_n7563 & new_n7581;
  assign new_n7583 = ~new_n7563 & ~new_n7581;
  assign new_n7584 = ~new_n7582 & ~new_n7583;
  assign new_n7585 = ~new_n7580 & ~new_n7584;
  assign new_n7586 = new_n7580 & new_n7584;
  assign new_n7587 = ~new_n4495 & ~new_n4546;
  assign new_n7588 = ~new_n4494 & ~new_n7587;
  assign new_n7589 = ~new_n7586 & new_n7588;
  assign new_n7590 = ~new_n7585 & ~new_n7589;
  assign new_n7591 = new_n7578 & new_n7590;
  assign new_n7592 = ~new_n7578 & ~new_n7590;
  assign new_n7593 = ~new_n7554 & ~new_n7555;
  assign new_n7594 = new_n7565 & ~new_n7593;
  assign new_n7595 = ~new_n7565 & new_n7593;
  assign new_n7596 = ~new_n7594 & ~new_n7595;
  assign new_n7597 = ~new_n7592 & new_n7596;
  assign new_n7598 = ~new_n7591 & ~new_n7597;
  assign new_n7599 = ~new_n7576 & ~new_n7598;
  assign new_n7600 = new_n7576 & new_n7598;
  assign new_n7601 = ~new_n7599 & ~new_n7600;
  assign new_n7602 = new_n7210 & ~new_n7601;
  assign new_n7603 = ~new_n7210 & new_n7601;
  assign new_n7604 = ~new_n7602 & ~new_n7603;
  assign new_n7605 = ~new_n7203 & ~new_n7205;
  assign new_n7606 = ~new_n7206 & ~new_n7605;
  assign new_n7607 = ~new_n7591 & ~new_n7592;
  assign new_n7608 = ~new_n7596 & ~new_n7607;
  assign new_n7609 = new_n7596 & new_n7607;
  assign new_n7610_1 = ~new_n7608 & ~new_n7609;
  assign new_n7611 = new_n7606 & new_n7610_1;
  assign new_n7612 = ~new_n7606 & ~new_n7610_1;
  assign new_n7613 = ~new_n4363 & ~new_n7202;
  assign new_n7614 = ~new_n7203 & ~new_n7613;
  assign new_n7615 = ~new_n7585 & ~new_n7586;
  assign new_n7616 = ~new_n7588 & ~new_n7615;
  assign new_n7617 = new_n7588 & new_n7615;
  assign new_n7618 = ~new_n7616 & ~new_n7617;
  assign new_n7619 = new_n7614 & ~new_n7618;
  assign new_n7620 = ~new_n7614 & new_n7618;
  assign new_n7621 = ~new_n4469 & new_n4549;
  assign new_n7622 = ~new_n4468 & ~new_n7621;
  assign new_n7623 = ~new_n7620 & ~new_n7622;
  assign new_n7624 = ~new_n7619 & ~new_n7623;
  assign new_n7625 = ~new_n7612 & ~new_n7624;
  assign new_n7626 = ~new_n7611 & ~new_n7625;
  assign new_n7627 = ~new_n7604 & ~new_n7626;
  assign new_n7628 = new_n7604 & new_n7626;
  assign n2301 = new_n7627 | new_n7628;
  assign new_n7630 = ~new_n4450 & ~new_n4451;
  assign new_n7631 = new_n4465 & ~new_n7630;
  assign new_n7632 = ~new_n4465 & new_n7630;
  assign n2316 = ~new_n7631 & ~new_n7632;
  assign new_n7634 = n7862 & n9195;
  assign new_n7635 = n1333 & n4634;
  assign new_n7636 = new_n6839 & ~new_n6842;
  assign new_n7637 = ~new_n6843 & ~new_n7636;
  assign new_n7638 = ~new_n7635 & new_n7637;
  assign new_n7639 = new_n7635 & ~new_n7637;
  assign new_n7640 = ~new_n7638 & ~new_n7639;
  assign new_n7641 = n5240 & n7265;
  assign new_n7642 = n3172 & n10223;
  assign new_n7643 = n2879 & n11757;
  assign new_n7644 = ~new_n7642 & ~new_n7643;
  assign new_n7645 = new_n7642 & new_n7643;
  assign new_n7646_1 = ~new_n7644 & ~new_n7645;
  assign new_n7647 = new_n7641 & ~new_n7646_1;
  assign new_n7648 = ~new_n7641 & new_n7646_1;
  assign new_n7649 = ~new_n7647 & ~new_n7648;
  assign new_n7650 = ~new_n7640 & new_n7649;
  assign new_n7651 = new_n7640 & ~new_n7649;
  assign new_n7652 = ~new_n7650 & ~new_n7651;
  assign new_n7653 = ~new_n7634 & ~new_n7652;
  assign new_n7654 = new_n7634 & new_n7652;
  assign new_n7655 = ~new_n6836 & ~new_n6847;
  assign new_n7656 = ~new_n6837 & ~new_n7655;
  assign new_n7657 = ~new_n7654 & new_n7656;
  assign new_n7658 = ~new_n7653 & ~new_n7657;
  assign new_n7659 = n3172 & n4634;
  assign new_n7660 = n1333 & n9195;
  assign new_n7661 = new_n7659 & new_n7660;
  assign new_n7662 = ~new_n7659 & ~new_n7660;
  assign new_n7663 = ~new_n7661 & ~new_n7662;
  assign new_n7664 = ~new_n7639 & new_n7649;
  assign new_n7665 = ~new_n7638 & ~new_n7664;
  assign new_n7666 = ~new_n7663 & ~new_n7665;
  assign new_n7667 = new_n7663 & new_n7665;
  assign new_n7668 = ~new_n7666 & ~new_n7667;
  assign new_n7669 = n10223 & n11757;
  assign new_n7670 = n2879 & n5240;
  assign new_n7671 = n7265 & n11821;
  assign new_n7672 = ~new_n7670 & ~new_n7671;
  assign new_n7673 = new_n7670 & new_n7671;
  assign new_n7674 = ~new_n7672 & ~new_n7673;
  assign new_n7675 = ~new_n7669 & ~new_n7674;
  assign new_n7676_1 = new_n7669 & new_n7674;
  assign new_n7677 = ~new_n7675 & ~new_n7676_1;
  assign new_n7678 = new_n7641 & ~new_n7644;
  assign new_n7679 = ~new_n7645 & ~new_n7678;
  assign new_n7680 = ~new_n7677 & ~new_n7679;
  assign new_n7681 = new_n7677 & new_n7679;
  assign new_n7682 = ~new_n7680 & ~new_n7681;
  assign new_n7683 = ~new_n7668 & new_n7682;
  assign new_n7684 = new_n7668 & ~new_n7682;
  assign new_n7685 = ~new_n7683 & ~new_n7684;
  assign new_n7686 = new_n7658 & new_n7685;
  assign new_n7687 = ~new_n7666 & ~new_n7682;
  assign new_n7688 = new_n7661 & new_n7687;
  assign new_n7689 = ~new_n7661 & ~new_n7687;
  assign new_n7690_1 = ~new_n7667 & new_n7689;
  assign new_n7691 = n3172 & n9195;
  assign new_n7692 = n3865 & n7862;
  assign new_n7693 = n1333 & n2253;
  assign new_n7694 = ~new_n7692 & ~new_n7693;
  assign new_n7695 = new_n7692 & new_n7693;
  assign new_n7696 = ~new_n7694 & ~new_n7695;
  assign new_n7697 = new_n7691 & ~new_n7696;
  assign new_n7698 = ~new_n7691 & new_n7696;
  assign new_n7699 = ~new_n7697 & ~new_n7698;
  assign new_n7700 = ~new_n7676_1 & new_n7679;
  assign new_n7701 = ~new_n7675 & ~new_n7700;
  assign new_n7702 = new_n7699 & ~new_n7701;
  assign new_n7703 = ~new_n7699 & new_n7701;
  assign new_n7704 = ~new_n7702 & ~new_n7703;
  assign new_n7705 = n4634 & n11757;
  assign new_n7706 = new_n7673 & new_n7705;
  assign new_n7707 = ~new_n7673 & ~new_n7705;
  assign new_n7708 = ~new_n7706 & ~new_n7707;
  assign new_n7709 = n2879 & n11821;
  assign new_n7710 = n5240 & n10223;
  assign new_n7711 = n7265 & n9080;
  assign new_n7712 = ~new_n7710 & ~new_n7711;
  assign new_n7713 = new_n7710 & new_n7711;
  assign new_n7714 = ~new_n7712 & ~new_n7713;
  assign new_n7715 = ~new_n7709 & ~new_n7714;
  assign new_n7716 = new_n7709 & new_n7714;
  assign new_n7717 = ~new_n7715 & ~new_n7716;
  assign new_n7718 = new_n7708 & ~new_n7717;
  assign new_n7719 = ~new_n7708 & new_n7717;
  assign new_n7720 = ~new_n7718 & ~new_n7719;
  assign new_n7721 = new_n7704 & new_n7720;
  assign new_n7722 = ~new_n7704 & ~new_n7720;
  assign new_n7723 = ~new_n7721 & ~new_n7722;
  assign new_n7724 = ~new_n7690_1 & ~new_n7723;
  assign new_n7725 = ~new_n7688 & ~new_n7724;
  assign new_n7726 = new_n7690_1 & new_n7723;
  assign new_n7727 = new_n7725 & ~new_n7726;
  assign new_n7728 = new_n7688 & ~new_n7723;
  assign new_n7729 = ~new_n7727 & ~new_n7728;
  assign new_n7730_1 = ~new_n7686 & new_n7729;
  assign new_n7731 = new_n7686 & ~new_n7729;
  assign new_n7732 = ~new_n7730_1 & ~new_n7731;
  assign new_n7733_1 = n2253 & n7862;
  assign new_n7734 = ~new_n7658 & ~new_n7685;
  assign new_n7735 = ~new_n7686 & ~new_n7734;
  assign new_n7736 = new_n7733_1 & new_n7735;
  assign new_n7737 = ~new_n7653 & ~new_n7654;
  assign new_n7738 = new_n7656 & ~new_n7737;
  assign new_n7739 = ~new_n7656 & new_n7737;
  assign new_n7740 = ~new_n7738 & ~new_n7739;
  assign new_n7741 = new_n6851 & new_n7740;
  assign new_n7742 = ~new_n7733_1 & ~new_n7735;
  assign new_n7743 = ~new_n7736 & ~new_n7742;
  assign new_n7744 = new_n7741 & new_n7743;
  assign new_n7745 = ~new_n7736 & ~new_n7744;
  assign new_n7746 = ~new_n7732 & new_n7745;
  assign new_n7747 = new_n7732 & ~new_n7745;
  assign new_n7748 = ~new_n7746 & ~new_n7747;
  assign new_n7749 = ~new_n7741 & ~new_n7743;
  assign new_n7750 = ~new_n7744 & ~new_n7749;
  assign new_n7751 = ~new_n6851 & ~new_n7740;
  assign new_n7752 = ~new_n7741 & ~new_n7751;
  assign new_n7753 = n6877 & n12145;
  assign new_n7754 = n2522 & n9400;
  assign new_n7755 = n4187 & n7946;
  assign new_n7756 = n2464 & n9189;
  assign new_n7757 = n2024 & n11311;
  assign new_n7758 = ~new_n7756 & ~new_n7757;
  assign new_n7759 = new_n7756 & new_n7757;
  assign new_n7760 = ~new_n7758 & ~new_n7759;
  assign new_n7761 = new_n7755 & ~new_n7760;
  assign new_n7762 = ~new_n7755 & new_n7760;
  assign new_n7763 = ~new_n7761 & ~new_n7762;
  assign new_n7764 = new_n7754 & ~new_n7763;
  assign new_n7765 = ~new_n7754 & new_n7763;
  assign new_n7766 = ~new_n7764 & ~new_n7765;
  assign new_n7767 = new_n6868 & ~new_n6871;
  assign new_n7768 = ~new_n6872 & ~new_n7767;
  assign new_n7769 = ~new_n7766 & ~new_n7768;
  assign new_n7770 = new_n7766 & new_n7768;
  assign new_n7771 = ~new_n7769 & ~new_n7770;
  assign new_n7772 = new_n7753 & ~new_n7771;
  assign new_n7773 = ~new_n7753 & new_n7771;
  assign new_n7774 = ~new_n7772 & ~new_n7773;
  assign new_n7775 = ~new_n6878 & ~new_n6881;
  assign new_n7776 = ~new_n6877_1 & ~new_n7775;
  assign new_n7777 = ~new_n7774 & ~new_n7776;
  assign new_n7778 = new_n7774 & new_n7776;
  assign new_n7779 = ~new_n7777 & ~new_n7778;
  assign new_n7780 = new_n6886 & ~new_n7779;
  assign new_n7781 = ~new_n6886 & new_n7779;
  assign new_n7782 = ~new_n7780 & ~new_n7781;
  assign new_n7783 = ~new_n6957 & ~new_n7009;
  assign new_n7784 = ~new_n6956 & ~new_n7783;
  assign new_n7785 = new_n7782 & ~new_n7784;
  assign new_n7786 = ~new_n7782 & new_n7784;
  assign new_n7787 = ~new_n7785 & ~new_n7786;
  assign new_n7788 = n4805 & n6016;
  assign new_n7789 = ~new_n6964 & ~new_n6974;
  assign new_n7790 = ~new_n6963 & ~new_n7789;
  assign new_n7791 = new_n7788 & ~new_n7790;
  assign new_n7792 = ~new_n7788 & new_n7790;
  assign new_n7793 = ~new_n7791 & ~new_n7792;
  assign new_n7794 = n2558 & n6294;
  assign new_n7795 = n137 & n2498;
  assign new_n7796 = ~new_n6928 & ~new_n7795;
  assign new_n7797 = new_n6928 & new_n7795;
  assign new_n7798 = ~new_n7796 & ~new_n7797;
  assign new_n7799 = new_n7794 & ~new_n7798;
  assign new_n7800 = ~new_n7794 & new_n7798;
  assign new_n7801 = ~new_n7799 & ~new_n7800;
  assign new_n7802 = n521 & n11478;
  assign new_n7803 = new_n6966 & ~new_n6969;
  assign new_n7804 = ~new_n6970 & ~new_n7803;
  assign new_n7805 = new_n7802 & ~new_n7804;
  assign new_n7806 = ~new_n7802 & new_n7804;
  assign new_n7807 = ~new_n7805 & ~new_n7806;
  assign new_n7808 = ~new_n7801 & ~new_n7807;
  assign new_n7809 = new_n7801 & new_n7807;
  assign new_n7810 = ~new_n7808 & ~new_n7809;
  assign new_n7811 = ~new_n7793 & ~new_n7810;
  assign new_n7812 = new_n7793 & new_n7810;
  assign new_n7813 = ~new_n7811 & ~new_n7812;
  assign new_n7814 = new_n6978 & ~new_n7813;
  assign new_n7815 = ~new_n6978 & new_n7813;
  assign new_n7816 = ~new_n7814 & ~new_n7815;
  assign new_n7817 = n7236 & n7270;
  assign new_n7818 = ~new_n6985 & ~new_n6995;
  assign new_n7819 = ~new_n6984 & ~new_n7818;
  assign new_n7820 = new_n7817 & ~new_n7819;
  assign new_n7821 = ~new_n7817 & new_n7819;
  assign new_n7822 = ~new_n7820 & ~new_n7821;
  assign new_n7823_1 = n806 & n3992;
  assign new_n7824 = new_n6987 & ~new_n6990;
  assign new_n7825 = ~new_n6991 & ~new_n7824;
  assign new_n7826 = new_n7823_1 & ~new_n7825;
  assign new_n7827 = ~new_n7823_1 & new_n7825;
  assign new_n7828 = ~new_n7826 & ~new_n7827;
  assign new_n7829 = n6358 & n9111;
  assign new_n7830 = n5198 & n9763;
  assign new_n7831 = ~new_n6938 & ~new_n7830;
  assign new_n7832 = n3342 & n5198;
  assign new_n7833 = new_n6935 & new_n7832;
  assign new_n7834 = ~new_n7831 & ~new_n7833;
  assign new_n7835 = ~new_n7829 & ~new_n7834;
  assign new_n7836 = new_n7829 & new_n7834;
  assign new_n7837 = ~new_n7835 & ~new_n7836;
  assign new_n7838 = ~new_n7828 & ~new_n7837;
  assign new_n7839 = new_n7828 & new_n7837;
  assign new_n7840 = ~new_n7838 & ~new_n7839;
  assign new_n7841 = new_n7822 & new_n7840;
  assign new_n7842 = ~new_n7822 & ~new_n7840;
  assign new_n7843 = ~new_n7841 & ~new_n7842;
  assign new_n7844 = new_n6999 & new_n7843;
  assign new_n7845 = ~new_n6999 & ~new_n7843;
  assign new_n7846 = ~new_n7844 & ~new_n7845;
  assign new_n7847 = ~new_n7816 & ~new_n7846;
  assign new_n7848 = new_n7816 & new_n7846;
  assign new_n7849 = ~new_n7847 & ~new_n7848;
  assign new_n7850 = new_n7006 & new_n7849;
  assign new_n7851 = ~new_n7006 & ~new_n7849;
  assign new_n7852 = ~new_n7850 & ~new_n7851;
  assign new_n7853 = ~new_n7787 & new_n7852;
  assign new_n7854 = new_n7787 & ~new_n7852;
  assign new_n7855 = ~new_n7853 & ~new_n7854;
  assign new_n7856 = ~new_n7752 & new_n7855;
  assign new_n7857 = new_n7752 & ~new_n7855;
  assign new_n7858 = ~new_n7013 & ~new_n7039;
  assign new_n7859 = ~new_n7014 & ~new_n7858;
  assign new_n7860 = ~new_n7857 & ~new_n7859;
  assign new_n7861 = ~new_n7856 & ~new_n7860;
  assign new_n7862_1 = new_n7750 & new_n7861;
  assign new_n7863 = ~new_n7750 & ~new_n7861;
  assign new_n7864 = n6877 & n12221;
  assign new_n7865 = n9400 & n12145;
  assign new_n7866 = n2464 & n2522;
  assign new_n7867 = ~new_n7865 & ~new_n7866;
  assign new_n7868 = new_n7865 & new_n7866;
  assign new_n7869 = ~new_n7867 & ~new_n7868;
  assign new_n7870 = n9189 & n11311;
  assign new_n7871 = n4203 & n7946;
  assign new_n7872 = n2024 & n4187;
  assign new_n7873 = ~new_n7871 & ~new_n7872;
  assign new_n7874 = new_n7871 & new_n7872;
  assign new_n7875 = ~new_n7873 & ~new_n7874;
  assign new_n7876 = ~new_n7870 & ~new_n7875;
  assign new_n7877 = new_n7870 & new_n7875;
  assign new_n7878 = ~new_n7876 & ~new_n7877;
  assign new_n7879 = new_n7755 & ~new_n7758;
  assign new_n7880 = ~new_n7759 & ~new_n7879;
  assign new_n7881 = ~new_n7878 & new_n7880;
  assign new_n7882 = new_n7878 & ~new_n7880;
  assign new_n7883 = ~new_n7881 & ~new_n7882;
  assign new_n7884 = new_n7869 & new_n7883;
  assign new_n7885 = ~new_n7869 & ~new_n7883;
  assign new_n7886 = ~new_n7884 & ~new_n7885;
  assign new_n7887 = ~new_n7765 & ~new_n7768;
  assign new_n7888 = ~new_n7764 & ~new_n7887;
  assign new_n7889 = new_n7886 & ~new_n7888;
  assign new_n7890 = ~new_n7886 & new_n7888;
  assign new_n7891_1 = ~new_n7889 & ~new_n7890;
  assign new_n7892 = ~new_n7773 & ~new_n7776;
  assign new_n7893 = ~new_n7772 & ~new_n7892;
  assign new_n7894 = new_n7891_1 & ~new_n7893;
  assign new_n7895 = ~new_n7891_1 & new_n7893;
  assign new_n7896 = ~new_n7894 & ~new_n7895;
  assign new_n7897 = new_n7864 & new_n7896;
  assign new_n7898 = ~new_n7864 & ~new_n7896;
  assign new_n7899 = ~new_n7897 & ~new_n7898;
  assign new_n7900 = new_n7780 & new_n7899;
  assign new_n7901 = ~new_n7780 & ~new_n7899;
  assign new_n7902 = ~new_n7900 & ~new_n7901;
  assign new_n7903 = ~new_n7786 & new_n7852;
  assign new_n7904 = ~new_n7785 & ~new_n7903;
  assign new_n7905 = new_n7902 & ~new_n7904;
  assign new_n7906 = ~new_n7902 & new_n7904;
  assign new_n7907 = ~new_n7905 & ~new_n7906;
  assign new_n7908 = n5153 & n7236;
  assign new_n7909 = ~new_n7820 & ~new_n7840;
  assign new_n7910 = ~new_n7821 & ~new_n7909;
  assign new_n7911 = n3992 & n7270;
  assign new_n7912 = n806 & n8384;
  assign new_n7913 = new_n7911 & new_n7912;
  assign new_n7914 = ~new_n7911 & ~new_n7912;
  assign new_n7915 = ~new_n7913 & ~new_n7914;
  assign new_n7916 = n3342 & n6358;
  assign new_n7917 = n5198 & n9111;
  assign new_n7918 = n1471 & n9763;
  assign new_n7919 = ~new_n7917 & ~new_n7918;
  assign new_n7920 = new_n7917 & new_n7918;
  assign new_n7921 = ~new_n7919 & ~new_n7920;
  assign new_n7922 = ~new_n7916 & ~new_n7921;
  assign new_n7923 = new_n7916 & new_n7921;
  assign new_n7924 = ~new_n7922 & ~new_n7923;
  assign new_n7925 = new_n7829 & ~new_n7831;
  assign new_n7926 = ~new_n7833 & ~new_n7925;
  assign new_n7927 = ~new_n7924 & new_n7926;
  assign new_n7928 = new_n7924 & ~new_n7926;
  assign new_n7929 = ~new_n7927 & ~new_n7928;
  assign new_n7930 = ~new_n7915 & ~new_n7929;
  assign new_n7931 = new_n7915 & new_n7929;
  assign new_n7932 = ~new_n7930 & ~new_n7931;
  assign new_n7933 = ~new_n7826 & ~new_n7837;
  assign new_n7934 = ~new_n7827 & ~new_n7933;
  assign new_n7935 = ~new_n7932 & new_n7934;
  assign new_n7936 = new_n7932 & ~new_n7934;
  assign new_n7937 = ~new_n7935 & ~new_n7936;
  assign new_n7938 = new_n7910 & ~new_n7937;
  assign new_n7939 = ~new_n7910 & new_n7937;
  assign new_n7940 = ~new_n7938 & ~new_n7939;
  assign new_n7941 = new_n7908 & new_n7940;
  assign new_n7942 = ~new_n7908 & ~new_n7940;
  assign new_n7943 = ~new_n7941 & ~new_n7942;
  assign new_n7944 = new_n7844 & new_n7943;
  assign new_n7945 = ~new_n7844 & ~new_n7943;
  assign new_n7946_1 = ~new_n7944 & ~new_n7945;
  assign new_n7947 = n4805 & n5798;
  assign new_n7948 = ~new_n7792 & ~new_n7810;
  assign new_n7949 = ~new_n7791 & ~new_n7948;
  assign new_n7950 = n6016 & n11478;
  assign new_n7951 = n521 & n5283;
  assign new_n7952 = ~new_n7950 & ~new_n7951;
  assign new_n7953 = new_n7950 & new_n7951;
  assign new_n7954 = ~new_n7952 & ~new_n7953;
  assign new_n7955 = n137 & n5579;
  assign new_n7956 = n2558 & n6797;
  assign new_n7957 = n2498 & n6294;
  assign new_n7958 = ~new_n7956 & ~new_n7957;
  assign new_n7959 = new_n7956 & new_n7957;
  assign new_n7960 = ~new_n7958 & ~new_n7959;
  assign new_n7961 = ~new_n7955 & ~new_n7960;
  assign new_n7962 = new_n7794 & ~new_n7796;
  assign new_n7963 = ~new_n7797 & ~new_n7962;
  assign new_n7964 = new_n7961 & new_n7963;
  assign new_n7965_1 = new_n7955 & new_n7960;
  assign new_n7966_1 = new_n7963 & ~new_n7965_1;
  assign new_n7967 = ~new_n7961 & ~new_n7966_1;
  assign new_n7968 = ~new_n7964 & ~new_n7967;
  assign new_n7969 = ~new_n7963 & new_n7965_1;
  assign new_n7970 = ~new_n7968 & ~new_n7969;
  assign new_n7971 = ~new_n7954 & new_n7970;
  assign new_n7972 = new_n7954 & ~new_n7970;
  assign new_n7973 = ~new_n7971 & ~new_n7972;
  assign new_n7974 = new_n7801 & ~new_n7805;
  assign new_n7975 = ~new_n7806 & ~new_n7974;
  assign new_n7976 = ~new_n7973 & ~new_n7975;
  assign new_n7977 = new_n7973 & new_n7975;
  assign new_n7978 = ~new_n7976 & ~new_n7977;
  assign new_n7979 = ~new_n7949 & new_n7978;
  assign new_n7980 = new_n7949 & ~new_n7978;
  assign new_n7981_1 = ~new_n7979 & ~new_n7980;
  assign new_n7982 = new_n7947 & new_n7981_1;
  assign new_n7983 = ~new_n7947 & ~new_n7981_1;
  assign new_n7984 = ~new_n7982 & ~new_n7983;
  assign new_n7985 = new_n7814 & new_n7984;
  assign new_n7986 = ~new_n7814 & ~new_n7984;
  assign new_n7987 = ~new_n7985 & ~new_n7986;
  assign new_n7988 = ~new_n7946_1 & ~new_n7987;
  assign new_n7989 = new_n7946_1 & new_n7987;
  assign new_n7990 = ~new_n7988 & ~new_n7989;
  assign new_n7991 = new_n7006 & ~new_n7847;
  assign new_n7992 = ~new_n7848 & ~new_n7991;
  assign new_n7993 = new_n7990 & new_n7992;
  assign new_n7994 = ~new_n7990 & ~new_n7992;
  assign new_n7995 = ~new_n7993 & ~new_n7994;
  assign new_n7996 = new_n7907 & ~new_n7995;
  assign new_n7997 = ~new_n7907 & new_n7995;
  assign new_n7998 = ~new_n7996 & ~new_n7997;
  assign new_n7999 = ~new_n7863 & new_n7998;
  assign new_n8000 = ~new_n7862_1 & ~new_n7999;
  assign new_n8001 = new_n7748 & ~new_n8000;
  assign new_n8002 = ~new_n7748 & new_n8000;
  assign new_n8003 = ~new_n7885 & ~new_n7888;
  assign new_n8004 = new_n7868 & new_n8003;
  assign new_n8005 = ~new_n7868 & ~new_n8003;
  assign new_n8006 = ~new_n7884 & new_n8005;
  assign new_n8007 = ~new_n8004 & ~new_n8006;
  assign new_n8008 = n9400 & n12221;
  assign new_n8009 = n2464 & n12145;
  assign new_n8010 = n6877 & n10217;
  assign new_n8011 = ~new_n8009 & ~new_n8010;
  assign new_n8012 = new_n8009 & new_n8010;
  assign new_n8013 = ~new_n8011 & ~new_n8012;
  assign new_n8014 = ~new_n8008 & ~new_n8013;
  assign new_n8015 = new_n8008 & new_n8013;
  assign new_n8016 = ~new_n8014 & ~new_n8015;
  assign new_n8017 = ~new_n7877 & new_n7880;
  assign new_n8018 = ~new_n7876 & ~new_n8017;
  assign new_n8019 = ~new_n8016 & ~new_n8018;
  assign new_n8020 = n2522 & n11311;
  assign new_n8021 = ~new_n7874 & ~new_n8020;
  assign new_n8022 = new_n7874 & new_n8020;
  assign new_n8023 = ~new_n8021 & ~new_n8022;
  assign new_n8024 = n7946 & n12753;
  assign new_n8025 = n2024 & n4203;
  assign new_n8026 = n4187 & n9189;
  assign new_n8027 = ~new_n8025 & ~new_n8026;
  assign new_n8028_1 = new_n8025 & new_n8026;
  assign new_n8029 = ~new_n8027 & ~new_n8028_1;
  assign new_n8030 = new_n8024 & ~new_n8029;
  assign new_n8031 = ~new_n8024 & new_n8029;
  assign new_n8032 = ~new_n8030 & ~new_n8031;
  assign new_n8033 = new_n8023 & new_n8032;
  assign new_n8034 = ~new_n8023 & ~new_n8032;
  assign new_n8035 = ~new_n8033 & ~new_n8034;
  assign new_n8036 = new_n8019 & new_n8035;
  assign new_n8037 = new_n8016 & new_n8018;
  assign new_n8038 = ~new_n8035 & new_n8037;
  assign new_n8039 = ~new_n8019 & ~new_n8035;
  assign new_n8040 = ~new_n8037 & ~new_n8039;
  assign new_n8041 = ~new_n8038 & ~new_n8040;
  assign new_n8042 = ~new_n8036 & ~new_n8041;
  assign new_n8043 = ~new_n8007 & new_n8042;
  assign new_n8044 = new_n8007 & ~new_n8042;
  assign new_n8045 = ~new_n8043 & ~new_n8044;
  assign new_n8046 = new_n7894 & ~new_n8045;
  assign new_n8047 = ~new_n7894 & new_n8045;
  assign new_n8048 = ~new_n8046 & ~new_n8047;
  assign new_n8049 = ~new_n7897 & ~new_n7900;
  assign new_n8050 = new_n8048 & ~new_n8049;
  assign new_n8051 = ~new_n8048 & new_n8049;
  assign new_n8052 = ~new_n8050 & ~new_n8051;
  assign new_n8053 = ~new_n7971 & new_n7975;
  assign new_n8054 = ~new_n7953 & ~new_n8053;
  assign new_n8055 = ~new_n7972 & new_n8054;
  assign new_n8056 = new_n7953 & new_n8053;
  assign new_n8057 = ~new_n8055 & ~new_n8056;
  assign new_n8058 = n2347 & n4805;
  assign new_n8059 = n5283 & n6016;
  assign new_n8060 = n5798 & n11478;
  assign new_n8061 = ~new_n8059 & ~new_n8060;
  assign new_n8062 = new_n8059 & new_n8060;
  assign new_n8063 = ~new_n8061 & ~new_n8062;
  assign new_n8064 = new_n8058 & ~new_n8063;
  assign new_n8065_1 = ~new_n8058 & new_n8063;
  assign new_n8066 = ~new_n8064 & ~new_n8065_1;
  assign new_n8067 = new_n7967 & ~new_n8066;
  assign new_n8068 = ~new_n7967 & new_n8066;
  assign new_n8069 = ~new_n8067 & ~new_n8068;
  assign new_n8070 = n137 & n521;
  assign new_n8071 = ~new_n7959 & ~new_n8070;
  assign new_n8072 = new_n7959 & new_n8070;
  assign new_n8073 = ~new_n8071 & ~new_n8072;
  assign new_n8074 = n2498 & n6797;
  assign new_n8075 = n2558 & n3146;
  assign new_n8076 = n5579 & n6294;
  assign new_n8077 = ~new_n8075 & ~new_n8076;
  assign new_n8078 = new_n8075 & new_n8076;
  assign new_n8079 = ~new_n8077 & ~new_n8078;
  assign new_n8080 = ~new_n8074 & ~new_n8079;
  assign new_n8081 = new_n8074 & new_n8079;
  assign new_n8082 = ~new_n8080 & ~new_n8081;
  assign new_n8083 = new_n8073 & ~new_n8082;
  assign new_n8084 = ~new_n8073 & new_n8082;
  assign new_n8085 = ~new_n8083 & ~new_n8084;
  assign new_n8086 = ~new_n8069 & ~new_n8085;
  assign new_n8087 = new_n8069 & new_n8085;
  assign new_n8088 = ~new_n8086 & ~new_n8087;
  assign new_n8089 = new_n8057 & ~new_n8088;
  assign new_n8090 = ~new_n8057 & new_n8088;
  assign new_n8091 = ~new_n8089 & ~new_n8090;
  assign new_n8092 = new_n7979 & new_n8091;
  assign new_n8093 = ~new_n7979 & ~new_n8091;
  assign new_n8094 = ~new_n8092 & ~new_n8093;
  assign new_n8095 = ~new_n7982 & ~new_n7985;
  assign new_n8096 = new_n8094 & ~new_n8095;
  assign new_n8097 = ~new_n8094 & new_n8095;
  assign new_n8098 = ~new_n8096 & ~new_n8097;
  assign new_n8099 = ~new_n7941 & ~new_n7944;
  assign new_n8100_1 = ~new_n7930 & new_n7934;
  assign new_n8101 = new_n7913 & new_n8100_1;
  assign new_n8102 = ~new_n7913 & ~new_n8100_1;
  assign new_n8103 = ~new_n7931 & new_n8102;
  assign new_n8104 = ~new_n8101 & ~new_n8103;
  assign new_n8105 = n3992 & n5153;
  assign new_n8106 = n7270 & n8384;
  assign new_n8107 = n2507 & n7236;
  assign new_n8108 = new_n8106 & new_n8107;
  assign new_n8109 = ~new_n8106 & ~new_n8107;
  assign new_n8110 = ~new_n8108 & ~new_n8109;
  assign new_n8111 = ~new_n8105 & ~new_n8110;
  assign new_n8112 = new_n8105 & new_n8110;
  assign new_n8113 = ~new_n8111 & ~new_n8112;
  assign new_n8114 = ~new_n7923 & new_n7926;
  assign new_n8115 = ~new_n7922 & ~new_n8114;
  assign new_n8116 = ~new_n8113 & ~new_n8115;
  assign new_n8117 = new_n8113 & new_n8115;
  assign new_n8118 = ~new_n8116 & ~new_n8117;
  assign new_n8119 = n806 & n6358;
  assign new_n8120 = ~new_n7920 & ~new_n8119;
  assign new_n8121 = new_n7920 & new_n8119;
  assign new_n8122 = ~new_n8120 & ~new_n8121;
  assign new_n8123 = n7646 & n9763;
  assign new_n8124 = n1471 & n9111;
  assign new_n8125 = ~new_n7832 & ~new_n8124;
  assign new_n8126 = new_n7832 & new_n8124;
  assign new_n8127 = ~new_n8125 & ~new_n8126;
  assign new_n8128 = new_n8123 & ~new_n8127;
  assign new_n8129 = ~new_n8123 & new_n8127;
  assign new_n8130 = ~new_n8128 & ~new_n8129;
  assign new_n8131 = ~new_n8122 & new_n8130;
  assign new_n8132 = new_n8122 & ~new_n8130;
  assign new_n8133 = ~new_n8131 & ~new_n8132;
  assign new_n8134 = new_n8118 & new_n8133;
  assign new_n8135 = ~new_n8118 & ~new_n8133;
  assign new_n8136 = ~new_n8134 & ~new_n8135;
  assign new_n8137 = new_n8104 & ~new_n8136;
  assign new_n8138_1 = ~new_n8104 & new_n8136;
  assign new_n8139 = ~new_n8137 & ~new_n8138_1;
  assign new_n8140 = new_n7938 & ~new_n8139;
  assign new_n8141 = ~new_n7938 & new_n8139;
  assign new_n8142 = ~new_n8140 & ~new_n8141;
  assign new_n8143 = ~new_n8099 & new_n8142;
  assign new_n8144 = new_n8099 & ~new_n8142;
  assign new_n8145 = ~new_n8143 & ~new_n8144;
  assign new_n8146 = ~new_n8098 & ~new_n8145;
  assign new_n8147 = new_n8098 & new_n8145;
  assign new_n8148 = ~new_n8146 & ~new_n8147;
  assign new_n8149 = ~new_n7988 & ~new_n7992;
  assign new_n8150 = ~new_n7989 & ~new_n8149;
  assign new_n8151 = ~new_n8148 & new_n8150;
  assign new_n8152 = new_n8148 & ~new_n8150;
  assign new_n8153 = ~new_n8151 & ~new_n8152;
  assign new_n8154 = new_n8052 & new_n8153;
  assign new_n8155 = ~new_n8052 & ~new_n8153;
  assign new_n8156 = ~new_n8154 & ~new_n8155;
  assign new_n8157 = ~new_n7906 & ~new_n7995;
  assign new_n8158 = ~new_n7905 & ~new_n8157;
  assign new_n8159 = ~new_n8156 & ~new_n8158;
  assign new_n8160 = new_n8156 & new_n8158;
  assign new_n8161 = ~new_n8159 & ~new_n8160;
  assign new_n8162 = ~new_n8002 & ~new_n8161;
  assign new_n8163 = ~new_n8001 & ~new_n8162;
  assign new_n8164 = ~new_n8092 & ~new_n8096;
  assign new_n8165 = ~new_n8116 & new_n8133;
  assign new_n8166 = ~new_n8117 & ~new_n8165;
  assign new_n8167 = n6358 & n7270;
  assign new_n8168 = n806 & n5198;
  assign new_n8169 = new_n8167 & ~new_n8168;
  assign new_n8170 = ~new_n8167 & new_n8168;
  assign new_n8171 = ~new_n8169 & ~new_n8170;
  assign new_n8172 = n2507 & n3992;
  assign new_n8173 = n5153 & n8384;
  assign new_n8174 = ~new_n8172 & ~new_n8173;
  assign new_n8175 = new_n8172 & new_n8173;
  assign new_n8176 = ~new_n8174 & ~new_n8175;
  assign new_n8177 = n1576 & n4805;
  assign new_n8178 = n2558 & n4938;
  assign new_n8179 = new_n8177 & new_n8178;
  assign new_n8180 = ~new_n8177 & ~new_n8178;
  assign new_n8181 = ~new_n8179 & ~new_n8180;
  assign new_n8182 = new_n8176 & ~new_n8181;
  assign new_n8183 = ~new_n8176 & new_n8181;
  assign new_n8184 = ~new_n8182 & ~new_n8183;
  assign new_n8185 = ~new_n8171 & new_n8184;
  assign new_n8186 = new_n8171 & ~new_n8184;
  assign new_n8187 = ~new_n8185 & ~new_n8186;
  assign new_n8188 = ~new_n8121 & new_n8130;
  assign new_n8189 = ~new_n8120 & ~new_n8188;
  assign new_n8190 = new_n8123 & ~new_n8125;
  assign new_n8191 = ~new_n8126 & ~new_n8190;
  assign new_n8192 = ~new_n8105 & ~new_n8108;
  assign new_n8193 = ~new_n8109 & ~new_n8192;
  assign new_n8194 = ~new_n8191 & new_n8193;
  assign new_n8195 = new_n8191 & ~new_n8193;
  assign new_n8196 = ~new_n8194 & ~new_n8195;
  assign new_n8197 = new_n8189 & new_n8196;
  assign new_n8198 = ~new_n8189 & ~new_n8196;
  assign new_n8199 = ~new_n8197 & ~new_n8198;
  assign new_n8200 = new_n8187 & new_n8199;
  assign new_n8201 = ~new_n8187 & ~new_n8199;
  assign new_n8202_1 = ~new_n8200 & ~new_n8201;
  assign new_n8203 = new_n8166 & ~new_n8202_1;
  assign new_n8204 = ~new_n8166 & new_n8202_1;
  assign new_n8205 = ~new_n8203 & ~new_n8204;
  assign new_n8206 = n137 & n6016;
  assign new_n8207 = n521 & n6294;
  assign new_n8208 = ~new_n8206 & ~new_n8207;
  assign new_n8209 = new_n8206 & new_n8207;
  assign new_n8210 = ~new_n8208 & ~new_n8209;
  assign new_n8211 = n5579 & n6797;
  assign new_n8212 = n2498 & n3146;
  assign new_n8213 = new_n8211 & ~new_n8212;
  assign new_n8214 = ~new_n8211 & new_n8212;
  assign new_n8215 = ~new_n8213 & ~new_n8214;
  assign new_n8216 = ~new_n8210 & ~new_n8215;
  assign new_n8217 = new_n8210 & new_n8215;
  assign new_n8218 = ~new_n8216 & ~new_n8217;
  assign new_n8219 = ~new_n8205 & new_n8218;
  assign new_n8220 = new_n8205 & ~new_n8218;
  assign new_n8221 = ~new_n8219 & ~new_n8220;
  assign new_n8222 = ~new_n8055 & ~new_n8088;
  assign new_n8223 = ~new_n8056 & ~new_n8222;
  assign new_n8224 = n5283 & n5798;
  assign new_n8225 = ~new_n8068 & ~new_n8085;
  assign new_n8226 = ~new_n8067 & ~new_n8225;
  assign new_n8227 = new_n8224 & ~new_n8226;
  assign new_n8228 = ~new_n8224 & new_n8226;
  assign new_n8229 = ~new_n8227 & ~new_n8228;
  assign new_n8230 = new_n8223 & new_n8229;
  assign new_n8231 = ~new_n8223 & ~new_n8229;
  assign new_n8232 = ~new_n8230 & ~new_n8231;
  assign new_n8233 = new_n8221 & new_n8232;
  assign new_n8234 = ~new_n8221 & ~new_n8232;
  assign new_n8235 = ~new_n8233 & ~new_n8234;
  assign new_n8236_1 = ~new_n8072 & ~new_n8082;
  assign new_n8237 = ~new_n8071 & ~new_n8236_1;
  assign new_n8238 = n2347 & n11478;
  assign new_n8239 = ~new_n8074 & ~new_n8078;
  assign new_n8240 = ~new_n8077 & ~new_n8239;
  assign new_n8241 = ~new_n8238 & new_n8240;
  assign new_n8242 = new_n8238 & ~new_n8240;
  assign new_n8243 = ~new_n8241 & ~new_n8242;
  assign new_n8244 = new_n8058 & ~new_n8061;
  assign new_n8245 = ~new_n8062 & ~new_n8244;
  assign new_n8246 = ~new_n8243 & new_n8245;
  assign new_n8247 = new_n8243 & ~new_n8245;
  assign new_n8248 = ~new_n8246 & ~new_n8247;
  assign new_n8249 = new_n8237 & ~new_n8248;
  assign new_n8250 = ~new_n8237 & new_n8248;
  assign new_n8251 = ~new_n8249 & ~new_n8250;
  assign new_n8252 = ~new_n8235 & new_n8251;
  assign new_n8253 = new_n8235 & ~new_n8251;
  assign new_n8254 = ~new_n8252 & ~new_n8253;
  assign new_n8255 = new_n8164 & new_n8254;
  assign new_n8256 = ~new_n8164 & ~new_n8254;
  assign new_n8257 = ~new_n8255 & ~new_n8256;
  assign new_n8258 = n6826 & n7265;
  assign new_n8259 = ~new_n7731 & ~new_n7747;
  assign new_n8260 = ~new_n8258 & new_n8259;
  assign new_n8261 = new_n8258 & ~new_n8259;
  assign new_n8262 = ~new_n8260 & ~new_n8261;
  assign new_n8263 = new_n8257 & ~new_n8262;
  assign new_n8264 = ~new_n8257 & new_n8262;
  assign new_n8265 = ~new_n8263 & ~new_n8264;
  assign new_n8266 = ~new_n8163 & new_n8265;
  assign new_n8267 = new_n8163 & ~new_n8265;
  assign new_n8268 = ~new_n8266 & ~new_n8267;
  assign new_n8269 = ~new_n8006 & new_n8042;
  assign new_n8270 = ~new_n8004 & ~new_n8269;
  assign new_n8271 = n2512 & n7862;
  assign new_n8272 = new_n8270 & new_n8271;
  assign new_n8273 = ~new_n8270 & ~new_n8271;
  assign new_n8274 = ~new_n8272 & ~new_n8273;
  assign new_n8275 = new_n7725 & ~new_n8274;
  assign new_n8276_1 = ~new_n7725 & new_n8274;
  assign new_n8277 = ~new_n8275 & ~new_n8276_1;
  assign new_n8278 = ~new_n8147 & new_n8150;
  assign new_n8279 = ~new_n8146 & ~new_n8278;
  assign new_n8280 = ~new_n7703 & new_n7720;
  assign new_n8281 = ~new_n7702 & ~new_n8280;
  assign new_n8282 = ~new_n8279 & new_n8281;
  assign new_n8283 = new_n8279 & ~new_n8281;
  assign new_n8284 = ~new_n8282 & ~new_n8283;
  assign new_n8285 = ~new_n8140 & ~new_n8143;
  assign new_n8286 = n7646 & n9111;
  assign new_n8287 = n4722 & n9763;
  assign new_n8288 = ~new_n8286 & new_n8287;
  assign new_n8289 = new_n8286 & ~new_n8287;
  assign new_n8290 = ~new_n8288 & ~new_n8289;
  assign new_n8291 = n1471 & n3342;
  assign new_n8292 = n6431 & n7236;
  assign new_n8293 = ~new_n8291 & new_n8292;
  assign new_n8294 = new_n8291 & ~new_n8292;
  assign new_n8295 = ~new_n8293 & ~new_n8294;
  assign new_n8296 = ~new_n8290 & ~new_n8295;
  assign new_n8297 = new_n8290 & new_n8295;
  assign new_n8298 = ~new_n8296 & ~new_n8297;
  assign new_n8299 = ~new_n8008 & ~new_n8012;
  assign new_n8300 = ~new_n8011 & ~new_n8299;
  assign new_n8301 = ~new_n8298 & ~new_n8300;
  assign new_n8302 = new_n8298 & new_n8300;
  assign new_n8303_1 = ~new_n8301 & ~new_n8302;
  assign new_n8304 = ~new_n8103 & new_n8136;
  assign new_n8305 = ~new_n8101 & ~new_n8304;
  assign new_n8306 = n4203 & n9189;
  assign new_n8307 = n2522 & n4187;
  assign new_n8308 = ~new_n8306 & new_n8307;
  assign new_n8309 = new_n8306 & ~new_n8307;
  assign new_n8310 = ~new_n8308 & ~new_n8309;
  assign new_n8311 = n2464 & n12221;
  assign new_n8312 = n9400 & n10217;
  assign new_n8313 = ~new_n8311 & new_n8312;
  assign new_n8314 = new_n8311 & ~new_n8312;
  assign new_n8315 = ~new_n8313 & ~new_n8314;
  assign new_n8316 = new_n8310 & ~new_n8315;
  assign new_n8317 = ~new_n8310 & new_n8315;
  assign new_n8318 = ~new_n8316 & ~new_n8317;
  assign new_n8319 = ~new_n8022 & new_n8032;
  assign new_n8320 = ~new_n8021 & ~new_n8319;
  assign new_n8321 = ~new_n8318 & new_n8320;
  assign new_n8322 = new_n8318 & ~new_n8320;
  assign new_n8323 = ~new_n8321 & ~new_n8322;
  assign new_n8324 = n11311 & n12145;
  assign new_n8325 = new_n8024 & ~new_n8027;
  assign new_n8326 = ~new_n8028_1 & ~new_n8325;
  assign new_n8327 = ~new_n8324 & new_n8326;
  assign new_n8328 = new_n8324 & ~new_n8326;
  assign new_n8329 = ~new_n8327 & ~new_n8328;
  assign new_n8330 = ~new_n8040 & new_n8329;
  assign new_n8331 = new_n8040 & ~new_n8329;
  assign new_n8332 = ~new_n8330 & ~new_n8331;
  assign new_n8333 = new_n8323 & new_n8332;
  assign new_n8334 = ~new_n8323 & ~new_n8332;
  assign new_n8335 = ~new_n8333 & ~new_n8334;
  assign new_n8336_1 = new_n8305 & ~new_n8335;
  assign new_n8337 = ~new_n8305 & new_n8335;
  assign new_n8338 = ~new_n8336_1 & ~new_n8337;
  assign new_n8339 = ~new_n8303_1 & new_n8338;
  assign new_n8340 = new_n8303_1 & ~new_n8338;
  assign new_n8341 = ~new_n8339 & ~new_n8340;
  assign new_n8342 = new_n8285 & new_n8341;
  assign new_n8343 = ~new_n8285 & ~new_n8341;
  assign new_n8344 = ~new_n8342 & ~new_n8343;
  assign new_n8345 = ~new_n8046 & ~new_n8050;
  assign new_n8346 = ~new_n7691 & ~new_n7695;
  assign new_n8347 = ~new_n7694 & ~new_n8346;
  assign new_n8348 = ~new_n7706 & ~new_n7717;
  assign new_n8349 = ~new_n7707 & ~new_n8348;
  assign new_n8350 = ~new_n7709 & ~new_n7713;
  assign new_n8351 = ~new_n7712 & ~new_n8350;
  assign new_n8352 = n1333 & n3865;
  assign new_n8353 = n4634 & n5240;
  assign new_n8354 = ~new_n8352 & new_n8353;
  assign new_n8355 = new_n8352 & ~new_n8353;
  assign new_n8356 = ~new_n8354 & ~new_n8355;
  assign new_n8357 = new_n8351 & ~new_n8356;
  assign new_n8358 = ~new_n8351 & new_n8356;
  assign new_n8359 = ~new_n8357 & ~new_n8358;
  assign new_n8360 = n9195 & n11757;
  assign new_n8361 = n2253 & n3172;
  assign new_n8362 = new_n8360 & ~new_n8361;
  assign new_n8363 = ~new_n8360 & new_n8361;
  assign new_n8364 = ~new_n8362 & ~new_n8363;
  assign new_n8365 = n10223 & n11821;
  assign new_n8366 = n2879 & n9080;
  assign new_n8367 = new_n8365 & ~new_n8366;
  assign new_n8368 = ~new_n8365 & new_n8366;
  assign new_n8369 = ~new_n8367 & ~new_n8368;
  assign new_n8370 = ~new_n8364 & ~new_n8369;
  assign new_n8371 = new_n8364 & new_n8369;
  assign new_n8372 = ~new_n8370 & ~new_n8371;
  assign new_n8373 = ~new_n8359 & new_n8372;
  assign new_n8374 = new_n8359 & ~new_n8372;
  assign new_n8375 = ~new_n8373 & ~new_n8374;
  assign new_n8376 = new_n8349 & new_n8375;
  assign new_n8377 = ~new_n8349 & ~new_n8375;
  assign new_n8378 = ~new_n8376 & ~new_n8377;
  assign new_n8379 = ~new_n8347 & new_n8378;
  assign new_n8380 = new_n8347 & ~new_n8378;
  assign new_n8381 = ~new_n8379 & ~new_n8380;
  assign new_n8382 = n2024 & n12753;
  assign new_n8383 = n7946 & n10174;
  assign new_n8384_1 = n6877 & n7823;
  assign new_n8385 = new_n8383 & ~new_n8384_1;
  assign new_n8386 = ~new_n8383 & new_n8384_1;
  assign new_n8387 = ~new_n8385 & ~new_n8386;
  assign new_n8388 = new_n8382 & ~new_n8387;
  assign new_n8389 = ~new_n8382 & new_n8387;
  assign new_n8390 = ~new_n8388 & ~new_n8389;
  assign new_n8391 = ~new_n8381 & new_n8390;
  assign new_n8392 = new_n8381 & ~new_n8390;
  assign new_n8393 = ~new_n8391 & ~new_n8392;
  assign new_n8394 = new_n8345 & ~new_n8393;
  assign new_n8395 = ~new_n8345 & new_n8393;
  assign new_n8396 = ~new_n8394 & ~new_n8395;
  assign new_n8397 = new_n8344 & new_n8396;
  assign new_n8398_1 = ~new_n8344 & ~new_n8396;
  assign new_n8399 = ~new_n8397 & ~new_n8398_1;
  assign new_n8400 = new_n8284 & new_n8399;
  assign new_n8401 = ~new_n8284 & ~new_n8399;
  assign new_n8402 = ~new_n8400 & ~new_n8401;
  assign new_n8403 = ~new_n8155 & ~new_n8158;
  assign new_n8404 = ~new_n8154 & ~new_n8403;
  assign new_n8405 = ~new_n8402 & new_n8404;
  assign new_n8406 = new_n8402 & ~new_n8404;
  assign new_n8407 = ~new_n8405 & ~new_n8406;
  assign new_n8408 = ~new_n8277 & ~new_n8407;
  assign new_n8409 = new_n8277 & new_n8407;
  assign new_n8410 = ~new_n8408 & ~new_n8409;
  assign new_n8411 = ~new_n8268 & new_n8410;
  assign new_n8412 = new_n8268 & ~new_n8410;
  assign n2383 = new_n8411 | new_n8412;
  assign new_n8414 = ~new_n6661 & ~new_n6662;
  assign new_n8415 = new_n6672 & ~new_n8414;
  assign new_n8416 = ~new_n6672 & new_n8414;
  assign n2425 = ~new_n8415 & ~new_n8416;
  assign new_n8418 = ~new_n3273 & ~new_n3274;
  assign new_n8419 = new_n3328 & ~new_n8418;
  assign new_n8420 = ~new_n3328 & new_n8418;
  assign n2431 = ~new_n8419 & ~new_n8420;
  assign new_n8422 = ~new_n2304 & ~new_n2305;
  assign new_n8423 = new_n2327 & ~new_n8422;
  assign new_n8424 = ~new_n2327 & new_n8422;
  assign n2434 = ~new_n8423 & ~new_n8424;
  assign new_n8426 = ~new_n5663 & ~new_n5664;
  assign new_n8427 = ~new_n5668 & new_n8426;
  assign new_n8428 = new_n5668 & ~new_n8426;
  assign n2581 = ~new_n8427 & ~new_n8428;
  assign new_n8430 = ~new_n7611 & ~new_n7612;
  assign new_n8431 = new_n7624 & ~new_n8430;
  assign new_n8432 = ~new_n7624 & new_n8430;
  assign n2624 = ~new_n8431 & ~new_n8432;
  assign new_n8434 = ~new_n4588 & new_n4608;
  assign new_n8435 = ~new_n4589 & ~new_n8434;
  assign new_n8436 = n2564 & n2577;
  assign new_n8437 = n3842 & n4189;
  assign new_n8438 = ~new_n8436 & ~new_n8437;
  assign new_n8439 = new_n8436 & new_n8437;
  assign new_n8440 = ~new_n8438 & ~new_n8439;
  assign new_n8441 = n6770 & n11917;
  assign new_n8442 = n4921 & n9920;
  assign new_n8443 = n3627 & n9956;
  assign new_n8444 = ~new_n8442 & ~new_n8443;
  assign new_n8445 = new_n8442 & new_n8443;
  assign new_n8446 = ~new_n8444 & ~new_n8445;
  assign new_n8447 = ~new_n8441 & ~new_n8446;
  assign new_n8448 = new_n8441 & new_n8446;
  assign new_n8449 = ~new_n8447 & ~new_n8448;
  assign new_n8450 = new_n4597 & ~new_n4600;
  assign new_n8451 = ~new_n4601 & ~new_n8450;
  assign new_n8452 = ~new_n8449 & new_n8451;
  assign new_n8453 = new_n8449 & ~new_n8451;
  assign new_n8454 = ~new_n8452 & ~new_n8453;
  assign new_n8455 = new_n8440 & new_n8454;
  assign new_n8456 = ~new_n8440 & ~new_n8454;
  assign new_n8457 = ~new_n8455 & ~new_n8456;
  assign new_n8458 = ~new_n4595 & ~new_n4605;
  assign new_n8459 = ~new_n4594 & ~new_n8458;
  assign new_n8460 = new_n8457 & new_n8459;
  assign new_n8461 = ~new_n8457 & ~new_n8459;
  assign new_n8462 = ~new_n8460 & ~new_n8461;
  assign new_n8463 = new_n8435 & ~new_n8462;
  assign new_n8464 = ~new_n8456 & ~new_n8459;
  assign new_n8465 = ~new_n8439 & ~new_n8464;
  assign new_n8466 = ~new_n8455 & new_n8465;
  assign new_n8467 = new_n8439 & new_n8464;
  assign new_n8468 = ~new_n8466 & ~new_n8467;
  assign new_n8469 = n2564 & n9637;
  assign new_n8470 = n2577 & n4189;
  assign new_n8471 = n1835 & n6687;
  assign new_n8472 = ~new_n8470 & ~new_n8471;
  assign new_n8473 = new_n8470 & new_n8471;
  assign new_n8474 = ~new_n8472 & ~new_n8473;
  assign new_n8475 = ~new_n8469 & ~new_n8474;
  assign new_n8476_1 = new_n8469 & new_n8474;
  assign new_n8477 = ~new_n8475 & ~new_n8476_1;
  assign new_n8478 = ~new_n8447 & ~new_n8451;
  assign new_n8479 = ~new_n8448 & ~new_n8478;
  assign new_n8480 = ~new_n8477 & new_n8479;
  assign new_n8481 = new_n8477 & ~new_n8479;
  assign new_n8482 = ~new_n8480 & ~new_n8481;
  assign new_n8483 = n3842 & n6770;
  assign new_n8484 = new_n8445 & new_n8483;
  assign new_n8485 = ~new_n8445 & ~new_n8483;
  assign new_n8486 = ~new_n8484 & ~new_n8485;
  assign new_n8487 = n3627 & n4921;
  assign new_n8488 = n9920 & n11917;
  assign new_n8489 = n4516 & n9956;
  assign new_n8490 = new_n8488 & new_n8489;
  assign new_n8491 = ~new_n8488 & ~new_n8489;
  assign new_n8492 = ~new_n8490 & ~new_n8491;
  assign new_n8493 = ~new_n8487 & ~new_n8492;
  assign new_n8494 = new_n8487 & new_n8492;
  assign new_n8495 = ~new_n8493 & ~new_n8494;
  assign new_n8496 = new_n8486 & ~new_n8495;
  assign new_n8497 = ~new_n8486 & new_n8495;
  assign new_n8498 = ~new_n8496 & ~new_n8497;
  assign new_n8499 = ~new_n8482 & ~new_n8498;
  assign new_n8500 = new_n8482 & new_n8498;
  assign new_n8501 = ~new_n8499 & ~new_n8500;
  assign new_n8502 = ~new_n8468 & new_n8501;
  assign new_n8503 = new_n8468 & ~new_n8501;
  assign new_n8504 = ~new_n8502 & ~new_n8503;
  assign new_n8505 = new_n8463 & new_n8504;
  assign new_n8506 = ~new_n8463 & ~new_n8504;
  assign new_n8507 = ~new_n8505 & ~new_n8506;
  assign new_n8508 = n6687 & n9637;
  assign new_n8509 = ~new_n8435 & new_n8462;
  assign new_n8510 = ~new_n8463 & ~new_n8509;
  assign new_n8511 = new_n8508 & new_n8510;
  assign new_n8512 = ~new_n8508 & ~new_n8510;
  assign new_n8513 = ~new_n8511 & ~new_n8512;
  assign new_n8514 = new_n4612 & new_n8513;
  assign new_n8515 = ~new_n8511 & ~new_n8514;
  assign new_n8516 = new_n8507 & ~new_n8515;
  assign new_n8517 = ~new_n8507 & new_n8515;
  assign new_n8518 = ~new_n8516 & ~new_n8517;
  assign new_n8519 = n8065 & n8336;
  assign new_n8520 = n10439 & n10928;
  assign new_n8521 = n6986 & n8595;
  assign new_n8522 = ~new_n8520 & ~new_n8521;
  assign new_n8523 = new_n8520 & new_n8521;
  assign new_n8524 = ~new_n8522 & ~new_n8523;
  assign new_n8525 = n2226 & n6126;
  assign new_n8526 = n1094 & n3602;
  assign new_n8527 = n3719 & n10678;
  assign new_n8528 = new_n8526 & new_n8527;
  assign new_n8529 = ~new_n8526 & ~new_n8527;
  assign new_n8530 = ~new_n8528 & ~new_n8529;
  assign new_n8531 = ~new_n8525 & ~new_n8530;
  assign new_n8532 = new_n8525 & new_n8530;
  assign new_n8533 = ~new_n8531 & ~new_n8532;
  assign new_n8534 = new_n4815 & ~new_n4818;
  assign new_n8535 = ~new_n4819 & ~new_n8534;
  assign new_n8536 = ~new_n8533 & new_n8535;
  assign new_n8537 = new_n8533 & ~new_n8535;
  assign new_n8538 = ~new_n8536 & ~new_n8537;
  assign new_n8539 = new_n8524 & new_n8538;
  assign new_n8540 = ~new_n8524 & ~new_n8538;
  assign new_n8541 = ~new_n8539 & ~new_n8540;
  assign new_n8542 = ~new_n4813 & ~new_n4823;
  assign new_n8543 = ~new_n4812 & ~new_n8542;
  assign new_n8544 = ~new_n8541 & new_n8543;
  assign new_n8545 = new_n8541 & ~new_n8543;
  assign new_n8546 = ~new_n8544 & ~new_n8545;
  assign new_n8547 = new_n4830 & new_n8546;
  assign new_n8548 = ~new_n4830 & ~new_n8546;
  assign new_n8549 = ~new_n8547 & ~new_n8548;
  assign new_n8550 = new_n8519 & new_n8549;
  assign new_n8551 = ~new_n8519 & ~new_n8549;
  assign new_n8552 = ~new_n8550 & ~new_n8551;
  assign new_n8553 = new_n4834 & new_n8552;
  assign new_n8554 = ~new_n8550 & ~new_n8553;
  assign new_n8555 = ~new_n8540 & ~new_n8543;
  assign new_n8556 = new_n8523 & new_n8555;
  assign new_n8557 = ~new_n8523 & ~new_n8555;
  assign new_n8558 = ~new_n8539 & new_n8557;
  assign new_n8559 = ~new_n8556 & ~new_n8558;
  assign new_n8560 = n8065 & n10928;
  assign new_n8561 = n6986 & n10439;
  assign new_n8562 = n8336 & n10391;
  assign new_n8563 = ~new_n8561 & ~new_n8562;
  assign new_n8564 = new_n8561 & new_n8562;
  assign new_n8565 = ~new_n8563 & ~new_n8564;
  assign new_n8566 = ~new_n8560 & ~new_n8565;
  assign new_n8567 = new_n8560 & new_n8565;
  assign new_n8568 = ~new_n8566 & ~new_n8567;
  assign new_n8569 = ~new_n8532 & new_n8535;
  assign new_n8570 = ~new_n8531 & ~new_n8569;
  assign new_n8571 = new_n8568 & new_n8570;
  assign new_n8572 = ~new_n8568 & ~new_n8570;
  assign new_n8573 = ~new_n8571 & ~new_n8572;
  assign new_n8574 = n2226 & n8595;
  assign new_n8575 = ~new_n8528 & ~new_n8574;
  assign new_n8576 = new_n8528 & new_n8574;
  assign new_n8577 = ~new_n8575 & ~new_n8576;
  assign new_n8578 = n3602 & n10678;
  assign new_n8579 = n1094 & n6126;
  assign new_n8580 = n3719 & n7320;
  assign new_n8581 = ~new_n8579 & ~new_n8580;
  assign new_n8582 = new_n8579 & new_n8580;
  assign new_n8583 = ~new_n8581 & ~new_n8582;
  assign new_n8584 = ~new_n8578 & ~new_n8583;
  assign new_n8585 = new_n8578 & new_n8583;
  assign new_n8586 = ~new_n8584 & ~new_n8585;
  assign new_n8587 = new_n8577 & ~new_n8586;
  assign new_n8588 = ~new_n8577 & new_n8586;
  assign new_n8589 = ~new_n8587 & ~new_n8588;
  assign new_n8590 = ~new_n8573 & ~new_n8589;
  assign new_n8591 = new_n8573 & new_n8589;
  assign new_n8592 = ~new_n8590 & ~new_n8591;
  assign new_n8593 = ~new_n8559 & new_n8592;
  assign new_n8594 = ~new_n8558 & ~new_n8592;
  assign new_n8595_1 = ~new_n8556 & new_n8594;
  assign new_n8596 = ~new_n8593 & ~new_n8595_1;
  assign new_n8597 = new_n8547 & new_n8596;
  assign new_n8598 = ~new_n8547 & ~new_n8596;
  assign new_n8599 = ~new_n8597 & ~new_n8598;
  assign new_n8600 = ~new_n8554 & new_n8599;
  assign new_n8601 = new_n8554 & ~new_n8599;
  assign new_n8602 = ~new_n8600 & ~new_n8601;
  assign new_n8603 = n4970 & n12391;
  assign new_n8604 = n7610 & n7891;
  assign new_n8605 = ~new_n8603 & ~new_n8604;
  assign new_n8606 = new_n8603 & new_n8604;
  assign new_n8607 = ~new_n8605 & ~new_n8606;
  assign new_n8608 = n4826 & n7160;
  assign new_n8609 = n4828 & n7733;
  assign new_n8610 = n2515 & n12925;
  assign new_n8611 = ~new_n8609 & ~new_n8610;
  assign new_n8612 = new_n8609 & new_n8610;
  assign new_n8613 = ~new_n8611 & ~new_n8612;
  assign new_n8614 = new_n8608 & new_n8613;
  assign new_n8615 = ~new_n8608 & ~new_n8613;
  assign new_n8616 = ~new_n8614 & ~new_n8615;
  assign new_n8617 = new_n4873 & ~new_n4876;
  assign new_n8618 = ~new_n4877 & ~new_n8617;
  assign new_n8619 = ~new_n8616 & ~new_n8618;
  assign new_n8620 = new_n8616 & new_n8618;
  assign new_n8621 = ~new_n8619 & ~new_n8620;
  assign new_n8622 = ~new_n8607 & new_n8621;
  assign new_n8623 = new_n8607 & ~new_n8621;
  assign new_n8624 = ~new_n8622 & ~new_n8623;
  assign new_n8625 = ~new_n4871 & ~new_n4881;
  assign new_n8626 = ~new_n4870 & ~new_n8625;
  assign new_n8627 = ~new_n8624 & new_n8626;
  assign new_n8628 = new_n8624 & ~new_n8626;
  assign new_n8629 = ~new_n8627 & ~new_n8628;
  assign new_n8630 = ~new_n4886 & ~new_n4889;
  assign new_n8631 = ~new_n4885 & ~new_n8630;
  assign new_n8632 = new_n8629 & ~new_n8631;
  assign new_n8633 = ~new_n8622 & ~new_n8626;
  assign new_n8634 = ~new_n8606 & ~new_n8633;
  assign new_n8635 = ~new_n8623 & new_n8634;
  assign new_n8636 = new_n8606 & new_n8633;
  assign new_n8637 = ~new_n8635 & ~new_n8636;
  assign new_n8638 = n503 & n12391;
  assign new_n8639 = n4970 & n7891;
  assign new_n8640 = n10965 & n12069;
  assign new_n8641 = ~new_n8639 & ~new_n8640;
  assign new_n8642 = new_n8639 & new_n8640;
  assign new_n8643 = ~new_n8641 & ~new_n8642;
  assign new_n8644 = ~new_n8638 & ~new_n8643;
  assign new_n8645 = new_n8638 & new_n8643;
  assign new_n8646 = ~new_n8644 & ~new_n8645;
  assign new_n8647 = ~new_n8615 & ~new_n8618;
  assign new_n8648 = ~new_n8614 & ~new_n8647;
  assign new_n8649 = new_n8646 & ~new_n8648;
  assign new_n8650 = ~new_n8646 & new_n8648;
  assign new_n8651 = ~new_n8649 & ~new_n8650;
  assign new_n8652 = n7160 & n7610;
  assign new_n8653 = ~new_n8612 & ~new_n8652;
  assign new_n8654 = new_n8612 & new_n8652;
  assign new_n8655 = ~new_n8653 & ~new_n8654;
  assign new_n8656 = n2515 & n7733;
  assign new_n8657 = n4826 & n4828;
  assign new_n8658 = n1199 & n12925;
  assign new_n8659 = ~new_n8657 & ~new_n8658;
  assign new_n8660 = new_n8657 & new_n8658;
  assign new_n8661 = ~new_n8659 & ~new_n8660;
  assign new_n8662 = ~new_n8656 & ~new_n8661;
  assign new_n8663 = new_n8656 & new_n8661;
  assign new_n8664 = ~new_n8662 & ~new_n8663;
  assign new_n8665_1 = new_n8655 & ~new_n8664;
  assign new_n8666 = ~new_n8655 & new_n8664;
  assign new_n8667 = ~new_n8665_1 & ~new_n8666;
  assign new_n8668 = ~new_n8651 & ~new_n8667;
  assign new_n8669 = new_n8651 & new_n8667;
  assign new_n8670 = ~new_n8668 & ~new_n8669;
  assign new_n8671 = ~new_n8637 & new_n8670;
  assign new_n8672 = new_n8637 & ~new_n8670;
  assign new_n8673 = ~new_n8671 & ~new_n8672;
  assign new_n8674 = new_n8632 & new_n8673;
  assign new_n8675 = ~new_n8632 & ~new_n8673;
  assign new_n8676 = ~new_n8674 & ~new_n8675;
  assign new_n8677 = n503 & n12069;
  assign new_n8678 = ~new_n8629 & new_n8631;
  assign new_n8679 = ~new_n8632 & ~new_n8678;
  assign new_n8680 = new_n8677 & new_n8679;
  assign new_n8681 = ~new_n8677 & ~new_n8679;
  assign new_n8682 = ~new_n8680 & ~new_n8681;
  assign new_n8683 = new_n4893 & new_n8682;
  assign new_n8684 = ~new_n8680 & ~new_n8683;
  assign new_n8685 = new_n8676 & ~new_n8684;
  assign new_n8686 = ~new_n8676 & new_n8684;
  assign new_n8687 = ~new_n8685 & ~new_n8686;
  assign new_n8688 = n6359 & n11222;
  assign new_n8689 = n6611 & n11153;
  assign new_n8690 = n217 & n5314;
  assign new_n8691 = new_n8689 & new_n8690;
  assign new_n8692 = ~new_n8689 & ~new_n8690;
  assign new_n8693 = ~new_n8691 & ~new_n8692;
  assign new_n8694 = n996 & n4086;
  assign new_n8695 = n405 & n5767;
  assign new_n8696 = n5319 & n8433;
  assign new_n8697 = ~new_n8695 & ~new_n8696;
  assign new_n8698 = new_n8695 & new_n8696;
  assign new_n8699 = ~new_n8697 & ~new_n8698;
  assign new_n8700 = ~new_n8694 & ~new_n8699;
  assign new_n8701 = new_n8694 & new_n8699;
  assign new_n8702 = ~new_n8700 & ~new_n8701;
  assign new_n8703 = new_n4839 & ~new_n4841;
  assign new_n8704 = ~new_n4842 & ~new_n8703;
  assign new_n8705 = ~new_n8702 & new_n8704;
  assign new_n8706 = new_n8702 & ~new_n8704;
  assign new_n8707 = ~new_n8705 & ~new_n8706;
  assign new_n8708 = ~new_n8693 & ~new_n8707;
  assign new_n8709 = new_n8693 & new_n8707;
  assign new_n8710 = ~new_n8708 & ~new_n8709;
  assign new_n8711 = ~new_n4847 & new_n4851;
  assign new_n8712 = ~new_n4848 & ~new_n8711;
  assign new_n8713 = ~new_n8710 & ~new_n8712;
  assign new_n8714 = new_n8710 & new_n8712;
  assign new_n8715 = ~new_n8713 & ~new_n8714;
  assign new_n8716 = ~new_n4856 & ~new_n4859;
  assign new_n8717_1 = ~new_n4855 & ~new_n8716;
  assign new_n8718 = new_n8715 & ~new_n8717_1;
  assign new_n8719 = ~new_n8715 & new_n8717_1;
  assign new_n8720 = ~new_n8718 & ~new_n8719;
  assign new_n8721 = new_n8688 & new_n8720;
  assign new_n8722 = ~new_n8688 & ~new_n8720;
  assign new_n8723 = ~new_n8721 & ~new_n8722;
  assign new_n8724 = new_n4864 & new_n8723;
  assign new_n8725 = ~new_n8721 & ~new_n8724;
  assign new_n8726 = ~new_n8708 & new_n8712;
  assign new_n8727 = new_n8691 & new_n8726;
  assign new_n8728 = ~new_n8691 & ~new_n8726;
  assign new_n8729 = ~new_n8709 & new_n8728;
  assign new_n8730 = ~new_n8727 & ~new_n8729;
  assign new_n8731 = n5314 & n6611;
  assign new_n8732 = n11222 & n11296;
  assign new_n8733 = n6359 & n11153;
  assign new_n8734 = ~new_n8732 & ~new_n8733;
  assign new_n8735 = new_n8732 & new_n8733;
  assign new_n8736 = ~new_n8734 & ~new_n8735;
  assign new_n8737 = new_n8731 & ~new_n8736;
  assign new_n8738 = ~new_n8731 & new_n8736;
  assign new_n8739 = ~new_n8737 & ~new_n8738;
  assign new_n8740 = ~new_n8701 & new_n8704;
  assign new_n8741 = ~new_n8700 & ~new_n8740;
  assign new_n8742 = new_n8739 & ~new_n8741;
  assign new_n8743 = ~new_n8739 & new_n8741;
  assign new_n8744 = ~new_n8742 & ~new_n8743;
  assign new_n8745 = n217 & n996;
  assign new_n8746 = ~new_n8698 & ~new_n8745;
  assign new_n8747 = new_n8698 & new_n8745;
  assign new_n8748 = n405 & n5319;
  assign new_n8749 = n8433 & n9457;
  assign new_n8750 = n4086 & n5767;
  assign new_n8751 = ~new_n8749 & ~new_n8750;
  assign new_n8752 = new_n8749 & new_n8750;
  assign new_n8753 = ~new_n8751 & ~new_n8752;
  assign new_n8754 = ~new_n8748 & ~new_n8753;
  assign new_n8755 = new_n8748 & new_n8753;
  assign new_n8756 = ~new_n8754 & ~new_n8755;
  assign new_n8757 = ~new_n8747 & ~new_n8756;
  assign new_n8758 = ~new_n8746 & new_n8757;
  assign new_n8759_1 = ~new_n8746 & ~new_n8747;
  assign new_n8760 = new_n8756 & ~new_n8759_1;
  assign new_n8761 = ~new_n8758 & ~new_n8760;
  assign new_n8762 = ~new_n8744 & new_n8761;
  assign new_n8763 = new_n8744 & ~new_n8761;
  assign new_n8764 = ~new_n8762 & ~new_n8763;
  assign new_n8765 = new_n8730 & ~new_n8764;
  assign new_n8766 = ~new_n8730 & new_n8764;
  assign new_n8767 = ~new_n8765 & ~new_n8766;
  assign new_n8768 = new_n8718 & ~new_n8767;
  assign new_n8769 = ~new_n8718 & new_n8767;
  assign new_n8770 = ~new_n8768 & ~new_n8769;
  assign new_n8771 = ~new_n8725 & new_n8770;
  assign new_n8772 = new_n8725 & ~new_n8770;
  assign new_n8773 = ~new_n8771 & ~new_n8772;
  assign new_n8774 = new_n8687 & new_n8773;
  assign new_n8775 = ~new_n8687 & ~new_n8773;
  assign new_n8776 = ~new_n8774 & ~new_n8775;
  assign new_n8777 = ~new_n4893 & ~new_n8682;
  assign new_n8778 = ~new_n8683 & ~new_n8777;
  assign new_n8779 = ~new_n4864 & ~new_n8723;
  assign new_n8780 = ~new_n8724 & ~new_n8779;
  assign new_n8781 = new_n8778 & new_n8780;
  assign new_n8782 = ~new_n8778 & ~new_n8780;
  assign new_n8783 = new_n4865 & ~new_n4899;
  assign new_n8784 = ~new_n4898 & ~new_n8783;
  assign new_n8785 = ~new_n8782 & ~new_n8784;
  assign new_n8786 = ~new_n8781 & ~new_n8785;
  assign new_n8787 = ~new_n8776 & ~new_n8786;
  assign new_n8788 = new_n8776 & new_n8786;
  assign new_n8789 = ~new_n8787 & ~new_n8788;
  assign new_n8790 = ~new_n8602 & new_n8789;
  assign new_n8791 = new_n8602 & ~new_n8789;
  assign new_n8792 = ~new_n8790 & ~new_n8791;
  assign new_n8793 = ~new_n4834 & ~new_n8552;
  assign new_n8794 = ~new_n8553 & ~new_n8793;
  assign new_n8795 = ~new_n8781 & ~new_n8782;
  assign new_n8796 = new_n8784 & ~new_n8795;
  assign new_n8797 = ~new_n8784 & new_n8795;
  assign new_n8798 = ~new_n8796 & ~new_n8797;
  assign new_n8799 = ~new_n8794 & ~new_n8798;
  assign new_n8800 = new_n8794 & new_n8798;
  assign new_n8801 = ~new_n4904 & ~new_n4908;
  assign new_n8802 = ~new_n4905 & ~new_n8801;
  assign new_n8803 = ~new_n8800 & ~new_n8802;
  assign new_n8804 = ~new_n8799 & ~new_n8803;
  assign new_n8805 = ~new_n8792 & ~new_n8804;
  assign new_n8806 = new_n8792 & new_n8804;
  assign new_n8807 = ~new_n8805 & ~new_n8806;
  assign new_n8808 = new_n8518 & new_n8807;
  assign new_n8809 = ~new_n8518 & ~new_n8807;
  assign new_n8810 = ~new_n4612 & ~new_n8513;
  assign new_n8811 = ~new_n8514 & ~new_n8810;
  assign new_n8812 = ~new_n4802 & ~new_n4911;
  assign new_n8813 = ~new_n4803 & ~new_n8812;
  assign new_n8814 = new_n8811 & ~new_n8813;
  assign new_n8815 = ~new_n8811 & new_n8813;
  assign new_n8816 = ~new_n8799 & ~new_n8800;
  assign new_n8817 = new_n8802 & ~new_n8816;
  assign new_n8818 = ~new_n8802 & new_n8816;
  assign new_n8819_1 = ~new_n8817 & ~new_n8818;
  assign new_n8820 = ~new_n8815 & ~new_n8819_1;
  assign new_n8821 = ~new_n8814 & ~new_n8820;
  assign new_n8822 = ~new_n8809 & ~new_n8821;
  assign new_n8823 = ~new_n8808 & ~new_n8822;
  assign new_n8824 = ~new_n8791 & ~new_n8804;
  assign new_n8825 = ~new_n8790 & ~new_n8824;
  assign new_n8826 = ~new_n8775 & ~new_n8786;
  assign new_n8827 = ~new_n8774 & ~new_n8826;
  assign new_n8828 = ~new_n8768 & ~new_n8771;
  assign new_n8829 = n4086 & n5319;
  assign new_n8830 = n405 & n9457;
  assign new_n8831 = ~new_n8829 & ~new_n8830;
  assign new_n8832 = new_n8829 & new_n8830;
  assign new_n8833 = ~new_n8831 & ~new_n8832;
  assign new_n8834 = n1357 & n11222;
  assign new_n8835 = n4817 & n8433;
  assign new_n8836 = new_n8834 & ~new_n8835;
  assign new_n8837 = ~new_n8834 & new_n8835;
  assign new_n8838 = ~new_n8836 & ~new_n8837;
  assign new_n8839 = ~new_n8833 & ~new_n8838;
  assign new_n8840 = new_n8833 & new_n8838;
  assign new_n8841 = ~new_n8839 & ~new_n8840;
  assign new_n8842 = ~new_n8560 & ~new_n8564;
  assign new_n8843 = ~new_n8563 & ~new_n8842;
  assign new_n8844 = ~new_n8841 & ~new_n8843;
  assign new_n8845 = new_n8841 & new_n8843;
  assign new_n8846 = ~new_n8844 & ~new_n8845;
  assign new_n8847 = ~new_n8729 & new_n8764;
  assign new_n8848 = ~new_n8727 & ~new_n8847;
  assign new_n8849 = n1094 & n8595;
  assign new_n8850 = n6126 & n10678;
  assign new_n8851 = ~new_n8849 & new_n8850;
  assign new_n8852 = new_n8849 & ~new_n8850;
  assign new_n8853 = ~new_n8851 & ~new_n8852;
  assign new_n8854 = n6986 & n8065;
  assign new_n8855 = n10391 & n10928;
  assign new_n8856 = ~new_n8854 & new_n8855;
  assign new_n8857 = new_n8854 & ~new_n8855;
  assign new_n8858 = ~new_n8856 & ~new_n8857;
  assign new_n8859 = ~new_n8853 & ~new_n8858;
  assign new_n8860 = new_n8853 & new_n8858;
  assign new_n8861 = ~new_n8859 & ~new_n8860;
  assign new_n8862 = ~new_n8572 & ~new_n8589;
  assign new_n8863 = ~new_n8571 & ~new_n8862;
  assign new_n8864 = n2226 & n10439;
  assign new_n8865 = ~new_n8578 & ~new_n8582;
  assign new_n8866 = ~new_n8581 & ~new_n8865;
  assign new_n8867 = ~new_n8864 & new_n8866;
  assign new_n8868 = new_n8864 & ~new_n8866;
  assign new_n8869 = ~new_n8867 & ~new_n8868;
  assign new_n8870 = ~new_n8576 & ~new_n8586;
  assign new_n8871 = ~new_n8575 & ~new_n8870;
  assign new_n8872 = ~new_n8869 & new_n8871;
  assign new_n8873 = new_n8869 & ~new_n8871;
  assign new_n8874 = ~new_n8872 & ~new_n8873;
  assign new_n8875 = ~new_n8863 & new_n8874;
  assign new_n8876 = new_n8863 & ~new_n8874;
  assign new_n8877 = ~new_n8875 & ~new_n8876;
  assign new_n8878 = new_n8861 & new_n8877;
  assign new_n8879 = ~new_n8861 & ~new_n8877;
  assign new_n8880 = ~new_n8878 & ~new_n8879;
  assign new_n8881 = new_n8848 & ~new_n8880;
  assign new_n8882 = ~new_n8848 & new_n8880;
  assign new_n8883 = ~new_n8881 & ~new_n8882;
  assign new_n8884 = ~new_n8846 & new_n8883;
  assign new_n8885 = new_n8846 & ~new_n8883;
  assign new_n8886 = ~new_n8884 & ~new_n8885;
  assign new_n8887 = new_n8828 & new_n8886;
  assign new_n8888 = ~new_n8828 & ~new_n8886;
  assign new_n8889 = ~new_n8887 & ~new_n8888;
  assign new_n8890 = ~new_n8597 & ~new_n8600;
  assign new_n8891 = n4189 & n9637;
  assign new_n8892 = ~new_n8484 & ~new_n8495;
  assign new_n8893 = ~new_n8485 & ~new_n8892;
  assign new_n8894 = new_n8891 & new_n8893;
  assign new_n8895 = ~new_n8891 & ~new_n8893;
  assign new_n8896 = ~new_n8894 & ~new_n8895;
  assign new_n8897 = ~new_n8481 & new_n8498;
  assign new_n8898 = ~new_n8480 & ~new_n8897;
  assign new_n8899 = ~new_n8896 & new_n8898;
  assign new_n8900 = new_n8896 & ~new_n8898;
  assign new_n8901 = ~new_n8899 & ~new_n8900;
  assign new_n8902 = n3627 & n11917;
  assign new_n8903 = n4516 & n4921;
  assign new_n8904 = ~new_n8902 & new_n8903;
  assign new_n8905 = new_n8902 & ~new_n8903;
  assign new_n8906 = ~new_n8904 & ~new_n8905;
  assign new_n8907 = n1835 & n2564;
  assign new_n8908 = n2577 & n6770;
  assign new_n8909 = n3842 & n9920;
  assign new_n8910 = new_n8908 & new_n8909;
  assign new_n8911 = ~new_n8908 & ~new_n8909;
  assign new_n8912 = ~new_n8910 & ~new_n8911;
  assign new_n8913 = new_n8907 & ~new_n8912;
  assign new_n8914 = ~new_n8907 & new_n8912;
  assign new_n8915 = ~new_n8913 & ~new_n8914;
  assign new_n8916 = ~new_n8906 & ~new_n8915;
  assign new_n8917 = new_n8906 & new_n8915;
  assign new_n8918 = ~new_n8916 & ~new_n8917;
  assign new_n8919 = ~new_n8487 & ~new_n8490;
  assign new_n8920 = ~new_n8491 & ~new_n8919;
  assign new_n8921 = ~new_n8469 & ~new_n8473;
  assign new_n8922 = ~new_n8472 & ~new_n8921;
  assign new_n8923 = ~new_n8920 & new_n8922;
  assign new_n8924 = new_n8920 & ~new_n8922;
  assign new_n8925 = ~new_n8923 & ~new_n8924;
  assign new_n8926 = ~new_n8918 & new_n8925;
  assign new_n8927 = new_n8918 & ~new_n8925;
  assign new_n8928 = ~new_n8926 & ~new_n8927;
  assign new_n8929 = n3602 & n7320;
  assign new_n8930 = n3719 & n7523;
  assign new_n8931 = n4190 & n8336;
  assign new_n8932 = ~new_n8930 & new_n8931;
  assign new_n8933 = new_n8930 & ~new_n8931;
  assign new_n8934 = ~new_n8932 & ~new_n8933;
  assign new_n8935 = new_n8929 & ~new_n8934;
  assign new_n8936 = ~new_n8929 & new_n8934;
  assign new_n8937 = ~new_n8935 & ~new_n8936;
  assign new_n8938 = ~new_n8928 & new_n8937;
  assign new_n8939 = new_n8928 & ~new_n8937;
  assign new_n8940 = ~new_n8938 & ~new_n8939;
  assign new_n8941 = ~new_n8901 & ~new_n8940;
  assign new_n8942 = new_n8901 & new_n8940;
  assign new_n8943 = ~new_n8941 & ~new_n8942;
  assign new_n8944 = ~new_n8556 & ~new_n8594;
  assign new_n8945 = ~new_n8943 & new_n8944;
  assign new_n8946 = new_n8943 & ~new_n8944;
  assign new_n8947 = ~new_n8945 & ~new_n8946;
  assign new_n8948 = ~new_n8890 & ~new_n8947;
  assign new_n8949 = new_n8890 & new_n8947;
  assign new_n8950 = ~new_n8948 & ~new_n8949;
  assign new_n8951 = ~new_n8889 & new_n8950;
  assign new_n8952 = new_n8889 & ~new_n8950;
  assign new_n8953 = ~new_n8951 & ~new_n8952;
  assign new_n8954 = ~new_n8827 & ~new_n8953;
  assign new_n8955 = new_n8827 & new_n8953;
  assign new_n8956 = ~new_n8954 & ~new_n8955;
  assign new_n8957 = ~new_n8649 & new_n8667;
  assign new_n8958 = ~new_n8650 & ~new_n8957;
  assign new_n8959 = n503 & n7891;
  assign new_n8960 = ~new_n8656 & ~new_n8660;
  assign new_n8961 = ~new_n8659 & ~new_n8960;
  assign new_n8962 = ~new_n8959 & new_n8961;
  assign new_n8963 = new_n8959 & ~new_n8961;
  assign new_n8964 = ~new_n8962 & ~new_n8963;
  assign new_n8965 = n10965 & n12391;
  assign new_n8966 = ~new_n8638 & ~new_n8642;
  assign new_n8967 = ~new_n8641 & ~new_n8966;
  assign new_n8968 = ~new_n8965 & new_n8967;
  assign new_n8969 = new_n8965 & ~new_n8967;
  assign new_n8970 = ~new_n8968 & ~new_n8969;
  assign new_n8971 = ~new_n8654 & ~new_n8664;
  assign new_n8972 = ~new_n8653 & ~new_n8971;
  assign new_n8973 = new_n8970 & new_n8972;
  assign new_n8974 = ~new_n8970 & ~new_n8972;
  assign new_n8975 = ~new_n8973 & ~new_n8974;
  assign new_n8976 = new_n8964 & ~new_n8975;
  assign new_n8977 = ~new_n8964 & new_n8975;
  assign new_n8978 = ~new_n8976 & ~new_n8977;
  assign new_n8979 = ~new_n8958 & ~new_n8978;
  assign new_n8980 = new_n8958 & new_n8978;
  assign new_n8981 = ~new_n8979 & ~new_n8980;
  assign new_n8982 = ~new_n8956 & new_n8981;
  assign new_n8983 = new_n8956 & ~new_n8981;
  assign new_n8984 = ~new_n8982 & ~new_n8983;
  assign new_n8985 = ~new_n8825 & ~new_n8984;
  assign new_n8986 = new_n8825 & new_n8984;
  assign new_n8987 = ~new_n8985 & ~new_n8986;
  assign new_n8988 = ~new_n8674 & ~new_n8685;
  assign new_n8989 = ~new_n8505 & ~new_n8516;
  assign new_n8990 = ~new_n8988 & new_n8989;
  assign new_n8991 = new_n8988 & ~new_n8989;
  assign new_n8992 = ~new_n8990 & ~new_n8991;
  assign new_n8993 = ~new_n8466 & ~new_n8501;
  assign new_n8994 = ~new_n8467 & ~new_n8993;
  assign new_n8995 = ~new_n8746 & ~new_n8757;
  assign new_n8996 = ~new_n8742 & ~new_n8761;
  assign new_n8997 = ~new_n8743 & ~new_n8996;
  assign new_n8998 = new_n8995 & new_n8997;
  assign new_n8999 = ~new_n8995 & ~new_n8997;
  assign new_n9000 = ~new_n8998 & ~new_n8999;
  assign new_n9001 = n4970 & n7160;
  assign new_n9002 = n4828 & n7610;
  assign new_n9003 = ~new_n9001 & ~new_n9002;
  assign new_n9004 = new_n9001 & new_n9002;
  assign new_n9005 = ~new_n9003 & ~new_n9004;
  assign new_n9006 = n2515 & n4826;
  assign new_n9007 = n1199 & n7733;
  assign new_n9008 = new_n9006 & ~new_n9007;
  assign new_n9009 = ~new_n9006 & new_n9007;
  assign new_n9010 = ~new_n9008 & ~new_n9009;
  assign new_n9011 = ~new_n9005 & ~new_n9010;
  assign new_n9012 = new_n9005 & new_n9010;
  assign new_n9013 = ~new_n9011 & ~new_n9012;
  assign new_n9014 = ~new_n9000 & new_n9013;
  assign new_n9015 = new_n9000 & ~new_n9013;
  assign new_n9016 = ~new_n9014 & ~new_n9015;
  assign new_n9017 = new_n8994 & new_n9016;
  assign new_n9018 = ~new_n8994 & ~new_n9016;
  assign new_n9019 = ~new_n9017 & ~new_n9018;
  assign new_n9020 = ~new_n8635 & ~new_n8670;
  assign new_n9021 = ~new_n8636 & ~new_n9020;
  assign new_n9022 = n11153 & n11296;
  assign new_n9023 = n996 & n6611;
  assign new_n9024 = n217 & n5767;
  assign new_n9025 = ~new_n9023 & new_n9024;
  assign new_n9026 = new_n9023 & ~new_n9024;
  assign new_n9027 = ~new_n9025 & ~new_n9026;
  assign new_n9028 = new_n9022 & new_n9027;
  assign new_n9029 = ~new_n9022 & ~new_n9027;
  assign new_n9030 = ~new_n9028 & ~new_n9029;
  assign new_n9031 = ~new_n8748 & ~new_n8752;
  assign new_n9032 = ~new_n8751 & ~new_n9031;
  assign new_n9033 = ~new_n9030 & new_n9032;
  assign new_n9034 = new_n9030 & ~new_n9032;
  assign new_n9035 = ~new_n9033 & ~new_n9034;
  assign new_n9036 = n5314 & n6359;
  assign new_n9037 = new_n8731 & ~new_n8734;
  assign new_n9038 = ~new_n8735 & ~new_n9037;
  assign new_n9039 = ~new_n9036 & new_n9038;
  assign new_n9040 = new_n9036 & ~new_n9038;
  assign new_n9041 = ~new_n9039 & ~new_n9040;
  assign new_n9042 = n7546 & n12069;
  assign new_n9043 = n6578 & n12925;
  assign new_n9044 = new_n9042 & new_n9043;
  assign new_n9045 = ~new_n9042 & ~new_n9043;
  assign new_n9046 = ~new_n9044 & ~new_n9045;
  assign new_n9047 = new_n9041 & ~new_n9046;
  assign new_n9048 = ~new_n9041 & new_n9046;
  assign new_n9049 = ~new_n9047 & ~new_n9048;
  assign new_n9050 = ~new_n9035 & new_n9049;
  assign new_n9051 = new_n9035 & ~new_n9049;
  assign new_n9052 = ~new_n9050 & ~new_n9051;
  assign new_n9053 = new_n9021 & new_n9052;
  assign new_n9054 = ~new_n9021 & ~new_n9052;
  assign new_n9055 = ~new_n9053 & ~new_n9054;
  assign new_n9056 = n6687 & n11536;
  assign new_n9057 = n2087 & n9956;
  assign new_n9058 = ~new_n9056 & new_n9057;
  assign new_n9059 = new_n9056 & ~new_n9057;
  assign new_n9060 = ~new_n9058 & ~new_n9059;
  assign new_n9061 = new_n9055 & new_n9060;
  assign new_n9062 = ~new_n9055 & ~new_n9060;
  assign new_n9063 = ~new_n9061 & ~new_n9062;
  assign new_n9064 = new_n9019 & ~new_n9063;
  assign new_n9065 = ~new_n9019 & new_n9063;
  assign new_n9066 = ~new_n9064 & ~new_n9065;
  assign new_n9067 = ~new_n8992 & ~new_n9066;
  assign new_n9068 = new_n8992 & new_n9066;
  assign new_n9069 = ~new_n9067 & ~new_n9068;
  assign new_n9070 = ~new_n8987 & new_n9069;
  assign new_n9071 = new_n8987 & ~new_n9069;
  assign new_n9072 = ~new_n9070 & ~new_n9071;
  assign new_n9073 = new_n8823 & ~new_n9072;
  assign new_n9074 = ~new_n8823 & new_n9072;
  assign n2679 = new_n9073 | new_n9074;
  assign new_n9076 = n2253 & n6687;
  assign new_n9077 = ~new_n6698 & ~new_n6701;
  assign new_n9078 = ~new_n6697 & ~new_n9077;
  assign new_n9079 = n2564 & n9195;
  assign new_n9080_1 = n4189 & n4634;
  assign new_n9081 = ~new_n9079 & ~new_n9080_1;
  assign new_n9082 = new_n9079 & new_n9080_1;
  assign new_n9083 = ~new_n9081 & ~new_n9082;
  assign new_n9084 = n6770 & n10223;
  assign new_n9085 = n2879 & n9920;
  assign new_n9086 = n3627 & n7265;
  assign new_n9087 = ~new_n9085 & ~new_n9086;
  assign new_n9088 = new_n9085 & new_n9086;
  assign new_n9089 = ~new_n9087 & ~new_n9088;
  assign new_n9090 = new_n9084 & new_n9089;
  assign new_n9091 = ~new_n9084 & ~new_n9089;
  assign new_n9092 = ~new_n9090 & ~new_n9091;
  assign new_n9093 = ~new_n6679 & ~new_n6684;
  assign new_n9094 = ~new_n6682 & ~new_n9093;
  assign new_n9095 = ~new_n9092 & new_n9094;
  assign new_n9096 = new_n9092 & ~new_n9094;
  assign new_n9097 = ~new_n9095 & ~new_n9096;
  assign new_n9098 = new_n9083 & ~new_n9097;
  assign new_n9099 = ~new_n9083 & new_n9097;
  assign new_n9100 = ~new_n9098 & ~new_n9099;
  assign new_n9101 = ~new_n6690 & ~new_n6693;
  assign new_n9102 = ~new_n6689_1 & ~new_n9101;
  assign new_n9103 = new_n9100 & new_n9102;
  assign new_n9104 = ~new_n9100 & ~new_n9102;
  assign new_n9105 = ~new_n9103 & ~new_n9104;
  assign new_n9106 = ~new_n9078 & ~new_n9105;
  assign new_n9107 = new_n9078 & new_n9105;
  assign new_n9108 = ~new_n9106 & ~new_n9107;
  assign new_n9109 = new_n9076 & new_n9108;
  assign new_n9110 = ~new_n9076 & ~new_n9108;
  assign new_n9111_1 = ~new_n9109 & ~new_n9110;
  assign new_n9112 = new_n6705 & new_n9111_1;
  assign new_n9113 = ~new_n6705 & ~new_n9111_1;
  assign new_n9114 = ~new_n9112 & ~new_n9113;
  assign new_n9115 = ~new_n6676 & ~new_n6814;
  assign new_n9116 = ~new_n6815 & ~new_n9115;
  assign new_n9117 = new_n9114 & ~new_n9116;
  assign new_n9118 = ~new_n9114 & new_n9116;
  assign new_n9119 = ~new_n9117 & ~new_n9118;
  assign new_n9120 = new_n6775 & ~new_n6809_1;
  assign new_n9121 = ~new_n6808 & ~new_n9120;
  assign new_n9122 = n8336 & n12221;
  assign new_n9123 = ~new_n6796 & new_n6799;
  assign new_n9124 = ~new_n6795 & ~new_n9123;
  assign new_n9125 = n10928 & n12145;
  assign new_n9126 = n2522 & n6986;
  assign new_n9127 = ~new_n9125 & ~new_n9126;
  assign new_n9128 = new_n9125 & new_n9126;
  assign new_n9129 = ~new_n9127 & ~new_n9128;
  assign new_n9130 = n2226 & n9189;
  assign new_n9131 = n1094 & n2024;
  assign new_n9132 = n7946 & n10678;
  assign new_n9133 = ~new_n9131 & ~new_n9132;
  assign new_n9134 = new_n9131 & new_n9132;
  assign new_n9135 = ~new_n9133 & ~new_n9134;
  assign new_n9136 = new_n9130 & new_n9135;
  assign new_n9137_1 = ~new_n9130 & ~new_n9135;
  assign new_n9138 = ~new_n9136 & ~new_n9137_1;
  assign new_n9139 = new_n6783 & ~new_n6786;
  assign new_n9140 = ~new_n6787 & ~new_n9139;
  assign new_n9141 = ~new_n9138 & ~new_n9140;
  assign new_n9142 = new_n9138 & new_n9140;
  assign new_n9143 = ~new_n9141 & ~new_n9142;
  assign new_n9144 = new_n9129 & ~new_n9143;
  assign new_n9145 = ~new_n9129 & new_n9143;
  assign new_n9146 = ~new_n9144 & ~new_n9145;
  assign new_n9147 = ~new_n6781 & ~new_n6791;
  assign new_n9148 = ~new_n6780 & ~new_n9147;
  assign new_n9149 = new_n9146 & new_n9148;
  assign new_n9150 = ~new_n9146 & ~new_n9148;
  assign new_n9151 = ~new_n9149 & ~new_n9150;
  assign new_n9152 = ~new_n9124 & ~new_n9151;
  assign new_n9153 = new_n9124 & new_n9151;
  assign new_n9154 = ~new_n9152 & ~new_n9153;
  assign new_n9155 = new_n9122 & new_n9154;
  assign new_n9156 = ~new_n9122 & ~new_n9154;
  assign new_n9157 = ~new_n9155 & ~new_n9156;
  assign new_n9158 = new_n6803 & new_n9157;
  assign new_n9159 = ~new_n6803 & ~new_n9157;
  assign new_n9160 = ~new_n9158 & ~new_n9159;
  assign new_n9161 = ~new_n9121 & ~new_n9160;
  assign new_n9162 = new_n9121 & new_n9160;
  assign new_n9163 = ~new_n9161 & ~new_n9162;
  assign new_n9164 = n5798 & n12069;
  assign new_n9165 = ~new_n6727 & new_n6731;
  assign new_n9166 = ~new_n6728 & ~new_n9165;
  assign new_n9167 = n6016 & n12391;
  assign new_n9168 = n521 & n7891;
  assign new_n9169 = ~new_n9167 & ~new_n9168;
  assign new_n9170 = new_n9167 & new_n9168;
  assign new_n9171 = ~new_n9169 & ~new_n9170;
  assign new_n9172 = n5579 & n7160;
  assign new_n9173 = new_n6709 & ~new_n6712;
  assign new_n9174 = ~new_n6558 & ~new_n9173;
  assign new_n9175 = new_n9172 & ~new_n9174;
  assign new_n9176 = ~new_n9172 & ~new_n9173;
  assign new_n9177 = ~new_n9175 & ~new_n9176;
  assign new_n9178 = n2498 & n4828;
  assign new_n9179 = n2515 & n2558;
  assign new_n9180 = ~new_n9178 & ~new_n9179;
  assign new_n9181 = new_n9178 & new_n9179;
  assign new_n9182 = ~new_n9180 & ~new_n9181;
  assign new_n9183 = new_n9177 & ~new_n9182;
  assign new_n9184 = ~new_n9177 & new_n9182;
  assign new_n9185 = ~new_n9183 & ~new_n9184;
  assign new_n9186 = new_n9171 & ~new_n9185;
  assign new_n9187 = ~new_n9171 & new_n9185;
  assign new_n9188 = ~new_n9186 & ~new_n9187;
  assign new_n9189_1 = ~new_n6717 & ~new_n6722;
  assign new_n9190 = ~new_n6721 & ~new_n9189_1;
  assign new_n9191 = new_n9188 & ~new_n9190;
  assign new_n9192 = ~new_n9188 & new_n9190;
  assign new_n9193 = ~new_n9191 & ~new_n9192;
  assign new_n9194 = new_n9166 & ~new_n9193;
  assign new_n9195_1 = ~new_n9166 & new_n9193;
  assign new_n9196 = ~new_n9194 & ~new_n9195_1;
  assign new_n9197 = new_n9164 & new_n9196;
  assign new_n9198 = ~new_n9164 & ~new_n9196;
  assign new_n9199 = ~new_n9197 & ~new_n9198;
  assign new_n9200 = new_n6735 & new_n9199;
  assign new_n9201 = ~new_n6735 & ~new_n9199;
  assign new_n9202 = ~new_n9200 & ~new_n9201;
  assign new_n9203 = n5153 & n11222;
  assign new_n9204 = ~new_n6758 & new_n6761;
  assign new_n9205 = ~new_n6757 & ~new_n9204;
  assign new_n9206 = n7270 & n11153;
  assign new_n9207 = n806 & n5314;
  assign new_n9208 = ~new_n9206 & ~new_n9207;
  assign new_n9209 = new_n9206 & new_n9207;
  assign new_n9210 = ~new_n9208 & ~new_n9209;
  assign new_n9211 = n996 & n3342;
  assign new_n9212 = n5767 & n9111;
  assign new_n9213 = n5319 & n9763;
  assign new_n9214 = ~new_n9212 & ~new_n9213;
  assign new_n9215 = new_n9212 & new_n9213;
  assign new_n9216 = ~new_n9214 & ~new_n9215;
  assign new_n9217 = new_n9211 & new_n9216;
  assign new_n9218 = ~new_n9211 & ~new_n9216;
  assign new_n9219 = ~new_n9217 & ~new_n9218;
  assign new_n9220 = ~new_n6745 & ~new_n6749;
  assign new_n9221 = ~new_n6748 & ~new_n9220;
  assign new_n9222 = ~new_n9219 & ~new_n9221;
  assign new_n9223 = new_n9219 & new_n9221;
  assign new_n9224 = ~new_n9222 & ~new_n9223;
  assign new_n9225 = new_n9210 & new_n9224;
  assign new_n9226 = ~new_n9210 & ~new_n9224;
  assign new_n9227 = ~new_n9225 & ~new_n9226;
  assign new_n9228 = ~new_n6742_1 & ~new_n6753;
  assign new_n9229 = ~new_n6743 & ~new_n9228;
  assign new_n9230 = new_n9227 & new_n9229;
  assign new_n9231 = ~new_n9227 & ~new_n9229;
  assign new_n9232 = ~new_n9230 & ~new_n9231;
  assign new_n9233 = ~new_n9205 & ~new_n9232;
  assign new_n9234 = new_n9205 & new_n9232;
  assign new_n9235 = ~new_n9233 & ~new_n9234;
  assign new_n9236 = new_n9203 & new_n9235;
  assign new_n9237 = ~new_n9203 & ~new_n9235;
  assign new_n9238 = ~new_n9236 & ~new_n9237;
  assign new_n9239 = new_n6765 & new_n9238;
  assign new_n9240 = ~new_n6765 & ~new_n9238;
  assign new_n9241_1 = ~new_n9239 & ~new_n9240;
  assign new_n9242 = new_n9202 & new_n9241_1;
  assign new_n9243 = ~new_n9202 & ~new_n9241_1;
  assign new_n9244 = ~new_n9242 & ~new_n9243;
  assign new_n9245 = ~new_n6769 & ~new_n6772;
  assign new_n9246 = ~new_n6768 & ~new_n9245;
  assign new_n9247 = ~new_n9244 & ~new_n9246;
  assign new_n9248 = new_n9244 & new_n9246;
  assign new_n9249 = ~new_n9247 & ~new_n9248;
  assign new_n9250 = new_n9163 & ~new_n9249;
  assign new_n9251 = ~new_n9163 & new_n9249;
  assign new_n9252 = ~new_n9250 & ~new_n9251;
  assign new_n9253 = new_n9119 & ~new_n9252;
  assign new_n9254 = ~new_n9119 & new_n9252;
  assign n2708 = new_n9253 | new_n9254;
  assign new_n9256 = ~new_n956 & ~new_n957;
  assign new_n9257 = ~new_n961 & ~new_n9256;
  assign new_n9258 = new_n961 & new_n9256;
  assign n2818 = ~new_n9257 & ~new_n9258;
  assign new_n9260 = ~new_n2296 & ~new_n2297;
  assign new_n9261 = new_n2329 & ~new_n9260;
  assign new_n9262 = ~new_n2329 & new_n9260;
  assign n2902 = ~new_n9261 & ~new_n9262;
  assign new_n9264 = n5305 & n11407;
  assign new_n9265 = n8759 & n12709;
  assign new_n9266 = n5331 & n12489;
  assign new_n9267 = n7965 & n10990;
  assign new_n9268 = new_n9266 & new_n9267;
  assign new_n9269 = ~new_n9266 & ~new_n9267;
  assign new_n9270 = ~new_n9268 & ~new_n9269;
  assign new_n9271 = new_n9265 & new_n9270;
  assign new_n9272 = ~new_n9265 & ~new_n9270;
  assign new_n9273 = ~new_n9271 & ~new_n9272;
  assign new_n9274 = new_n9264 & new_n9273;
  assign new_n9275 = ~new_n9264 & ~new_n9273;
  assign n3071 = ~new_n9274 & ~new_n9275;
  assign new_n9277 = ~new_n3297 & ~new_n3298;
  assign new_n9278 = new_n3322 & ~new_n9277;
  assign new_n9279 = ~new_n3322 & new_n9277;
  assign n3124 = ~new_n9278 & ~new_n9279;
  assign new_n9281 = n1097 & n11407;
  assign new_n9282 = n5305 & n11877;
  assign new_n9283 = ~new_n9281 & ~new_n9282;
  assign new_n9284 = n1097 & n11877;
  assign new_n9285 = new_n9264 & new_n9284;
  assign new_n9286 = ~new_n9283 & ~new_n9285;
  assign new_n9287 = n5212 & n5964;
  assign new_n9288 = ~new_n9264 & new_n9287;
  assign new_n9289 = ~new_n9286 & ~new_n9288;
  assign new_n9290 = ~new_n9283 & new_n9287;
  assign new_n9291 = ~new_n9264 & new_n9290;
  assign new_n9292 = ~new_n9289 & ~new_n9291;
  assign new_n9293 = n5964 & n11407;
  assign new_n9294 = n5212 & n5305;
  assign new_n9295 = ~new_n9293 & ~new_n9294;
  assign new_n9296 = new_n9293 & new_n9294;
  assign new_n9297 = ~new_n9295 & ~new_n9296;
  assign new_n9298 = new_n9274 & new_n9297;
  assign new_n9299 = ~new_n9274 & ~new_n9297;
  assign new_n9300 = n8759 & n11728;
  assign new_n9301 = n6776 & n12709;
  assign new_n9302 = ~new_n9300 & ~new_n9301;
  assign new_n9303 = new_n9300 & new_n9301;
  assign new_n9304 = ~new_n9302 & ~new_n9303;
  assign new_n9305 = new_n9271 & new_n9304;
  assign new_n9306 = ~new_n9271 & ~new_n9304;
  assign new_n9307 = ~new_n9305 & ~new_n9306;
  assign new_n9308 = n5760 & n7965;
  assign new_n9309 = n7388 & n10990;
  assign new_n9310 = ~new_n9308 & ~new_n9309;
  assign new_n9311 = new_n9308 & new_n9309;
  assign new_n9312 = ~new_n9310 & ~new_n9311;
  assign new_n9313 = n5331 & n7159;
  assign new_n9314 = n8476 & n12489;
  assign new_n9315 = ~new_n9313 & ~new_n9314;
  assign new_n9316 = new_n9313 & new_n9314;
  assign new_n9317 = ~new_n9315 & ~new_n9316;
  assign new_n9318 = new_n9268 & new_n9317;
  assign new_n9319 = ~new_n9268 & ~new_n9317;
  assign new_n9320 = ~new_n9318 & ~new_n9319;
  assign new_n9321 = new_n9312 & ~new_n9320;
  assign new_n9322 = ~new_n9312 & new_n9320;
  assign new_n9323 = ~new_n9321 & ~new_n9322;
  assign new_n9324 = new_n9307 & new_n9323;
  assign new_n9325 = ~new_n9307 & ~new_n9323;
  assign new_n9326 = ~new_n9324 & ~new_n9325;
  assign new_n9327 = ~new_n9299 & ~new_n9326;
  assign new_n9328 = ~new_n9298 & ~new_n9327;
  assign new_n9329 = new_n9292 & ~new_n9328;
  assign new_n9330 = ~new_n9292 & new_n9328;
  assign new_n9331 = ~new_n9329 & ~new_n9330;
  assign new_n9332 = ~new_n9305 & new_n9323;
  assign new_n9333 = ~new_n9306 & ~new_n9332;
  assign new_n9334 = n12299 & n12709;
  assign new_n9335 = n6429 & n8759;
  assign new_n9336 = ~new_n9334 & ~new_n9335;
  assign new_n9337 = n6776 & n11728;
  assign new_n9338 = ~new_n9265 & new_n9337;
  assign new_n9339 = ~new_n9336 & new_n9338;
  assign new_n9340 = n6429 & n12299;
  assign new_n9341 = new_n9265 & new_n9340;
  assign new_n9342 = ~new_n9336 & ~new_n9341;
  assign new_n9343 = ~new_n9338 & ~new_n9342;
  assign new_n9344 = ~new_n9339 & ~new_n9343;
  assign new_n9345 = new_n9333 & new_n9344;
  assign new_n9346 = ~new_n9333 & ~new_n9344;
  assign new_n9347 = ~new_n9345 & ~new_n9346;
  assign new_n9348 = n2530 & n12489;
  assign new_n9349 = n7159 & n8476;
  assign new_n9350 = n5331 & n12777;
  assign new_n9351 = ~new_n9349 & ~new_n9350;
  assign new_n9352 = new_n9349 & new_n9350;
  assign new_n9353 = ~new_n9351 & ~new_n9352;
  assign new_n9354 = new_n9348 & ~new_n9353;
  assign new_n9355 = ~new_n9348 & new_n9353;
  assign new_n9356 = ~new_n9354 & ~new_n9355;
  assign new_n9357 = new_n9316 & ~new_n9356;
  assign new_n9358 = ~new_n9316 & new_n9356;
  assign new_n9359 = ~new_n9357 & ~new_n9358;
  assign new_n9360 = n10990 & n11892;
  assign new_n9361 = n1478 & n7965;
  assign new_n9362 = ~new_n9360 & ~new_n9361;
  assign new_n9363 = n1478 & n11892;
  assign new_n9364 = new_n9267 & new_n9363;
  assign new_n9365 = ~new_n9362 & ~new_n9364;
  assign new_n9366 = n5760 & n7388;
  assign new_n9367 = ~new_n9267 & new_n9366;
  assign new_n9368 = ~new_n9365 & ~new_n9367;
  assign new_n9369 = ~new_n9362 & new_n9366;
  assign new_n9370 = ~new_n9267 & new_n9369;
  assign new_n9371 = ~new_n9368 & ~new_n9370;
  assign new_n9372 = new_n9359 & new_n9371;
  assign new_n9373 = ~new_n9359 & ~new_n9371;
  assign new_n9374 = ~new_n9372 & ~new_n9373;
  assign new_n9375 = ~new_n9312 & ~new_n9318;
  assign new_n9376 = ~new_n9319 & ~new_n9375;
  assign new_n9377 = ~new_n9374 & new_n9376;
  assign new_n9378 = new_n9374 & ~new_n9376;
  assign new_n9379 = ~new_n9377 & ~new_n9378;
  assign new_n9380 = new_n9347 & new_n9379;
  assign new_n9381 = ~new_n9347 & ~new_n9379;
  assign new_n9382 = ~new_n9380 & ~new_n9381;
  assign new_n9383 = new_n9331 & ~new_n9382;
  assign new_n9384 = ~new_n9331 & new_n9382;
  assign n3214 = ~new_n9383 & ~new_n9384;
  assign new_n9386 = ~new_n6294_1 & ~new_n6295;
  assign new_n9387_1 = ~new_n6297 & ~new_n9386;
  assign new_n9388 = ~new_n6294_1 & new_n6298;
  assign n3230 = new_n9387_1 | new_n9388;
  assign new_n9390 = ~new_n5629 & ~new_n5630;
  assign new_n9391 = new_n5684 & ~new_n9390;
  assign new_n9392 = ~new_n5684 & new_n9390;
  assign n3272 = new_n9391 | new_n9392;
  assign new_n9394 = n5320 & n5964;
  assign new_n9395 = n1097 & n4370;
  assign new_n9396 = ~new_n9394 & ~new_n9395;
  assign new_n9397 = new_n9394 & new_n9395;
  assign new_n9398 = ~new_n9396 & ~new_n9397;
  assign new_n9399 = n4370 & n5964;
  assign new_n9400_1 = n1097 & n5212;
  assign new_n9401 = n5964 & n11877;
  assign new_n9402 = new_n9400_1 & new_n9401;
  assign new_n9403 = ~new_n9400_1 & ~new_n9401;
  assign new_n9404 = n4312 & n11407;
  assign new_n9405 = ~new_n9403 & new_n9404;
  assign new_n9406 = ~new_n9402 & ~new_n9405;
  assign new_n9407 = ~new_n9399 & new_n9406;
  assign new_n9408 = new_n9399 & ~new_n9406;
  assign new_n9409 = n11407 & n12705;
  assign new_n9410 = n4312 & n5212;
  assign new_n9411 = ~new_n9284 & ~new_n9410;
  assign new_n9412 = new_n9284 & new_n9410;
  assign new_n9413 = ~new_n9411 & ~new_n9412;
  assign new_n9414 = new_n9409 & ~new_n9413;
  assign new_n9415 = ~new_n9409 & new_n9413;
  assign new_n9416 = ~new_n9414 & ~new_n9415;
  assign new_n9417 = ~new_n9408 & new_n9416;
  assign new_n9418 = ~new_n9407 & ~new_n9417;
  assign new_n9419 = new_n9398 & new_n9418;
  assign new_n9420 = ~new_n9398 & ~new_n9418;
  assign new_n9421 = ~new_n9419 & ~new_n9420;
  assign new_n9422 = n4312 & n11877;
  assign new_n9423 = n5212 & n12705;
  assign new_n9424 = n11407 & n12025;
  assign new_n9425 = new_n9423 & new_n9424;
  assign new_n9426 = ~new_n9423 & ~new_n9424;
  assign new_n9427 = ~new_n9425 & ~new_n9426;
  assign new_n9428 = ~new_n9422 & ~new_n9427;
  assign new_n9429 = new_n9422 & new_n9427;
  assign new_n9430 = ~new_n9428 & ~new_n9429;
  assign new_n9431 = new_n9409 & ~new_n9411;
  assign new_n9432 = ~new_n9412 & ~new_n9431;
  assign new_n9433 = ~new_n9430 & ~new_n9432;
  assign new_n9434 = new_n9430 & new_n9432;
  assign new_n9435 = ~new_n9433 & ~new_n9434;
  assign new_n9436 = ~new_n9421 & new_n9435;
  assign new_n9437 = new_n9421 & ~new_n9435;
  assign new_n9438 = ~new_n9436 & ~new_n9437;
  assign new_n9439 = n5305 & n5320;
  assign new_n9440 = ~new_n9407 & ~new_n9408;
  assign new_n9441 = ~new_n9416 & ~new_n9440;
  assign new_n9442 = new_n9416 & new_n9440;
  assign new_n9443 = ~new_n9441 & ~new_n9442;
  assign new_n9444 = new_n9439 & ~new_n9443;
  assign new_n9445 = ~new_n9439 & new_n9443;
  assign new_n9446 = n4370 & n5305;
  assign new_n9447 = ~new_n9285 & ~new_n9290;
  assign new_n9448 = ~new_n9446 & new_n9447;
  assign new_n9449 = new_n9446 & ~new_n9447;
  assign new_n9450 = ~new_n9402 & ~new_n9403;
  assign new_n9451 = ~new_n9404 & ~new_n9450;
  assign new_n9452 = new_n9404 & new_n9450;
  assign new_n9453 = ~new_n9451 & ~new_n9452;
  assign new_n9454 = ~new_n9449 & ~new_n9453;
  assign new_n9455 = ~new_n9448 & ~new_n9454;
  assign new_n9456 = ~new_n9445 & new_n9455;
  assign new_n9457_1 = ~new_n9444 & ~new_n9456;
  assign new_n9458 = new_n9438 & ~new_n9457_1;
  assign new_n9459 = n5212 & n12025;
  assign new_n9460 = n11877 & n12705;
  assign new_n9461 = n11257 & n11407;
  assign new_n9462 = ~new_n9460 & ~new_n9461;
  assign new_n9463 = new_n9460 & new_n9461;
  assign new_n9464 = ~new_n9462 & ~new_n9463;
  assign new_n9465 = ~new_n9459 & ~new_n9464;
  assign new_n9466 = new_n9459 & new_n9464;
  assign new_n9467 = ~new_n9465 & ~new_n9466;
  assign new_n9468 = n4312 & n4370;
  assign new_n9469 = new_n9425 & new_n9468;
  assign new_n9470 = ~new_n9425 & ~new_n9468;
  assign new_n9471 = ~new_n9469 & ~new_n9470;
  assign new_n9472 = new_n9467 & new_n9471;
  assign new_n9473 = ~new_n9467 & ~new_n9471;
  assign new_n9474 = ~new_n9472 & ~new_n9473;
  assign new_n9475 = n5964 & n12000;
  assign new_n9476 = n1097 & n5320;
  assign new_n9477 = n5305 & n9725;
  assign new_n9478 = ~new_n9476 & ~new_n9477;
  assign new_n9479 = new_n9476 & new_n9477;
  assign new_n9480 = ~new_n9478 & ~new_n9479;
  assign new_n9481 = ~new_n9475 & ~new_n9480;
  assign new_n9482 = new_n9475 & new_n9480;
  assign new_n9483 = ~new_n9481 & ~new_n9482;
  assign new_n9484 = ~new_n9429 & new_n9432;
  assign new_n9485 = ~new_n9428 & ~new_n9484;
  assign new_n9486 = ~new_n9483 & ~new_n9485;
  assign new_n9487 = new_n9483 & new_n9485;
  assign new_n9488 = ~new_n9486 & ~new_n9487;
  assign new_n9489 = ~new_n9474 & ~new_n9488;
  assign new_n9490 = new_n9474 & new_n9488;
  assign new_n9491 = ~new_n9489 & ~new_n9490;
  assign new_n9492 = ~new_n9420 & ~new_n9435;
  assign new_n9493 = ~new_n9397 & ~new_n9492;
  assign new_n9494 = ~new_n9419 & new_n9493;
  assign new_n9495 = new_n9397 & new_n9492;
  assign new_n9496 = ~new_n9494 & ~new_n9495;
  assign new_n9497 = ~new_n9491 & new_n9496;
  assign new_n9498 = new_n9491 & ~new_n9496;
  assign new_n9499 = ~new_n9497 & ~new_n9498;
  assign new_n9500 = new_n9458 & ~new_n9499;
  assign new_n9501 = ~new_n9458 & new_n9499;
  assign new_n9502 = ~new_n9500 & ~new_n9501;
  assign new_n9503 = n5305 & n12000;
  assign new_n9504 = ~new_n9438 & new_n9457_1;
  assign new_n9505 = ~new_n9458 & ~new_n9504;
  assign new_n9506 = new_n9503 & new_n9505;
  assign new_n9507 = ~new_n9286 & new_n9296;
  assign new_n9508 = ~new_n9448 & ~new_n9449;
  assign new_n9509 = new_n9453 & ~new_n9508;
  assign new_n9510 = ~new_n9453 & new_n9508;
  assign new_n9511 = ~new_n9509 & ~new_n9510;
  assign new_n9512 = new_n9507 & ~new_n9511;
  assign new_n9513 = ~new_n9444 & ~new_n9445;
  assign new_n9514 = ~new_n9455 & ~new_n9513;
  assign new_n9515 = new_n9455 & new_n9513;
  assign new_n9516 = ~new_n9514 & ~new_n9515;
  assign new_n9517 = new_n9512 & new_n9516;
  assign new_n9518 = ~new_n9503 & ~new_n9505;
  assign new_n9519 = ~new_n9506 & ~new_n9518;
  assign new_n9520 = new_n9517 & new_n9519;
  assign new_n9521 = ~new_n9506 & ~new_n9520;
  assign new_n9522 = new_n9502 & ~new_n9521;
  assign new_n9523 = ~new_n9502 & new_n9521;
  assign new_n9524 = ~new_n9522 & ~new_n9523;
  assign new_n9525 = n8717 & n8759;
  assign new_n9526 = n2433 & n8759;
  assign new_n9527 = n8276 & n12709;
  assign new_n9528 = n7436 & n11728;
  assign new_n9529 = ~new_n9340 & ~new_n9528;
  assign new_n9530 = new_n9340 & new_n9528;
  assign new_n9531 = ~new_n9529 & ~new_n9530;
  assign new_n9532 = new_n9527 & ~new_n9531;
  assign new_n9533 = ~new_n9527 & new_n9531;
  assign new_n9534 = ~new_n9532 & ~new_n9533;
  assign new_n9535 = n6776 & n8819;
  assign new_n9536 = n11728 & n12299;
  assign new_n9537 = n6429 & n6776;
  assign new_n9538 = new_n9536 & new_n9537;
  assign new_n9539 = ~new_n9536 & ~new_n9537;
  assign new_n9540 = n7436 & n12709;
  assign new_n9541 = ~new_n9539 & new_n9540;
  assign new_n9542 = ~new_n9538 & ~new_n9541;
  assign new_n9543 = new_n9535 & ~new_n9542;
  assign new_n9544 = ~new_n9535 & new_n9542;
  assign new_n9545 = ~new_n9543 & ~new_n9544;
  assign new_n9546 = ~new_n9534 & new_n9545;
  assign new_n9547 = new_n9534 & ~new_n9545;
  assign new_n9548 = ~new_n9546 & ~new_n9547;
  assign new_n9549 = ~new_n9526 & ~new_n9548;
  assign new_n9550 = new_n9526 & new_n9548;
  assign new_n9551 = n8759 & n8819;
  assign new_n9552 = ~new_n9337 & ~new_n9341;
  assign new_n9553 = ~new_n9336 & ~new_n9552;
  assign new_n9554 = new_n9551 & new_n9553;
  assign new_n9555 = ~new_n9551 & ~new_n9553;
  assign new_n9556 = ~new_n9538 & ~new_n9539;
  assign new_n9557 = ~new_n9540 & ~new_n9556;
  assign new_n9558 = new_n9540 & new_n9556;
  assign new_n9559 = ~new_n9557 & ~new_n9558;
  assign new_n9560 = ~new_n9555 & new_n9559;
  assign new_n9561 = ~new_n9554 & ~new_n9560;
  assign new_n9562 = ~new_n9550 & new_n9561;
  assign new_n9563 = ~new_n9549 & ~new_n9562;
  assign new_n9564 = n2433 & n6776;
  assign new_n9565 = n8819 & n12299;
  assign new_n9566 = new_n9564 & new_n9565;
  assign new_n9567 = ~new_n9564 & ~new_n9565;
  assign new_n9568 = ~new_n9566 & ~new_n9567;
  assign new_n9569 = n6429 & n7436;
  assign new_n9570 = n9241 & n12709;
  assign new_n9571_1 = n8276 & n11728;
  assign new_n9572 = new_n9570 & new_n9571_1;
  assign new_n9573 = ~new_n9570 & ~new_n9571_1;
  assign new_n9574 = ~new_n9572 & ~new_n9573;
  assign new_n9575 = ~new_n9569 & ~new_n9574;
  assign new_n9576 = new_n9569 & new_n9574;
  assign new_n9577 = ~new_n9575 & ~new_n9576;
  assign new_n9578_1 = new_n9527 & ~new_n9529;
  assign new_n9579 = ~new_n9530 & ~new_n9578_1;
  assign new_n9580 = ~new_n9577 & new_n9579;
  assign new_n9581 = new_n9577 & ~new_n9579;
  assign new_n9582 = ~new_n9580 & ~new_n9581;
  assign new_n9583_1 = ~new_n9568 & ~new_n9582;
  assign new_n9584 = new_n9568 & new_n9582;
  assign new_n9585 = ~new_n9583_1 & ~new_n9584;
  assign new_n9586 = new_n9534 & ~new_n9543;
  assign new_n9587 = ~new_n9544 & ~new_n9586;
  assign new_n9588 = ~new_n9585 & ~new_n9587;
  assign new_n9589 = new_n9585 & new_n9587;
  assign new_n9590 = ~new_n9588 & ~new_n9589;
  assign new_n9591 = new_n9563 & new_n9590;
  assign new_n9592 = ~new_n9563 & ~new_n9590;
  assign new_n9593 = ~new_n9591 & ~new_n9592;
  assign new_n9594 = new_n9525 & new_n9593;
  assign new_n9595 = new_n9303 & ~new_n9342;
  assign new_n9596 = ~new_n9554 & new_n9560;
  assign new_n9597 = ~new_n9554 & ~new_n9555;
  assign new_n9598 = ~new_n9559 & ~new_n9597;
  assign new_n9599 = ~new_n9596 & ~new_n9598;
  assign new_n9600 = new_n9595 & new_n9599;
  assign new_n9601 = ~new_n9549 & ~new_n9550;
  assign new_n9602 = ~new_n9561 & ~new_n9601;
  assign new_n9603 = new_n9561 & new_n9601;
  assign new_n9604 = ~new_n9602 & ~new_n9603;
  assign new_n9605 = new_n9600 & ~new_n9604;
  assign new_n9606 = ~new_n9525 & ~new_n9593;
  assign new_n9607 = ~new_n9594 & ~new_n9606;
  assign new_n9608 = new_n9605 & new_n9607;
  assign new_n9609 = ~new_n9594 & ~new_n9608;
  assign new_n9610 = ~new_n9575 & ~new_n9579;
  assign new_n9611 = ~new_n9576 & ~new_n9610;
  assign new_n9612 = n2433 & n12299;
  assign new_n9613 = n7730 & n8759;
  assign new_n9614 = n6776 & n8717;
  assign new_n9615 = ~new_n9613 & ~new_n9614;
  assign new_n9616 = new_n9613 & new_n9614;
  assign new_n9617 = ~new_n9615 & ~new_n9616;
  assign new_n9618 = new_n9612 & ~new_n9617;
  assign new_n9619 = ~new_n9612 & new_n9617;
  assign new_n9620 = ~new_n9618 & ~new_n9619;
  assign new_n9621 = ~new_n9611 & ~new_n9620;
  assign new_n9622 = new_n9611 & new_n9620;
  assign new_n9623 = ~new_n9621 & ~new_n9622;
  assign new_n9624 = n7436 & n8819;
  assign new_n9625 = ~new_n9572 & ~new_n9624;
  assign new_n9626 = new_n9572 & new_n9624;
  assign new_n9627 = ~new_n9625 & ~new_n9626;
  assign new_n9628 = n9241 & n11728;
  assign new_n9629 = n10510 & n12709;
  assign new_n9630 = n6429 & n8276;
  assign new_n9631 = ~new_n9629 & ~new_n9630;
  assign new_n9632 = new_n9629 & new_n9630;
  assign new_n9633 = ~new_n9631 & ~new_n9632;
  assign new_n9634 = ~new_n9628 & ~new_n9633;
  assign new_n9635 = new_n9628 & new_n9633;
  assign new_n9636 = ~new_n9634 & ~new_n9635;
  assign new_n9637_1 = ~new_n9627 & new_n9636;
  assign new_n9638 = ~new_n9626 & ~new_n9636;
  assign new_n9639 = ~new_n9625 & new_n9638;
  assign new_n9640_1 = ~new_n9637_1 & ~new_n9639;
  assign new_n9641 = ~new_n9623 & ~new_n9640_1;
  assign new_n9642 = new_n9623 & new_n9640_1;
  assign new_n9643 = ~new_n9641 & ~new_n9642;
  assign new_n9644 = ~new_n9583_1 & new_n9587;
  assign new_n9645 = new_n9566 & new_n9644;
  assign new_n9646 = ~new_n9566 & ~new_n9644;
  assign new_n9647 = ~new_n9584 & new_n9646;
  assign new_n9648 = ~new_n9645 & ~new_n9647;
  assign new_n9649 = new_n9643 & ~new_n9648;
  assign new_n9650 = ~new_n9643 & new_n9648;
  assign new_n9651 = ~new_n9649 & ~new_n9650;
  assign new_n9652 = new_n9591 & new_n9651;
  assign new_n9653 = ~new_n9591 & ~new_n9651;
  assign new_n9654 = ~new_n9652 & ~new_n9653;
  assign new_n9655 = ~new_n9609 & new_n9654;
  assign new_n9656 = new_n9609 & ~new_n9654;
  assign new_n9657 = ~new_n9655 & ~new_n9656;
  assign new_n9658 = n6441 & n7965;
  assign new_n9659 = n7965 & n12947;
  assign new_n9660 = n7965 & n11791;
  assign new_n9661 = ~new_n9364 & ~new_n9369;
  assign new_n9662 = new_n9660 & ~new_n9661;
  assign new_n9663 = ~new_n9660 & new_n9661;
  assign new_n9664 = n2393 & n10990;
  assign new_n9665 = n5760 & n11892;
  assign new_n9666 = n1478 & n7388;
  assign new_n9667 = ~new_n9665 & ~new_n9666;
  assign new_n9668 = new_n9665 & new_n9666;
  assign new_n9669 = ~new_n9667 & ~new_n9668;
  assign new_n9670 = new_n9664 & ~new_n9669;
  assign new_n9671 = ~new_n9664 & new_n9669;
  assign new_n9672 = ~new_n9670 & ~new_n9671;
  assign new_n9673 = ~new_n9663 & ~new_n9672;
  assign new_n9674 = ~new_n9662 & ~new_n9673;
  assign new_n9675 = new_n9659 & ~new_n9674;
  assign new_n9676 = ~new_n9659 & new_n9674;
  assign new_n9677 = n7388 & n11791;
  assign new_n9678 = new_n9664 & ~new_n9667;
  assign new_n9679 = ~new_n9668 & ~new_n9678;
  assign new_n9680 = ~new_n9677 & new_n9679;
  assign new_n9681 = new_n9677 & ~new_n9679;
  assign new_n9682 = ~new_n9680 & ~new_n9681;
  assign new_n9683 = n5860 & n10990;
  assign new_n9684 = n2393 & n5760;
  assign new_n9685 = ~new_n9363 & ~new_n9684;
  assign new_n9686 = new_n9363 & new_n9684;
  assign new_n9687 = ~new_n9685 & ~new_n9686;
  assign new_n9688 = new_n9683 & ~new_n9687;
  assign new_n9689 = ~new_n9683 & new_n9687;
  assign new_n9690 = ~new_n9688 & ~new_n9689;
  assign new_n9691 = ~new_n9682 & new_n9690;
  assign new_n9692 = new_n9682 & ~new_n9690;
  assign new_n9693 = ~new_n9691 & ~new_n9692;
  assign new_n9694 = ~new_n9676 & new_n9693;
  assign new_n9695 = ~new_n9675 & ~new_n9694;
  assign new_n9696 = n7388 & n12947;
  assign new_n9697 = n11791 & n11892;
  assign new_n9698 = new_n9696 & new_n9697;
  assign new_n9699 = ~new_n9696 & ~new_n9697;
  assign new_n9700 = ~new_n9698 & ~new_n9699;
  assign new_n9701 = n1478 & n2393;
  assign new_n9702 = n5760 & n5860;
  assign new_n9703 = n3986 & n10990;
  assign new_n9704 = ~new_n9702 & ~new_n9703;
  assign new_n9705 = new_n9702 & new_n9703;
  assign new_n9706_1 = ~new_n9704 & ~new_n9705;
  assign new_n9707 = ~new_n9701 & ~new_n9706_1;
  assign new_n9708 = new_n9701 & new_n9706_1;
  assign new_n9709 = ~new_n9707 & ~new_n9708;
  assign new_n9710 = new_n9683 & ~new_n9685;
  assign new_n9711 = ~new_n9686 & ~new_n9710;
  assign new_n9712 = ~new_n9709 & new_n9711;
  assign new_n9713 = new_n9709 & ~new_n9711;
  assign new_n9714 = ~new_n9712 & ~new_n9713;
  assign new_n9715 = ~new_n9700 & ~new_n9714;
  assign new_n9716 = new_n9700 & new_n9714;
  assign new_n9717 = ~new_n9715 & ~new_n9716;
  assign new_n9718 = ~new_n9680 & ~new_n9690;
  assign new_n9719 = ~new_n9681 & ~new_n9718;
  assign new_n9720 = ~new_n9717 & ~new_n9719;
  assign new_n9721 = new_n9717 & new_n9719;
  assign new_n9722 = ~new_n9720 & ~new_n9721;
  assign new_n9723 = ~new_n9695 & ~new_n9722;
  assign new_n9724 = new_n9695 & new_n9722;
  assign new_n9725_1 = ~new_n9723 & ~new_n9724;
  assign new_n9726 = new_n9658 & new_n9725_1;
  assign new_n9727 = new_n9311 & ~new_n9365;
  assign new_n9728 = ~new_n9662 & ~new_n9663;
  assign new_n9729 = new_n9672 & ~new_n9728;
  assign new_n9730 = ~new_n9672 & new_n9728;
  assign new_n9731 = ~new_n9729 & ~new_n9730;
  assign new_n9732 = new_n9727 & new_n9731;
  assign new_n9733 = ~new_n9675 & ~new_n9676;
  assign new_n9734 = ~new_n9693 & ~new_n9733;
  assign new_n9735 = new_n9693 & new_n9733;
  assign new_n9736 = ~new_n9734 & ~new_n9735;
  assign new_n9737 = new_n9732 & new_n9736;
  assign new_n9738 = ~new_n9658 & ~new_n9725_1;
  assign new_n9739 = ~new_n9726 & ~new_n9738;
  assign new_n9740 = new_n9737 & new_n9739;
  assign new_n9741 = ~new_n9726 & ~new_n9740;
  assign new_n9742 = ~new_n9715 & ~new_n9719;
  assign new_n9743 = new_n9698 & new_n9742;
  assign new_n9744 = ~new_n9698 & ~new_n9742;
  assign new_n9745 = ~new_n9716 & new_n9744;
  assign new_n9746 = ~new_n9743 & ~new_n9745;
  assign new_n9747 = ~new_n9708 & new_n9711;
  assign new_n9748 = ~new_n9707 & ~new_n9747;
  assign new_n9749 = n11892 & n12947;
  assign new_n9750 = n7965 & n11999;
  assign new_n9751 = n6441 & n7388;
  assign new_n9752 = ~new_n9750 & ~new_n9751;
  assign new_n9753 = new_n9750 & new_n9751;
  assign new_n9754 = ~new_n9752 & ~new_n9753;
  assign new_n9755 = new_n9749 & ~new_n9754;
  assign new_n9756_1 = ~new_n9749 & new_n9754;
  assign new_n9757 = ~new_n9755 & ~new_n9756_1;
  assign new_n9758 = ~new_n9748 & new_n9757;
  assign new_n9759 = new_n9748 & ~new_n9757;
  assign new_n9760 = ~new_n9758 & ~new_n9759;
  assign new_n9761 = n2393 & n11791;
  assign new_n9762 = ~new_n9705 & ~new_n9761;
  assign new_n9763_1 = new_n9705 & new_n9761;
  assign new_n9764 = ~new_n9762 & ~new_n9763_1;
  assign new_n9765 = n5857 & n10990;
  assign new_n9766 = n3986 & n5760;
  assign new_n9767_1 = n1478 & n5860;
  assign new_n9768 = ~new_n9766 & ~new_n9767_1;
  assign new_n9769 = new_n9766 & new_n9767_1;
  assign new_n9770 = ~new_n9768 & ~new_n9769;
  assign new_n9771 = new_n9765 & ~new_n9770;
  assign new_n9772 = ~new_n9765 & new_n9770;
  assign new_n9773 = ~new_n9771 & ~new_n9772;
  assign new_n9774 = ~new_n9764 & new_n9773;
  assign new_n9775 = new_n9764 & ~new_n9773;
  assign new_n9776 = ~new_n9774 & ~new_n9775;
  assign new_n9777 = new_n9760 & new_n9776;
  assign new_n9778 = ~new_n9760 & ~new_n9776;
  assign new_n9779 = ~new_n9777 & ~new_n9778;
  assign new_n9780 = new_n9746 & ~new_n9779;
  assign new_n9781 = ~new_n9746 & new_n9779;
  assign new_n9782 = ~new_n9780 & ~new_n9781;
  assign new_n9783 = new_n9723 & ~new_n9782;
  assign new_n9784 = ~new_n9723 & new_n9782;
  assign new_n9785 = ~new_n9783 & ~new_n9784;
  assign new_n9786 = ~new_n9741 & new_n9785;
  assign new_n9787 = new_n9741 & ~new_n9785;
  assign new_n9788 = ~new_n9786 & ~new_n9787;
  assign new_n9789 = n2530 & n6254;
  assign new_n9790 = n8476 & n11967;
  assign new_n9791 = ~new_n9789 & ~new_n9790;
  assign new_n9792 = new_n9789 & new_n9790;
  assign new_n9793 = ~new_n9791 & ~new_n9792;
  assign new_n9794 = n12648 & n12777;
  assign new_n9795 = n7159 & n10545;
  assign new_n9796 = n7690 & n12489;
  assign new_n9797 = ~new_n9795 & ~new_n9796;
  assign new_n9798 = new_n9795 & new_n9796;
  assign new_n9799 = ~new_n9797 & ~new_n9798;
  assign new_n9800 = new_n9794 & new_n9799;
  assign new_n9801 = ~new_n9794 & ~new_n9799;
  assign new_n9802 = ~new_n9800 & ~new_n9801;
  assign new_n9803 = n2530 & n12777;
  assign new_n9804 = n7159 & n12648;
  assign new_n9805 = new_n9803 & new_n9804;
  assign new_n9806 = n10545 & n12489;
  assign new_n9807 = ~new_n9803 & ~new_n9804;
  assign new_n9808 = new_n9806 & ~new_n9807;
  assign new_n9809 = ~new_n9805 & ~new_n9808;
  assign new_n9810 = ~new_n9802 & ~new_n9809;
  assign new_n9811 = new_n9802 & new_n9809;
  assign new_n9812 = ~new_n9810 & ~new_n9811;
  assign new_n9813 = ~new_n9793 & new_n9812;
  assign new_n9814 = new_n9793 & ~new_n9812;
  assign new_n9815 = ~new_n9813 & ~new_n9814;
  assign new_n9816 = n6254 & n8476;
  assign new_n9817 = n8476 & n12777;
  assign new_n9818 = n2530 & n7159;
  assign new_n9819 = new_n9817 & new_n9818;
  assign new_n9820_1 = ~new_n9817 & ~new_n9818;
  assign new_n9821 = n12489 & n12648;
  assign new_n9822 = ~new_n9820_1 & new_n9821;
  assign new_n9823 = ~new_n9819 & ~new_n9822;
  assign new_n9824 = ~new_n9816 & new_n9823;
  assign new_n9825 = new_n9816 & ~new_n9823;
  assign new_n9826 = ~new_n9805 & ~new_n9807;
  assign new_n9827 = ~new_n9806 & ~new_n9826;
  assign new_n9828 = new_n9806 & new_n9826;
  assign new_n9829 = ~new_n9827 & ~new_n9828;
  assign new_n9830 = ~new_n9825 & ~new_n9829;
  assign new_n9831 = ~new_n9824 & ~new_n9830;
  assign new_n9832 = new_n9815 & ~new_n9831;
  assign new_n9833 = ~new_n9815 & new_n9831;
  assign new_n9834 = ~new_n9832 & ~new_n9833;
  assign new_n9835 = n5331 & n11967;
  assign new_n9836 = ~new_n9824 & ~new_n9825;
  assign new_n9837 = new_n9829 & ~new_n9836;
  assign new_n9838 = ~new_n9829 & new_n9836;
  assign new_n9839 = ~new_n9837 & ~new_n9838;
  assign new_n9840 = new_n9835 & ~new_n9839;
  assign new_n9841 = ~new_n9835 & new_n9839;
  assign new_n9842 = n5331 & n6254;
  assign new_n9843 = ~new_n9348 & ~new_n9352;
  assign new_n9844 = ~new_n9351 & ~new_n9843;
  assign new_n9845 = new_n9842 & new_n9844;
  assign new_n9846 = ~new_n9842 & ~new_n9844;
  assign new_n9847 = ~new_n9819 & ~new_n9820_1;
  assign new_n9848 = ~new_n9821 & ~new_n9847;
  assign new_n9849 = new_n9821 & new_n9847;
  assign new_n9850 = ~new_n9848 & ~new_n9849;
  assign new_n9851 = ~new_n9846 & new_n9850;
  assign new_n9852 = ~new_n9845 & ~new_n9851;
  assign new_n9853 = ~new_n9841 & ~new_n9852;
  assign new_n9854 = ~new_n9840 & ~new_n9853;
  assign new_n9855 = ~new_n9834 & ~new_n9854;
  assign new_n9856 = ~new_n9813 & new_n9831;
  assign new_n9857 = ~new_n9792 & ~new_n9856;
  assign new_n9858 = ~new_n9814 & new_n9857;
  assign new_n9859 = new_n9792 & new_n9856;
  assign new_n9860 = ~new_n9858 & ~new_n9859;
  assign new_n9861 = ~new_n9800 & new_n9809;
  assign new_n9862 = ~new_n9801 & ~new_n9861;
  assign new_n9863 = n1353 & n5331;
  assign new_n9864 = n2530 & n11967;
  assign new_n9865 = n447 & n8476;
  assign new_n9866 = ~new_n9864 & ~new_n9865;
  assign new_n9867 = new_n9864 & new_n9865;
  assign new_n9868 = ~new_n9866 & ~new_n9867;
  assign new_n9869 = new_n9863 & ~new_n9868;
  assign new_n9870 = ~new_n9863 & new_n9868;
  assign new_n9871 = ~new_n9869 & ~new_n9870;
  assign new_n9872 = new_n9862 & ~new_n9871;
  assign new_n9873 = ~new_n9862 & new_n9871;
  assign new_n9874 = ~new_n9872 & ~new_n9873;
  assign new_n9875 = n6254 & n12648;
  assign new_n9876 = new_n9798 & new_n9875;
  assign new_n9877 = ~new_n9798 & ~new_n9875;
  assign new_n9878 = ~new_n9876 & ~new_n9877;
  assign new_n9879 = n7159 & n7690;
  assign new_n9880 = n3616 & n12489;
  assign new_n9881 = n10545 & n12777;
  assign new_n9882 = ~new_n9880 & ~new_n9881;
  assign new_n9883 = new_n9880 & new_n9881;
  assign new_n9884 = ~new_n9882 & ~new_n9883;
  assign new_n9885 = ~new_n9879 & ~new_n9884;
  assign new_n9886 = new_n9879 & new_n9884;
  assign new_n9887 = ~new_n9885 & ~new_n9886;
  assign new_n9888 = new_n9878 & ~new_n9887;
  assign new_n9889 = ~new_n9878 & new_n9887;
  assign new_n9890 = ~new_n9888 & ~new_n9889;
  assign new_n9891 = new_n9874 & new_n9890;
  assign new_n9892 = ~new_n9874 & ~new_n9890;
  assign new_n9893 = ~new_n9891 & ~new_n9892;
  assign new_n9894 = ~new_n9860 & new_n9893;
  assign new_n9895 = new_n9860 & ~new_n9893;
  assign new_n9896 = ~new_n9894 & ~new_n9895;
  assign new_n9897 = new_n9855 & new_n9896;
  assign new_n9898 = ~new_n9855 & ~new_n9896;
  assign new_n9899 = ~new_n9897 & ~new_n9898;
  assign new_n9900 = n447 & n5331;
  assign new_n9901 = new_n9834 & new_n9854;
  assign new_n9902 = ~new_n9855 & ~new_n9901;
  assign new_n9903 = new_n9900 & new_n9902;
  assign new_n9904 = ~new_n9845 & ~new_n9846;
  assign new_n9905 = ~new_n9850 & new_n9904;
  assign new_n9906 = new_n9850 & ~new_n9904;
  assign new_n9907 = ~new_n9905 & ~new_n9906;
  assign new_n9908 = new_n9357 & ~new_n9907;
  assign new_n9909 = ~new_n9840 & ~new_n9841;
  assign new_n9910 = new_n9852 & ~new_n9909;
  assign new_n9911 = ~new_n9852 & new_n9909;
  assign new_n9912 = ~new_n9910 & ~new_n9911;
  assign new_n9913 = new_n9908 & new_n9912;
  assign new_n9914 = ~new_n9900 & ~new_n9902;
  assign new_n9915 = ~new_n9903 & ~new_n9914;
  assign new_n9916 = new_n9913 & new_n9915;
  assign new_n9917 = ~new_n9903 & ~new_n9916;
  assign new_n9918 = new_n9899 & ~new_n9917;
  assign new_n9919 = ~new_n9899 & new_n9917;
  assign new_n9920_1 = ~new_n9918 & ~new_n9919;
  assign new_n9921 = new_n9788 & new_n9920_1;
  assign new_n9922 = ~new_n9737 & ~new_n9739;
  assign new_n9923 = ~new_n9740 & ~new_n9922;
  assign new_n9924 = ~new_n9913 & ~new_n9915;
  assign new_n9925 = ~new_n9916 & ~new_n9924;
  assign new_n9926 = ~new_n9923 & ~new_n9925;
  assign new_n9927 = new_n9923 & new_n9925;
  assign new_n9928 = ~new_n9908 & ~new_n9912;
  assign new_n9929 = ~new_n9913 & ~new_n9928;
  assign new_n9930 = ~new_n9732 & ~new_n9736;
  assign new_n9931 = ~new_n9737 & ~new_n9930;
  assign new_n9932 = ~new_n9929 & ~new_n9931;
  assign new_n9933 = new_n9929 & new_n9931;
  assign new_n9934 = ~new_n9357 & new_n9907;
  assign new_n9935 = ~new_n9908 & ~new_n9934;
  assign new_n9936 = ~new_n9727 & ~new_n9731;
  assign new_n9937 = ~new_n9732 & ~new_n9936;
  assign new_n9938_1 = new_n9935 & new_n9937;
  assign new_n9939 = ~new_n9935 & ~new_n9937;
  assign new_n9940 = ~new_n9372 & ~new_n9376;
  assign new_n9941 = ~new_n9373 & ~new_n9940;
  assign new_n9942 = ~new_n9939 & new_n9941;
  assign new_n9943 = ~new_n9938_1 & ~new_n9942;
  assign new_n9944 = ~new_n9933 & new_n9943;
  assign new_n9945 = ~new_n9932 & ~new_n9944;
  assign new_n9946 = ~new_n9927 & ~new_n9945;
  assign new_n9947 = ~new_n9926 & ~new_n9946;
  assign new_n9948 = new_n9921 & new_n9947;
  assign new_n9949 = ~new_n9788 & ~new_n9920_1;
  assign new_n9950 = ~new_n9947 & new_n9949;
  assign new_n9951 = ~new_n9921 & ~new_n9947;
  assign new_n9952 = ~new_n9949 & ~new_n9951;
  assign new_n9953 = ~new_n9950 & ~new_n9952;
  assign new_n9954 = ~new_n9948 & ~new_n9953;
  assign new_n9955 = new_n9657 & ~new_n9954;
  assign new_n9956_1 = ~new_n9657 & new_n9954;
  assign new_n9957 = ~new_n9955 & ~new_n9956_1;
  assign new_n9958 = ~new_n9605 & ~new_n9607;
  assign new_n9959 = ~new_n9608 & ~new_n9958;
  assign new_n9960 = ~new_n9926 & ~new_n9927;
  assign new_n9961 = new_n9945 & ~new_n9960;
  assign new_n9962 = ~new_n9945 & new_n9960;
  assign new_n9963 = ~new_n9961 & ~new_n9962;
  assign new_n9964 = new_n9959 & ~new_n9963;
  assign new_n9965 = ~new_n9959 & new_n9963;
  assign new_n9966 = ~new_n9600 & new_n9604;
  assign new_n9967 = ~new_n9605 & ~new_n9966;
  assign new_n9968 = ~new_n9932 & ~new_n9933;
  assign new_n9969 = new_n9943 & new_n9968;
  assign new_n9970 = ~new_n9943 & ~new_n9968;
  assign new_n9971 = ~new_n9969 & ~new_n9970;
  assign new_n9972 = new_n9967 & ~new_n9971;
  assign new_n9973 = ~new_n9967 & new_n9971;
  assign new_n9974 = ~new_n9595 & ~new_n9599;
  assign new_n9975 = ~new_n9600 & ~new_n9974;
  assign new_n9976 = ~new_n9938_1 & ~new_n9939;
  assign new_n9977 = ~new_n9941 & ~new_n9976;
  assign new_n9978 = new_n9941 & new_n9976;
  assign new_n9979 = ~new_n9977 & ~new_n9978;
  assign new_n9980 = new_n9975 & new_n9979;
  assign new_n9981 = ~new_n9975 & ~new_n9979;
  assign new_n9982 = ~new_n9346 & ~new_n9379;
  assign new_n9983 = ~new_n9345 & ~new_n9982;
  assign new_n9984 = ~new_n9981 & ~new_n9983;
  assign new_n9985 = ~new_n9980 & ~new_n9984;
  assign new_n9986 = ~new_n9973 & ~new_n9985;
  assign new_n9987 = ~new_n9972 & ~new_n9986;
  assign new_n9988 = ~new_n9965 & ~new_n9987;
  assign new_n9989 = ~new_n9964 & ~new_n9988;
  assign new_n9990 = ~new_n9957 & ~new_n9989;
  assign new_n9991 = ~new_n9955 & new_n9989;
  assign new_n9992 = ~new_n9956_1 & new_n9991;
  assign new_n9993 = ~new_n9990 & ~new_n9992;
  assign new_n9994 = new_n9524 & ~new_n9993;
  assign new_n9995 = ~new_n9524 & new_n9993;
  assign new_n9996 = ~new_n9517 & ~new_n9519;
  assign new_n9997 = ~new_n9520 & ~new_n9996;
  assign new_n9998 = ~new_n9964 & ~new_n9965;
  assign new_n9999 = new_n9987 & ~new_n9998;
  assign new_n10000 = ~new_n9987 & new_n9998;
  assign new_n10001 = ~new_n9999 & ~new_n10000;
  assign new_n10002 = ~new_n9997 & ~new_n10001;
  assign new_n10003 = new_n9997 & new_n10001;
  assign new_n10004 = ~new_n9512 & ~new_n9516;
  assign new_n10005 = ~new_n9517 & ~new_n10004;
  assign new_n10006 = ~new_n9972 & ~new_n9973;
  assign new_n10007 = ~new_n9985 & ~new_n10006;
  assign new_n10008 = new_n9985 & new_n10006;
  assign new_n10009 = ~new_n10007 & ~new_n10008;
  assign new_n10010 = new_n10005 & ~new_n10009;
  assign new_n10011 = ~new_n10005 & new_n10009;
  assign new_n10012 = ~new_n9507 & new_n9511;
  assign new_n10013 = ~new_n9512 & ~new_n10012;
  assign new_n10014 = ~new_n9980 & ~new_n9981;
  assign new_n10015 = ~new_n9983 & ~new_n10014;
  assign new_n10016 = new_n9983 & new_n10014;
  assign new_n10017 = ~new_n10015 & ~new_n10016;
  assign new_n10018 = new_n10013 & ~new_n10017;
  assign new_n10019 = ~new_n10013 & new_n10017;
  assign new_n10020 = ~new_n9330 & ~new_n9382;
  assign new_n10021 = ~new_n9329 & ~new_n10020;
  assign new_n10022_1 = ~new_n10019 & ~new_n10021;
  assign new_n10023 = ~new_n10018 & ~new_n10022_1;
  assign new_n10024 = ~new_n10011 & ~new_n10023;
  assign new_n10025 = ~new_n10010 & ~new_n10024;
  assign new_n10026 = ~new_n10003 & new_n10025;
  assign new_n10027 = ~new_n10002 & ~new_n10026;
  assign new_n10028 = ~new_n9995 & new_n10027;
  assign new_n10029 = ~new_n9994 & ~new_n10028;
  assign new_n10030 = ~new_n9652 & ~new_n9655;
  assign new_n10031 = ~new_n9467 & ~new_n9469;
  assign new_n10032 = ~new_n9470 & ~new_n10031;
  assign new_n10033 = n11877 & n12025;
  assign new_n10034 = n5212 & n11257;
  assign new_n10035 = ~new_n10033 & new_n10034;
  assign new_n10036 = new_n10033 & ~new_n10034;
  assign new_n10037 = ~new_n10035 & ~new_n10036;
  assign new_n10038 = n5964 & n9725;
  assign new_n10039 = n4312 & n5320;
  assign new_n10040 = n4370 & n12705;
  assign new_n10041 = new_n10039 & new_n10040;
  assign new_n10042 = ~new_n10039 & ~new_n10040;
  assign new_n10043 = ~new_n10041 & ~new_n10042;
  assign new_n10044 = new_n10038 & ~new_n10043;
  assign new_n10045 = ~new_n10038 & new_n10043;
  assign new_n10046 = ~new_n10044 & ~new_n10045;
  assign new_n10047 = ~new_n10037 & ~new_n10046;
  assign new_n10048 = new_n10037 & new_n10046;
  assign new_n10049 = ~new_n10047 & ~new_n10048;
  assign new_n10050 = ~new_n10032 & ~new_n10049;
  assign new_n10051 = new_n10032 & new_n10049;
  assign new_n10052 = ~new_n10050 & ~new_n10051;
  assign new_n10053 = ~new_n9475 & ~new_n9479;
  assign new_n10054 = ~new_n9478 & ~new_n10053;
  assign new_n10055 = n1097 & n12000;
  assign new_n10056 = ~new_n9459 & ~new_n9463;
  assign new_n10057 = ~new_n9462 & ~new_n10056;
  assign new_n10058 = ~new_n10055 & new_n10057;
  assign new_n10059 = new_n10055 & ~new_n10057;
  assign new_n10060 = ~new_n10058 & ~new_n10059;
  assign new_n10061 = ~new_n10054 & new_n10060;
  assign new_n10062 = new_n10054 & ~new_n10060;
  assign new_n10063 = ~new_n10061 & ~new_n10062;
  assign new_n10064 = ~new_n10052 & new_n10063;
  assign new_n10065 = new_n10052 & ~new_n10063;
  assign new_n10066 = ~new_n10064 & ~new_n10065;
  assign new_n10067 = ~new_n9474 & ~new_n9487;
  assign new_n10068 = ~new_n9486 & ~new_n10067;
  assign new_n10069 = ~new_n10066 & new_n10068;
  assign new_n10070 = new_n10066 & ~new_n10068;
  assign new_n10071 = ~new_n10069 & ~new_n10070;
  assign new_n10072 = ~new_n9872 & new_n9890;
  assign new_n10073 = ~new_n9873 & ~new_n10072;
  assign new_n10074 = ~new_n10071 & new_n10073;
  assign new_n10075 = new_n10071 & ~new_n10073;
  assign new_n10076 = ~new_n10074 & ~new_n10075;
  assign new_n10077 = new_n10030 & ~new_n10076;
  assign new_n10078 = ~new_n10030 & new_n10076;
  assign new_n10079 = ~new_n10077 & ~new_n10078;
  assign new_n10080 = ~new_n9783 & ~new_n9786;
  assign new_n10081 = n6776 & n7730;
  assign new_n10082 = ~new_n9625 & ~new_n9638;
  assign new_n10083 = ~new_n10081 & new_n10082;
  assign new_n10084 = new_n10081 & ~new_n10082;
  assign new_n10085 = ~new_n10083 & ~new_n10084;
  assign new_n10086 = n8717 & n12299;
  assign new_n10087 = n8276 & n8819;
  assign new_n10088 = n6429 & n9241;
  assign new_n10089 = ~new_n10087 & new_n10088;
  assign new_n10090 = new_n10087 & ~new_n10088;
  assign new_n10091 = ~new_n10089 & ~new_n10090;
  assign new_n10092 = new_n10086 & new_n10091;
  assign new_n10093 = ~new_n10086 & ~new_n10091;
  assign new_n10094 = ~new_n10092 & ~new_n10093;
  assign new_n10095 = ~new_n10085 & new_n10094;
  assign new_n10096 = new_n10085 & ~new_n10094;
  assign new_n10097 = ~new_n10095 & ~new_n10096;
  assign new_n10098 = n2433 & n7436;
  assign new_n10099 = new_n9612 & ~new_n9615;
  assign new_n10100 = ~new_n9616 & ~new_n10099;
  assign new_n10101 = ~new_n9628 & ~new_n9632;
  assign new_n10102 = ~new_n9631 & ~new_n10101;
  assign new_n10103 = ~new_n10100 & new_n10102;
  assign new_n10104 = new_n10100 & ~new_n10102;
  assign new_n10105 = ~new_n10103 & ~new_n10104;
  assign new_n10106 = new_n10098 & ~new_n10105;
  assign new_n10107 = ~new_n10098 & new_n10105;
  assign new_n10108 = ~new_n10106 & ~new_n10107;
  assign new_n10109 = ~new_n9622 & ~new_n9640_1;
  assign new_n10110 = ~new_n9621 & ~new_n10109;
  assign new_n10111 = new_n10108 & ~new_n10110;
  assign new_n10112 = ~new_n10108 & new_n10110;
  assign new_n10113 = ~new_n10111 & ~new_n10112;
  assign new_n10114 = ~new_n10097 & ~new_n10113;
  assign new_n10115 = new_n10097 & new_n10113;
  assign new_n10116 = ~new_n10114 & ~new_n10115;
  assign new_n10117 = ~new_n9745 & new_n9779;
  assign new_n10118 = ~new_n9743 & ~new_n10117;
  assign new_n10119 = n5760 & n5857;
  assign new_n10120 = n45 & n10990;
  assign new_n10121 = ~new_n10119 & new_n10120;
  assign new_n10122 = new_n10119 & ~new_n10120;
  assign new_n10123 = ~new_n10121 & ~new_n10122;
  assign new_n10124 = n1478 & n3986;
  assign new_n10125 = n7965 & n10022;
  assign new_n10126 = ~new_n10124 & ~new_n10125;
  assign new_n10127 = new_n10124 & new_n10125;
  assign new_n10128 = ~new_n10126 & ~new_n10127;
  assign new_n10129 = ~new_n10123 & new_n10128;
  assign new_n10130 = new_n10123 & ~new_n10128;
  assign new_n10131 = ~new_n10129 & ~new_n10130;
  assign new_n10132 = new_n10118 & new_n10131;
  assign new_n10133 = ~new_n10118 & ~new_n10131;
  assign new_n10134 = ~new_n10132 & ~new_n10133;
  assign new_n10135 = ~new_n10116 & new_n10134;
  assign new_n10136 = new_n10116 & ~new_n10134;
  assign new_n10137 = ~new_n10135 & ~new_n10136;
  assign new_n10138 = new_n10080 & new_n10137;
  assign new_n10139 = ~new_n10080 & ~new_n10137;
  assign new_n10140 = ~new_n10138 & ~new_n10139;
  assign new_n10141 = ~new_n9643 & ~new_n9647;
  assign new_n10142 = ~new_n9645 & ~new_n10141;
  assign new_n10143 = n10510 & n11728;
  assign new_n10144 = n10644 & n12709;
  assign new_n10145 = n1198 & n8759;
  assign new_n10146 = new_n10144 & ~new_n10145;
  assign new_n10147 = ~new_n10144 & new_n10145;
  assign new_n10148 = ~new_n10146 & ~new_n10147;
  assign new_n10149 = new_n10143 & ~new_n10148;
  assign new_n10150 = ~new_n10143 & new_n10148;
  assign new_n10151 = ~new_n10149 & ~new_n10150;
  assign new_n10152 = new_n10142 & new_n10151;
  assign new_n10153 = ~new_n10142 & ~new_n10151;
  assign new_n10154 = ~new_n10152 & ~new_n10153;
  assign new_n10155 = ~new_n10140 & new_n10154;
  assign new_n10156 = new_n10140 & ~new_n10154;
  assign new_n10157 = ~new_n10155 & ~new_n10156;
  assign new_n10158 = ~new_n9952 & ~new_n10157;
  assign new_n10159 = new_n9952 & new_n10157;
  assign new_n10160 = ~new_n10158 & ~new_n10159;
  assign new_n10161 = ~new_n10079 & new_n10160;
  assign new_n10162 = new_n10079 & ~new_n10160;
  assign new_n10163 = ~new_n10161 & ~new_n10162;
  assign new_n10164 = ~new_n9956_1 & ~new_n9991;
  assign new_n10165 = n5305 & n6604;
  assign new_n10166 = new_n9491 & ~new_n9494;
  assign new_n10167 = ~new_n9495 & ~new_n10166;
  assign new_n10168 = n10547 & n11407;
  assign new_n10169 = new_n9863 & ~new_n9866;
  assign new_n10170 = ~new_n9867 & ~new_n10169;
  assign new_n10171 = ~new_n10168 & new_n10170;
  assign new_n10172 = new_n10168 & ~new_n10170;
  assign new_n10173 = ~new_n10171 & ~new_n10172;
  assign new_n10174_1 = new_n10167 & ~new_n10173;
  assign new_n10175 = ~new_n10167 & new_n10173;
  assign new_n10176 = ~new_n10174_1 & ~new_n10175;
  assign new_n10177 = ~new_n10165 & new_n10176;
  assign new_n10178 = new_n10165 & ~new_n10176;
  assign new_n10179 = ~new_n10177 & ~new_n10178;
  assign new_n10180 = ~new_n9858 & ~new_n9893;
  assign new_n10181 = ~new_n9859 & ~new_n10180;
  assign new_n10182 = n4436 & n5331;
  assign new_n10183 = n4499 & n12489;
  assign new_n10184 = ~new_n10182 & new_n10183;
  assign new_n10185 = new_n10182 & ~new_n10183;
  assign new_n10186 = ~new_n10184 & ~new_n10185;
  assign new_n10187 = ~new_n9758 & new_n9776;
  assign new_n10188 = ~new_n9759 & ~new_n10187;
  assign new_n10189 = ~new_n10186 & new_n10188;
  assign new_n10190 = new_n10186 & ~new_n10188;
  assign new_n10191 = ~new_n10189 & ~new_n10190;
  assign new_n10192 = new_n10181 & new_n10191;
  assign new_n10193 = ~new_n10181 & ~new_n10191;
  assign new_n10194 = ~new_n10192 & ~new_n10193;
  assign new_n10195 = ~new_n9876 & ~new_n9887;
  assign new_n10196 = ~new_n9877 & ~new_n10195;
  assign new_n10197 = n447 & n2530;
  assign new_n10198 = ~new_n9879 & ~new_n9883;
  assign new_n10199 = ~new_n9882 & ~new_n10198;
  assign new_n10200 = ~new_n10197 & new_n10199;
  assign new_n10201 = new_n10197 & ~new_n10199;
  assign new_n10202 = ~new_n10200 & ~new_n10201;
  assign new_n10203 = new_n10196 & ~new_n10202;
  assign new_n10204 = ~new_n10196 & new_n10202;
  assign new_n10205 = ~new_n10203 & ~new_n10204;
  assign new_n10206 = ~new_n9763_1 & new_n9773;
  assign new_n10207 = ~new_n9762 & ~new_n10206;
  assign new_n10208 = new_n9765 & ~new_n9768;
  assign new_n10209 = ~new_n9769 & ~new_n10208;
  assign new_n10210 = new_n9749 & ~new_n9752;
  assign new_n10211 = ~new_n9753 & ~new_n10210;
  assign new_n10212 = ~new_n10209 & ~new_n10211;
  assign new_n10213 = new_n10209 & new_n10211;
  assign new_n10214 = ~new_n10212 & ~new_n10213;
  assign new_n10215 = n6441 & n11892;
  assign new_n10216 = n5860 & n11791;
  assign new_n10217_1 = new_n10215 & ~new_n10216;
  assign new_n10218 = ~new_n10215 & new_n10216;
  assign new_n10219 = ~new_n10217_1 & ~new_n10218;
  assign new_n10220 = n7388 & n11999;
  assign new_n10221 = n2393 & n12947;
  assign new_n10222 = ~new_n10220 & ~new_n10221;
  assign new_n10223_1 = new_n10220 & new_n10221;
  assign new_n10224 = ~new_n10222 & ~new_n10223_1;
  assign new_n10225 = ~new_n10219 & new_n10224;
  assign new_n10226 = new_n10219 & ~new_n10224;
  assign new_n10227 = ~new_n10225 & ~new_n10226;
  assign new_n10228 = ~new_n10214 & new_n10227;
  assign new_n10229 = new_n10214 & ~new_n10227;
  assign new_n10230 = ~new_n10228 & ~new_n10229;
  assign new_n10231 = new_n10207 & new_n10230;
  assign new_n10232 = ~new_n10207 & ~new_n10230;
  assign new_n10233 = ~new_n10231 & ~new_n10232;
  assign new_n10234 = n11967 & n12648;
  assign new_n10235 = n6254 & n10545;
  assign new_n10236 = ~new_n10234 & ~new_n10235;
  assign new_n10237 = new_n10234 & new_n10235;
  assign new_n10238 = ~new_n10236 & ~new_n10237;
  assign new_n10239 = n7690 & n12777;
  assign new_n10240 = n3616 & n7159;
  assign new_n10241 = new_n10239 & ~new_n10240;
  assign new_n10242 = ~new_n10239 & new_n10240;
  assign new_n10243 = ~new_n10241 & ~new_n10242;
  assign new_n10244 = ~new_n10238 & ~new_n10243;
  assign new_n10245 = new_n10238 & new_n10243;
  assign new_n10246 = ~new_n10244 & ~new_n10245;
  assign new_n10247 = new_n10233 & new_n10246;
  assign new_n10248 = ~new_n10233 & ~new_n10246;
  assign new_n10249 = ~new_n10247 & ~new_n10248;
  assign new_n10250 = new_n10205 & ~new_n10249;
  assign new_n10251 = ~new_n10205 & new_n10249;
  assign new_n10252 = ~new_n10250 & ~new_n10251;
  assign new_n10253 = ~new_n10194 & ~new_n10252;
  assign new_n10254 = new_n10194 & new_n10252;
  assign new_n10255 = ~new_n10253 & ~new_n10254;
  assign new_n10256 = n1353 & n8476;
  assign new_n10257 = new_n10255 & ~new_n10256;
  assign new_n10258 = ~new_n10255 & new_n10256;
  assign new_n10259 = ~new_n10257 & ~new_n10258;
  assign new_n10260 = ~new_n10179 & new_n10259;
  assign new_n10261 = new_n10179 & ~new_n10259;
  assign new_n10262 = ~new_n10260 & ~new_n10261;
  assign new_n10263 = ~new_n9500 & ~new_n9522;
  assign new_n10264 = ~new_n9897 & ~new_n9918;
  assign new_n10265 = new_n10263 & new_n10264;
  assign new_n10266 = ~new_n10263 & ~new_n10264;
  assign new_n10267 = ~new_n10265 & ~new_n10266;
  assign new_n10268 = new_n10262 & new_n10267;
  assign new_n10269 = ~new_n10262 & ~new_n10267;
  assign new_n10270 = ~new_n10268 & ~new_n10269;
  assign new_n10271 = new_n10164 & new_n10270;
  assign new_n10272 = ~new_n10164 & ~new_n10270;
  assign new_n10273 = ~new_n10271 & ~new_n10272;
  assign new_n10274 = new_n10163 & ~new_n10273;
  assign new_n10275 = ~new_n10163 & new_n10273;
  assign new_n10276 = ~new_n10274 & ~new_n10275;
  assign new_n10277 = ~new_n10029 & ~new_n10276;
  assign new_n10278_1 = new_n10029 & new_n10276;
  assign n3287 = new_n10277 | new_n10278_1;
  assign new_n10280 = ~new_n10002 & ~new_n10003;
  assign new_n10281 = new_n10025 & new_n10280;
  assign new_n10282 = ~new_n10025 & ~new_n10280;
  assign n3339 = new_n10281 | new_n10282;
  assign new_n10284 = ~new_n4458 & ~new_n4459;
  assign new_n10285 = ~new_n4463 & ~new_n10284;
  assign new_n10286 = new_n4463 & new_n10284;
  assign n3456 = ~new_n10285 & ~new_n10286;
  assign new_n10288 = n4005 & n6687;
  assign new_n10289 = n2585 & n6687;
  assign new_n10290 = n2508 & n6687;
  assign new_n10291 = n6687 & n12720;
  assign new_n10292 = n2509 & n2564;
  assign new_n10293 = new_n10291 & new_n10292;
  assign new_n10294 = n4189 & n6038;
  assign new_n10295 = ~new_n10291 & ~new_n10292;
  assign new_n10296 = new_n10294 & ~new_n10295;
  assign new_n10297 = ~new_n10293 & ~new_n10296;
  assign new_n10298 = ~new_n10290 & new_n10297;
  assign new_n10299 = new_n10290 & ~new_n10297;
  assign new_n10300 = n2564 & n12720;
  assign new_n10301 = n6038 & n6770;
  assign new_n10302 = n2509 & n4189;
  assign new_n10303 = ~new_n10301 & ~new_n10302;
  assign new_n10304 = n2509 & n6770;
  assign new_n10305 = new_n10294 & new_n10304;
  assign new_n10306 = ~new_n10303 & ~new_n10305;
  assign new_n10307 = ~new_n10300 & ~new_n10306;
  assign new_n10308 = new_n10300 & new_n10306;
  assign new_n10309 = ~new_n10307 & ~new_n10308;
  assign new_n10310 = ~new_n10299 & ~new_n10309;
  assign new_n10311 = ~new_n10298 & ~new_n10310;
  assign new_n10312 = ~new_n10289 & ~new_n10311;
  assign new_n10313 = new_n10289 & new_n10311;
  assign new_n10314 = n2508 & n2564;
  assign new_n10315 = new_n10300 & ~new_n10303;
  assign new_n10316 = ~new_n10305 & ~new_n10315;
  assign new_n10317 = ~new_n10314 & new_n10316;
  assign new_n10318 = new_n10314 & ~new_n10316;
  assign new_n10319 = ~new_n10317 & ~new_n10318;
  assign new_n10320 = n6038 & n9920;
  assign new_n10321 = n4189 & n12720;
  assign new_n10322 = ~new_n10320 & ~new_n10321;
  assign new_n10323 = new_n10320 & new_n10321;
  assign new_n10324 = ~new_n10322 & ~new_n10323;
  assign new_n10325 = ~new_n10304 & ~new_n10324;
  assign new_n10326 = new_n10304 & new_n10324;
  assign new_n10327_1 = ~new_n10325 & ~new_n10326;
  assign new_n10328 = ~new_n10319 & new_n10327_1;
  assign new_n10329 = ~new_n10318 & ~new_n10327_1;
  assign new_n10330 = ~new_n10317 & new_n10329;
  assign new_n10331 = ~new_n10328 & ~new_n10330;
  assign new_n10332 = ~new_n10313 & new_n10331;
  assign new_n10333 = ~new_n10312 & ~new_n10332;
  assign new_n10334 = n2564 & n2585;
  assign new_n10335 = n2508 & n4189;
  assign new_n10336 = ~new_n10334 & ~new_n10335;
  assign new_n10337 = new_n10334 & new_n10335;
  assign new_n10338 = ~new_n10336 & ~new_n10337;
  assign new_n10339 = ~new_n10317 & ~new_n10329;
  assign new_n10340 = ~new_n10338 & ~new_n10339;
  assign new_n10341 = new_n10338 & new_n10339;
  assign new_n10342 = ~new_n10340 & ~new_n10341;
  assign new_n10343 = new_n10304 & ~new_n10322;
  assign new_n10344 = ~new_n10323 & ~new_n10343;
  assign new_n10345 = n6770 & n12720;
  assign new_n10346 = n2509 & n9920;
  assign new_n10347 = n3627 & n6038;
  assign new_n10348 = ~new_n10346 & ~new_n10347;
  assign new_n10349 = new_n10346 & new_n10347;
  assign new_n10350 = ~new_n10348 & ~new_n10349;
  assign new_n10351 = new_n10345 & new_n10350;
  assign new_n10352 = ~new_n10345 & ~new_n10350;
  assign new_n10353 = ~new_n10351 & ~new_n10352;
  assign new_n10354 = new_n10344 & ~new_n10353;
  assign new_n10355 = ~new_n10344 & new_n10353;
  assign new_n10356 = ~new_n10354 & ~new_n10355;
  assign new_n10357 = new_n10342 & ~new_n10356;
  assign new_n10358 = ~new_n10342 & new_n10356;
  assign new_n10359 = ~new_n10357 & ~new_n10358;
  assign new_n10360 = new_n10333 & ~new_n10359;
  assign new_n10361 = ~new_n10333 & new_n10359;
  assign new_n10362 = ~new_n10360 & ~new_n10361;
  assign new_n10363 = new_n10288 & new_n10362;
  assign new_n10364 = n2509 & n6687;
  assign new_n10365 = n2564 & n6038;
  assign new_n10366 = new_n10364 & new_n10365;
  assign new_n10367 = ~new_n10293 & ~new_n10295;
  assign new_n10368 = ~new_n10294 & ~new_n10367;
  assign new_n10369 = new_n10294 & new_n10367;
  assign new_n10370 = ~new_n10368 & ~new_n10369;
  assign new_n10371 = new_n10366 & new_n10370;
  assign new_n10372 = ~new_n10298 & new_n10310;
  assign new_n10373 = ~new_n10298 & ~new_n10299;
  assign new_n10374 = new_n10309 & ~new_n10373;
  assign new_n10375 = ~new_n10372 & ~new_n10374;
  assign new_n10376 = new_n10371 & ~new_n10375;
  assign new_n10377 = ~new_n10312 & ~new_n10313;
  assign new_n10378 = ~new_n10331 & ~new_n10377;
  assign new_n10379 = new_n10331 & new_n10377;
  assign new_n10380 = ~new_n10378 & ~new_n10379;
  assign new_n10381 = new_n10376 & ~new_n10380;
  assign new_n10382 = ~new_n10288 & ~new_n10362;
  assign new_n10383 = ~new_n10363 & ~new_n10382;
  assign new_n10384 = new_n10381 & new_n10383;
  assign new_n10385 = ~new_n10363 & ~new_n10384;
  assign new_n10386 = ~new_n10340 & new_n10356;
  assign new_n10387 = ~new_n10337 & ~new_n10386;
  assign new_n10388 = ~new_n10341 & new_n10387;
  assign new_n10389 = new_n10337 & new_n10386;
  assign new_n10390 = ~new_n10388 & ~new_n10389;
  assign new_n10391_1 = n2564 & n4005;
  assign new_n10392 = n2585 & n4189;
  assign new_n10393 = n6687 & n12706;
  assign new_n10394 = ~new_n10392 & ~new_n10393;
  assign new_n10395 = new_n10392 & new_n10393;
  assign new_n10396 = ~new_n10394 & ~new_n10395;
  assign new_n10397 = ~new_n10391_1 & ~new_n10396;
  assign new_n10398 = new_n10391_1 & new_n10396;
  assign new_n10399 = ~new_n10397 & ~new_n10398;
  assign new_n10400 = new_n10344 & ~new_n10351;
  assign new_n10401 = ~new_n10352 & ~new_n10400;
  assign new_n10402 = ~new_n10399 & ~new_n10401;
  assign new_n10403 = n2508 & n6770;
  assign new_n10404 = new_n10349 & new_n10403;
  assign new_n10405 = ~new_n10349 & ~new_n10403;
  assign new_n10406 = ~new_n10404 & ~new_n10405;
  assign new_n10407 = n4516 & n6038;
  assign new_n10408 = n2509 & n3627;
  assign new_n10409 = n9920 & n12720;
  assign new_n10410 = ~new_n10408 & ~new_n10409;
  assign new_n10411 = new_n10408 & new_n10409;
  assign new_n10412 = ~new_n10410 & ~new_n10411;
  assign new_n10413 = new_n10407 & ~new_n10412;
  assign new_n10414 = ~new_n10407 & new_n10412;
  assign new_n10415 = ~new_n10413 & ~new_n10414;
  assign new_n10416 = new_n10406 & new_n10415;
  assign new_n10417 = ~new_n10406 & ~new_n10415;
  assign new_n10418 = ~new_n10416 & ~new_n10417;
  assign new_n10419 = new_n10402 & new_n10418;
  assign new_n10420 = new_n10399 & new_n10401;
  assign new_n10421 = new_n10418 & ~new_n10420;
  assign new_n10422 = ~new_n10402 & ~new_n10421;
  assign new_n10423 = ~new_n10418 & new_n10420;
  assign new_n10424 = new_n10422 & ~new_n10423;
  assign new_n10425 = ~new_n10419 & ~new_n10424;
  assign new_n10426 = ~new_n10390 & ~new_n10425;
  assign new_n10427 = new_n10390 & new_n10425;
  assign new_n10428 = ~new_n10426 & ~new_n10427;
  assign new_n10429 = new_n10360 & new_n10428;
  assign new_n10430 = ~new_n10360 & ~new_n10428;
  assign new_n10431 = ~new_n10429 & ~new_n10430;
  assign new_n10432 = ~new_n10385 & new_n10431;
  assign new_n10433 = new_n10385 & ~new_n10431;
  assign new_n10434 = ~new_n10432 & ~new_n10433;
  assign new_n10435 = n4928 & n8336;
  assign new_n10436 = n5105 & n10928;
  assign new_n10437 = n1209 & n10928;
  assign new_n10438 = n6986 & n7500;
  assign new_n10439_1 = new_n10437 & new_n10438;
  assign new_n10440 = n2226 & n7354;
  assign new_n10441 = ~new_n10437 & ~new_n10438;
  assign new_n10442 = new_n10440 & ~new_n10441;
  assign new_n10443 = ~new_n10439_1 & ~new_n10442;
  assign new_n10444 = ~new_n10436 & new_n10443;
  assign new_n10445 = new_n10436 & ~new_n10443;
  assign new_n10446 = n1209 & n6986;
  assign new_n10447 = n1094 & n7354;
  assign new_n10448 = n2226 & n7500;
  assign new_n10449 = ~new_n10447 & ~new_n10448;
  assign new_n10450 = new_n10447 & new_n10448;
  assign new_n10451_1 = ~new_n10449 & ~new_n10450;
  assign new_n10452 = ~new_n10446 & ~new_n10451_1;
  assign new_n10453 = new_n10446 & new_n10451_1;
  assign new_n10454 = ~new_n10452 & ~new_n10453;
  assign new_n10455 = ~new_n10445 & ~new_n10454;
  assign new_n10456 = ~new_n10444 & ~new_n10455;
  assign new_n10457 = n4141 & n10928;
  assign new_n10458 = n5105 & n6986;
  assign new_n10459 = ~new_n10457 & ~new_n10458;
  assign new_n10460 = new_n10457 & new_n10458;
  assign new_n10461 = ~new_n10459 & ~new_n10460;
  assign new_n10462 = n1094 & n7500;
  assign new_n10463 = n7354 & n10678;
  assign new_n10464 = new_n10462 & new_n10463;
  assign new_n10465 = ~new_n10462 & ~new_n10463;
  assign new_n10466 = ~new_n10464 & ~new_n10465;
  assign new_n10467 = n1209 & n2226;
  assign new_n10468 = new_n10446 & ~new_n10449;
  assign new_n10469 = ~new_n10450 & ~new_n10468;
  assign new_n10470 = ~new_n10467 & new_n10469;
  assign new_n10471 = new_n10467 & ~new_n10469;
  assign new_n10472 = ~new_n10470 & ~new_n10471;
  assign new_n10473 = ~new_n10466 & ~new_n10472;
  assign new_n10474 = new_n10466 & new_n10472;
  assign new_n10475 = ~new_n10473 & ~new_n10474;
  assign new_n10476_1 = new_n10461 & new_n10475;
  assign new_n10477 = ~new_n10461 & ~new_n10475;
  assign new_n10478 = ~new_n10476_1 & ~new_n10477;
  assign new_n10479 = ~new_n10456 & new_n10478;
  assign new_n10480 = new_n10456 & ~new_n10478;
  assign new_n10481 = ~new_n10479 & ~new_n10480;
  assign new_n10482 = n4141 & n8336;
  assign new_n10483 = n5105 & n8336;
  assign new_n10484 = n7500 & n10928;
  assign new_n10485 = n1209 & n8336;
  assign new_n10486 = n6986 & n7354;
  assign new_n10487 = ~new_n10485 & ~new_n10486;
  assign new_n10488 = new_n10484 & ~new_n10487;
  assign new_n10489 = new_n378 & new_n10446;
  assign new_n10490 = ~new_n10488 & ~new_n10489;
  assign new_n10491 = ~new_n10483 & new_n10490;
  assign new_n10492 = new_n10483 & ~new_n10490;
  assign new_n10493 = ~new_n10439_1 & ~new_n10441;
  assign new_n10494 = ~new_n10440 & ~new_n10493;
  assign new_n10495 = new_n10440 & new_n10493;
  assign new_n10496 = ~new_n10494 & ~new_n10495;
  assign new_n10497 = ~new_n10492 & ~new_n10496;
  assign new_n10498 = ~new_n10491 & ~new_n10497;
  assign new_n10499 = new_n10482 & new_n10498;
  assign new_n10500 = ~new_n10482 & ~new_n10498;
  assign new_n10501 = ~new_n10444 & ~new_n10445;
  assign new_n10502 = new_n10454 & ~new_n10501;
  assign new_n10503 = ~new_n10454 & new_n10501;
  assign new_n10504 = ~new_n10502 & ~new_n10503;
  assign new_n10505 = ~new_n10500 & ~new_n10504;
  assign new_n10506 = ~new_n10499 & ~new_n10505;
  assign new_n10507 = ~new_n10481 & ~new_n10506;
  assign new_n10508 = new_n10481 & new_n10506;
  assign new_n10509 = ~new_n10507 & ~new_n10508;
  assign new_n10510_1 = new_n10435 & new_n10509;
  assign new_n10511 = ~new_n10487 & ~new_n10489;
  assign new_n10512 = n7500 & n8336;
  assign new_n10513 = n7354 & n10928;
  assign new_n10514 = new_n10512 & new_n10513;
  assign new_n10515 = ~new_n10511 & new_n10514;
  assign new_n10516 = ~new_n10491 & ~new_n10492;
  assign new_n10517 = ~new_n10496 & new_n10516;
  assign new_n10518 = new_n10496 & ~new_n10516;
  assign new_n10519 = ~new_n10517 & ~new_n10518;
  assign new_n10520 = new_n10515 & ~new_n10519;
  assign new_n10521 = ~new_n10499 & ~new_n10500;
  assign new_n10522 = ~new_n10504 & new_n10521;
  assign new_n10523 = new_n10504 & ~new_n10521;
  assign new_n10524 = ~new_n10522 & ~new_n10523;
  assign new_n10525 = new_n10520 & new_n10524;
  assign new_n10526 = ~new_n10435 & ~new_n10509;
  assign new_n10527 = ~new_n10510_1 & ~new_n10526;
  assign new_n10528 = new_n10525 & new_n10527;
  assign new_n10529 = ~new_n10510_1 & ~new_n10528;
  assign new_n10530 = new_n10456 & ~new_n10477;
  assign new_n10531 = new_n10460 & new_n10530;
  assign new_n10532 = ~new_n10460 & ~new_n10530;
  assign new_n10533 = ~new_n10476_1 & new_n10532;
  assign new_n10534 = ~new_n10531 & ~new_n10533;
  assign new_n10535 = n7500 & n10678;
  assign new_n10536 = n7320 & n7354;
  assign new_n10537 = n1094 & n1209;
  assign new_n10538 = ~new_n10536 & ~new_n10537;
  assign new_n10539 = new_n10536 & new_n10537;
  assign new_n10540 = ~new_n10538 & ~new_n10539;
  assign new_n10541 = ~new_n10535 & ~new_n10540;
  assign new_n10542 = new_n10535 & new_n10540;
  assign new_n10543 = ~new_n10541 & ~new_n10542;
  assign new_n10544 = n2226 & n5105;
  assign new_n10545_1 = new_n10464 & new_n10544;
  assign new_n10546 = ~new_n10464 & ~new_n10544;
  assign new_n10547_1 = ~new_n10545_1 & ~new_n10546;
  assign new_n10548 = new_n10543 & ~new_n10547_1;
  assign new_n10549 = ~new_n10543 & new_n10547_1;
  assign new_n10550 = ~new_n10548 & ~new_n10549;
  assign new_n10551 = n4928 & n10928;
  assign new_n10552 = n4141 & n6986;
  assign new_n10553 = n8236 & n8336;
  assign new_n10554 = ~new_n10552 & ~new_n10553;
  assign new_n10555 = new_n10552 & new_n10553;
  assign new_n10556 = ~new_n10554 & ~new_n10555;
  assign new_n10557 = ~new_n10551 & ~new_n10556;
  assign new_n10558 = new_n10551 & new_n10556;
  assign new_n10559 = ~new_n10557 & ~new_n10558;
  assign new_n10560 = new_n10466 & ~new_n10470;
  assign new_n10561 = ~new_n10471 & ~new_n10560;
  assign new_n10562 = ~new_n10559 & new_n10561;
  assign new_n10563 = new_n10559 & ~new_n10561;
  assign new_n10564 = ~new_n10562 & ~new_n10563;
  assign new_n10565 = new_n10550 & new_n10564;
  assign new_n10566 = ~new_n10550 & ~new_n10564;
  assign new_n10567 = ~new_n10565 & ~new_n10566;
  assign new_n10568 = new_n10534 & new_n10567;
  assign new_n10569 = ~new_n10534 & ~new_n10567;
  assign new_n10570 = ~new_n10568 & ~new_n10569;
  assign new_n10571 = new_n10507 & ~new_n10570;
  assign new_n10572 = ~new_n10507 & new_n10570;
  assign new_n10573 = ~new_n10571 & ~new_n10572;
  assign new_n10574 = ~new_n10529 & new_n10573;
  assign new_n10575 = new_n10529 & ~new_n10573;
  assign new_n10576 = ~new_n10574 & ~new_n10575;
  assign new_n10577 = n5814 & n11222;
  assign new_n10578 = n11222 & n12704;
  assign new_n10579 = n7294 & n11153;
  assign new_n10580 = n1980 & n11153;
  assign new_n10581 = n5314 & n10848;
  assign new_n10582 = new_n10580 & new_n10581;
  assign new_n10583 = n996 & n8028;
  assign new_n10584 = ~new_n10580 & ~new_n10581;
  assign new_n10585 = new_n10583 & ~new_n10584;
  assign new_n10586 = ~new_n10582 & ~new_n10585;
  assign new_n10587 = ~new_n10579 & new_n10586;
  assign new_n10588 = new_n10579 & ~new_n10586;
  assign new_n10589_1 = ~new_n10587 & ~new_n10588;
  assign new_n10590 = n5767 & n8028;
  assign new_n10591 = n1980 & n5314;
  assign new_n10592 = n996 & n10848;
  assign new_n10593 = ~new_n10591 & ~new_n10592;
  assign new_n10594 = new_n10591 & new_n10592;
  assign new_n10595 = ~new_n10593 & ~new_n10594;
  assign new_n10596 = new_n10590 & ~new_n10595;
  assign new_n10597 = ~new_n10590 & new_n10595;
  assign new_n10598 = ~new_n10596 & ~new_n10597;
  assign new_n10599 = ~new_n10589_1 & new_n10598;
  assign new_n10600 = new_n10589_1 & ~new_n10598;
  assign new_n10601 = ~new_n10599 & ~new_n10600;
  assign new_n10602 = new_n10578 & new_n10601;
  assign new_n10603 = ~new_n10578 & ~new_n10601;
  assign new_n10604 = n7294 & n11222;
  assign new_n10605 = n10848 & n11153;
  assign new_n10606 = n1980 & n11222;
  assign new_n10607 = new_n10605 & new_n10606;
  assign new_n10608 = n5314 & n8028;
  assign new_n10609 = ~new_n10605 & ~new_n10606;
  assign new_n10610 = new_n10608 & ~new_n10609;
  assign new_n10611 = ~new_n10607 & ~new_n10610;
  assign new_n10612 = ~new_n10604 & new_n10611;
  assign new_n10613 = new_n10604 & ~new_n10611;
  assign new_n10614 = ~new_n10582 & ~new_n10584;
  assign new_n10615 = new_n10583 & ~new_n10614;
  assign new_n10616 = ~new_n10583 & new_n10614;
  assign new_n10617 = ~new_n10615 & ~new_n10616;
  assign new_n10618 = ~new_n10613 & new_n10617;
  assign new_n10619 = ~new_n10612 & ~new_n10618;
  assign new_n10620 = ~new_n10603 & new_n10619;
  assign new_n10621 = ~new_n10602 & ~new_n10620;
  assign new_n10622 = n11153 & n12704;
  assign new_n10623 = n5314 & n7294;
  assign new_n10624 = ~new_n10622 & ~new_n10623;
  assign new_n10625 = new_n10622 & new_n10623;
  assign new_n10626 = ~new_n10624 & ~new_n10625;
  assign new_n10627 = n996 & n1980;
  assign new_n10628 = n5319 & n8028;
  assign new_n10629 = n5767 & n10848;
  assign new_n10630 = ~new_n10628 & ~new_n10629;
  assign new_n10631 = new_n10628 & new_n10629;
  assign new_n10632 = ~new_n10630 & ~new_n10631;
  assign new_n10633 = ~new_n10627 & ~new_n10632;
  assign new_n10634 = new_n10590 & ~new_n10593;
  assign new_n10635 = ~new_n10594 & ~new_n10634;
  assign new_n10636 = new_n10633 & new_n10635;
  assign new_n10637 = new_n10627 & new_n10632;
  assign new_n10638 = new_n10635 & ~new_n10637;
  assign new_n10639 = ~new_n10633 & ~new_n10638;
  assign new_n10640 = ~new_n10636 & ~new_n10639;
  assign new_n10641 = ~new_n10635 & new_n10637;
  assign new_n10642 = ~new_n10640 & ~new_n10641;
  assign new_n10643 = new_n10626 & ~new_n10642;
  assign new_n10644_1 = ~new_n10626 & new_n10642;
  assign new_n10645 = ~new_n10643 & ~new_n10644_1;
  assign new_n10646 = ~new_n10587 & ~new_n10598;
  assign new_n10647 = ~new_n10588 & ~new_n10646;
  assign new_n10648 = new_n10645 & new_n10647;
  assign new_n10649 = ~new_n10645 & ~new_n10647;
  assign new_n10650 = ~new_n10648 & ~new_n10649;
  assign new_n10651 = ~new_n10621 & ~new_n10650;
  assign new_n10652 = new_n10621 & new_n10650;
  assign new_n10653 = ~new_n10651 & ~new_n10652;
  assign new_n10654 = new_n10577 & new_n10653;
  assign new_n10655 = n10848 & n11222;
  assign new_n10656 = n8028 & n11153;
  assign new_n10657 = new_n10655 & new_n10656;
  assign new_n10658 = ~new_n10607 & ~new_n10609;
  assign new_n10659 = new_n10608 & ~new_n10658;
  assign new_n10660 = ~new_n10608 & new_n10658;
  assign new_n10661 = ~new_n10659 & ~new_n10660;
  assign new_n10662 = new_n10657 & ~new_n10661;
  assign new_n10663 = ~new_n10612 & ~new_n10613;
  assign new_n10664 = new_n10617 & new_n10663;
  assign new_n10665 = ~new_n10617 & ~new_n10663;
  assign new_n10666 = ~new_n10664 & ~new_n10665;
  assign new_n10667 = new_n10662 & ~new_n10666;
  assign new_n10668 = new_n10603 & ~new_n10619;
  assign new_n10669 = new_n10602 & new_n10619;
  assign new_n10670 = ~new_n10621 & ~new_n10669;
  assign new_n10671 = ~new_n10668 & ~new_n10670;
  assign new_n10672 = new_n10667 & new_n10671;
  assign new_n10673 = ~new_n10577 & ~new_n10653;
  assign new_n10674 = ~new_n10654 & ~new_n10673;
  assign new_n10675 = new_n10672 & new_n10674;
  assign new_n10676 = ~new_n10654 & ~new_n10675;
  assign new_n10677 = ~new_n10644_1 & ~new_n10647;
  assign new_n10678_1 = ~new_n10625 & ~new_n10677;
  assign new_n10679 = ~new_n10643 & new_n10678_1;
  assign new_n10680 = new_n10625 & new_n10677;
  assign new_n10681 = ~new_n10679 & ~new_n10680;
  assign new_n10682 = n5814 & n11153;
  assign new_n10683 = n5314 & n12704;
  assign new_n10684 = n4903 & n11222;
  assign new_n10685_1 = ~new_n10683 & ~new_n10684;
  assign new_n10686 = new_n10683 & new_n10684;
  assign new_n10687 = ~new_n10685_1 & ~new_n10686;
  assign new_n10688 = ~new_n10682 & ~new_n10687;
  assign new_n10689 = new_n10682 & new_n10687;
  assign new_n10690 = ~new_n10688 & ~new_n10689;
  assign new_n10691 = new_n10639 & new_n10690;
  assign new_n10692 = ~new_n10639 & ~new_n10690;
  assign new_n10693 = ~new_n10691 & ~new_n10692;
  assign new_n10694 = n996 & n7294;
  assign new_n10695_1 = new_n10631 & new_n10694;
  assign new_n10696 = ~new_n10631 & ~new_n10694;
  assign new_n10697 = ~new_n10695_1 & ~new_n10696;
  assign new_n10698 = n5319 & n10848;
  assign new_n10699 = n8028 & n9457;
  assign new_n10700 = n1980 & n5767;
  assign new_n10701 = ~new_n10699 & ~new_n10700;
  assign new_n10702 = new_n10699 & new_n10700;
  assign new_n10703 = ~new_n10701 & ~new_n10702;
  assign new_n10704 = ~new_n10698 & ~new_n10703;
  assign new_n10705 = new_n10698 & new_n10703;
  assign new_n10706 = ~new_n10704 & ~new_n10705;
  assign new_n10707 = new_n10697 & ~new_n10706;
  assign new_n10708 = ~new_n10697 & new_n10706;
  assign new_n10709 = ~new_n10707 & ~new_n10708;
  assign new_n10710 = new_n10693 & new_n10709;
  assign new_n10711 = ~new_n10693 & ~new_n10709;
  assign new_n10712 = ~new_n10710 & ~new_n10711;
  assign new_n10713 = ~new_n10681 & new_n10712;
  assign new_n10714 = new_n10681 & ~new_n10712;
  assign new_n10715 = ~new_n10713 & ~new_n10714;
  assign new_n10716 = ~new_n10651 & ~new_n10715;
  assign new_n10717 = new_n10651 & new_n10715;
  assign new_n10718 = ~new_n10716 & ~new_n10717;
  assign new_n10719 = ~new_n10676 & new_n10718;
  assign new_n10720 = new_n10676 & ~new_n10718;
  assign new_n10721 = ~new_n10719 & ~new_n10720;
  assign new_n10722 = n5069 & n12069;
  assign new_n10723 = n6806 & n12069;
  assign new_n10724 = n2802 & n12391;
  assign new_n10725 = n1564 & n7160;
  assign new_n10726 = n533 & n12391;
  assign new_n10727 = new_n10725 & new_n10726;
  assign new_n10728 = ~new_n10725 & ~new_n10726;
  assign new_n10729 = n1512 & n7891;
  assign new_n10730 = ~new_n10728 & new_n10729;
  assign new_n10731 = ~new_n10727 & ~new_n10730;
  assign new_n10732 = new_n10724 & ~new_n10731;
  assign new_n10733 = ~new_n10724 & new_n10731;
  assign new_n10734 = ~new_n10732 & ~new_n10733;
  assign new_n10735 = n533 & n7891;
  assign new_n10736 = n1564 & n4828;
  assign new_n10737 = n1512 & n7160;
  assign new_n10738 = ~new_n10736 & ~new_n10737;
  assign new_n10739 = n1512 & n4828;
  assign new_n10740 = new_n10725 & new_n10739;
  assign new_n10741 = ~new_n10738 & ~new_n10740;
  assign new_n10742 = ~new_n10735 & ~new_n10741;
  assign new_n10743 = new_n10735 & new_n10741;
  assign new_n10744 = ~new_n10742 & ~new_n10743;
  assign new_n10745 = ~new_n10734 & ~new_n10744;
  assign new_n10746 = new_n10734 & new_n10744;
  assign new_n10747 = ~new_n10745 & ~new_n10746;
  assign new_n10748 = new_n10723 & new_n10747;
  assign new_n10749 = ~new_n10723 & ~new_n10747;
  assign new_n10750 = n2802 & n12069;
  assign new_n10751 = n1512 & n12391;
  assign new_n10752 = n1564 & n7891;
  assign new_n10753 = n533 & n12069;
  assign new_n10754 = ~new_n10752 & ~new_n10753;
  assign new_n10755 = new_n10751 & ~new_n10754;
  assign new_n10756 = new_n380 & new_n10735;
  assign new_n10757 = ~new_n10755 & ~new_n10756;
  assign new_n10758 = ~new_n10750 & new_n10757;
  assign new_n10759 = new_n10750 & ~new_n10757;
  assign new_n10760 = ~new_n10727 & ~new_n10728;
  assign new_n10761 = ~new_n10729 & ~new_n10760;
  assign new_n10762 = new_n10729 & new_n10760;
  assign new_n10763 = ~new_n10761 & ~new_n10762;
  assign new_n10764 = ~new_n10759 & ~new_n10763;
  assign new_n10765 = ~new_n10758 & ~new_n10764;
  assign new_n10766 = ~new_n10749 & new_n10765;
  assign new_n10767 = ~new_n10748 & ~new_n10766;
  assign new_n10768 = n2802 & n7891;
  assign new_n10769 = n6806 & n12391;
  assign new_n10770 = ~new_n10768 & ~new_n10769;
  assign new_n10771 = new_n10768 & new_n10769;
  assign new_n10772 = ~new_n10770 & ~new_n10771;
  assign new_n10773 = n533 & n7160;
  assign new_n10774 = n1564 & n2515;
  assign new_n10775 = ~new_n10739 & ~new_n10774;
  assign new_n10776 = new_n10739 & new_n10774;
  assign new_n10777 = ~new_n10775 & ~new_n10776;
  assign new_n10778 = ~new_n10773 & ~new_n10777;
  assign new_n10779 = new_n10773 & new_n10777;
  assign new_n10780 = ~new_n10778 & ~new_n10779;
  assign new_n10781 = new_n10735 & ~new_n10738;
  assign new_n10782 = ~new_n10740 & ~new_n10781;
  assign new_n10783 = ~new_n10780 & new_n10782;
  assign new_n10784 = new_n10780 & ~new_n10782;
  assign new_n10785 = ~new_n10783 & ~new_n10784;
  assign new_n10786 = new_n10772 & new_n10785;
  assign new_n10787 = ~new_n10772 & ~new_n10785;
  assign new_n10788 = ~new_n10786 & ~new_n10787;
  assign new_n10789_1 = ~new_n10732 & ~new_n10744;
  assign new_n10790 = ~new_n10733 & ~new_n10789_1;
  assign new_n10791 = ~new_n10788 & new_n10790;
  assign new_n10792 = new_n10788 & ~new_n10790;
  assign new_n10793 = ~new_n10791 & ~new_n10792;
  assign new_n10794 = ~new_n10767 & ~new_n10793;
  assign new_n10795 = new_n10767 & new_n10793;
  assign new_n10796 = ~new_n10794 & ~new_n10795;
  assign new_n10797 = new_n10722 & new_n10796;
  assign new_n10798 = ~new_n10754 & ~new_n10756;
  assign new_n10799 = n1564 & n12391;
  assign new_n10800 = n1512 & n12069;
  assign new_n10801 = new_n10799 & new_n10800;
  assign new_n10802 = ~new_n10798 & new_n10801;
  assign new_n10803 = ~new_n10758 & ~new_n10759;
  assign new_n10804 = new_n10763 & ~new_n10803;
  assign new_n10805 = ~new_n10763 & new_n10803;
  assign new_n10806 = ~new_n10804 & ~new_n10805;
  assign new_n10807 = new_n10802 & ~new_n10806;
  assign new_n10808 = ~new_n10748 & ~new_n10749;
  assign new_n10809 = new_n10765 & new_n10808;
  assign new_n10810 = ~new_n10765 & ~new_n10808;
  assign new_n10811 = ~new_n10809 & ~new_n10810;
  assign new_n10812 = new_n10807 & new_n10811;
  assign new_n10813 = ~new_n10722 & ~new_n10796;
  assign new_n10814 = ~new_n10797 & ~new_n10813;
  assign new_n10815 = new_n10812 & new_n10814;
  assign new_n10816 = ~new_n10797 & ~new_n10815;
  assign new_n10817 = ~new_n10787 & new_n10790;
  assign new_n10818 = ~new_n10771 & ~new_n10817;
  assign new_n10819 = ~new_n10786 & new_n10818;
  assign new_n10820 = new_n10771 & new_n10817;
  assign new_n10821 = ~new_n10819 & ~new_n10820;
  assign new_n10822 = n5069 & n12391;
  assign new_n10823 = n6806 & n7891;
  assign new_n10824 = n12044 & n12069;
  assign new_n10825 = ~new_n10823 & ~new_n10824;
  assign new_n10826 = new_n10823 & new_n10824;
  assign new_n10827 = ~new_n10825 & ~new_n10826;
  assign new_n10828 = ~new_n10822 & ~new_n10827;
  assign new_n10829 = new_n10822 & new_n10827;
  assign new_n10830 = ~new_n10828 & ~new_n10829;
  assign new_n10831 = ~new_n10779 & new_n10782;
  assign new_n10832 = ~new_n10778 & ~new_n10831;
  assign new_n10833 = new_n10830 & new_n10832;
  assign new_n10834 = ~new_n10830 & ~new_n10832;
  assign new_n10835 = ~new_n10833 & ~new_n10834;
  assign new_n10836 = n2802 & n7160;
  assign new_n10837 = new_n10776 & new_n10836;
  assign new_n10838 = ~new_n10776 & ~new_n10836;
  assign new_n10839 = ~new_n10837 & ~new_n10838;
  assign new_n10840 = n1199 & n1564;
  assign new_n10841 = n1512 & n2515;
  assign new_n10842 = n533 & n4828;
  assign new_n10843 = ~new_n10841 & ~new_n10842;
  assign new_n10844 = new_n10841 & new_n10842;
  assign new_n10845 = ~new_n10843 & ~new_n10844;
  assign new_n10846 = new_n10840 & ~new_n10845;
  assign new_n10847 = ~new_n10840 & new_n10845;
  assign new_n10848_1 = ~new_n10846 & ~new_n10847;
  assign new_n10849 = new_n10839 & new_n10848_1;
  assign new_n10850 = ~new_n10839 & ~new_n10848_1;
  assign new_n10851_1 = ~new_n10849 & ~new_n10850;
  assign new_n10852 = ~new_n10835 & new_n10851_1;
  assign new_n10853 = new_n10835 & ~new_n10851_1;
  assign new_n10854 = ~new_n10852 & ~new_n10853;
  assign new_n10855 = new_n10821 & ~new_n10854;
  assign new_n10856 = ~new_n10821 & new_n10854;
  assign new_n10857 = ~new_n10855 & ~new_n10856;
  assign new_n10858 = ~new_n10794 & new_n10857;
  assign new_n10859 = new_n10794 & ~new_n10857;
  assign new_n10860 = ~new_n10858 & ~new_n10859;
  assign new_n10861 = ~new_n10816 & new_n10860;
  assign new_n10862 = new_n10816 & ~new_n10860;
  assign new_n10863 = ~new_n10861 & ~new_n10862;
  assign new_n10864 = ~new_n10672 & ~new_n10674;
  assign new_n10865 = ~new_n10675 & ~new_n10864;
  assign new_n10866 = ~new_n10812 & ~new_n10814;
  assign new_n10867 = ~new_n10815 & ~new_n10866;
  assign new_n10868 = new_n10865 & new_n10867;
  assign new_n10869 = ~new_n10865 & ~new_n10867;
  assign new_n10870 = ~new_n10667 & ~new_n10671;
  assign new_n10871 = ~new_n10672 & ~new_n10870;
  assign new_n10872 = ~new_n10802 & new_n10806;
  assign new_n10873 = ~new_n10807 & ~new_n10872;
  assign new_n10874 = ~new_n10662 & new_n10666;
  assign new_n10875 = ~new_n10667 & ~new_n10874;
  assign new_n10876 = new_n10873 & new_n10875;
  assign new_n10877 = ~new_n10873 & ~new_n10875;
  assign new_n10878 = ~new_n10657 & new_n10661;
  assign new_n10879 = ~new_n10662 & ~new_n10878;
  assign new_n10880 = ~new_n380 & new_n10751;
  assign new_n10881 = ~new_n10798 & ~new_n10880;
  assign new_n10882 = ~new_n10754 & new_n10880;
  assign new_n10883 = ~new_n10881 & ~new_n10882;
  assign new_n10884 = ~new_n10879 & ~new_n10883;
  assign new_n10885 = new_n10879 & new_n10883;
  assign new_n10886 = ~new_n10655 & ~new_n10656;
  assign new_n10887 = ~new_n10657 & ~new_n10886;
  assign new_n10888 = new_n381_1 & new_n10887;
  assign new_n10889 = ~new_n381_1 & ~new_n10887;
  assign new_n10890 = ~new_n10799 & ~new_n10800;
  assign new_n10891 = ~new_n10801 & ~new_n10890;
  assign new_n10892 = ~new_n10889 & new_n10891;
  assign new_n10893 = ~new_n10888 & ~new_n10892;
  assign new_n10894 = ~new_n10885 & new_n10893;
  assign new_n10895 = ~new_n10884 & ~new_n10894;
  assign new_n10896 = ~new_n10877 & new_n10895;
  assign new_n10897 = ~new_n10876 & ~new_n10896;
  assign new_n10898_1 = new_n10871 & ~new_n10897;
  assign new_n10899 = ~new_n10871 & new_n10897;
  assign new_n10900 = ~new_n10807 & ~new_n10811;
  assign new_n10901 = ~new_n10812 & ~new_n10900;
  assign new_n10902 = ~new_n10899 & new_n10901;
  assign new_n10903 = ~new_n10898_1 & ~new_n10902;
  assign new_n10904 = ~new_n10869 & ~new_n10903;
  assign new_n10905 = ~new_n10868 & ~new_n10904;
  assign new_n10906 = ~new_n10863 & new_n10905;
  assign new_n10907 = new_n10863 & ~new_n10905;
  assign new_n10908 = ~new_n10906 & ~new_n10907;
  assign new_n10909 = ~new_n10721 & ~new_n10908;
  assign new_n10910 = new_n10721 & ~new_n10906;
  assign new_n10911 = ~new_n10907 & new_n10910;
  assign new_n10912 = ~new_n10909 & ~new_n10911;
  assign new_n10913_1 = new_n10576 & new_n10912;
  assign new_n10914 = ~new_n10576 & ~new_n10912;
  assign new_n10915 = ~new_n10913_1 & ~new_n10914;
  assign new_n10916 = ~new_n10525 & ~new_n10527;
  assign new_n10917 = ~new_n10528 & ~new_n10916;
  assign new_n10918 = ~new_n10868 & ~new_n10869;
  assign new_n10919 = new_n10903 & ~new_n10918;
  assign new_n10920 = ~new_n10903 & new_n10918;
  assign new_n10921 = ~new_n10919 & ~new_n10920;
  assign new_n10922 = ~new_n10917 & ~new_n10921;
  assign new_n10923 = new_n10917 & new_n10921;
  assign new_n10924 = ~new_n10520 & ~new_n10524;
  assign new_n10925 = ~new_n10525 & ~new_n10924;
  assign new_n10926 = ~new_n10898_1 & ~new_n10899;
  assign new_n10927 = ~new_n10901 & ~new_n10926;
  assign new_n10928_1 = new_n10901 & new_n10926;
  assign new_n10929 = ~new_n10927 & ~new_n10928_1;
  assign new_n10930 = ~new_n10925 & ~new_n10929;
  assign new_n10931 = new_n10925 & new_n10929;
  assign new_n10932 = ~new_n10515 & new_n10519;
  assign new_n10933 = ~new_n10520 & ~new_n10932;
  assign new_n10934 = ~new_n10876 & ~new_n10877;
  assign new_n10935 = ~new_n10895 & ~new_n10934;
  assign new_n10936 = new_n10895 & new_n10934;
  assign new_n10937 = ~new_n10935 & ~new_n10936;
  assign new_n10938 = ~new_n10933 & ~new_n10937;
  assign new_n10939 = new_n10933 & new_n10937;
  assign new_n10940 = ~new_n10884 & ~new_n10885;
  assign new_n10941 = ~new_n10893 & ~new_n10940;
  assign new_n10942 = ~new_n10884 & new_n10894;
  assign new_n10943 = ~new_n10941 & ~new_n10942;
  assign new_n10944 = ~new_n378 & new_n10484;
  assign new_n10945 = ~new_n10511 & ~new_n10944;
  assign new_n10946 = ~new_n10487 & new_n10944;
  assign new_n10947 = ~new_n10945 & ~new_n10946;
  assign new_n10948 = ~new_n10943 & new_n10947;
  assign new_n10949_1 = new_n10943 & ~new_n10947;
  assign new_n10950 = ~new_n10512 & ~new_n10513;
  assign new_n10951 = ~new_n10514 & ~new_n10950;
  assign new_n10952 = ~new_n10888 & ~new_n10889;
  assign new_n10953 = new_n10891 & ~new_n10952;
  assign new_n10954 = ~new_n10891 & new_n10952;
  assign new_n10955 = ~new_n10953 & ~new_n10954;
  assign new_n10956 = new_n10951 & ~new_n10955;
  assign new_n10957 = ~new_n10951 & new_n10955;
  assign new_n10958 = new_n384 & ~new_n10957;
  assign new_n10959 = ~new_n10956 & ~new_n10958;
  assign new_n10960 = ~new_n10949_1 & ~new_n10959;
  assign new_n10961 = ~new_n10948 & ~new_n10960;
  assign new_n10962 = ~new_n10939 & new_n10961;
  assign new_n10963 = ~new_n10938 & ~new_n10962;
  assign new_n10964 = ~new_n10931 & ~new_n10963;
  assign new_n10965_1 = ~new_n10930 & ~new_n10964;
  assign new_n10966 = ~new_n10923 & ~new_n10965_1;
  assign new_n10967 = ~new_n10922 & ~new_n10966;
  assign new_n10968 = ~new_n10915 & new_n10967;
  assign new_n10969 = new_n10915 & ~new_n10967;
  assign new_n10970 = ~new_n10968 & ~new_n10969;
  assign new_n10971 = ~new_n10434 & new_n10970;
  assign new_n10972 = new_n10434 & ~new_n10970;
  assign new_n10973 = ~new_n10381 & ~new_n10383;
  assign new_n10974 = ~new_n10384 & ~new_n10973;
  assign new_n10975 = ~new_n10376 & new_n10380;
  assign new_n10976 = ~new_n10381 & ~new_n10975;
  assign new_n10977 = ~new_n10930 & ~new_n10931;
  assign new_n10978 = new_n10963 & ~new_n10977;
  assign new_n10979 = ~new_n10963 & new_n10977;
  assign new_n10980 = ~new_n10978 & ~new_n10979;
  assign new_n10981 = new_n10976 & ~new_n10980;
  assign new_n10982 = ~new_n10976 & new_n10980;
  assign new_n10983 = ~new_n10371 & new_n10375;
  assign new_n10984 = ~new_n10376 & ~new_n10983;
  assign new_n10985 = ~new_n10938 & ~new_n10939;
  assign new_n10986 = new_n10961 & new_n10985;
  assign new_n10987 = ~new_n10961 & ~new_n10985;
  assign new_n10988 = ~new_n10986 & ~new_n10987;
  assign new_n10989 = new_n10984 & ~new_n10988;
  assign new_n10990_1 = ~new_n10984 & new_n10988;
  assign new_n10991 = ~new_n10366 & ~new_n10370;
  assign new_n10992 = ~new_n10371 & ~new_n10991;
  assign new_n10993 = ~new_n10948 & ~new_n10949_1;
  assign new_n10994 = new_n10959 & ~new_n10993;
  assign new_n10995 = ~new_n10959 & new_n10993;
  assign new_n10996 = ~new_n10994 & ~new_n10995;
  assign new_n10997 = new_n10992 & new_n10996;
  assign new_n10998 = ~new_n10992 & ~new_n10996;
  assign new_n10999 = ~new_n10364 & ~new_n10365;
  assign new_n11000 = ~new_n10366 & ~new_n10999;
  assign new_n11001 = new_n387 & new_n11000;
  assign new_n11002 = ~new_n387 & ~new_n11000;
  assign new_n11003 = ~new_n10956 & ~new_n10957;
  assign new_n11004 = ~new_n384 & ~new_n11003;
  assign new_n11005 = new_n384 & new_n11003;
  assign new_n11006 = ~new_n11004 & ~new_n11005;
  assign new_n11007 = ~new_n11002 & new_n11006;
  assign new_n11008 = ~new_n11001 & ~new_n11007;
  assign new_n11009 = ~new_n10998 & ~new_n11008;
  assign new_n11010 = ~new_n10997 & ~new_n11009;
  assign new_n11011 = ~new_n10990_1 & ~new_n11010;
  assign new_n11012 = ~new_n10989 & ~new_n11011;
  assign new_n11013 = ~new_n10982 & ~new_n11012;
  assign new_n11014 = ~new_n10981 & ~new_n11013;
  assign new_n11015 = ~new_n10974 & new_n11014;
  assign new_n11016 = new_n10974 & ~new_n11014;
  assign new_n11017 = ~new_n10922 & ~new_n10923;
  assign new_n11018 = ~new_n10965_1 & ~new_n11017;
  assign new_n11019 = new_n10965_1 & new_n11017;
  assign new_n11020 = ~new_n11018 & ~new_n11019;
  assign new_n11021 = ~new_n11016 & ~new_n11020;
  assign new_n11022 = ~new_n11015 & ~new_n11021;
  assign new_n11023_1 = ~new_n10972 & ~new_n11022;
  assign new_n11024 = ~new_n10971 & ~new_n11023_1;
  assign new_n11025 = ~new_n10907 & ~new_n10910;
  assign new_n11026 = ~new_n10571 & ~new_n10574;
  assign new_n11027 = n4005 & n4189;
  assign new_n11028 = n2508 & n9920;
  assign new_n11029 = n2564 & n12706;
  assign new_n11030 = ~new_n11028 & new_n11029;
  assign new_n11031 = new_n11028 & ~new_n11029;
  assign new_n11032 = ~new_n11030 & ~new_n11031;
  assign new_n11033 = new_n11027 & ~new_n11032;
  assign new_n11034 = ~new_n11027 & new_n11032;
  assign new_n11035 = ~new_n11033 & ~new_n11034;
  assign new_n11036 = n2585 & n6770;
  assign new_n11037 = n3627 & n12720;
  assign new_n11038 = n2509 & n4516;
  assign new_n11039 = ~new_n11037 & new_n11038;
  assign new_n11040 = new_n11037 & ~new_n11038;
  assign new_n11041 = ~new_n11039 & ~new_n11040;
  assign new_n11042 = new_n11036 & new_n11041;
  assign new_n11043 = ~new_n11036 & ~new_n11041;
  assign new_n11044 = ~new_n11042 & ~new_n11043;
  assign new_n11045 = new_n10407 & ~new_n10410;
  assign new_n11046 = ~new_n10411 & ~new_n11045;
  assign new_n11047 = ~new_n11044 & ~new_n11046;
  assign new_n11048 = new_n11044 & new_n11046;
  assign new_n11049 = ~new_n11047 & ~new_n11048;
  assign new_n11050 = ~new_n11035 & ~new_n11049;
  assign new_n11051 = new_n11035 & new_n11049;
  assign new_n11052 = ~new_n11050 & ~new_n11051;
  assign new_n11053 = ~new_n10405 & ~new_n10415;
  assign new_n11054 = ~new_n10404 & ~new_n11053;
  assign new_n11055 = ~new_n10391_1 & ~new_n10395;
  assign new_n11056 = ~new_n10394 & ~new_n11055;
  assign new_n11057 = ~new_n11054 & new_n11056;
  assign new_n11058 = new_n11054 & ~new_n11056;
  assign new_n11059 = ~new_n11057 & ~new_n11058;
  assign new_n11060 = new_n11052 & new_n11059;
  assign new_n11061 = ~new_n11052 & ~new_n11059;
  assign new_n11062 = ~new_n11060 & ~new_n11061;
  assign new_n11063 = ~new_n10422 & new_n11062;
  assign new_n11064 = new_n10422 & ~new_n11062;
  assign new_n11065 = ~new_n11063 & ~new_n11064;
  assign new_n11066 = new_n11026 & new_n11065;
  assign new_n11067 = ~new_n11026 & ~new_n11065;
  assign new_n11068 = ~new_n11066 & ~new_n11067;
  assign new_n11069 = new_n11025 & new_n11068;
  assign new_n11070 = ~new_n11025 & ~new_n11068;
  assign new_n11071 = ~new_n11069 & ~new_n11070;
  assign new_n11072 = ~new_n10679 & ~new_n10712;
  assign new_n11073 = ~new_n10680 & ~new_n11072;
  assign new_n11074 = n1980 & n5319;
  assign new_n11075 = n9457 & n10848;
  assign new_n11076 = ~new_n11074 & ~new_n11075;
  assign new_n11077 = new_n11074 & new_n11075;
  assign new_n11078 = ~new_n11076 & ~new_n11077;
  assign new_n11079 = n1906 & n11222;
  assign new_n11080 = n4817 & n8028;
  assign new_n11081 = new_n11079 & ~new_n11080;
  assign new_n11082 = ~new_n11079 & new_n11080;
  assign new_n11083 = ~new_n11081 & ~new_n11082;
  assign new_n11084 = ~new_n11078 & ~new_n11083;
  assign new_n11085 = new_n11078 & new_n11083;
  assign new_n11086 = ~new_n11084 & ~new_n11085;
  assign new_n11087 = ~new_n11073 & ~new_n11086;
  assign new_n11088 = new_n11073 & new_n11086;
  assign new_n11089 = ~new_n11087 & ~new_n11088;
  assign new_n11090 = ~new_n10692 & ~new_n10709;
  assign new_n11091 = ~new_n10691 & ~new_n11090;
  assign new_n11092 = ~new_n10695_1 & ~new_n10706;
  assign new_n11093 = ~new_n10696 & ~new_n11092;
  assign new_n11094 = new_n11091 & new_n11093;
  assign new_n11095 = ~new_n11091 & ~new_n11093;
  assign new_n11096 = ~new_n11094 & ~new_n11095;
  assign new_n11097 = n1564 & n6578;
  assign new_n11098 = n4903 & n11153;
  assign new_n11099 = n996 & n12704;
  assign new_n11100 = n5767 & n7294;
  assign new_n11101 = ~new_n11099 & new_n11100;
  assign new_n11102 = new_n11099 & ~new_n11100;
  assign new_n11103 = ~new_n11101 & ~new_n11102;
  assign new_n11104 = new_n11098 & new_n11103;
  assign new_n11105 = ~new_n11098 & ~new_n11103;
  assign new_n11106 = ~new_n11104 & ~new_n11105;
  assign new_n11107 = ~new_n10682 & ~new_n10686;
  assign new_n11108 = ~new_n10685_1 & ~new_n11107;
  assign new_n11109 = ~new_n11106 & new_n11108;
  assign new_n11110 = new_n11106 & ~new_n11108;
  assign new_n11111 = ~new_n11109 & ~new_n11110;
  assign new_n11112 = ~new_n10698 & ~new_n10702;
  assign new_n11113 = ~new_n10701 & ~new_n11112;
  assign new_n11114 = n5694 & n12069;
  assign new_n11115 = n5314 & n5814;
  assign new_n11116 = new_n11114 & ~new_n11115;
  assign new_n11117 = ~new_n11114 & new_n11115;
  assign new_n11118 = ~new_n11116 & ~new_n11117;
  assign new_n11119 = ~new_n11113 & ~new_n11118;
  assign new_n11120 = new_n11113 & new_n11118;
  assign new_n11121 = ~new_n11119 & ~new_n11120;
  assign new_n11122 = ~new_n11111 & new_n11121;
  assign new_n11123 = new_n11111 & ~new_n11121;
  assign new_n11124 = ~new_n11122 & ~new_n11123;
  assign new_n11125 = ~new_n11097 & new_n11124;
  assign new_n11126 = new_n11097 & ~new_n11124;
  assign new_n11127 = ~new_n11125 & ~new_n11126;
  assign new_n11128 = new_n11096 & ~new_n11127;
  assign new_n11129 = ~new_n11096 & new_n11127;
  assign new_n11130 = ~new_n11128 & ~new_n11129;
  assign new_n11131 = ~new_n10717 & ~new_n10719;
  assign new_n11132 = ~new_n10535 & ~new_n10539;
  assign new_n11133 = ~new_n10538 & ~new_n11132;
  assign new_n11134 = n1094 & n5105;
  assign new_n11135 = n1209 & n10678;
  assign new_n11136 = ~new_n11134 & new_n11135;
  assign new_n11137 = new_n11134 & ~new_n11135;
  assign new_n11138 = ~new_n11136 & ~new_n11137;
  assign new_n11139 = n4928 & n6986;
  assign new_n11140 = n2226 & n4141;
  assign new_n11141 = new_n11139 & new_n11140;
  assign new_n11142 = ~new_n11139 & ~new_n11140;
  assign new_n11143 = ~new_n11141 & ~new_n11142;
  assign new_n11144 = new_n11138 & ~new_n11143;
  assign new_n11145 = ~new_n11138 & new_n11143;
  assign new_n11146 = ~new_n11144 & ~new_n11145;
  assign new_n11147 = ~new_n11133 & new_n11146;
  assign new_n11148 = new_n11133 & ~new_n11146;
  assign new_n11149 = ~new_n11147 & ~new_n11148;
  assign new_n11150 = n8236 & n10928;
  assign new_n11151 = ~new_n10543 & ~new_n10545_1;
  assign new_n11152 = ~new_n10546 & ~new_n11151;
  assign new_n11153_1 = new_n11150 & new_n11152;
  assign new_n11154 = ~new_n11150 & ~new_n11152;
  assign new_n11155 = ~new_n11153_1 & ~new_n11154;
  assign new_n11156 = new_n11149 & new_n11155;
  assign new_n11157 = ~new_n11149 & ~new_n11155;
  assign new_n11158 = ~new_n11156 & ~new_n11157;
  assign new_n11159 = ~new_n10550 & ~new_n10562;
  assign new_n11160 = ~new_n10563 & ~new_n11159;
  assign new_n11161 = ~new_n10551 & ~new_n10555;
  assign new_n11162 = ~new_n10554 & ~new_n11161;
  assign new_n11163 = ~new_n11160 & new_n11162;
  assign new_n11164 = new_n11160 & ~new_n11162;
  assign new_n11165 = ~new_n11163 & ~new_n11164;
  assign new_n11166 = new_n11158 & new_n11165;
  assign new_n11167 = ~new_n11158 & ~new_n11165;
  assign new_n11168 = ~new_n11166 & ~new_n11167;
  assign new_n11169 = new_n11131 & new_n11168;
  assign new_n11170 = ~new_n11131 & ~new_n11168;
  assign new_n11171 = ~new_n11169 & ~new_n11170;
  assign new_n11172 = new_n11130 & new_n11171;
  assign new_n11173 = ~new_n11130 & ~new_n11171;
  assign new_n11174 = ~new_n11172 & ~new_n11173;
  assign new_n11175 = new_n11089 & ~new_n11174;
  assign new_n11176 = ~new_n11089 & new_n11174;
  assign new_n11177 = ~new_n11175 & ~new_n11176;
  assign new_n11178 = ~new_n11071 & ~new_n11177;
  assign new_n11179 = new_n11071 & new_n11177;
  assign new_n11180 = ~new_n11178 & ~new_n11179;
  assign new_n11181 = ~new_n10913_1 & ~new_n10967;
  assign new_n11182 = ~new_n10914 & ~new_n11181;
  assign new_n11183 = new_n11180 & new_n11182;
  assign new_n11184 = ~new_n11180 & ~new_n11182;
  assign new_n11185 = ~new_n11183 & ~new_n11184;
  assign new_n11186 = ~new_n10429 & ~new_n10432;
  assign new_n11187 = ~new_n10838 & ~new_n10848_1;
  assign new_n11188 = ~new_n10837 & ~new_n11187;
  assign new_n11189 = ~new_n10822 & ~new_n10826;
  assign new_n11190 = ~new_n10825 & ~new_n11189;
  assign new_n11191 = ~new_n11188 & new_n11190;
  assign new_n11192 = new_n11188 & ~new_n11190;
  assign new_n11193 = ~new_n11191 & ~new_n11192;
  assign new_n11194 = n5069 & n7891;
  assign new_n11195 = n12044 & n12391;
  assign new_n11196 = ~new_n11194 & new_n11195;
  assign new_n11197 = new_n11194 & ~new_n11195;
  assign new_n11198 = ~new_n11196 & ~new_n11197;
  assign new_n11199 = ~new_n11193 & new_n11198;
  assign new_n11200 = new_n11193 & ~new_n11198;
  assign new_n11201 = ~new_n11199 & ~new_n11200;
  assign new_n11202 = ~new_n10840 & ~new_n10844;
  assign new_n11203 = ~new_n10843 & ~new_n11202;
  assign new_n11204 = ~new_n10833 & new_n10851_1;
  assign new_n11205 = ~new_n10834 & ~new_n11204;
  assign new_n11206 = new_n11203 & new_n11205;
  assign new_n11207 = ~new_n11203 & ~new_n11205;
  assign new_n11208 = ~new_n11206 & ~new_n11207;
  assign new_n11209 = new_n11201 & new_n11208;
  assign new_n11210 = ~new_n11201 & ~new_n11208;
  assign new_n11211 = ~new_n11209 & ~new_n11210;
  assign new_n11212 = ~new_n10388 & new_n10425;
  assign new_n11213 = ~new_n10389 & ~new_n11212;
  assign new_n11214 = n615 & n6687;
  assign new_n11215 = n2087 & n6038;
  assign new_n11216_1 = ~new_n11214 & new_n11215;
  assign new_n11217 = new_n11214 & ~new_n11215;
  assign new_n11218 = ~new_n11216_1 & ~new_n11217;
  assign new_n11219 = new_n11213 & new_n11218;
  assign new_n11220 = ~new_n11213 & ~new_n11218;
  assign new_n11221 = ~new_n11219 & ~new_n11220;
  assign new_n11222_1 = ~new_n11211 & new_n11221;
  assign new_n11223 = new_n11211 & ~new_n11221;
  assign new_n11224 = ~new_n11222_1 & ~new_n11223;
  assign new_n11225 = ~new_n10819 & new_n10854;
  assign new_n11226 = ~new_n10820 & ~new_n11225;
  assign new_n11227 = n6806 & n7160;
  assign new_n11228 = n2802 & n4828;
  assign new_n11229 = ~new_n11227 & ~new_n11228;
  assign new_n11230 = new_n11227 & new_n11228;
  assign new_n11231 = ~new_n11229 & ~new_n11230;
  assign new_n11232 = n533 & n2515;
  assign new_n11233 = n1199 & n1512;
  assign new_n11234 = new_n11232 & ~new_n11233;
  assign new_n11235 = ~new_n11232 & new_n11233;
  assign new_n11236 = ~new_n11234 & ~new_n11235;
  assign new_n11237 = ~new_n11231 & ~new_n11236;
  assign new_n11238 = new_n11231 & new_n11236;
  assign new_n11239 = ~new_n11237 & ~new_n11238;
  assign new_n11240 = new_n11226 & new_n11239;
  assign new_n11241 = ~new_n11226 & ~new_n11239;
  assign new_n11242 = ~new_n11240 & ~new_n11241;
  assign new_n11243 = ~new_n11224 & new_n11242;
  assign new_n11244 = new_n11224 & ~new_n11242;
  assign new_n11245 = ~new_n11243 & ~new_n11244;
  assign new_n11246 = new_n11186 & new_n11245;
  assign new_n11247 = ~new_n11186 & ~new_n11245;
  assign new_n11248 = ~new_n11246 & ~new_n11247;
  assign new_n11249 = n7320 & n7500;
  assign new_n11250 = n7354 & n7523;
  assign new_n11251 = n783 & n8336;
  assign new_n11252 = ~new_n11250 & new_n11251;
  assign new_n11253 = new_n11250 & ~new_n11251;
  assign new_n11254 = ~new_n11252 & ~new_n11253;
  assign new_n11255 = ~new_n11249 & new_n11254;
  assign new_n11256 = new_n11249 & ~new_n11254;
  assign new_n11257_1 = ~new_n11255 & ~new_n11256;
  assign new_n11258 = ~new_n10859 & ~new_n10861;
  assign new_n11259 = ~new_n10533 & ~new_n10567;
  assign new_n11260 = ~new_n10531 & ~new_n11259;
  assign new_n11261 = new_n11258 & new_n11260;
  assign new_n11262 = ~new_n11258 & ~new_n11260;
  assign new_n11263 = ~new_n11261 & ~new_n11262;
  assign new_n11264 = new_n11257_1 & ~new_n11263;
  assign new_n11265 = ~new_n11257_1 & new_n11263;
  assign new_n11266 = ~new_n11264 & ~new_n11265;
  assign new_n11267 = new_n11248 & new_n11266;
  assign new_n11268 = ~new_n11248 & ~new_n11266;
  assign new_n11269 = ~new_n11267 & ~new_n11268;
  assign new_n11270 = new_n11185 & ~new_n11269;
  assign new_n11271 = ~new_n11185 & new_n11269;
  assign new_n11272 = ~new_n11270 & ~new_n11271;
  assign new_n11273 = ~new_n11024 & ~new_n11272;
  assign new_n11274 = new_n11024 & new_n11272;
  assign n3654 = ~new_n11273 & ~new_n11274;
  assign new_n11276 = ~new_n11015 & ~new_n11016;
  assign new_n11277 = new_n11020 & ~new_n11276;
  assign new_n11278 = ~new_n11020 & new_n11276;
  assign n3661 = new_n11277 | new_n11278;
  assign new_n11280 = n6703 & n12299;
  assign new_n11281 = n6776 & n9640;
  assign new_n11282 = n3022 & n8759;
  assign new_n11283 = ~new_n11281 & ~new_n11282;
  assign new_n11284 = new_n11281 & new_n11282;
  assign new_n11285 = ~new_n11283 & ~new_n11284;
  assign new_n11286 = new_n11280 & ~new_n11285;
  assign new_n11287 = ~new_n11280 & new_n11285;
  assign new_n11288 = ~new_n11286 & ~new_n11287;
  assign new_n11289 = new_n7065 & ~new_n11288;
  assign new_n11290 = n8759 & n11023;
  assign new_n11291 = new_n11280 & ~new_n11283;
  assign new_n11292 = ~new_n11284 & ~new_n11291;
  assign new_n11293 = ~new_n11290 & new_n11292;
  assign new_n11294 = new_n11290 & ~new_n11292;
  assign new_n11295 = ~new_n11293 & ~new_n11294;
  assign new_n11296_1 = n6703 & n7436;
  assign new_n11297 = n3022 & n6776;
  assign new_n11298 = n9640 & n12299;
  assign new_n11299 = ~new_n11297 & ~new_n11298;
  assign new_n11300 = new_n11297 & new_n11298;
  assign new_n11301 = ~new_n11299 & ~new_n11300;
  assign new_n11302 = new_n11296_1 & ~new_n11301;
  assign new_n11303 = ~new_n11296_1 & new_n11301;
  assign new_n11304 = ~new_n11302 & ~new_n11303;
  assign new_n11305 = ~new_n11295 & new_n11304;
  assign new_n11306 = new_n11295 & ~new_n11304;
  assign new_n11307 = ~new_n11305 & ~new_n11306;
  assign new_n11308 = new_n11289 & new_n11307;
  assign new_n11309 = n8759 & n10451;
  assign new_n11310 = n6776 & n11023;
  assign new_n11311_1 = new_n11296_1 & ~new_n11299;
  assign new_n11312 = ~new_n11300 & ~new_n11311_1;
  assign new_n11313 = ~new_n11310 & new_n11312;
  assign new_n11314 = new_n11310 & ~new_n11312;
  assign new_n11315 = ~new_n11313 & ~new_n11314;
  assign new_n11316 = n6703 & n8276;
  assign new_n11317 = n3022 & n12299;
  assign new_n11318 = n7436 & n9640;
  assign new_n11319 = ~new_n11317 & ~new_n11318;
  assign new_n11320 = new_n11317 & new_n11318;
  assign new_n11321 = ~new_n11319 & ~new_n11320;
  assign new_n11322 = new_n11316 & ~new_n11321;
  assign new_n11323 = ~new_n11316 & new_n11321;
  assign new_n11324 = ~new_n11322 & ~new_n11323;
  assign new_n11325 = ~new_n11315 & new_n11324;
  assign new_n11326_1 = new_n11315 & ~new_n11324;
  assign new_n11327 = ~new_n11325 & ~new_n11326_1;
  assign new_n11328 = new_n11309 & new_n11327;
  assign new_n11329 = ~new_n11309 & ~new_n11327;
  assign new_n11330 = ~new_n11328 & ~new_n11329;
  assign new_n11331 = ~new_n11293 & ~new_n11304;
  assign new_n11332 = ~new_n11294 & ~new_n11331;
  assign new_n11333 = ~new_n11330 & ~new_n11332;
  assign new_n11334 = new_n11330 & new_n11332;
  assign new_n11335 = ~new_n11333 & ~new_n11334;
  assign new_n11336 = new_n11308 & ~new_n11335;
  assign new_n11337 = ~new_n11308 & new_n11335;
  assign new_n11338 = ~new_n11336 & ~new_n11337;
  assign new_n11339 = n11876 & n11892;
  assign new_n11340 = n7388 & n10898;
  assign new_n11341 = n3754 & n7965;
  assign new_n11342 = ~new_n11340 & ~new_n11341;
  assign new_n11343 = new_n11340 & new_n11341;
  assign new_n11344 = ~new_n11342 & ~new_n11343;
  assign new_n11345 = new_n11339 & ~new_n11344;
  assign new_n11346 = ~new_n11339 & new_n11344;
  assign new_n11347 = ~new_n11345 & ~new_n11346;
  assign new_n11348 = new_n7073 & ~new_n11347;
  assign new_n11349 = n2749 & n7965;
  assign new_n11350 = new_n11339 & ~new_n11342;
  assign new_n11351 = ~new_n11343 & ~new_n11350;
  assign new_n11352 = new_n11349 & ~new_n11351;
  assign new_n11353 = ~new_n11349 & new_n11351;
  assign new_n11354 = ~new_n11352 & ~new_n11353;
  assign new_n11355 = n10898 & n11892;
  assign new_n11356 = n3754 & n7388;
  assign new_n11357 = n2393 & n11876;
  assign new_n11358 = ~new_n11356 & ~new_n11357;
  assign new_n11359 = new_n11356 & new_n11357;
  assign new_n11360 = ~new_n11358 & ~new_n11359;
  assign new_n11361 = new_n11355 & ~new_n11360;
  assign new_n11362 = ~new_n11355 & new_n11360;
  assign new_n11363 = ~new_n11361 & ~new_n11362;
  assign new_n11364 = ~new_n11354 & ~new_n11363;
  assign new_n11365 = new_n11354 & new_n11363;
  assign new_n11366 = ~new_n11364 & ~new_n11365;
  assign new_n11367 = new_n11348 & ~new_n11366;
  assign new_n11368 = n159 & n7965;
  assign new_n11369 = ~new_n11353 & ~new_n11363;
  assign new_n11370 = ~new_n11352 & ~new_n11369;
  assign new_n11371 = ~new_n11368 & new_n11370;
  assign new_n11372 = n2749 & n7388;
  assign new_n11373 = new_n11355 & ~new_n11358;
  assign new_n11374 = ~new_n11359 & ~new_n11373;
  assign new_n11375 = new_n11372 & ~new_n11374;
  assign new_n11376 = ~new_n11372 & new_n11374;
  assign new_n11377 = ~new_n11375 & ~new_n11376;
  assign new_n11378 = n3754 & n11892;
  assign new_n11379 = n5860 & n11876;
  assign new_n11380 = n2393 & n10898;
  assign new_n11381 = ~new_n11379 & ~new_n11380;
  assign new_n11382 = new_n11379 & new_n11380;
  assign new_n11383 = ~new_n11381 & ~new_n11382;
  assign new_n11384 = new_n11378 & ~new_n11383;
  assign new_n11385 = ~new_n11378 & new_n11383;
  assign new_n11386 = ~new_n11384 & ~new_n11385;
  assign new_n11387 = ~new_n11377 & ~new_n11386;
  assign new_n11388 = new_n11377 & new_n11386;
  assign new_n11389 = ~new_n11387 & ~new_n11388;
  assign new_n11390 = new_n11371 & new_n11389;
  assign new_n11391 = new_n11368 & ~new_n11370;
  assign new_n11392 = ~new_n11389 & new_n11391;
  assign new_n11393 = ~new_n11371 & ~new_n11389;
  assign new_n11394 = ~new_n11391 & ~new_n11393;
  assign new_n11395 = ~new_n11392 & ~new_n11394;
  assign new_n11396 = ~new_n11390 & ~new_n11395;
  assign new_n11397 = new_n11367 & new_n11396;
  assign new_n11398 = ~new_n11367 & ~new_n11396;
  assign new_n11399 = ~new_n11397 & ~new_n11398;
  assign new_n11400 = n2530 & n5645;
  assign new_n11401 = n1067 & n8476;
  assign new_n11402 = n5331 & n8665;
  assign new_n11403 = ~new_n11401 & ~new_n11402;
  assign new_n11404 = new_n11401 & new_n11402;
  assign new_n11405 = ~new_n11403 & ~new_n11404;
  assign new_n11406 = new_n11400 & ~new_n11405;
  assign new_n11407_1 = ~new_n11400 & new_n11405;
  assign new_n11408 = ~new_n11406 & ~new_n11407_1;
  assign new_n11409 = new_n7081 & ~new_n11408;
  assign new_n11410 = n5331 & n11922;
  assign new_n11411 = n5645 & n12648;
  assign new_n11412 = n8476 & n8665;
  assign new_n11413 = n1067 & n2530;
  assign new_n11414 = ~new_n11412 & ~new_n11413;
  assign new_n11415 = new_n11412 & new_n11413;
  assign new_n11416 = ~new_n11414 & ~new_n11415;
  assign new_n11417 = new_n11411 & ~new_n11416;
  assign new_n11418 = ~new_n11411 & new_n11416;
  assign new_n11419 = ~new_n11417 & ~new_n11418;
  assign new_n11420 = new_n11410 & ~new_n11419;
  assign new_n11421 = ~new_n11410 & new_n11419;
  assign new_n11422 = ~new_n11420 & ~new_n11421;
  assign new_n11423_1 = ~new_n11400 & ~new_n11404;
  assign new_n11424 = ~new_n11403 & ~new_n11423_1;
  assign new_n11425 = ~new_n11422 & new_n11424;
  assign new_n11426 = new_n11422 & ~new_n11424;
  assign new_n11427 = ~new_n11425 & ~new_n11426;
  assign new_n11428 = new_n11409 & ~new_n11427;
  assign new_n11429 = n2551 & n5331;
  assign new_n11430 = n8476 & n11922;
  assign new_n11431 = new_n11411 & ~new_n11414;
  assign new_n11432 = ~new_n11415 & ~new_n11431;
  assign new_n11433 = ~new_n11430 & new_n11432;
  assign new_n11434 = new_n11430 & ~new_n11432;
  assign new_n11435 = ~new_n11433 & ~new_n11434;
  assign new_n11436 = n5645 & n10545;
  assign new_n11437 = n2530 & n8665;
  assign new_n11438 = n1067 & n12648;
  assign new_n11439 = ~new_n11437 & ~new_n11438;
  assign new_n11440 = new_n11437 & new_n11438;
  assign new_n11441 = ~new_n11439 & ~new_n11440;
  assign new_n11442 = new_n11436 & ~new_n11441;
  assign new_n11443 = ~new_n11436 & new_n11441;
  assign new_n11444 = ~new_n11442 & ~new_n11443;
  assign new_n11445 = ~new_n11435 & new_n11444;
  assign new_n11446 = new_n11435 & ~new_n11444;
  assign new_n11447 = ~new_n11445 & ~new_n11446;
  assign new_n11448 = new_n11429 & new_n11447;
  assign new_n11449 = ~new_n11429 & ~new_n11447;
  assign new_n11450 = ~new_n11448 & ~new_n11449;
  assign new_n11451 = ~new_n11420 & ~new_n11424;
  assign new_n11452 = ~new_n11421 & ~new_n11451;
  assign new_n11453 = ~new_n11450 & new_n11452;
  assign new_n11454 = new_n11450 & ~new_n11452;
  assign new_n11455 = ~new_n11453 & ~new_n11454;
  assign new_n11456 = new_n11428 & ~new_n11455;
  assign new_n11457 = ~new_n11428 & new_n11455;
  assign new_n11458 = ~new_n11456 & ~new_n11457;
  assign new_n11459 = new_n11399 & new_n11458;
  assign new_n11460 = ~new_n11399 & ~new_n11458;
  assign new_n11461 = ~new_n11459 & ~new_n11460;
  assign new_n11462 = ~new_n11409 & new_n11427;
  assign new_n11463 = ~new_n11428 & ~new_n11462;
  assign new_n11464 = ~new_n11348 & new_n11366;
  assign new_n11465 = ~new_n11367 & ~new_n11464;
  assign new_n11466 = new_n11463 & new_n11465;
  assign new_n11467 = ~new_n11463 & ~new_n11465;
  assign new_n11468 = ~new_n7073 & new_n11347;
  assign new_n11469 = ~new_n11348 & ~new_n11468;
  assign new_n11470 = ~new_n7076 & new_n7082;
  assign new_n11471 = ~new_n7075 & ~new_n11470;
  assign new_n11472 = new_n11469 & ~new_n11471;
  assign new_n11473 = ~new_n11469 & new_n11471;
  assign new_n11474 = ~new_n7081 & new_n11408;
  assign new_n11475 = ~new_n11409 & ~new_n11474;
  assign new_n11476 = ~new_n11473 & new_n11475;
  assign new_n11477 = ~new_n11472 & ~new_n11476;
  assign new_n11478_1 = ~new_n11467 & ~new_n11477;
  assign new_n11479 = ~new_n11466 & ~new_n11478_1;
  assign new_n11480 = new_n11461 & new_n11479;
  assign new_n11481 = ~new_n11461 & ~new_n11479;
  assign new_n11482 = ~new_n11480 & ~new_n11481;
  assign new_n11483 = new_n11338 & ~new_n11482;
  assign new_n11484 = ~new_n11338 & new_n11482;
  assign new_n11485 = ~new_n11483 & ~new_n11484;
  assign new_n11486 = ~new_n11289 & ~new_n11307;
  assign new_n11487 = ~new_n11308 & ~new_n11486;
  assign new_n11488 = ~new_n11466 & ~new_n11467;
  assign new_n11489 = ~new_n11477 & ~new_n11488;
  assign new_n11490 = new_n11477 & new_n11488;
  assign new_n11491 = ~new_n11489 & ~new_n11490;
  assign new_n11492 = new_n11487 & ~new_n11491;
  assign new_n11493 = ~new_n11487 & new_n11491;
  assign new_n11494 = ~new_n7065 & new_n11288;
  assign new_n11495 = ~new_n11289 & ~new_n11494;
  assign new_n11496 = ~new_n7068 & ~new_n7085;
  assign new_n11497 = ~new_n7067 & ~new_n11496;
  assign new_n11498 = new_n11495 & ~new_n11497;
  assign new_n11499 = ~new_n11495 & new_n11497;
  assign new_n11500 = ~new_n11472 & ~new_n11473;
  assign new_n11501 = new_n11475 & new_n11500;
  assign new_n11502 = ~new_n11475 & ~new_n11500;
  assign new_n11503 = ~new_n11501 & ~new_n11502;
  assign new_n11504 = ~new_n11499 & new_n11503;
  assign new_n11505 = ~new_n11498 & ~new_n11504;
  assign new_n11506 = ~new_n11493 & ~new_n11505;
  assign new_n11507 = ~new_n11492 & ~new_n11506;
  assign new_n11508 = new_n11485 & new_n11507;
  assign new_n11509 = ~new_n11485 & ~new_n11507;
  assign new_n11510 = ~new_n11508 & ~new_n11509;
  assign new_n11511 = n1097 & n1798;
  assign new_n11512 = n5305 & n12591;
  assign new_n11513 = ~new_n11511 & ~new_n11512;
  assign new_n11514 = n1097 & n12591;
  assign new_n11515 = new_n7043 & new_n11514;
  assign new_n11516 = ~new_n11513 & ~new_n11515;
  assign new_n11517 = new_n7057 & ~new_n11516;
  assign new_n11518 = n5305 & n7456;
  assign new_n11519 = n3932 & n5964;
  assign new_n11520 = ~new_n11513 & new_n11519;
  assign new_n11521 = ~new_n11515 & ~new_n11520;
  assign new_n11522 = new_n11518 & ~new_n11521;
  assign new_n11523 = ~new_n11518 & new_n11521;
  assign new_n11524 = ~new_n11522 & ~new_n11523;
  assign new_n11525 = n1097 & n3932;
  assign new_n11526 = n1798 & n4312;
  assign new_n11527 = n5964 & n12591;
  assign new_n11528 = ~new_n11526 & ~new_n11527;
  assign new_n11529 = new_n11526 & new_n11527;
  assign new_n11530 = ~new_n11528 & ~new_n11529;
  assign new_n11531 = new_n11525 & ~new_n11530;
  assign new_n11532 = ~new_n11525 & new_n11530;
  assign new_n11533 = ~new_n11531 & ~new_n11532;
  assign new_n11534 = ~new_n11524 & ~new_n11533;
  assign new_n11535 = new_n11524 & new_n11533;
  assign new_n11536_1 = ~new_n11534 & ~new_n11535;
  assign new_n11537 = new_n11517 & ~new_n11536_1;
  assign new_n11538 = n5305 & n11662;
  assign new_n11539 = n5964 & n7456;
  assign new_n11540 = n3932 & n4312;
  assign new_n11541 = n1798 & n12705;
  assign new_n11542 = ~new_n11514 & ~new_n11541;
  assign new_n11543 = n12591 & n12705;
  assign new_n11544 = new_n11511 & new_n11543;
  assign new_n11545 = ~new_n11542 & ~new_n11544;
  assign new_n11546 = ~new_n11540 & new_n11545;
  assign new_n11547 = new_n11540 & ~new_n11545;
  assign new_n11548 = ~new_n11546 & ~new_n11547;
  assign new_n11549 = new_n11539 & ~new_n11548;
  assign new_n11550 = ~new_n11539 & new_n11548;
  assign new_n11551 = ~new_n11549 & ~new_n11550;
  assign new_n11552 = new_n11525 & ~new_n11528;
  assign new_n11553 = ~new_n11529 & ~new_n11552;
  assign new_n11554 = ~new_n11551 & ~new_n11553;
  assign new_n11555 = new_n11551 & new_n11553;
  assign new_n11556 = ~new_n11554 & ~new_n11555;
  assign new_n11557 = new_n11538 & ~new_n11556;
  assign new_n11558 = ~new_n11538 & new_n11556;
  assign new_n11559 = ~new_n11557 & ~new_n11558;
  assign new_n11560 = ~new_n11523 & ~new_n11533;
  assign new_n11561 = ~new_n11522 & ~new_n11560;
  assign new_n11562 = ~new_n11559 & ~new_n11561;
  assign new_n11563 = new_n11559 & new_n11561;
  assign new_n11564 = ~new_n11562 & ~new_n11563;
  assign new_n11565 = new_n11537 & ~new_n11564;
  assign new_n11566 = ~new_n11537 & new_n11564;
  assign new_n11567 = ~new_n11565 & ~new_n11566;
  assign new_n11568 = ~new_n11517 & new_n11536_1;
  assign new_n11569 = ~new_n11537 & ~new_n11568;
  assign new_n11570 = ~new_n11492 & ~new_n11493;
  assign new_n11571 = ~new_n11505 & ~new_n11570;
  assign new_n11572 = new_n11505 & new_n11570;
  assign new_n11573 = ~new_n11571 & ~new_n11572;
  assign new_n11574 = ~new_n11569 & new_n11573;
  assign new_n11575 = new_n11569 & ~new_n11573;
  assign new_n11576 = ~new_n11498 & ~new_n11499;
  assign new_n11577 = ~new_n11503 & new_n11576;
  assign new_n11578 = new_n11503 & ~new_n11576;
  assign new_n11579 = ~new_n11577 & ~new_n11578;
  assign new_n11580 = ~new_n7043 & new_n11519;
  assign new_n11581 = ~new_n11516 & ~new_n11580;
  assign new_n11582 = ~new_n11513 & new_n11580;
  assign new_n11583 = ~new_n11581 & ~new_n11582;
  assign new_n11584 = new_n11579 & ~new_n11583;
  assign new_n11585 = ~new_n11579 & new_n11583;
  assign new_n11586 = ~new_n7060 & ~new_n7088;
  assign new_n11587 = ~new_n7059 & ~new_n11586;
  assign new_n11588 = ~new_n11585 & new_n11587;
  assign new_n11589 = ~new_n11584 & ~new_n11588;
  assign new_n11590 = ~new_n11575 & ~new_n11589;
  assign new_n11591 = ~new_n11574 & ~new_n11590;
  assign new_n11592 = ~new_n11567 & ~new_n11591;
  assign new_n11593 = new_n11567 & new_n11591;
  assign new_n11594 = ~new_n11592 & ~new_n11593;
  assign new_n11595 = new_n11510 & ~new_n11594;
  assign new_n11596 = ~new_n11510 & new_n11594;
  assign n3677 = ~new_n11595 & ~new_n11596;
  assign new_n11598 = ~new_n10018 & ~new_n10019;
  assign new_n11599 = new_n10021 & ~new_n11598;
  assign new_n11600 = ~new_n10021 & new_n11598;
  assign n3849 = ~new_n11599 & ~new_n11600;
  assign new_n11602 = ~new_n7022 & ~new_n7023;
  assign new_n11603 = new_n7037 & new_n11602;
  assign new_n11604 = ~new_n7037 & ~new_n11602;
  assign n4088 = new_n11603 | new_n11604;
  assign new_n11606 = ~new_n1262 & ~new_n1264;
  assign n4155 = ~new_n1265 & ~new_n11606;
  assign new_n11608 = ~new_n3281 & ~new_n3282;
  assign new_n11609 = new_n3326 & ~new_n11608;
  assign new_n11610 = ~new_n3326 & new_n11608;
  assign n4159 = ~new_n11609 & ~new_n11610;
  assign new_n11612 = ~new_n7024 & ~new_n7026;
  assign n4226 = ~new_n7027 & ~new_n11612;
  assign new_n11614 = n7690 & n8665;
  assign new_n11615 = n1067 & n3616;
  assign new_n11616 = new_n11614 & ~new_n11615;
  assign new_n11617 = ~new_n11614 & new_n11615;
  assign new_n11618 = ~new_n11616 & ~new_n11617;
  assign new_n11619 = n2551 & n8476;
  assign new_n11620 = n2530 & n11922;
  assign new_n11621 = new_n11619 & new_n11620;
  assign new_n11622 = ~new_n11619 & ~new_n11620;
  assign new_n11623 = ~new_n11621 & ~new_n11622;
  assign new_n11624 = ~new_n11436 & ~new_n11440;
  assign new_n11625 = ~new_n11439 & ~new_n11624;
  assign new_n11626 = n8665 & n12648;
  assign new_n11627 = n1067 & n10545;
  assign new_n11628 = n5645 & n7690;
  assign new_n11629 = new_n11627 & new_n11628;
  assign new_n11630 = ~new_n11627 & ~new_n11628;
  assign new_n11631 = ~new_n11629 & ~new_n11630;
  assign new_n11632 = ~new_n11626 & ~new_n11631;
  assign new_n11633 = new_n11626 & new_n11631;
  assign new_n11634 = ~new_n11632 & ~new_n11633;
  assign new_n11635 = ~new_n11625 & ~new_n11634;
  assign new_n11636 = new_n11625 & new_n11634;
  assign new_n11637 = ~new_n11635 & ~new_n11636;
  assign new_n11638 = ~new_n11623 & ~new_n11637;
  assign new_n11639 = ~new_n11433 & ~new_n11444;
  assign new_n11640 = ~new_n11434 & ~new_n11639;
  assign new_n11641 = ~new_n11638 & ~new_n11640;
  assign new_n11642 = new_n11621 & new_n11641;
  assign new_n11643 = new_n11623 & new_n11637;
  assign new_n11644 = ~new_n11621 & ~new_n11641;
  assign new_n11645 = ~new_n11643 & new_n11644;
  assign new_n11646 = n8476 & n12826;
  assign new_n11647 = n2530 & n2551;
  assign new_n11648 = n4094 & n5331;
  assign new_n11649 = ~new_n11647 & ~new_n11648;
  assign new_n11650 = new_n11647 & new_n11648;
  assign new_n11651 = ~new_n11649 & ~new_n11650;
  assign new_n11652 = ~new_n11646 & ~new_n11651;
  assign new_n11653 = new_n11646 & new_n11651;
  assign new_n11654 = ~new_n11652 & ~new_n11653;
  assign new_n11655 = new_n11625 & ~new_n11632;
  assign new_n11656 = ~new_n11633 & ~new_n11655;
  assign new_n11657 = new_n11654 & ~new_n11656;
  assign new_n11658 = ~new_n11654 & new_n11656;
  assign new_n11659 = ~new_n11657 & ~new_n11658;
  assign new_n11660 = n1067 & n7690;
  assign new_n11661 = n3616 & n5645;
  assign new_n11662_1 = n8665 & n10545;
  assign new_n11663 = ~new_n11661 & ~new_n11662_1;
  assign new_n11664 = new_n11661 & new_n11662_1;
  assign new_n11665 = ~new_n11663 & ~new_n11664;
  assign new_n11666 = ~new_n11660 & ~new_n11665;
  assign new_n11667 = new_n11660 & new_n11665;
  assign new_n11668 = ~new_n11666 & ~new_n11667;
  assign new_n11669 = n11922 & n12648;
  assign new_n11670 = new_n11629 & new_n11669;
  assign new_n11671 = ~new_n11629 & ~new_n11669;
  assign new_n11672 = ~new_n11670 & ~new_n11671;
  assign new_n11673 = new_n11668 & ~new_n11672;
  assign new_n11674 = ~new_n11668 & new_n11672;
  assign new_n11675 = ~new_n11673 & ~new_n11674;
  assign new_n11676 = ~new_n11659 & ~new_n11675;
  assign new_n11677 = new_n11659 & new_n11675;
  assign new_n11678 = ~new_n11676 & ~new_n11677;
  assign new_n11679 = ~new_n11645 & ~new_n11678;
  assign new_n11680 = ~new_n11642 & ~new_n11679;
  assign new_n11681 = n5964 & n11662;
  assign new_n11682 = n1097 & n7456;
  assign new_n11683 = new_n11681 & new_n11682;
  assign new_n11684 = ~new_n11681 & ~new_n11682;
  assign new_n11685 = ~new_n11683 & ~new_n11684;
  assign new_n11686 = n3932 & n12705;
  assign new_n11687 = n1798 & n12025;
  assign new_n11688 = ~new_n11686 & ~new_n11687;
  assign new_n11689 = new_n11686 & new_n11687;
  assign new_n11690 = ~new_n11688 & ~new_n11689;
  assign new_n11691 = n4312 & n12591;
  assign new_n11692 = ~new_n11540 & ~new_n11544;
  assign new_n11693 = ~new_n11542 & ~new_n11692;
  assign new_n11694 = new_n11691 & new_n11693;
  assign new_n11695 = ~new_n11691 & ~new_n11693;
  assign new_n11696 = ~new_n11694 & ~new_n11695;
  assign new_n11697 = ~new_n11690 & new_n11696;
  assign new_n11698 = new_n11690 & ~new_n11696;
  assign new_n11699 = ~new_n11697 & ~new_n11698;
  assign new_n11700 = ~new_n11685 & new_n11699;
  assign new_n11701 = ~new_n11550 & ~new_n11553;
  assign new_n11702 = ~new_n11549 & ~new_n11701;
  assign new_n11703 = ~new_n11700 & ~new_n11702;
  assign new_n11704 = new_n11683 & new_n11703;
  assign new_n11705 = new_n11685 & ~new_n11699;
  assign new_n11706 = ~new_n11683 & ~new_n11703;
  assign new_n11707_1 = ~new_n11705 & new_n11706;
  assign new_n11708 = n5964 & n10327;
  assign new_n11709 = n1097 & n11662;
  assign new_n11710 = n5305 & n9583;
  assign new_n11711 = ~new_n11709 & ~new_n11710;
  assign new_n11712 = new_n11709 & new_n11710;
  assign new_n11713 = ~new_n11711 & ~new_n11712;
  assign new_n11714 = ~new_n11708 & ~new_n11713;
  assign new_n11715 = new_n11708 & new_n11713;
  assign new_n11716 = ~new_n11714 & ~new_n11715;
  assign new_n11717 = new_n11690 & ~new_n11695;
  assign new_n11718 = ~new_n11694 & ~new_n11717;
  assign new_n11719 = new_n11716 & ~new_n11718;
  assign new_n11720 = ~new_n11716 & new_n11718;
  assign new_n11721 = ~new_n11719 & ~new_n11720;
  assign new_n11722 = n4312 & n7456;
  assign new_n11723 = new_n11689 & new_n11722;
  assign new_n11724 = ~new_n11689 & ~new_n11722;
  assign new_n11725 = ~new_n11723 & ~new_n11724;
  assign new_n11726 = n3932 & n12025;
  assign new_n11727 = n1798 & n11257;
  assign new_n11728_1 = ~new_n11543 & ~new_n11727;
  assign new_n11729 = new_n11543 & new_n11727;
  assign new_n11730 = ~new_n11728_1 & ~new_n11729;
  assign new_n11731 = ~new_n11726 & ~new_n11730;
  assign new_n11732 = new_n11726 & new_n11730;
  assign new_n11733 = ~new_n11731 & ~new_n11732;
  assign new_n11734 = new_n11725 & ~new_n11733;
  assign new_n11735 = ~new_n11725 & new_n11733;
  assign new_n11736 = ~new_n11734 & ~new_n11735;
  assign new_n11737 = new_n11721 & new_n11736;
  assign new_n11738 = ~new_n11721 & ~new_n11736;
  assign new_n11739 = ~new_n11737 & ~new_n11738;
  assign new_n11740 = ~new_n11707_1 & ~new_n11739;
  assign new_n11741 = ~new_n11704 & ~new_n11740;
  assign new_n11742 = n753 & n5305;
  assign new_n11743 = n1798 & n10547;
  assign new_n11744 = ~new_n11742 & new_n11743;
  assign new_n11745 = new_n11742 & ~new_n11743;
  assign new_n11746 = ~new_n11744 & ~new_n11745;
  assign new_n11747 = new_n11741 & new_n11746;
  assign new_n11748 = ~new_n11741 & ~new_n11746;
  assign new_n11749 = ~new_n11747 & ~new_n11748;
  assign new_n11750 = n4094 & n8476;
  assign new_n11751 = ~new_n11646 & ~new_n11650;
  assign new_n11752 = ~new_n11649 & ~new_n11751;
  assign new_n11753 = ~new_n11750 & new_n11752;
  assign new_n11754 = new_n11750 & ~new_n11752;
  assign new_n11755_1 = ~new_n11753 & ~new_n11754;
  assign new_n11756 = ~new_n11668 & ~new_n11670;
  assign new_n11757_1 = ~new_n11671 & ~new_n11756;
  assign new_n11758 = n2530 & n12826;
  assign new_n11759 = ~new_n11660 & ~new_n11664;
  assign new_n11760 = ~new_n11663 & ~new_n11759;
  assign new_n11761 = ~new_n11758 & new_n11760;
  assign new_n11762 = new_n11758 & ~new_n11760;
  assign new_n11763 = ~new_n11761 & ~new_n11762;
  assign new_n11764 = new_n11757_1 & ~new_n11763;
  assign new_n11765 = ~new_n11757_1 & new_n11763;
  assign new_n11766 = ~new_n11764 & ~new_n11765;
  assign new_n11767 = ~new_n11657 & new_n11675;
  assign new_n11768 = ~new_n11658 & ~new_n11767;
  assign new_n11769 = ~new_n11766 & ~new_n11768;
  assign new_n11770 = new_n11766 & new_n11768;
  assign new_n11771 = ~new_n11769 & ~new_n11770;
  assign new_n11772 = ~new_n11755_1 & ~new_n11771;
  assign new_n11773 = new_n11755_1 & new_n11771;
  assign new_n11774 = ~new_n11772 & ~new_n11773;
  assign new_n11775 = ~new_n11749 & new_n11774;
  assign new_n11776 = new_n11749 & ~new_n11774;
  assign new_n11777 = ~new_n11775 & ~new_n11776;
  assign new_n11778 = ~new_n11680 & new_n11777;
  assign new_n11779 = new_n11680 & ~new_n11777;
  assign new_n11780_1 = ~new_n11778 & ~new_n11779;
  assign new_n11781 = ~new_n11618 & new_n11780_1;
  assign new_n11782 = new_n11618 & ~new_n11780_1;
  assign new_n11783 = ~new_n11781 & ~new_n11782;
  assign new_n11784 = ~new_n11700 & ~new_n11705;
  assign new_n11785 = new_n11702 & new_n11784;
  assign new_n11786 = ~new_n11702 & ~new_n11784;
  assign new_n11787 = ~new_n11785 & ~new_n11786;
  assign new_n11788 = ~new_n11558 & ~new_n11561;
  assign new_n11789 = ~new_n11557 & ~new_n11788;
  assign new_n11790 = ~new_n11787 & ~new_n11789;
  assign new_n11791_1 = ~new_n11704 & ~new_n11707_1;
  assign new_n11792 = new_n11739 & new_n11791_1;
  assign new_n11793 = ~new_n11739 & ~new_n11791_1;
  assign new_n11794 = ~new_n11792 & ~new_n11793;
  assign new_n11795 = new_n11790 & ~new_n11794;
  assign new_n11796 = n5305 & n10327;
  assign new_n11797 = new_n11787 & new_n11789;
  assign new_n11798 = ~new_n11790 & ~new_n11797;
  assign new_n11799 = new_n11796 & new_n11798;
  assign new_n11800 = ~new_n11796 & ~new_n11798;
  assign new_n11801 = ~new_n11799 & ~new_n11800;
  assign new_n11802 = new_n11565 & new_n11801;
  assign new_n11803 = ~new_n11799 & ~new_n11802;
  assign new_n11804 = ~new_n11790 & new_n11794;
  assign new_n11805 = ~new_n11795 & ~new_n11804;
  assign new_n11806 = ~new_n11803 & new_n11805;
  assign new_n11807 = ~new_n11795 & ~new_n11806;
  assign new_n11808 = n2551 & n12648;
  assign new_n11809 = n10545 & n11922;
  assign new_n11810 = ~new_n11808 & ~new_n11809;
  assign new_n11811 = new_n11808 & new_n11809;
  assign new_n11812 = ~new_n11810 & ~new_n11811;
  assign new_n11813 = new_n11807 & new_n11812;
  assign new_n11814 = ~new_n11807 & ~new_n11812;
  assign new_n11815 = ~new_n11813 & ~new_n11814;
  assign new_n11816 = ~new_n11783 & new_n11815;
  assign new_n11817 = new_n11783 & ~new_n11815;
  assign new_n11818 = ~new_n11816 & ~new_n11817;
  assign new_n11819 = ~new_n11638 & ~new_n11643;
  assign new_n11820 = new_n11640 & ~new_n11819;
  assign new_n11821_1 = ~new_n11640 & new_n11819;
  assign new_n11822 = ~new_n11820 & ~new_n11821_1;
  assign new_n11823 = ~new_n11449 & new_n11452;
  assign new_n11824 = ~new_n11448 & ~new_n11823;
  assign new_n11825 = new_n11822 & ~new_n11824;
  assign new_n11826 = ~new_n11642 & ~new_n11645;
  assign new_n11827 = new_n11678 & ~new_n11826;
  assign new_n11828 = ~new_n11678 & new_n11826;
  assign new_n11829 = ~new_n11827 & ~new_n11828;
  assign new_n11830 = new_n11825 & new_n11829;
  assign new_n11831 = ~new_n11825 & ~new_n11829;
  assign new_n11832 = ~new_n11830 & ~new_n11831;
  assign new_n11833 = n5331 & n12826;
  assign new_n11834 = ~new_n11822 & new_n11824;
  assign new_n11835 = ~new_n11825 & ~new_n11834;
  assign new_n11836 = new_n11833 & new_n11835;
  assign new_n11837 = ~new_n11833 & ~new_n11835;
  assign new_n11838 = ~new_n11836 & ~new_n11837;
  assign new_n11839 = new_n11456 & new_n11838;
  assign new_n11840 = ~new_n11836 & ~new_n11839;
  assign new_n11841 = new_n11832 & ~new_n11840;
  assign new_n11842 = ~new_n11830 & ~new_n11841;
  assign new_n11843 = ~new_n11329 & ~new_n11332;
  assign new_n11844 = ~new_n11328 & ~new_n11843;
  assign new_n11845 = n6776 & n10451;
  assign new_n11846 = n11023 & n12299;
  assign new_n11847 = ~new_n11845 & ~new_n11846;
  assign new_n11848 = new_n11845 & new_n11846;
  assign new_n11849 = ~new_n11847 & ~new_n11848;
  assign new_n11850 = ~new_n11313 & ~new_n11324;
  assign new_n11851 = ~new_n11314 & ~new_n11850;
  assign new_n11852 = new_n11849 & ~new_n11851;
  assign new_n11853 = ~new_n11849 & new_n11851;
  assign new_n11854 = ~new_n11852 & ~new_n11853;
  assign new_n11855 = n3022 & n7436;
  assign new_n11856 = n8276 & n9640;
  assign new_n11857 = n6703 & n9241;
  assign new_n11858 = ~new_n11856 & ~new_n11857;
  assign new_n11859 = new_n11856 & new_n11857;
  assign new_n11860 = ~new_n11858 & ~new_n11859;
  assign new_n11861 = new_n11855 & new_n11860;
  assign new_n11862 = ~new_n11855 & ~new_n11860;
  assign new_n11863 = ~new_n11861 & ~new_n11862;
  assign new_n11864 = ~new_n11316 & ~new_n11320;
  assign new_n11865 = ~new_n11319 & ~new_n11864;
  assign new_n11866 = ~new_n11863 & new_n11865;
  assign new_n11867 = new_n11863 & ~new_n11865;
  assign new_n11868 = ~new_n11866 & ~new_n11867;
  assign new_n11869 = new_n11854 & new_n11868;
  assign new_n11870 = ~new_n11854 & ~new_n11868;
  assign new_n11871 = ~new_n11869 & ~new_n11870;
  assign new_n11872 = ~new_n11844 & ~new_n11871;
  assign new_n11873 = ~new_n11853 & ~new_n11868;
  assign new_n11874 = new_n11848 & new_n11873;
  assign new_n11875 = ~new_n11848 & ~new_n11873;
  assign new_n11876_1 = ~new_n11852 & new_n11875;
  assign new_n11877_1 = ~new_n11874 & ~new_n11876_1;
  assign new_n11878 = n6776 & n10278;
  assign new_n11879 = n10451 & n12299;
  assign new_n11880 = n8759 & n11423;
  assign new_n11881 = ~new_n11879 & ~new_n11880;
  assign new_n11882 = new_n11879 & new_n11880;
  assign new_n11883 = ~new_n11881 & ~new_n11882;
  assign new_n11884 = ~new_n11878 & ~new_n11883;
  assign new_n11885 = new_n11878 & new_n11883;
  assign new_n11886 = ~new_n11884 & ~new_n11885;
  assign new_n11887 = ~new_n11861 & ~new_n11865;
  assign new_n11888 = ~new_n11862 & ~new_n11887;
  assign new_n11889 = new_n11886 & new_n11888;
  assign new_n11890 = ~new_n11886 & ~new_n11888;
  assign new_n11891 = ~new_n11889 & ~new_n11890;
  assign new_n11892_1 = n7436 & n11023;
  assign new_n11893 = ~new_n11859 & ~new_n11892_1;
  assign new_n11894 = new_n11859 & new_n11892_1;
  assign new_n11895 = ~new_n11893 & ~new_n11894;
  assign new_n11896 = n9241 & n9640;
  assign new_n11897 = n6703 & n10510;
  assign new_n11898 = n3022 & n8276;
  assign new_n11899 = ~new_n11897 & ~new_n11898;
  assign new_n11900 = new_n11897 & new_n11898;
  assign new_n11901 = ~new_n11899 & ~new_n11900;
  assign new_n11902 = ~new_n11896 & ~new_n11901;
  assign new_n11903 = new_n11896 & new_n11901;
  assign new_n11904 = ~new_n11902 & ~new_n11903;
  assign new_n11905 = ~new_n11895 & new_n11904;
  assign new_n11906 = ~new_n11894 & ~new_n11904;
  assign new_n11907 = ~new_n11893 & new_n11906;
  assign new_n11908 = ~new_n11905 & ~new_n11907;
  assign new_n11909 = new_n11891 & new_n11908;
  assign new_n11910 = ~new_n11891 & ~new_n11908;
  assign new_n11911 = ~new_n11909 & ~new_n11910;
  assign new_n11912 = ~new_n11877_1 & ~new_n11911;
  assign new_n11913 = new_n11877_1 & new_n11911;
  assign new_n11914 = ~new_n11912 & ~new_n11913;
  assign new_n11915 = new_n11872 & ~new_n11914;
  assign new_n11916 = ~new_n11872 & new_n11914;
  assign new_n11917_1 = ~new_n11915 & ~new_n11916;
  assign new_n11918 = n8759 & n10278;
  assign new_n11919_1 = new_n11844 & new_n11871;
  assign new_n11920 = ~new_n11872 & ~new_n11919_1;
  assign new_n11921 = new_n11918 & new_n11920;
  assign new_n11922_1 = ~new_n11918 & ~new_n11920;
  assign new_n11923 = ~new_n11921 & ~new_n11922_1;
  assign new_n11924 = new_n11336 & new_n11923;
  assign new_n11925 = ~new_n11921 & ~new_n11924;
  assign new_n11926 = new_n11917_1 & ~new_n11925;
  assign new_n11927 = ~new_n11917_1 & new_n11925;
  assign new_n11928 = ~new_n11926 & ~new_n11927;
  assign new_n11929 = n1510 & n7965;
  assign new_n11930 = n159 & n7388;
  assign new_n11931 = n2749 & n11892;
  assign new_n11932 = ~new_n11930 & ~new_n11931;
  assign new_n11933 = new_n11930 & new_n11931;
  assign new_n11934 = ~new_n11932 & ~new_n11933;
  assign new_n11935 = ~new_n11376 & ~new_n11386;
  assign new_n11936 = ~new_n11375 & ~new_n11935;
  assign new_n11937 = new_n11934 & ~new_n11936;
  assign new_n11938 = ~new_n11934 & new_n11936;
  assign new_n11939 = ~new_n11937 & ~new_n11938;
  assign new_n11940 = n2393 & n3754;
  assign new_n11941 = n5860 & n10898;
  assign new_n11942 = n3986 & n11876;
  assign new_n11943 = ~new_n11941 & ~new_n11942;
  assign new_n11944 = new_n11941 & new_n11942;
  assign new_n11945 = ~new_n11943 & ~new_n11944;
  assign new_n11946 = new_n11940 & new_n11945;
  assign new_n11947 = ~new_n11940 & ~new_n11945;
  assign new_n11948 = ~new_n11946 & ~new_n11947;
  assign new_n11949 = new_n11378 & ~new_n11381;
  assign new_n11950 = ~new_n11382 & ~new_n11949;
  assign new_n11951 = ~new_n11948 & ~new_n11950;
  assign new_n11952 = new_n11948 & new_n11950;
  assign new_n11953 = ~new_n11951 & ~new_n11952;
  assign new_n11954 = ~new_n11939 & new_n11953;
  assign new_n11955 = new_n11939 & ~new_n11953;
  assign new_n11956 = ~new_n11954 & ~new_n11955;
  assign new_n11957 = ~new_n11394 & new_n11956;
  assign new_n11958 = new_n11394 & ~new_n11956;
  assign new_n11959 = ~new_n11957 & ~new_n11958;
  assign new_n11960 = new_n11929 & new_n11959;
  assign new_n11961 = ~new_n11929 & ~new_n11959;
  assign new_n11962 = ~new_n11960 & ~new_n11961;
  assign new_n11963 = new_n11397 & new_n11962;
  assign new_n11964 = ~new_n11397 & ~new_n11962;
  assign new_n11965 = ~new_n11963 & ~new_n11964;
  assign new_n11966 = ~new_n11456 & ~new_n11838;
  assign new_n11967_1 = ~new_n11839 & ~new_n11966;
  assign new_n11968 = ~new_n11965 & ~new_n11967_1;
  assign new_n11969 = new_n11965 & new_n11967_1;
  assign new_n11970 = ~new_n11460 & ~new_n11479;
  assign new_n11971 = ~new_n11459 & ~new_n11970;
  assign new_n11972 = ~new_n11969 & new_n11971;
  assign new_n11973 = ~new_n11968 & ~new_n11972;
  assign new_n11974 = ~new_n11832 & new_n11840;
  assign new_n11975 = ~new_n11841 & ~new_n11974;
  assign new_n11976 = ~new_n11960 & ~new_n11963;
  assign new_n11977 = ~new_n11938 & ~new_n11953;
  assign new_n11978 = new_n11933 & new_n11977;
  assign new_n11979 = ~new_n11933 & ~new_n11977;
  assign new_n11980 = ~new_n11937 & new_n11979;
  assign new_n11981 = ~new_n11978 & ~new_n11980;
  assign new_n11982 = n159 & n11892;
  assign new_n11983 = n7965 & n12247;
  assign new_n11984 = n1510 & n7388;
  assign new_n11985 = ~new_n11983 & ~new_n11984;
  assign new_n11986 = new_n11983 & new_n11984;
  assign new_n11987 = ~new_n11985 & ~new_n11986;
  assign new_n11988 = new_n11982 & ~new_n11987;
  assign new_n11989 = ~new_n11982 & new_n11987;
  assign new_n11990 = ~new_n11988 & ~new_n11989;
  assign new_n11991 = ~new_n11946 & new_n11950;
  assign new_n11992 = ~new_n11947 & ~new_n11991;
  assign new_n11993 = ~new_n11990 & new_n11992;
  assign new_n11994 = new_n11990 & ~new_n11992;
  assign new_n11995 = ~new_n11993 & ~new_n11994;
  assign new_n11996 = n2393 & n2749;
  assign new_n11997 = ~new_n11944 & ~new_n11996;
  assign new_n11998 = new_n11944 & new_n11996;
  assign new_n11999_1 = ~new_n11997 & ~new_n11998;
  assign new_n12000_1 = n3986 & n10898;
  assign new_n12001 = n5857 & n11876;
  assign new_n12002 = n3754 & n5860;
  assign new_n12003 = ~new_n12001 & ~new_n12002;
  assign new_n12004 = new_n12001 & new_n12002;
  assign new_n12005_1 = ~new_n12003 & ~new_n12004;
  assign new_n12006 = ~new_n12000_1 & ~new_n12005_1;
  assign new_n12007 = new_n12000_1 & new_n12005_1;
  assign new_n12008 = ~new_n12006 & ~new_n12007;
  assign new_n12009 = new_n11999_1 & ~new_n12008;
  assign new_n12010 = ~new_n11999_1 & new_n12008;
  assign new_n12011 = ~new_n12009 & ~new_n12010;
  assign new_n12012 = new_n11995 & new_n12011;
  assign new_n12013 = ~new_n11995 & ~new_n12011;
  assign new_n12014_1 = ~new_n12012 & ~new_n12013;
  assign new_n12015 = new_n11981 & new_n12014_1;
  assign new_n12016 = ~new_n11981 & ~new_n12014_1;
  assign new_n12017 = ~new_n12015 & ~new_n12016;
  assign new_n12018 = new_n11957 & ~new_n12017;
  assign new_n12019 = ~new_n11957 & new_n12017;
  assign new_n12020_1 = ~new_n12018 & ~new_n12019;
  assign new_n12021 = ~new_n11976 & new_n12020_1;
  assign new_n12022 = new_n11976 & ~new_n12020_1;
  assign new_n12023 = ~new_n12021 & ~new_n12022;
  assign new_n12024 = new_n11975 & new_n12023;
  assign new_n12025_1 = ~new_n11975 & ~new_n12023;
  assign new_n12026 = ~new_n12024 & ~new_n12025_1;
  assign new_n12027 = ~new_n11973 & ~new_n12026;
  assign new_n12028 = new_n11973 & new_n12026;
  assign new_n12029 = ~new_n12027 & ~new_n12028;
  assign new_n12030 = ~new_n11928 & ~new_n12029;
  assign new_n12031 = new_n11928 & new_n12029;
  assign new_n12032 = ~new_n11336 & ~new_n11923;
  assign new_n12033 = ~new_n11924 & ~new_n12032;
  assign new_n12034 = ~new_n11968 & ~new_n11969;
  assign new_n12035 = new_n11971 & new_n12034;
  assign new_n12036 = ~new_n11971 & ~new_n12034;
  assign new_n12037 = ~new_n12035 & ~new_n12036;
  assign new_n12038 = ~new_n12033 & new_n12037;
  assign new_n12039 = new_n12033 & ~new_n12037;
  assign new_n12040 = ~new_n11484 & ~new_n11507;
  assign new_n12041 = ~new_n11483 & ~new_n12040;
  assign new_n12042 = ~new_n12039 & new_n12041;
  assign new_n12043 = ~new_n12038 & ~new_n12042;
  assign new_n12044_1 = ~new_n12031 & ~new_n12043;
  assign new_n12045 = ~new_n12030 & ~new_n12044_1;
  assign new_n12046 = ~new_n11842 & new_n12045;
  assign new_n12047 = new_n11842 & ~new_n12045;
  assign new_n12048 = ~new_n12046 & ~new_n12047;
  assign new_n12049 = ~new_n11818 & new_n12048;
  assign new_n12050 = new_n11818 & ~new_n12048;
  assign new_n12051 = ~new_n12049 & ~new_n12050;
  assign new_n12052 = ~new_n11915 & ~new_n11926;
  assign new_n12053 = ~new_n11708 & ~new_n11712;
  assign new_n12054 = ~new_n11711 & ~new_n12053;
  assign new_n12055 = n1097 & n10327;
  assign new_n12056 = ~new_n11726 & ~new_n11729;
  assign new_n12057 = ~new_n11728_1 & ~new_n12056;
  assign new_n12058 = ~new_n12055 & new_n12057;
  assign new_n12059 = new_n12055 & ~new_n12057;
  assign new_n12060 = ~new_n12058 & ~new_n12059;
  assign new_n12061 = ~new_n12054 & new_n12060;
  assign new_n12062 = new_n12054 & ~new_n12060;
  assign new_n12063 = ~new_n12061 & ~new_n12062;
  assign new_n12064 = ~new_n11876_1 & ~new_n11911;
  assign new_n12065 = ~new_n11874 & ~new_n12064;
  assign new_n12066 = n9640 & n10510;
  assign new_n12067 = n6703 & n10644;
  assign new_n12068 = n2278 & n8759;
  assign new_n12069_1 = new_n12067 & ~new_n12068;
  assign new_n12070 = ~new_n12067 & new_n12068;
  assign new_n12071 = ~new_n12069_1 & ~new_n12070;
  assign new_n12072 = new_n12066 & ~new_n12071;
  assign new_n12073 = ~new_n12066 & new_n12071;
  assign new_n12074 = ~new_n12072 & ~new_n12073;
  assign new_n12075 = ~new_n12065 & ~new_n12074;
  assign new_n12076_1 = new_n12065 & new_n12074;
  assign new_n12077 = ~new_n12075 & ~new_n12076_1;
  assign new_n12078 = ~new_n11723 & ~new_n11733;
  assign new_n12079 = ~new_n11724 & ~new_n12078;
  assign new_n12080 = n12025 & n12591;
  assign new_n12081 = n3932 & n11257;
  assign new_n12082 = ~new_n12080 & new_n12081;
  assign new_n12083 = new_n12080 & ~new_n12081;
  assign new_n12084 = ~new_n12082 & ~new_n12083;
  assign new_n12085 = n5964 & n9583;
  assign new_n12086 = n4312 & n11662;
  assign new_n12087 = n7456 & n12705;
  assign new_n12088 = new_n12086 & new_n12087;
  assign new_n12089 = ~new_n12086 & ~new_n12087;
  assign new_n12090 = ~new_n12088 & ~new_n12089;
  assign new_n12091 = new_n12085 & ~new_n12090;
  assign new_n12092 = ~new_n12085 & new_n12090;
  assign new_n12093 = ~new_n12091 & ~new_n12092;
  assign new_n12094 = ~new_n12084 & ~new_n12093;
  assign new_n12095 = new_n12084 & new_n12093;
  assign new_n12096 = ~new_n12094 & ~new_n12095;
  assign new_n12097 = ~new_n12079 & new_n12096;
  assign new_n12098 = new_n12079 & ~new_n12096;
  assign new_n12099 = ~new_n12097 & ~new_n12098;
  assign new_n12100 = new_n12077 & new_n12099;
  assign new_n12101 = ~new_n12077 & ~new_n12099;
  assign new_n12102 = ~new_n12100 & ~new_n12101;
  assign new_n12103 = ~new_n12063 & new_n12102;
  assign new_n12104 = new_n12063 & ~new_n12102;
  assign new_n12105 = ~new_n12103 & ~new_n12104;
  assign new_n12106 = new_n12052 & new_n12105;
  assign new_n12107 = ~new_n12052 & ~new_n12105;
  assign new_n12108 = ~new_n12106 & ~new_n12107;
  assign new_n12109 = new_n11973 & ~new_n12025_1;
  assign new_n12110 = ~new_n12024 & ~new_n12109;
  assign new_n12111_1 = ~new_n12108 & new_n12110;
  assign new_n12112 = new_n12108 & ~new_n12110;
  assign new_n12113 = ~new_n12111_1 & ~new_n12112;
  assign new_n12114 = ~new_n12000_1 & ~new_n12004;
  assign new_n12115 = ~new_n12003 & ~new_n12114;
  assign new_n12116 = n2749 & n5860;
  assign new_n12117 = n7388 & n12247;
  assign new_n12118 = n159 & n2393;
  assign new_n12119 = ~new_n12117 & new_n12118;
  assign new_n12120 = new_n12117 & ~new_n12118;
  assign new_n12121 = ~new_n12119 & ~new_n12120;
  assign new_n12122 = ~new_n12116 & new_n12121;
  assign new_n12123 = new_n12116 & ~new_n12121;
  assign new_n12124 = ~new_n12122 & ~new_n12123;
  assign new_n12125 = new_n12115 & ~new_n12124;
  assign new_n12126 = ~new_n12115 & new_n12124;
  assign new_n12127 = ~new_n12125 & ~new_n12126;
  assign new_n12128 = ~new_n11994 & ~new_n12011;
  assign new_n12129 = ~new_n11993 & ~new_n12128;
  assign new_n12130 = new_n12127 & new_n12129;
  assign new_n12131 = ~new_n12127 & ~new_n12129;
  assign new_n12132 = ~new_n12130 & ~new_n12131;
  assign new_n12133 = ~new_n11998 & ~new_n12008;
  assign new_n12134 = ~new_n11997 & ~new_n12133;
  assign new_n12135 = n5331 & n10685;
  assign new_n12136 = n4499 & n5645;
  assign new_n12137 = new_n12135 & ~new_n12136;
  assign new_n12138 = ~new_n12135 & new_n12136;
  assign new_n12139 = ~new_n12137 & ~new_n12138;
  assign new_n12140 = n1510 & n11892;
  assign new_n12141 = ~new_n11982 & ~new_n11986;
  assign new_n12142 = ~new_n11985 & ~new_n12141;
  assign new_n12143 = new_n12140 & new_n12142;
  assign new_n12144 = ~new_n12140 & ~new_n12142;
  assign new_n12145_1 = ~new_n12143 & ~new_n12144;
  assign new_n12146 = new_n12139 & ~new_n12145_1;
  assign new_n12147 = ~new_n12139 & new_n12145_1;
  assign new_n12148 = ~new_n12146 & ~new_n12147;
  assign new_n12149 = ~new_n12134 & new_n12148;
  assign new_n12150 = new_n12134 & ~new_n12148;
  assign new_n12151 = ~new_n12149 & ~new_n12150;
  assign new_n12152 = new_n12132 & ~new_n12151;
  assign new_n12153 = ~new_n12132 & new_n12151;
  assign new_n12154 = ~new_n12152 & ~new_n12153;
  assign new_n12155 = ~new_n12018 & ~new_n12021;
  assign new_n12156 = ~new_n11878 & ~new_n11882;
  assign new_n12157 = ~new_n11881 & ~new_n12156;
  assign new_n12158 = n3754 & n3986;
  assign new_n12159 = n5857 & n10898;
  assign new_n12160 = ~new_n12158 & ~new_n12159;
  assign new_n12161 = new_n12158 & new_n12159;
  assign new_n12162 = ~new_n12160 & ~new_n12161;
  assign new_n12163 = n7965 & n12511;
  assign new_n12164 = n45 & n11876;
  assign new_n12165 = new_n12163 & ~new_n12164;
  assign new_n12166 = ~new_n12163 & new_n12164;
  assign new_n12167 = ~new_n12165 & ~new_n12166;
  assign new_n12168 = ~new_n12162 & ~new_n12167;
  assign new_n12169 = new_n12162 & new_n12167;
  assign new_n12170 = ~new_n12168 & ~new_n12169;
  assign new_n12171 = ~new_n12157 & new_n12170;
  assign new_n12172 = new_n12157 & ~new_n12170;
  assign new_n12173 = ~new_n12171 & ~new_n12172;
  assign new_n12174 = ~new_n11980 & ~new_n12014_1;
  assign new_n12175 = ~new_n11978 & ~new_n12174;
  assign new_n12176 = n10278 & n12299;
  assign new_n12177 = n8276 & n11023;
  assign new_n12178 = n3022 & n9241;
  assign new_n12179 = ~new_n12177 & new_n12178;
  assign new_n12180 = new_n12177 & ~new_n12178;
  assign new_n12181 = ~new_n12179 & ~new_n12180;
  assign new_n12182 = new_n12176 & new_n12181;
  assign new_n12183 = ~new_n12176 & ~new_n12181;
  assign new_n12184 = ~new_n12182 & ~new_n12183;
  assign new_n12185 = ~new_n11893 & ~new_n11906;
  assign new_n12186 = n6776 & n11423;
  assign new_n12187 = new_n12185 & new_n12186;
  assign new_n12188 = ~new_n12185 & ~new_n12186;
  assign new_n12189 = ~new_n12187 & ~new_n12188;
  assign new_n12190 = new_n12184 & ~new_n12189;
  assign new_n12191 = ~new_n12184 & new_n12189;
  assign new_n12192 = ~new_n12190 & ~new_n12191;
  assign new_n12193 = n7436 & n10451;
  assign new_n12194 = ~new_n11896 & ~new_n11900;
  assign new_n12195 = ~new_n11899 & ~new_n12194;
  assign new_n12196 = ~new_n12193 & new_n12195;
  assign new_n12197 = new_n12193 & ~new_n12195;
  assign new_n12198 = ~new_n12196 & ~new_n12197;
  assign new_n12199 = ~new_n11890 & ~new_n11908;
  assign new_n12200 = ~new_n11889 & ~new_n12199;
  assign new_n12201 = new_n12198 & ~new_n12200;
  assign new_n12202 = ~new_n12198 & new_n12200;
  assign new_n12203 = ~new_n12201 & ~new_n12202;
  assign new_n12204 = ~new_n12192 & ~new_n12203;
  assign new_n12205 = new_n12192 & new_n12203;
  assign new_n12206 = ~new_n12204 & ~new_n12205;
  assign new_n12207 = new_n12175 & ~new_n12206;
  assign new_n12208 = ~new_n12175 & new_n12206;
  assign new_n12209 = ~new_n12207 & ~new_n12208;
  assign new_n12210 = ~new_n12173 & new_n12209;
  assign new_n12211 = new_n12173 & ~new_n12209;
  assign new_n12212 = ~new_n12210 & ~new_n12211;
  assign new_n12213 = new_n12155 & new_n12212;
  assign new_n12214 = ~new_n12155 & ~new_n12212;
  assign new_n12215 = ~new_n12213 & ~new_n12214;
  assign new_n12216 = ~new_n11720 & ~new_n11736;
  assign new_n12217 = ~new_n11719 & ~new_n12216;
  assign new_n12218 = ~new_n12215 & new_n12217;
  assign new_n12219 = new_n12215 & ~new_n12217;
  assign new_n12220 = ~new_n12218 & ~new_n12219;
  assign new_n12221_1 = ~new_n12154 & new_n12220;
  assign new_n12222 = new_n12154 & ~new_n12220;
  assign new_n12223 = ~new_n12221_1 & ~new_n12222;
  assign new_n12224 = new_n12113 & ~new_n12223;
  assign new_n12225 = ~new_n12113 & new_n12223;
  assign new_n12226 = ~new_n12224 & ~new_n12225;
  assign new_n12227 = new_n11803 & ~new_n11805;
  assign new_n12228 = ~new_n11806 & ~new_n12227;
  assign new_n12229 = ~new_n12030 & ~new_n12031;
  assign new_n12230 = new_n12043 & ~new_n12229;
  assign new_n12231 = ~new_n12043 & new_n12229;
  assign new_n12232 = ~new_n12230 & ~new_n12231;
  assign new_n12233 = new_n12228 & ~new_n12232;
  assign new_n12234 = ~new_n12228 & new_n12232;
  assign new_n12235 = ~new_n11565 & ~new_n11801;
  assign new_n12236 = ~new_n11802 & ~new_n12235;
  assign new_n12237 = ~new_n12038 & ~new_n12039;
  assign new_n12238 = new_n12041 & ~new_n12237;
  assign new_n12239 = ~new_n12041 & new_n12237;
  assign new_n12240 = ~new_n12238 & ~new_n12239;
  assign new_n12241 = new_n12236 & new_n12240;
  assign new_n12242 = ~new_n12236 & ~new_n12240;
  assign new_n12243 = ~new_n11510 & ~new_n11592;
  assign new_n12244 = ~new_n11593 & ~new_n12243;
  assign new_n12245 = ~new_n12242 & ~new_n12244;
  assign new_n12246 = ~new_n12241 & ~new_n12245;
  assign new_n12247_1 = ~new_n12234 & ~new_n12246;
  assign new_n12248 = ~new_n12233 & ~new_n12247_1;
  assign new_n12249 = new_n12226 & new_n12248;
  assign new_n12250 = ~new_n12226 & ~new_n12248;
  assign new_n12251 = ~new_n12249 & ~new_n12250;
  assign new_n12252 = new_n12051 & new_n12251;
  assign new_n12253 = ~new_n12051 & ~new_n12251;
  assign n4230 = new_n12252 | new_n12253;
  assign new_n12255 = ~new_n6653 & ~new_n6654;
  assign new_n12256 = new_n6674 & ~new_n12255;
  assign new_n12257 = ~new_n6674 & new_n12255;
  assign n4300 = ~new_n12256 & ~new_n12257;
  assign new_n12259 = ~new_n4013 & ~new_n4014;
  assign new_n12260 = new_n4018 & ~new_n12259;
  assign new_n12261 = ~new_n4018 & new_n12259;
  assign n4326 = new_n12260 | new_n12261;
  assign new_n12263 = n5320 & n6687;
  assign new_n12264 = ~new_n1394 & ~new_n1404;
  assign new_n12265 = ~new_n1393 & ~new_n12264;
  assign new_n12266 = new_n12263 & ~new_n12265;
  assign new_n12267 = ~new_n12263 & new_n12265;
  assign new_n12268 = ~new_n12266 & ~new_n12267;
  assign new_n12269 = n2564 & n4370;
  assign new_n12270 = new_n1396 & ~new_n1399;
  assign new_n12271 = ~new_n1400 & ~new_n12270;
  assign new_n12272 = new_n12269 & ~new_n12271;
  assign new_n12273 = ~new_n12269 & new_n12271;
  assign new_n12274 = ~new_n12272 & ~new_n12273;
  assign new_n12275 = n5212 & n6770;
  assign new_n12276 = n9920 & n11407;
  assign new_n12277 = ~new_n1382 & ~new_n12276;
  assign new_n12278 = new_n1382 & new_n12276;
  assign new_n12279 = ~new_n12277 & ~new_n12278;
  assign new_n12280 = new_n12275 & ~new_n12279;
  assign new_n12281 = ~new_n12275 & new_n12279;
  assign new_n12282 = ~new_n12280 & ~new_n12281;
  assign new_n12283 = ~new_n12274 & ~new_n12282;
  assign new_n12284 = new_n12274 & new_n12282;
  assign new_n12285 = ~new_n12283 & ~new_n12284;
  assign new_n12286 = ~new_n12268 & ~new_n12285;
  assign new_n12287 = new_n12268 & new_n12285;
  assign new_n12288 = ~new_n12286 & ~new_n12287;
  assign new_n12289 = new_n1408 & ~new_n12288;
  assign new_n12290 = ~new_n1408 & new_n12288;
  assign new_n12291 = ~new_n12289 & ~new_n12290;
  assign new_n12292 = n2433 & n8336;
  assign new_n12293 = n8819 & n10928;
  assign new_n12294 = new_n1516 & ~new_n1519;
  assign new_n12295 = ~new_n1520 & ~new_n12294;
  assign new_n12296 = ~new_n12293 & new_n12295;
  assign new_n12297 = new_n12293 & ~new_n12295;
  assign new_n12298 = ~new_n12296 & ~new_n12297;
  assign new_n12299_1 = n1094 & n12709;
  assign new_n12300 = n6429 & n6986;
  assign new_n12301 = n2226 & n11728;
  assign new_n12302 = ~new_n12300 & ~new_n12301;
  assign new_n12303 = new_n12300 & new_n12301;
  assign new_n12304 = ~new_n12302 & ~new_n12303;
  assign new_n12305 = new_n12299_1 & ~new_n12304;
  assign new_n12306 = ~new_n12299_1 & new_n12304;
  assign new_n12307 = ~new_n12305 & ~new_n12306;
  assign new_n12308 = ~new_n12298 & new_n12307;
  assign new_n12309 = new_n12298 & ~new_n12307;
  assign new_n12310 = ~new_n12308 & ~new_n12309;
  assign new_n12311 = new_n12292 & new_n12310;
  assign new_n12312 = ~new_n12292 & ~new_n12310;
  assign new_n12313 = ~new_n12311 & ~new_n12312;
  assign new_n12314 = ~new_n1525 & new_n1529;
  assign new_n12315 = ~new_n1526 & ~new_n12314;
  assign new_n12316 = ~new_n12313 & new_n12315;
  assign new_n12317 = new_n12313 & ~new_n12315;
  assign new_n12318 = ~new_n12316 & ~new_n12317;
  assign new_n12319 = new_n1534 & ~new_n12318;
  assign new_n12320 = ~new_n1534 & new_n12318;
  assign new_n12321 = ~new_n12319 & ~new_n12320;
  assign new_n12322 = ~new_n1588 & ~new_n1591;
  assign new_n12323 = ~new_n1587 & ~new_n12322;
  assign new_n12324 = new_n12321 & ~new_n12323;
  assign new_n12325 = ~new_n12321 & new_n12323;
  assign new_n12326 = ~new_n12324 & ~new_n12325;
  assign new_n12327 = n11967 & n12069;
  assign new_n12328 = n6254 & n12391;
  assign new_n12329 = new_n1543 & ~new_n1546;
  assign new_n12330 = ~new_n1547 & ~new_n12329;
  assign new_n12331 = ~new_n12328 & new_n12330;
  assign new_n12332 = new_n12328 & ~new_n12330;
  assign new_n12333 = ~new_n12331 & ~new_n12332;
  assign new_n12334 = n4828 & n12489;
  assign new_n12335 = n7159 & n7160;
  assign new_n12336 = ~new_n1429 & ~new_n12335;
  assign new_n12337 = new_n1429 & new_n12335;
  assign new_n12338 = ~new_n12336 & ~new_n12337;
  assign new_n12339 = new_n12334 & ~new_n12338;
  assign new_n12340 = ~new_n12334 & new_n12338;
  assign new_n12341 = ~new_n12339 & ~new_n12340;
  assign new_n12342 = ~new_n12333 & new_n12341;
  assign new_n12343 = new_n12333 & ~new_n12341;
  assign new_n12344 = ~new_n12342 & ~new_n12343;
  assign new_n12345 = new_n12327 & new_n12344;
  assign new_n12346 = ~new_n12327 & ~new_n12344;
  assign new_n12347 = ~new_n12345 & ~new_n12346;
  assign new_n12348 = ~new_n1541 & ~new_n1551;
  assign new_n12349 = ~new_n1540 & ~new_n12348;
  assign new_n12350 = ~new_n12347 & ~new_n12349;
  assign new_n12351 = new_n12347 & new_n12349;
  assign new_n12352 = ~new_n12350 & ~new_n12351;
  assign new_n12353 = new_n1556 & ~new_n12352;
  assign new_n12354 = ~new_n1556 & new_n12352;
  assign new_n12355 = ~new_n12353 & ~new_n12354;
  assign new_n12356 = n11222 & n12947;
  assign new_n12357 = n11153 & n11791;
  assign new_n12358 = new_n1564_1 & ~new_n1567;
  assign new_n12359 = ~new_n1568 & ~new_n12358;
  assign new_n12360 = ~new_n12357 & new_n12359;
  assign new_n12361 = new_n12357 & ~new_n12359;
  assign new_n12362 = ~new_n12360 & ~new_n12361;
  assign new_n12363 = n5767 & n10990;
  assign new_n12364 = n1478 & n5314;
  assign new_n12365 = n996 & n5760;
  assign new_n12366 = ~new_n12364 & ~new_n12365;
  assign new_n12367 = new_n12364 & new_n12365;
  assign new_n12368 = ~new_n12366 & ~new_n12367;
  assign new_n12369 = new_n12363 & ~new_n12368;
  assign new_n12370 = ~new_n12363 & new_n12368;
  assign new_n12371 = ~new_n12369 & ~new_n12370;
  assign new_n12372 = ~new_n12362 & new_n12371;
  assign new_n12373 = new_n12362 & ~new_n12371;
  assign new_n12374 = ~new_n12372 & ~new_n12373;
  assign new_n12375 = new_n12356 & new_n12374;
  assign new_n12376 = ~new_n12356 & ~new_n12374;
  assign new_n12377 = ~new_n12375 & ~new_n12376;
  assign new_n12378 = ~new_n1562 & ~new_n1572;
  assign new_n12379 = ~new_n1561 & ~new_n12378;
  assign new_n12380 = ~new_n12377 & ~new_n12379;
  assign new_n12381 = new_n12377 & new_n12379;
  assign new_n12382 = ~new_n12380 & ~new_n12381;
  assign new_n12383 = ~new_n1576_1 & new_n12382;
  assign new_n12384 = new_n1576_1 & ~new_n12382;
  assign new_n12385 = ~new_n12383 & ~new_n12384;
  assign new_n12386 = ~new_n1580 & ~new_n1583;
  assign new_n12387 = ~new_n1579 & ~new_n12386;
  assign new_n12388 = new_n12385 & ~new_n12387;
  assign new_n12389 = ~new_n12385 & new_n12387;
  assign new_n12390 = ~new_n12388 & ~new_n12389;
  assign new_n12391_1 = new_n12355 & new_n12390;
  assign new_n12392 = ~new_n12355 & ~new_n12390;
  assign new_n12393 = ~new_n12391_1 & ~new_n12392;
  assign new_n12394 = ~new_n12326 & new_n12393;
  assign new_n12395 = new_n12326 & ~new_n12393;
  assign new_n12396 = ~new_n12394 & ~new_n12395;
  assign new_n12397 = ~new_n12291 & new_n12396;
  assign new_n12398 = new_n12291 & ~new_n12396;
  assign new_n12399 = ~new_n12397 & ~new_n12398;
  assign new_n12400 = ~new_n1513 & ~new_n1594;
  assign new_n12401 = ~new_n1512_1 & ~new_n12400;
  assign new_n12402 = ~new_n12399 & new_n12401;
  assign new_n12403 = new_n12399 & ~new_n12401;
  assign n4333 = ~new_n12402 & ~new_n12403;
  assign new_n12405 = n7862 & n12000;
  assign new_n12406 = n1333 & n5320;
  assign new_n12407 = n3172 & n4370;
  assign new_n12408 = ~new_n12406 & ~new_n12407;
  assign new_n12409 = new_n12406 & new_n12407;
  assign new_n12410 = ~new_n12408 & ~new_n12409;
  assign new_n12411 = n5240 & n11877;
  assign new_n12412 = n3172 & n11407;
  assign new_n12413 = new_n12411 & new_n12412;
  assign new_n12414 = n5212 & n11757;
  assign new_n12415 = n5240 & n11407;
  assign new_n12416 = n3172 & n11877;
  assign new_n12417 = ~new_n12415 & ~new_n12416;
  assign new_n12418 = new_n12414 & ~new_n12417;
  assign new_n12419 = ~new_n12413 & ~new_n12418;
  assign new_n12420 = n11757 & n11877;
  assign new_n12421 = n5212 & n5240;
  assign new_n12422 = n11407 & n11821;
  assign new_n12423 = ~new_n12421 & ~new_n12422;
  assign new_n12424 = new_n12421 & new_n12422;
  assign new_n12425 = ~new_n12423 & ~new_n12424;
  assign new_n12426 = new_n12420 & new_n12425;
  assign new_n12427 = ~new_n12420 & ~new_n12425;
  assign new_n12428 = ~new_n12426 & ~new_n12427;
  assign new_n12429 = new_n12419 & ~new_n12428;
  assign new_n12430 = ~new_n12419 & new_n12428;
  assign new_n12431 = ~new_n12429 & ~new_n12430;
  assign new_n12432 = ~new_n12410 & ~new_n12431;
  assign new_n12433 = new_n12410 & new_n12431;
  assign new_n12434 = ~new_n12432 & ~new_n12433;
  assign new_n12435 = n1333 & n4370;
  assign new_n12436 = n1333 & n11407;
  assign new_n12437 = new_n12420 & new_n12436;
  assign new_n12438 = n1333 & n11877;
  assign new_n12439 = n11407 & n11757;
  assign new_n12440 = ~new_n12438 & ~new_n12439;
  assign new_n12441 = n3172 & n5212;
  assign new_n12442 = ~new_n12440 & new_n12441;
  assign new_n12443 = ~new_n12437 & ~new_n12442;
  assign new_n12444_1 = ~new_n12435 & new_n12443;
  assign new_n12445 = new_n12435 & ~new_n12443;
  assign new_n12446 = ~new_n12413 & ~new_n12417;
  assign new_n12447 = ~new_n12414 & ~new_n12446;
  assign new_n12448 = new_n12414 & new_n12446;
  assign new_n12449 = ~new_n12447 & ~new_n12448;
  assign new_n12450 = ~new_n12445 & ~new_n12449;
  assign new_n12451 = ~new_n12444_1 & ~new_n12450;
  assign new_n12452 = ~new_n12434 & ~new_n12451;
  assign new_n12453 = new_n12434 & new_n12451;
  assign new_n12454 = ~new_n12452 & ~new_n12453;
  assign new_n12455 = n5320 & n7862;
  assign new_n12456 = ~new_n12444_1 & ~new_n12445;
  assign new_n12457 = ~new_n12449 & ~new_n12456;
  assign new_n12458 = new_n12449 & new_n12456;
  assign new_n12459 = ~new_n12457 & ~new_n12458;
  assign new_n12460 = new_n12455 & new_n12459;
  assign new_n12461 = ~new_n12455 & ~new_n12459;
  assign new_n12462 = n4370 & n7862;
  assign new_n12463 = n7862 & n11877;
  assign new_n12464 = n1333 & n5212;
  assign new_n12465 = new_n12463 & new_n12464;
  assign new_n12466 = ~new_n12463 & ~new_n12464;
  assign new_n12467 = new_n12412 & ~new_n12466;
  assign new_n12468 = ~new_n12465 & ~new_n12467;
  assign new_n12469 = ~new_n12462 & new_n12468;
  assign new_n12470 = new_n12462 & ~new_n12468;
  assign new_n12471 = ~new_n12437 & ~new_n12440;
  assign new_n12472 = ~new_n12441 & ~new_n12471;
  assign new_n12473 = new_n12441 & new_n12471;
  assign new_n12474 = ~new_n12472 & ~new_n12473;
  assign new_n12475 = ~new_n12470 & ~new_n12474;
  assign new_n12476 = ~new_n12469 & ~new_n12475;
  assign new_n12477 = ~new_n12461 & new_n12476;
  assign new_n12478 = ~new_n12460 & ~new_n12477;
  assign new_n12479 = new_n12454 & ~new_n12478;
  assign new_n12480 = ~new_n12454 & new_n12478;
  assign new_n12481 = ~new_n12479 & ~new_n12480;
  assign new_n12482 = new_n12405 & new_n12481;
  assign new_n12483 = n5212 & n7862;
  assign new_n12484 = new_n12436 & new_n12483;
  assign new_n12485 = ~new_n12465 & ~new_n12466;
  assign new_n12486 = ~new_n12412 & ~new_n12485;
  assign new_n12487 = new_n12412 & new_n12485;
  assign new_n12488 = ~new_n12486 & ~new_n12487;
  assign new_n12489_1 = new_n12484 & new_n12488;
  assign new_n12490 = ~new_n12469 & new_n12475;
  assign new_n12491 = ~new_n12469 & ~new_n12470;
  assign new_n12492 = new_n12474 & ~new_n12491;
  assign new_n12493 = ~new_n12490 & ~new_n12492;
  assign new_n12494 = new_n12489_1 & ~new_n12493;
  assign new_n12495 = ~new_n12460 & ~new_n12461;
  assign new_n12496 = ~new_n12476 & ~new_n12495;
  assign new_n12497 = new_n12476 & new_n12495;
  assign new_n12498 = ~new_n12496 & ~new_n12497;
  assign new_n12499 = new_n12494 & new_n12498;
  assign new_n12500 = ~new_n12405 & ~new_n12481;
  assign new_n12501 = ~new_n12482 & ~new_n12500;
  assign new_n12502 = new_n12499 & new_n12501;
  assign new_n12503 = ~new_n12482 & ~new_n12502;
  assign new_n12504 = ~new_n12432 & new_n12451;
  assign new_n12505 = ~new_n12409 & ~new_n12504;
  assign new_n12506 = ~new_n12433 & new_n12505;
  assign new_n12507 = new_n12409 & new_n12504;
  assign new_n12508 = ~new_n12506 & ~new_n12507;
  assign new_n12509 = n1333 & n12000;
  assign new_n12510 = n7862 & n9725;
  assign new_n12511_1 = n3172 & n5320;
  assign new_n12512 = ~new_n12510 & ~new_n12511_1;
  assign new_n12513 = new_n12510 & new_n12511_1;
  assign new_n12514 = ~new_n12512 & ~new_n12513;
  assign new_n12515 = ~new_n12509 & ~new_n12514;
  assign new_n12516 = new_n12509 & new_n12514;
  assign new_n12517 = ~new_n12515 & ~new_n12516;
  assign new_n12518 = new_n12419 & ~new_n12426;
  assign new_n12519 = ~new_n12427 & ~new_n12518;
  assign new_n12520 = ~new_n12517 & ~new_n12519;
  assign new_n12521 = new_n12517 & new_n12519;
  assign new_n12522 = ~new_n12520 & ~new_n12521;
  assign new_n12523 = n4370 & n11757;
  assign new_n12524 = new_n12424 & new_n12523;
  assign new_n12525 = ~new_n12424 & ~new_n12523;
  assign new_n12526 = ~new_n12524 & ~new_n12525;
  assign new_n12527 = n5212 & n11821;
  assign new_n12528 = n9080 & n11407;
  assign new_n12529 = new_n12411 & new_n12528;
  assign new_n12530 = ~new_n12411 & ~new_n12528;
  assign new_n12531 = ~new_n12529 & ~new_n12530;
  assign new_n12532 = ~new_n12527 & ~new_n12531;
  assign new_n12533 = new_n12527 & new_n12531;
  assign new_n12534 = ~new_n12532 & ~new_n12533;
  assign new_n12535 = new_n12526 & ~new_n12534;
  assign new_n12536 = ~new_n12526 & new_n12534;
  assign new_n12537 = ~new_n12535 & ~new_n12536;
  assign new_n12538 = new_n12522 & ~new_n12537;
  assign new_n12539 = ~new_n12522 & new_n12537;
  assign new_n12540 = ~new_n12538 & ~new_n12539;
  assign new_n12541 = new_n12508 & ~new_n12540;
  assign new_n12542 = ~new_n12508 & new_n12540;
  assign new_n12543 = ~new_n12541 & ~new_n12542;
  assign new_n12544 = new_n12479 & ~new_n12543;
  assign new_n12545 = ~new_n12479 & new_n12543;
  assign new_n12546 = ~new_n12544 & ~new_n12545;
  assign new_n12547 = ~new_n12503 & new_n12546;
  assign new_n12548 = new_n12503 & ~new_n12546;
  assign new_n12549 = ~new_n12547 & ~new_n12548;
  assign new_n12550 = n2464 & n6429;
  assign new_n12551 = n6877 & n12709;
  assign new_n12552 = new_n12550 & new_n12551;
  assign new_n12553 = n2464 & n12709;
  assign new_n12554 = n6429 & n6877;
  assign new_n12555 = ~new_n12553 & ~new_n12554;
  assign new_n12556 = ~new_n12552 & ~new_n12555;
  assign new_n12557 = n9400 & n12709;
  assign new_n12558 = n6877 & n11728;
  assign new_n12559 = new_n12557 & new_n12558;
  assign new_n12560 = ~new_n12556 & new_n12559;
  assign new_n12561 = n2464 & n11728;
  assign new_n12562 = n6429 & n11311;
  assign new_n12563 = new_n12557 & new_n12562;
  assign new_n12564 = n11311 & n12709;
  assign new_n12565 = n6429 & n9400;
  assign new_n12566 = ~new_n12564 & ~new_n12565;
  assign new_n12567 = ~new_n12563 & ~new_n12566;
  assign new_n12568 = ~new_n12561 & ~new_n12567;
  assign new_n12569 = new_n12561 & new_n12567;
  assign new_n12570 = ~new_n12568 & ~new_n12569;
  assign new_n12571 = n6877 & n8819;
  assign new_n12572 = n9400 & n11728;
  assign new_n12573 = ~new_n12555 & new_n12572;
  assign new_n12574 = ~new_n12552 & ~new_n12573;
  assign new_n12575 = ~new_n12571 & new_n12574;
  assign new_n12576 = new_n12571 & ~new_n12574;
  assign new_n12577 = ~new_n12575 & ~new_n12576;
  assign new_n12578 = ~new_n12570 & ~new_n12577;
  assign new_n12579 = new_n12570 & new_n12577;
  assign new_n12580 = ~new_n12578 & ~new_n12579;
  assign new_n12581 = new_n12560 & new_n12580;
  assign new_n12582 = ~new_n12570 & ~new_n12576;
  assign new_n12583 = ~new_n12575 & ~new_n12582;
  assign new_n12584 = n2433 & n6877;
  assign new_n12585 = n11311 & n11728;
  assign new_n12586 = n4187 & n6429;
  assign new_n12587 = new_n12553 & new_n12586;
  assign new_n12588 = n4187 & n12709;
  assign new_n12589 = ~new_n12550 & ~new_n12588;
  assign new_n12590 = ~new_n12587 & ~new_n12589;
  assign new_n12591_1 = ~new_n12585 & ~new_n12590;
  assign new_n12592 = new_n12585 & new_n12590;
  assign new_n12593 = ~new_n12591_1 & ~new_n12592;
  assign new_n12594 = n8819 & n9400;
  assign new_n12595 = new_n12561 & ~new_n12566;
  assign new_n12596 = ~new_n12563 & ~new_n12595;
  assign new_n12597 = ~new_n12594 & new_n12596;
  assign new_n12598 = new_n12594 & ~new_n12596;
  assign new_n12599 = ~new_n12597 & ~new_n12598;
  assign new_n12600 = ~new_n12593 & ~new_n12599;
  assign new_n12601 = new_n12593 & new_n12599;
  assign new_n12602 = ~new_n12600 & ~new_n12601;
  assign new_n12603 = ~new_n12584 & ~new_n12602;
  assign new_n12604 = new_n12584 & new_n12602;
  assign new_n12605 = ~new_n12603 & ~new_n12604;
  assign new_n12606 = new_n12583 & new_n12605;
  assign new_n12607 = ~new_n12583 & ~new_n12605;
  assign new_n12608 = ~new_n12606 & ~new_n12607;
  assign new_n12609 = new_n12581 & new_n12608;
  assign new_n12610 = n6877 & n8717;
  assign new_n12611 = n2433 & n9400;
  assign new_n12612 = n2464 & n8819;
  assign new_n12613 = ~new_n12611 & ~new_n12612;
  assign new_n12614 = new_n12611 & new_n12612;
  assign new_n12615 = ~new_n12613 & ~new_n12614;
  assign new_n12616 = n4203 & n12709;
  assign new_n12617 = n4187 & n11728;
  assign new_n12618 = ~new_n12616 & ~new_n12617;
  assign new_n12619 = new_n12616 & new_n12617;
  assign new_n12620 = ~new_n12618 & ~new_n12619;
  assign new_n12621 = new_n12562 & new_n12620;
  assign new_n12622 = ~new_n12562 & ~new_n12620;
  assign new_n12623 = ~new_n12621 & ~new_n12622;
  assign new_n12624 = new_n12585 & ~new_n12589;
  assign new_n12625 = ~new_n12587 & ~new_n12624;
  assign new_n12626 = new_n12623 & new_n12625;
  assign new_n12627 = ~new_n12623 & ~new_n12625;
  assign new_n12628 = ~new_n12626 & ~new_n12627;
  assign new_n12629 = ~new_n12615 & new_n12628;
  assign new_n12630 = new_n12615 & ~new_n12628;
  assign new_n12631 = ~new_n12629 & ~new_n12630;
  assign new_n12632 = ~new_n12593 & ~new_n12598;
  assign new_n12633 = ~new_n12597 & ~new_n12632;
  assign new_n12634 = ~new_n12631 & ~new_n12633;
  assign new_n12635 = new_n12631 & new_n12633;
  assign new_n12636 = ~new_n12634 & ~new_n12635;
  assign new_n12637 = new_n12583 & ~new_n12603;
  assign new_n12638 = ~new_n12604 & ~new_n12637;
  assign new_n12639 = new_n12636 & ~new_n12638;
  assign new_n12640 = ~new_n12636 & new_n12638;
  assign new_n12641 = ~new_n12639 & ~new_n12640;
  assign new_n12642 = new_n12610 & new_n12641;
  assign new_n12643 = ~new_n12610 & ~new_n12641;
  assign new_n12644 = ~new_n12642 & ~new_n12643;
  assign new_n12645 = new_n12609 & new_n12644;
  assign new_n12646 = ~new_n12609 & ~new_n12644;
  assign new_n12647 = ~new_n12645 & ~new_n12646;
  assign new_n12648_1 = ~new_n12581 & ~new_n12608;
  assign new_n12649 = ~new_n12609 & ~new_n12648_1;
  assign new_n12650 = ~new_n12560 & ~new_n12580;
  assign new_n12651 = ~new_n12581 & ~new_n12650;
  assign new_n12652 = n5283 & n12777;
  assign new_n12653 = n4805 & n12489;
  assign new_n12654 = new_n12652 & new_n12653;
  assign new_n12655 = n5283 & n12489;
  assign new_n12656 = n4805 & n12777;
  assign new_n12657 = ~new_n12655 & ~new_n12656;
  assign new_n12658 = ~new_n12654 & ~new_n12657;
  assign new_n12659 = n11478 & n12489;
  assign new_n12660 = n4805 & n7159;
  assign new_n12661 = new_n12659 & new_n12660;
  assign new_n12662 = ~new_n12658 & new_n12661;
  assign new_n12663 = n5283 & n7159;
  assign new_n12664 = n137 & n12777;
  assign new_n12665 = new_n12659 & new_n12664;
  assign new_n12666 = n137 & n12489;
  assign new_n12667 = n11478 & n12777;
  assign new_n12668 = ~new_n12666 & ~new_n12667;
  assign new_n12669 = ~new_n12665 & ~new_n12668;
  assign new_n12670 = ~new_n12663 & ~new_n12669;
  assign new_n12671 = new_n12663 & new_n12669;
  assign new_n12672 = ~new_n12670 & ~new_n12671;
  assign new_n12673 = n4805 & n6254;
  assign new_n12674 = n7159 & n11478;
  assign new_n12675 = ~new_n12657 & new_n12674;
  assign new_n12676 = ~new_n12654 & ~new_n12675;
  assign new_n12677 = ~new_n12673 & new_n12676;
  assign new_n12678 = new_n12673 & ~new_n12676;
  assign new_n12679 = ~new_n12677 & ~new_n12678;
  assign new_n12680 = ~new_n12672 & ~new_n12679;
  assign new_n12681 = new_n12672 & new_n12679;
  assign new_n12682 = ~new_n12680 & ~new_n12681;
  assign new_n12683 = new_n12662 & new_n12682;
  assign new_n12684 = ~new_n12662 & ~new_n12682;
  assign new_n12685 = ~new_n12683 & ~new_n12684;
  assign new_n12686 = n1478 & n8384;
  assign new_n12687 = n7236 & n10990;
  assign new_n12688 = new_n12686 & new_n12687;
  assign new_n12689 = n8384 & n10990;
  assign new_n12690 = n1478 & n7236;
  assign new_n12691 = ~new_n12689 & ~new_n12690;
  assign new_n12692 = ~new_n12688 & ~new_n12691;
  assign new_n12693 = n3992 & n10990;
  assign new_n12694 = n5760 & n7236;
  assign new_n12695 = new_n12693 & new_n12694;
  assign new_n12696 = ~new_n12692 & new_n12695;
  assign new_n12697 = n5760 & n8384;
  assign new_n12698 = n1478 & n6358;
  assign new_n12699 = new_n12693 & new_n12698;
  assign new_n12700 = n6358 & n10990;
  assign new_n12701 = n1478 & n3992;
  assign new_n12702 = ~new_n12700 & ~new_n12701;
  assign new_n12703 = ~new_n12699 & ~new_n12702;
  assign new_n12704_1 = ~new_n12697 & ~new_n12703;
  assign new_n12705_1 = new_n12697 & new_n12703;
  assign new_n12706_1 = ~new_n12704_1 & ~new_n12705_1;
  assign new_n12707 = n7236 & n11791;
  assign new_n12708 = n3992 & n5760;
  assign new_n12709_1 = ~new_n12691 & new_n12708;
  assign new_n12710 = ~new_n12688 & ~new_n12709_1;
  assign new_n12711 = ~new_n12707 & new_n12710;
  assign new_n12712 = new_n12707 & ~new_n12710;
  assign new_n12713 = ~new_n12711 & ~new_n12712;
  assign new_n12714 = ~new_n12706_1 & ~new_n12713;
  assign new_n12715 = new_n12706_1 & new_n12713;
  assign new_n12716 = ~new_n12714 & ~new_n12715;
  assign new_n12717 = new_n12696 & new_n12716;
  assign new_n12718 = ~new_n12696 & ~new_n12716;
  assign new_n12719 = ~new_n12717 & ~new_n12718;
  assign new_n12720_1 = ~new_n12685 & ~new_n12719;
  assign new_n12721 = new_n12685 & new_n12719;
  assign new_n12722 = ~new_n12720_1 & ~new_n12721;
  assign new_n12723 = new_n12653 & new_n12687;
  assign new_n12724 = ~new_n12659 & ~new_n12660;
  assign new_n12725 = ~new_n12661 & ~new_n12724;
  assign new_n12726 = new_n12723 & new_n12725;
  assign new_n12727 = ~new_n12723 & ~new_n12725;
  assign new_n12728 = ~new_n12693 & ~new_n12694;
  assign new_n12729 = ~new_n12695 & ~new_n12728;
  assign new_n12730 = ~new_n12727 & new_n12729;
  assign new_n12731 = ~new_n12726 & ~new_n12730;
  assign new_n12732 = ~new_n12687 & new_n12708;
  assign new_n12733 = new_n12691 & new_n12732;
  assign new_n12734 = new_n12692 & ~new_n12732;
  assign new_n12735 = ~new_n12733 & ~new_n12734;
  assign new_n12736 = ~new_n12731 & ~new_n12735;
  assign new_n12737 = new_n12731 & new_n12735;
  assign new_n12738 = ~new_n12653 & new_n12674;
  assign new_n12739 = ~new_n12658 & ~new_n12738;
  assign new_n12740 = ~new_n12657 & new_n12738;
  assign new_n12741 = ~new_n12739 & ~new_n12740;
  assign new_n12742 = ~new_n12737 & new_n12741;
  assign new_n12743 = ~new_n12736 & ~new_n12742;
  assign new_n12744 = ~new_n12722 & new_n12743;
  assign new_n12745 = new_n12722 & ~new_n12743;
  assign new_n12746 = ~new_n12744 & ~new_n12745;
  assign new_n12747 = ~new_n12651 & ~new_n12746;
  assign new_n12748 = new_n12651 & new_n12746;
  assign new_n12749 = ~new_n12551 & new_n12572;
  assign new_n12750 = new_n12555 & new_n12749;
  assign new_n12751 = new_n12556 & ~new_n12749;
  assign new_n12752 = ~new_n12750 & ~new_n12751;
  assign new_n12753_1 = ~new_n12736 & ~new_n12737;
  assign new_n12754 = new_n12741 & new_n12753_1;
  assign new_n12755 = ~new_n12741 & ~new_n12753_1;
  assign new_n12756 = ~new_n12754 & ~new_n12755;
  assign new_n12757 = new_n12752 & ~new_n12756;
  assign new_n12758 = ~new_n12752 & new_n12756;
  assign new_n12759 = ~new_n12557 & ~new_n12558;
  assign new_n12760 = ~new_n12559 & ~new_n12759;
  assign new_n12761 = ~new_n12726 & ~new_n12727;
  assign new_n12762 = new_n12729 & ~new_n12761;
  assign new_n12763 = ~new_n12729 & new_n12761;
  assign new_n12764 = ~new_n12762 & ~new_n12763;
  assign new_n12765 = new_n12760 & ~new_n12764;
  assign new_n12766 = ~new_n12760 & new_n12764;
  assign new_n12767 = ~new_n12653 & ~new_n12687;
  assign new_n12768 = ~new_n12723 & ~new_n12767;
  assign new_n12769 = new_n12551 & new_n12768;
  assign new_n12770 = ~new_n12766 & new_n12769;
  assign new_n12771 = ~new_n12765 & ~new_n12770;
  assign new_n12772 = ~new_n12758 & new_n12771;
  assign new_n12773 = ~new_n12757 & ~new_n12772;
  assign new_n12774 = ~new_n12748 & ~new_n12773;
  assign new_n12775 = ~new_n12747 & ~new_n12774;
  assign new_n12776 = new_n12649 & new_n12775;
  assign new_n12777_1 = ~new_n12649 & ~new_n12775;
  assign new_n12778 = n4805 & n11967;
  assign new_n12779 = ~new_n12672 & ~new_n12678;
  assign new_n12780 = ~new_n12677 & ~new_n12779;
  assign new_n12781 = ~new_n12778 & ~new_n12780;
  assign new_n12782 = new_n12778 & new_n12780;
  assign new_n12783 = ~new_n12781 & ~new_n12782;
  assign new_n12784 = n6254 & n11478;
  assign new_n12785 = new_n12663 & ~new_n12668;
  assign new_n12786 = ~new_n12665 & ~new_n12785;
  assign new_n12787 = ~new_n12784 & new_n12786;
  assign new_n12788 = new_n12784 & ~new_n12786;
  assign new_n12789 = ~new_n12787 & ~new_n12788;
  assign new_n12790 = n137 & n7159;
  assign new_n12791 = n6294 & n12489;
  assign new_n12792 = ~new_n12652 & ~new_n12791;
  assign new_n12793 = new_n12652 & new_n12791;
  assign new_n12794 = ~new_n12792 & ~new_n12793;
  assign new_n12795 = new_n12790 & ~new_n12794;
  assign new_n12796 = ~new_n12790 & new_n12794;
  assign new_n12797 = ~new_n12795 & ~new_n12796;
  assign new_n12798 = ~new_n12789 & new_n12797;
  assign new_n12799 = new_n12789 & ~new_n12797;
  assign new_n12800 = ~new_n12798 & ~new_n12799;
  assign new_n12801 = new_n12783 & new_n12800;
  assign new_n12802 = ~new_n12783 & ~new_n12800;
  assign new_n12803 = ~new_n12801 & ~new_n12802;
  assign new_n12804 = new_n12683 & new_n12803;
  assign new_n12805 = ~new_n12683 & ~new_n12803;
  assign new_n12806 = ~new_n12804 & ~new_n12805;
  assign new_n12807_1 = n7236 & n12947;
  assign new_n12808 = ~new_n12706_1 & ~new_n12712;
  assign new_n12809 = ~new_n12711 & ~new_n12808;
  assign new_n12810 = new_n12807_1 & new_n12809;
  assign new_n12811 = ~new_n12807_1 & ~new_n12809;
  assign new_n12812 = ~new_n12810 & ~new_n12811;
  assign new_n12813 = n3992 & n11791;
  assign new_n12814 = new_n12697 & ~new_n12702;
  assign new_n12815 = ~new_n12699 & ~new_n12814;
  assign new_n12816 = ~new_n12813 & new_n12815;
  assign new_n12817 = new_n12813 & ~new_n12815;
  assign new_n12818 = ~new_n12816 & ~new_n12817;
  assign new_n12819 = n5760 & n6358;
  assign new_n12820 = n5198 & n10990;
  assign new_n12821 = ~new_n12686 & ~new_n12820;
  assign new_n12822 = new_n12686 & new_n12820;
  assign new_n12823 = ~new_n12821 & ~new_n12822;
  assign new_n12824 = new_n12819 & ~new_n12823;
  assign new_n12825 = ~new_n12819 & new_n12823;
  assign new_n12826_1 = ~new_n12824 & ~new_n12825;
  assign new_n12827 = ~new_n12818 & new_n12826_1;
  assign new_n12828 = new_n12818 & ~new_n12826_1;
  assign new_n12829 = ~new_n12827 & ~new_n12828;
  assign new_n12830 = ~new_n12812 & new_n12829;
  assign new_n12831 = new_n12812 & ~new_n12829;
  assign new_n12832 = ~new_n12830 & ~new_n12831;
  assign new_n12833 = new_n12717 & ~new_n12832;
  assign new_n12834 = ~new_n12717 & new_n12832;
  assign new_n12835 = ~new_n12833 & ~new_n12834;
  assign new_n12836 = ~new_n12806 & ~new_n12835;
  assign new_n12837 = new_n12806 & new_n12835;
  assign new_n12838 = ~new_n12836 & ~new_n12837;
  assign new_n12839 = ~new_n12720_1 & ~new_n12743;
  assign new_n12840 = ~new_n12721 & ~new_n12839;
  assign new_n12841 = ~new_n12838 & new_n12840;
  assign new_n12842 = new_n12838 & ~new_n12840;
  assign new_n12843 = ~new_n12841 & ~new_n12842;
  assign new_n12844 = ~new_n12777_1 & new_n12843;
  assign new_n12845 = ~new_n12776 & ~new_n12844;
  assign new_n12846 = ~new_n12647 & new_n12845;
  assign new_n12847 = new_n12647 & ~new_n12845;
  assign new_n12848 = n6441 & n7236;
  assign new_n12849 = n3992 & n12947;
  assign new_n12850 = n8384 & n11791;
  assign new_n12851 = new_n12849 & new_n12850;
  assign new_n12852 = ~new_n12849 & ~new_n12850;
  assign new_n12853 = ~new_n12851 & ~new_n12852;
  assign new_n12854 = ~new_n12816 & ~new_n12826_1;
  assign new_n12855 = ~new_n12817 & ~new_n12854;
  assign new_n12856 = ~new_n12853 & new_n12855;
  assign new_n12857 = new_n12853 & ~new_n12855;
  assign new_n12858 = ~new_n12856 & ~new_n12857;
  assign new_n12859 = n5198 & n5760;
  assign new_n12860 = n1471 & n10990;
  assign new_n12861 = ~new_n12859 & ~new_n12860;
  assign new_n12862 = new_n12859 & new_n12860;
  assign new_n12863 = ~new_n12861 & ~new_n12862;
  assign new_n12864 = new_n12698 & new_n12863;
  assign new_n12865 = ~new_n12698 & ~new_n12863;
  assign new_n12866 = ~new_n12864 & ~new_n12865;
  assign new_n12867 = new_n12819 & ~new_n12821;
  assign new_n12868 = ~new_n12822 & ~new_n12867;
  assign new_n12869 = ~new_n12866 & ~new_n12868;
  assign new_n12870 = new_n12866 & new_n12868;
  assign new_n12871 = ~new_n12869 & ~new_n12870;
  assign new_n12872 = new_n12858 & ~new_n12871;
  assign new_n12873 = ~new_n12858 & new_n12871;
  assign new_n12874 = ~new_n12872 & ~new_n12873;
  assign new_n12875 = ~new_n12810 & ~new_n12829;
  assign new_n12876 = ~new_n12811 & ~new_n12875;
  assign new_n12877 = new_n12874 & new_n12876;
  assign new_n12878 = ~new_n12874 & ~new_n12876;
  assign new_n12879 = ~new_n12877 & ~new_n12878;
  assign new_n12880 = new_n12848 & new_n12879;
  assign new_n12881 = ~new_n12848 & ~new_n12879;
  assign new_n12882 = ~new_n12880 & ~new_n12881;
  assign new_n12883 = new_n12833 & new_n12882;
  assign new_n12884 = ~new_n12833 & ~new_n12882;
  assign new_n12885 = ~new_n12883 & ~new_n12884;
  assign new_n12886 = n447 & n4805;
  assign new_n12887 = n11478 & n11967;
  assign new_n12888 = n5283 & n6254;
  assign new_n12889 = ~new_n12887 & ~new_n12888;
  assign new_n12890 = new_n12887 & new_n12888;
  assign new_n12891 = ~new_n12889 & ~new_n12890;
  assign new_n12892 = ~new_n12787 & ~new_n12797;
  assign new_n12893 = ~new_n12788 & ~new_n12892;
  assign new_n12894 = new_n12891 & ~new_n12893;
  assign new_n12895 = ~new_n12891 & new_n12893;
  assign new_n12896 = ~new_n12894 & ~new_n12895;
  assign new_n12897 = n6294 & n7159;
  assign new_n12898 = n6797 & n12489;
  assign new_n12899 = new_n12897 & new_n12898;
  assign new_n12900 = ~new_n12897 & ~new_n12898;
  assign new_n12901 = ~new_n12899 & ~new_n12900;
  assign new_n12902 = ~new_n12664 & ~new_n12901;
  assign new_n12903 = new_n12664 & new_n12901;
  assign new_n12904 = ~new_n12902 & ~new_n12903;
  assign new_n12905 = new_n12790 & ~new_n12792;
  assign new_n12906 = ~new_n12793 & ~new_n12905;
  assign new_n12907 = ~new_n12904 & new_n12906;
  assign new_n12908 = new_n12904 & ~new_n12906;
  assign new_n12909 = ~new_n12907 & ~new_n12908;
  assign new_n12910 = new_n12896 & ~new_n12909;
  assign new_n12911 = ~new_n12896 & new_n12909;
  assign new_n12912 = ~new_n12910 & ~new_n12911;
  assign new_n12913 = ~new_n12781 & new_n12800;
  assign new_n12914 = ~new_n12782 & ~new_n12913;
  assign new_n12915 = ~new_n12912 & ~new_n12914;
  assign new_n12916 = new_n12912 & new_n12914;
  assign new_n12917 = ~new_n12915 & ~new_n12916;
  assign new_n12918 = new_n12886 & new_n12917;
  assign new_n12919 = ~new_n12886 & ~new_n12917;
  assign new_n12920 = ~new_n12918 & ~new_n12919;
  assign new_n12921 = new_n12804 & new_n12920;
  assign new_n12922 = ~new_n12804 & ~new_n12920;
  assign new_n12923 = ~new_n12921 & ~new_n12922;
  assign new_n12924 = ~new_n12836 & ~new_n12840;
  assign new_n12925_1 = ~new_n12837 & ~new_n12924;
  assign new_n12926 = ~new_n12923 & new_n12925_1;
  assign new_n12927 = new_n12923 & ~new_n12925_1;
  assign new_n12928 = ~new_n12926 & ~new_n12927;
  assign new_n12929 = ~new_n12885 & ~new_n12928;
  assign new_n12930 = new_n12885 & new_n12928;
  assign new_n12931 = ~new_n12929 & ~new_n12930;
  assign new_n12932 = ~new_n12847 & ~new_n12931;
  assign new_n12933 = ~new_n12846 & ~new_n12932;
  assign new_n12934 = ~new_n12629 & new_n12633;
  assign new_n12935 = ~new_n12614 & ~new_n12934;
  assign new_n12936 = ~new_n12630 & new_n12935;
  assign new_n12937 = new_n12614 & new_n12934;
  assign new_n12938 = ~new_n12936 & ~new_n12937;
  assign new_n12939 = n8717 & n9400;
  assign new_n12940 = n2433 & n2464;
  assign new_n12941 = n6877 & n7730;
  assign new_n12942 = ~new_n12940 & ~new_n12941;
  assign new_n12943 = new_n12940 & new_n12941;
  assign new_n12944 = ~new_n12942 & ~new_n12943;
  assign new_n12945 = ~new_n12939 & ~new_n12944;
  assign new_n12946 = new_n12939 & new_n12944;
  assign new_n12947_1 = ~new_n12945 & ~new_n12946;
  assign new_n12948 = ~new_n12621 & new_n12625;
  assign new_n12949 = ~new_n12622 & ~new_n12948;
  assign new_n12950 = new_n12947_1 & new_n12949;
  assign new_n12951 = ~new_n12947_1 & ~new_n12949;
  assign new_n12952 = ~new_n12950 & ~new_n12951;
  assign new_n12953 = n8819 & n11311;
  assign new_n12954 = ~new_n12619 & ~new_n12953;
  assign new_n12955 = new_n12619 & new_n12953;
  assign new_n12956 = ~new_n12954 & ~new_n12955;
  assign new_n12957 = n4203 & n11728;
  assign new_n12958 = n12709 & n12753;
  assign new_n12959 = ~new_n12586 & ~new_n12958;
  assign new_n12960 = new_n12586 & new_n12958;
  assign new_n12961 = ~new_n12959 & ~new_n12960;
  assign new_n12962 = ~new_n12957 & ~new_n12961;
  assign new_n12963 = new_n12957 & new_n12961;
  assign new_n12964 = ~new_n12962 & ~new_n12963;
  assign new_n12965 = new_n12956 & ~new_n12964;
  assign new_n12966 = ~new_n12956 & new_n12964;
  assign new_n12967 = ~new_n12965 & ~new_n12966;
  assign new_n12968 = new_n12952 & new_n12967;
  assign new_n12969 = ~new_n12952 & ~new_n12967;
  assign new_n12970 = ~new_n12968 & ~new_n12969;
  assign new_n12971 = new_n12938 & new_n12970;
  assign new_n12972 = ~new_n12938 & ~new_n12970;
  assign new_n12973 = ~new_n12971 & ~new_n12972;
  assign new_n12974 = new_n12639 & ~new_n12973;
  assign new_n12975 = ~new_n12639 & new_n12973;
  assign new_n12976 = ~new_n12974 & ~new_n12975;
  assign new_n12977 = ~new_n12642 & ~new_n12645;
  assign new_n12978 = new_n12976 & ~new_n12977;
  assign new_n12979 = ~new_n12976 & new_n12977;
  assign new_n12980 = ~new_n12978 & ~new_n12979;
  assign new_n12981 = ~new_n12895 & new_n12909;
  assign new_n12982 = ~new_n12890 & ~new_n12981;
  assign new_n12983 = ~new_n12894 & new_n12982;
  assign new_n12984 = new_n12890 & new_n12981;
  assign new_n12985 = ~new_n12983 & ~new_n12984;
  assign new_n12986 = ~new_n12902 & ~new_n12906;
  assign new_n12987 = ~new_n12903 & ~new_n12986;
  assign new_n12988 = n5283 & n11967;
  assign new_n12989 = n1353 & n4805;
  assign new_n12990 = n447 & n11478;
  assign new_n12991 = ~new_n12989 & ~new_n12990;
  assign new_n12992 = new_n12989 & new_n12990;
  assign new_n12993 = ~new_n12991 & ~new_n12992;
  assign new_n12994 = new_n12988 & ~new_n12993;
  assign new_n12995 = ~new_n12988 & new_n12993;
  assign new_n12996 = ~new_n12994 & ~new_n12995;
  assign new_n12997 = ~new_n12987 & ~new_n12996;
  assign new_n12998 = new_n12987 & new_n12996;
  assign new_n12999 = ~new_n12997 & ~new_n12998;
  assign new_n13000 = n3146 & n12489;
  assign new_n13001 = n6294 & n12777;
  assign new_n13002 = n6797 & n7159;
  assign new_n13003 = ~new_n13001 & ~new_n13002;
  assign new_n13004 = new_n13001 & new_n13002;
  assign new_n13005 = ~new_n13003 & ~new_n13004;
  assign new_n13006 = new_n13000 & ~new_n13005;
  assign new_n13007 = ~new_n13000 & new_n13005;
  assign new_n13008 = ~new_n13006 & ~new_n13007;
  assign new_n13009 = n137 & n6254;
  assign new_n13010 = new_n12899 & new_n13009;
  assign new_n13011 = ~new_n12899 & ~new_n13009;
  assign new_n13012 = ~new_n13010 & ~new_n13011;
  assign new_n13013 = ~new_n13008 & new_n13012;
  assign new_n13014 = new_n13008 & ~new_n13012;
  assign new_n13015 = ~new_n13013 & ~new_n13014;
  assign new_n13016 = new_n12999 & ~new_n13015;
  assign new_n13017 = ~new_n12999 & new_n13015;
  assign new_n13018 = ~new_n13016 & ~new_n13017;
  assign new_n13019 = new_n12985 & new_n13018;
  assign new_n13020 = ~new_n12985 & ~new_n13018;
  assign new_n13021 = ~new_n13019 & ~new_n13020;
  assign new_n13022 = ~new_n12915 & new_n13021;
  assign new_n13023 = new_n12915 & ~new_n13021;
  assign new_n13024 = ~new_n13022 & ~new_n13023;
  assign new_n13025 = ~new_n12918 & ~new_n12921;
  assign new_n13026 = ~new_n13024 & new_n13025;
  assign new_n13027 = new_n13024 & ~new_n13025;
  assign new_n13028 = ~new_n13026 & ~new_n13027;
  assign new_n13029 = ~new_n12856 & ~new_n12871;
  assign new_n13030 = new_n12851 & new_n13029;
  assign new_n13031 = ~new_n12851 & ~new_n13029;
  assign new_n13032 = ~new_n12857 & new_n13031;
  assign new_n13033 = ~new_n13030 & ~new_n13032;
  assign new_n13034 = n3992 & n6441;
  assign new_n13035 = n8384 & n12947;
  assign new_n13036 = n7236 & n11999;
  assign new_n13037 = ~new_n13035 & ~new_n13036;
  assign new_n13038 = new_n13035 & new_n13036;
  assign new_n13039 = ~new_n13037 & ~new_n13038;
  assign new_n13040 = ~new_n13034 & ~new_n13039;
  assign new_n13041 = new_n13034 & new_n13039;
  assign new_n13042 = ~new_n13040 & ~new_n13041;
  assign new_n13043 = ~new_n12864 & new_n12868;
  assign new_n13044 = ~new_n12865 & ~new_n13043;
  assign new_n13045 = new_n13042 & new_n13044;
  assign new_n13046 = ~new_n13042 & ~new_n13044;
  assign new_n13047 = ~new_n13045 & ~new_n13046;
  assign new_n13048 = n6358 & n11791;
  assign new_n13049 = ~new_n12862 & ~new_n13048;
  assign new_n13050 = new_n12862 & new_n13048;
  assign new_n13051 = ~new_n13049 & ~new_n13050;
  assign new_n13052 = n1471 & n5760;
  assign new_n13053 = n1478 & n5198;
  assign new_n13054 = n7646 & n10990;
  assign new_n13055 = ~new_n13053 & ~new_n13054;
  assign new_n13056 = new_n13053 & new_n13054;
  assign new_n13057 = ~new_n13055 & ~new_n13056;
  assign new_n13058 = ~new_n13052 & ~new_n13057;
  assign new_n13059 = new_n13052 & new_n13057;
  assign new_n13060 = ~new_n13058 & ~new_n13059;
  assign new_n13061 = new_n13051 & ~new_n13060;
  assign new_n13062 = ~new_n13051 & new_n13060;
  assign new_n13063 = ~new_n13061 & ~new_n13062;
  assign new_n13064 = new_n13047 & new_n13063;
  assign new_n13065 = ~new_n13047 & ~new_n13063;
  assign new_n13066 = ~new_n13064 & ~new_n13065;
  assign new_n13067 = ~new_n13033 & ~new_n13066;
  assign new_n13068 = new_n13033 & new_n13066;
  assign new_n13069 = ~new_n13067 & ~new_n13068;
  assign new_n13070 = new_n12877 & ~new_n13069;
  assign new_n13071 = ~new_n12877 & new_n13069;
  assign new_n13072 = ~new_n13070 & ~new_n13071;
  assign new_n13073 = ~new_n12880 & ~new_n12883;
  assign new_n13074 = new_n13072 & ~new_n13073;
  assign new_n13075 = ~new_n13072 & new_n13073;
  assign new_n13076 = ~new_n13074 & ~new_n13075;
  assign new_n13077 = ~new_n13028 & ~new_n13076;
  assign new_n13078 = new_n13028 & new_n13076;
  assign new_n13079 = ~new_n13077 & ~new_n13078;
  assign new_n13080 = new_n12885 & ~new_n12926;
  assign new_n13081 = ~new_n12927 & ~new_n13080;
  assign new_n13082 = ~new_n13079 & ~new_n13081;
  assign new_n13083 = new_n13079 & new_n13081;
  assign new_n13084 = ~new_n13082 & ~new_n13083;
  assign new_n13085 = ~new_n12980 & new_n13084;
  assign new_n13086 = new_n12980 & ~new_n13084;
  assign new_n13087 = ~new_n13085 & ~new_n13086;
  assign new_n13088 = ~new_n12933 & ~new_n13087;
  assign new_n13089 = new_n12933 & new_n13087;
  assign new_n13090 = ~new_n13088 & ~new_n13089;
  assign new_n13091 = ~new_n12549 & ~new_n13090;
  assign new_n13092 = new_n12549 & new_n13090;
  assign new_n13093 = ~new_n12499 & ~new_n12501;
  assign new_n13094 = ~new_n12502 & ~new_n13093;
  assign new_n13095 = ~new_n12494 & ~new_n12498;
  assign new_n13096 = ~new_n12499 & ~new_n13095;
  assign new_n13097 = ~new_n12776 & ~new_n12777_1;
  assign new_n13098 = new_n12843 & new_n13097;
  assign new_n13099 = ~new_n12843 & ~new_n13097;
  assign new_n13100 = ~new_n13098 & ~new_n13099;
  assign new_n13101 = ~new_n13096 & ~new_n13100;
  assign new_n13102 = new_n13096 & new_n13100;
  assign new_n13103 = ~new_n12489_1 & new_n12493;
  assign new_n13104 = ~new_n12494 & ~new_n13103;
  assign new_n13105 = ~new_n12747 & ~new_n12748;
  assign new_n13106 = new_n12773 & ~new_n13105;
  assign new_n13107 = ~new_n12773 & new_n13105;
  assign new_n13108 = ~new_n13106 & ~new_n13107;
  assign new_n13109 = new_n13104 & ~new_n13108;
  assign new_n13110 = ~new_n13104 & new_n13108;
  assign new_n13111 = ~new_n12484 & ~new_n12488;
  assign new_n13112 = ~new_n12489_1 & ~new_n13111;
  assign new_n13113 = ~new_n12757 & ~new_n12758;
  assign new_n13114 = ~new_n12771 & ~new_n13113;
  assign new_n13115 = new_n12771 & new_n13113;
  assign new_n13116 = ~new_n13114 & ~new_n13115;
  assign new_n13117 = new_n13112 & ~new_n13116;
  assign new_n13118 = ~new_n13112 & new_n13116;
  assign new_n13119 = n7862 & n11407;
  assign new_n13120 = ~new_n12551 & ~new_n12768;
  assign new_n13121 = ~new_n12769 & ~new_n13120;
  assign new_n13122 = new_n13119 & new_n13121;
  assign new_n13123 = ~new_n12436 & ~new_n12483;
  assign new_n13124 = ~new_n12484 & ~new_n13123;
  assign new_n13125 = new_n13122 & new_n13124;
  assign new_n13126 = ~new_n13122 & ~new_n13124;
  assign new_n13127 = ~new_n12765 & ~new_n12766;
  assign new_n13128 = ~new_n12769 & ~new_n13127;
  assign new_n13129 = new_n12769 & new_n13127;
  assign new_n13130 = ~new_n13128 & ~new_n13129;
  assign new_n13131 = ~new_n13126 & new_n13130;
  assign new_n13132 = ~new_n13125 & ~new_n13131;
  assign new_n13133 = ~new_n13118 & ~new_n13132;
  assign new_n13134 = ~new_n13117 & ~new_n13133;
  assign new_n13135 = ~new_n13110 & ~new_n13134;
  assign new_n13136 = ~new_n13109 & ~new_n13135;
  assign new_n13137 = ~new_n13102 & new_n13136;
  assign new_n13138 = ~new_n13101 & ~new_n13137;
  assign new_n13139 = ~new_n13094 & ~new_n13138;
  assign new_n13140 = new_n13094 & new_n13138;
  assign new_n13141 = ~new_n12846 & ~new_n12847;
  assign new_n13142 = ~new_n12931 & ~new_n13141;
  assign new_n13143 = new_n12931 & new_n13141;
  assign new_n13144 = ~new_n13142 & ~new_n13143;
  assign new_n13145 = ~new_n13140 & ~new_n13144;
  assign new_n13146 = ~new_n13139 & ~new_n13145;
  assign new_n13147 = ~new_n13092 & ~new_n13146;
  assign new_n13148 = ~new_n13091 & ~new_n13147;
  assign new_n13149 = new_n12933 & ~new_n13085;
  assign new_n13150 = ~new_n13086 & ~new_n13149;
  assign new_n13151 = ~new_n13077 & ~new_n13081;
  assign new_n13152 = ~new_n13078 & ~new_n13151;
  assign new_n13153 = ~new_n13070 & ~new_n13074;
  assign new_n13154 = n1471 & n1478;
  assign new_n13155 = n5760 & n7646;
  assign new_n13156 = ~new_n13154 & ~new_n13155;
  assign new_n13157 = new_n13154 & new_n13155;
  assign new_n13158 = ~new_n13156 & ~new_n13157;
  assign new_n13159 = n7236 & n10022;
  assign new_n13160 = n4722 & n10990;
  assign new_n13161 = new_n13159 & ~new_n13160;
  assign new_n13162 = ~new_n13159 & new_n13160;
  assign new_n13163 = ~new_n13161 & ~new_n13162;
  assign new_n13164 = ~new_n13158 & ~new_n13163;
  assign new_n13165 = new_n13158 & new_n13163;
  assign new_n13166 = ~new_n13164 & ~new_n13165;
  assign new_n13167 = ~new_n12939 & ~new_n12943;
  assign new_n13168 = ~new_n12942 & ~new_n13167;
  assign new_n13169 = ~new_n13166 & ~new_n13168;
  assign new_n13170 = new_n13166 & new_n13168;
  assign new_n13171 = ~new_n13169 & ~new_n13170;
  assign new_n13172 = new_n13153 & new_n13171;
  assign new_n13173 = ~new_n13153 & ~new_n13171;
  assign new_n13174 = ~new_n13172 & ~new_n13173;
  assign new_n13175 = new_n13152 & ~new_n13174;
  assign new_n13176 = ~new_n13152 & new_n13174;
  assign new_n13177 = ~new_n13175 & ~new_n13176;
  assign new_n13178 = ~new_n12974 & ~new_n12978;
  assign new_n13179 = ~new_n12521 & new_n12537;
  assign new_n13180 = ~new_n12520 & ~new_n13179;
  assign new_n13181 = ~new_n12524 & ~new_n12534;
  assign new_n13182 = ~new_n12525 & ~new_n13181;
  assign new_n13183 = n11821 & n11877;
  assign new_n13184 = n5212 & n9080;
  assign new_n13185 = ~new_n13183 & new_n13184;
  assign new_n13186 = new_n13183 & ~new_n13184;
  assign new_n13187 = ~new_n13185 & ~new_n13186;
  assign new_n13188 = n1333 & n9725;
  assign new_n13189 = n5320 & n11757;
  assign new_n13190 = n4370 & n5240;
  assign new_n13191 = new_n13189 & new_n13190;
  assign new_n13192 = ~new_n13189 & ~new_n13190;
  assign new_n13193 = ~new_n13191 & ~new_n13192;
  assign new_n13194 = new_n13188 & ~new_n13193;
  assign new_n13195 = ~new_n13188 & new_n13193;
  assign new_n13196 = ~new_n13194 & ~new_n13195;
  assign new_n13197 = ~new_n13187 & ~new_n13196;
  assign new_n13198 = new_n13187 & new_n13196;
  assign new_n13199 = ~new_n13197 & ~new_n13198;
  assign new_n13200 = ~new_n13182 & ~new_n13199;
  assign new_n13201 = new_n13182 & new_n13199;
  assign new_n13202 = ~new_n13200 & ~new_n13201;
  assign new_n13203 = n3172 & n12000;
  assign new_n13204 = ~new_n12527 & ~new_n12529;
  assign new_n13205 = ~new_n12530 & ~new_n13204;
  assign new_n13206 = ~new_n13203 & new_n13205;
  assign new_n13207 = new_n13203 & ~new_n13205;
  assign new_n13208 = ~new_n13206 & ~new_n13207;
  assign new_n13209 = ~new_n12509 & ~new_n12513;
  assign new_n13210 = ~new_n12512 & ~new_n13209;
  assign new_n13211 = ~new_n13208 & new_n13210;
  assign new_n13212 = new_n13208 & ~new_n13210;
  assign new_n13213 = ~new_n13211 & ~new_n13212;
  assign new_n13214 = new_n13202 & ~new_n13213;
  assign new_n13215 = ~new_n13202 & new_n13213;
  assign new_n13216 = ~new_n13214 & ~new_n13215;
  assign new_n13217 = ~new_n12936 & ~new_n12970;
  assign new_n13218 = ~new_n12937 & ~new_n13217;
  assign new_n13219 = n11728 & n12753;
  assign new_n13220 = n10174 & n12709;
  assign new_n13221 = n1198 & n6877;
  assign new_n13222 = new_n13220 & ~new_n13221;
  assign new_n13223 = ~new_n13220 & new_n13221;
  assign new_n13224 = ~new_n13222 & ~new_n13223;
  assign new_n13225 = new_n13219 & ~new_n13224;
  assign new_n13226 = ~new_n13219 & new_n13224;
  assign new_n13227 = ~new_n13225 & ~new_n13226;
  assign new_n13228 = new_n13218 & new_n13227;
  assign new_n13229 = ~new_n13218 & ~new_n13227;
  assign new_n13230 = ~new_n13228 & ~new_n13229;
  assign new_n13231 = ~new_n13216 & new_n13230;
  assign new_n13232 = new_n13216 & ~new_n13230;
  assign new_n13233 = ~new_n13231 & ~new_n13232;
  assign new_n13234 = ~new_n13180 & new_n13233;
  assign new_n13235 = new_n13180 & ~new_n13233;
  assign new_n13236 = ~new_n13234 & ~new_n13235;
  assign new_n13237 = ~new_n12955 & ~new_n12964;
  assign new_n13238 = ~new_n12954 & ~new_n13237;
  assign new_n13239 = ~new_n12957 & ~new_n12960;
  assign new_n13240 = ~new_n12959 & ~new_n13239;
  assign new_n13241 = n7730 & n9400;
  assign new_n13242 = n2433 & n11311;
  assign new_n13243 = new_n13241 & ~new_n13242;
  assign new_n13244 = ~new_n13241 & new_n13242;
  assign new_n13245 = ~new_n13243 & ~new_n13244;
  assign new_n13246 = ~new_n13240 & new_n13245;
  assign new_n13247 = new_n13240 & ~new_n13245;
  assign new_n13248 = ~new_n13246 & ~new_n13247;
  assign new_n13249 = new_n13238 & ~new_n13248;
  assign new_n13250 = ~new_n13238 & new_n13248;
  assign new_n13251 = ~new_n13249 & ~new_n13250;
  assign new_n13252 = ~new_n12951 & ~new_n12967;
  assign new_n13253 = ~new_n12950 & ~new_n13252;
  assign new_n13254 = n2464 & n8717;
  assign new_n13255 = n4187 & n8819;
  assign new_n13256 = n4203 & n6429;
  assign new_n13257 = ~new_n13255 & new_n13256;
  assign new_n13258 = new_n13255 & ~new_n13256;
  assign new_n13259 = ~new_n13257 & ~new_n13258;
  assign new_n13260 = new_n13254 & new_n13259;
  assign new_n13261 = ~new_n13254 & ~new_n13259;
  assign new_n13262 = ~new_n13260 & ~new_n13261;
  assign new_n13263 = new_n13253 & ~new_n13262;
  assign new_n13264 = ~new_n13253 & new_n13262;
  assign new_n13265 = ~new_n13263 & ~new_n13264;
  assign new_n13266 = ~new_n13251 & ~new_n13265;
  assign new_n13267 = new_n13251 & new_n13265;
  assign new_n13268 = ~new_n13266 & ~new_n13267;
  assign new_n13269 = ~new_n13032 & ~new_n13066;
  assign new_n13270 = ~new_n13030 & ~new_n13269;
  assign new_n13271 = ~new_n13268 & new_n13270;
  assign new_n13272 = new_n13268 & ~new_n13270;
  assign new_n13273 = ~new_n13271 & ~new_n13272;
  assign new_n13274 = ~new_n13236 & new_n13273;
  assign new_n13275 = new_n13236 & ~new_n13273;
  assign new_n13276 = ~new_n13274 & ~new_n13275;
  assign new_n13277 = new_n13178 & new_n13276;
  assign new_n13278 = ~new_n13178 & ~new_n13276;
  assign new_n13279 = ~new_n13277 & ~new_n13278;
  assign new_n13280 = new_n13177 & ~new_n13279;
  assign new_n13281 = ~new_n13177 & new_n13279;
  assign new_n13282 = ~new_n13280 & ~new_n13281;
  assign new_n13283 = ~new_n13150 & new_n13282;
  assign new_n13284 = new_n13150 & ~new_n13282;
  assign new_n13285 = ~new_n13283 & ~new_n13284;
  assign new_n13286 = ~new_n12544 & ~new_n12547;
  assign new_n13287 = n6604 & n7862;
  assign new_n13288 = n6826 & n11407;
  assign new_n13289 = ~new_n13287 & new_n13288;
  assign new_n13290 = new_n13287 & ~new_n13288;
  assign new_n13291 = ~new_n13289 & ~new_n13290;
  assign new_n13292 = new_n13000 & ~new_n13003;
  assign new_n13293 = ~new_n13004 & ~new_n13292;
  assign new_n13294 = n1353 & n11478;
  assign new_n13295 = n447 & n5283;
  assign new_n13296 = ~new_n13294 & new_n13295;
  assign new_n13297 = new_n13294 & ~new_n13295;
  assign new_n13298 = ~new_n13296 & ~new_n13297;
  assign new_n13299 = new_n13293 & ~new_n13298;
  assign new_n13300 = ~new_n13293 & new_n13298;
  assign new_n13301 = ~new_n13299 & ~new_n13300;
  assign new_n13302 = ~new_n13291 & new_n13301;
  assign new_n13303 = new_n13291 & ~new_n13301;
  assign new_n13304 = ~new_n13302 & ~new_n13303;
  assign new_n13305 = ~new_n12506 & new_n12540;
  assign new_n13306 = ~new_n12507 & ~new_n13305;
  assign new_n13307 = new_n13008 & ~new_n13010;
  assign new_n13308 = ~new_n13011 & ~new_n13307;
  assign new_n13309 = new_n13306 & new_n13308;
  assign new_n13310 = ~new_n13306 & ~new_n13308;
  assign new_n13311 = ~new_n13309 & ~new_n13310;
  assign new_n13312 = new_n13304 & new_n13311;
  assign new_n13313 = ~new_n13304 & ~new_n13311;
  assign new_n13314 = ~new_n13312 & ~new_n13313;
  assign new_n13315 = ~new_n13286 & new_n13314;
  assign new_n13316 = new_n13286 & ~new_n13314;
  assign new_n13317 = ~new_n13315 & ~new_n13316;
  assign new_n13318 = ~new_n12998 & new_n13015;
  assign new_n13319 = ~new_n12997 & ~new_n13318;
  assign new_n13320 = ~new_n13023 & ~new_n13027;
  assign new_n13321 = ~new_n12988 & ~new_n12992;
  assign new_n13322 = ~new_n12991 & ~new_n13321;
  assign new_n13323 = ~new_n13045 & new_n13063;
  assign new_n13324 = ~new_n13046 & ~new_n13323;
  assign new_n13325 = n4436 & n4805;
  assign new_n13326 = n137 & n11967;
  assign new_n13327 = n6254 & n6294;
  assign new_n13328 = ~new_n13326 & ~new_n13327;
  assign new_n13329 = new_n13326 & new_n13327;
  assign new_n13330 = ~new_n13328 & ~new_n13329;
  assign new_n13331 = n6797 & n12777;
  assign new_n13332 = n3146 & n7159;
  assign new_n13333 = new_n13331 & ~new_n13332;
  assign new_n13334 = ~new_n13331 & new_n13332;
  assign new_n13335 = ~new_n13333 & ~new_n13334;
  assign new_n13336 = ~new_n13330 & ~new_n13335;
  assign new_n13337 = new_n13330 & new_n13335;
  assign new_n13338 = ~new_n13336 & ~new_n13337;
  assign new_n13339 = new_n13325 & ~new_n13338;
  assign new_n13340 = ~new_n13325 & new_n13338;
  assign new_n13341 = ~new_n13339 & ~new_n13340;
  assign new_n13342 = ~new_n13324 & ~new_n13341;
  assign new_n13343 = new_n13324 & new_n13341;
  assign new_n13344 = ~new_n13342 & ~new_n13343;
  assign new_n13345 = ~new_n12983 & ~new_n13018;
  assign new_n13346 = ~new_n12984 & ~new_n13345;
  assign new_n13347 = new_n13344 & new_n13346;
  assign new_n13348 = ~new_n13344 & ~new_n13346;
  assign new_n13349 = ~new_n13347 & ~new_n13348;
  assign new_n13350 = n4938 & n12489;
  assign new_n13351 = n3992 & n11999;
  assign new_n13352 = n6441 & n8384;
  assign new_n13353 = ~new_n13351 & ~new_n13352;
  assign new_n13354 = new_n13351 & new_n13352;
  assign new_n13355 = ~new_n13353 & ~new_n13354;
  assign new_n13356 = n6358 & n12947;
  assign new_n13357 = n5198 & n11791;
  assign new_n13358 = new_n13356 & ~new_n13357;
  assign new_n13359 = ~new_n13356 & new_n13357;
  assign new_n13360 = ~new_n13358 & ~new_n13359;
  assign new_n13361 = ~new_n13355 & ~new_n13360;
  assign new_n13362 = new_n13355 & new_n13360;
  assign new_n13363 = ~new_n13361 & ~new_n13362;
  assign new_n13364 = ~new_n13052 & ~new_n13056;
  assign new_n13365 = ~new_n13055 & ~new_n13364;
  assign new_n13366 = ~new_n13034 & ~new_n13038;
  assign new_n13367 = ~new_n13037 & ~new_n13366;
  assign new_n13368 = ~new_n13365 & new_n13367;
  assign new_n13369 = new_n13365 & ~new_n13367;
  assign new_n13370 = ~new_n13368 & ~new_n13369;
  assign new_n13371 = new_n13363 & new_n13370;
  assign new_n13372 = ~new_n13363 & ~new_n13370;
  assign new_n13373 = ~new_n13371 & ~new_n13372;
  assign new_n13374 = ~new_n13049 & new_n13060;
  assign new_n13375 = ~new_n13050 & ~new_n13374;
  assign new_n13376 = ~new_n13373 & new_n13375;
  assign new_n13377 = new_n13373 & ~new_n13375;
  assign new_n13378 = ~new_n13376 & ~new_n13377;
  assign new_n13379 = ~new_n13350 & new_n13378;
  assign new_n13380 = new_n13350 & ~new_n13378;
  assign new_n13381 = ~new_n13379 & ~new_n13380;
  assign new_n13382 = new_n13349 & ~new_n13381;
  assign new_n13383 = ~new_n13349 & new_n13381;
  assign new_n13384 = ~new_n13382 & ~new_n13383;
  assign new_n13385 = ~new_n13322 & new_n13384;
  assign new_n13386 = new_n13322 & ~new_n13384;
  assign new_n13387 = ~new_n13385 & ~new_n13386;
  assign new_n13388 = new_n13320 & new_n13387;
  assign new_n13389 = ~new_n13320 & ~new_n13387;
  assign new_n13390 = ~new_n13388 & ~new_n13389;
  assign new_n13391 = ~new_n13319 & ~new_n13390;
  assign new_n13392 = new_n13319 & new_n13390;
  assign new_n13393 = ~new_n13391 & ~new_n13392;
  assign new_n13394 = ~new_n13317 & ~new_n13393;
  assign new_n13395 = new_n13317 & new_n13393;
  assign new_n13396 = ~new_n13394 & ~new_n13395;
  assign new_n13397 = ~new_n13285 & new_n13396;
  assign new_n13398 = new_n13285 & ~new_n13396;
  assign new_n13399 = ~new_n13397 & ~new_n13398;
  assign new_n13400 = new_n13148 & ~new_n13399;
  assign new_n13401 = ~new_n13148 & new_n13399;
  assign n4378 = new_n13400 | new_n13401;
  assign new_n13403 = ~new_n4452 & ~new_n4454;
  assign n4397 = ~new_n4455 & ~new_n13403;
  assign new_n13405 = ~new_n4784 & ~new_n4786;
  assign n4553 = ~new_n4787 & ~new_n13405;
  assign new_n13407 = ~new_n950 & ~new_n952;
  assign n4686 = ~new_n953 & ~new_n13407;
  assign new_n13409 = ~new_n10989 & ~new_n10990_1;
  assign new_n13410 = new_n11010 & ~new_n13409;
  assign new_n13411 = ~new_n11010 & new_n13409;
  assign n4689 = ~new_n13410 & ~new_n13411;
  assign new_n13413 = ~new_n5677 & ~new_n5678;
  assign new_n13414 = ~new_n5682 & new_n13413;
  assign new_n13415 = new_n5682 & ~new_n13413;
  assign n4733 = new_n13414 | new_n13415;
  assign new_n13417 = ~new_n2314 & ~new_n2315;
  assign new_n13418 = new_n2325 & ~new_n13417;
  assign new_n13419 = ~new_n2325 & new_n13417;
  assign n4757 = ~new_n13418 & ~new_n13419;
  assign new_n13421 = ~new_n5647 & ~new_n5648;
  assign new_n13422 = new_n5672 & ~new_n13421;
  assign new_n13423 = ~new_n5672 & new_n13421;
  assign n4971 = ~new_n13422 & ~new_n13423;
  assign new_n13425 = ~new_n7619 & ~new_n7620;
  assign new_n13426 = new_n7622 & ~new_n13425;
  assign new_n13427 = ~new_n7622 & new_n13425;
  assign n5030 = ~new_n13426 & ~new_n13427;
  assign new_n13429 = ~new_n3289 & ~new_n3290;
  assign new_n13430 = new_n3324 & ~new_n13429;
  assign new_n13431 = ~new_n3324 & new_n13429;
  assign n5034 = ~new_n13430 & ~new_n13431;
  assign new_n13433 = ~new_n3305 & ~new_n3306;
  assign new_n13434 = new_n3320 & ~new_n13433;
  assign new_n13435 = ~new_n3320 & new_n13433;
  assign n5094 = ~new_n13434 & ~new_n13435;
  assign new_n13437 = ~new_n12266 & new_n12285;
  assign new_n13438 = ~new_n12267 & ~new_n13437;
  assign new_n13439 = n2564 & n5320;
  assign new_n13440 = n4189 & n4370;
  assign new_n13441 = ~new_n13439 & ~new_n13440;
  assign new_n13442 = new_n13439 & new_n13440;
  assign new_n13443 = ~new_n13441 & ~new_n13442;
  assign new_n13444 = ~new_n12273 & ~new_n12282;
  assign new_n13445 = ~new_n12272 & ~new_n13444;
  assign new_n13446 = new_n13443 & ~new_n13445;
  assign new_n13447 = ~new_n13443 & new_n13445;
  assign new_n13448 = ~new_n13446 & ~new_n13447;
  assign new_n13449 = n6770 & n11877;
  assign new_n13450 = new_n12275 & ~new_n12277;
  assign new_n13451 = ~new_n12278 & ~new_n13450;
  assign new_n13452 = ~new_n13449 & new_n13451;
  assign new_n13453 = new_n13449 & ~new_n13451;
  assign new_n13454 = n5212 & n9920;
  assign new_n13455 = n3627 & n11407;
  assign new_n13456 = ~new_n13454 & ~new_n13455;
  assign new_n13457 = new_n13454 & new_n13455;
  assign new_n13458 = ~new_n13456 & ~new_n13457;
  assign new_n13459 = ~new_n13453 & ~new_n13458;
  assign new_n13460 = ~new_n13452 & new_n13459;
  assign new_n13461 = ~new_n13452 & ~new_n13453;
  assign new_n13462 = new_n13458 & ~new_n13461;
  assign new_n13463 = ~new_n13460 & ~new_n13462;
  assign new_n13464 = new_n13448 & new_n13463;
  assign new_n13465 = ~new_n13448 & ~new_n13463;
  assign new_n13466 = ~new_n13464 & ~new_n13465;
  assign new_n13467 = new_n13438 & ~new_n13466;
  assign new_n13468 = ~new_n13447 & ~new_n13463;
  assign new_n13469 = ~new_n13442 & ~new_n13468;
  assign new_n13470 = ~new_n13446 & new_n13469;
  assign new_n13471 = new_n13442 & new_n13468;
  assign new_n13472 = ~new_n13470 & ~new_n13471;
  assign new_n13473 = ~new_n13452 & ~new_n13459;
  assign new_n13474 = n4189 & n5320;
  assign new_n13475 = n6687 & n9725;
  assign new_n13476 = n2564 & n12000;
  assign new_n13477 = ~new_n13475 & ~new_n13476;
  assign new_n13478 = new_n13475 & new_n13476;
  assign new_n13479 = ~new_n13477 & ~new_n13478;
  assign new_n13480 = new_n13474 & ~new_n13479;
  assign new_n13481 = ~new_n13474 & new_n13479;
  assign new_n13482 = ~new_n13480 & ~new_n13481;
  assign new_n13483 = new_n13473 & ~new_n13482;
  assign new_n13484 = ~new_n13473 & new_n13482;
  assign new_n13485 = ~new_n13483 & ~new_n13484;
  assign new_n13486 = n4370 & n6770;
  assign new_n13487 = ~new_n13457 & ~new_n13486;
  assign new_n13488 = new_n13457 & new_n13486;
  assign new_n13489 = ~new_n13487 & ~new_n13488;
  assign new_n13490 = n4516 & n11407;
  assign new_n13491 = n9920 & n11877;
  assign new_n13492 = n3627 & n5212;
  assign new_n13493 = ~new_n13491 & ~new_n13492;
  assign new_n13494 = new_n13491 & new_n13492;
  assign new_n13495 = ~new_n13493 & ~new_n13494;
  assign new_n13496 = new_n13490 & ~new_n13495;
  assign new_n13497 = ~new_n13490 & new_n13495;
  assign new_n13498 = ~new_n13496 & ~new_n13497;
  assign new_n13499 = new_n13489 & new_n13498;
  assign new_n13500 = ~new_n13489 & ~new_n13498;
  assign new_n13501 = ~new_n13499 & ~new_n13500;
  assign new_n13502 = new_n13485 & ~new_n13501;
  assign new_n13503 = ~new_n13485 & new_n13501;
  assign new_n13504 = ~new_n13502 & ~new_n13503;
  assign new_n13505 = new_n13472 & ~new_n13504;
  assign new_n13506 = ~new_n13472 & new_n13504;
  assign new_n13507 = ~new_n13505 & ~new_n13506;
  assign new_n13508 = ~new_n13467 & new_n13507;
  assign new_n13509 = new_n13467 & ~new_n13507;
  assign new_n13510 = ~new_n13508 & ~new_n13509;
  assign new_n13511 = n6687 & n12000;
  assign new_n13512 = ~new_n13438 & new_n13466;
  assign new_n13513 = ~new_n13467 & ~new_n13512;
  assign new_n13514 = new_n13511 & new_n13513;
  assign new_n13515 = ~new_n13511 & ~new_n13513;
  assign new_n13516 = ~new_n13514 & ~new_n13515;
  assign new_n13517 = new_n12289 & new_n13516;
  assign new_n13518 = ~new_n13514 & ~new_n13517;
  assign new_n13519 = ~new_n13510 & new_n13518;
  assign new_n13520 = new_n13510 & ~new_n13518;
  assign new_n13521 = ~new_n13519 & ~new_n13520;
  assign new_n13522 = n8336 & n8717;
  assign new_n13523 = ~new_n12312 & new_n12315;
  assign new_n13524 = ~new_n12311 & ~new_n13523;
  assign new_n13525 = n2433 & n10928;
  assign new_n13526 = n6986 & n8819;
  assign new_n13527 = ~new_n13525 & ~new_n13526;
  assign new_n13528 = new_n13525 & new_n13526;
  assign new_n13529 = ~new_n13527 & ~new_n13528;
  assign new_n13530 = n2226 & n6429;
  assign new_n13531 = n1094 & n11728;
  assign new_n13532 = n10678 & n12709;
  assign new_n13533 = ~new_n13531 & ~new_n13532;
  assign new_n13534 = new_n13531 & new_n13532;
  assign new_n13535 = ~new_n13533 & ~new_n13534;
  assign new_n13536 = new_n13530 & new_n13535;
  assign new_n13537 = ~new_n13530 & ~new_n13535;
  assign new_n13538 = ~new_n13536 & ~new_n13537;
  assign new_n13539 = new_n12299_1 & ~new_n12302;
  assign new_n13540 = ~new_n12303 & ~new_n13539;
  assign new_n13541 = ~new_n13538 & ~new_n13540;
  assign new_n13542 = new_n13538 & new_n13540;
  assign new_n13543 = ~new_n13541 & ~new_n13542;
  assign new_n13544 = new_n13529 & ~new_n13543;
  assign new_n13545 = ~new_n13529 & new_n13543;
  assign new_n13546 = ~new_n13544 & ~new_n13545;
  assign new_n13547 = ~new_n12296 & ~new_n12307;
  assign new_n13548 = ~new_n12297 & ~new_n13547;
  assign new_n13549 = new_n13546 & new_n13548;
  assign new_n13550 = ~new_n13546 & ~new_n13548;
  assign new_n13551 = ~new_n13549 & ~new_n13550;
  assign new_n13552 = ~new_n13524 & ~new_n13551;
  assign new_n13553 = new_n13524 & new_n13551;
  assign new_n13554 = ~new_n13552 & ~new_n13553;
  assign new_n13555 = new_n13522 & new_n13554;
  assign new_n13556 = ~new_n13522 & ~new_n13554;
  assign new_n13557 = ~new_n13555 & ~new_n13556;
  assign new_n13558 = new_n12319 & new_n13557;
  assign new_n13559 = ~new_n13555 & ~new_n13558;
  assign new_n13560 = ~new_n13545 & ~new_n13548;
  assign new_n13561 = ~new_n13528 & ~new_n13560;
  assign new_n13562 = ~new_n13544 & new_n13561;
  assign new_n13563 = new_n13528 & new_n13560;
  assign new_n13564 = ~new_n13562 & ~new_n13563;
  assign new_n13565 = n8717 & n10928;
  assign new_n13566 = n2433 & n6986;
  assign new_n13567 = n7730 & n8336;
  assign new_n13568 = ~new_n13566 & ~new_n13567;
  assign new_n13569 = new_n13566 & new_n13567;
  assign new_n13570 = ~new_n13568 & ~new_n13569;
  assign new_n13571 = ~new_n13565 & ~new_n13570;
  assign new_n13572 = new_n13565 & new_n13570;
  assign new_n13573 = ~new_n13571 & ~new_n13572;
  assign new_n13574 = ~new_n13537 & ~new_n13540;
  assign new_n13575 = ~new_n13536 & ~new_n13574;
  assign new_n13576 = new_n13573 & ~new_n13575;
  assign new_n13577 = ~new_n13573 & new_n13575;
  assign new_n13578 = ~new_n13576 & ~new_n13577;
  assign new_n13579 = n2226 & n8819;
  assign new_n13580 = ~new_n13534 & ~new_n13579;
  assign new_n13581 = new_n13534 & new_n13579;
  assign new_n13582 = ~new_n13580 & ~new_n13581;
  assign new_n13583 = n10678 & n11728;
  assign new_n13584 = n7320 & n12709;
  assign new_n13585 = n1094 & n6429;
  assign new_n13586 = ~new_n13584 & ~new_n13585;
  assign new_n13587 = new_n13584 & new_n13585;
  assign new_n13588 = ~new_n13586 & ~new_n13587;
  assign new_n13589 = ~new_n13583 & ~new_n13588;
  assign new_n13590 = new_n13583 & new_n13588;
  assign new_n13591 = ~new_n13589 & ~new_n13590;
  assign new_n13592 = ~new_n13582 & new_n13591;
  assign new_n13593 = ~new_n13581 & ~new_n13591;
  assign new_n13594 = ~new_n13580 & new_n13593;
  assign new_n13595 = ~new_n13592 & ~new_n13594;
  assign new_n13596 = ~new_n13578 & ~new_n13595;
  assign new_n13597 = new_n13578 & new_n13595;
  assign new_n13598 = ~new_n13596 & ~new_n13597;
  assign new_n13599 = ~new_n13564 & new_n13598;
  assign new_n13600 = new_n13564 & ~new_n13598;
  assign new_n13601 = ~new_n13599 & ~new_n13600;
  assign new_n13602 = ~new_n13552 & ~new_n13601;
  assign new_n13603 = new_n13552 & new_n13601;
  assign new_n13604 = ~new_n13602 & ~new_n13603;
  assign new_n13605 = ~new_n13559 & new_n13604;
  assign new_n13606 = new_n13559 & ~new_n13604;
  assign new_n13607 = ~new_n13605 & ~new_n13606;
  assign new_n13608 = ~new_n12319 & ~new_n13557;
  assign new_n13609 = ~new_n13558 & ~new_n13608;
  assign new_n13610 = ~new_n12325 & new_n12393;
  assign new_n13611 = ~new_n12324 & ~new_n13610;
  assign new_n13612 = ~new_n13609 & new_n13611;
  assign new_n13613 = new_n13609 & ~new_n13611;
  assign new_n13614 = n6441 & n11222;
  assign new_n13615 = ~new_n12375 & new_n12379;
  assign new_n13616 = ~new_n12376 & ~new_n13615;
  assign new_n13617 = n11153 & n12947;
  assign new_n13618 = n5314 & n11791;
  assign new_n13619 = ~new_n13617 & ~new_n13618;
  assign new_n13620 = new_n13617 & new_n13618;
  assign new_n13621 = ~new_n13619 & ~new_n13620;
  assign new_n13622 = ~new_n12360 & ~new_n12371;
  assign new_n13623 = ~new_n12361 & ~new_n13622;
  assign new_n13624 = new_n13621 & ~new_n13623;
  assign new_n13625 = ~new_n13621 & new_n13623;
  assign new_n13626 = ~new_n13624 & ~new_n13625;
  assign new_n13627 = n996 & n1478;
  assign new_n13628 = n5319 & n10990;
  assign new_n13629 = n5760 & n5767;
  assign new_n13630 = ~new_n13628 & ~new_n13629;
  assign new_n13631 = new_n13628 & new_n13629;
  assign new_n13632 = ~new_n13630 & ~new_n13631;
  assign new_n13633 = ~new_n13627 & ~new_n13632;
  assign new_n13634 = new_n12363 & ~new_n12366;
  assign new_n13635 = ~new_n12367 & ~new_n13634;
  assign new_n13636 = new_n13633 & new_n13635;
  assign new_n13637 = new_n13627 & new_n13632;
  assign new_n13638 = new_n13635 & ~new_n13637;
  assign new_n13639 = ~new_n13633 & ~new_n13638;
  assign new_n13640 = ~new_n13636 & ~new_n13639;
  assign new_n13641 = ~new_n13635 & new_n13637;
  assign new_n13642 = ~new_n13640 & ~new_n13641;
  assign new_n13643 = new_n13626 & new_n13642;
  assign new_n13644 = ~new_n13626 & ~new_n13642;
  assign new_n13645 = ~new_n13643 & ~new_n13644;
  assign new_n13646 = new_n13616 & ~new_n13645;
  assign new_n13647 = ~new_n13616 & new_n13645;
  assign new_n13648 = ~new_n13646 & ~new_n13647;
  assign new_n13649 = new_n13614 & new_n13648;
  assign new_n13650 = ~new_n13614 & ~new_n13648;
  assign new_n13651 = ~new_n13649 & ~new_n13650;
  assign new_n13652 = new_n12384 & new_n13651;
  assign new_n13653 = ~new_n12384 & ~new_n13651;
  assign new_n13654 = ~new_n13652 & ~new_n13653;
  assign new_n13655 = n447 & n12069;
  assign new_n13656 = ~new_n12346 & ~new_n12349;
  assign new_n13657 = ~new_n12345 & ~new_n13656;
  assign new_n13658 = n11967 & n12391;
  assign new_n13659 = n6254 & n7891;
  assign new_n13660 = ~new_n13658 & ~new_n13659;
  assign new_n13661 = new_n13658 & new_n13659;
  assign new_n13662 = ~new_n13660 & ~new_n13661;
  assign new_n13663 = n7160 & n12777;
  assign new_n13664 = n4828 & n7159;
  assign new_n13665 = n2515 & n12489;
  assign new_n13666 = ~new_n13664 & ~new_n13665;
  assign new_n13667 = new_n13664 & new_n13665;
  assign new_n13668 = ~new_n13666 & ~new_n13667;
  assign new_n13669 = new_n13663 & new_n13668;
  assign new_n13670 = ~new_n13663 & ~new_n13668;
  assign new_n13671 = ~new_n13669 & ~new_n13670;
  assign new_n13672 = new_n12334 & ~new_n12336;
  assign new_n13673 = ~new_n12337 & ~new_n13672;
  assign new_n13674 = ~new_n13671 & ~new_n13673;
  assign new_n13675 = new_n13671 & new_n13673;
  assign new_n13676 = ~new_n13674 & ~new_n13675;
  assign new_n13677 = new_n13662 & ~new_n13676;
  assign new_n13678 = ~new_n13662 & new_n13676;
  assign new_n13679 = ~new_n13677 & ~new_n13678;
  assign new_n13680 = ~new_n12331 & ~new_n12341;
  assign new_n13681 = ~new_n12332 & ~new_n13680;
  assign new_n13682 = new_n13679 & new_n13681;
  assign new_n13683 = ~new_n13679 & ~new_n13681;
  assign new_n13684 = ~new_n13682 & ~new_n13683;
  assign new_n13685 = ~new_n13657 & ~new_n13684;
  assign new_n13686 = new_n13657 & new_n13684;
  assign new_n13687 = ~new_n13685 & ~new_n13686;
  assign new_n13688 = new_n13655 & new_n13687;
  assign new_n13689 = ~new_n13655 & ~new_n13687;
  assign new_n13690 = ~new_n13688 & ~new_n13689;
  assign new_n13691 = new_n12353 & new_n13690;
  assign new_n13692 = ~new_n12353 & ~new_n13690;
  assign new_n13693 = ~new_n13691 & ~new_n13692;
  assign new_n13694 = new_n12355 & ~new_n12389;
  assign new_n13695 = ~new_n12388 & ~new_n13694;
  assign new_n13696 = new_n13693 & ~new_n13695;
  assign new_n13697 = ~new_n13693 & new_n13695;
  assign new_n13698 = ~new_n13696 & ~new_n13697;
  assign new_n13699 = new_n13654 & new_n13698;
  assign new_n13700 = ~new_n13654 & ~new_n13698;
  assign new_n13701 = ~new_n13699 & ~new_n13700;
  assign new_n13702 = ~new_n13613 & ~new_n13701;
  assign new_n13703 = ~new_n13612 & ~new_n13702;
  assign new_n13704 = ~new_n13607 & ~new_n13703;
  assign new_n13705 = new_n13607 & new_n13703;
  assign new_n13706 = ~new_n13704 & ~new_n13705;
  assign new_n13707 = ~new_n13625 & ~new_n13642;
  assign new_n13708 = ~new_n13620 & ~new_n13707;
  assign new_n13709 = ~new_n13624 & new_n13708;
  assign new_n13710 = new_n13620 & new_n13707;
  assign new_n13711 = ~new_n13709 & ~new_n13710;
  assign new_n13712 = n6441 & n11153;
  assign new_n13713 = n5314 & n12947;
  assign new_n13714 = n11222 & n11999;
  assign new_n13715 = ~new_n13713 & ~new_n13714;
  assign new_n13716 = new_n13713 & new_n13714;
  assign new_n13717 = ~new_n13715 & ~new_n13716;
  assign new_n13718 = ~new_n13712 & ~new_n13717;
  assign new_n13719 = new_n13712 & new_n13717;
  assign new_n13720 = ~new_n13718 & ~new_n13719;
  assign new_n13721 = new_n13639 & new_n13720;
  assign new_n13722 = ~new_n13639 & ~new_n13720;
  assign new_n13723 = ~new_n13721 & ~new_n13722;
  assign new_n13724 = n996 & n11791;
  assign new_n13725 = ~new_n13631 & ~new_n13724;
  assign new_n13726 = new_n13631 & new_n13724;
  assign new_n13727 = ~new_n13725 & ~new_n13726;
  assign new_n13728 = n5319 & n5760;
  assign new_n13729 = n9457 & n10990;
  assign new_n13730 = n1478 & n5767;
  assign new_n13731 = ~new_n13729 & ~new_n13730;
  assign new_n13732 = new_n13729 & new_n13730;
  assign new_n13733 = ~new_n13731 & ~new_n13732;
  assign new_n13734 = ~new_n13728 & ~new_n13733;
  assign new_n13735 = new_n13728 & new_n13733;
  assign new_n13736 = ~new_n13734 & ~new_n13735;
  assign new_n13737 = new_n13727 & ~new_n13736;
  assign new_n13738 = ~new_n13727 & new_n13736;
  assign new_n13739 = ~new_n13737 & ~new_n13738;
  assign new_n13740 = new_n13723 & new_n13739;
  assign new_n13741 = ~new_n13723 & ~new_n13739;
  assign new_n13742 = ~new_n13740 & ~new_n13741;
  assign new_n13743 = ~new_n13711 & new_n13742;
  assign new_n13744 = new_n13711 & ~new_n13742;
  assign new_n13745 = ~new_n13743 & ~new_n13744;
  assign new_n13746 = ~new_n13646 & ~new_n13745;
  assign new_n13747 = new_n13646 & new_n13745;
  assign new_n13748 = ~new_n13746 & ~new_n13747;
  assign new_n13749 = ~new_n13649 & ~new_n13652;
  assign new_n13750 = ~new_n13748 & new_n13749;
  assign new_n13751 = new_n13748 & ~new_n13749;
  assign new_n13752 = ~new_n13750 & ~new_n13751;
  assign new_n13753 = ~new_n13678 & ~new_n13681;
  assign new_n13754 = ~new_n13661 & ~new_n13753;
  assign new_n13755 = ~new_n13677 & new_n13754;
  assign new_n13756 = new_n13661 & new_n13753;
  assign new_n13757 = ~new_n13755 & ~new_n13756;
  assign new_n13758 = n7891 & n11967;
  assign new_n13759 = n1353 & n12069;
  assign new_n13760 = n447 & n12391;
  assign new_n13761 = ~new_n13759 & ~new_n13760;
  assign new_n13762 = new_n13759 & new_n13760;
  assign new_n13763 = ~new_n13761 & ~new_n13762;
  assign new_n13764 = new_n13758 & ~new_n13763;
  assign new_n13765 = ~new_n13758 & new_n13763;
  assign new_n13766 = ~new_n13764 & ~new_n13765;
  assign new_n13767 = ~new_n13669 & new_n13673;
  assign new_n13768 = ~new_n13670 & ~new_n13767;
  assign new_n13769 = new_n13766 & ~new_n13768;
  assign new_n13770 = n6254 & n7160;
  assign new_n13771 = new_n13667 & new_n13770;
  assign new_n13772 = ~new_n13667 & ~new_n13770;
  assign new_n13773 = ~new_n13771 & ~new_n13772;
  assign new_n13774 = n1199 & n12489;
  assign new_n13775 = n2515 & n7159;
  assign new_n13776 = n4828 & n12777;
  assign new_n13777 = ~new_n13775 & ~new_n13776;
  assign new_n13778 = new_n13775 & new_n13776;
  assign new_n13779 = ~new_n13777 & ~new_n13778;
  assign new_n13780 = new_n13774 & ~new_n13779;
  assign new_n13781 = ~new_n13774 & new_n13779;
  assign new_n13782 = ~new_n13780 & ~new_n13781;
  assign new_n13783 = new_n13773 & new_n13782;
  assign new_n13784 = ~new_n13773 & ~new_n13782;
  assign new_n13785 = ~new_n13783 & ~new_n13784;
  assign new_n13786 = new_n13769 & new_n13785;
  assign new_n13787 = ~new_n13766 & new_n13768;
  assign new_n13788 = new_n13785 & ~new_n13787;
  assign new_n13789 = ~new_n13769 & ~new_n13788;
  assign new_n13790 = ~new_n13786 & ~new_n13789;
  assign new_n13791 = ~new_n13785 & new_n13787;
  assign new_n13792 = ~new_n13790 & ~new_n13791;
  assign new_n13793 = ~new_n13757 & new_n13792;
  assign new_n13794 = new_n13757 & ~new_n13792;
  assign new_n13795 = ~new_n13793 & ~new_n13794;
  assign new_n13796 = ~new_n13685 & ~new_n13795;
  assign new_n13797 = new_n13685 & new_n13795;
  assign new_n13798 = ~new_n13796 & ~new_n13797;
  assign new_n13799 = ~new_n13688 & ~new_n13691;
  assign new_n13800 = ~new_n13798 & new_n13799;
  assign new_n13801 = new_n13798 & ~new_n13799;
  assign new_n13802 = ~new_n13800 & ~new_n13801;
  assign new_n13803 = new_n13752 & new_n13802;
  assign new_n13804 = ~new_n13752 & ~new_n13802;
  assign new_n13805 = ~new_n13803 & ~new_n13804;
  assign new_n13806 = new_n13654 & ~new_n13697;
  assign new_n13807 = ~new_n13696 & ~new_n13806;
  assign new_n13808 = ~new_n13805 & ~new_n13807;
  assign new_n13809 = new_n13805 & new_n13807;
  assign new_n13810 = ~new_n13808 & ~new_n13809;
  assign new_n13811 = new_n13706 & ~new_n13810;
  assign new_n13812 = ~new_n13706 & new_n13810;
  assign new_n13813 = ~new_n13811 & ~new_n13812;
  assign new_n13814 = ~new_n13521 & ~new_n13813;
  assign new_n13815 = new_n13521 & new_n13813;
  assign new_n13816 = ~new_n13814 & ~new_n13815;
  assign new_n13817 = ~new_n12289 & ~new_n13516;
  assign new_n13818 = ~new_n13517 & ~new_n13817;
  assign new_n13819 = ~new_n12397 & ~new_n12401;
  assign new_n13820 = ~new_n12398 & ~new_n13819;
  assign new_n13821 = new_n13818 & ~new_n13820;
  assign new_n13822 = ~new_n13818 & new_n13820;
  assign new_n13823 = ~new_n13612 & ~new_n13613;
  assign new_n13824 = new_n13701 & ~new_n13823;
  assign new_n13825 = ~new_n13701 & new_n13823;
  assign new_n13826 = ~new_n13824 & ~new_n13825;
  assign new_n13827 = ~new_n13822 & ~new_n13826;
  assign new_n13828 = ~new_n13821 & ~new_n13827;
  assign new_n13829 = ~new_n13816 & new_n13828;
  assign new_n13830 = new_n13816 & ~new_n13828;
  assign n5132 = ~new_n13829 & ~new_n13830;
  assign new_n13832 = ~new_n13119 & ~new_n13121;
  assign n5191 = ~new_n13122 & ~new_n13832;
  assign new_n13834 = ~new_n4166 & new_n4328;
  assign new_n13835 = ~new_n4165 & ~new_n13834;
  assign new_n13836 = ~new_n4322 & new_n4325;
  assign new_n13837 = ~new_n4321 & ~new_n13836;
  assign new_n13838 = new_n3664 & ~new_n3667;
  assign new_n13839 = ~new_n3668 & ~new_n13838;
  assign new_n13840 = ~new_n3674 & ~new_n3691;
  assign new_n13841 = ~new_n3673 & ~new_n13840;
  assign new_n13842 = ~new_n13839 & new_n13841;
  assign new_n13843 = new_n13839 & ~new_n13841;
  assign new_n13844 = ~new_n13842 & ~new_n13843;
  assign new_n13845 = n2577 & n11757;
  assign new_n13846 = n3172 & n9637;
  assign new_n13847 = new_n13845 & ~new_n13846;
  assign new_n13848 = ~new_n13845 & new_n13846;
  assign new_n13849 = ~new_n13847 & ~new_n13848;
  assign new_n13850 = n11821 & n11917;
  assign new_n13851 = n4921 & n9080;
  assign new_n13852 = new_n13850 & ~new_n13851;
  assign new_n13853 = ~new_n13850 & new_n13851;
  assign new_n13854 = ~new_n13852 & ~new_n13853;
  assign new_n13855 = ~new_n13849 & new_n13854;
  assign new_n13856 = new_n13849 & ~new_n13854;
  assign new_n13857 = ~new_n13855 & ~new_n13856;
  assign new_n13858 = ~new_n3680 & ~new_n3684;
  assign new_n13859 = ~new_n3683 & ~new_n13858;
  assign new_n13860 = n1333 & n1835;
  assign new_n13861 = n3842 & n5240;
  assign new_n13862 = ~new_n13860 & new_n13861;
  assign new_n13863 = new_n13860 & ~new_n13861;
  assign new_n13864 = ~new_n13862 & ~new_n13863;
  assign new_n13865 = new_n13859 & new_n13864;
  assign new_n13866 = ~new_n13859 & ~new_n13864;
  assign new_n13867 = ~new_n13865 & ~new_n13866;
  assign new_n13868 = new_n13857 & new_n13867;
  assign new_n13869 = ~new_n13857 & ~new_n13867;
  assign new_n13870 = ~new_n13868 & ~new_n13869;
  assign new_n13871 = ~new_n3678 & new_n3688;
  assign new_n13872 = ~new_n3677_1 & ~new_n13871;
  assign new_n13873 = ~new_n13870 & new_n13872;
  assign new_n13874 = new_n13870 & ~new_n13872;
  assign new_n13875 = ~new_n13873 & ~new_n13874;
  assign new_n13876 = ~new_n13844 & ~new_n13875;
  assign new_n13877 = new_n13844 & new_n13875;
  assign new_n13878 = ~new_n13876 & ~new_n13877;
  assign new_n13879 = n3719 & n10174;
  assign new_n13880 = n4190 & n6877;
  assign new_n13881 = new_n13879 & ~new_n13880;
  assign new_n13882 = ~new_n13879 & new_n13880;
  assign new_n13883 = ~new_n13881 & ~new_n13882;
  assign new_n13884 = ~new_n13878 & new_n13883;
  assign new_n13885 = new_n13878 & ~new_n13883;
  assign new_n13886 = ~new_n13884 & ~new_n13885;
  assign new_n13887 = ~new_n4171 & ~new_n4206;
  assign new_n13888 = ~new_n4172 & ~new_n13887;
  assign new_n13889 = n3602 & n12753;
  assign new_n13890 = new_n13888 & new_n13889;
  assign new_n13891 = ~new_n13888 & ~new_n13889;
  assign new_n13892 = ~new_n13890 & ~new_n13891;
  assign new_n13893 = new_n13886 & new_n13892;
  assign new_n13894 = ~new_n13886 & ~new_n13892;
  assign new_n13895 = ~new_n13893 & ~new_n13894;
  assign new_n13896 = ~new_n4307 & ~new_n4311;
  assign new_n13897 = ~new_n4268 & new_n4302;
  assign new_n13898 = ~new_n4269 & ~new_n13897;
  assign new_n13899 = ~new_n4176 & ~new_n4180;
  assign new_n13900 = ~new_n4179 & ~new_n13899;
  assign new_n13901 = n405 & n7646;
  assign new_n13902 = n4722 & n8433;
  assign new_n13903 = ~new_n13901 & new_n13902;
  assign new_n13904 = new_n13901 & ~new_n13902;
  assign new_n13905 = ~new_n13903 & ~new_n13904;
  assign new_n13906 = n1471 & n4086;
  assign new_n13907 = n1357 & n7236;
  assign new_n13908 = ~new_n13906 & ~new_n13907;
  assign new_n13909 = new_n13906 & new_n13907;
  assign new_n13910 = ~new_n13908 & ~new_n13909;
  assign new_n13911 = ~new_n13905 & new_n13910;
  assign new_n13912 = new_n13905 & ~new_n13910;
  assign new_n13913 = ~new_n13911 & ~new_n13912;
  assign new_n13914 = ~new_n13900 & new_n13913;
  assign new_n13915 = new_n13900 & ~new_n13913;
  assign new_n13916 = ~new_n13914 & ~new_n13915;
  assign new_n13917 = new_n13898 & ~new_n13916;
  assign new_n13918 = ~new_n13898 & new_n13916;
  assign new_n13919 = ~new_n13917 & ~new_n13918;
  assign new_n13920 = ~new_n4185 & new_n4203_1;
  assign new_n13921 = ~new_n4186 & ~new_n13920;
  assign new_n13922 = ~new_n4189_1 & ~new_n4200;
  assign new_n13923 = ~new_n4190_1 & ~new_n13922;
  assign new_n13924 = n4187 & n8595;
  assign new_n13925 = n4203 & n6126;
  assign new_n13926 = new_n13924 & ~new_n13925;
  assign new_n13927 = ~new_n13924 & new_n13925;
  assign new_n13928 = ~new_n13926 & ~new_n13927;
  assign new_n13929 = ~new_n4192 & ~new_n4196;
  assign new_n13930 = ~new_n4195 & ~new_n13929;
  assign new_n13931 = ~new_n13928 & new_n13930;
  assign new_n13932 = new_n13928 & ~new_n13930;
  assign new_n13933 = ~new_n13931 & ~new_n13932;
  assign new_n13934 = n9400 & n10391;
  assign new_n13935 = n2464 & n8065;
  assign new_n13936 = n10439 & n11311;
  assign new_n13937 = ~new_n13935 & ~new_n13936;
  assign new_n13938 = new_n13935 & new_n13936;
  assign new_n13939 = ~new_n13937 & ~new_n13938;
  assign new_n13940 = new_n13934 & new_n13939;
  assign new_n13941 = ~new_n13934 & ~new_n13939;
  assign new_n13942 = ~new_n13940 & ~new_n13941;
  assign new_n13943 = new_n13933 & new_n13942;
  assign new_n13944 = ~new_n13933 & ~new_n13942;
  assign new_n13945 = ~new_n13943 & ~new_n13944;
  assign new_n13946 = ~new_n13923 & new_n13945;
  assign new_n13947 = new_n13923 & ~new_n13945;
  assign new_n13948 = ~new_n13946 & ~new_n13947;
  assign new_n13949 = new_n13921 & ~new_n13948;
  assign new_n13950 = ~new_n13921 & new_n13948;
  assign new_n13951 = ~new_n13949 & ~new_n13950;
  assign new_n13952 = ~new_n13919 & new_n13951;
  assign new_n13953 = new_n13919 & ~new_n13951;
  assign new_n13954 = ~new_n13952 & ~new_n13953;
  assign new_n13955 = ~new_n13896 & new_n13954;
  assign new_n13956 = new_n13896 & ~new_n13954;
  assign new_n13957 = ~new_n13955 & ~new_n13956;
  assign new_n13958 = ~new_n13895 & new_n13957;
  assign new_n13959 = new_n13895 & ~new_n13957;
  assign new_n13960 = ~new_n13958 & ~new_n13959;
  assign new_n13961 = ~new_n4211 & ~new_n4213;
  assign new_n13962 = ~new_n4314 & ~new_n4317;
  assign new_n13963 = ~new_n4313 & ~new_n13962;
  assign new_n13964 = new_n13961 & new_n13963;
  assign new_n13965 = ~new_n13961 & ~new_n13963;
  assign new_n13966 = ~new_n13964 & ~new_n13965;
  assign new_n13967 = new_n13960 & ~new_n13966;
  assign new_n13968 = ~new_n13960 & new_n13966;
  assign new_n13969 = ~new_n13967 & ~new_n13968;
  assign new_n13970 = ~new_n13837 & ~new_n13969;
  assign new_n13971 = new_n13837 & new_n13969;
  assign new_n13972 = ~new_n13970 & ~new_n13971;
  assign new_n13973 = n4805 & n7546;
  assign new_n13974 = n4938 & n12925;
  assign new_n13975 = ~new_n13973 & new_n13974;
  assign new_n13976 = new_n13973 & ~new_n13974;
  assign new_n13977 = ~new_n13975 & ~new_n13976;
  assign new_n13978 = ~new_n4282 & new_n4299;
  assign new_n13979 = ~new_n4281 & ~new_n13978;
  assign new_n13980 = ~new_n13977 & new_n13979;
  assign new_n13981 = new_n13977 & ~new_n13979;
  assign new_n13982 = ~new_n13980 & ~new_n13981;
  assign new_n13983 = n137 & n4970;
  assign new_n13984 = n6294 & n7610;
  assign new_n13985 = ~new_n13983 & ~new_n13984;
  assign new_n13986 = new_n13983 & new_n13984;
  assign new_n13987 = ~new_n13985 & ~new_n13986;
  assign new_n13988 = n4826 & n6797;
  assign new_n13989 = n3146 & n7733;
  assign new_n13990 = new_n13988 & ~new_n13989;
  assign new_n13991 = ~new_n13988 & new_n13989;
  assign new_n13992 = ~new_n13990 & ~new_n13991;
  assign new_n13993 = ~new_n13987 & ~new_n13992;
  assign new_n13994 = new_n13987 & new_n13992;
  assign new_n13995 = ~new_n13993 & ~new_n13994;
  assign new_n13996 = ~new_n13982 & new_n13995;
  assign new_n13997 = new_n13982 & ~new_n13995;
  assign new_n13998 = ~new_n13996 & ~new_n13997;
  assign new_n13999 = ~new_n4218 & ~new_n4255;
  assign new_n14000 = ~new_n4219 & ~new_n13999;
  assign new_n14001 = new_n4272 & ~new_n4275;
  assign new_n14002 = ~new_n4276 & ~new_n14001;
  assign new_n14003 = new_n4288 & ~new_n4291;
  assign new_n14004 = ~new_n4292 & ~new_n14003;
  assign new_n14005 = ~new_n14002 & new_n14004;
  assign new_n14006 = new_n14002 & ~new_n14004;
  assign new_n14007 = ~new_n14005 & ~new_n14006;
  assign new_n14008 = ~new_n4286 & new_n4296;
  assign new_n14009 = ~new_n4285 & ~new_n14008;
  assign new_n14010 = n6359 & n8384;
  assign new_n14011 = n3992 & n11296;
  assign new_n14012 = n6358 & n6611;
  assign new_n14013 = n217 & n5198;
  assign new_n14014 = ~new_n14012 & new_n14013;
  assign new_n14015 = new_n14012 & ~new_n14013;
  assign new_n14016 = ~new_n14014 & ~new_n14015;
  assign new_n14017 = new_n14011 & new_n14016;
  assign new_n14018 = ~new_n14011 & ~new_n14016;
  assign new_n14019 = ~new_n14017 & ~new_n14018;
  assign new_n14020 = new_n14010 & new_n14019;
  assign new_n14021 = ~new_n14010 & ~new_n14019;
  assign new_n14022 = ~new_n14020 & ~new_n14021;
  assign new_n14023 = new_n14009 & ~new_n14022;
  assign new_n14024 = ~new_n14009 & new_n14022;
  assign new_n14025 = ~new_n14023 & ~new_n14024;
  assign new_n14026 = ~new_n14007 & ~new_n14025;
  assign new_n14027 = new_n14007 & new_n14025;
  assign new_n14028 = ~new_n14026 & ~new_n14027;
  assign new_n14029 = new_n14000 & new_n14028;
  assign new_n14030 = ~new_n14000 & ~new_n14028;
  assign new_n14031 = ~new_n14029 & ~new_n14030;
  assign new_n14032 = new_n13998 & new_n14031;
  assign new_n14033 = ~new_n13998 & ~new_n14031;
  assign new_n14034 = ~new_n14032 & ~new_n14033;
  assign new_n14035 = new_n4223 & ~new_n4226_1;
  assign new_n14036 = ~new_n4227 & ~new_n14035;
  assign new_n14037 = new_n4252 & ~new_n14036;
  assign new_n14038 = ~new_n4252 & new_n14036;
  assign new_n14039 = ~new_n14037 & ~new_n14038;
  assign new_n14040 = n503 & n5283;
  assign new_n14041 = n10965 & n11478;
  assign new_n14042 = ~new_n14040 & new_n14041;
  assign new_n14043 = new_n14040 & ~new_n14041;
  assign new_n14044 = ~new_n14042 & ~new_n14043;
  assign new_n14045 = ~new_n4237 & ~new_n4241;
  assign new_n14046 = ~new_n4240 & ~new_n14045;
  assign new_n14047 = ~new_n4235 & new_n4245;
  assign new_n14048 = ~new_n4234 & ~new_n14047;
  assign new_n14049 = new_n14046 & new_n14048;
  assign new_n14050 = ~new_n14046 & ~new_n14048;
  assign new_n14051 = ~new_n14049 & ~new_n14050;
  assign new_n14052 = new_n14044 & ~new_n14051;
  assign new_n14053 = ~new_n14044 & new_n14051;
  assign new_n14054 = ~new_n14052 & ~new_n14053;
  assign new_n14055 = ~new_n14039 & ~new_n14054;
  assign new_n14056 = new_n14039 & new_n14054;
  assign new_n14057 = ~new_n14055 & ~new_n14056;
  assign new_n14058 = ~new_n3660 & new_n3694;
  assign new_n14059 = ~new_n3659 & ~new_n14058;
  assign new_n14060 = n6826 & n9956;
  assign new_n14061 = n7862 & n11536;
  assign new_n14062 = ~new_n14060 & new_n14061;
  assign new_n14063 = new_n14060 & ~new_n14061;
  assign new_n14064 = ~new_n14062 & ~new_n14063;
  assign new_n14065 = ~new_n14059 & ~new_n14064;
  assign new_n14066 = new_n14059 & new_n14064;
  assign new_n14067 = ~new_n14065 & ~new_n14066;
  assign new_n14068 = ~new_n14057 & new_n14067;
  assign new_n14069 = new_n14057 & ~new_n14067;
  assign new_n14070 = ~new_n14068 & ~new_n14069;
  assign new_n14071 = ~new_n14034 & new_n14070;
  assign new_n14072 = new_n14034 & ~new_n14070;
  assign new_n14073 = ~new_n14071 & ~new_n14072;
  assign new_n14074 = ~new_n4260 & ~new_n4264;
  assign new_n14075 = ~new_n3699 & ~new_n3725;
  assign new_n14076 = new_n14074 & new_n14075;
  assign new_n14077 = ~new_n14074 & ~new_n14075;
  assign new_n14078 = ~new_n14076 & ~new_n14077;
  assign new_n14079 = ~new_n14073 & new_n14078;
  assign new_n14080 = new_n14073 & ~new_n14078;
  assign new_n14081 = ~new_n14079 & ~new_n14080;
  assign new_n14082 = ~new_n13972 & new_n14081;
  assign new_n14083 = new_n13972 & ~new_n14081;
  assign new_n14084 = ~new_n14082 & ~new_n14083;
  assign new_n14085 = new_n13835 & ~new_n14084;
  assign new_n14086 = ~new_n13835 & new_n14084;
  assign n5257 = ~new_n14085 & ~new_n14086;
  assign new_n14088 = ~new_n13117 & ~new_n13118;
  assign new_n14089 = new_n13132 & ~new_n14088;
  assign new_n14090 = ~new_n13132 & new_n14088;
  assign n5411 = ~new_n14089 & ~new_n14090;
  assign new_n14092 = ~new_n4006 & ~new_n4007;
  assign new_n14093 = ~new_n4020 & ~new_n14092;
  assign new_n14094 = new_n4020 & new_n14092;
  assign n5435 = ~new_n14093 & ~new_n14094;
  assign new_n14096 = ~new_n7043 & ~new_n7052;
  assign n5641 = ~new_n7053 & ~new_n14096;
  assign new_n14098 = ~new_n10010 & ~new_n10011;
  assign new_n14099 = new_n10023 & ~new_n14098;
  assign new_n14100 = ~new_n10023 & new_n14098;
  assign n5670 = ~new_n14099 & ~new_n14100;
  assign new_n14102 = ~new_n5639 & ~new_n5640;
  assign new_n14103 = new_n5674 & new_n14102;
  assign new_n14104 = ~new_n5674 & ~new_n14102;
  assign n5693 = new_n14103 | new_n14104;
  assign new_n14106 = ~new_n1495 & ~new_n1496;
  assign new_n14107 = new_n1509 & ~new_n14106;
  assign new_n14108 = ~new_n1509 & new_n14106;
  assign n5934 = ~new_n14107 & ~new_n14108;
  assign new_n14110 = ~new_n13109 & ~new_n13110;
  assign new_n14111 = new_n13134 & ~new_n14110;
  assign new_n14112 = ~new_n13134 & new_n14110;
  assign n6089 = ~new_n14111 & ~new_n14112;
  assign new_n14114 = ~new_n9109 & ~new_n9112;
  assign new_n14115 = ~new_n9099 & ~new_n9102;
  assign new_n14116 = ~new_n9082 & ~new_n14115;
  assign new_n14117 = ~new_n9098 & new_n14116;
  assign new_n14118 = new_n9082 & new_n14115;
  assign new_n14119 = ~new_n14117 & ~new_n14118;
  assign new_n14120 = n4189 & n9195;
  assign new_n14121 = n3865 & n6687;
  assign new_n14122 = n2253 & n2564;
  assign new_n14123 = ~new_n14121 & ~new_n14122;
  assign new_n14124 = new_n14121 & new_n14122;
  assign new_n14125 = ~new_n14123 & ~new_n14124;
  assign new_n14126 = new_n14120 & ~new_n14125;
  assign new_n14127 = ~new_n14120 & new_n14125;
  assign new_n14128 = ~new_n14126 & ~new_n14127;
  assign new_n14129 = ~new_n9091 & new_n9094;
  assign new_n14130 = ~new_n9090 & ~new_n14129;
  assign new_n14131 = ~new_n14128 & ~new_n14130;
  assign new_n14132 = new_n14128 & new_n14130;
  assign new_n14133 = ~new_n14131 & ~new_n14132;
  assign new_n14134 = n4634 & n6770;
  assign new_n14135 = new_n9088 & new_n14134;
  assign new_n14136 = ~new_n9088 & ~new_n14134;
  assign new_n14137 = ~new_n14135 & ~new_n14136;
  assign new_n14138 = n2879 & n3627;
  assign new_n14139 = n4516 & n7265;
  assign new_n14140 = ~new_n6683 & ~new_n14139;
  assign new_n14141 = new_n6683 & new_n14139;
  assign new_n14142 = ~new_n14140 & ~new_n14141;
  assign new_n14143 = ~new_n14138 & ~new_n14142;
  assign new_n14144 = new_n14138 & new_n14142;
  assign new_n14145 = ~new_n14143 & ~new_n14144;
  assign new_n14146 = new_n14137 & ~new_n14145;
  assign new_n14147 = ~new_n14137 & new_n14145;
  assign new_n14148 = ~new_n14146 & ~new_n14147;
  assign new_n14149 = new_n14133 & new_n14148;
  assign new_n14150 = ~new_n14133 & ~new_n14148;
  assign new_n14151 = ~new_n14149 & ~new_n14150;
  assign new_n14152 = ~new_n14119 & new_n14151;
  assign new_n14153 = new_n14119 & ~new_n14151;
  assign new_n14154 = ~new_n14152 & ~new_n14153;
  assign new_n14155 = new_n9106 & new_n14154;
  assign new_n14156 = ~new_n9106 & ~new_n14154;
  assign new_n14157 = ~new_n14155 & ~new_n14156;
  assign new_n14158 = ~new_n14114 & new_n14157;
  assign new_n14159 = new_n14114 & ~new_n14157;
  assign new_n14160 = ~new_n14158 & ~new_n14159;
  assign new_n14161 = ~new_n9155 & ~new_n9158;
  assign new_n14162 = ~new_n9145 & ~new_n9148;
  assign new_n14163 = new_n9128 & new_n14162;
  assign new_n14164 = ~new_n9128 & ~new_n14162;
  assign new_n14165 = ~new_n9144 & new_n14164;
  assign new_n14166 = ~new_n14163 & ~new_n14165;
  assign new_n14167 = ~new_n9137_1 & ~new_n9140;
  assign new_n14168 = ~new_n9136 & ~new_n14167;
  assign new_n14169 = n6986 & n12145;
  assign new_n14170 = n8336 & n10217;
  assign new_n14171 = n10928 & n12221;
  assign new_n14172 = ~new_n14170 & ~new_n14171;
  assign new_n14173 = new_n14170 & new_n14171;
  assign new_n14174 = ~new_n14172 & ~new_n14173;
  assign new_n14175 = new_n14169 & ~new_n14174;
  assign new_n14176 = ~new_n14169 & new_n14174;
  assign new_n14177 = ~new_n14175 & ~new_n14176;
  assign new_n14178 = ~new_n14168 & ~new_n14177;
  assign new_n14179 = new_n14168 & new_n14177;
  assign new_n14180 = ~new_n14178 & ~new_n14179;
  assign new_n14181 = n2226 & n2522;
  assign new_n14182 = new_n9134 & new_n14181;
  assign new_n14183 = ~new_n9134 & ~new_n14181;
  assign new_n14184 = ~new_n14182 & ~new_n14183;
  assign new_n14185 = n2024 & n10678;
  assign new_n14186 = n1094 & n9189;
  assign new_n14187 = n7320 & n7946;
  assign new_n14188 = ~new_n14186 & ~new_n14187;
  assign new_n14189 = new_n14186 & new_n14187;
  assign new_n14190 = ~new_n14188 & ~new_n14189;
  assign new_n14191 = ~new_n14185 & ~new_n14190;
  assign new_n14192 = new_n14185 & new_n14190;
  assign new_n14193 = ~new_n14191 & ~new_n14192;
  assign new_n14194 = new_n14184 & ~new_n14193;
  assign new_n14195 = ~new_n14184 & new_n14193;
  assign new_n14196 = ~new_n14194 & ~new_n14195;
  assign new_n14197 = new_n14180 & new_n14196;
  assign new_n14198 = ~new_n14180 & ~new_n14196;
  assign new_n14199 = ~new_n14197 & ~new_n14198;
  assign new_n14200 = new_n14166 & new_n14199;
  assign new_n14201 = ~new_n14166 & ~new_n14199;
  assign new_n14202 = ~new_n14200 & ~new_n14201;
  assign new_n14203 = new_n9152 & ~new_n14202;
  assign new_n14204 = ~new_n9152 & new_n14202;
  assign new_n14205 = ~new_n14203 & ~new_n14204;
  assign new_n14206 = ~new_n14161 & new_n14205;
  assign new_n14207 = new_n14161 & ~new_n14205;
  assign new_n14208 = ~new_n14206 & ~new_n14207;
  assign new_n14209 = ~new_n9186 & ~new_n9190;
  assign new_n14210 = ~new_n9187 & ~new_n14209;
  assign new_n14211 = ~new_n9170 & ~new_n14210;
  assign new_n14212 = new_n9170 & new_n14210;
  assign new_n14213 = ~new_n14211 & ~new_n14212;
  assign new_n14214 = n5798 & n12391;
  assign new_n14215 = n6016 & n7891;
  assign new_n14216 = n2347 & n12069;
  assign new_n14217 = ~new_n14215 & ~new_n14216;
  assign new_n14218 = new_n14215 & new_n14216;
  assign new_n14219 = ~new_n14217 & ~new_n14218;
  assign new_n14220 = ~new_n14214 & ~new_n14219;
  assign new_n14221 = new_n14214 & new_n14219;
  assign new_n14222 = ~new_n14220 & ~new_n14221;
  assign new_n14223 = ~new_n9176 & new_n9182;
  assign new_n14224 = ~new_n9175 & ~new_n14223;
  assign new_n14225 = new_n14222 & ~new_n14224;
  assign new_n14226 = ~new_n14222 & new_n14224;
  assign new_n14227 = ~new_n14225 & ~new_n14226;
  assign new_n14228 = n521 & n7160;
  assign new_n14229 = new_n9181 & new_n14228;
  assign new_n14230 = ~new_n9181 & ~new_n14228;
  assign new_n14231 = ~new_n14229 & ~new_n14230;
  assign new_n14232 = n1199 & n2558;
  assign new_n14233 = n2498 & n2515;
  assign new_n14234 = n4828 & n5579;
  assign new_n14235 = ~new_n14233 & ~new_n14234;
  assign new_n14236 = new_n14233 & new_n14234;
  assign new_n14237 = ~new_n14235 & ~new_n14236;
  assign new_n14238 = new_n14232 & ~new_n14237;
  assign new_n14239 = ~new_n14232 & new_n14237;
  assign new_n14240 = ~new_n14238 & ~new_n14239;
  assign new_n14241 = new_n14231 & new_n14240;
  assign new_n14242 = ~new_n14231 & ~new_n14240;
  assign new_n14243 = ~new_n14241 & ~new_n14242;
  assign new_n14244 = new_n14227 & ~new_n14243;
  assign new_n14245 = ~new_n14227 & new_n14243;
  assign new_n14246 = ~new_n14244 & ~new_n14245;
  assign new_n14247 = ~new_n14213 & new_n14246;
  assign new_n14248 = ~new_n14212 & ~new_n14246;
  assign new_n14249 = ~new_n14211 & new_n14248;
  assign new_n14250 = ~new_n14247 & ~new_n14249;
  assign new_n14251 = ~new_n9194 & new_n14250;
  assign new_n14252 = new_n9194 & ~new_n14250;
  assign new_n14253 = ~new_n14251 & ~new_n14252;
  assign new_n14254 = ~new_n9197 & ~new_n9200;
  assign new_n14255 = ~new_n14253 & new_n14254;
  assign new_n14256 = new_n14253 & ~new_n14254;
  assign new_n14257 = ~new_n14255 & ~new_n14256;
  assign new_n14258 = ~new_n9236 & ~new_n9239;
  assign new_n14259 = ~new_n9226 & ~new_n9229;
  assign new_n14260 = ~new_n9209 & ~new_n14259;
  assign new_n14261 = ~new_n9225 & new_n14260;
  assign new_n14262 = new_n9209 & new_n14259;
  assign new_n14263 = ~new_n14261 & ~new_n14262;
  assign new_n14264 = n5153 & n11153;
  assign new_n14265 = n5314 & n7270;
  assign new_n14266 = n2507 & n11222;
  assign new_n14267 = ~new_n14265 & ~new_n14266;
  assign new_n14268 = new_n14265 & new_n14266;
  assign new_n14269 = ~new_n14267 & ~new_n14268;
  assign new_n14270 = ~new_n14264 & ~new_n14269;
  assign new_n14271 = new_n14264 & new_n14269;
  assign new_n14272 = ~new_n14270 & ~new_n14271;
  assign new_n14273 = ~new_n9218 & new_n9221;
  assign new_n14274 = ~new_n9217 & ~new_n14273;
  assign new_n14275 = new_n14272 & ~new_n14274;
  assign new_n14276 = ~new_n14272 & new_n14274;
  assign new_n14277 = ~new_n14275 & ~new_n14276;
  assign new_n14278 = n806 & n996;
  assign new_n14279 = new_n9215 & new_n14278;
  assign new_n14280 = ~new_n9215 & ~new_n14278;
  assign new_n14281 = ~new_n14279 & ~new_n14280;
  assign new_n14282 = n5319 & n9111;
  assign new_n14283 = n9457 & n9763;
  assign new_n14284 = n3342 & n5767;
  assign new_n14285 = ~new_n14283 & ~new_n14284;
  assign new_n14286 = new_n14283 & new_n14284;
  assign new_n14287 = ~new_n14285 & ~new_n14286;
  assign new_n14288 = ~new_n14282 & ~new_n14287;
  assign new_n14289 = new_n14282 & new_n14287;
  assign new_n14290 = ~new_n14288 & ~new_n14289;
  assign new_n14291 = new_n14281 & ~new_n14290;
  assign new_n14292 = ~new_n14281 & new_n14290;
  assign new_n14293 = ~new_n14291 & ~new_n14292;
  assign new_n14294 = ~new_n14277 & ~new_n14293;
  assign new_n14295 = new_n14277 & new_n14293;
  assign new_n14296 = ~new_n14294 & ~new_n14295;
  assign new_n14297 = ~new_n14263 & new_n14296;
  assign new_n14298 = new_n14263 & ~new_n14296;
  assign new_n14299 = ~new_n14297 & ~new_n14298;
  assign new_n14300 = ~new_n9233 & ~new_n14299;
  assign new_n14301 = new_n9233 & new_n14299;
  assign new_n14302 = ~new_n14300 & ~new_n14301;
  assign new_n14303 = ~new_n14258 & new_n14302;
  assign new_n14304 = new_n14258 & ~new_n14302;
  assign new_n14305 = ~new_n14303 & ~new_n14304;
  assign new_n14306 = ~new_n14257 & ~new_n14305;
  assign new_n14307 = new_n14257 & new_n14305;
  assign new_n14308 = ~new_n14306 & ~new_n14307;
  assign new_n14309 = ~new_n9243 & ~new_n9246;
  assign new_n14310 = ~new_n9242 & ~new_n14309;
  assign new_n14311 = ~new_n14308 & new_n14310;
  assign new_n14312 = new_n14308 & ~new_n14310;
  assign new_n14313 = ~new_n14311 & ~new_n14312;
  assign new_n14314 = ~new_n14208 & ~new_n14313;
  assign new_n14315 = new_n14208 & new_n14313;
  assign new_n14316 = ~new_n14314 & ~new_n14315;
  assign new_n14317 = ~new_n9162 & new_n9249;
  assign new_n14318 = ~new_n9161 & ~new_n14317;
  assign new_n14319 = ~new_n14316 & ~new_n14318;
  assign new_n14320 = new_n14316 & new_n14318;
  assign new_n14321 = ~new_n14319 & ~new_n14320;
  assign new_n14322 = new_n14160 & new_n14321;
  assign new_n14323 = ~new_n14160 & ~new_n14321;
  assign new_n14324 = ~new_n9118 & new_n9252;
  assign new_n14325 = ~new_n9117 & ~new_n14324;
  assign new_n14326 = ~new_n14323 & ~new_n14325;
  assign new_n14327 = ~new_n14322 & ~new_n14326;
  assign new_n14328 = ~new_n14155 & ~new_n14158;
  assign new_n14329 = ~new_n14211 & ~new_n14248;
  assign new_n14330 = ~new_n14226 & ~new_n14243;
  assign new_n14331 = ~new_n14225 & ~new_n14330;
  assign new_n14332 = ~new_n14230 & ~new_n14240;
  assign new_n14333 = ~new_n14229 & ~new_n14332;
  assign new_n14334 = new_n14232 & ~new_n14235;
  assign new_n14335 = ~new_n14236 & ~new_n14334;
  assign new_n14336 = n5798 & n7891;
  assign new_n14337 = n2347 & n12391;
  assign new_n14338 = ~new_n14336 & new_n14337;
  assign new_n14339 = new_n14336 & ~new_n14337;
  assign new_n14340 = ~new_n14338 & ~new_n14339;
  assign new_n14341 = new_n14335 & ~new_n14340;
  assign new_n14342 = ~new_n14335 & new_n14340;
  assign new_n14343 = ~new_n14341 & ~new_n14342;
  assign new_n14344 = ~new_n14214 & ~new_n14218;
  assign new_n14345 = ~new_n14217 & ~new_n14344;
  assign new_n14346 = ~new_n14343 & new_n14345;
  assign new_n14347 = new_n14343 & ~new_n14345;
  assign new_n14348 = ~new_n14346 & ~new_n14347;
  assign new_n14349 = ~new_n14333 & new_n14348;
  assign new_n14350 = new_n14333 & ~new_n14348;
  assign new_n14351 = ~new_n14349 & ~new_n14350;
  assign new_n14352 = new_n14331 & ~new_n14351;
  assign new_n14353 = ~new_n14331 & new_n14351;
  assign new_n14354 = ~new_n14352 & ~new_n14353;
  assign new_n14355 = ~new_n14117 & ~new_n14151;
  assign new_n14356 = ~new_n14118 & ~new_n14355;
  assign new_n14357 = n2512 & n6687;
  assign new_n14358 = n2087 & n7265;
  assign new_n14359 = ~new_n14357 & new_n14358;
  assign new_n14360 = new_n14357 & ~new_n14358;
  assign new_n14361 = ~new_n14359 & ~new_n14360;
  assign new_n14362 = new_n14356 & new_n14361;
  assign new_n14363 = ~new_n14356 & ~new_n14361;
  assign new_n14364 = ~new_n14362 & ~new_n14363;
  assign new_n14365 = ~new_n14354 & new_n14364;
  assign new_n14366 = new_n14354 & ~new_n14364;
  assign new_n14367 = ~new_n14365 & ~new_n14366;
  assign new_n14368 = ~new_n14329 & new_n14367;
  assign new_n14369 = new_n14329 & ~new_n14367;
  assign new_n14370 = ~new_n14368 & ~new_n14369;
  assign new_n14371 = new_n14328 & new_n14370;
  assign new_n14372 = ~new_n14328 & ~new_n14370;
  assign new_n14373 = ~new_n14371 & ~new_n14372;
  assign new_n14374 = new_n14327 & new_n14373;
  assign new_n14375 = ~new_n14327 & ~new_n14373;
  assign new_n14376 = ~new_n14374 & ~new_n14375;
  assign new_n14377 = ~new_n14314 & new_n14318;
  assign new_n14378 = ~new_n14315 & ~new_n14377;
  assign new_n14379 = n6016 & n7160;
  assign new_n14380 = n521 & n4828;
  assign new_n14381 = ~new_n14379 & ~new_n14380;
  assign new_n14382 = new_n14379 & new_n14380;
  assign new_n14383 = ~new_n14381 & ~new_n14382;
  assign new_n14384 = n2515 & n5579;
  assign new_n14385 = n1199 & n2498;
  assign new_n14386 = new_n14384 & ~new_n14385;
  assign new_n14387 = ~new_n14384 & new_n14385;
  assign new_n14388 = ~new_n14386 & ~new_n14387;
  assign new_n14389 = ~new_n14383 & ~new_n14388;
  assign new_n14390 = new_n14383 & new_n14388;
  assign new_n14391 = ~new_n14389 & ~new_n14390;
  assign new_n14392 = ~new_n14378 & new_n14391;
  assign new_n14393 = new_n14378 & ~new_n14391;
  assign new_n14394 = ~new_n14392 & ~new_n14393;
  assign new_n14395 = ~new_n14282 & ~new_n14286;
  assign new_n14396 = ~new_n14285 & ~new_n14395;
  assign new_n14397 = n1576 & n12069;
  assign new_n14398 = n5153 & n5314;
  assign new_n14399 = new_n14397 & ~new_n14398;
  assign new_n14400 = ~new_n14397 & new_n14398;
  assign new_n14401 = ~new_n14399 & ~new_n14400;
  assign new_n14402 = ~new_n14396 & ~new_n14401;
  assign new_n14403 = new_n14396 & new_n14401;
  assign new_n14404 = ~new_n14402 & ~new_n14403;
  assign new_n14405 = ~new_n14275 & new_n14293;
  assign new_n14406 = ~new_n14276 & ~new_n14405;
  assign new_n14407 = ~new_n14279 & ~new_n14290;
  assign new_n14408 = ~new_n14280 & ~new_n14407;
  assign new_n14409 = n2507 & n11153;
  assign new_n14410 = n996 & n7270;
  assign new_n14411 = n806 & n5767;
  assign new_n14412 = ~new_n14410 & new_n14411;
  assign new_n14413 = new_n14410 & ~new_n14411;
  assign new_n14414 = ~new_n14412 & ~new_n14413;
  assign new_n14415 = new_n14409 & new_n14414;
  assign new_n14416 = ~new_n14409 & ~new_n14414;
  assign new_n14417 = ~new_n14415 & ~new_n14416;
  assign new_n14418 = ~new_n14264 & ~new_n14268;
  assign new_n14419 = ~new_n14267 & ~new_n14418;
  assign new_n14420 = ~new_n14417 & new_n14419;
  assign new_n14421 = new_n14417 & ~new_n14419;
  assign new_n14422 = ~new_n14420 & ~new_n14421;
  assign new_n14423 = new_n14408 & new_n14422;
  assign new_n14424 = ~new_n14408 & ~new_n14422;
  assign new_n14425 = ~new_n14423 & ~new_n14424;
  assign new_n14426 = new_n14406 & ~new_n14425;
  assign new_n14427 = ~new_n14406 & new_n14425;
  assign new_n14428 = ~new_n14426 & ~new_n14427;
  assign new_n14429 = ~new_n14404 & ~new_n14428;
  assign new_n14430 = new_n14404 & new_n14428;
  assign new_n14431 = ~new_n14429 & ~new_n14430;
  assign new_n14432 = ~new_n14306 & ~new_n14310;
  assign new_n14433 = ~new_n14307 & ~new_n14432;
  assign new_n14434 = ~new_n14261 & ~new_n14296;
  assign new_n14435 = ~new_n14262 & ~new_n14434;
  assign new_n14436 = ~new_n14178 & new_n14196;
  assign new_n14437 = ~new_n14179 & ~new_n14436;
  assign new_n14438 = ~new_n14185 & ~new_n14189;
  assign new_n14439 = ~new_n14188 & ~new_n14438;
  assign new_n14440 = n1094 & n2522;
  assign new_n14441 = n9189 & n10678;
  assign new_n14442 = ~new_n14440 & new_n14441;
  assign new_n14443 = new_n14440 & ~new_n14441;
  assign new_n14444 = ~new_n14442 & ~new_n14443;
  assign new_n14445 = n10217 & n10928;
  assign new_n14446 = n6986 & n12221;
  assign new_n14447 = new_n14445 & new_n14446;
  assign new_n14448 = ~new_n14445 & ~new_n14446;
  assign new_n14449 = ~new_n14447 & ~new_n14448;
  assign new_n14450 = new_n14444 & ~new_n14449;
  assign new_n14451 = ~new_n14444 & new_n14449;
  assign new_n14452 = ~new_n14450 & ~new_n14451;
  assign new_n14453 = ~new_n14439 & new_n14452;
  assign new_n14454 = new_n14439 & ~new_n14452;
  assign new_n14455 = ~new_n14453 & ~new_n14454;
  assign new_n14456 = new_n14437 & new_n14455;
  assign new_n14457 = ~new_n14437 & ~new_n14455;
  assign new_n14458 = ~new_n14456 & ~new_n14457;
  assign new_n14459 = ~new_n14183 & new_n14193;
  assign new_n14460 = ~new_n14182 & ~new_n14459;
  assign new_n14461 = n2226 & n12145;
  assign new_n14462 = new_n14169 & ~new_n14172;
  assign new_n14463 = ~new_n14173 & ~new_n14462;
  assign new_n14464 = ~new_n14461 & new_n14463;
  assign new_n14465 = new_n14461 & ~new_n14463;
  assign new_n14466 = ~new_n14464 & ~new_n14465;
  assign new_n14467 = ~new_n14460 & new_n14466;
  assign new_n14468 = new_n14460 & ~new_n14466;
  assign new_n14469 = ~new_n14467 & ~new_n14468;
  assign new_n14470 = n3342 & n5319;
  assign new_n14471 = n9111 & n9457;
  assign new_n14472 = ~new_n14470 & ~new_n14471;
  assign new_n14473 = new_n14470 & new_n14471;
  assign new_n14474 = ~new_n14472 & ~new_n14473;
  assign new_n14475 = n6431 & n11222;
  assign new_n14476 = n4817 & n9763;
  assign new_n14477 = new_n14475 & ~new_n14476;
  assign new_n14478 = ~new_n14475 & new_n14476;
  assign new_n14479 = ~new_n14477 & ~new_n14478;
  assign new_n14480 = ~new_n14474 & ~new_n14479;
  assign new_n14481 = new_n14474 & new_n14479;
  assign new_n14482 = ~new_n14480 & ~new_n14481;
  assign new_n14483 = ~new_n14469 & new_n14482;
  assign new_n14484 = new_n14469 & ~new_n14482;
  assign new_n14485 = ~new_n14483 & ~new_n14484;
  assign new_n14486 = new_n14458 & ~new_n14485;
  assign new_n14487 = ~new_n14458 & new_n14485;
  assign new_n14488 = ~new_n14486 & ~new_n14487;
  assign new_n14489 = ~new_n14435 & new_n14488;
  assign new_n14490 = new_n14435 & ~new_n14488;
  assign new_n14491 = ~new_n14489 & ~new_n14490;
  assign new_n14492 = ~new_n14301 & ~new_n14303;
  assign new_n14493 = ~new_n14165 & ~new_n14199;
  assign new_n14494 = ~new_n14163 & ~new_n14493;
  assign new_n14495 = n2024 & n7320;
  assign new_n14496 = n7523 & n7946;
  assign new_n14497 = n7823 & n8336;
  assign new_n14498 = ~new_n14496 & new_n14497;
  assign new_n14499 = new_n14496 & ~new_n14497;
  assign new_n14500 = ~new_n14498 & ~new_n14499;
  assign new_n14501 = new_n14495 & ~new_n14500;
  assign new_n14502 = ~new_n14495 & new_n14500;
  assign new_n14503 = ~new_n14501 & ~new_n14502;
  assign new_n14504 = new_n14494 & new_n14503;
  assign new_n14505 = ~new_n14494 & ~new_n14503;
  assign new_n14506 = ~new_n14504 & ~new_n14505;
  assign new_n14507 = ~new_n14135 & ~new_n14145;
  assign new_n14508 = ~new_n14136 & ~new_n14507;
  assign new_n14509 = ~new_n14138 & ~new_n14141;
  assign new_n14510 = ~new_n14140 & ~new_n14509;
  assign new_n14511 = n2564 & n3865;
  assign new_n14512 = n4634 & n9920;
  assign new_n14513 = ~new_n14511 & new_n14512;
  assign new_n14514 = new_n14511 & ~new_n14512;
  assign new_n14515 = ~new_n14513 & ~new_n14514;
  assign new_n14516 = new_n14510 & ~new_n14515;
  assign new_n14517 = ~new_n14510 & new_n14515;
  assign new_n14518 = ~new_n14516 & ~new_n14517;
  assign new_n14519 = n6770 & n9195;
  assign new_n14520 = n2253 & n4189;
  assign new_n14521 = new_n14519 & ~new_n14520;
  assign new_n14522 = ~new_n14519 & new_n14520;
  assign new_n14523 = ~new_n14521 & ~new_n14522;
  assign new_n14524 = n3627 & n10223;
  assign new_n14525 = n2879 & n4516;
  assign new_n14526 = new_n14524 & ~new_n14525;
  assign new_n14527 = ~new_n14524 & new_n14525;
  assign new_n14528 = ~new_n14526 & ~new_n14527;
  assign new_n14529 = ~new_n14523 & ~new_n14528;
  assign new_n14530 = new_n14523 & new_n14528;
  assign new_n14531 = ~new_n14529 & ~new_n14530;
  assign new_n14532 = ~new_n14518 & new_n14531;
  assign new_n14533 = new_n14518 & ~new_n14531;
  assign new_n14534 = ~new_n14532 & ~new_n14533;
  assign new_n14535 = ~new_n14508 & new_n14534;
  assign new_n14536 = new_n14508 & ~new_n14534;
  assign new_n14537 = ~new_n14535 & ~new_n14536;
  assign new_n14538 = ~new_n14120 & ~new_n14124;
  assign new_n14539 = ~new_n14123 & ~new_n14538;
  assign new_n14540 = ~new_n14132 & ~new_n14148;
  assign new_n14541 = ~new_n14131 & ~new_n14540;
  assign new_n14542 = new_n14539 & new_n14541;
  assign new_n14543 = ~new_n14539 & ~new_n14541;
  assign new_n14544 = ~new_n14542 & ~new_n14543;
  assign new_n14545 = ~new_n14537 & new_n14544;
  assign new_n14546 = new_n14537 & ~new_n14544;
  assign new_n14547 = ~new_n14545 & ~new_n14546;
  assign new_n14548 = new_n14506 & new_n14547;
  assign new_n14549 = ~new_n14506 & ~new_n14547;
  assign new_n14550 = ~new_n14548 & ~new_n14549;
  assign new_n14551 = new_n14492 & new_n14550;
  assign new_n14552 = ~new_n14492 & ~new_n14550;
  assign new_n14553 = ~new_n14551 & ~new_n14552;
  assign new_n14554 = new_n14491 & ~new_n14553;
  assign new_n14555 = ~new_n14491 & new_n14553;
  assign new_n14556 = ~new_n14554 & ~new_n14555;
  assign new_n14557 = ~new_n14433 & new_n14556;
  assign new_n14558 = new_n14433 & ~new_n14556;
  assign new_n14559 = ~new_n14557 & ~new_n14558;
  assign new_n14560 = new_n14431 & new_n14559;
  assign new_n14561 = ~new_n14431 & ~new_n14559;
  assign new_n14562 = ~new_n14560 & ~new_n14561;
  assign new_n14563 = ~new_n14252 & ~new_n14256;
  assign new_n14564 = ~new_n14203 & ~new_n14206;
  assign new_n14565 = n2558 & n6578;
  assign new_n14566 = new_n14564 & ~new_n14565;
  assign new_n14567 = ~new_n14564 & new_n14565;
  assign new_n14568 = ~new_n14566 & ~new_n14567;
  assign new_n14569 = ~new_n14563 & ~new_n14568;
  assign new_n14570 = new_n14563 & new_n14568;
  assign new_n14571 = ~new_n14569 & ~new_n14570;
  assign new_n14572 = new_n14562 & new_n14571;
  assign new_n14573 = ~new_n14562 & ~new_n14571;
  assign new_n14574 = ~new_n14572 & ~new_n14573;
  assign new_n14575 = ~new_n14394 & new_n14574;
  assign new_n14576 = new_n14394 & ~new_n14574;
  assign new_n14577 = ~new_n14575 & ~new_n14576;
  assign new_n14578 = new_n14376 & new_n14577;
  assign new_n14579 = ~new_n14376 & ~new_n14577;
  assign n6192 = ~new_n14578 & ~new_n14579;
  assign new_n14581 = ~new_n932 & ~new_n933;
  assign new_n14582 = new_n967 & ~new_n14581;
  assign new_n14583 = ~new_n967 & new_n14581;
  assign n6273 = new_n14582 | new_n14583;
  assign new_n14585 = ~new_n8814 & ~new_n8815;
  assign new_n14586 = ~new_n8819_1 & new_n14585;
  assign new_n14587 = new_n8819_1 & ~new_n14585;
  assign n6445 = ~new_n14586 & ~new_n14587;
  assign new_n14589 = ~new_n10981 & ~new_n10982;
  assign new_n14590 = new_n11012 & ~new_n14589;
  assign new_n14591 = ~new_n11012 & new_n14589;
  assign n6645 = ~new_n14590 & ~new_n14591;
  assign new_n14593 = ~new_n9298 & ~new_n9299;
  assign new_n14594 = new_n9326 & ~new_n14593;
  assign new_n14595 = ~new_n9326 & new_n14593;
  assign n6689 = ~new_n14594 & ~new_n14595;
  assign new_n14597 = ~new_n1381 & ~new_n1498;
  assign n6742 = ~new_n1499 & ~new_n14597;
  assign new_n14599 = ~new_n2280 & ~new_n2281;
  assign new_n14600 = new_n2333 & ~new_n14599;
  assign new_n14601 = ~new_n2333 & new_n14599;
  assign n6809 = ~new_n14600 & ~new_n14601;
  assign new_n14603 = ~new_n7856 & ~new_n7857;
  assign new_n14604 = new_n7859 & new_n14603;
  assign new_n14605 = ~new_n7859 & ~new_n14603;
  assign n6822 = ~new_n14604 & ~new_n14605;
  assign new_n14607 = ~new_n13125 & ~new_n13126;
  assign new_n14608 = ~new_n13130 & new_n14607;
  assign new_n14609 = new_n13130 & ~new_n14607;
  assign n6860 = new_n14608 | new_n14609;
  assign new_n14611 = ~new_n10997 & ~new_n10998;
  assign new_n14612 = new_n11008 & ~new_n14611;
  assign new_n14613 = ~new_n11008 & new_n14611;
  assign n7193 = ~new_n14612 & ~new_n14613;
  assign new_n14615 = ~new_n8808 & ~new_n8809;
  assign new_n14616 = new_n8821 & ~new_n14615;
  assign new_n14617 = ~new_n8821 & new_n14615;
  assign n7568 = ~new_n14616 & ~new_n14617;
  assign new_n14619 = ~new_n1502 & ~new_n1503;
  assign new_n14620 = ~new_n1507 & ~new_n14619;
  assign new_n14621 = new_n1507 & new_n14619;
  assign n7676 = ~new_n14620 & ~new_n14621;
  assign new_n14623 = ~new_n1066 & ~new_n1070;
  assign new_n14624 = ~new_n530 & ~new_n532;
  assign new_n14625 = new_n14623 & new_n14624;
  assign new_n14626 = ~new_n14623 & ~new_n14624;
  assign new_n14627 = ~new_n14625 & ~new_n14626;
  assign new_n14628 = ~new_n1077 & ~new_n1081;
  assign new_n14629 = ~new_n1080 & ~new_n14628;
  assign new_n14630 = ~new_n1090 & ~new_n1103;
  assign new_n14631 = ~new_n1093 & ~new_n1097_1;
  assign new_n14632 = ~new_n1096 & ~new_n14631;
  assign new_n14633 = n2393 & n12704;
  assign new_n14634 = n5860 & n7294;
  assign new_n14635 = ~new_n14633 & new_n14634;
  assign new_n14636 = new_n14633 & ~new_n14634;
  assign new_n14637 = ~new_n14635 & ~new_n14636;
  assign new_n14638 = n4903 & n7388;
  assign new_n14639 = n5814 & n11892;
  assign new_n14640 = new_n14638 & new_n14639;
  assign new_n14641 = ~new_n14638 & ~new_n14639;
  assign new_n14642 = ~new_n14640 & ~new_n14641;
  assign new_n14643 = new_n14637 & ~new_n14642;
  assign new_n14644 = ~new_n14637 & new_n14642;
  assign new_n14645 = ~new_n14643 & ~new_n14644;
  assign new_n14646 = ~new_n14632 & ~new_n14645;
  assign new_n14647 = new_n14632 & new_n14645;
  assign new_n14648 = ~new_n14646 & ~new_n14647;
  assign new_n14649 = new_n14630 & new_n14648;
  assign new_n14650 = ~new_n14630 & ~new_n14648;
  assign new_n14651 = ~new_n14649 & ~new_n14650;
  assign new_n14652 = new_n14629 & ~new_n14651;
  assign new_n14653 = ~new_n14629 & new_n14651;
  assign new_n14654 = ~new_n14652 & ~new_n14653;
  assign new_n14655 = n5331 & n5694;
  assign new_n14656 = n1564 & n4499;
  assign new_n14657 = new_n14655 & new_n14656;
  assign new_n14658 = ~new_n14655 & ~new_n14656;
  assign new_n14659 = ~new_n14657 & ~new_n14658;
  assign new_n14660 = new_n1110 & ~new_n14659;
  assign new_n14661 = ~new_n1110 & new_n14659;
  assign new_n14662 = ~new_n14660 & ~new_n14661;
  assign new_n14663 = ~new_n14654 & ~new_n14662;
  assign new_n14664 = new_n14654 & new_n14662;
  assign new_n14665 = ~new_n14663 & ~new_n14664;
  assign new_n14666 = ~new_n1046 & ~new_n1055;
  assign new_n14667 = ~new_n1045 & ~new_n14666;
  assign new_n14668 = n2530 & n5069;
  assign new_n14669 = ~new_n1048 & ~new_n1051;
  assign new_n14670 = ~new_n1050 & ~new_n14669;
  assign new_n14671 = ~new_n14668 & new_n14670;
  assign new_n14672 = new_n14668 & ~new_n14670;
  assign new_n14673 = ~new_n14671 & ~new_n14672;
  assign new_n14674 = new_n14667 & ~new_n14673;
  assign new_n14675 = ~new_n14667 & new_n14673;
  assign new_n14676 = ~new_n14674 & ~new_n14675;
  assign new_n14677 = ~new_n1042 & ~new_n1058;
  assign new_n14678 = ~new_n1041 & ~new_n14677;
  assign new_n14679 = new_n14676 & new_n14678;
  assign new_n14680 = ~new_n14676 & ~new_n14678;
  assign new_n14681 = ~new_n14679 & ~new_n14680;
  assign new_n14682 = ~new_n492 & ~new_n525;
  assign new_n14683 = ~new_n493 & ~new_n14682;
  assign new_n14684 = n615 & n5305;
  assign new_n14685 = n6038 & n10547;
  assign new_n14686 = ~new_n14684 & new_n14685;
  assign new_n14687 = new_n14684 & ~new_n14685;
  assign new_n14688 = ~new_n14686 & ~new_n14687;
  assign new_n14689 = ~new_n14683 & ~new_n14688;
  assign new_n14690 = new_n14683 & new_n14688;
  assign new_n14691 = ~new_n14689 & ~new_n14690;
  assign new_n14692 = n8476 & n12044;
  assign new_n14693 = ~new_n1030 & ~new_n1034;
  assign new_n14694 = ~new_n1033 & ~new_n14693;
  assign new_n14695 = ~new_n14692 & new_n14694;
  assign new_n14696 = new_n14692 & ~new_n14694;
  assign new_n14697 = ~new_n14695 & ~new_n14696;
  assign new_n14698 = ~new_n14691 & new_n14697;
  assign new_n14699 = new_n14691 & ~new_n14697;
  assign new_n14700 = ~new_n14698 & ~new_n14699;
  assign new_n14701 = ~new_n14681 & new_n14700;
  assign new_n14702 = new_n14681 & ~new_n14700;
  assign new_n14703 = ~new_n14701 & ~new_n14702;
  assign new_n14704 = ~new_n14665 & new_n14703;
  assign new_n14705 = new_n14665 & ~new_n14703;
  assign new_n14706 = ~new_n14704 & ~new_n14705;
  assign new_n14707 = ~new_n1027 & ~new_n1061;
  assign new_n14708 = ~new_n1028 & ~new_n14707;
  assign new_n14709 = n6806 & n12648;
  assign new_n14710 = n2802 & n10545;
  assign new_n14711 = ~new_n14709 & ~new_n14710;
  assign new_n14712 = new_n14709 & new_n14710;
  assign new_n14713 = ~new_n14711 & ~new_n14712;
  assign new_n14714 = n533 & n7690;
  assign new_n14715 = n1512 & n3616;
  assign new_n14716 = new_n14714 & ~new_n14715;
  assign new_n14717 = ~new_n14714 & new_n14715;
  assign new_n14718 = ~new_n14716 & ~new_n14717;
  assign new_n14719 = ~new_n14713 & ~new_n14718;
  assign new_n14720 = new_n14713 & new_n14718;
  assign new_n14721 = ~new_n14719 & ~new_n14720;
  assign new_n14722 = new_n14708 & new_n14721;
  assign new_n14723 = ~new_n14708 & ~new_n14721;
  assign new_n14724 = ~new_n14722 & ~new_n14723;
  assign new_n14725 = new_n14706 & ~new_n14724;
  assign new_n14726 = ~new_n14706 & new_n14724;
  assign new_n14727 = ~new_n14725 & ~new_n14726;
  assign new_n14728 = ~new_n14627 & new_n14727;
  assign new_n14729 = new_n14627 & ~new_n14727;
  assign new_n14730 = ~new_n14728 & ~new_n14729;
  assign new_n14731 = ~new_n1131 & ~new_n1135;
  assign new_n14732 = ~new_n1132 & ~new_n14731;
  assign new_n14733 = ~new_n1124 & ~new_n1127;
  assign new_n14734 = ~new_n1123 & ~new_n14733;
  assign new_n14735 = ~new_n1117 & ~new_n1121;
  assign new_n14736 = n1980 & n3986;
  assign new_n14737 = n5857 & n10848;
  assign new_n14738 = ~new_n14736 & ~new_n14737;
  assign new_n14739 = new_n14736 & new_n14737;
  assign new_n14740 = ~new_n14738 & ~new_n14739;
  assign new_n14741 = n1906 & n7965;
  assign new_n14742 = n45 & n8028;
  assign new_n14743 = new_n14741 & ~new_n14742;
  assign new_n14744 = ~new_n14741 & new_n14742;
  assign new_n14745 = ~new_n14743 & ~new_n14744;
  assign new_n14746 = ~new_n14740 & ~new_n14745;
  assign new_n14747 = new_n14740 & new_n14745;
  assign new_n14748 = ~new_n14746 & ~new_n14747;
  assign new_n14749 = ~new_n980 & ~new_n984;
  assign new_n14750 = ~new_n983 & ~new_n14749;
  assign new_n14751 = ~new_n14748 & ~new_n14750;
  assign new_n14752 = new_n14748 & new_n14750;
  assign new_n14753 = ~new_n14751 & ~new_n14752;
  assign new_n14754 = ~new_n1074 & new_n1112;
  assign new_n14755 = ~new_n1075 & ~new_n14754;
  assign new_n14756 = ~new_n993 & new_n1004;
  assign new_n14757 = ~new_n994 & ~new_n14756;
  assign new_n14758 = n1209 & n9241;
  assign new_n14759 = n5105 & n8276;
  assign new_n14760 = new_n14758 & ~new_n14759;
  assign new_n14761 = ~new_n14758 & new_n14759;
  assign new_n14762 = ~new_n14760 & ~new_n14761;
  assign new_n14763 = new_n996_1 & ~new_n999;
  assign new_n14764 = ~new_n1000 & ~new_n14763;
  assign new_n14765 = ~new_n14762 & new_n14764;
  assign new_n14766 = new_n14762 & ~new_n14764;
  assign new_n14767 = ~new_n14765 & ~new_n14766;
  assign new_n14768 = n6776 & n8236;
  assign new_n14769 = n4928 & n12299;
  assign new_n14770 = n4141 & n7436;
  assign new_n14771 = ~new_n14769 & ~new_n14770;
  assign new_n14772 = new_n14769 & new_n14770;
  assign new_n14773 = ~new_n14771 & ~new_n14772;
  assign new_n14774 = new_n14768 & new_n14773;
  assign new_n14775 = ~new_n14768 & ~new_n14773;
  assign new_n14776 = ~new_n14774 & ~new_n14775;
  assign new_n14777 = ~new_n14767 & new_n14776;
  assign new_n14778 = new_n14767 & ~new_n14776;
  assign new_n14779 = ~new_n14777 & ~new_n14778;
  assign new_n14780 = new_n14757 & ~new_n14779;
  assign new_n14781 = ~new_n14757 & new_n14779;
  assign new_n14782 = ~new_n14780 & ~new_n14781;
  assign new_n14783 = new_n1011 & ~new_n14782;
  assign new_n14784 = ~new_n1011 & new_n14782;
  assign new_n14785 = ~new_n14783 & ~new_n14784;
  assign new_n14786 = new_n14755 & ~new_n14785;
  assign new_n14787 = ~new_n14755 & new_n14785;
  assign new_n14788 = ~new_n14786 & ~new_n14787;
  assign new_n14789 = ~new_n14753 & new_n14788;
  assign new_n14790 = new_n14753 & ~new_n14788;
  assign new_n14791 = ~new_n14789 & ~new_n14790;
  assign new_n14792 = new_n14735 & new_n14791;
  assign new_n14793 = ~new_n14735 & ~new_n14791;
  assign new_n14794 = ~new_n14792 & ~new_n14793;
  assign new_n14795 = ~new_n1019 & ~new_n1023;
  assign new_n14796 = ~new_n977 & ~new_n1014;
  assign new_n14797 = ~new_n978 & ~new_n14796;
  assign new_n14798 = n7500 & n10510;
  assign new_n14799 = n7354 & n10644;
  assign new_n14800 = n783 & n8759;
  assign new_n14801 = new_n14799 & ~new_n14800;
  assign new_n14802 = ~new_n14799 & new_n14800;
  assign new_n14803 = ~new_n14801 & ~new_n14802;
  assign new_n14804 = new_n14798 & ~new_n14803;
  assign new_n14805 = ~new_n14798 & new_n14803;
  assign new_n14806 = ~new_n14804 & ~new_n14805;
  assign new_n14807 = new_n14797 & new_n14806;
  assign new_n14808 = ~new_n14797 & ~new_n14806;
  assign new_n14809 = ~new_n14807 & ~new_n14808;
  assign new_n14810 = ~new_n509 & new_n519;
  assign new_n14811 = ~new_n508 & ~new_n14810;
  assign new_n14812 = ~new_n504 & new_n522;
  assign new_n14813 = ~new_n505 & ~new_n14812;
  assign new_n14814 = ~new_n14811 & new_n14813;
  assign new_n14815 = new_n14811 & ~new_n14813;
  assign new_n14816 = ~new_n14814 & ~new_n14815;
  assign new_n14817 = new_n495 & ~new_n498;
  assign new_n14818 = ~new_n499 & ~new_n14817;
  assign new_n14819 = n2585 & n4312;
  assign new_n14820 = n1097 & n4005;
  assign new_n14821 = new_n14819 & ~new_n14820;
  assign new_n14822 = ~new_n14819 & new_n14820;
  assign new_n14823 = ~new_n14821 & ~new_n14822;
  assign new_n14824 = n12025 & n12720;
  assign new_n14825 = n2509 & n11257;
  assign new_n14826 = new_n14824 & ~new_n14825;
  assign new_n14827 = ~new_n14824 & new_n14825;
  assign new_n14828 = ~new_n14826 & ~new_n14827;
  assign new_n14829 = ~new_n14823 & new_n14828;
  assign new_n14830 = new_n14823 & ~new_n14828;
  assign new_n14831 = ~new_n14829 & ~new_n14830;
  assign new_n14832 = ~new_n511 & ~new_n515;
  assign new_n14833 = ~new_n514 & ~new_n14832;
  assign new_n14834 = n5964 & n12706;
  assign new_n14835 = n2508 & n12705;
  assign new_n14836 = ~new_n14834 & new_n14835;
  assign new_n14837 = new_n14834 & ~new_n14835;
  assign new_n14838 = ~new_n14836 & ~new_n14837;
  assign new_n14839 = new_n14833 & new_n14838;
  assign new_n14840 = ~new_n14833 & ~new_n14838;
  assign new_n14841 = ~new_n14839 & ~new_n14840;
  assign new_n14842 = new_n14831 & new_n14841;
  assign new_n14843 = ~new_n14831 & ~new_n14841;
  assign new_n14844 = ~new_n14842 & ~new_n14843;
  assign new_n14845 = new_n14818 & new_n14844;
  assign new_n14846 = ~new_n14818 & ~new_n14844;
  assign new_n14847 = ~new_n14845 & ~new_n14846;
  assign new_n14848 = ~new_n14816 & new_n14847;
  assign new_n14849 = new_n14816 & ~new_n14847;
  assign new_n14850 = ~new_n14848 & ~new_n14849;
  assign new_n14851 = new_n14809 & new_n14850;
  assign new_n14852 = ~new_n14809 & ~new_n14850;
  assign new_n14853 = ~new_n14851 & ~new_n14852;
  assign new_n14854 = ~new_n14795 & new_n14853;
  assign new_n14855 = new_n14795 & ~new_n14853;
  assign new_n14856 = ~new_n14854 & ~new_n14855;
  assign new_n14857 = ~new_n14794 & new_n14856;
  assign new_n14858 = new_n14794 & ~new_n14856;
  assign new_n14859 = ~new_n14857 & ~new_n14858;
  assign new_n14860 = ~new_n14734 & ~new_n14859;
  assign new_n14861 = new_n14734 & new_n14859;
  assign new_n14862 = ~new_n14860 & ~new_n14861;
  assign new_n14863 = new_n14732 & new_n14862;
  assign new_n14864 = ~new_n14732 & ~new_n14862;
  assign new_n14865 = ~new_n14863 & ~new_n14864;
  assign new_n14866 = new_n14730 & new_n14865;
  assign new_n14867 = ~new_n14730 & ~new_n14865;
  assign new_n14868 = ~new_n14866 & ~new_n14867;
  assign new_n14869 = ~new_n972 & ~new_n1138_1;
  assign new_n14870 = ~new_n973 & ~new_n14869;
  assign new_n14871 = ~new_n14868 & new_n14870;
  assign new_n14872 = new_n14868 & ~new_n14870;
  assign n7966 = new_n14871 | new_n14872;
  assign new_n14874 = ~new_n14322 & ~new_n14323;
  assign new_n14875 = ~new_n14325 & new_n14874;
  assign new_n14876 = new_n14325 & ~new_n14874;
  assign n7981 = ~new_n14875 & ~new_n14876;
  assign new_n14878 = ~new_n13814 & ~new_n13828;
  assign new_n14879 = ~new_n13815 & ~new_n14878;
  assign new_n14880 = new_n13758 & ~new_n13761;
  assign new_n14881 = ~new_n13762 & ~new_n14880;
  assign new_n14882 = new_n13789 & new_n14881;
  assign new_n14883 = ~new_n13789 & ~new_n14881;
  assign new_n14884 = ~new_n14882 & ~new_n14883;
  assign new_n14885 = new_n14879 & ~new_n14884;
  assign new_n14886 = ~new_n14879 & new_n14884;
  assign new_n14887 = ~new_n14885 & ~new_n14886;
  assign new_n14888 = ~new_n13509 & ~new_n13520;
  assign new_n14889 = ~new_n13603 & ~new_n13605;
  assign new_n14890 = ~new_n13488 & new_n13498;
  assign new_n14891 = ~new_n13487 & ~new_n14890;
  assign new_n14892 = n5320 & n6770;
  assign new_n14893 = n3627 & n11877;
  assign new_n14894 = n4516 & n5212;
  assign new_n14895 = ~new_n14893 & new_n14894;
  assign new_n14896 = new_n14893 & ~new_n14894;
  assign new_n14897 = ~new_n14895 & ~new_n14896;
  assign new_n14898 = new_n14892 & new_n14897;
  assign new_n14899 = ~new_n14892 & ~new_n14897;
  assign new_n14900 = ~new_n14898 & ~new_n14899;
  assign new_n14901 = n2564 & n9725;
  assign new_n14902 = n4370 & n9920;
  assign new_n14903 = ~new_n14901 & new_n14902;
  assign new_n14904 = new_n14901 & ~new_n14902;
  assign new_n14905 = ~new_n14903 & ~new_n14904;
  assign new_n14906 = ~new_n14900 & new_n14905;
  assign new_n14907 = new_n14900 & ~new_n14905;
  assign new_n14908 = ~new_n14906 & ~new_n14907;
  assign new_n14909 = n4189 & n12000;
  assign new_n14910 = ~new_n13490 & ~new_n13494;
  assign new_n14911 = ~new_n13493 & ~new_n14910;
  assign new_n14912 = new_n14909 & new_n14911;
  assign new_n14913 = ~new_n14909 & ~new_n14911;
  assign new_n14914 = ~new_n14912 & ~new_n14913;
  assign new_n14915 = ~new_n14908 & new_n14914;
  assign new_n14916 = new_n14908 & ~new_n14914;
  assign new_n14917 = ~new_n14915 & ~new_n14916;
  assign new_n14918 = new_n14891 & ~new_n14917;
  assign new_n14919 = ~new_n14891 & new_n14917;
  assign new_n14920 = ~new_n14918 & ~new_n14919;
  assign new_n14921 = ~new_n13562 & ~new_n13598;
  assign new_n14922 = ~new_n13563 & ~new_n14921;
  assign new_n14923 = n7320 & n11728;
  assign new_n14924 = n7523 & n12709;
  assign new_n14925 = n1198 & n8336;
  assign new_n14926 = new_n14924 & ~new_n14925;
  assign new_n14927 = ~new_n14924 & new_n14925;
  assign new_n14928 = ~new_n14926 & ~new_n14927;
  assign new_n14929 = new_n14923 & ~new_n14928;
  assign new_n14930 = ~new_n14923 & new_n14928;
  assign new_n14931 = ~new_n14929 & ~new_n14930;
  assign new_n14932 = new_n14922 & new_n14931;
  assign new_n14933 = ~new_n14922 & ~new_n14931;
  assign new_n14934 = ~new_n14932 & ~new_n14933;
  assign new_n14935 = new_n13474 & ~new_n13477;
  assign new_n14936 = ~new_n13478 & ~new_n14935;
  assign new_n14937 = ~new_n14934 & new_n14936;
  assign new_n14938 = new_n14934 & ~new_n14936;
  assign new_n14939 = ~new_n14937 & ~new_n14938;
  assign new_n14940 = ~new_n14920 & new_n14939;
  assign new_n14941 = new_n14920 & ~new_n14939;
  assign new_n14942 = ~new_n14940 & ~new_n14941;
  assign new_n14943 = new_n14889 & ~new_n14942;
  assign new_n14944 = ~new_n14889 & new_n14942;
  assign new_n14945 = ~new_n14943 & ~new_n14944;
  assign new_n14946 = ~new_n13804 & ~new_n13807;
  assign new_n14947 = ~new_n13803 & ~new_n14946;
  assign new_n14948 = ~new_n13747 & ~new_n13751;
  assign new_n14949 = n1478 & n5319;
  assign new_n14950 = n5760 & n9457;
  assign new_n14951 = ~new_n14949 & ~new_n14950;
  assign new_n14952 = new_n14949 & new_n14950;
  assign new_n14953 = ~new_n14951 & ~new_n14952;
  assign new_n14954 = n10022 & n11222;
  assign new_n14955 = n4817 & n10990;
  assign new_n14956 = new_n14954 & ~new_n14955;
  assign new_n14957 = ~new_n14954 & new_n14955;
  assign new_n14958 = ~new_n14956 & ~new_n14957;
  assign new_n14959 = ~new_n14953 & ~new_n14958;
  assign new_n14960 = new_n14953 & new_n14958;
  assign new_n14961 = ~new_n14959 & ~new_n14960;
  assign new_n14962 = ~new_n13565 & ~new_n13569;
  assign new_n14963 = ~new_n13568 & ~new_n14962;
  assign new_n14964 = ~new_n14961 & ~new_n14963;
  assign new_n14965 = new_n14961 & new_n14963;
  assign new_n14966 = ~new_n14964 & ~new_n14965;
  assign new_n14967 = ~new_n13709 & ~new_n13742;
  assign new_n14968 = ~new_n13710 & ~new_n14967;
  assign new_n14969 = ~new_n13576 & new_n13595;
  assign new_n14970 = ~new_n13577 & ~new_n14969;
  assign new_n14971 = ~new_n13580 & ~new_n13593;
  assign new_n14972 = n1094 & n8819;
  assign new_n14973 = n6429 & n10678;
  assign new_n14974 = new_n14972 & ~new_n14973;
  assign new_n14975 = ~new_n14972 & new_n14973;
  assign new_n14976 = ~new_n14974 & ~new_n14975;
  assign new_n14977 = ~new_n13583 & ~new_n13587;
  assign new_n14978 = ~new_n13586 & ~new_n14977;
  assign new_n14979 = ~new_n14976 & new_n14978;
  assign new_n14980 = new_n14976 & ~new_n14978;
  assign new_n14981 = ~new_n14979 & ~new_n14980;
  assign new_n14982 = n7730 & n10928;
  assign new_n14983 = n6986 & n8717;
  assign new_n14984 = n2226 & n2433;
  assign new_n14985 = ~new_n14983 & ~new_n14984;
  assign new_n14986 = new_n14983 & new_n14984;
  assign new_n14987 = ~new_n14985 & ~new_n14986;
  assign new_n14988 = new_n14982 & new_n14987;
  assign new_n14989 = ~new_n14982 & ~new_n14987;
  assign new_n14990 = ~new_n14988 & ~new_n14989;
  assign new_n14991 = new_n14981 & new_n14990;
  assign new_n14992 = ~new_n14981 & ~new_n14990;
  assign new_n14993 = ~new_n14991 & ~new_n14992;
  assign new_n14994 = ~new_n14971 & new_n14993;
  assign new_n14995 = new_n14971 & ~new_n14993;
  assign new_n14996 = ~new_n14994 & ~new_n14995;
  assign new_n14997 = new_n14970 & new_n14996;
  assign new_n14998 = ~new_n14970 & ~new_n14996;
  assign new_n14999 = ~new_n14997 & ~new_n14998;
  assign new_n15000 = ~new_n14968 & new_n14999;
  assign new_n15001 = new_n14968 & ~new_n14999;
  assign new_n15002 = ~new_n15000 & ~new_n15001;
  assign new_n15003 = ~new_n14966 & new_n15002;
  assign new_n15004 = new_n14966 & ~new_n15002;
  assign new_n15005 = ~new_n15003 & ~new_n15004;
  assign new_n15006 = new_n14948 & new_n15005;
  assign new_n15007 = ~new_n14948 & ~new_n15005;
  assign new_n15008 = ~new_n15006 & ~new_n15007;
  assign new_n15009 = ~new_n13484 & ~new_n13501;
  assign new_n15010 = ~new_n13483 & ~new_n15009;
  assign new_n15011 = ~new_n15008 & new_n15010;
  assign new_n15012 = new_n15008 & ~new_n15010;
  assign new_n15013 = ~new_n15011 & ~new_n15012;
  assign new_n15014 = ~new_n14947 & ~new_n15013;
  assign new_n15015 = new_n14947 & new_n15013;
  assign new_n15016 = ~new_n15014 & ~new_n15015;
  assign new_n15017 = ~new_n14945 & new_n15016;
  assign new_n15018 = new_n14945 & ~new_n15016;
  assign new_n15019 = ~new_n15017 & ~new_n15018;
  assign new_n15020 = ~new_n13797 & ~new_n13801;
  assign new_n15021 = ~new_n13722 & ~new_n13739;
  assign new_n15022 = ~new_n13721 & ~new_n15021;
  assign new_n15023 = ~new_n13726 & ~new_n13736;
  assign new_n15024 = ~new_n13725 & ~new_n15023;
  assign new_n15025 = n11153 & n11999;
  assign new_n15026 = n996 & n12947;
  assign new_n15027 = n5767 & n11791;
  assign new_n15028 = ~new_n15026 & new_n15027;
  assign new_n15029 = new_n15026 & ~new_n15027;
  assign new_n15030 = ~new_n15028 & ~new_n15029;
  assign new_n15031 = new_n15025 & new_n15030;
  assign new_n15032 = ~new_n15025 & ~new_n15030;
  assign new_n15033 = ~new_n15031 & ~new_n15032;
  assign new_n15034 = ~new_n13712 & ~new_n13716;
  assign new_n15035 = ~new_n13715 & ~new_n15034;
  assign new_n15036 = ~new_n15033 & new_n15035;
  assign new_n15037 = new_n15033 & ~new_n15035;
  assign new_n15038 = ~new_n15036 & ~new_n15037;
  assign new_n15039 = new_n15024 & ~new_n15038;
  assign new_n15040 = ~new_n15024 & new_n15038;
  assign new_n15041 = ~new_n15039 & ~new_n15040;
  assign new_n15042 = new_n15022 & new_n15041;
  assign new_n15043 = ~new_n15022 & ~new_n15041;
  assign new_n15044 = ~new_n15042 & ~new_n15043;
  assign new_n15045 = n7160 & n11967;
  assign new_n15046 = n4828 & n6254;
  assign new_n15047 = ~new_n15045 & ~new_n15046;
  assign new_n15048 = new_n15045 & new_n15046;
  assign new_n15049 = ~new_n15047 & ~new_n15048;
  assign new_n15050 = n2515 & n12777;
  assign new_n15051 = n1199 & n7159;
  assign new_n15052 = new_n15050 & ~new_n15051;
  assign new_n15053 = ~new_n15050 & new_n15051;
  assign new_n15054 = ~new_n15052 & ~new_n15053;
  assign new_n15055 = ~new_n15049 & ~new_n15054;
  assign new_n15056 = new_n15049 & new_n15054;
  assign new_n15057 = ~new_n15055 & ~new_n15056;
  assign new_n15058 = ~new_n13728 & ~new_n13732;
  assign new_n15059 = ~new_n13731 & ~new_n15058;
  assign new_n15060 = n4436 & n12069;
  assign new_n15061 = n5314 & n6441;
  assign new_n15062 = new_n15060 & ~new_n15061;
  assign new_n15063 = ~new_n15060 & new_n15061;
  assign new_n15064 = ~new_n15062 & ~new_n15063;
  assign new_n15065 = ~new_n15059 & new_n15064;
  assign new_n15066 = new_n15059 & ~new_n15064;
  assign new_n15067 = ~new_n15065 & ~new_n15066;
  assign new_n15068 = ~new_n15057 & new_n15067;
  assign new_n15069 = new_n15057 & ~new_n15067;
  assign new_n15070 = ~new_n15068 & ~new_n15069;
  assign new_n15071 = ~new_n15044 & new_n15070;
  assign new_n15072 = new_n15044 & ~new_n15070;
  assign new_n15073 = ~new_n15071 & ~new_n15072;
  assign new_n15074 = n6578 & n12489;
  assign new_n15075 = ~new_n13755 & ~new_n13792;
  assign new_n15076 = ~new_n13756 & ~new_n15075;
  assign new_n15077 = new_n15074 & new_n15076;
  assign new_n15078 = ~new_n15074 & ~new_n15076;
  assign new_n15079 = ~new_n15077 & ~new_n15078;
  assign new_n15080 = new_n15073 & new_n15079;
  assign new_n15081 = ~new_n15073 & ~new_n15079;
  assign new_n15082 = ~new_n15080 & ~new_n15081;
  assign new_n15083 = ~new_n13470 & new_n13504;
  assign new_n15084 = ~new_n13471 & ~new_n15083;
  assign new_n15085 = ~new_n13772 & ~new_n13782;
  assign new_n15086 = ~new_n13771 & ~new_n15085;
  assign new_n15087 = ~new_n13774 & ~new_n13778;
  assign new_n15088 = ~new_n13777 & ~new_n15087;
  assign new_n15089 = n1353 & n12391;
  assign new_n15090 = n447 & n7891;
  assign new_n15091 = new_n15089 & ~new_n15090;
  assign new_n15092 = ~new_n15089 & new_n15090;
  assign new_n15093 = ~new_n15091 & ~new_n15092;
  assign new_n15094 = new_n15088 & ~new_n15093;
  assign new_n15095 = ~new_n15088 & new_n15093;
  assign new_n15096 = ~new_n15094 & ~new_n15095;
  assign new_n15097 = ~new_n15086 & new_n15096;
  assign new_n15098 = new_n15086 & ~new_n15096;
  assign new_n15099 = ~new_n15097 & ~new_n15098;
  assign new_n15100 = n2087 & n11407;
  assign new_n15101 = n6604 & n6687;
  assign new_n15102 = new_n15100 & new_n15101;
  assign new_n15103 = ~new_n15100 & ~new_n15101;
  assign new_n15104 = ~new_n15102 & ~new_n15103;
  assign new_n15105 = new_n15099 & ~new_n15104;
  assign new_n15106 = ~new_n15099 & new_n15104;
  assign new_n15107 = ~new_n15105 & ~new_n15106;
  assign new_n15108 = ~new_n15084 & new_n15107;
  assign new_n15109 = new_n15084 & ~new_n15107;
  assign new_n15110 = ~new_n15108 & ~new_n15109;
  assign new_n15111 = ~new_n15082 & new_n15110;
  assign new_n15112 = new_n15082 & ~new_n15110;
  assign new_n15113 = ~new_n15111 & ~new_n15112;
  assign new_n15114 = new_n15020 & new_n15113;
  assign new_n15115 = ~new_n15020 & ~new_n15113;
  assign new_n15116 = ~new_n15114 & ~new_n15115;
  assign new_n15117 = ~new_n13705 & new_n13810;
  assign new_n15118 = ~new_n13704 & ~new_n15117;
  assign new_n15119 = new_n15116 & new_n15118;
  assign new_n15120 = ~new_n15116 & ~new_n15118;
  assign new_n15121 = ~new_n15119 & ~new_n15120;
  assign new_n15122 = new_n15019 & new_n15121;
  assign new_n15123 = ~new_n15019 & ~new_n15121;
  assign new_n15124 = ~new_n15122 & ~new_n15123;
  assign new_n15125 = ~new_n14888 & new_n15124;
  assign new_n15126 = new_n14888 & ~new_n15124;
  assign new_n15127 = ~new_n15125 & ~new_n15126;
  assign new_n15128 = new_n14887 & ~new_n15127;
  assign new_n15129 = ~new_n14887 & new_n15127;
  assign n8100 = ~new_n15128 & ~new_n15129;
  assign new_n15131 = ~new_n11001 & ~new_n11002;
  assign new_n15132 = ~new_n11006 & new_n15131;
  assign new_n15133 = new_n11006 & ~new_n15131;
  assign n8138 = new_n15132 | new_n15133;
  assign new_n15135 = ~new_n6665 & ~new_n6666;
  assign new_n15136 = ~new_n6670 & new_n15135;
  assign new_n15137 = new_n6670 & ~new_n15135;
  assign n8202 = new_n15136 | new_n15137;
  assign new_n15139 = ~new_n3611 & ~new_n4009;
  assign n8303 = ~new_n4010 & ~new_n15139;
  assign new_n15141 = ~new_n3313 & ~new_n3314;
  assign new_n15142 = ~new_n3318 & new_n15141;
  assign new_n15143 = new_n3318 & ~new_n15141;
  assign n8398 = new_n15142 | new_n15143;
  assign new_n15145 = ~new_n4790 & ~new_n4791;
  assign new_n15146 = ~new_n4795 & new_n15145;
  assign new_n15147 = new_n4795 & ~new_n15145;
  assign n9137 = new_n15146 | new_n15147;
  assign new_n15149 = ~new_n7862_1 & ~new_n7863;
  assign new_n15150 = new_n7998 & new_n15149;
  assign new_n15151 = ~new_n7998 & ~new_n15149;
  assign n9387 = ~new_n15150 & ~new_n15151;
  assign new_n15153 = ~new_n13139 & ~new_n13140;
  assign new_n15154 = ~new_n13144 & new_n15153;
  assign new_n15155 = new_n13144 & ~new_n15153;
  assign n9571 = new_n15154 | new_n15155;
  assign new_n15157 = ~new_n924 & ~new_n925;
  assign new_n15158 = new_n969 & new_n15157;
  assign new_n15159 = ~new_n969 & ~new_n15157;
  assign n9578 = ~new_n15158 & ~new_n15159;
  assign new_n15161 = ~new_n1260 & ~new_n1261;
  assign new_n15162 = new_n1275 & ~new_n15161;
  assign new_n15163 = ~new_n1275 & new_n15161;
  assign n9706 = ~new_n15162 & ~new_n15163;
  assign new_n15165 = ~new_n4782 & ~new_n4783;
  assign new_n15166 = new_n4797 & ~new_n15165;
  assign new_n15167 = ~new_n4797 & new_n15165;
  assign n9756 = ~new_n15166 & ~new_n15167;
  assign new_n15169 = ~new_n7602 & new_n7626;
  assign new_n15170 = ~new_n7603 & ~new_n15169;
  assign new_n15171 = ~new_n7151 & ~new_n7188;
  assign new_n15172 = ~new_n7152 & ~new_n15171;
  assign new_n15173 = ~new_n7411 & new_n7421;
  assign new_n15174 = ~new_n7410 & ~new_n15173;
  assign new_n15175 = new_n7413 & ~new_n7416;
  assign new_n15176 = ~new_n7417 & ~new_n15175;
  assign new_n15177 = n4094 & n12391;
  assign new_n15178 = n7891 & n12826;
  assign new_n15179 = ~new_n15177 & new_n15178;
  assign new_n15180 = new_n15177 & ~new_n15178;
  assign new_n15181 = ~new_n15179 & ~new_n15180;
  assign new_n15182 = new_n15176 & ~new_n15181;
  assign new_n15183 = ~new_n15176 & new_n15181;
  assign new_n15184 = ~new_n15182 & ~new_n15183;
  assign new_n15185 = ~new_n15174 & ~new_n15184;
  assign new_n15186 = new_n15174 & new_n15184;
  assign new_n15187 = ~new_n15185 & ~new_n15186;
  assign new_n15188 = n1798 & n2087;
  assign new_n15189 = n753 & n6687;
  assign new_n15190 = new_n15188 & new_n15189;
  assign new_n15191 = ~new_n15188 & ~new_n15189;
  assign new_n15192 = ~new_n15190 & ~new_n15191;
  assign new_n15193 = new_n15187 & ~new_n15192;
  assign new_n15194 = ~new_n15187 & new_n15192;
  assign new_n15195 = ~new_n15193 & ~new_n15194;
  assign new_n15196 = ~new_n15172 & ~new_n15195;
  assign new_n15197 = new_n15172 & new_n15195;
  assign new_n15198 = ~new_n15196 & ~new_n15197;
  assign new_n15199 = ~new_n7392 & ~new_n7427;
  assign new_n15200 = ~new_n7393 & ~new_n15199;
  assign new_n15201 = n2551 & n7160;
  assign new_n15202 = n4828 & n11922;
  assign new_n15203 = ~new_n15201 & ~new_n15202;
  assign new_n15204 = new_n15201 & new_n15202;
  assign new_n15205 = ~new_n15203 & ~new_n15204;
  assign new_n15206 = n2515 & n8665;
  assign new_n15207 = n1067 & n1199;
  assign new_n15208 = new_n15206 & ~new_n15207;
  assign new_n15209 = ~new_n15206 & new_n15207;
  assign new_n15210 = ~new_n15208 & ~new_n15209;
  assign new_n15211 = ~new_n15205 & ~new_n15210;
  assign new_n15212 = new_n15205 & new_n15210;
  assign new_n15213 = ~new_n15211 & ~new_n15212;
  assign new_n15214 = ~new_n15200 & new_n15213;
  assign new_n15215 = new_n15200 & ~new_n15213;
  assign new_n15216 = ~new_n15214 & ~new_n15215;
  assign new_n15217 = ~new_n7520 & ~new_n7537;
  assign new_n15218 = ~new_n7519 & ~new_n15217;
  assign new_n15219 = ~new_n7523_1 & ~new_n7534;
  assign new_n15220 = ~new_n7524 & ~new_n15219;
  assign new_n15221 = new_n15218 & new_n15220;
  assign new_n15222 = ~new_n15218 & ~new_n15220;
  assign new_n15223 = ~new_n15221 & ~new_n15222;
  assign new_n15224 = n5645 & n6578;
  assign new_n15225 = n11153 & n12247;
  assign new_n15226 = n159 & n996;
  assign new_n15227 = n2749 & n5767;
  assign new_n15228 = ~new_n15226 & new_n15227;
  assign new_n15229 = new_n15226 & ~new_n15227;
  assign new_n15230 = ~new_n15228 & ~new_n15229;
  assign new_n15231 = new_n15225 & new_n15230;
  assign new_n15232 = ~new_n15225 & ~new_n15230;
  assign new_n15233 = ~new_n15231 & ~new_n15232;
  assign new_n15234 = ~new_n7508 & ~new_n7512;
  assign new_n15235 = ~new_n7511 & ~new_n15234;
  assign new_n15236 = ~new_n15233 & new_n15235;
  assign new_n15237 = new_n15233 & ~new_n15235;
  assign new_n15238 = ~new_n15236 & ~new_n15237;
  assign new_n15239 = ~new_n7526 & ~new_n7530;
  assign new_n15240 = ~new_n7529 & ~new_n15239;
  assign new_n15241 = n10685 & n12069;
  assign new_n15242 = n1510 & n5314;
  assign new_n15243 = new_n15241 & ~new_n15242;
  assign new_n15244 = ~new_n15241 & new_n15242;
  assign new_n15245 = ~new_n15243 & ~new_n15244;
  assign new_n15246 = ~new_n15240 & ~new_n15245;
  assign new_n15247 = new_n15240 & new_n15245;
  assign new_n15248 = ~new_n15246 & ~new_n15247;
  assign new_n15249 = ~new_n15238 & new_n15248;
  assign new_n15250 = new_n15238 & ~new_n15248;
  assign new_n15251 = ~new_n15249 & ~new_n15250;
  assign new_n15252 = new_n15224 & new_n15251;
  assign new_n15253 = ~new_n15224 & ~new_n15251;
  assign new_n15254 = ~new_n15252 & ~new_n15253;
  assign new_n15255 = new_n15223 & ~new_n15254;
  assign new_n15256 = ~new_n15223 & new_n15254;
  assign new_n15257 = ~new_n15255 & ~new_n15256;
  assign new_n15258 = ~new_n15216 & ~new_n15257;
  assign new_n15259 = new_n15216 & new_n15257;
  assign new_n15260 = ~new_n15258 & ~new_n15259;
  assign new_n15261 = ~new_n7407 & ~new_n7424;
  assign new_n15262 = ~new_n7406 & ~new_n15261;
  assign new_n15263 = ~new_n7395 & ~new_n7399;
  assign new_n15264 = ~new_n7398 & ~new_n15263;
  assign new_n15265 = ~new_n15262 & ~new_n15264;
  assign new_n15266 = new_n15262 & new_n15264;
  assign new_n15267 = ~new_n15265 & ~new_n15266;
  assign new_n15268 = ~new_n15260 & new_n15267;
  assign new_n15269 = new_n15260 & ~new_n15267;
  assign new_n15270 = ~new_n15268 & ~new_n15269;
  assign new_n15271 = ~new_n15198 & new_n15270;
  assign new_n15272 = new_n15198 & ~new_n15270;
  assign new_n15273 = ~new_n15271 & ~new_n15272;
  assign new_n15274 = ~new_n7432 & ~new_n7434;
  assign new_n15275 = ~new_n7193_1 & ~new_n7209;
  assign new_n15276 = new_n15274 & new_n15275;
  assign new_n15277 = ~new_n15274 & ~new_n15275;
  assign new_n15278 = ~new_n15276 & ~new_n15277;
  assign new_n15279 = new_n15273 & new_n15278;
  assign new_n15280 = ~new_n15273 & ~new_n15278;
  assign new_n15281 = ~new_n15279 & ~new_n15280;
  assign new_n15282 = ~new_n7574 & new_n7598;
  assign new_n15283 = ~new_n7575 & ~new_n15282;
  assign new_n15284 = ~new_n7505 & ~new_n7540;
  assign new_n15285 = ~new_n7506 & ~new_n15284;
  assign new_n15286 = new_n7436_1 & ~new_n7569;
  assign new_n15287 = ~new_n7568_1 & ~new_n15286;
  assign new_n15288 = new_n15285 & new_n15287;
  assign new_n15289 = ~new_n15285 & ~new_n15287;
  assign new_n15290 = ~new_n15288 & ~new_n15289;
  assign new_n15291 = n3754 & n5319;
  assign new_n15292 = n9457 & n10898;
  assign new_n15293 = ~new_n15291 & ~new_n15292;
  assign new_n15294 = new_n15291 & new_n15292;
  assign new_n15295 = ~new_n15293 & ~new_n15294;
  assign new_n15296 = n11222 & n12511;
  assign new_n15297 = n4817 & n11876;
  assign new_n15298 = new_n15296 & ~new_n15297;
  assign new_n15299 = ~new_n15296 & new_n15297;
  assign new_n15300 = ~new_n15298 & ~new_n15299;
  assign new_n15301 = ~new_n15295 & ~new_n15300;
  assign new_n15302 = new_n15295 & new_n15300;
  assign new_n15303 = ~new_n15301 & ~new_n15302;
  assign new_n15304 = ~new_n7545 & ~new_n7547;
  assign new_n15305 = ~new_n7297 & ~new_n7308;
  assign new_n15306 = ~new_n7298 & ~new_n15305;
  assign new_n15307 = n1094 & n11023;
  assign new_n15308 = n3022 & n10678;
  assign new_n15309 = ~new_n15307 & new_n15308;
  assign new_n15310 = new_n15307 & ~new_n15308;
  assign new_n15311 = ~new_n15309 & ~new_n15310;
  assign new_n15312 = n6986 & n10278;
  assign new_n15313 = n10928 & n11423;
  assign new_n15314 = ~new_n15312 & new_n15313;
  assign new_n15315 = new_n15312 & ~new_n15313;
  assign new_n15316 = ~new_n15314 & ~new_n15315;
  assign new_n15317 = ~new_n15311 & ~new_n15316;
  assign new_n15318 = new_n15311 & new_n15316;
  assign new_n15319 = ~new_n15317 & ~new_n15318;
  assign new_n15320 = ~new_n7282 & ~new_n7286;
  assign new_n15321 = ~new_n7285 & ~new_n15320;
  assign new_n15322 = ~new_n15319 & new_n15321;
  assign new_n15323 = new_n15319 & ~new_n15321;
  assign new_n15324 = ~new_n15322 & ~new_n15323;
  assign new_n15325 = new_n15306 & ~new_n15324;
  assign new_n15326 = ~new_n15306 & new_n15324;
  assign new_n15327 = ~new_n15325 & ~new_n15326;
  assign new_n15328 = ~new_n7294_1 & ~new_n7311;
  assign new_n15329 = ~new_n7293 & ~new_n15328;
  assign new_n15330 = n2226 & n10451;
  assign new_n15331 = ~new_n7300 & ~new_n7304;
  assign new_n15332 = ~new_n7303 & ~new_n15331;
  assign new_n15333 = ~new_n15330 & new_n15332;
  assign new_n15334 = new_n15330 & ~new_n15332;
  assign new_n15335 = ~new_n15333 & ~new_n15334;
  assign new_n15336 = new_n15329 & new_n15335;
  assign new_n15337 = ~new_n15329 & ~new_n15335;
  assign new_n15338 = ~new_n15336 & ~new_n15337;
  assign new_n15339 = ~new_n15327 & new_n15338;
  assign new_n15340 = new_n15327 & ~new_n15338;
  assign new_n15341 = ~new_n15339 & ~new_n15340;
  assign new_n15342 = new_n15304 & new_n15341;
  assign new_n15343 = ~new_n15304 & ~new_n15341;
  assign new_n15344 = ~new_n15342 & ~new_n15343;
  assign new_n15345 = ~new_n7319 & ~new_n7321;
  assign new_n15346 = ~new_n7154 & ~new_n7158;
  assign new_n15347 = ~new_n7157 & ~new_n15346;
  assign new_n15348 = ~new_n7185 & ~new_n15347;
  assign new_n15349 = new_n7185 & new_n15347;
  assign new_n15350 = ~new_n15348 & ~new_n15349;
  assign new_n15351 = ~new_n7279 & ~new_n7314;
  assign new_n15352 = ~new_n7280 & ~new_n15351;
  assign new_n15353 = n7320 & n9640;
  assign new_n15354 = n6703 & n7523;
  assign new_n15355 = n2278 & n8336;
  assign new_n15356 = ~new_n15354 & new_n15355;
  assign new_n15357 = new_n15354 & ~new_n15355;
  assign new_n15358 = ~new_n15356 & ~new_n15357;
  assign new_n15359 = new_n15353 & ~new_n15358;
  assign new_n15360 = ~new_n15353 & new_n15358;
  assign new_n15361 = ~new_n15359 & ~new_n15360;
  assign new_n15362 = new_n15352 & new_n15361;
  assign new_n15363 = ~new_n15352 & ~new_n15361;
  assign new_n15364 = ~new_n15362 & ~new_n15363;
  assign new_n15365 = ~new_n15350 & new_n15364;
  assign new_n15366 = new_n15350 & ~new_n15364;
  assign new_n15367 = ~new_n15365 & ~new_n15366;
  assign new_n15368 = new_n7170 & ~new_n7173;
  assign new_n15369 = ~new_n7174 & ~new_n15368;
  assign new_n15370 = n2564 & n9583;
  assign new_n15371 = n7456 & n9920;
  assign new_n15372 = n4189 & n10327;
  assign new_n15373 = new_n15371 & new_n15372;
  assign new_n15374 = ~new_n15371 & ~new_n15372;
  assign new_n15375 = ~new_n15373 & ~new_n15374;
  assign new_n15376 = new_n15370 & ~new_n15375;
  assign new_n15377 = ~new_n15370 & new_n15375;
  assign new_n15378 = ~new_n15376 & ~new_n15377;
  assign new_n15379 = ~new_n15369 & new_n15378;
  assign new_n15380 = new_n15369 & ~new_n15378;
  assign new_n15381 = ~new_n15379 & ~new_n15380;
  assign new_n15382 = n3627 & n12591;
  assign new_n15383 = n3932 & n4516;
  assign new_n15384 = ~new_n15382 & new_n15383;
  assign new_n15385 = new_n15382 & ~new_n15383;
  assign new_n15386 = ~new_n15384 & ~new_n15385;
  assign new_n15387 = ~new_n15381 & new_n15386;
  assign new_n15388 = new_n15381 & ~new_n15386;
  assign new_n15389 = ~new_n15387 & ~new_n15388;
  assign new_n15390 = n6770 & n11662;
  assign new_n15391 = ~new_n7167 & new_n7178;
  assign new_n15392 = ~new_n7168 & ~new_n15391;
  assign new_n15393 = new_n15390 & new_n15392;
  assign new_n15394 = ~new_n15390 & ~new_n15392;
  assign new_n15395 = ~new_n15393 & ~new_n15394;
  assign new_n15396 = new_n15389 & new_n15395;
  assign new_n15397 = ~new_n15389 & ~new_n15395;
  assign new_n15398 = ~new_n15396 & ~new_n15397;
  assign new_n15399 = ~new_n15367 & new_n15398;
  assign new_n15400 = new_n15367 & ~new_n15398;
  assign new_n15401 = ~new_n15399 & ~new_n15400;
  assign new_n15402 = new_n15345 & new_n15401;
  assign new_n15403 = ~new_n15345 & ~new_n15401;
  assign new_n15404 = ~new_n15402 & ~new_n15403;
  assign new_n15405 = ~new_n15344 & new_n15404;
  assign new_n15406 = new_n15344 & ~new_n15404;
  assign new_n15407 = ~new_n15405 & ~new_n15406;
  assign new_n15408 = new_n15303 & new_n15407;
  assign new_n15409 = ~new_n15303 & ~new_n15407;
  assign new_n15410 = ~new_n15408 & ~new_n15409;
  assign new_n15411 = new_n15290 & ~new_n15410;
  assign new_n15412 = ~new_n15290 & new_n15410;
  assign new_n15413 = ~new_n15411 & ~new_n15412;
  assign new_n15414 = ~new_n15283 & ~new_n15413;
  assign new_n15415 = new_n15283 & new_n15413;
  assign new_n15416 = ~new_n15414 & ~new_n15415;
  assign new_n15417 = ~new_n15281 & new_n15416;
  assign new_n15418 = new_n15281 & ~new_n15416;
  assign new_n15419 = ~new_n15417 & ~new_n15418;
  assign new_n15420 = ~new_n15170 & ~new_n15419;
  assign new_n15421 = new_n15170 & new_n15419;
  assign n9767 = ~new_n15420 & ~new_n15421;
  assign new_n15423 = ~new_n2318 & ~new_n2319;
  assign new_n15424 = ~new_n2323 & new_n15423;
  assign new_n15425 = new_n2323 & ~new_n15423;
  assign n9820 = new_n15424 | new_n15425;
  assign new_n15427 = ~new_n10971 & ~new_n10972;
  assign new_n15428 = ~new_n11022 & new_n15427;
  assign new_n15429 = new_n11022 & ~new_n15427;
  assign n9938 = new_n15428 | new_n15429;
  assign new_n15431 = ~new_n940 & ~new_n941;
  assign new_n15432 = new_n965 & new_n15431;
  assign new_n15433 = ~new_n965 & ~new_n15431;
  assign n10476 = new_n15432 | new_n15433;
  assign new_n15435 = ~new_n948 & ~new_n949;
  assign new_n15436 = new_n963 & ~new_n15435;
  assign new_n15437 = ~new_n963 & new_n15435;
  assign n10589 = ~new_n15436 & ~new_n15437;
  assign new_n15439 = ~new_n1268 & ~new_n1269_1;
  assign new_n15440 = ~new_n1273 & ~new_n15439;
  assign new_n15441 = new_n1273 & new_n15439;
  assign n10695 = ~new_n15440 & ~new_n15441;
  assign new_n15443 = ~new_n4027 & ~new_n4028;
  assign new_n15444 = ~new_n4162 & ~new_n15443;
  assign new_n15445 = new_n4162 & new_n15443;
  assign n10789 = ~new_n15444 & ~new_n15445;
  assign new_n15447 = ~new_n3307 & ~new_n3309;
  assign n10851 = ~new_n3310 & ~new_n15447;
  assign new_n15449 = ~new_n5655 & ~new_n5656;
  assign new_n15450 = new_n5670_1 & ~new_n15449;
  assign new_n15451 = ~new_n5670_1 & new_n15449;
  assign n10913 = ~new_n15450 & ~new_n15451;
  assign new_n15453 = ~new_n8001 & ~new_n8002;
  assign new_n15454 = ~new_n8161 & new_n15453;
  assign new_n15455 = new_n8161 & ~new_n15453;
  assign n10949 = ~new_n15454 & ~new_n15455;
  assign new_n15457 = ~new_n13091 & ~new_n13092;
  assign new_n15458 = new_n13146 & ~new_n15457;
  assign new_n15459 = ~new_n13146 & new_n15457;
  assign n11216 = new_n15458 | new_n15459;
  assign new_n15461 = ~new_n5657 & ~new_n5659;
  assign n11326 = ~new_n5660 & ~new_n15461;
  assign new_n15463 = ~new_n6303 & new_n6465;
  assign new_n15464 = ~new_n6302 & ~new_n15463;
  assign new_n15465 = ~new_n6355 & new_n6462;
  assign new_n15466 = ~new_n6356 & ~new_n15465;
  assign new_n15467 = n4312 & n9195;
  assign new_n15468 = ~new_n6012 & ~new_n6016_1;
  assign new_n15469 = ~new_n6015 & ~new_n15468;
  assign new_n15470 = new_n15467 & new_n15469;
  assign new_n15471 = ~new_n15467 & ~new_n15469;
  assign new_n15472 = ~new_n15470 & ~new_n15471;
  assign new_n15473 = n1097 & n2253;
  assign new_n15474 = n4634 & n12705;
  assign new_n15475 = n3865 & n5964;
  assign new_n15476 = new_n15474 & ~new_n15475;
  assign new_n15477 = ~new_n15474 & new_n15475;
  assign new_n15478 = ~new_n15476 & ~new_n15477;
  assign new_n15479 = new_n15473 & ~new_n15478;
  assign new_n15480 = ~new_n15473 & new_n15478;
  assign new_n15481 = ~new_n15479 & ~new_n15480;
  assign new_n15482 = ~new_n6009 & new_n6020;
  assign new_n15483 = ~new_n6010 & ~new_n15482;
  assign new_n15484 = new_n15481 & new_n15483;
  assign new_n15485 = ~new_n15481 & ~new_n15483;
  assign new_n15486 = ~new_n15484 & ~new_n15485;
  assign new_n15487 = new_n15472 & ~new_n15486;
  assign new_n15488 = ~new_n15472 & new_n15486;
  assign new_n15489 = ~new_n15487 & ~new_n15488;
  assign new_n15490 = ~new_n6449 & ~new_n6453;
  assign new_n15491 = ~new_n6323 & ~new_n6340;
  assign new_n15492 = ~new_n6322 & ~new_n15491;
  assign new_n15493 = ~new_n6326 & new_n6337;
  assign new_n15494 = ~new_n6327 & ~new_n15493;
  assign new_n15495 = n9189 & n9241;
  assign new_n15496 = n2522 & n8276;
  assign new_n15497 = ~new_n15495 & new_n15496;
  assign new_n15498 = new_n15495 & ~new_n15496;
  assign new_n15499 = ~new_n15497 & ~new_n15498;
  assign new_n15500 = n12221 & n12299;
  assign new_n15501 = n6776 & n10217;
  assign new_n15502 = new_n15500 & ~new_n15501;
  assign new_n15503 = ~new_n15500 & new_n15501;
  assign new_n15504 = ~new_n15502 & ~new_n15503;
  assign new_n15505 = ~new_n15499 & ~new_n15504;
  assign new_n15506 = new_n15499 & new_n15504;
  assign new_n15507 = ~new_n15505 & ~new_n15506;
  assign new_n15508 = n7436 & n12145;
  assign new_n15509 = ~new_n6329 & ~new_n6333;
  assign new_n15510 = ~new_n6332 & ~new_n15509;
  assign new_n15511 = new_n15508 & new_n15510;
  assign new_n15512 = ~new_n15508 & ~new_n15510;
  assign new_n15513 = ~new_n15511 & ~new_n15512;
  assign new_n15514 = new_n15507 & ~new_n15513;
  assign new_n15515 = ~new_n15507 & new_n15513;
  assign new_n15516 = ~new_n15514 & ~new_n15515;
  assign new_n15517 = ~new_n15494 & new_n15516;
  assign new_n15518 = new_n15494 & ~new_n15516;
  assign new_n15519 = ~new_n15517 & ~new_n15518;
  assign new_n15520 = new_n15492 & new_n15519;
  assign new_n15521 = ~new_n15492 & ~new_n15519;
  assign new_n15522 = ~new_n15520 & ~new_n15521;
  assign new_n15523 = ~new_n6311 & ~new_n6315;
  assign new_n15524 = ~new_n6314 & ~new_n15523;
  assign new_n15525 = ~new_n15522 & new_n15524;
  assign new_n15526 = new_n15522 & ~new_n15524;
  assign new_n15527 = ~new_n15525 & ~new_n15526;
  assign new_n15528 = ~new_n6409 & ~new_n6444;
  assign new_n15529 = ~new_n6410 & ~new_n15528;
  assign new_n15530 = n3342 & n3986;
  assign new_n15531 = n5857 & n9111;
  assign new_n15532 = ~new_n15530 & ~new_n15531;
  assign new_n15533 = new_n15530 & new_n15531;
  assign new_n15534 = ~new_n15532 & ~new_n15533;
  assign new_n15535 = n6431 & n7965;
  assign new_n15536 = n45 & n9763;
  assign new_n15537 = new_n15535 & ~new_n15536;
  assign new_n15538 = ~new_n15535 & new_n15536;
  assign new_n15539 = ~new_n15537 & ~new_n15538;
  assign new_n15540 = ~new_n15534 & ~new_n15539;
  assign new_n15541 = new_n15534 & new_n15539;
  assign new_n15542 = ~new_n15540 & ~new_n15541;
  assign new_n15543 = ~new_n15529 & new_n15542;
  assign new_n15544 = new_n15529 & ~new_n15542;
  assign new_n15545 = ~new_n15543 & ~new_n15544;
  assign new_n15546 = new_n15527 & ~new_n15545;
  assign new_n15547 = ~new_n15527 & new_n15545;
  assign new_n15548 = ~new_n15546 & ~new_n15547;
  assign new_n15549 = new_n15490 & ~new_n15548;
  assign new_n15550 = ~new_n15490 & new_n15548;
  assign new_n15551 = ~new_n15549 & ~new_n15550;
  assign new_n15552 = ~new_n15489 & new_n15551;
  assign new_n15553 = new_n15489 & ~new_n15551;
  assign new_n15554 = ~new_n15552 & ~new_n15553;
  assign new_n15555 = new_n6460 & new_n15554;
  assign new_n15556 = ~new_n6460 & ~new_n15554;
  assign new_n15557 = ~new_n15555 & ~new_n15556;
  assign new_n15558 = ~new_n6401 & ~new_n6405;
  assign new_n15559 = ~new_n6424 & ~new_n6441_1;
  assign new_n15560 = ~new_n6423 & ~new_n15559;
  assign new_n15561 = ~new_n6427 & ~new_n6438;
  assign new_n15562 = ~new_n6428 & ~new_n15561;
  assign new_n15563 = n2507 & n7388;
  assign new_n15564 = n2393 & n7270;
  assign new_n15565 = n806 & n5860;
  assign new_n15566 = ~new_n15564 & new_n15565;
  assign new_n15567 = new_n15564 & ~new_n15565;
  assign new_n15568 = ~new_n15566 & ~new_n15567;
  assign new_n15569 = new_n15563 & new_n15568;
  assign new_n15570 = ~new_n15563 & ~new_n15568;
  assign new_n15571 = ~new_n15569 & ~new_n15570;
  assign new_n15572 = ~new_n6412 & ~new_n6416;
  assign new_n15573 = ~new_n6415 & ~new_n15572;
  assign new_n15574 = ~new_n15571 & new_n15573;
  assign new_n15575 = new_n15571 & ~new_n15573;
  assign new_n15576 = ~new_n15574 & ~new_n15575;
  assign new_n15577 = new_n15562 & ~new_n15576;
  assign new_n15578 = ~new_n15562 & new_n15576;
  assign new_n15579 = ~new_n15577 & ~new_n15578;
  assign new_n15580 = new_n15560 & new_n15579;
  assign new_n15581 = ~new_n15560 & ~new_n15579;
  assign new_n15582 = ~new_n15580 & ~new_n15581;
  assign new_n15583 = n6016 & n12648;
  assign new_n15584 = n521 & n10545;
  assign new_n15585 = ~new_n15583 & ~new_n15584;
  assign new_n15586 = new_n15583 & new_n15584;
  assign new_n15587 = ~new_n15585 & ~new_n15586;
  assign new_n15588 = n5579 & n7690;
  assign new_n15589 = n2498 & n3616;
  assign new_n15590 = new_n15588 & ~new_n15589;
  assign new_n15591 = ~new_n15588 & new_n15589;
  assign new_n15592 = ~new_n15590 & ~new_n15591;
  assign new_n15593 = ~new_n15587 & ~new_n15592;
  assign new_n15594 = new_n15587 & new_n15592;
  assign new_n15595 = ~new_n15593 & ~new_n15594;
  assign new_n15596 = ~new_n6430 & ~new_n6434;
  assign new_n15597 = ~new_n6433 & ~new_n15596;
  assign new_n15598 = n1576 & n5331;
  assign new_n15599 = n5153 & n11892;
  assign new_n15600 = new_n15598 & ~new_n15599;
  assign new_n15601 = ~new_n15598 & new_n15599;
  assign new_n15602 = ~new_n15600 & ~new_n15601;
  assign new_n15603 = ~new_n15597 & new_n15602;
  assign new_n15604 = new_n15597 & ~new_n15602;
  assign new_n15605 = ~new_n15603 & ~new_n15604;
  assign new_n15606 = ~new_n15595 & new_n15605;
  assign new_n15607 = new_n15595 & ~new_n15605;
  assign new_n15608 = ~new_n15606 & ~new_n15607;
  assign new_n15609 = ~new_n15582 & new_n15608;
  assign new_n15610 = new_n15582 & ~new_n15608;
  assign new_n15611 = ~new_n15609 & ~new_n15610;
  assign new_n15612 = n2558 & n4499;
  assign new_n15613 = ~new_n6360 & ~new_n6396;
  assign new_n15614 = ~new_n6361 & ~new_n15613;
  assign new_n15615 = new_n15612 & new_n15614;
  assign new_n15616 = ~new_n15612 & ~new_n15614;
  assign new_n15617 = ~new_n15615 & ~new_n15616;
  assign new_n15618 = new_n15611 & new_n15617;
  assign new_n15619 = ~new_n15611 & ~new_n15617;
  assign new_n15620 = ~new_n15618 & ~new_n15619;
  assign new_n15621 = ~new_n15558 & ~new_n15620;
  assign new_n15622 = new_n15558 & new_n15620;
  assign new_n15623 = ~new_n15621 & ~new_n15622;
  assign new_n15624 = ~new_n6348 & ~new_n6350;
  assign new_n15625 = ~new_n6308 & new_n6343;
  assign new_n15626 = ~new_n6309 & ~new_n15625;
  assign new_n15627 = ~new_n5994 & ~new_n5998;
  assign new_n15628 = ~new_n5997 & ~new_n15627;
  assign new_n15629 = ~new_n6005 & new_n6023;
  assign new_n15630 = ~new_n6006 & ~new_n15629;
  assign new_n15631 = ~new_n15628 & ~new_n15630;
  assign new_n15632 = new_n15628 & new_n15630;
  assign new_n15633 = ~new_n15631 & ~new_n15632;
  assign new_n15634 = n7946 & n10644;
  assign new_n15635 = n7823 & n8759;
  assign new_n15636 = n2024 & n10510;
  assign new_n15637 = ~new_n15635 & new_n15636;
  assign new_n15638 = new_n15635 & ~new_n15636;
  assign new_n15639 = ~new_n15637 & ~new_n15638;
  assign new_n15640 = new_n15634 & ~new_n15639;
  assign new_n15641 = ~new_n15634 & new_n15639;
  assign new_n15642 = ~new_n15640 & ~new_n15641;
  assign new_n15643 = ~new_n15633 & new_n15642;
  assign new_n15644 = new_n15633 & ~new_n15642;
  assign new_n15645 = ~new_n15643 & ~new_n15644;
  assign new_n15646 = ~new_n15626 & ~new_n15645;
  assign new_n15647 = new_n15626 & new_n15645;
  assign new_n15648 = ~new_n15646 & ~new_n15647;
  assign new_n15649 = n10223 & n12025;
  assign new_n15650 = n2879 & n11257;
  assign new_n15651 = new_n15649 & ~new_n15650;
  assign new_n15652 = ~new_n15649 & new_n15650;
  assign new_n15653 = ~new_n15651 & ~new_n15652;
  assign new_n15654 = ~new_n15648 & new_n15653;
  assign new_n15655 = new_n15648 & ~new_n15653;
  assign new_n15656 = ~new_n15654 & ~new_n15655;
  assign new_n15657 = new_n15624 & ~new_n15656;
  assign new_n15658 = ~new_n15624 & new_n15656;
  assign new_n15659 = ~new_n15657 & ~new_n15658;
  assign new_n15660 = new_n15623 & new_n15659;
  assign new_n15661 = ~new_n15623 & ~new_n15659;
  assign new_n15662 = ~new_n15660 & ~new_n15661;
  assign new_n15663 = new_n15557 & ~new_n15662;
  assign new_n15664 = ~new_n15557 & new_n15662;
  assign new_n15665 = ~new_n15663 & ~new_n15664;
  assign new_n15666 = ~new_n15466 & ~new_n15665;
  assign new_n15667 = new_n15466 & new_n15665;
  assign new_n15668 = ~new_n15666 & ~new_n15667;
  assign new_n15669 = ~new_n6032 & ~new_n6048;
  assign new_n15670 = ~new_n6374 & ~new_n6393;
  assign new_n15671 = ~new_n6375 & ~new_n15670;
  assign new_n15672 = ~new_n6379 & ~new_n6391;
  assign new_n15673 = ~new_n6381 & ~new_n6385;
  assign new_n15674 = ~new_n6384 & ~new_n15673;
  assign new_n15675 = n2347 & n8476;
  assign new_n15676 = n2530 & n5798;
  assign new_n15677 = new_n15675 & ~new_n15676;
  assign new_n15678 = ~new_n15675 & new_n15676;
  assign new_n15679 = ~new_n15677 & ~new_n15678;
  assign new_n15680 = ~new_n15674 & new_n15679;
  assign new_n15681 = new_n15674 & ~new_n15679;
  assign new_n15682 = ~new_n15680 & ~new_n15681;
  assign new_n15683 = new_n15672 & new_n15682;
  assign new_n15684 = ~new_n15672 & ~new_n15682;
  assign new_n15685 = ~new_n15683 & ~new_n15684;
  assign new_n15686 = ~new_n6363 & ~new_n6367;
  assign new_n15687 = ~new_n6366 & ~new_n15686;
  assign new_n15688 = new_n15685 & ~new_n15687;
  assign new_n15689 = ~new_n15685 & new_n15687;
  assign new_n15690 = ~new_n15688 & ~new_n15689;
  assign new_n15691 = ~new_n15671 & ~new_n15690;
  assign new_n15692 = new_n15671 & new_n15690;
  assign new_n15693 = ~new_n15691 & ~new_n15692;
  assign new_n15694 = ~new_n5991 & ~new_n6028;
  assign new_n15695 = n7265 & n10547;
  assign new_n15696 = n2512 & n5305;
  assign new_n15697 = ~new_n15695 & new_n15696;
  assign new_n15698 = new_n15695 & ~new_n15696;
  assign new_n15699 = ~new_n15697 & ~new_n15698;
  assign new_n15700 = ~new_n15694 & ~new_n15699;
  assign new_n15701 = new_n15694 & new_n15699;
  assign new_n15702 = ~new_n15700 & ~new_n15701;
  assign new_n15703 = ~new_n15693 & new_n15702;
  assign new_n15704 = new_n15693 & ~new_n15702;
  assign new_n15705 = ~new_n15703 & ~new_n15704;
  assign new_n15706 = new_n15669 & new_n15705;
  assign new_n15707 = ~new_n15669 & ~new_n15705;
  assign new_n15708 = ~new_n15706 & ~new_n15707;
  assign new_n15709 = ~new_n15668 & new_n15708;
  assign new_n15710 = new_n15668 & ~new_n15708;
  assign new_n15711 = ~new_n15709 & ~new_n15710;
  assign new_n15712 = ~new_n15464 & ~new_n15711;
  assign new_n15713 = new_n15464 & new_n15711;
  assign n11707 = ~new_n15712 & ~new_n15713;
  assign new_n15715 = ~new_n7030 & ~new_n7031;
  assign new_n15716 = ~new_n7035 & ~new_n15715;
  assign new_n15717 = new_n7035 & new_n15715;
  assign n11755 = ~new_n15716 & ~new_n15717;
  assign new_n15719 = ~new_n3996 & ~new_n3997;
  assign new_n15720 = new_n4022 & ~new_n15719;
  assign new_n15721 = ~new_n4022 & new_n15719;
  assign n11780 = ~new_n15720 & ~new_n15721;
  assign new_n15723 = ~new_n11584 & ~new_n11585;
  assign new_n15724 = new_n11587 & new_n15723;
  assign new_n15725 = ~new_n11587 & ~new_n15723;
  assign n11919 = new_n15724 | new_n15725;
  assign new_n15727 = ~new_n11574 & ~new_n11575;
  assign new_n15728 = new_n11589 & ~new_n15727;
  assign new_n15729 = ~new_n11589 & new_n15727;
  assign n12005 = new_n15728 | new_n15729;
  assign new_n15731 = ~new_n12241 & ~new_n12242;
  assign new_n15732 = new_n12244 & ~new_n15731;
  assign new_n15733 = ~new_n12244 & new_n15731;
  assign n12014 = ~new_n15732 & ~new_n15733;
  assign new_n15735 = new_n9995 & ~new_n10027;
  assign new_n15736 = new_n10029 & ~new_n15735;
  assign new_n15737 = new_n9994 & new_n10027;
  assign n12020 = new_n15736 | new_n15737;
  assign new_n15739 = ~new_n13101 & ~new_n13102;
  assign new_n15740 = new_n13136 & new_n15739;
  assign new_n15741 = ~new_n13136 & ~new_n15739;
  assign n12076 = new_n15740 | new_n15741;
  assign new_n15743 = ~new_n13821 & ~new_n13822;
  assign new_n15744 = new_n13826 & new_n15743;
  assign new_n15745 = ~new_n13826 & ~new_n15743;
  assign n12111 = new_n15744 | new_n15745;
  assign new_n15747 = ~new_n12233 & ~new_n12234;
  assign new_n15748 = new_n12246 & ~new_n15747;
  assign new_n15749 = ~new_n12246 & new_n15747;
  assign n12444 = ~new_n15748 & ~new_n15749;
  assign new_n15751 = ~new_n6286 & ~new_n6287;
  assign new_n15752 = ~new_n6299 & ~new_n15751;
  assign new_n15753 = new_n6299 & new_n15751;
  assign n12807 = ~new_n15752 & ~new_n15753;
endmodule


