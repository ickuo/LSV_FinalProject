// Benchmark "top" written by ABC on Sun Dec 21 18:08:13 2025

module top ( 
    n2, n11, n13, n16, n21, n45, n46, n55, n74, n75, n81, n84, n85, n93,
    n96, n98, n101, n111, n128, n131, n134, n139, n153, n159, n177, n199,
    n206, n211, n216, n223, n243, n264, n266, n280, n282, n287, n290, n309,
    n336, n346, n349, n360, n368, n369, n377, n388, n394, n409, n428, n435,
    n447, n454, n457, n468, n471, n481, n494, n500, n507, n511, n519, n525,
    n557, n561, n569, n571, n575, n581, n582, n583, n587, n600, n603, n609,
    n613, n614, n616, n646, n659, n661, n664, n673,
    n44, n87, n105, n123, n148, n163, n191, n196, n226, n240, n254, n260,
    n283, n291, n299, n442, n449, n484, n518, n534, n542, n547, n568, n627,
    n635, n672  );
  input  n2, n11, n13, n16, n21, n45, n46, n55, n74, n75, n81, n84, n85,
    n93, n96, n98, n101, n111, n128, n131, n134, n139, n153, n159, n177,
    n199, n206, n211, n216, n223, n243, n264, n266, n280, n282, n287, n290,
    n309, n336, n346, n349, n360, n368, n369, n377, n388, n394, n409, n428,
    n435, n447, n454, n457, n468, n471, n481, n494, n500, n507, n511, n519,
    n525, n557, n561, n569, n571, n575, n581, n582, n583, n587, n600, n603,
    n609, n613, n614, n616, n646, n659, n661, n664, n673;
  output n44, n87, n105, n123, n148, n163, n191, n196, n226, n240, n254, n260,
    n283, n291, n299, n442, n449, n484, n518, n534, n542, n547, n568, n627,
    n635, n672;
  wire new_n109, new_n110, new_n111_1, new_n112, new_n113, new_n114,
    new_n115, new_n116, new_n117, new_n118, new_n119, new_n120, new_n121,
    new_n122, new_n123_1, new_n124, new_n125, new_n126, new_n127,
    new_n128_1, new_n129, new_n130, new_n131_1, new_n132, new_n133,
    new_n134_1, new_n135, new_n136, new_n137, new_n138, new_n139_1,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148_1, new_n149, new_n150, new_n151, new_n152,
    new_n153_1, new_n154, new_n155, new_n156, new_n157, new_n158,
    new_n159_1, new_n160, new_n161, new_n162, new_n163_1, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177_1, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191_1, new_n192,
    new_n193, new_n194, new_n195, new_n196_1, new_n197, new_n198,
    new_n199_1, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206_1, new_n207, new_n208, new_n209, new_n210, new_n211_1,
    new_n212, new_n213, new_n214, new_n215, new_n216_1, new_n217, new_n218,
    new_n219, new_n220, new_n221, new_n222, new_n223_1, new_n224, new_n225,
    new_n226_1, new_n227, new_n228, new_n229, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240_1, new_n241, new_n242, new_n243_1, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254_1, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260_1, new_n261, new_n262, new_n263, new_n264_1, new_n265,
    new_n266_1, new_n267, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280_1, new_n281, new_n282_1, new_n283_1, new_n284, new_n285,
    new_n286, new_n287_1, new_n288, new_n289, new_n290_1, new_n291_1,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299_1, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309_1, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336_1, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346_1, new_n347,
    new_n348, new_n349_1, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360_1, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368_1,
    new_n369_1, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377_1, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388_1, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394_1, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409_1, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428_1, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435_1, new_n436, new_n438, new_n439,
    new_n440, new_n442_1, new_n443, new_n444, new_n446, new_n447_1,
    new_n448, new_n449_1, new_n450, new_n451, new_n452, new_n453,
    new_n454_1, new_n455, new_n456, new_n457_1, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468_1, new_n469, new_n470, new_n471_1, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481_1, new_n482, new_n483, new_n484_1, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494_1, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500_1, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507_1, new_n508, new_n509, new_n510, new_n511_1, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518_1,
    new_n519_1, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525_1, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534_1, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542_1, new_n543, new_n544, new_n546,
    new_n547_1, new_n548, new_n549, new_n550, new_n551, new_n553, new_n554,
    new_n555, new_n557_1, new_n558, new_n559, new_n561_1, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568_1, new_n569_1,
    new_n570, new_n571_1, new_n572, new_n573, new_n575_1, new_n576,
    new_n577, new_n579, new_n580, new_n581_1, new_n583_1, new_n584,
    new_n585, new_n587_1, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600_1, new_n602,
    new_n603_1, new_n604, new_n606, new_n608, new_n609_1, new_n610,
    new_n612, new_n613_1, new_n614_1, new_n616_1, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627_1,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635_1,
    new_n636, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n646_1, new_n647, new_n648;
  assign new_n109 = ~n206 & ~n368;
  assign new_n110 = ~n85 & ~n349;
  assign new_n111_1 = ~n93 & new_n110;
  assign new_n112 = new_n109 & new_n111_1;
  assign new_n113 = n98 & new_n112;
  assign new_n114 = n409 & n468;
  assign new_n115 = n409 & n428;
  assign new_n116 = ~n468 & ~new_n115;
  assign new_n117 = ~new_n114 & ~new_n116;
  assign new_n118 = ~n616 & ~new_n117;
  assign new_n119 = n409 & ~n428;
  assign new_n120 = n468 & ~new_n119;
  assign new_n121 = ~n468 & new_n119;
  assign new_n122 = ~new_n120 & ~new_n121;
  assign new_n123_1 = ~n616 & ~new_n122;
  assign new_n124 = n616 & new_n122;
  assign new_n125 = ~n409 & ~n428;
  assign new_n126 = ~new_n115 & ~new_n125;
  assign new_n127 = ~n216 & ~new_n126;
  assign new_n128_1 = n216 & new_n126;
  assign new_n129 = n428 & n454;
  assign new_n130 = ~new_n128_1 & ~new_n129;
  assign new_n131_1 = ~new_n127 & ~new_n130;
  assign new_n132 = ~new_n124 & new_n131_1;
  assign new_n133 = ~new_n123_1 & ~new_n132;
  assign new_n134_1 = ~new_n118 & ~new_n133;
  assign new_n135 = new_n114 & new_n134_1;
  assign new_n136 = n93 & new_n135;
  assign new_n137 = ~new_n113 & ~new_n136;
  assign new_n138 = ~n266 & ~n519;
  assign new_n139_1 = ~n454 & ~n659;
  assign new_n140 = ~n216 & ~n616;
  assign new_n141 = new_n139_1 & new_n140;
  assign new_n142 = n511 & ~new_n141;
  assign new_n143 = n16 & new_n142;
  assign new_n144 = ~n45 & ~new_n143;
  assign new_n145 = n45 & new_n143;
  assign new_n146 = ~new_n144 & ~new_n145;
  assign new_n147 = n266 & ~new_n146;
  assign new_n148_1 = ~new_n138 & ~new_n147;
  assign new_n149 = ~new_n137 & ~new_n148_1;
  assign new_n150 = ~n266 & n377;
  assign new_n151 = n266 & ~new_n143;
  assign new_n152 = n511 & new_n151;
  assign new_n153_1 = ~new_n150 & ~new_n152;
  assign new_n154 = n21 & new_n112;
  assign new_n155 = n616 & new_n117;
  assign new_n156 = ~new_n114 & ~new_n134_1;
  assign new_n157 = ~new_n155 & new_n156;
  assign new_n158 = n93 & ~new_n135;
  assign new_n159_1 = ~new_n157 & new_n158;
  assign new_n160 = ~new_n154 & ~new_n159_1;
  assign new_n161 = ~new_n153_1 & new_n160;
  assign new_n162 = new_n153_1 & ~new_n160;
  assign new_n163_1 = n81 & ~n266;
  assign new_n164 = ~n16 & ~new_n142;
  assign new_n165 = new_n151 & ~new_n164;
  assign new_n166 = ~new_n163_1 & ~new_n165;
  assign new_n167 = n264 & new_n112;
  assign new_n168 = n454 & n659;
  assign new_n169 = n216 & new_n168;
  assign new_n170 = n616 & new_n169;
  assign new_n171 = ~n93 & n206;
  assign new_n172 = new_n170 & new_n171;
  assign new_n173 = ~new_n167 & ~new_n172;
  assign new_n174 = ~new_n118 & ~new_n155;
  assign new_n175 = new_n133 & ~new_n174;
  assign new_n176 = new_n134_1 & ~new_n155;
  assign new_n177_1 = n93 & ~new_n176;
  assign new_n178 = ~new_n175 & new_n177_1;
  assign new_n179 = new_n173 & ~new_n178;
  assign new_n180 = ~new_n166 & new_n179;
  assign new_n181 = ~n616 & ~new_n169;
  assign new_n182 = ~new_n170 & ~new_n181;
  assign new_n183 = n206 & new_n182;
  assign new_n184 = n75 & n435;
  assign new_n185 = ~n75 & ~n435;
  assign new_n186 = ~n2 & ~n582;
  assign new_n187 = n2 & n582;
  assign new_n188 = n287 & n600;
  assign new_n189 = ~new_n187 & ~new_n188;
  assign new_n190 = ~new_n186 & ~new_n189;
  assign new_n191_1 = ~new_n185 & new_n190;
  assign new_n192 = n349 & ~new_n191_1;
  assign new_n193 = ~new_n184 & new_n192;
  assign new_n194 = ~n85 & n199;
  assign new_n195 = ~n349 & ~new_n194;
  assign new_n196_1 = n75 & n177;
  assign new_n197 = ~n2 & ~n13;
  assign new_n198 = n2 & n13;
  assign new_n199_1 = n280 & n287;
  assign new_n200 = ~new_n198 & ~new_n199_1;
  assign new_n201 = ~new_n197 & ~new_n200;
  assign new_n202 = ~new_n196_1 & ~new_n201;
  assign new_n203 = ~n75 & ~n177;
  assign new_n204 = n85 & ~new_n203;
  assign new_n205 = ~new_n202 & new_n204;
  assign new_n206_1 = new_n195 & ~new_n205;
  assign new_n207 = new_n109 & ~new_n206_1;
  assign new_n208 = ~new_n193 & new_n207;
  assign new_n209 = ~new_n183 & ~new_n208;
  assign new_n210 = n75 & n131;
  assign new_n211_1 = ~n2 & ~n159;
  assign new_n212 = n2 & n159;
  assign new_n213 = n96 & n287;
  assign new_n214 = ~new_n212 & ~new_n213;
  assign new_n215 = ~new_n211_1 & ~new_n214;
  assign new_n216_1 = ~new_n210 & ~new_n215;
  assign new_n217 = ~n75 & ~n131;
  assign new_n218 = ~n206 & n368;
  assign new_n219 = ~new_n217 & new_n218;
  assign new_n220 = ~new_n216_1 & new_n219;
  assign new_n221 = ~n93 & ~new_n220;
  assign new_n222 = new_n209 & new_n221;
  assign new_n223_1 = ~new_n123_1 & ~new_n124;
  assign new_n224 = new_n131_1 & new_n223_1;
  assign new_n225 = ~new_n131_1 & ~new_n223_1;
  assign new_n226_1 = ~new_n224 & ~new_n225;
  assign new_n227 = n93 & ~new_n226_1;
  assign new_n228 = ~new_n222 & ~new_n227;
  assign new_n229 = ~n266 & ~n507;
  assign new_n230 = n511 & new_n139_1;
  assign new_n231 = ~n216 & new_n230;
  assign new_n232 = n616 & new_n231;
  assign new_n233 = ~n616 & ~new_n231;
  assign new_n234 = ~new_n232 & ~new_n233;
  assign new_n235 = n266 & ~new_n234;
  assign new_n236 = ~new_n229 & ~new_n235;
  assign new_n237 = ~new_n228 & new_n236;
  assign new_n238 = new_n228 & ~new_n236;
  assign new_n239 = n85 & ~n349;
  assign new_n240_1 = ~new_n196_1 & ~new_n203;
  assign new_n241 = new_n201 & new_n240_1;
  assign new_n242 = ~new_n201 & ~new_n240_1;
  assign new_n243_1 = ~new_n241 & ~new_n242;
  assign new_n244 = new_n239 & new_n243_1;
  assign new_n245 = n211 & new_n110;
  assign new_n246 = ~new_n184 & ~new_n185;
  assign new_n247 = new_n190 & new_n246;
  assign new_n248 = ~new_n190 & ~new_n246;
  assign new_n249 = n349 & ~new_n248;
  assign new_n250 = ~new_n247 & new_n249;
  assign new_n251 = ~new_n245 & ~new_n250;
  assign new_n252 = ~new_n244 & new_n251;
  assign new_n253 = new_n109 & ~new_n252;
  assign new_n254_1 = ~n216 & ~new_n168;
  assign new_n255 = ~new_n169 & ~new_n254_1;
  assign new_n256 = n206 & new_n255;
  assign new_n257 = ~new_n253 & ~new_n256;
  assign new_n258 = ~new_n210 & ~new_n217;
  assign new_n259 = new_n215 & new_n258;
  assign new_n260_1 = ~new_n215 & ~new_n258;
  assign new_n261 = ~new_n259 & ~new_n260_1;
  assign new_n262 = new_n218 & new_n261;
  assign new_n263 = ~n93 & ~new_n262;
  assign new_n264_1 = new_n257 & new_n263;
  assign new_n265 = ~new_n127 & ~new_n128_1;
  assign new_n266_1 = new_n129 & new_n265;
  assign new_n267 = ~new_n129 & ~new_n265;
  assign new_n268 = ~new_n266_1 & ~new_n267;
  assign new_n269 = n93 & ~new_n268;
  assign new_n270 = ~new_n264_1 & ~new_n269;
  assign new_n271 = ~n266 & ~n457;
  assign new_n272 = n216 & ~new_n230;
  assign new_n273 = ~new_n231 & ~new_n272;
  assign new_n274 = n266 & new_n273;
  assign new_n275 = ~new_n271 & ~new_n274;
  assign new_n276 = new_n270 & ~new_n275;
  assign new_n277 = ~new_n270 & new_n275;
  assign new_n278 = ~n428 & ~n454;
  assign new_n279 = ~new_n129 & ~new_n278;
  assign new_n280_1 = n93 & ~new_n279;
  assign new_n281 = ~new_n186 & ~new_n187;
  assign new_n282_1 = new_n188 & ~new_n281;
  assign new_n283_1 = ~new_n188 & new_n281;
  assign new_n284 = ~new_n282_1 & ~new_n283_1;
  assign new_n285 = n349 & ~new_n284;
  assign new_n286 = ~new_n197 & ~new_n198;
  assign new_n287_1 = new_n199_1 & new_n286;
  assign new_n288 = ~new_n199_1 & ~new_n286;
  assign new_n289 = ~new_n287_1 & ~new_n288;
  assign new_n290_1 = new_n239 & new_n289;
  assign new_n291_1 = n525 & new_n110;
  assign new_n292 = ~new_n290_1 & ~new_n291_1;
  assign new_n293 = ~new_n285 & new_n292;
  assign new_n294 = new_n109 & ~new_n293;
  assign new_n295 = ~new_n211_1 & ~new_n212;
  assign new_n296 = new_n213 & new_n295;
  assign new_n297 = ~new_n213 & ~new_n295;
  assign new_n298 = ~new_n296 & ~new_n297;
  assign new_n299_1 = new_n218 & new_n298;
  assign new_n300 = n206 & ~new_n168;
  assign new_n301 = ~new_n139_1 & new_n300;
  assign new_n302 = ~new_n299_1 & ~new_n301;
  assign new_n303 = ~new_n294 & new_n302;
  assign new_n304 = ~n93 & new_n303;
  assign new_n305 = ~new_n280_1 & ~new_n304;
  assign new_n306 = n93 & ~n659;
  assign new_n307 = ~n280 & ~n287;
  assign new_n308 = ~new_n199_1 & new_n239;
  assign new_n309_1 = ~new_n307 & new_n308;
  assign new_n310 = n664 & new_n110;
  assign new_n311 = ~n287 & ~n600;
  assign new_n312 = n349 & ~new_n188;
  assign new_n313 = ~new_n311 & new_n312;
  assign new_n314 = ~new_n310 & ~new_n313;
  assign new_n315 = ~new_n309_1 & new_n314;
  assign new_n316 = new_n109 & ~new_n315;
  assign new_n317 = n206 & ~n659;
  assign new_n318 = ~n96 & ~n287;
  assign new_n319 = ~new_n213 & ~new_n318;
  assign new_n320 = new_n218 & new_n319;
  assign new_n321 = ~new_n317 & ~new_n320;
  assign new_n322 = ~new_n316 & new_n321;
  assign new_n323 = ~n93 & new_n322;
  assign new_n324 = ~new_n306 & ~new_n323;
  assign new_n325 = n511 & ~n659;
  assign new_n326 = ~n511 & n659;
  assign new_n327 = ~new_n325 & ~new_n326;
  assign new_n328 = n266 & ~new_n327;
  assign new_n329 = ~n266 & n673;
  assign new_n330 = ~new_n328 & ~new_n329;
  assign new_n331 = new_n324 & new_n330;
  assign new_n332 = n454 & ~new_n325;
  assign new_n333 = ~new_n230 & ~new_n332;
  assign new_n334 = n266 & new_n333;
  assign new_n335 = ~n46 & ~n266;
  assign new_n336_1 = ~new_n334 & ~new_n335;
  assign new_n337 = new_n331 & ~new_n336_1;
  assign new_n338 = ~new_n305 & ~new_n337;
  assign new_n339 = ~new_n331 & new_n336_1;
  assign new_n340 = ~new_n338 & ~new_n339;
  assign new_n341 = ~new_n277 & new_n340;
  assign new_n342 = ~new_n276 & ~new_n341;
  assign new_n343 = ~new_n238 & new_n342;
  assign new_n344 = ~new_n237 & ~new_n343;
  assign new_n345 = new_n166 & ~new_n179;
  assign new_n346_1 = ~new_n344 & ~new_n345;
  assign new_n347 = ~new_n180 & ~new_n346_1;
  assign new_n348 = ~new_n162 & ~new_n347;
  assign new_n349_1 = ~new_n161 & ~new_n348;
  assign new_n350 = ~new_n149 & ~new_n349_1;
  assign new_n351 = new_n137 & new_n146;
  assign new_n352 = n266 & ~new_n351;
  assign new_n353 = ~new_n350 & new_n352;
  assign new_n354 = n84 & ~n266;
  assign new_n355 = n111 & new_n145;
  assign new_n356 = ~n111 & ~new_n145;
  assign new_n357 = ~new_n355 & ~new_n356;
  assign new_n358 = n266 & new_n357;
  assign new_n359 = ~new_n354 & ~new_n358;
  assign new_n360_1 = new_n353 & new_n359;
  assign new_n361 = n11 & ~n266;
  assign new_n362 = n282 & new_n355;
  assign new_n363 = ~n282 & ~new_n355;
  assign new_n364 = ~new_n362 & ~new_n363;
  assign new_n365 = n266 & new_n364;
  assign new_n366 = ~new_n361 & ~new_n365;
  assign new_n367 = new_n360_1 & new_n366;
  assign new_n368_1 = n646 & new_n362;
  assign new_n369_1 = ~n646 & ~new_n362;
  assign new_n370 = ~new_n368_1 & ~new_n369_1;
  assign new_n371 = n266 & ~new_n370;
  assign new_n372 = ~n266 & ~n571;
  assign new_n373 = ~new_n371 & ~new_n372;
  assign new_n374 = new_n367 & ~new_n373;
  assign new_n375 = n243 & new_n368_1;
  assign new_n376 = ~n243 & ~new_n368_1;
  assign new_n377_1 = ~new_n375 & ~new_n376;
  assign new_n378 = n266 & ~new_n377_1;
  assign new_n379 = ~n266 & ~n500;
  assign new_n380 = ~new_n378 & ~new_n379;
  assign new_n381 = new_n374 & ~new_n380;
  assign new_n382 = n557 & new_n375;
  assign new_n383 = ~n557 & ~new_n375;
  assign new_n384 = ~new_n382 & ~new_n383;
  assign new_n385 = n266 & ~new_n384;
  assign new_n386 = ~n139 & ~n266;
  assign new_n387 = ~new_n385 & ~new_n386;
  assign new_n388_1 = new_n381 & ~new_n387;
  assign new_n389 = n561 & new_n382;
  assign new_n390 = ~n561 & ~new_n382;
  assign new_n391 = ~new_n389 & ~new_n390;
  assign new_n392 = n266 & ~new_n391;
  assign new_n393 = ~n266 & ~n346;
  assign new_n394_1 = ~new_n392 & ~new_n393;
  assign new_n395 = new_n388_1 & ~new_n394_1;
  assign new_n396 = new_n137 & ~new_n148_1;
  assign new_n397 = ~new_n137 & new_n148_1;
  assign new_n398 = ~new_n153_1 & ~new_n160;
  assign new_n399 = new_n153_1 & new_n160;
  assign new_n400 = ~new_n166 & ~new_n179;
  assign new_n401 = new_n166 & new_n179;
  assign new_n402 = ~new_n305 & ~new_n336_1;
  assign new_n403 = new_n305 & new_n336_1;
  assign new_n404 = new_n324 & ~new_n330;
  assign new_n405 = ~new_n403 & ~new_n404;
  assign new_n406 = ~new_n402 & ~new_n405;
  assign new_n407 = new_n270 & new_n275;
  assign new_n408 = ~new_n406 & ~new_n407;
  assign new_n409_1 = ~new_n270 & ~new_n275;
  assign new_n410 = ~new_n408 & ~new_n409_1;
  assign new_n411 = new_n228 & new_n236;
  assign new_n412 = ~new_n410 & ~new_n411;
  assign new_n413 = ~new_n228 & ~new_n236;
  assign new_n414 = ~new_n412 & ~new_n413;
  assign new_n415 = ~new_n401 & new_n414;
  assign new_n416 = ~new_n400 & ~new_n415;
  assign new_n417 = ~new_n399 & ~new_n416;
  assign new_n418 = ~new_n398 & ~new_n417;
  assign new_n419 = ~new_n397 & new_n418;
  assign new_n420 = ~n266 & ~new_n419;
  assign new_n421 = ~new_n396 & new_n420;
  assign new_n422 = ~new_n359 & new_n421;
  assign new_n423 = ~new_n366 & new_n422;
  assign new_n424 = new_n373 & new_n423;
  assign new_n425 = new_n380 & new_n424;
  assign new_n426 = new_n387 & new_n425;
  assign new_n427 = new_n394_1 & new_n426;
  assign new_n428_1 = ~new_n395 & ~new_n427;
  assign new_n429 = ~n471 & ~new_n389;
  assign new_n430 = n471 & new_n389;
  assign new_n431 = ~new_n429 & ~new_n430;
  assign new_n432 = n266 & ~new_n431;
  assign new_n433 = ~n266 & ~n614;
  assign new_n434 = ~new_n432 & ~new_n433;
  assign new_n435_1 = new_n428_1 & new_n434;
  assign new_n436 = ~new_n428_1 & ~new_n434;
  assign n44 = new_n435_1 | new_n436;
  assign new_n438 = ~new_n381 & ~new_n425;
  assign new_n439 = new_n387 & new_n438;
  assign new_n440 = ~new_n387 & ~new_n438;
  assign n87 = new_n439 | new_n440;
  assign new_n442_1 = ~new_n353 & ~new_n421;
  assign new_n443 = new_n359 & ~new_n442_1;
  assign new_n444 = ~new_n359 & new_n442_1;
  assign n105 = new_n443 | new_n444;
  assign new_n446 = new_n427 & new_n434;
  assign new_n447_1 = n613 & new_n430;
  assign new_n448 = ~n613 & ~new_n430;
  assign new_n449_1 = ~new_n447_1 & ~new_n448;
  assign new_n450 = n266 & ~new_n449_1;
  assign new_n451 = ~n266 & ~n609;
  assign new_n452 = ~new_n450 & ~new_n451;
  assign new_n453 = new_n446 & new_n452;
  assign new_n454_1 = n583 & new_n447_1;
  assign new_n455 = ~n583 & ~new_n447_1;
  assign new_n456 = ~new_n454_1 & ~new_n455;
  assign new_n457_1 = n266 & ~new_n456;
  assign new_n458 = ~n266 & ~n603;
  assign new_n459 = ~new_n457_1 & ~new_n458;
  assign new_n460 = new_n453 & new_n459;
  assign new_n461 = n55 & new_n454_1;
  assign new_n462 = ~n55 & ~new_n454_1;
  assign new_n463 = ~new_n461 & ~new_n462;
  assign new_n464 = n266 & ~new_n463;
  assign new_n465 = ~n266 & ~n447;
  assign new_n466 = ~new_n464 & ~new_n465;
  assign new_n467 = new_n460 & new_n466;
  assign new_n468_1 = n128 & new_n461;
  assign new_n469 = ~n128 & ~new_n461;
  assign new_n470 = ~new_n468_1 & ~new_n469;
  assign new_n471_1 = n266 & ~new_n470;
  assign new_n472 = ~n266 & ~n394;
  assign new_n473 = ~new_n471_1 & ~new_n472;
  assign new_n474 = new_n467 & new_n473;
  assign new_n475 = n388 & new_n468_1;
  assign new_n476 = ~n388 & ~new_n468_1;
  assign new_n477 = ~new_n475 & ~new_n476;
  assign new_n478 = n266 & ~new_n477;
  assign new_n479 = ~n266 & ~n360;
  assign new_n480 = ~new_n478 & ~new_n479;
  assign new_n481_1 = new_n474 & new_n480;
  assign new_n482 = n661 & new_n475;
  assign new_n483 = ~n661 & ~new_n475;
  assign new_n484_1 = ~new_n482 & ~new_n483;
  assign new_n485 = n266 & ~new_n484_1;
  assign new_n486 = ~n266 & ~n581;
  assign new_n487 = ~new_n485 & ~new_n486;
  assign new_n488 = new_n481_1 & new_n487;
  assign new_n489 = n575 & new_n482;
  assign new_n490 = ~n575 & ~new_n482;
  assign new_n491 = ~new_n489 & ~new_n490;
  assign new_n492 = n266 & ~new_n491;
  assign new_n493 = ~n134 & ~n266;
  assign new_n494_1 = ~new_n492 & ~new_n493;
  assign new_n495 = new_n488 & new_n494_1;
  assign new_n496 = n369 & new_n489;
  assign new_n497 = ~n369 & ~new_n489;
  assign new_n498 = ~new_n496 & ~new_n497;
  assign new_n499 = n266 & ~new_n498;
  assign new_n500_1 = ~n101 & ~n266;
  assign new_n501 = ~new_n499 & ~new_n500_1;
  assign new_n502 = new_n495 & new_n501;
  assign new_n503 = n336 & new_n496;
  assign new_n504 = ~n336 & ~new_n496;
  assign new_n505 = ~new_n503 & ~new_n504;
  assign new_n506 = n266 & ~new_n505;
  assign new_n507_1 = ~n266 & ~n569;
  assign new_n508 = ~new_n506 & ~new_n507_1;
  assign new_n509 = new_n502 & new_n508;
  assign new_n510 = n494 & new_n503;
  assign new_n511_1 = ~n494 & ~new_n503;
  assign new_n512 = ~new_n510 & ~new_n511_1;
  assign new_n513 = n266 & ~new_n512;
  assign new_n514 = ~n153 & ~n266;
  assign new_n515 = ~new_n513 & ~new_n514;
  assign new_n516 = new_n509 & new_n515;
  assign new_n517 = n223 & new_n510;
  assign new_n518_1 = ~n223 & ~new_n510;
  assign new_n519_1 = ~new_n517 & ~new_n518_1;
  assign new_n520 = n266 & ~new_n519_1;
  assign new_n521 = ~n266 & ~n309;
  assign new_n522 = ~new_n520 & ~new_n521;
  assign new_n523 = ~new_n516 & new_n522;
  assign new_n524 = new_n395 & ~new_n434;
  assign new_n525_1 = ~new_n452 & new_n524;
  assign new_n526 = ~new_n459 & new_n525_1;
  assign new_n527 = ~new_n466 & new_n526;
  assign new_n528 = ~new_n473 & new_n527;
  assign new_n529 = ~new_n480 & new_n528;
  assign new_n530 = ~new_n487 & new_n529;
  assign new_n531 = ~new_n494_1 & new_n530;
  assign new_n532 = ~new_n501 & new_n531;
  assign new_n533 = ~new_n508 & new_n532;
  assign new_n534_1 = ~new_n515 & new_n533;
  assign new_n535 = ~new_n522 & ~new_n534_1;
  assign new_n536 = ~new_n523 & ~new_n535;
  assign new_n537 = n290 & ~new_n517;
  assign new_n538 = ~n290 & new_n517;
  assign new_n539 = ~new_n537 & ~new_n538;
  assign new_n540 = n266 & ~new_n539;
  assign new_n541 = n74 & ~n266;
  assign new_n542_1 = ~new_n540 & ~new_n541;
  assign new_n543 = new_n536 & new_n542_1;
  assign new_n544 = ~new_n536 & ~new_n542_1;
  assign n123 = new_n543 | new_n544;
  assign new_n546 = ~new_n180 & ~new_n345;
  assign new_n547_1 = ~n266 & new_n414;
  assign new_n548 = n266 & new_n344;
  assign new_n549 = ~new_n547_1 & ~new_n548;
  assign new_n550 = ~new_n546 & new_n549;
  assign new_n551 = new_n546 & ~new_n549;
  assign n148 = new_n550 | new_n551;
  assign new_n553 = ~new_n388_1 & ~new_n426;
  assign new_n554 = new_n394_1 & new_n553;
  assign new_n555 = ~new_n394_1 & ~new_n553;
  assign n163 = new_n554 | new_n555;
  assign new_n557_1 = ~new_n481_1 & ~new_n529;
  assign new_n558 = new_n487 & new_n557_1;
  assign new_n559 = ~new_n487 & ~new_n557_1;
  assign n191 = new_n558 | new_n559;
  assign new_n561_1 = ~new_n402 & ~new_n403;
  assign new_n562 = ~n266 & ~n673;
  assign new_n563 = ~new_n328 & ~new_n562;
  assign new_n564 = new_n324 & new_n563;
  assign new_n565 = ~new_n561_1 & new_n564;
  assign new_n566 = new_n561_1 & ~new_n564;
  assign n196 = new_n565 | new_n566;
  assign new_n568_1 = ~new_n407 & ~new_n409_1;
  assign new_n569_1 = ~n266 & ~new_n406;
  assign new_n570 = n266 & ~new_n340;
  assign new_n571_1 = ~new_n569_1 & ~new_n570;
  assign new_n572 = new_n568_1 & new_n571_1;
  assign new_n573 = ~new_n568_1 & ~new_n571_1;
  assign n226 = ~new_n572 & ~new_n573;
  assign new_n575_1 = ~new_n474 & ~new_n528;
  assign new_n576 = new_n480 & new_n575_1;
  assign new_n577 = ~new_n480 & ~new_n575_1;
  assign n240 = new_n576 | new_n577;
  assign new_n579 = ~new_n509 & ~new_n533;
  assign new_n580 = new_n515 & new_n579;
  assign new_n581_1 = ~new_n515 & ~new_n579;
  assign n254 = new_n580 | new_n581_1;
  assign new_n583_1 = ~new_n367 & ~new_n423;
  assign new_n584 = new_n373 & new_n583_1;
  assign new_n585 = ~new_n373 & ~new_n583_1;
  assign n260 = new_n584 | new_n585;
  assign new_n587_1 = ~new_n446 & ~new_n524;
  assign new_n588 = new_n452 & new_n587_1;
  assign new_n589 = ~new_n452 & ~new_n587_1;
  assign n283 = new_n588 | new_n589;
  assign new_n591 = ~new_n374 & ~new_n424;
  assign new_n592 = new_n380 & new_n591;
  assign new_n593 = ~new_n380 & ~new_n591;
  assign n291 = new_n592 | new_n593;
  assign new_n595 = ~new_n396 & ~new_n397;
  assign new_n596 = ~n266 & ~new_n418;
  assign new_n597 = n266 & new_n349_1;
  assign new_n598 = ~new_n596 & ~new_n597;
  assign new_n599 = new_n595 & new_n598;
  assign new_n600_1 = ~new_n595 & ~new_n598;
  assign n299 = new_n599 | new_n600_1;
  assign new_n602 = ~new_n453 & ~new_n525_1;
  assign new_n603_1 = new_n459 & new_n602;
  assign new_n604 = ~new_n459 & ~new_n602;
  assign n442 = new_n603_1 | new_n604;
  assign new_n606 = ~new_n324 & ~new_n330;
  assign n449 = new_n331 | new_n606;
  assign new_n608 = ~new_n502 & ~new_n532;
  assign new_n609_1 = new_n508 & new_n608;
  assign new_n610 = ~new_n508 & ~new_n608;
  assign n484 = new_n609_1 | new_n610;
  assign new_n612 = ~new_n516 & ~new_n534_1;
  assign new_n613_1 = new_n522 & ~new_n612;
  assign new_n614_1 = ~new_n522 & new_n612;
  assign n518 = ~new_n613_1 & ~new_n614_1;
  assign new_n616_1 = ~new_n360_1 & ~new_n366;
  assign new_n617 = ~new_n422 & ~new_n616_1;
  assign new_n618 = ~new_n367 & new_n617;
  assign n534 = ~new_n423 & ~new_n618;
  assign new_n620 = ~new_n488 & ~new_n530;
  assign new_n621 = new_n494_1 & new_n620;
  assign new_n622 = ~new_n494_1 & ~new_n620;
  assign n542 = new_n621 | new_n622;
  assign new_n624 = ~new_n161 & ~new_n162;
  assign new_n625 = ~n266 & ~new_n416;
  assign new_n626 = n266 & new_n347;
  assign new_n627_1 = ~new_n625 & ~new_n626;
  assign new_n628 = ~new_n624 & new_n627_1;
  assign new_n629 = new_n624 & ~new_n627_1;
  assign n547 = new_n628 | new_n629;
  assign new_n631 = ~new_n411 & ~new_n413;
  assign new_n632 = ~n266 & ~new_n410;
  assign new_n633 = n266 & new_n342;
  assign new_n634 = ~new_n632 & ~new_n633;
  assign new_n635_1 = new_n631 & new_n634;
  assign new_n636 = ~new_n631 & ~new_n634;
  assign n568 = ~new_n635_1 & ~new_n636;
  assign new_n638 = ~new_n467 & ~new_n527;
  assign new_n639 = new_n473 & new_n638;
  assign new_n640 = ~new_n473 & ~new_n638;
  assign n627 = new_n639 | new_n640;
  assign new_n642 = ~new_n495 & ~new_n531;
  assign new_n643 = new_n501 & new_n642;
  assign new_n644 = ~new_n501 & ~new_n642;
  assign n635 = new_n643 | new_n644;
  assign new_n646_1 = ~new_n460 & ~new_n526;
  assign new_n647 = new_n466 & new_n646_1;
  assign new_n648 = ~new_n466 & ~new_n646_1;
  assign n672 = new_n647 | new_n648;
endmodule


